module top(in1, in2, in3, in4, in5, out1, out2, out3);
  input [15:0] in1, in2, in3, in4, in5;
  output [16:0] out1, out2;
  output [33:0] out3;
  wire [15:0] in1, in2, in3, in4, in5;
  wire [16:0] out1, out2;
  wire [33:0] out3;
  wire add_10_21_n_1, add_10_21_n_2, add_10_21_n_3, add_10_21_n_4, add_10_21_n_5, add_10_21_n_6, add_10_21_n_7, add_10_21_n_8;
  wire add_10_21_n_9, add_10_21_n_10, add_10_21_n_11, add_10_21_n_12, add_10_21_n_13, add_10_21_n_14, add_10_21_n_15, add_10_21_n_16;
  wire add_10_21_n_17, add_10_21_n_18, add_10_21_n_19, add_10_21_n_20, add_10_21_n_21, add_10_21_n_22, add_10_21_n_23, add_10_21_n_24;
  wire add_10_21_n_25, add_10_21_n_26, add_10_21_n_27, add_10_21_n_28, add_10_21_n_29, add_10_21_n_30, add_10_21_n_31, add_10_21_n_32;
  wire add_10_21_n_33, add_10_21_n_34, add_10_21_n_35, add_10_21_n_36, add_10_21_n_37, add_10_21_n_38, add_10_21_n_39, add_10_21_n_40;
  wire add_10_21_n_41, add_10_21_n_42, add_10_21_n_43, add_10_21_n_44, add_10_21_n_45, add_10_21_n_46, add_10_21_n_47, add_10_21_n_48;
  wire add_10_21_n_49, add_10_21_n_50, add_10_21_n_51, add_10_21_n_52, add_10_21_n_54, add_10_21_n_56, add_10_21_n_57, add_10_21_n_59;
  wire add_10_21_n_60, add_10_21_n_62, add_10_21_n_63, add_10_21_n_65, add_10_21_n_66, add_10_21_n_68, add_10_21_n_69, add_10_21_n_71;
  wire add_10_21_n_72, add_10_21_n_74, add_10_21_n_75, add_10_21_n_77, add_10_21_n_78, add_10_21_n_80, add_10_21_n_81, add_10_21_n_83;
  wire add_10_21_n_84, add_10_21_n_86, add_10_21_n_87, add_10_21_n_89, add_10_21_n_90, add_10_21_n_92, add_10_21_n_93, csa_tree_add_12_51_groupi_n_0;
  wire csa_tree_add_12_51_groupi_n_1, csa_tree_add_12_51_groupi_n_2, csa_tree_add_12_51_groupi_n_3, csa_tree_add_12_51_groupi_n_4, csa_tree_add_12_51_groupi_n_5, csa_tree_add_12_51_groupi_n_6, csa_tree_add_12_51_groupi_n_7, csa_tree_add_12_51_groupi_n_8;
  wire csa_tree_add_12_51_groupi_n_9, csa_tree_add_12_51_groupi_n_10, csa_tree_add_12_51_groupi_n_11, csa_tree_add_12_51_groupi_n_12, csa_tree_add_12_51_groupi_n_13, csa_tree_add_12_51_groupi_n_14, csa_tree_add_12_51_groupi_n_15, csa_tree_add_12_51_groupi_n_16;
  wire csa_tree_add_12_51_groupi_n_17, csa_tree_add_12_51_groupi_n_18, csa_tree_add_12_51_groupi_n_19, csa_tree_add_12_51_groupi_n_20, csa_tree_add_12_51_groupi_n_21, csa_tree_add_12_51_groupi_n_22, csa_tree_add_12_51_groupi_n_23, csa_tree_add_12_51_groupi_n_24;
  wire csa_tree_add_12_51_groupi_n_25, csa_tree_add_12_51_groupi_n_26, csa_tree_add_12_51_groupi_n_27, csa_tree_add_12_51_groupi_n_28, csa_tree_add_12_51_groupi_n_29, csa_tree_add_12_51_groupi_n_30, csa_tree_add_12_51_groupi_n_31, csa_tree_add_12_51_groupi_n_32;
  wire csa_tree_add_12_51_groupi_n_33, csa_tree_add_12_51_groupi_n_34, csa_tree_add_12_51_groupi_n_35, csa_tree_add_12_51_groupi_n_36, csa_tree_add_12_51_groupi_n_37, csa_tree_add_12_51_groupi_n_38, csa_tree_add_12_51_groupi_n_39, csa_tree_add_12_51_groupi_n_40;
  wire csa_tree_add_12_51_groupi_n_41, csa_tree_add_12_51_groupi_n_42, csa_tree_add_12_51_groupi_n_43, csa_tree_add_12_51_groupi_n_44, csa_tree_add_12_51_groupi_n_45, csa_tree_add_12_51_groupi_n_46, csa_tree_add_12_51_groupi_n_47, csa_tree_add_12_51_groupi_n_48;
  wire csa_tree_add_12_51_groupi_n_49, csa_tree_add_12_51_groupi_n_50, csa_tree_add_12_51_groupi_n_51, csa_tree_add_12_51_groupi_n_52, csa_tree_add_12_51_groupi_n_53, csa_tree_add_12_51_groupi_n_54, csa_tree_add_12_51_groupi_n_55, csa_tree_add_12_51_groupi_n_56;
  wire csa_tree_add_12_51_groupi_n_57, csa_tree_add_12_51_groupi_n_58, csa_tree_add_12_51_groupi_n_59, csa_tree_add_12_51_groupi_n_60, csa_tree_add_12_51_groupi_n_61, csa_tree_add_12_51_groupi_n_62, csa_tree_add_12_51_groupi_n_63, csa_tree_add_12_51_groupi_n_64;
  wire csa_tree_add_12_51_groupi_n_65, csa_tree_add_12_51_groupi_n_66, csa_tree_add_12_51_groupi_n_67, csa_tree_add_12_51_groupi_n_68, csa_tree_add_12_51_groupi_n_69, csa_tree_add_12_51_groupi_n_70, csa_tree_add_12_51_groupi_n_71, csa_tree_add_12_51_groupi_n_72;
  wire csa_tree_add_12_51_groupi_n_73, csa_tree_add_12_51_groupi_n_74, csa_tree_add_12_51_groupi_n_75, csa_tree_add_12_51_groupi_n_76, csa_tree_add_12_51_groupi_n_77, csa_tree_add_12_51_groupi_n_78, csa_tree_add_12_51_groupi_n_79, csa_tree_add_12_51_groupi_n_80;
  wire csa_tree_add_12_51_groupi_n_81, csa_tree_add_12_51_groupi_n_82, csa_tree_add_12_51_groupi_n_83, csa_tree_add_12_51_groupi_n_84, csa_tree_add_12_51_groupi_n_85, csa_tree_add_12_51_groupi_n_86, csa_tree_add_12_51_groupi_n_87, csa_tree_add_12_51_groupi_n_88;
  wire csa_tree_add_12_51_groupi_n_89, csa_tree_add_12_51_groupi_n_90, csa_tree_add_12_51_groupi_n_91, csa_tree_add_12_51_groupi_n_92, csa_tree_add_12_51_groupi_n_93, csa_tree_add_12_51_groupi_n_94, csa_tree_add_12_51_groupi_n_95, csa_tree_add_12_51_groupi_n_96;
  wire csa_tree_add_12_51_groupi_n_97, csa_tree_add_12_51_groupi_n_98, csa_tree_add_12_51_groupi_n_99, csa_tree_add_12_51_groupi_n_100, csa_tree_add_12_51_groupi_n_101, csa_tree_add_12_51_groupi_n_102, csa_tree_add_12_51_groupi_n_103, csa_tree_add_12_51_groupi_n_104;
  wire csa_tree_add_12_51_groupi_n_105, csa_tree_add_12_51_groupi_n_106, csa_tree_add_12_51_groupi_n_107, csa_tree_add_12_51_groupi_n_108, csa_tree_add_12_51_groupi_n_109, csa_tree_add_12_51_groupi_n_110, csa_tree_add_12_51_groupi_n_111, csa_tree_add_12_51_groupi_n_112;
  wire csa_tree_add_12_51_groupi_n_113, csa_tree_add_12_51_groupi_n_114, csa_tree_add_12_51_groupi_n_115, csa_tree_add_12_51_groupi_n_116, csa_tree_add_12_51_groupi_n_117, csa_tree_add_12_51_groupi_n_118, csa_tree_add_12_51_groupi_n_119, csa_tree_add_12_51_groupi_n_120;
  wire csa_tree_add_12_51_groupi_n_121, csa_tree_add_12_51_groupi_n_122, csa_tree_add_12_51_groupi_n_123, csa_tree_add_12_51_groupi_n_124, csa_tree_add_12_51_groupi_n_125, csa_tree_add_12_51_groupi_n_126, csa_tree_add_12_51_groupi_n_127, csa_tree_add_12_51_groupi_n_128;
  wire csa_tree_add_12_51_groupi_n_129, csa_tree_add_12_51_groupi_n_130, csa_tree_add_12_51_groupi_n_131, csa_tree_add_12_51_groupi_n_132, csa_tree_add_12_51_groupi_n_133, csa_tree_add_12_51_groupi_n_134, csa_tree_add_12_51_groupi_n_135, csa_tree_add_12_51_groupi_n_136;
  wire csa_tree_add_12_51_groupi_n_137, csa_tree_add_12_51_groupi_n_138, csa_tree_add_12_51_groupi_n_139, csa_tree_add_12_51_groupi_n_140, csa_tree_add_12_51_groupi_n_141, csa_tree_add_12_51_groupi_n_142, csa_tree_add_12_51_groupi_n_143, csa_tree_add_12_51_groupi_n_144;
  wire csa_tree_add_12_51_groupi_n_145, csa_tree_add_12_51_groupi_n_146, csa_tree_add_12_51_groupi_n_147, csa_tree_add_12_51_groupi_n_148, csa_tree_add_12_51_groupi_n_149, csa_tree_add_12_51_groupi_n_150, csa_tree_add_12_51_groupi_n_151, csa_tree_add_12_51_groupi_n_152;
  wire csa_tree_add_12_51_groupi_n_153, csa_tree_add_12_51_groupi_n_154, csa_tree_add_12_51_groupi_n_155, csa_tree_add_12_51_groupi_n_156, csa_tree_add_12_51_groupi_n_157, csa_tree_add_12_51_groupi_n_158, csa_tree_add_12_51_groupi_n_159, csa_tree_add_12_51_groupi_n_160;
  wire csa_tree_add_12_51_groupi_n_161, csa_tree_add_12_51_groupi_n_162, csa_tree_add_12_51_groupi_n_163, csa_tree_add_12_51_groupi_n_164, csa_tree_add_12_51_groupi_n_165, csa_tree_add_12_51_groupi_n_166, csa_tree_add_12_51_groupi_n_167, csa_tree_add_12_51_groupi_n_168;
  wire csa_tree_add_12_51_groupi_n_169, csa_tree_add_12_51_groupi_n_170, csa_tree_add_12_51_groupi_n_171, csa_tree_add_12_51_groupi_n_172, csa_tree_add_12_51_groupi_n_173, csa_tree_add_12_51_groupi_n_174, csa_tree_add_12_51_groupi_n_175, csa_tree_add_12_51_groupi_n_176;
  wire csa_tree_add_12_51_groupi_n_177, csa_tree_add_12_51_groupi_n_178, csa_tree_add_12_51_groupi_n_179, csa_tree_add_12_51_groupi_n_180, csa_tree_add_12_51_groupi_n_181, csa_tree_add_12_51_groupi_n_182, csa_tree_add_12_51_groupi_n_183, csa_tree_add_12_51_groupi_n_184;
  wire csa_tree_add_12_51_groupi_n_185, csa_tree_add_12_51_groupi_n_186, csa_tree_add_12_51_groupi_n_187, csa_tree_add_12_51_groupi_n_188, csa_tree_add_12_51_groupi_n_189, csa_tree_add_12_51_groupi_n_190, csa_tree_add_12_51_groupi_n_191, csa_tree_add_12_51_groupi_n_192;
  wire csa_tree_add_12_51_groupi_n_193, csa_tree_add_12_51_groupi_n_194, csa_tree_add_12_51_groupi_n_195, csa_tree_add_12_51_groupi_n_196, csa_tree_add_12_51_groupi_n_197, csa_tree_add_12_51_groupi_n_198, csa_tree_add_12_51_groupi_n_199, csa_tree_add_12_51_groupi_n_200;
  wire csa_tree_add_12_51_groupi_n_201, csa_tree_add_12_51_groupi_n_202, csa_tree_add_12_51_groupi_n_203, csa_tree_add_12_51_groupi_n_204, csa_tree_add_12_51_groupi_n_205, csa_tree_add_12_51_groupi_n_206, csa_tree_add_12_51_groupi_n_207, csa_tree_add_12_51_groupi_n_208;
  wire csa_tree_add_12_51_groupi_n_209, csa_tree_add_12_51_groupi_n_210, csa_tree_add_12_51_groupi_n_211, csa_tree_add_12_51_groupi_n_212, csa_tree_add_12_51_groupi_n_213, csa_tree_add_12_51_groupi_n_214, csa_tree_add_12_51_groupi_n_215, csa_tree_add_12_51_groupi_n_216;
  wire csa_tree_add_12_51_groupi_n_217, csa_tree_add_12_51_groupi_n_218, csa_tree_add_12_51_groupi_n_219, csa_tree_add_12_51_groupi_n_220, csa_tree_add_12_51_groupi_n_221, csa_tree_add_12_51_groupi_n_222, csa_tree_add_12_51_groupi_n_223, csa_tree_add_12_51_groupi_n_224;
  wire csa_tree_add_12_51_groupi_n_225, csa_tree_add_12_51_groupi_n_226, csa_tree_add_12_51_groupi_n_227, csa_tree_add_12_51_groupi_n_228, csa_tree_add_12_51_groupi_n_229, csa_tree_add_12_51_groupi_n_230, csa_tree_add_12_51_groupi_n_231, csa_tree_add_12_51_groupi_n_232;
  wire csa_tree_add_12_51_groupi_n_233, csa_tree_add_12_51_groupi_n_234, csa_tree_add_12_51_groupi_n_235, csa_tree_add_12_51_groupi_n_236, csa_tree_add_12_51_groupi_n_237, csa_tree_add_12_51_groupi_n_238, csa_tree_add_12_51_groupi_n_239, csa_tree_add_12_51_groupi_n_240;
  wire csa_tree_add_12_51_groupi_n_241, csa_tree_add_12_51_groupi_n_242, csa_tree_add_12_51_groupi_n_243, csa_tree_add_12_51_groupi_n_244, csa_tree_add_12_51_groupi_n_245, csa_tree_add_12_51_groupi_n_246, csa_tree_add_12_51_groupi_n_247, csa_tree_add_12_51_groupi_n_248;
  wire csa_tree_add_12_51_groupi_n_249, csa_tree_add_12_51_groupi_n_250, csa_tree_add_12_51_groupi_n_251, csa_tree_add_12_51_groupi_n_252, csa_tree_add_12_51_groupi_n_253, csa_tree_add_12_51_groupi_n_254, csa_tree_add_12_51_groupi_n_255, csa_tree_add_12_51_groupi_n_256;
  wire csa_tree_add_12_51_groupi_n_257, csa_tree_add_12_51_groupi_n_258, csa_tree_add_12_51_groupi_n_259, csa_tree_add_12_51_groupi_n_260, csa_tree_add_12_51_groupi_n_261, csa_tree_add_12_51_groupi_n_262, csa_tree_add_12_51_groupi_n_263, csa_tree_add_12_51_groupi_n_264;
  wire csa_tree_add_12_51_groupi_n_265, csa_tree_add_12_51_groupi_n_266, csa_tree_add_12_51_groupi_n_267, csa_tree_add_12_51_groupi_n_268, csa_tree_add_12_51_groupi_n_269, csa_tree_add_12_51_groupi_n_270, csa_tree_add_12_51_groupi_n_271, csa_tree_add_12_51_groupi_n_272;
  wire csa_tree_add_12_51_groupi_n_273, csa_tree_add_12_51_groupi_n_274, csa_tree_add_12_51_groupi_n_275, csa_tree_add_12_51_groupi_n_276, csa_tree_add_12_51_groupi_n_277, csa_tree_add_12_51_groupi_n_278, csa_tree_add_12_51_groupi_n_279, csa_tree_add_12_51_groupi_n_280;
  wire csa_tree_add_12_51_groupi_n_281, csa_tree_add_12_51_groupi_n_282, csa_tree_add_12_51_groupi_n_283, csa_tree_add_12_51_groupi_n_284, csa_tree_add_12_51_groupi_n_285, csa_tree_add_12_51_groupi_n_286, csa_tree_add_12_51_groupi_n_287, csa_tree_add_12_51_groupi_n_288;
  wire csa_tree_add_12_51_groupi_n_289, csa_tree_add_12_51_groupi_n_290, csa_tree_add_12_51_groupi_n_291, csa_tree_add_12_51_groupi_n_292, csa_tree_add_12_51_groupi_n_293, csa_tree_add_12_51_groupi_n_294, csa_tree_add_12_51_groupi_n_295, csa_tree_add_12_51_groupi_n_296;
  wire csa_tree_add_12_51_groupi_n_297, csa_tree_add_12_51_groupi_n_298, csa_tree_add_12_51_groupi_n_299, csa_tree_add_12_51_groupi_n_300, csa_tree_add_12_51_groupi_n_301, csa_tree_add_12_51_groupi_n_302, csa_tree_add_12_51_groupi_n_303, csa_tree_add_12_51_groupi_n_304;
  wire csa_tree_add_12_51_groupi_n_305, csa_tree_add_12_51_groupi_n_306, csa_tree_add_12_51_groupi_n_307, csa_tree_add_12_51_groupi_n_308, csa_tree_add_12_51_groupi_n_309, csa_tree_add_12_51_groupi_n_310, csa_tree_add_12_51_groupi_n_311, csa_tree_add_12_51_groupi_n_312;
  wire csa_tree_add_12_51_groupi_n_313, csa_tree_add_12_51_groupi_n_314, csa_tree_add_12_51_groupi_n_315, csa_tree_add_12_51_groupi_n_316, csa_tree_add_12_51_groupi_n_317, csa_tree_add_12_51_groupi_n_318, csa_tree_add_12_51_groupi_n_319, csa_tree_add_12_51_groupi_n_320;
  wire csa_tree_add_12_51_groupi_n_321, csa_tree_add_12_51_groupi_n_322, csa_tree_add_12_51_groupi_n_323, csa_tree_add_12_51_groupi_n_324, csa_tree_add_12_51_groupi_n_325, csa_tree_add_12_51_groupi_n_326, csa_tree_add_12_51_groupi_n_327, csa_tree_add_12_51_groupi_n_328;
  wire csa_tree_add_12_51_groupi_n_329, csa_tree_add_12_51_groupi_n_330, csa_tree_add_12_51_groupi_n_331, csa_tree_add_12_51_groupi_n_332, csa_tree_add_12_51_groupi_n_333, csa_tree_add_12_51_groupi_n_334, csa_tree_add_12_51_groupi_n_335, csa_tree_add_12_51_groupi_n_336;
  wire csa_tree_add_12_51_groupi_n_337, csa_tree_add_12_51_groupi_n_338, csa_tree_add_12_51_groupi_n_339, csa_tree_add_12_51_groupi_n_340, csa_tree_add_12_51_groupi_n_341, csa_tree_add_12_51_groupi_n_342, csa_tree_add_12_51_groupi_n_343, csa_tree_add_12_51_groupi_n_344;
  wire csa_tree_add_12_51_groupi_n_345, csa_tree_add_12_51_groupi_n_346, csa_tree_add_12_51_groupi_n_347, csa_tree_add_12_51_groupi_n_348, csa_tree_add_12_51_groupi_n_349, csa_tree_add_12_51_groupi_n_350, csa_tree_add_12_51_groupi_n_351, csa_tree_add_12_51_groupi_n_352;
  wire csa_tree_add_12_51_groupi_n_353, csa_tree_add_12_51_groupi_n_354, csa_tree_add_12_51_groupi_n_355, csa_tree_add_12_51_groupi_n_356, csa_tree_add_12_51_groupi_n_357, csa_tree_add_12_51_groupi_n_358, csa_tree_add_12_51_groupi_n_359, csa_tree_add_12_51_groupi_n_360;
  wire csa_tree_add_12_51_groupi_n_361, csa_tree_add_12_51_groupi_n_362, csa_tree_add_12_51_groupi_n_363, csa_tree_add_12_51_groupi_n_364, csa_tree_add_12_51_groupi_n_365, csa_tree_add_12_51_groupi_n_366, csa_tree_add_12_51_groupi_n_367, csa_tree_add_12_51_groupi_n_368;
  wire csa_tree_add_12_51_groupi_n_369, csa_tree_add_12_51_groupi_n_370, csa_tree_add_12_51_groupi_n_371, csa_tree_add_12_51_groupi_n_372, csa_tree_add_12_51_groupi_n_373, csa_tree_add_12_51_groupi_n_374, csa_tree_add_12_51_groupi_n_375, csa_tree_add_12_51_groupi_n_376;
  wire csa_tree_add_12_51_groupi_n_377, csa_tree_add_12_51_groupi_n_378, csa_tree_add_12_51_groupi_n_379, csa_tree_add_12_51_groupi_n_380, csa_tree_add_12_51_groupi_n_381, csa_tree_add_12_51_groupi_n_382, csa_tree_add_12_51_groupi_n_383, csa_tree_add_12_51_groupi_n_384;
  wire csa_tree_add_12_51_groupi_n_385, csa_tree_add_12_51_groupi_n_386, csa_tree_add_12_51_groupi_n_387, csa_tree_add_12_51_groupi_n_388, csa_tree_add_12_51_groupi_n_389, csa_tree_add_12_51_groupi_n_390, csa_tree_add_12_51_groupi_n_391, csa_tree_add_12_51_groupi_n_392;
  wire csa_tree_add_12_51_groupi_n_393, csa_tree_add_12_51_groupi_n_394, csa_tree_add_12_51_groupi_n_395, csa_tree_add_12_51_groupi_n_396, csa_tree_add_12_51_groupi_n_397, csa_tree_add_12_51_groupi_n_398, csa_tree_add_12_51_groupi_n_399, csa_tree_add_12_51_groupi_n_400;
  wire csa_tree_add_12_51_groupi_n_401, csa_tree_add_12_51_groupi_n_402, csa_tree_add_12_51_groupi_n_403, csa_tree_add_12_51_groupi_n_404, csa_tree_add_12_51_groupi_n_405, csa_tree_add_12_51_groupi_n_406, csa_tree_add_12_51_groupi_n_407, csa_tree_add_12_51_groupi_n_408;
  wire csa_tree_add_12_51_groupi_n_409, csa_tree_add_12_51_groupi_n_410, csa_tree_add_12_51_groupi_n_411, csa_tree_add_12_51_groupi_n_412, csa_tree_add_12_51_groupi_n_413, csa_tree_add_12_51_groupi_n_414, csa_tree_add_12_51_groupi_n_415, csa_tree_add_12_51_groupi_n_416;
  wire csa_tree_add_12_51_groupi_n_417, csa_tree_add_12_51_groupi_n_418, csa_tree_add_12_51_groupi_n_419, csa_tree_add_12_51_groupi_n_420, csa_tree_add_12_51_groupi_n_421, csa_tree_add_12_51_groupi_n_422, csa_tree_add_12_51_groupi_n_423, csa_tree_add_12_51_groupi_n_424;
  wire csa_tree_add_12_51_groupi_n_425, csa_tree_add_12_51_groupi_n_426, csa_tree_add_12_51_groupi_n_427, csa_tree_add_12_51_groupi_n_428, csa_tree_add_12_51_groupi_n_429, csa_tree_add_12_51_groupi_n_430, csa_tree_add_12_51_groupi_n_431, csa_tree_add_12_51_groupi_n_432;
  wire csa_tree_add_12_51_groupi_n_433, csa_tree_add_12_51_groupi_n_434, csa_tree_add_12_51_groupi_n_435, csa_tree_add_12_51_groupi_n_436, csa_tree_add_12_51_groupi_n_437, csa_tree_add_12_51_groupi_n_438, csa_tree_add_12_51_groupi_n_439, csa_tree_add_12_51_groupi_n_440;
  wire csa_tree_add_12_51_groupi_n_441, csa_tree_add_12_51_groupi_n_442, csa_tree_add_12_51_groupi_n_443, csa_tree_add_12_51_groupi_n_444, csa_tree_add_12_51_groupi_n_445, csa_tree_add_12_51_groupi_n_446, csa_tree_add_12_51_groupi_n_447, csa_tree_add_12_51_groupi_n_448;
  wire csa_tree_add_12_51_groupi_n_449, csa_tree_add_12_51_groupi_n_450, csa_tree_add_12_51_groupi_n_451, csa_tree_add_12_51_groupi_n_452, csa_tree_add_12_51_groupi_n_453, csa_tree_add_12_51_groupi_n_454, csa_tree_add_12_51_groupi_n_455, csa_tree_add_12_51_groupi_n_456;
  wire csa_tree_add_12_51_groupi_n_457, csa_tree_add_12_51_groupi_n_458, csa_tree_add_12_51_groupi_n_459, csa_tree_add_12_51_groupi_n_460, csa_tree_add_12_51_groupi_n_461, csa_tree_add_12_51_groupi_n_462, csa_tree_add_12_51_groupi_n_463, csa_tree_add_12_51_groupi_n_464;
  wire csa_tree_add_12_51_groupi_n_465, csa_tree_add_12_51_groupi_n_466, csa_tree_add_12_51_groupi_n_467, csa_tree_add_12_51_groupi_n_468, csa_tree_add_12_51_groupi_n_469, csa_tree_add_12_51_groupi_n_470, csa_tree_add_12_51_groupi_n_471, csa_tree_add_12_51_groupi_n_472;
  wire csa_tree_add_12_51_groupi_n_473, csa_tree_add_12_51_groupi_n_474, csa_tree_add_12_51_groupi_n_475, csa_tree_add_12_51_groupi_n_476, csa_tree_add_12_51_groupi_n_477, csa_tree_add_12_51_groupi_n_478, csa_tree_add_12_51_groupi_n_479, csa_tree_add_12_51_groupi_n_480;
  wire csa_tree_add_12_51_groupi_n_481, csa_tree_add_12_51_groupi_n_482, csa_tree_add_12_51_groupi_n_483, csa_tree_add_12_51_groupi_n_484, csa_tree_add_12_51_groupi_n_485, csa_tree_add_12_51_groupi_n_486, csa_tree_add_12_51_groupi_n_487, csa_tree_add_12_51_groupi_n_488;
  wire csa_tree_add_12_51_groupi_n_489, csa_tree_add_12_51_groupi_n_490, csa_tree_add_12_51_groupi_n_491, csa_tree_add_12_51_groupi_n_492, csa_tree_add_12_51_groupi_n_493, csa_tree_add_12_51_groupi_n_494, csa_tree_add_12_51_groupi_n_495, csa_tree_add_12_51_groupi_n_496;
  wire csa_tree_add_12_51_groupi_n_497, csa_tree_add_12_51_groupi_n_498, csa_tree_add_12_51_groupi_n_499, csa_tree_add_12_51_groupi_n_500, csa_tree_add_12_51_groupi_n_501, csa_tree_add_12_51_groupi_n_502, csa_tree_add_12_51_groupi_n_503, csa_tree_add_12_51_groupi_n_504;
  wire csa_tree_add_12_51_groupi_n_505, csa_tree_add_12_51_groupi_n_506, csa_tree_add_12_51_groupi_n_507, csa_tree_add_12_51_groupi_n_508, csa_tree_add_12_51_groupi_n_509, csa_tree_add_12_51_groupi_n_510, csa_tree_add_12_51_groupi_n_511, csa_tree_add_12_51_groupi_n_512;
  wire csa_tree_add_12_51_groupi_n_513, csa_tree_add_12_51_groupi_n_514, csa_tree_add_12_51_groupi_n_515, csa_tree_add_12_51_groupi_n_516, csa_tree_add_12_51_groupi_n_517, csa_tree_add_12_51_groupi_n_518, csa_tree_add_12_51_groupi_n_519, csa_tree_add_12_51_groupi_n_520;
  wire csa_tree_add_12_51_groupi_n_521, csa_tree_add_12_51_groupi_n_522, csa_tree_add_12_51_groupi_n_523, csa_tree_add_12_51_groupi_n_524, csa_tree_add_12_51_groupi_n_525, csa_tree_add_12_51_groupi_n_526, csa_tree_add_12_51_groupi_n_527, csa_tree_add_12_51_groupi_n_528;
  wire csa_tree_add_12_51_groupi_n_529, csa_tree_add_12_51_groupi_n_530, csa_tree_add_12_51_groupi_n_531, csa_tree_add_12_51_groupi_n_532, csa_tree_add_12_51_groupi_n_533, csa_tree_add_12_51_groupi_n_534, csa_tree_add_12_51_groupi_n_535, csa_tree_add_12_51_groupi_n_536;
  wire csa_tree_add_12_51_groupi_n_537, csa_tree_add_12_51_groupi_n_538, csa_tree_add_12_51_groupi_n_539, csa_tree_add_12_51_groupi_n_540, csa_tree_add_12_51_groupi_n_541, csa_tree_add_12_51_groupi_n_542, csa_tree_add_12_51_groupi_n_543, csa_tree_add_12_51_groupi_n_544;
  wire csa_tree_add_12_51_groupi_n_545, csa_tree_add_12_51_groupi_n_546, csa_tree_add_12_51_groupi_n_547, csa_tree_add_12_51_groupi_n_548, csa_tree_add_12_51_groupi_n_549, csa_tree_add_12_51_groupi_n_550, csa_tree_add_12_51_groupi_n_551, csa_tree_add_12_51_groupi_n_552;
  wire csa_tree_add_12_51_groupi_n_553, csa_tree_add_12_51_groupi_n_554, csa_tree_add_12_51_groupi_n_555, csa_tree_add_12_51_groupi_n_556, csa_tree_add_12_51_groupi_n_557, csa_tree_add_12_51_groupi_n_558, csa_tree_add_12_51_groupi_n_559, csa_tree_add_12_51_groupi_n_560;
  wire csa_tree_add_12_51_groupi_n_561, csa_tree_add_12_51_groupi_n_562, csa_tree_add_12_51_groupi_n_563, csa_tree_add_12_51_groupi_n_564, csa_tree_add_12_51_groupi_n_565, csa_tree_add_12_51_groupi_n_566, csa_tree_add_12_51_groupi_n_567, csa_tree_add_12_51_groupi_n_568;
  wire csa_tree_add_12_51_groupi_n_569, csa_tree_add_12_51_groupi_n_570, csa_tree_add_12_51_groupi_n_571, csa_tree_add_12_51_groupi_n_572, csa_tree_add_12_51_groupi_n_573, csa_tree_add_12_51_groupi_n_574, csa_tree_add_12_51_groupi_n_575, csa_tree_add_12_51_groupi_n_576;
  wire csa_tree_add_12_51_groupi_n_577, csa_tree_add_12_51_groupi_n_578, csa_tree_add_12_51_groupi_n_579, csa_tree_add_12_51_groupi_n_580, csa_tree_add_12_51_groupi_n_581, csa_tree_add_12_51_groupi_n_582, csa_tree_add_12_51_groupi_n_583, csa_tree_add_12_51_groupi_n_584;
  wire csa_tree_add_12_51_groupi_n_585, csa_tree_add_12_51_groupi_n_586, csa_tree_add_12_51_groupi_n_587, csa_tree_add_12_51_groupi_n_588, csa_tree_add_12_51_groupi_n_589, csa_tree_add_12_51_groupi_n_590, csa_tree_add_12_51_groupi_n_591, csa_tree_add_12_51_groupi_n_592;
  wire csa_tree_add_12_51_groupi_n_593, csa_tree_add_12_51_groupi_n_594, csa_tree_add_12_51_groupi_n_595, csa_tree_add_12_51_groupi_n_596, csa_tree_add_12_51_groupi_n_597, csa_tree_add_12_51_groupi_n_598, csa_tree_add_12_51_groupi_n_599, csa_tree_add_12_51_groupi_n_600;
  wire csa_tree_add_12_51_groupi_n_601, csa_tree_add_12_51_groupi_n_602, csa_tree_add_12_51_groupi_n_603, csa_tree_add_12_51_groupi_n_604, csa_tree_add_12_51_groupi_n_605, csa_tree_add_12_51_groupi_n_606, csa_tree_add_12_51_groupi_n_607, csa_tree_add_12_51_groupi_n_608;
  wire csa_tree_add_12_51_groupi_n_609, csa_tree_add_12_51_groupi_n_610, csa_tree_add_12_51_groupi_n_611, csa_tree_add_12_51_groupi_n_612, csa_tree_add_12_51_groupi_n_613, csa_tree_add_12_51_groupi_n_614, csa_tree_add_12_51_groupi_n_615, csa_tree_add_12_51_groupi_n_616;
  wire csa_tree_add_12_51_groupi_n_617, csa_tree_add_12_51_groupi_n_618, csa_tree_add_12_51_groupi_n_619, csa_tree_add_12_51_groupi_n_620, csa_tree_add_12_51_groupi_n_621, csa_tree_add_12_51_groupi_n_622, csa_tree_add_12_51_groupi_n_623, csa_tree_add_12_51_groupi_n_624;
  wire csa_tree_add_12_51_groupi_n_625, csa_tree_add_12_51_groupi_n_626, csa_tree_add_12_51_groupi_n_627, csa_tree_add_12_51_groupi_n_628, csa_tree_add_12_51_groupi_n_629, csa_tree_add_12_51_groupi_n_630, csa_tree_add_12_51_groupi_n_631, csa_tree_add_12_51_groupi_n_632;
  wire csa_tree_add_12_51_groupi_n_633, csa_tree_add_12_51_groupi_n_634, csa_tree_add_12_51_groupi_n_635, csa_tree_add_12_51_groupi_n_636, csa_tree_add_12_51_groupi_n_637, csa_tree_add_12_51_groupi_n_638, csa_tree_add_12_51_groupi_n_639, csa_tree_add_12_51_groupi_n_640;
  wire csa_tree_add_12_51_groupi_n_641, csa_tree_add_12_51_groupi_n_642, csa_tree_add_12_51_groupi_n_643, csa_tree_add_12_51_groupi_n_644, csa_tree_add_12_51_groupi_n_645, csa_tree_add_12_51_groupi_n_646, csa_tree_add_12_51_groupi_n_647, csa_tree_add_12_51_groupi_n_648;
  wire csa_tree_add_12_51_groupi_n_649, csa_tree_add_12_51_groupi_n_650, csa_tree_add_12_51_groupi_n_651, csa_tree_add_12_51_groupi_n_652, csa_tree_add_12_51_groupi_n_653, csa_tree_add_12_51_groupi_n_654, csa_tree_add_12_51_groupi_n_655, csa_tree_add_12_51_groupi_n_656;
  wire csa_tree_add_12_51_groupi_n_657, csa_tree_add_12_51_groupi_n_658, csa_tree_add_12_51_groupi_n_659, csa_tree_add_12_51_groupi_n_660, csa_tree_add_12_51_groupi_n_661, csa_tree_add_12_51_groupi_n_662, csa_tree_add_12_51_groupi_n_663, csa_tree_add_12_51_groupi_n_664;
  wire csa_tree_add_12_51_groupi_n_665, csa_tree_add_12_51_groupi_n_666, csa_tree_add_12_51_groupi_n_667, csa_tree_add_12_51_groupi_n_668, csa_tree_add_12_51_groupi_n_669, csa_tree_add_12_51_groupi_n_670, csa_tree_add_12_51_groupi_n_671, csa_tree_add_12_51_groupi_n_672;
  wire csa_tree_add_12_51_groupi_n_673, csa_tree_add_12_51_groupi_n_674, csa_tree_add_12_51_groupi_n_675, csa_tree_add_12_51_groupi_n_676, csa_tree_add_12_51_groupi_n_677, csa_tree_add_12_51_groupi_n_678, csa_tree_add_12_51_groupi_n_679, csa_tree_add_12_51_groupi_n_680;
  wire csa_tree_add_12_51_groupi_n_681, csa_tree_add_12_51_groupi_n_682, csa_tree_add_12_51_groupi_n_683, csa_tree_add_12_51_groupi_n_684, csa_tree_add_12_51_groupi_n_685, csa_tree_add_12_51_groupi_n_686, csa_tree_add_12_51_groupi_n_687, csa_tree_add_12_51_groupi_n_688;
  wire csa_tree_add_12_51_groupi_n_689, csa_tree_add_12_51_groupi_n_690, csa_tree_add_12_51_groupi_n_691, csa_tree_add_12_51_groupi_n_692, csa_tree_add_12_51_groupi_n_693, csa_tree_add_12_51_groupi_n_694, csa_tree_add_12_51_groupi_n_695, csa_tree_add_12_51_groupi_n_696;
  wire csa_tree_add_12_51_groupi_n_697, csa_tree_add_12_51_groupi_n_698, csa_tree_add_12_51_groupi_n_699, csa_tree_add_12_51_groupi_n_700, csa_tree_add_12_51_groupi_n_701, csa_tree_add_12_51_groupi_n_702, csa_tree_add_12_51_groupi_n_703, csa_tree_add_12_51_groupi_n_704;
  wire csa_tree_add_12_51_groupi_n_705, csa_tree_add_12_51_groupi_n_706, csa_tree_add_12_51_groupi_n_707, csa_tree_add_12_51_groupi_n_708, csa_tree_add_12_51_groupi_n_709, csa_tree_add_12_51_groupi_n_710, csa_tree_add_12_51_groupi_n_711, csa_tree_add_12_51_groupi_n_712;
  wire csa_tree_add_12_51_groupi_n_713, csa_tree_add_12_51_groupi_n_714, csa_tree_add_12_51_groupi_n_715, csa_tree_add_12_51_groupi_n_716, csa_tree_add_12_51_groupi_n_717, csa_tree_add_12_51_groupi_n_718, csa_tree_add_12_51_groupi_n_719, csa_tree_add_12_51_groupi_n_720;
  wire csa_tree_add_12_51_groupi_n_721, csa_tree_add_12_51_groupi_n_722, csa_tree_add_12_51_groupi_n_723, csa_tree_add_12_51_groupi_n_724, csa_tree_add_12_51_groupi_n_725, csa_tree_add_12_51_groupi_n_726, csa_tree_add_12_51_groupi_n_727, csa_tree_add_12_51_groupi_n_728;
  wire csa_tree_add_12_51_groupi_n_729, csa_tree_add_12_51_groupi_n_730, csa_tree_add_12_51_groupi_n_731, csa_tree_add_12_51_groupi_n_732, csa_tree_add_12_51_groupi_n_733, csa_tree_add_12_51_groupi_n_734, csa_tree_add_12_51_groupi_n_735, csa_tree_add_12_51_groupi_n_736;
  wire csa_tree_add_12_51_groupi_n_737, csa_tree_add_12_51_groupi_n_738, csa_tree_add_12_51_groupi_n_739, csa_tree_add_12_51_groupi_n_740, csa_tree_add_12_51_groupi_n_741, csa_tree_add_12_51_groupi_n_742, csa_tree_add_12_51_groupi_n_743, csa_tree_add_12_51_groupi_n_744;
  wire csa_tree_add_12_51_groupi_n_745, csa_tree_add_12_51_groupi_n_746, csa_tree_add_12_51_groupi_n_747, csa_tree_add_12_51_groupi_n_748, csa_tree_add_12_51_groupi_n_749, csa_tree_add_12_51_groupi_n_750, csa_tree_add_12_51_groupi_n_751, csa_tree_add_12_51_groupi_n_752;
  wire csa_tree_add_12_51_groupi_n_753, csa_tree_add_12_51_groupi_n_754, csa_tree_add_12_51_groupi_n_755, csa_tree_add_12_51_groupi_n_756, csa_tree_add_12_51_groupi_n_757, csa_tree_add_12_51_groupi_n_758, csa_tree_add_12_51_groupi_n_759, csa_tree_add_12_51_groupi_n_760;
  wire csa_tree_add_12_51_groupi_n_761, csa_tree_add_12_51_groupi_n_762, csa_tree_add_12_51_groupi_n_763, csa_tree_add_12_51_groupi_n_764, csa_tree_add_12_51_groupi_n_765, csa_tree_add_12_51_groupi_n_766, csa_tree_add_12_51_groupi_n_767, csa_tree_add_12_51_groupi_n_768;
  wire csa_tree_add_12_51_groupi_n_769, csa_tree_add_12_51_groupi_n_770, csa_tree_add_12_51_groupi_n_771, csa_tree_add_12_51_groupi_n_772, csa_tree_add_12_51_groupi_n_773, csa_tree_add_12_51_groupi_n_774, csa_tree_add_12_51_groupi_n_775, csa_tree_add_12_51_groupi_n_776;
  wire csa_tree_add_12_51_groupi_n_777, csa_tree_add_12_51_groupi_n_778, csa_tree_add_12_51_groupi_n_779, csa_tree_add_12_51_groupi_n_780, csa_tree_add_12_51_groupi_n_781, csa_tree_add_12_51_groupi_n_782, csa_tree_add_12_51_groupi_n_783, csa_tree_add_12_51_groupi_n_784;
  wire csa_tree_add_12_51_groupi_n_785, csa_tree_add_12_51_groupi_n_786, csa_tree_add_12_51_groupi_n_787, csa_tree_add_12_51_groupi_n_788, csa_tree_add_12_51_groupi_n_789, csa_tree_add_12_51_groupi_n_790, csa_tree_add_12_51_groupi_n_791, csa_tree_add_12_51_groupi_n_792;
  wire csa_tree_add_12_51_groupi_n_793, csa_tree_add_12_51_groupi_n_794, csa_tree_add_12_51_groupi_n_795, csa_tree_add_12_51_groupi_n_796, csa_tree_add_12_51_groupi_n_797, csa_tree_add_12_51_groupi_n_798, csa_tree_add_12_51_groupi_n_799, csa_tree_add_12_51_groupi_n_800;
  wire csa_tree_add_12_51_groupi_n_801, csa_tree_add_12_51_groupi_n_802, csa_tree_add_12_51_groupi_n_803, csa_tree_add_12_51_groupi_n_804, csa_tree_add_12_51_groupi_n_805, csa_tree_add_12_51_groupi_n_806, csa_tree_add_12_51_groupi_n_807, csa_tree_add_12_51_groupi_n_808;
  wire csa_tree_add_12_51_groupi_n_809, csa_tree_add_12_51_groupi_n_810, csa_tree_add_12_51_groupi_n_811, csa_tree_add_12_51_groupi_n_812, csa_tree_add_12_51_groupi_n_813, csa_tree_add_12_51_groupi_n_814, csa_tree_add_12_51_groupi_n_815, csa_tree_add_12_51_groupi_n_816;
  wire csa_tree_add_12_51_groupi_n_817, csa_tree_add_12_51_groupi_n_818, csa_tree_add_12_51_groupi_n_819, csa_tree_add_12_51_groupi_n_820, csa_tree_add_12_51_groupi_n_821, csa_tree_add_12_51_groupi_n_822, csa_tree_add_12_51_groupi_n_823, csa_tree_add_12_51_groupi_n_824;
  wire csa_tree_add_12_51_groupi_n_825, csa_tree_add_12_51_groupi_n_826, csa_tree_add_12_51_groupi_n_827, csa_tree_add_12_51_groupi_n_828, csa_tree_add_12_51_groupi_n_829, csa_tree_add_12_51_groupi_n_830, csa_tree_add_12_51_groupi_n_831, csa_tree_add_12_51_groupi_n_832;
  wire csa_tree_add_12_51_groupi_n_833, csa_tree_add_12_51_groupi_n_834, csa_tree_add_12_51_groupi_n_835, csa_tree_add_12_51_groupi_n_836, csa_tree_add_12_51_groupi_n_837, csa_tree_add_12_51_groupi_n_838, csa_tree_add_12_51_groupi_n_839, csa_tree_add_12_51_groupi_n_840;
  wire csa_tree_add_12_51_groupi_n_841, csa_tree_add_12_51_groupi_n_842, csa_tree_add_12_51_groupi_n_843, csa_tree_add_12_51_groupi_n_844, csa_tree_add_12_51_groupi_n_845, csa_tree_add_12_51_groupi_n_846, csa_tree_add_12_51_groupi_n_847, csa_tree_add_12_51_groupi_n_848;
  wire csa_tree_add_12_51_groupi_n_849, csa_tree_add_12_51_groupi_n_850, csa_tree_add_12_51_groupi_n_851, csa_tree_add_12_51_groupi_n_852, csa_tree_add_12_51_groupi_n_853, csa_tree_add_12_51_groupi_n_854, csa_tree_add_12_51_groupi_n_855, csa_tree_add_12_51_groupi_n_856;
  wire csa_tree_add_12_51_groupi_n_857, csa_tree_add_12_51_groupi_n_858, csa_tree_add_12_51_groupi_n_859, csa_tree_add_12_51_groupi_n_860, csa_tree_add_12_51_groupi_n_861, csa_tree_add_12_51_groupi_n_862, csa_tree_add_12_51_groupi_n_863, csa_tree_add_12_51_groupi_n_864;
  wire csa_tree_add_12_51_groupi_n_865, csa_tree_add_12_51_groupi_n_866, csa_tree_add_12_51_groupi_n_867, csa_tree_add_12_51_groupi_n_868, csa_tree_add_12_51_groupi_n_869, csa_tree_add_12_51_groupi_n_870, csa_tree_add_12_51_groupi_n_871, csa_tree_add_12_51_groupi_n_872;
  wire csa_tree_add_12_51_groupi_n_873, csa_tree_add_12_51_groupi_n_874, csa_tree_add_12_51_groupi_n_875, csa_tree_add_12_51_groupi_n_876, csa_tree_add_12_51_groupi_n_877, csa_tree_add_12_51_groupi_n_878, csa_tree_add_12_51_groupi_n_879, csa_tree_add_12_51_groupi_n_880;
  wire csa_tree_add_12_51_groupi_n_881, csa_tree_add_12_51_groupi_n_882, csa_tree_add_12_51_groupi_n_883, csa_tree_add_12_51_groupi_n_884, csa_tree_add_12_51_groupi_n_885, csa_tree_add_12_51_groupi_n_886, csa_tree_add_12_51_groupi_n_887, csa_tree_add_12_51_groupi_n_888;
  wire csa_tree_add_12_51_groupi_n_889, csa_tree_add_12_51_groupi_n_890, csa_tree_add_12_51_groupi_n_891, csa_tree_add_12_51_groupi_n_892, csa_tree_add_12_51_groupi_n_893, csa_tree_add_12_51_groupi_n_894, csa_tree_add_12_51_groupi_n_895, csa_tree_add_12_51_groupi_n_896;
  wire csa_tree_add_12_51_groupi_n_897, csa_tree_add_12_51_groupi_n_898, csa_tree_add_12_51_groupi_n_899, csa_tree_add_12_51_groupi_n_900, csa_tree_add_12_51_groupi_n_901, csa_tree_add_12_51_groupi_n_902, csa_tree_add_12_51_groupi_n_903, csa_tree_add_12_51_groupi_n_904;
  wire csa_tree_add_12_51_groupi_n_905, csa_tree_add_12_51_groupi_n_906, csa_tree_add_12_51_groupi_n_907, csa_tree_add_12_51_groupi_n_908, csa_tree_add_12_51_groupi_n_909, csa_tree_add_12_51_groupi_n_910, csa_tree_add_12_51_groupi_n_911, csa_tree_add_12_51_groupi_n_912;
  wire csa_tree_add_12_51_groupi_n_913, csa_tree_add_12_51_groupi_n_914, csa_tree_add_12_51_groupi_n_915, csa_tree_add_12_51_groupi_n_916, csa_tree_add_12_51_groupi_n_917, csa_tree_add_12_51_groupi_n_918, csa_tree_add_12_51_groupi_n_919, csa_tree_add_12_51_groupi_n_920;
  wire csa_tree_add_12_51_groupi_n_921, csa_tree_add_12_51_groupi_n_922, csa_tree_add_12_51_groupi_n_923, csa_tree_add_12_51_groupi_n_924, csa_tree_add_12_51_groupi_n_925, csa_tree_add_12_51_groupi_n_926, csa_tree_add_12_51_groupi_n_927, csa_tree_add_12_51_groupi_n_928;
  wire csa_tree_add_12_51_groupi_n_929, csa_tree_add_12_51_groupi_n_930, csa_tree_add_12_51_groupi_n_931, csa_tree_add_12_51_groupi_n_932, csa_tree_add_12_51_groupi_n_933, csa_tree_add_12_51_groupi_n_934, csa_tree_add_12_51_groupi_n_935, csa_tree_add_12_51_groupi_n_936;
  wire csa_tree_add_12_51_groupi_n_937, csa_tree_add_12_51_groupi_n_938, csa_tree_add_12_51_groupi_n_939, csa_tree_add_12_51_groupi_n_940, csa_tree_add_12_51_groupi_n_941, csa_tree_add_12_51_groupi_n_942, csa_tree_add_12_51_groupi_n_943, csa_tree_add_12_51_groupi_n_944;
  wire csa_tree_add_12_51_groupi_n_945, csa_tree_add_12_51_groupi_n_946, csa_tree_add_12_51_groupi_n_947, csa_tree_add_12_51_groupi_n_948, csa_tree_add_12_51_groupi_n_949, csa_tree_add_12_51_groupi_n_950, csa_tree_add_12_51_groupi_n_951, csa_tree_add_12_51_groupi_n_952;
  wire csa_tree_add_12_51_groupi_n_953, csa_tree_add_12_51_groupi_n_954, csa_tree_add_12_51_groupi_n_955, csa_tree_add_12_51_groupi_n_956, csa_tree_add_12_51_groupi_n_957, csa_tree_add_12_51_groupi_n_958, csa_tree_add_12_51_groupi_n_959, csa_tree_add_12_51_groupi_n_960;
  wire csa_tree_add_12_51_groupi_n_961, csa_tree_add_12_51_groupi_n_962, csa_tree_add_12_51_groupi_n_963, csa_tree_add_12_51_groupi_n_964, csa_tree_add_12_51_groupi_n_965, csa_tree_add_12_51_groupi_n_966, csa_tree_add_12_51_groupi_n_967, csa_tree_add_12_51_groupi_n_968;
  wire csa_tree_add_12_51_groupi_n_969, csa_tree_add_12_51_groupi_n_970, csa_tree_add_12_51_groupi_n_971, csa_tree_add_12_51_groupi_n_972, csa_tree_add_12_51_groupi_n_973, csa_tree_add_12_51_groupi_n_974, csa_tree_add_12_51_groupi_n_975, csa_tree_add_12_51_groupi_n_976;
  wire csa_tree_add_12_51_groupi_n_977, csa_tree_add_12_51_groupi_n_978, csa_tree_add_12_51_groupi_n_979, csa_tree_add_12_51_groupi_n_980, csa_tree_add_12_51_groupi_n_981, csa_tree_add_12_51_groupi_n_982, csa_tree_add_12_51_groupi_n_983, csa_tree_add_12_51_groupi_n_984;
  wire csa_tree_add_12_51_groupi_n_985, csa_tree_add_12_51_groupi_n_986, csa_tree_add_12_51_groupi_n_987, csa_tree_add_12_51_groupi_n_988, csa_tree_add_12_51_groupi_n_989, csa_tree_add_12_51_groupi_n_990, csa_tree_add_12_51_groupi_n_991, csa_tree_add_12_51_groupi_n_992;
  wire csa_tree_add_12_51_groupi_n_993, csa_tree_add_12_51_groupi_n_994, csa_tree_add_12_51_groupi_n_995, csa_tree_add_12_51_groupi_n_996, csa_tree_add_12_51_groupi_n_997, csa_tree_add_12_51_groupi_n_998, csa_tree_add_12_51_groupi_n_999, csa_tree_add_12_51_groupi_n_1000;
  wire csa_tree_add_12_51_groupi_n_1001, csa_tree_add_12_51_groupi_n_1002, csa_tree_add_12_51_groupi_n_1003, csa_tree_add_12_51_groupi_n_1004, csa_tree_add_12_51_groupi_n_1005, csa_tree_add_12_51_groupi_n_1006, csa_tree_add_12_51_groupi_n_1007, csa_tree_add_12_51_groupi_n_1008;
  wire csa_tree_add_12_51_groupi_n_1009, csa_tree_add_12_51_groupi_n_1010, csa_tree_add_12_51_groupi_n_1011, csa_tree_add_12_51_groupi_n_1012, csa_tree_add_12_51_groupi_n_1013, csa_tree_add_12_51_groupi_n_1014, csa_tree_add_12_51_groupi_n_1015, csa_tree_add_12_51_groupi_n_1016;
  wire csa_tree_add_12_51_groupi_n_1017, csa_tree_add_12_51_groupi_n_1018, csa_tree_add_12_51_groupi_n_1019, csa_tree_add_12_51_groupi_n_1020, csa_tree_add_12_51_groupi_n_1021, csa_tree_add_12_51_groupi_n_1022, csa_tree_add_12_51_groupi_n_1023, csa_tree_add_12_51_groupi_n_1024;
  wire csa_tree_add_12_51_groupi_n_1025, csa_tree_add_12_51_groupi_n_1026, csa_tree_add_12_51_groupi_n_1027, csa_tree_add_12_51_groupi_n_1028, csa_tree_add_12_51_groupi_n_1029, csa_tree_add_12_51_groupi_n_1030, csa_tree_add_12_51_groupi_n_1031, csa_tree_add_12_51_groupi_n_1032;
  wire csa_tree_add_12_51_groupi_n_1033, csa_tree_add_12_51_groupi_n_1034, csa_tree_add_12_51_groupi_n_1035, csa_tree_add_12_51_groupi_n_1036, csa_tree_add_12_51_groupi_n_1037, csa_tree_add_12_51_groupi_n_1038, csa_tree_add_12_51_groupi_n_1039, csa_tree_add_12_51_groupi_n_1040;
  wire csa_tree_add_12_51_groupi_n_1041, csa_tree_add_12_51_groupi_n_1042, csa_tree_add_12_51_groupi_n_1043, csa_tree_add_12_51_groupi_n_1044, csa_tree_add_12_51_groupi_n_1045, csa_tree_add_12_51_groupi_n_1046, csa_tree_add_12_51_groupi_n_1047, csa_tree_add_12_51_groupi_n_1048;
  wire csa_tree_add_12_51_groupi_n_1049, csa_tree_add_12_51_groupi_n_1050, csa_tree_add_12_51_groupi_n_1051, csa_tree_add_12_51_groupi_n_1052, csa_tree_add_12_51_groupi_n_1053, csa_tree_add_12_51_groupi_n_1054, csa_tree_add_12_51_groupi_n_1055, csa_tree_add_12_51_groupi_n_1056;
  wire csa_tree_add_12_51_groupi_n_1057, csa_tree_add_12_51_groupi_n_1058, csa_tree_add_12_51_groupi_n_1059, csa_tree_add_12_51_groupi_n_1060, csa_tree_add_12_51_groupi_n_1061, csa_tree_add_12_51_groupi_n_1062, csa_tree_add_12_51_groupi_n_1063, csa_tree_add_12_51_groupi_n_1064;
  wire csa_tree_add_12_51_groupi_n_1065, csa_tree_add_12_51_groupi_n_1066, csa_tree_add_12_51_groupi_n_1067, csa_tree_add_12_51_groupi_n_1068, csa_tree_add_12_51_groupi_n_1069, csa_tree_add_12_51_groupi_n_1070, csa_tree_add_12_51_groupi_n_1071, csa_tree_add_12_51_groupi_n_1072;
  wire csa_tree_add_12_51_groupi_n_1073, csa_tree_add_12_51_groupi_n_1074, csa_tree_add_12_51_groupi_n_1075, csa_tree_add_12_51_groupi_n_1076, csa_tree_add_12_51_groupi_n_1077, csa_tree_add_12_51_groupi_n_1078, csa_tree_add_12_51_groupi_n_1079, csa_tree_add_12_51_groupi_n_1080;
  wire csa_tree_add_12_51_groupi_n_1081, csa_tree_add_12_51_groupi_n_1082, csa_tree_add_12_51_groupi_n_1083, csa_tree_add_12_51_groupi_n_1084, csa_tree_add_12_51_groupi_n_1085, csa_tree_add_12_51_groupi_n_1086, csa_tree_add_12_51_groupi_n_1087, csa_tree_add_12_51_groupi_n_1088;
  wire csa_tree_add_12_51_groupi_n_1089, csa_tree_add_12_51_groupi_n_1090, csa_tree_add_12_51_groupi_n_1091, csa_tree_add_12_51_groupi_n_1092, csa_tree_add_12_51_groupi_n_1093, csa_tree_add_12_51_groupi_n_1094, csa_tree_add_12_51_groupi_n_1095, csa_tree_add_12_51_groupi_n_1096;
  wire csa_tree_add_12_51_groupi_n_1097, csa_tree_add_12_51_groupi_n_1098, csa_tree_add_12_51_groupi_n_1099, csa_tree_add_12_51_groupi_n_1100, csa_tree_add_12_51_groupi_n_1101, csa_tree_add_12_51_groupi_n_1102, csa_tree_add_12_51_groupi_n_1103, csa_tree_add_12_51_groupi_n_1104;
  wire csa_tree_add_12_51_groupi_n_1105, csa_tree_add_12_51_groupi_n_1106, csa_tree_add_12_51_groupi_n_1107, csa_tree_add_12_51_groupi_n_1108, csa_tree_add_12_51_groupi_n_1109, csa_tree_add_12_51_groupi_n_1110, csa_tree_add_12_51_groupi_n_1111, csa_tree_add_12_51_groupi_n_1112;
  wire csa_tree_add_12_51_groupi_n_1113, csa_tree_add_12_51_groupi_n_1114, csa_tree_add_12_51_groupi_n_1115, csa_tree_add_12_51_groupi_n_1116, csa_tree_add_12_51_groupi_n_1117, csa_tree_add_12_51_groupi_n_1118, csa_tree_add_12_51_groupi_n_1119, csa_tree_add_12_51_groupi_n_1120;
  wire csa_tree_add_12_51_groupi_n_1121, csa_tree_add_12_51_groupi_n_1122, csa_tree_add_12_51_groupi_n_1123, csa_tree_add_12_51_groupi_n_1124, csa_tree_add_12_51_groupi_n_1125, csa_tree_add_12_51_groupi_n_1126, csa_tree_add_12_51_groupi_n_1127, csa_tree_add_12_51_groupi_n_1128;
  wire csa_tree_add_12_51_groupi_n_1129, csa_tree_add_12_51_groupi_n_1130, csa_tree_add_12_51_groupi_n_1131, csa_tree_add_12_51_groupi_n_1132, csa_tree_add_12_51_groupi_n_1133, csa_tree_add_12_51_groupi_n_1134, csa_tree_add_12_51_groupi_n_1135, csa_tree_add_12_51_groupi_n_1136;
  wire csa_tree_add_12_51_groupi_n_1137, csa_tree_add_12_51_groupi_n_1138, csa_tree_add_12_51_groupi_n_1139, csa_tree_add_12_51_groupi_n_1140, csa_tree_add_12_51_groupi_n_1141, csa_tree_add_12_51_groupi_n_1142, csa_tree_add_12_51_groupi_n_1143, csa_tree_add_12_51_groupi_n_1144;
  wire csa_tree_add_12_51_groupi_n_1145, csa_tree_add_12_51_groupi_n_1146, csa_tree_add_12_51_groupi_n_1147, csa_tree_add_12_51_groupi_n_1148, csa_tree_add_12_51_groupi_n_1149, csa_tree_add_12_51_groupi_n_1150, csa_tree_add_12_51_groupi_n_1151, csa_tree_add_12_51_groupi_n_1152;
  wire csa_tree_add_12_51_groupi_n_1153, csa_tree_add_12_51_groupi_n_1154, csa_tree_add_12_51_groupi_n_1155, csa_tree_add_12_51_groupi_n_1156, csa_tree_add_12_51_groupi_n_1157, csa_tree_add_12_51_groupi_n_1158, csa_tree_add_12_51_groupi_n_1159, csa_tree_add_12_51_groupi_n_1160;
  wire csa_tree_add_12_51_groupi_n_1161, csa_tree_add_12_51_groupi_n_1162, csa_tree_add_12_51_groupi_n_1163, csa_tree_add_12_51_groupi_n_1164, csa_tree_add_12_51_groupi_n_1165, csa_tree_add_12_51_groupi_n_1166, csa_tree_add_12_51_groupi_n_1167, csa_tree_add_12_51_groupi_n_1168;
  wire csa_tree_add_12_51_groupi_n_1169, csa_tree_add_12_51_groupi_n_1170, csa_tree_add_12_51_groupi_n_1171, csa_tree_add_12_51_groupi_n_1172, csa_tree_add_12_51_groupi_n_1173, csa_tree_add_12_51_groupi_n_1174, csa_tree_add_12_51_groupi_n_1175, csa_tree_add_12_51_groupi_n_1176;
  wire csa_tree_add_12_51_groupi_n_1177, csa_tree_add_12_51_groupi_n_1178, csa_tree_add_12_51_groupi_n_1179, csa_tree_add_12_51_groupi_n_1180, csa_tree_add_12_51_groupi_n_1181, csa_tree_add_12_51_groupi_n_1182, csa_tree_add_12_51_groupi_n_1183, csa_tree_add_12_51_groupi_n_1184;
  wire csa_tree_add_12_51_groupi_n_1185, csa_tree_add_12_51_groupi_n_1186, csa_tree_add_12_51_groupi_n_1187, csa_tree_add_12_51_groupi_n_1188, csa_tree_add_12_51_groupi_n_1189, csa_tree_add_12_51_groupi_n_1190, csa_tree_add_12_51_groupi_n_1191, csa_tree_add_12_51_groupi_n_1192;
  wire csa_tree_add_12_51_groupi_n_1193, csa_tree_add_12_51_groupi_n_1194, csa_tree_add_12_51_groupi_n_1195, csa_tree_add_12_51_groupi_n_1196, csa_tree_add_12_51_groupi_n_1197, csa_tree_add_12_51_groupi_n_1198, csa_tree_add_12_51_groupi_n_1199, csa_tree_add_12_51_groupi_n_1200;
  wire csa_tree_add_12_51_groupi_n_1201, csa_tree_add_12_51_groupi_n_1202, csa_tree_add_12_51_groupi_n_1203, csa_tree_add_12_51_groupi_n_1204, csa_tree_add_12_51_groupi_n_1205, csa_tree_add_12_51_groupi_n_1206, csa_tree_add_12_51_groupi_n_1207, csa_tree_add_12_51_groupi_n_1208;
  wire csa_tree_add_12_51_groupi_n_1209, csa_tree_add_12_51_groupi_n_1210, csa_tree_add_12_51_groupi_n_1211, csa_tree_add_12_51_groupi_n_1212, csa_tree_add_12_51_groupi_n_1213, csa_tree_add_12_51_groupi_n_1214, csa_tree_add_12_51_groupi_n_1215, csa_tree_add_12_51_groupi_n_1216;
  wire csa_tree_add_12_51_groupi_n_1217, csa_tree_add_12_51_groupi_n_1218, csa_tree_add_12_51_groupi_n_1219, csa_tree_add_12_51_groupi_n_1220, csa_tree_add_12_51_groupi_n_1221, csa_tree_add_12_51_groupi_n_1222, csa_tree_add_12_51_groupi_n_1223, csa_tree_add_12_51_groupi_n_1224;
  wire csa_tree_add_12_51_groupi_n_1225, csa_tree_add_12_51_groupi_n_1226, csa_tree_add_12_51_groupi_n_1227, csa_tree_add_12_51_groupi_n_1228, csa_tree_add_12_51_groupi_n_1229, csa_tree_add_12_51_groupi_n_1230, csa_tree_add_12_51_groupi_n_1231, csa_tree_add_12_51_groupi_n_1232;
  wire csa_tree_add_12_51_groupi_n_1233, csa_tree_add_12_51_groupi_n_1234, csa_tree_add_12_51_groupi_n_1235, csa_tree_add_12_51_groupi_n_1236, csa_tree_add_12_51_groupi_n_1237, csa_tree_add_12_51_groupi_n_1238, csa_tree_add_12_51_groupi_n_1239, csa_tree_add_12_51_groupi_n_1240;
  wire csa_tree_add_12_51_groupi_n_1241, csa_tree_add_12_51_groupi_n_1242, csa_tree_add_12_51_groupi_n_1243, csa_tree_add_12_51_groupi_n_1244, csa_tree_add_12_51_groupi_n_1245, csa_tree_add_12_51_groupi_n_1246, csa_tree_add_12_51_groupi_n_1247, csa_tree_add_12_51_groupi_n_1248;
  wire csa_tree_add_12_51_groupi_n_1249, csa_tree_add_12_51_groupi_n_1250, csa_tree_add_12_51_groupi_n_1251, csa_tree_add_12_51_groupi_n_1252, csa_tree_add_12_51_groupi_n_1253, csa_tree_add_12_51_groupi_n_1254, csa_tree_add_12_51_groupi_n_1255, csa_tree_add_12_51_groupi_n_1256;
  wire csa_tree_add_12_51_groupi_n_1257, csa_tree_add_12_51_groupi_n_1258, csa_tree_add_12_51_groupi_n_1259, csa_tree_add_12_51_groupi_n_1260, csa_tree_add_12_51_groupi_n_1261, csa_tree_add_12_51_groupi_n_1262, csa_tree_add_12_51_groupi_n_1263, csa_tree_add_12_51_groupi_n_1264;
  wire csa_tree_add_12_51_groupi_n_1265, csa_tree_add_12_51_groupi_n_1266, csa_tree_add_12_51_groupi_n_1267, csa_tree_add_12_51_groupi_n_1268, csa_tree_add_12_51_groupi_n_1269, csa_tree_add_12_51_groupi_n_1270, csa_tree_add_12_51_groupi_n_1271, csa_tree_add_12_51_groupi_n_1272;
  wire csa_tree_add_12_51_groupi_n_1273, csa_tree_add_12_51_groupi_n_1274, csa_tree_add_12_51_groupi_n_1275, csa_tree_add_12_51_groupi_n_1276, csa_tree_add_12_51_groupi_n_1277, csa_tree_add_12_51_groupi_n_1278, csa_tree_add_12_51_groupi_n_1279, csa_tree_add_12_51_groupi_n_1280;
  wire csa_tree_add_12_51_groupi_n_1281, csa_tree_add_12_51_groupi_n_1282, csa_tree_add_12_51_groupi_n_1283, csa_tree_add_12_51_groupi_n_1284, csa_tree_add_12_51_groupi_n_1285, csa_tree_add_12_51_groupi_n_1286, csa_tree_add_12_51_groupi_n_1287, csa_tree_add_12_51_groupi_n_1288;
  wire csa_tree_add_12_51_groupi_n_1289, csa_tree_add_12_51_groupi_n_1290, csa_tree_add_12_51_groupi_n_1291, csa_tree_add_12_51_groupi_n_1292, csa_tree_add_12_51_groupi_n_1293, csa_tree_add_12_51_groupi_n_1294, csa_tree_add_12_51_groupi_n_1295, csa_tree_add_12_51_groupi_n_1296;
  wire csa_tree_add_12_51_groupi_n_1297, csa_tree_add_12_51_groupi_n_1298, csa_tree_add_12_51_groupi_n_1299, csa_tree_add_12_51_groupi_n_1300, csa_tree_add_12_51_groupi_n_1301, csa_tree_add_12_51_groupi_n_1302, csa_tree_add_12_51_groupi_n_1303, csa_tree_add_12_51_groupi_n_1304;
  wire csa_tree_add_12_51_groupi_n_1305, csa_tree_add_12_51_groupi_n_1306, csa_tree_add_12_51_groupi_n_1307, csa_tree_add_12_51_groupi_n_1308, csa_tree_add_12_51_groupi_n_1309, csa_tree_add_12_51_groupi_n_1310, csa_tree_add_12_51_groupi_n_1311, csa_tree_add_12_51_groupi_n_1312;
  wire csa_tree_add_12_51_groupi_n_1313, csa_tree_add_12_51_groupi_n_1314, csa_tree_add_12_51_groupi_n_1315, csa_tree_add_12_51_groupi_n_1316, csa_tree_add_12_51_groupi_n_1317, csa_tree_add_12_51_groupi_n_1318, csa_tree_add_12_51_groupi_n_1319, csa_tree_add_12_51_groupi_n_1320;
  wire csa_tree_add_12_51_groupi_n_1321, csa_tree_add_12_51_groupi_n_1322, csa_tree_add_12_51_groupi_n_1323, csa_tree_add_12_51_groupi_n_1324, csa_tree_add_12_51_groupi_n_1325, csa_tree_add_12_51_groupi_n_1326, csa_tree_add_12_51_groupi_n_1327, csa_tree_add_12_51_groupi_n_1328;
  wire csa_tree_add_12_51_groupi_n_1329, csa_tree_add_12_51_groupi_n_1330, csa_tree_add_12_51_groupi_n_1331, csa_tree_add_12_51_groupi_n_1332, csa_tree_add_12_51_groupi_n_1333, csa_tree_add_12_51_groupi_n_1334, csa_tree_add_12_51_groupi_n_1335, csa_tree_add_12_51_groupi_n_1336;
  wire csa_tree_add_12_51_groupi_n_1337, csa_tree_add_12_51_groupi_n_1338, csa_tree_add_12_51_groupi_n_1339, csa_tree_add_12_51_groupi_n_1340, csa_tree_add_12_51_groupi_n_1341, csa_tree_add_12_51_groupi_n_1342, csa_tree_add_12_51_groupi_n_1343, csa_tree_add_12_51_groupi_n_1344;
  wire csa_tree_add_12_51_groupi_n_1345, csa_tree_add_12_51_groupi_n_1346, csa_tree_add_12_51_groupi_n_1347, csa_tree_add_12_51_groupi_n_1348, csa_tree_add_12_51_groupi_n_1349, csa_tree_add_12_51_groupi_n_1350, csa_tree_add_12_51_groupi_n_1351, csa_tree_add_12_51_groupi_n_1352;
  wire csa_tree_add_12_51_groupi_n_1353, csa_tree_add_12_51_groupi_n_1354, csa_tree_add_12_51_groupi_n_1355, csa_tree_add_12_51_groupi_n_1356, csa_tree_add_12_51_groupi_n_1357, csa_tree_add_12_51_groupi_n_1358, csa_tree_add_12_51_groupi_n_1359, csa_tree_add_12_51_groupi_n_1360;
  wire csa_tree_add_12_51_groupi_n_1361, csa_tree_add_12_51_groupi_n_1362, csa_tree_add_12_51_groupi_n_1363, csa_tree_add_12_51_groupi_n_1364, csa_tree_add_12_51_groupi_n_1365, csa_tree_add_12_51_groupi_n_1366, csa_tree_add_12_51_groupi_n_1367, csa_tree_add_12_51_groupi_n_1368;
  wire csa_tree_add_12_51_groupi_n_1369, csa_tree_add_12_51_groupi_n_1370, csa_tree_add_12_51_groupi_n_1371, csa_tree_add_12_51_groupi_n_1372, csa_tree_add_12_51_groupi_n_1373, csa_tree_add_12_51_groupi_n_1374, csa_tree_add_12_51_groupi_n_1375, csa_tree_add_12_51_groupi_n_1376;
  wire csa_tree_add_12_51_groupi_n_1377, csa_tree_add_12_51_groupi_n_1378, csa_tree_add_12_51_groupi_n_1379, csa_tree_add_12_51_groupi_n_1380, csa_tree_add_12_51_groupi_n_1381, csa_tree_add_12_51_groupi_n_1382, csa_tree_add_12_51_groupi_n_1383, csa_tree_add_12_51_groupi_n_1384;
  wire csa_tree_add_12_51_groupi_n_1385, csa_tree_add_12_51_groupi_n_1386, csa_tree_add_12_51_groupi_n_1387, csa_tree_add_12_51_groupi_n_1388, csa_tree_add_12_51_groupi_n_1389, csa_tree_add_12_51_groupi_n_1390, csa_tree_add_12_51_groupi_n_1391, csa_tree_add_12_51_groupi_n_1392;
  wire csa_tree_add_12_51_groupi_n_1393, csa_tree_add_12_51_groupi_n_1394, csa_tree_add_12_51_groupi_n_1395, csa_tree_add_12_51_groupi_n_1396, csa_tree_add_12_51_groupi_n_1397, csa_tree_add_12_51_groupi_n_1398, csa_tree_add_12_51_groupi_n_1399, csa_tree_add_12_51_groupi_n_1400;
  wire csa_tree_add_12_51_groupi_n_1401, csa_tree_add_12_51_groupi_n_1402, csa_tree_add_12_51_groupi_n_1403, csa_tree_add_12_51_groupi_n_1404, csa_tree_add_12_51_groupi_n_1405, csa_tree_add_12_51_groupi_n_1406, csa_tree_add_12_51_groupi_n_1407, csa_tree_add_12_51_groupi_n_1408;
  wire csa_tree_add_12_51_groupi_n_1409, csa_tree_add_12_51_groupi_n_1410, csa_tree_add_12_51_groupi_n_1411, csa_tree_add_12_51_groupi_n_1412, csa_tree_add_12_51_groupi_n_1413, csa_tree_add_12_51_groupi_n_1414, csa_tree_add_12_51_groupi_n_1415, csa_tree_add_12_51_groupi_n_1416;
  wire csa_tree_add_12_51_groupi_n_1417, csa_tree_add_12_51_groupi_n_1418, csa_tree_add_12_51_groupi_n_1419, csa_tree_add_12_51_groupi_n_1420, csa_tree_add_12_51_groupi_n_1421, csa_tree_add_12_51_groupi_n_1422, csa_tree_add_12_51_groupi_n_1423, csa_tree_add_12_51_groupi_n_1424;
  wire csa_tree_add_12_51_groupi_n_1425, csa_tree_add_12_51_groupi_n_1426, csa_tree_add_12_51_groupi_n_1427, csa_tree_add_12_51_groupi_n_1428, csa_tree_add_12_51_groupi_n_1429, csa_tree_add_12_51_groupi_n_1430, csa_tree_add_12_51_groupi_n_1431, csa_tree_add_12_51_groupi_n_1432;
  wire csa_tree_add_12_51_groupi_n_1433, csa_tree_add_12_51_groupi_n_1434, csa_tree_add_12_51_groupi_n_1435, csa_tree_add_12_51_groupi_n_1436, csa_tree_add_12_51_groupi_n_1437, csa_tree_add_12_51_groupi_n_1438, csa_tree_add_12_51_groupi_n_1439, csa_tree_add_12_51_groupi_n_1440;
  wire csa_tree_add_12_51_groupi_n_1441, csa_tree_add_12_51_groupi_n_1442, csa_tree_add_12_51_groupi_n_1443, csa_tree_add_12_51_groupi_n_1444, csa_tree_add_12_51_groupi_n_1445, csa_tree_add_12_51_groupi_n_1446, csa_tree_add_12_51_groupi_n_1447, csa_tree_add_12_51_groupi_n_1448;
  wire csa_tree_add_12_51_groupi_n_1449, csa_tree_add_12_51_groupi_n_1450, csa_tree_add_12_51_groupi_n_1451, csa_tree_add_12_51_groupi_n_1452, csa_tree_add_12_51_groupi_n_1453, csa_tree_add_12_51_groupi_n_1454, csa_tree_add_12_51_groupi_n_1455, csa_tree_add_12_51_groupi_n_1456;
  wire csa_tree_add_12_51_groupi_n_1457, csa_tree_add_12_51_groupi_n_1458, csa_tree_add_12_51_groupi_n_1459, csa_tree_add_12_51_groupi_n_1460, csa_tree_add_12_51_groupi_n_1461, csa_tree_add_12_51_groupi_n_1462, csa_tree_add_12_51_groupi_n_1463, csa_tree_add_12_51_groupi_n_1464;
  wire csa_tree_add_12_51_groupi_n_1465, csa_tree_add_12_51_groupi_n_1466, csa_tree_add_12_51_groupi_n_1467, csa_tree_add_12_51_groupi_n_1468, csa_tree_add_12_51_groupi_n_1469, csa_tree_add_12_51_groupi_n_1470, csa_tree_add_12_51_groupi_n_1471, csa_tree_add_12_51_groupi_n_1472;
  wire csa_tree_add_12_51_groupi_n_1473, csa_tree_add_12_51_groupi_n_1474, csa_tree_add_12_51_groupi_n_1475, csa_tree_add_12_51_groupi_n_1476, csa_tree_add_12_51_groupi_n_1477, csa_tree_add_12_51_groupi_n_1478, csa_tree_add_12_51_groupi_n_1479, csa_tree_add_12_51_groupi_n_1480;
  wire csa_tree_add_12_51_groupi_n_1481, csa_tree_add_12_51_groupi_n_1482, csa_tree_add_12_51_groupi_n_1483, csa_tree_add_12_51_groupi_n_1484, csa_tree_add_12_51_groupi_n_1485, csa_tree_add_12_51_groupi_n_1486, csa_tree_add_12_51_groupi_n_1487, csa_tree_add_12_51_groupi_n_1488;
  wire csa_tree_add_12_51_groupi_n_1489, csa_tree_add_12_51_groupi_n_1490, csa_tree_add_12_51_groupi_n_1491, csa_tree_add_12_51_groupi_n_1492, csa_tree_add_12_51_groupi_n_1493, csa_tree_add_12_51_groupi_n_1494, csa_tree_add_12_51_groupi_n_1495, csa_tree_add_12_51_groupi_n_1496;
  wire csa_tree_add_12_51_groupi_n_1497, csa_tree_add_12_51_groupi_n_1498, csa_tree_add_12_51_groupi_n_1499, csa_tree_add_12_51_groupi_n_1500, csa_tree_add_12_51_groupi_n_1501, csa_tree_add_12_51_groupi_n_1502, csa_tree_add_12_51_groupi_n_1503, csa_tree_add_12_51_groupi_n_1504;
  wire csa_tree_add_12_51_groupi_n_1505, csa_tree_add_12_51_groupi_n_1506, csa_tree_add_12_51_groupi_n_1507, csa_tree_add_12_51_groupi_n_1508, csa_tree_add_12_51_groupi_n_1509, csa_tree_add_12_51_groupi_n_1510, csa_tree_add_12_51_groupi_n_1511, csa_tree_add_12_51_groupi_n_1512;
  wire csa_tree_add_12_51_groupi_n_1513, csa_tree_add_12_51_groupi_n_1514, csa_tree_add_12_51_groupi_n_1515, csa_tree_add_12_51_groupi_n_1516, csa_tree_add_12_51_groupi_n_1517, csa_tree_add_12_51_groupi_n_1518, csa_tree_add_12_51_groupi_n_1519, csa_tree_add_12_51_groupi_n_1520;
  wire csa_tree_add_12_51_groupi_n_1521, csa_tree_add_12_51_groupi_n_1522, csa_tree_add_12_51_groupi_n_1523, csa_tree_add_12_51_groupi_n_1524, csa_tree_add_12_51_groupi_n_1525, csa_tree_add_12_51_groupi_n_1526, csa_tree_add_12_51_groupi_n_1527, csa_tree_add_12_51_groupi_n_1528;
  wire csa_tree_add_12_51_groupi_n_1529, csa_tree_add_12_51_groupi_n_1530, csa_tree_add_12_51_groupi_n_1531, csa_tree_add_12_51_groupi_n_1532, csa_tree_add_12_51_groupi_n_1533, csa_tree_add_12_51_groupi_n_1534, csa_tree_add_12_51_groupi_n_1535, csa_tree_add_12_51_groupi_n_1536;
  wire csa_tree_add_12_51_groupi_n_1537, csa_tree_add_12_51_groupi_n_1538, csa_tree_add_12_51_groupi_n_1539, csa_tree_add_12_51_groupi_n_1540, csa_tree_add_12_51_groupi_n_1541, csa_tree_add_12_51_groupi_n_1542, csa_tree_add_12_51_groupi_n_1543, csa_tree_add_12_51_groupi_n_1544;
  wire csa_tree_add_12_51_groupi_n_1545, csa_tree_add_12_51_groupi_n_1546, csa_tree_add_12_51_groupi_n_1547, csa_tree_add_12_51_groupi_n_1548, csa_tree_add_12_51_groupi_n_1549, csa_tree_add_12_51_groupi_n_1550, csa_tree_add_12_51_groupi_n_1551, csa_tree_add_12_51_groupi_n_1552;
  wire csa_tree_add_12_51_groupi_n_1553, csa_tree_add_12_51_groupi_n_1554, csa_tree_add_12_51_groupi_n_1555, csa_tree_add_12_51_groupi_n_1556, csa_tree_add_12_51_groupi_n_1557, csa_tree_add_12_51_groupi_n_1558, csa_tree_add_12_51_groupi_n_1559, csa_tree_add_12_51_groupi_n_1560;
  wire csa_tree_add_12_51_groupi_n_1561, csa_tree_add_12_51_groupi_n_1562, csa_tree_add_12_51_groupi_n_1563, csa_tree_add_12_51_groupi_n_1564, csa_tree_add_12_51_groupi_n_1565, csa_tree_add_12_51_groupi_n_1566, csa_tree_add_12_51_groupi_n_1567, csa_tree_add_12_51_groupi_n_1568;
  wire csa_tree_add_12_51_groupi_n_1569, csa_tree_add_12_51_groupi_n_1570, csa_tree_add_12_51_groupi_n_1571, csa_tree_add_12_51_groupi_n_1572, csa_tree_add_12_51_groupi_n_1573, csa_tree_add_12_51_groupi_n_1574, csa_tree_add_12_51_groupi_n_1575, csa_tree_add_12_51_groupi_n_1576;
  wire csa_tree_add_12_51_groupi_n_1577, csa_tree_add_12_51_groupi_n_1578, csa_tree_add_12_51_groupi_n_1579, csa_tree_add_12_51_groupi_n_1580, csa_tree_add_12_51_groupi_n_1581, csa_tree_add_12_51_groupi_n_1582, csa_tree_add_12_51_groupi_n_1583, csa_tree_add_12_51_groupi_n_1584;
  wire csa_tree_add_12_51_groupi_n_1585, csa_tree_add_12_51_groupi_n_1586, csa_tree_add_12_51_groupi_n_1587, csa_tree_add_12_51_groupi_n_1588, csa_tree_add_12_51_groupi_n_1589, csa_tree_add_12_51_groupi_n_1590, csa_tree_add_12_51_groupi_n_1591, csa_tree_add_12_51_groupi_n_1592;
  wire csa_tree_add_12_51_groupi_n_1593, csa_tree_add_12_51_groupi_n_1594, csa_tree_add_12_51_groupi_n_1595, csa_tree_add_12_51_groupi_n_1596, csa_tree_add_12_51_groupi_n_1597, csa_tree_add_12_51_groupi_n_1598, csa_tree_add_12_51_groupi_n_1599, csa_tree_add_12_51_groupi_n_1600;
  wire csa_tree_add_12_51_groupi_n_1601, csa_tree_add_12_51_groupi_n_1602, csa_tree_add_12_51_groupi_n_1603, csa_tree_add_12_51_groupi_n_1604, csa_tree_add_12_51_groupi_n_1605, csa_tree_add_12_51_groupi_n_1606, csa_tree_add_12_51_groupi_n_1607, csa_tree_add_12_51_groupi_n_1608;
  wire csa_tree_add_12_51_groupi_n_1609, csa_tree_add_12_51_groupi_n_1610, csa_tree_add_12_51_groupi_n_1611, csa_tree_add_12_51_groupi_n_1612, csa_tree_add_12_51_groupi_n_1613, csa_tree_add_12_51_groupi_n_1614, csa_tree_add_12_51_groupi_n_1615, csa_tree_add_12_51_groupi_n_1616;
  wire csa_tree_add_12_51_groupi_n_1617, csa_tree_add_12_51_groupi_n_1618, csa_tree_add_12_51_groupi_n_1619, csa_tree_add_12_51_groupi_n_1620, csa_tree_add_12_51_groupi_n_1621, csa_tree_add_12_51_groupi_n_1622, csa_tree_add_12_51_groupi_n_1623, csa_tree_add_12_51_groupi_n_1624;
  wire csa_tree_add_12_51_groupi_n_1625, csa_tree_add_12_51_groupi_n_1626, csa_tree_add_12_51_groupi_n_1627, csa_tree_add_12_51_groupi_n_1628, csa_tree_add_12_51_groupi_n_1629, csa_tree_add_12_51_groupi_n_1630, csa_tree_add_12_51_groupi_n_1631, csa_tree_add_12_51_groupi_n_1632;
  wire csa_tree_add_12_51_groupi_n_1633, csa_tree_add_12_51_groupi_n_1634, csa_tree_add_12_51_groupi_n_1635, csa_tree_add_12_51_groupi_n_1636, csa_tree_add_12_51_groupi_n_1637, csa_tree_add_12_51_groupi_n_1638, csa_tree_add_12_51_groupi_n_1639, csa_tree_add_12_51_groupi_n_1640;
  wire csa_tree_add_12_51_groupi_n_1641, csa_tree_add_12_51_groupi_n_1642, csa_tree_add_12_51_groupi_n_1643, csa_tree_add_12_51_groupi_n_1644, csa_tree_add_12_51_groupi_n_1645, csa_tree_add_12_51_groupi_n_1646, csa_tree_add_12_51_groupi_n_1647, csa_tree_add_12_51_groupi_n_1648;
  wire csa_tree_add_12_51_groupi_n_1649, csa_tree_add_12_51_groupi_n_1650, csa_tree_add_12_51_groupi_n_1651, csa_tree_add_12_51_groupi_n_1652, csa_tree_add_12_51_groupi_n_1653, csa_tree_add_12_51_groupi_n_1654, csa_tree_add_12_51_groupi_n_1655, csa_tree_add_12_51_groupi_n_1656;
  wire csa_tree_add_12_51_groupi_n_1657, csa_tree_add_12_51_groupi_n_1658, csa_tree_add_12_51_groupi_n_1659, csa_tree_add_12_51_groupi_n_1660, csa_tree_add_12_51_groupi_n_1661, csa_tree_add_12_51_groupi_n_1662, csa_tree_add_12_51_groupi_n_1663, csa_tree_add_12_51_groupi_n_1664;
  wire csa_tree_add_12_51_groupi_n_1665, csa_tree_add_12_51_groupi_n_1666, csa_tree_add_12_51_groupi_n_1667, csa_tree_add_12_51_groupi_n_1668, csa_tree_add_12_51_groupi_n_1669, csa_tree_add_12_51_groupi_n_1670, csa_tree_add_12_51_groupi_n_1671, csa_tree_add_12_51_groupi_n_1672;
  wire csa_tree_add_12_51_groupi_n_1673, csa_tree_add_12_51_groupi_n_1674, csa_tree_add_12_51_groupi_n_1675, csa_tree_add_12_51_groupi_n_1676, csa_tree_add_12_51_groupi_n_1677, csa_tree_add_12_51_groupi_n_1678, csa_tree_add_12_51_groupi_n_1679, csa_tree_add_12_51_groupi_n_1680;
  wire csa_tree_add_12_51_groupi_n_1681, csa_tree_add_12_51_groupi_n_1682, csa_tree_add_12_51_groupi_n_1683, csa_tree_add_12_51_groupi_n_1684, csa_tree_add_12_51_groupi_n_1685, csa_tree_add_12_51_groupi_n_1686, csa_tree_add_12_51_groupi_n_1687, csa_tree_add_12_51_groupi_n_1688;
  wire csa_tree_add_12_51_groupi_n_1689, csa_tree_add_12_51_groupi_n_1690, csa_tree_add_12_51_groupi_n_1691, csa_tree_add_12_51_groupi_n_1692, csa_tree_add_12_51_groupi_n_1693, csa_tree_add_12_51_groupi_n_1694, csa_tree_add_12_51_groupi_n_1695, csa_tree_add_12_51_groupi_n_1696;
  wire csa_tree_add_12_51_groupi_n_1697, csa_tree_add_12_51_groupi_n_1698, csa_tree_add_12_51_groupi_n_1699, csa_tree_add_12_51_groupi_n_1700, csa_tree_add_12_51_groupi_n_1701, csa_tree_add_12_51_groupi_n_1702, csa_tree_add_12_51_groupi_n_1703, csa_tree_add_12_51_groupi_n_1704;
  wire csa_tree_add_12_51_groupi_n_1705, csa_tree_add_12_51_groupi_n_1706, csa_tree_add_12_51_groupi_n_1707, csa_tree_add_12_51_groupi_n_1708, csa_tree_add_12_51_groupi_n_1709, csa_tree_add_12_51_groupi_n_1710, csa_tree_add_12_51_groupi_n_1711, csa_tree_add_12_51_groupi_n_1712;
  wire csa_tree_add_12_51_groupi_n_1713, csa_tree_add_12_51_groupi_n_1714, csa_tree_add_12_51_groupi_n_1715, csa_tree_add_12_51_groupi_n_1716, csa_tree_add_12_51_groupi_n_1717, csa_tree_add_12_51_groupi_n_1718, csa_tree_add_12_51_groupi_n_1719, csa_tree_add_12_51_groupi_n_1720;
  wire csa_tree_add_12_51_groupi_n_1721, csa_tree_add_12_51_groupi_n_1722, csa_tree_add_12_51_groupi_n_1723, csa_tree_add_12_51_groupi_n_1724, csa_tree_add_12_51_groupi_n_1725, csa_tree_add_12_51_groupi_n_1726, csa_tree_add_12_51_groupi_n_1727, csa_tree_add_12_51_groupi_n_1728;
  wire csa_tree_add_12_51_groupi_n_1729, csa_tree_add_12_51_groupi_n_1730, csa_tree_add_12_51_groupi_n_1731, csa_tree_add_12_51_groupi_n_1732, csa_tree_add_12_51_groupi_n_1733, csa_tree_add_12_51_groupi_n_1734, csa_tree_add_12_51_groupi_n_1735, csa_tree_add_12_51_groupi_n_1736;
  wire csa_tree_add_12_51_groupi_n_1737, csa_tree_add_12_51_groupi_n_1738, csa_tree_add_12_51_groupi_n_1739, csa_tree_add_12_51_groupi_n_1740, csa_tree_add_12_51_groupi_n_1741, csa_tree_add_12_51_groupi_n_1742, csa_tree_add_12_51_groupi_n_1743, csa_tree_add_12_51_groupi_n_1744;
  wire csa_tree_add_12_51_groupi_n_1745, csa_tree_add_12_51_groupi_n_1746, csa_tree_add_12_51_groupi_n_1747, csa_tree_add_12_51_groupi_n_1748, csa_tree_add_12_51_groupi_n_1749, csa_tree_add_12_51_groupi_n_1750, csa_tree_add_12_51_groupi_n_1751, csa_tree_add_12_51_groupi_n_1752;
  wire csa_tree_add_12_51_groupi_n_1753, csa_tree_add_12_51_groupi_n_1754, csa_tree_add_12_51_groupi_n_1755, csa_tree_add_12_51_groupi_n_1756, csa_tree_add_12_51_groupi_n_1757, csa_tree_add_12_51_groupi_n_1758, csa_tree_add_12_51_groupi_n_1759, csa_tree_add_12_51_groupi_n_1760;
  wire csa_tree_add_12_51_groupi_n_1761, csa_tree_add_12_51_groupi_n_1762, csa_tree_add_12_51_groupi_n_1763, csa_tree_add_12_51_groupi_n_1764, csa_tree_add_12_51_groupi_n_1765, csa_tree_add_12_51_groupi_n_1766, csa_tree_add_12_51_groupi_n_1767, csa_tree_add_12_51_groupi_n_1768;
  wire csa_tree_add_12_51_groupi_n_1769, csa_tree_add_12_51_groupi_n_1770, csa_tree_add_12_51_groupi_n_1771, csa_tree_add_12_51_groupi_n_1772, csa_tree_add_12_51_groupi_n_1773, csa_tree_add_12_51_groupi_n_1774, csa_tree_add_12_51_groupi_n_1775, csa_tree_add_12_51_groupi_n_1776;
  wire csa_tree_add_12_51_groupi_n_1777, csa_tree_add_12_51_groupi_n_1778, csa_tree_add_12_51_groupi_n_1779, csa_tree_add_12_51_groupi_n_1780, csa_tree_add_12_51_groupi_n_1781, csa_tree_add_12_51_groupi_n_1782, csa_tree_add_12_51_groupi_n_1783, csa_tree_add_12_51_groupi_n_1784;
  wire csa_tree_add_12_51_groupi_n_1785, csa_tree_add_12_51_groupi_n_1786, csa_tree_add_12_51_groupi_n_1787, csa_tree_add_12_51_groupi_n_1788, csa_tree_add_12_51_groupi_n_1789, csa_tree_add_12_51_groupi_n_1790, csa_tree_add_12_51_groupi_n_1791, csa_tree_add_12_51_groupi_n_1792;
  wire csa_tree_add_12_51_groupi_n_1793, csa_tree_add_12_51_groupi_n_1794, csa_tree_add_12_51_groupi_n_1795, csa_tree_add_12_51_groupi_n_1796, csa_tree_add_12_51_groupi_n_1797, csa_tree_add_12_51_groupi_n_1798, csa_tree_add_12_51_groupi_n_1799, csa_tree_add_12_51_groupi_n_1800;
  wire csa_tree_add_12_51_groupi_n_1801, csa_tree_add_12_51_groupi_n_1802, csa_tree_add_12_51_groupi_n_1803, csa_tree_add_12_51_groupi_n_1804, csa_tree_add_12_51_groupi_n_1805, csa_tree_add_12_51_groupi_n_1806, csa_tree_add_12_51_groupi_n_1807, csa_tree_add_12_51_groupi_n_1808;
  wire csa_tree_add_12_51_groupi_n_1809, csa_tree_add_12_51_groupi_n_1810, csa_tree_add_12_51_groupi_n_1811, csa_tree_add_12_51_groupi_n_1812, csa_tree_add_12_51_groupi_n_1813, csa_tree_add_12_51_groupi_n_1814, csa_tree_add_12_51_groupi_n_1815, csa_tree_add_12_51_groupi_n_1816;
  wire csa_tree_add_12_51_groupi_n_1817, csa_tree_add_12_51_groupi_n_1818, csa_tree_add_12_51_groupi_n_1819, csa_tree_add_12_51_groupi_n_1820, csa_tree_add_12_51_groupi_n_1821, csa_tree_add_12_51_groupi_n_1822, csa_tree_add_12_51_groupi_n_1823, csa_tree_add_12_51_groupi_n_1824;
  wire csa_tree_add_12_51_groupi_n_1825, csa_tree_add_12_51_groupi_n_1826, csa_tree_add_12_51_groupi_n_1827, csa_tree_add_12_51_groupi_n_1828, csa_tree_add_12_51_groupi_n_1829, csa_tree_add_12_51_groupi_n_1830, csa_tree_add_12_51_groupi_n_1831, csa_tree_add_12_51_groupi_n_1832;
  wire csa_tree_add_12_51_groupi_n_1833, csa_tree_add_12_51_groupi_n_1834, csa_tree_add_12_51_groupi_n_1835, csa_tree_add_12_51_groupi_n_1836, csa_tree_add_12_51_groupi_n_1837, csa_tree_add_12_51_groupi_n_1838, csa_tree_add_12_51_groupi_n_1839, csa_tree_add_12_51_groupi_n_1840;
  wire csa_tree_add_12_51_groupi_n_1841, csa_tree_add_12_51_groupi_n_1842, csa_tree_add_12_51_groupi_n_1843, csa_tree_add_12_51_groupi_n_1844, csa_tree_add_12_51_groupi_n_1845, csa_tree_add_12_51_groupi_n_1846, csa_tree_add_12_51_groupi_n_1847, csa_tree_add_12_51_groupi_n_1848;
  wire csa_tree_add_12_51_groupi_n_1849, csa_tree_add_12_51_groupi_n_1850, csa_tree_add_12_51_groupi_n_1851, csa_tree_add_12_51_groupi_n_1852, csa_tree_add_12_51_groupi_n_1853, csa_tree_add_12_51_groupi_n_1854, csa_tree_add_12_51_groupi_n_1855, csa_tree_add_12_51_groupi_n_1856;
  wire csa_tree_add_12_51_groupi_n_1857, csa_tree_add_12_51_groupi_n_1858, csa_tree_add_12_51_groupi_n_1859, csa_tree_add_12_51_groupi_n_1860, csa_tree_add_12_51_groupi_n_1861, csa_tree_add_12_51_groupi_n_1862, csa_tree_add_12_51_groupi_n_1863, csa_tree_add_12_51_groupi_n_1864;
  wire csa_tree_add_12_51_groupi_n_1865, csa_tree_add_12_51_groupi_n_1866, csa_tree_add_12_51_groupi_n_1867, csa_tree_add_12_51_groupi_n_1868, csa_tree_add_12_51_groupi_n_1869, csa_tree_add_12_51_groupi_n_1870, csa_tree_add_12_51_groupi_n_1871, csa_tree_add_12_51_groupi_n_1872;
  wire csa_tree_add_12_51_groupi_n_1873, csa_tree_add_12_51_groupi_n_1874, csa_tree_add_12_51_groupi_n_1875, csa_tree_add_12_51_groupi_n_1876, csa_tree_add_12_51_groupi_n_1877, csa_tree_add_12_51_groupi_n_1878, csa_tree_add_12_51_groupi_n_1879, csa_tree_add_12_51_groupi_n_1880;
  wire csa_tree_add_12_51_groupi_n_1881, csa_tree_add_12_51_groupi_n_1882, csa_tree_add_12_51_groupi_n_1883, csa_tree_add_12_51_groupi_n_1884, csa_tree_add_12_51_groupi_n_1885, csa_tree_add_12_51_groupi_n_1886, csa_tree_add_12_51_groupi_n_1887, csa_tree_add_12_51_groupi_n_1888;
  wire csa_tree_add_12_51_groupi_n_1889, csa_tree_add_12_51_groupi_n_1890, csa_tree_add_12_51_groupi_n_1891, csa_tree_add_12_51_groupi_n_1892, csa_tree_add_12_51_groupi_n_1893, csa_tree_add_12_51_groupi_n_1894, csa_tree_add_12_51_groupi_n_1895, csa_tree_add_12_51_groupi_n_1896;
  wire csa_tree_add_12_51_groupi_n_1897, csa_tree_add_12_51_groupi_n_1898, csa_tree_add_12_51_groupi_n_1899, csa_tree_add_12_51_groupi_n_1900, csa_tree_add_12_51_groupi_n_1901, csa_tree_add_12_51_groupi_n_1902, csa_tree_add_12_51_groupi_n_1903, csa_tree_add_12_51_groupi_n_1904;
  wire csa_tree_add_12_51_groupi_n_1905, csa_tree_add_12_51_groupi_n_1906, csa_tree_add_12_51_groupi_n_1907, csa_tree_add_12_51_groupi_n_1908, csa_tree_add_12_51_groupi_n_1909, csa_tree_add_12_51_groupi_n_1910, csa_tree_add_12_51_groupi_n_1911, csa_tree_add_12_51_groupi_n_1912;
  wire csa_tree_add_12_51_groupi_n_1913, csa_tree_add_12_51_groupi_n_1914, csa_tree_add_12_51_groupi_n_1915, csa_tree_add_12_51_groupi_n_1916, csa_tree_add_12_51_groupi_n_1917, csa_tree_add_12_51_groupi_n_1918, csa_tree_add_12_51_groupi_n_1919, csa_tree_add_12_51_groupi_n_1920;
  wire csa_tree_add_12_51_groupi_n_1921, csa_tree_add_12_51_groupi_n_1922, csa_tree_add_12_51_groupi_n_1923, csa_tree_add_12_51_groupi_n_1924, csa_tree_add_12_51_groupi_n_1925, csa_tree_add_12_51_groupi_n_1926, csa_tree_add_12_51_groupi_n_1927, csa_tree_add_12_51_groupi_n_1928;
  wire csa_tree_add_12_51_groupi_n_1929, csa_tree_add_12_51_groupi_n_1930, csa_tree_add_12_51_groupi_n_1931, csa_tree_add_12_51_groupi_n_1932, csa_tree_add_12_51_groupi_n_1933, csa_tree_add_12_51_groupi_n_1934, csa_tree_add_12_51_groupi_n_1935, csa_tree_add_12_51_groupi_n_1936;
  wire csa_tree_add_12_51_groupi_n_1937, csa_tree_add_12_51_groupi_n_1938, csa_tree_add_12_51_groupi_n_1939, csa_tree_add_12_51_groupi_n_1940, csa_tree_add_12_51_groupi_n_1941, csa_tree_add_12_51_groupi_n_1942, csa_tree_add_12_51_groupi_n_1943, csa_tree_add_12_51_groupi_n_1944;
  wire csa_tree_add_12_51_groupi_n_1945, csa_tree_add_12_51_groupi_n_1946, csa_tree_add_12_51_groupi_n_1947, csa_tree_add_12_51_groupi_n_1948, csa_tree_add_12_51_groupi_n_1949, csa_tree_add_12_51_groupi_n_1950, csa_tree_add_12_51_groupi_n_1951, csa_tree_add_12_51_groupi_n_1952;
  wire csa_tree_add_12_51_groupi_n_1953, csa_tree_add_12_51_groupi_n_1954, csa_tree_add_12_51_groupi_n_1955, csa_tree_add_12_51_groupi_n_1956, csa_tree_add_12_51_groupi_n_1957, csa_tree_add_12_51_groupi_n_1958, csa_tree_add_12_51_groupi_n_1959, csa_tree_add_12_51_groupi_n_1960;
  wire csa_tree_add_12_51_groupi_n_1961, csa_tree_add_12_51_groupi_n_1962, csa_tree_add_12_51_groupi_n_1963, csa_tree_add_12_51_groupi_n_1964, csa_tree_add_12_51_groupi_n_1965, csa_tree_add_12_51_groupi_n_1966, csa_tree_add_12_51_groupi_n_1967, csa_tree_add_12_51_groupi_n_1968;
  wire csa_tree_add_12_51_groupi_n_1969, csa_tree_add_12_51_groupi_n_1970, csa_tree_add_12_51_groupi_n_1971, csa_tree_add_12_51_groupi_n_1972, csa_tree_add_12_51_groupi_n_1973, csa_tree_add_12_51_groupi_n_1974, csa_tree_add_12_51_groupi_n_1975, csa_tree_add_12_51_groupi_n_1976;
  wire csa_tree_add_12_51_groupi_n_1977, csa_tree_add_12_51_groupi_n_1978, csa_tree_add_12_51_groupi_n_1979, csa_tree_add_12_51_groupi_n_1980, csa_tree_add_12_51_groupi_n_1981, csa_tree_add_12_51_groupi_n_1982, csa_tree_add_12_51_groupi_n_1983, csa_tree_add_12_51_groupi_n_1984;
  wire csa_tree_add_12_51_groupi_n_1985, csa_tree_add_12_51_groupi_n_1986, csa_tree_add_12_51_groupi_n_1987, csa_tree_add_12_51_groupi_n_1988, csa_tree_add_12_51_groupi_n_1989, csa_tree_add_12_51_groupi_n_1990, csa_tree_add_12_51_groupi_n_1991, csa_tree_add_12_51_groupi_n_1992;
  wire csa_tree_add_12_51_groupi_n_1993, csa_tree_add_12_51_groupi_n_1994, csa_tree_add_12_51_groupi_n_1995, csa_tree_add_12_51_groupi_n_1996, csa_tree_add_12_51_groupi_n_1997, csa_tree_add_12_51_groupi_n_1998, csa_tree_add_12_51_groupi_n_1999, csa_tree_add_12_51_groupi_n_2000;
  wire csa_tree_add_12_51_groupi_n_2001, csa_tree_add_12_51_groupi_n_2002, csa_tree_add_12_51_groupi_n_2003, csa_tree_add_12_51_groupi_n_2004, csa_tree_add_12_51_groupi_n_2005, csa_tree_add_12_51_groupi_n_2006, csa_tree_add_12_51_groupi_n_2007, csa_tree_add_12_51_groupi_n_2008;
  wire csa_tree_add_12_51_groupi_n_2009, csa_tree_add_12_51_groupi_n_2010, csa_tree_add_12_51_groupi_n_2011, csa_tree_add_12_51_groupi_n_2012, csa_tree_add_12_51_groupi_n_2013, csa_tree_add_12_51_groupi_n_2014, csa_tree_add_12_51_groupi_n_2015, csa_tree_add_12_51_groupi_n_2016;
  wire csa_tree_add_12_51_groupi_n_2017, csa_tree_add_12_51_groupi_n_2018, csa_tree_add_12_51_groupi_n_2019, csa_tree_add_12_51_groupi_n_2020, csa_tree_add_12_51_groupi_n_2021, csa_tree_add_12_51_groupi_n_2022, csa_tree_add_12_51_groupi_n_2023, csa_tree_add_12_51_groupi_n_2024;
  wire csa_tree_add_12_51_groupi_n_2025, csa_tree_add_12_51_groupi_n_2026, csa_tree_add_12_51_groupi_n_2027, csa_tree_add_12_51_groupi_n_2028, csa_tree_add_12_51_groupi_n_2029, csa_tree_add_12_51_groupi_n_2030, csa_tree_add_12_51_groupi_n_2031, csa_tree_add_12_51_groupi_n_2032;
  wire csa_tree_add_12_51_groupi_n_2033, csa_tree_add_12_51_groupi_n_2034, csa_tree_add_12_51_groupi_n_2035, csa_tree_add_12_51_groupi_n_2036, csa_tree_add_12_51_groupi_n_2037, csa_tree_add_12_51_groupi_n_2038, csa_tree_add_12_51_groupi_n_2039, csa_tree_add_12_51_groupi_n_2040;
  wire csa_tree_add_12_51_groupi_n_2041, csa_tree_add_12_51_groupi_n_2042, csa_tree_add_12_51_groupi_n_2043, csa_tree_add_12_51_groupi_n_2044, csa_tree_add_12_51_groupi_n_2045, csa_tree_add_12_51_groupi_n_2046, csa_tree_add_12_51_groupi_n_2047, csa_tree_add_12_51_groupi_n_2048;
  wire csa_tree_add_12_51_groupi_n_2049, csa_tree_add_12_51_groupi_n_2050, csa_tree_add_12_51_groupi_n_2051, csa_tree_add_12_51_groupi_n_2052, csa_tree_add_12_51_groupi_n_2053, csa_tree_add_12_51_groupi_n_2054, csa_tree_add_12_51_groupi_n_2055, csa_tree_add_12_51_groupi_n_2056;
  wire csa_tree_add_12_51_groupi_n_2057, csa_tree_add_12_51_groupi_n_2058, csa_tree_add_12_51_groupi_n_2059, csa_tree_add_12_51_groupi_n_2060, csa_tree_add_12_51_groupi_n_2061, csa_tree_add_12_51_groupi_n_2062, csa_tree_add_12_51_groupi_n_2063, csa_tree_add_12_51_groupi_n_2064;
  wire csa_tree_add_12_51_groupi_n_2065, csa_tree_add_12_51_groupi_n_2066, csa_tree_add_12_51_groupi_n_2067, csa_tree_add_12_51_groupi_n_2068, csa_tree_add_12_51_groupi_n_2069, csa_tree_add_12_51_groupi_n_2070, csa_tree_add_12_51_groupi_n_2071, csa_tree_add_12_51_groupi_n_2072;
  wire csa_tree_add_12_51_groupi_n_2073, csa_tree_add_12_51_groupi_n_2074, csa_tree_add_12_51_groupi_n_2075, csa_tree_add_12_51_groupi_n_2076, csa_tree_add_12_51_groupi_n_2077, csa_tree_add_12_51_groupi_n_2078, csa_tree_add_12_51_groupi_n_2079, csa_tree_add_12_51_groupi_n_2080;
  wire csa_tree_add_12_51_groupi_n_2081, csa_tree_add_12_51_groupi_n_2082, csa_tree_add_12_51_groupi_n_2083, csa_tree_add_12_51_groupi_n_2084, csa_tree_add_12_51_groupi_n_2085, csa_tree_add_12_51_groupi_n_2086, csa_tree_add_12_51_groupi_n_2087, csa_tree_add_12_51_groupi_n_2088;
  wire csa_tree_add_12_51_groupi_n_2089, csa_tree_add_12_51_groupi_n_2090, csa_tree_add_12_51_groupi_n_2091, csa_tree_add_12_51_groupi_n_2092, csa_tree_add_12_51_groupi_n_2093, csa_tree_add_12_51_groupi_n_2094, csa_tree_add_12_51_groupi_n_2095, csa_tree_add_12_51_groupi_n_2096;
  wire csa_tree_add_12_51_groupi_n_2097, csa_tree_add_12_51_groupi_n_2098, csa_tree_add_12_51_groupi_n_2099, csa_tree_add_12_51_groupi_n_2100, csa_tree_add_12_51_groupi_n_2101, csa_tree_add_12_51_groupi_n_2102, csa_tree_add_12_51_groupi_n_2103, csa_tree_add_12_51_groupi_n_2104;
  wire csa_tree_add_12_51_groupi_n_2105, csa_tree_add_12_51_groupi_n_2106, csa_tree_add_12_51_groupi_n_2107, csa_tree_add_12_51_groupi_n_2108, csa_tree_add_12_51_groupi_n_2109, csa_tree_add_12_51_groupi_n_2110, csa_tree_add_12_51_groupi_n_2111, csa_tree_add_12_51_groupi_n_2112;
  wire csa_tree_add_12_51_groupi_n_2113, csa_tree_add_12_51_groupi_n_2114, csa_tree_add_12_51_groupi_n_2115, csa_tree_add_12_51_groupi_n_2116, csa_tree_add_12_51_groupi_n_2117, csa_tree_add_12_51_groupi_n_2118, csa_tree_add_12_51_groupi_n_2119, csa_tree_add_12_51_groupi_n_2120;
  wire csa_tree_add_12_51_groupi_n_2121, csa_tree_add_12_51_groupi_n_2122, csa_tree_add_12_51_groupi_n_2123, csa_tree_add_12_51_groupi_n_2124, csa_tree_add_12_51_groupi_n_2125, csa_tree_add_12_51_groupi_n_2126, csa_tree_add_12_51_groupi_n_2127, csa_tree_add_12_51_groupi_n_2128;
  wire csa_tree_add_12_51_groupi_n_2129, csa_tree_add_12_51_groupi_n_2130, csa_tree_add_12_51_groupi_n_2131, csa_tree_add_12_51_groupi_n_2132, csa_tree_add_12_51_groupi_n_2133, csa_tree_add_12_51_groupi_n_2134, csa_tree_add_12_51_groupi_n_2135, csa_tree_add_12_51_groupi_n_2136;
  wire csa_tree_add_12_51_groupi_n_2137, csa_tree_add_12_51_groupi_n_2138, csa_tree_add_12_51_groupi_n_2139, csa_tree_add_12_51_groupi_n_2140, csa_tree_add_12_51_groupi_n_2141, csa_tree_add_12_51_groupi_n_2142, csa_tree_add_12_51_groupi_n_2143, csa_tree_add_12_51_groupi_n_2144;
  wire csa_tree_add_12_51_groupi_n_2145, csa_tree_add_12_51_groupi_n_2146, csa_tree_add_12_51_groupi_n_2147, csa_tree_add_12_51_groupi_n_2148, csa_tree_add_12_51_groupi_n_2149, csa_tree_add_12_51_groupi_n_2150, csa_tree_add_12_51_groupi_n_2151, csa_tree_add_12_51_groupi_n_2152;
  wire csa_tree_add_12_51_groupi_n_2153, csa_tree_add_12_51_groupi_n_2154, csa_tree_add_12_51_groupi_n_2155, csa_tree_add_12_51_groupi_n_2156, csa_tree_add_12_51_groupi_n_2157, csa_tree_add_12_51_groupi_n_2158, csa_tree_add_12_51_groupi_n_2159, csa_tree_add_12_51_groupi_n_2160;
  wire csa_tree_add_12_51_groupi_n_2161, csa_tree_add_12_51_groupi_n_2162, csa_tree_add_12_51_groupi_n_2163, csa_tree_add_12_51_groupi_n_2164, csa_tree_add_12_51_groupi_n_2165, csa_tree_add_12_51_groupi_n_2166, csa_tree_add_12_51_groupi_n_2167, csa_tree_add_12_51_groupi_n_2168;
  wire csa_tree_add_12_51_groupi_n_2169, csa_tree_add_12_51_groupi_n_2170, csa_tree_add_12_51_groupi_n_2171, csa_tree_add_12_51_groupi_n_2172, csa_tree_add_12_51_groupi_n_2173, csa_tree_add_12_51_groupi_n_2174, csa_tree_add_12_51_groupi_n_2175, csa_tree_add_12_51_groupi_n_2176;
  wire csa_tree_add_12_51_groupi_n_2177, csa_tree_add_12_51_groupi_n_2178, csa_tree_add_12_51_groupi_n_2179, csa_tree_add_12_51_groupi_n_2180, csa_tree_add_12_51_groupi_n_2181, csa_tree_add_12_51_groupi_n_2182, csa_tree_add_12_51_groupi_n_2183, csa_tree_add_12_51_groupi_n_2184;
  wire csa_tree_add_12_51_groupi_n_2185, csa_tree_add_12_51_groupi_n_2186, csa_tree_add_12_51_groupi_n_2187, csa_tree_add_12_51_groupi_n_2188, csa_tree_add_12_51_groupi_n_2189, csa_tree_add_12_51_groupi_n_2190, csa_tree_add_12_51_groupi_n_2191, csa_tree_add_12_51_groupi_n_2192;
  wire csa_tree_add_12_51_groupi_n_2193, csa_tree_add_12_51_groupi_n_2194, csa_tree_add_12_51_groupi_n_2195, csa_tree_add_12_51_groupi_n_2196, csa_tree_add_12_51_groupi_n_2197, csa_tree_add_12_51_groupi_n_2198, csa_tree_add_12_51_groupi_n_2199, csa_tree_add_12_51_groupi_n_2200;
  wire csa_tree_add_12_51_groupi_n_2201, csa_tree_add_12_51_groupi_n_2202, csa_tree_add_12_51_groupi_n_2203, csa_tree_add_12_51_groupi_n_2204, csa_tree_add_12_51_groupi_n_2205, csa_tree_add_12_51_groupi_n_2206, csa_tree_add_12_51_groupi_n_2207, csa_tree_add_12_51_groupi_n_2208;
  wire csa_tree_add_12_51_groupi_n_2209, csa_tree_add_12_51_groupi_n_2210, csa_tree_add_12_51_groupi_n_2211, csa_tree_add_12_51_groupi_n_2212, csa_tree_add_12_51_groupi_n_2213, csa_tree_add_12_51_groupi_n_2214, csa_tree_add_12_51_groupi_n_2215, csa_tree_add_12_51_groupi_n_2216;
  wire csa_tree_add_12_51_groupi_n_2217, csa_tree_add_12_51_groupi_n_2218, csa_tree_add_12_51_groupi_n_2219, csa_tree_add_12_51_groupi_n_2220, csa_tree_add_12_51_groupi_n_2221, csa_tree_add_12_51_groupi_n_2222, csa_tree_add_12_51_groupi_n_2223, csa_tree_add_12_51_groupi_n_2224;
  wire csa_tree_add_12_51_groupi_n_2225, csa_tree_add_12_51_groupi_n_2226, csa_tree_add_12_51_groupi_n_2227, csa_tree_add_12_51_groupi_n_2228, csa_tree_add_12_51_groupi_n_2229, csa_tree_add_12_51_groupi_n_2230, csa_tree_add_12_51_groupi_n_2231, csa_tree_add_12_51_groupi_n_2232;
  wire csa_tree_add_12_51_groupi_n_2233, csa_tree_add_12_51_groupi_n_2234, csa_tree_add_12_51_groupi_n_2235, csa_tree_add_12_51_groupi_n_2236, csa_tree_add_12_51_groupi_n_2237, csa_tree_add_12_51_groupi_n_2238, csa_tree_add_12_51_groupi_n_2239, csa_tree_add_12_51_groupi_n_2240;
  wire csa_tree_add_12_51_groupi_n_2241, csa_tree_add_12_51_groupi_n_2242, csa_tree_add_12_51_groupi_n_2243, csa_tree_add_12_51_groupi_n_2244, csa_tree_add_12_51_groupi_n_2245, csa_tree_add_12_51_groupi_n_2246, csa_tree_add_12_51_groupi_n_2247, csa_tree_add_12_51_groupi_n_2248;
  wire csa_tree_add_12_51_groupi_n_2249, csa_tree_add_12_51_groupi_n_2250, csa_tree_add_12_51_groupi_n_2251, csa_tree_add_12_51_groupi_n_2252, csa_tree_add_12_51_groupi_n_2253, csa_tree_add_12_51_groupi_n_2254, csa_tree_add_12_51_groupi_n_2255, csa_tree_add_12_51_groupi_n_2256;
  wire csa_tree_add_12_51_groupi_n_2257, csa_tree_add_12_51_groupi_n_2258, csa_tree_add_12_51_groupi_n_2259, csa_tree_add_12_51_groupi_n_2260, csa_tree_add_12_51_groupi_n_2261, csa_tree_add_12_51_groupi_n_2262, csa_tree_add_12_51_groupi_n_2263, csa_tree_add_12_51_groupi_n_2264;
  wire csa_tree_add_12_51_groupi_n_2265, csa_tree_add_12_51_groupi_n_2266, csa_tree_add_12_51_groupi_n_2267, csa_tree_add_12_51_groupi_n_2268, csa_tree_add_12_51_groupi_n_2269, csa_tree_add_12_51_groupi_n_2270, csa_tree_add_12_51_groupi_n_2271, csa_tree_add_12_51_groupi_n_2272;
  wire csa_tree_add_12_51_groupi_n_2273, csa_tree_add_12_51_groupi_n_2274, csa_tree_add_12_51_groupi_n_2275, csa_tree_add_12_51_groupi_n_2276, csa_tree_add_12_51_groupi_n_2277, csa_tree_add_12_51_groupi_n_2278, csa_tree_add_12_51_groupi_n_2279, csa_tree_add_12_51_groupi_n_2280;
  wire csa_tree_add_12_51_groupi_n_2281, csa_tree_add_12_51_groupi_n_2282, csa_tree_add_12_51_groupi_n_2283, csa_tree_add_12_51_groupi_n_2284, csa_tree_add_12_51_groupi_n_2285, csa_tree_add_12_51_groupi_n_2286, csa_tree_add_12_51_groupi_n_2287, csa_tree_add_12_51_groupi_n_2288;
  wire csa_tree_add_12_51_groupi_n_2289, csa_tree_add_12_51_groupi_n_2290, csa_tree_add_12_51_groupi_n_2291, csa_tree_add_12_51_groupi_n_2292, csa_tree_add_12_51_groupi_n_2293, csa_tree_add_12_51_groupi_n_2294, csa_tree_add_12_51_groupi_n_2295, csa_tree_add_12_51_groupi_n_2296;
  wire csa_tree_add_12_51_groupi_n_2297, csa_tree_add_12_51_groupi_n_2298, csa_tree_add_12_51_groupi_n_2299, csa_tree_add_12_51_groupi_n_2300, csa_tree_add_12_51_groupi_n_2301, csa_tree_add_12_51_groupi_n_2302, csa_tree_add_12_51_groupi_n_2303, csa_tree_add_12_51_groupi_n_2304;
  wire csa_tree_add_12_51_groupi_n_2305, csa_tree_add_12_51_groupi_n_2306, csa_tree_add_12_51_groupi_n_2307, csa_tree_add_12_51_groupi_n_2308, csa_tree_add_12_51_groupi_n_2309, csa_tree_add_12_51_groupi_n_2310, csa_tree_add_12_51_groupi_n_2311, csa_tree_add_12_51_groupi_n_2312;
  wire csa_tree_add_12_51_groupi_n_2313, csa_tree_add_12_51_groupi_n_2314, csa_tree_add_12_51_groupi_n_2315, csa_tree_add_12_51_groupi_n_2316, csa_tree_add_12_51_groupi_n_2317, csa_tree_add_12_51_groupi_n_2318, csa_tree_add_12_51_groupi_n_2319, csa_tree_add_12_51_groupi_n_2320;
  wire csa_tree_add_12_51_groupi_n_2321, csa_tree_add_12_51_groupi_n_2322, csa_tree_add_12_51_groupi_n_2323, csa_tree_add_12_51_groupi_n_2324, csa_tree_add_12_51_groupi_n_2325, csa_tree_add_12_51_groupi_n_2326, csa_tree_add_12_51_groupi_n_2327, csa_tree_add_12_51_groupi_n_2328;
  wire csa_tree_add_12_51_groupi_n_2329, csa_tree_add_12_51_groupi_n_2330, csa_tree_add_12_51_groupi_n_2331, csa_tree_add_12_51_groupi_n_2332, csa_tree_add_12_51_groupi_n_2333, csa_tree_add_12_51_groupi_n_2334, csa_tree_add_12_51_groupi_n_2335, csa_tree_add_12_51_groupi_n_2336;
  wire csa_tree_add_12_51_groupi_n_2337, csa_tree_add_12_51_groupi_n_2338, csa_tree_add_12_51_groupi_n_2339, csa_tree_add_12_51_groupi_n_2340, csa_tree_add_12_51_groupi_n_2341, csa_tree_add_12_51_groupi_n_2342, csa_tree_add_12_51_groupi_n_2343, csa_tree_add_12_51_groupi_n_2344;
  wire csa_tree_add_12_51_groupi_n_2345, csa_tree_add_12_51_groupi_n_2346, csa_tree_add_12_51_groupi_n_2347, csa_tree_add_12_51_groupi_n_2348, csa_tree_add_12_51_groupi_n_2349, csa_tree_add_12_51_groupi_n_2350, csa_tree_add_12_51_groupi_n_2351, csa_tree_add_12_51_groupi_n_2352;
  wire csa_tree_add_12_51_groupi_n_2353, csa_tree_add_12_51_groupi_n_2354, csa_tree_add_12_51_groupi_n_2355, csa_tree_add_12_51_groupi_n_2356, csa_tree_add_12_51_groupi_n_2357, csa_tree_add_12_51_groupi_n_2358, csa_tree_add_12_51_groupi_n_2359, csa_tree_add_12_51_groupi_n_2360;
  wire csa_tree_add_12_51_groupi_n_2361, csa_tree_add_12_51_groupi_n_2362, csa_tree_add_12_51_groupi_n_2363, csa_tree_add_12_51_groupi_n_2364, csa_tree_add_12_51_groupi_n_2365, csa_tree_add_12_51_groupi_n_2366, csa_tree_add_12_51_groupi_n_2367, csa_tree_add_12_51_groupi_n_2368;
  wire csa_tree_add_12_51_groupi_n_2369, csa_tree_add_12_51_groupi_n_2370, csa_tree_add_12_51_groupi_n_2371, csa_tree_add_12_51_groupi_n_2372, csa_tree_add_12_51_groupi_n_2373, csa_tree_add_12_51_groupi_n_2374, csa_tree_add_12_51_groupi_n_2375, csa_tree_add_12_51_groupi_n_2376;
  wire csa_tree_add_12_51_groupi_n_2377, csa_tree_add_12_51_groupi_n_2378, csa_tree_add_12_51_groupi_n_2379, csa_tree_add_12_51_groupi_n_2380, csa_tree_add_12_51_groupi_n_2381, csa_tree_add_12_51_groupi_n_2382, csa_tree_add_12_51_groupi_n_2383, csa_tree_add_12_51_groupi_n_2384;
  wire csa_tree_add_12_51_groupi_n_2385, csa_tree_add_12_51_groupi_n_2386, csa_tree_add_12_51_groupi_n_2387, csa_tree_add_12_51_groupi_n_2388, csa_tree_add_12_51_groupi_n_2389, csa_tree_add_12_51_groupi_n_2390, csa_tree_add_12_51_groupi_n_2391, csa_tree_add_12_51_groupi_n_2392;
  wire csa_tree_add_12_51_groupi_n_2393, csa_tree_add_12_51_groupi_n_2394, csa_tree_add_12_51_groupi_n_2395, csa_tree_add_12_51_groupi_n_2396, csa_tree_add_12_51_groupi_n_2397, csa_tree_add_12_51_groupi_n_2398, csa_tree_add_12_51_groupi_n_2399, csa_tree_add_12_51_groupi_n_2400;
  wire csa_tree_add_12_51_groupi_n_2401, csa_tree_add_12_51_groupi_n_2402, csa_tree_add_12_51_groupi_n_2403, csa_tree_add_12_51_groupi_n_2404, csa_tree_add_12_51_groupi_n_2405, csa_tree_add_12_51_groupi_n_2406, csa_tree_add_12_51_groupi_n_2407, csa_tree_add_12_51_groupi_n_2408;
  wire csa_tree_add_12_51_groupi_n_2409, csa_tree_add_12_51_groupi_n_2410, csa_tree_add_12_51_groupi_n_2411, csa_tree_add_12_51_groupi_n_2412, csa_tree_add_12_51_groupi_n_2413, csa_tree_add_12_51_groupi_n_2414, csa_tree_add_12_51_groupi_n_2415, csa_tree_add_12_51_groupi_n_2416;
  wire csa_tree_add_12_51_groupi_n_2417, csa_tree_add_12_51_groupi_n_2418, csa_tree_add_12_51_groupi_n_2419, csa_tree_add_12_51_groupi_n_2420, csa_tree_add_12_51_groupi_n_2421, csa_tree_add_12_51_groupi_n_2422, csa_tree_add_12_51_groupi_n_2423, csa_tree_add_12_51_groupi_n_2424;
  wire csa_tree_add_12_51_groupi_n_2425, csa_tree_add_12_51_groupi_n_2426, csa_tree_add_12_51_groupi_n_2427, csa_tree_add_12_51_groupi_n_2428, csa_tree_add_12_51_groupi_n_2429, csa_tree_add_12_51_groupi_n_2430, csa_tree_add_12_51_groupi_n_2431, csa_tree_add_12_51_groupi_n_2432;
  wire csa_tree_add_12_51_groupi_n_2433, csa_tree_add_12_51_groupi_n_2434, csa_tree_add_12_51_groupi_n_2435, csa_tree_add_12_51_groupi_n_2436, csa_tree_add_12_51_groupi_n_2437, csa_tree_add_12_51_groupi_n_2438, csa_tree_add_12_51_groupi_n_2439, csa_tree_add_12_51_groupi_n_2440;
  wire csa_tree_add_12_51_groupi_n_2441, csa_tree_add_12_51_groupi_n_2442, csa_tree_add_12_51_groupi_n_2443, csa_tree_add_12_51_groupi_n_2444, csa_tree_add_12_51_groupi_n_2445, csa_tree_add_12_51_groupi_n_2446, csa_tree_add_12_51_groupi_n_2447, csa_tree_add_12_51_groupi_n_2448;
  wire csa_tree_add_12_51_groupi_n_2449, csa_tree_add_12_51_groupi_n_2450, csa_tree_add_12_51_groupi_n_2451, csa_tree_add_12_51_groupi_n_2452, csa_tree_add_12_51_groupi_n_2453, csa_tree_add_12_51_groupi_n_2454, csa_tree_add_12_51_groupi_n_2455, csa_tree_add_12_51_groupi_n_2456;
  wire csa_tree_add_12_51_groupi_n_2457, csa_tree_add_12_51_groupi_n_2458, csa_tree_add_12_51_groupi_n_2459, csa_tree_add_12_51_groupi_n_2460, csa_tree_add_12_51_groupi_n_2461, csa_tree_add_12_51_groupi_n_2462, csa_tree_add_12_51_groupi_n_2463, csa_tree_add_12_51_groupi_n_2464;
  wire csa_tree_add_12_51_groupi_n_2465, csa_tree_add_12_51_groupi_n_2466, csa_tree_add_12_51_groupi_n_2467, csa_tree_add_12_51_groupi_n_2468, csa_tree_add_12_51_groupi_n_2469, csa_tree_add_12_51_groupi_n_2470, csa_tree_add_12_51_groupi_n_2471, csa_tree_add_12_51_groupi_n_2472;
  wire csa_tree_add_12_51_groupi_n_2473, csa_tree_add_12_51_groupi_n_2474, csa_tree_add_12_51_groupi_n_2475, csa_tree_add_12_51_groupi_n_2476, csa_tree_add_12_51_groupi_n_2477, csa_tree_add_12_51_groupi_n_2478, csa_tree_add_12_51_groupi_n_2479, csa_tree_add_12_51_groupi_n_2480;
  wire csa_tree_add_12_51_groupi_n_2481, csa_tree_add_12_51_groupi_n_2482, csa_tree_add_12_51_groupi_n_2483, csa_tree_add_12_51_groupi_n_2484, csa_tree_add_12_51_groupi_n_2485, csa_tree_add_12_51_groupi_n_2486, csa_tree_add_12_51_groupi_n_2487, csa_tree_add_12_51_groupi_n_2488;
  wire csa_tree_add_12_51_groupi_n_2489, csa_tree_add_12_51_groupi_n_2490, csa_tree_add_12_51_groupi_n_2491, csa_tree_add_12_51_groupi_n_2492, csa_tree_add_12_51_groupi_n_2493, csa_tree_add_12_51_groupi_n_2494, csa_tree_add_12_51_groupi_n_2495, csa_tree_add_12_51_groupi_n_2496;
  wire csa_tree_add_12_51_groupi_n_2497, csa_tree_add_12_51_groupi_n_2498, csa_tree_add_12_51_groupi_n_2499, csa_tree_add_12_51_groupi_n_2500, csa_tree_add_12_51_groupi_n_2501, csa_tree_add_12_51_groupi_n_2502, csa_tree_add_12_51_groupi_n_2503, csa_tree_add_12_51_groupi_n_2504;
  wire csa_tree_add_12_51_groupi_n_2505, csa_tree_add_12_51_groupi_n_2506, csa_tree_add_12_51_groupi_n_2507, csa_tree_add_12_51_groupi_n_2508, csa_tree_add_12_51_groupi_n_2509, csa_tree_add_12_51_groupi_n_2510, csa_tree_add_12_51_groupi_n_2511, csa_tree_add_12_51_groupi_n_2512;
  wire csa_tree_add_12_51_groupi_n_2513, csa_tree_add_12_51_groupi_n_2514, csa_tree_add_12_51_groupi_n_2515, csa_tree_add_12_51_groupi_n_2516, csa_tree_add_12_51_groupi_n_2517, csa_tree_add_12_51_groupi_n_2518, csa_tree_add_12_51_groupi_n_2519, csa_tree_add_12_51_groupi_n_2520;
  wire csa_tree_add_12_51_groupi_n_2521, csa_tree_add_12_51_groupi_n_2522, csa_tree_add_12_51_groupi_n_2523, csa_tree_add_12_51_groupi_n_2524, csa_tree_add_12_51_groupi_n_2525, csa_tree_add_12_51_groupi_n_2526, csa_tree_add_12_51_groupi_n_2527, csa_tree_add_12_51_groupi_n_2528;
  wire csa_tree_add_12_51_groupi_n_2529, csa_tree_add_12_51_groupi_n_2530, csa_tree_add_12_51_groupi_n_2531, csa_tree_add_12_51_groupi_n_2532, csa_tree_add_12_51_groupi_n_2533, csa_tree_add_12_51_groupi_n_2534, csa_tree_add_12_51_groupi_n_2535, csa_tree_add_12_51_groupi_n_2536;
  wire csa_tree_add_12_51_groupi_n_2537, csa_tree_add_12_51_groupi_n_2538, csa_tree_add_12_51_groupi_n_2539, csa_tree_add_12_51_groupi_n_2540, csa_tree_add_12_51_groupi_n_2541, csa_tree_add_12_51_groupi_n_2542, csa_tree_add_12_51_groupi_n_2543, csa_tree_add_12_51_groupi_n_2544;
  wire csa_tree_add_12_51_groupi_n_2545, csa_tree_add_12_51_groupi_n_2546, csa_tree_add_12_51_groupi_n_2547, csa_tree_add_12_51_groupi_n_2548, csa_tree_add_12_51_groupi_n_2549, csa_tree_add_12_51_groupi_n_2550, csa_tree_add_12_51_groupi_n_2551, csa_tree_add_12_51_groupi_n_2552;
  wire csa_tree_add_12_51_groupi_n_2553, csa_tree_add_12_51_groupi_n_2554, csa_tree_add_12_51_groupi_n_2555, csa_tree_add_12_51_groupi_n_2556, csa_tree_add_12_51_groupi_n_2557, csa_tree_add_12_51_groupi_n_2558, csa_tree_add_12_51_groupi_n_2559, csa_tree_add_12_51_groupi_n_2560;
  wire csa_tree_add_12_51_groupi_n_2561, csa_tree_add_12_51_groupi_n_2562, csa_tree_add_12_51_groupi_n_2563, csa_tree_add_12_51_groupi_n_2564, csa_tree_add_12_51_groupi_n_2565, csa_tree_add_12_51_groupi_n_2566, csa_tree_add_12_51_groupi_n_2567, csa_tree_add_12_51_groupi_n_2568;
  wire csa_tree_add_12_51_groupi_n_2569, csa_tree_add_12_51_groupi_n_2570, csa_tree_add_12_51_groupi_n_2571, csa_tree_add_12_51_groupi_n_2572, csa_tree_add_12_51_groupi_n_2573, csa_tree_add_12_51_groupi_n_2574, csa_tree_add_12_51_groupi_n_2575, csa_tree_add_12_51_groupi_n_2576;
  wire csa_tree_add_12_51_groupi_n_2577, csa_tree_add_12_51_groupi_n_2578, csa_tree_add_12_51_groupi_n_2579, csa_tree_add_12_51_groupi_n_2580, csa_tree_add_12_51_groupi_n_2581, csa_tree_add_12_51_groupi_n_2582, csa_tree_add_12_51_groupi_n_2583, csa_tree_add_12_51_groupi_n_2584;
  wire csa_tree_add_12_51_groupi_n_2585, csa_tree_add_12_51_groupi_n_2586, csa_tree_add_12_51_groupi_n_2587, csa_tree_add_12_51_groupi_n_2588, csa_tree_add_12_51_groupi_n_2589, csa_tree_add_12_51_groupi_n_2590, csa_tree_add_12_51_groupi_n_2591, csa_tree_add_12_51_groupi_n_2592;
  wire csa_tree_add_12_51_groupi_n_2593, csa_tree_add_12_51_groupi_n_2594, csa_tree_add_12_51_groupi_n_2595, csa_tree_add_12_51_groupi_n_2596, csa_tree_add_12_51_groupi_n_2597, csa_tree_add_12_51_groupi_n_2598, csa_tree_add_12_51_groupi_n_2599, csa_tree_add_12_51_groupi_n_2600;
  wire csa_tree_add_12_51_groupi_n_2601, csa_tree_add_12_51_groupi_n_2602, csa_tree_add_12_51_groupi_n_2603, csa_tree_add_12_51_groupi_n_2604, csa_tree_add_12_51_groupi_n_2605, csa_tree_add_12_51_groupi_n_2606, csa_tree_add_12_51_groupi_n_2607, csa_tree_add_12_51_groupi_n_2608;
  wire csa_tree_add_12_51_groupi_n_2609, csa_tree_add_12_51_groupi_n_2610, csa_tree_add_12_51_groupi_n_2611, csa_tree_add_12_51_groupi_n_2612, csa_tree_add_12_51_groupi_n_2613, csa_tree_add_12_51_groupi_n_2614, csa_tree_add_12_51_groupi_n_2615, csa_tree_add_12_51_groupi_n_2616;
  wire csa_tree_add_12_51_groupi_n_2617, csa_tree_add_12_51_groupi_n_2618, csa_tree_add_12_51_groupi_n_2619, csa_tree_add_12_51_groupi_n_2620, csa_tree_add_12_51_groupi_n_2621, csa_tree_add_12_51_groupi_n_2622, csa_tree_add_12_51_groupi_n_2623, csa_tree_add_12_51_groupi_n_2624;
  wire csa_tree_add_12_51_groupi_n_2625, csa_tree_add_12_51_groupi_n_2626, csa_tree_add_12_51_groupi_n_2627, csa_tree_add_12_51_groupi_n_2628, csa_tree_add_12_51_groupi_n_2629, csa_tree_add_12_51_groupi_n_2630, csa_tree_add_12_51_groupi_n_2631, csa_tree_add_12_51_groupi_n_2632;
  wire csa_tree_add_12_51_groupi_n_2633, csa_tree_add_12_51_groupi_n_2634, csa_tree_add_12_51_groupi_n_2635, csa_tree_add_12_51_groupi_n_2636, csa_tree_add_12_51_groupi_n_2637, csa_tree_add_12_51_groupi_n_2638, csa_tree_add_12_51_groupi_n_2639, csa_tree_add_12_51_groupi_n_2640;
  wire csa_tree_add_12_51_groupi_n_2641, csa_tree_add_12_51_groupi_n_2642, csa_tree_add_12_51_groupi_n_2643, csa_tree_add_12_51_groupi_n_2644, csa_tree_add_12_51_groupi_n_2645, csa_tree_add_12_51_groupi_n_2646, csa_tree_add_12_51_groupi_n_2647, csa_tree_add_12_51_groupi_n_2648;
  wire csa_tree_add_12_51_groupi_n_2649, csa_tree_add_12_51_groupi_n_2650, csa_tree_add_12_51_groupi_n_2651, csa_tree_add_12_51_groupi_n_2652, csa_tree_add_12_51_groupi_n_2653, csa_tree_add_12_51_groupi_n_2654, csa_tree_add_12_51_groupi_n_2655, csa_tree_add_12_51_groupi_n_2656;
  wire csa_tree_add_12_51_groupi_n_2657, csa_tree_add_12_51_groupi_n_2658, csa_tree_add_12_51_groupi_n_2659, csa_tree_add_12_51_groupi_n_2660, csa_tree_add_12_51_groupi_n_2661, csa_tree_add_12_51_groupi_n_2662, csa_tree_add_12_51_groupi_n_2663, csa_tree_add_12_51_groupi_n_2664;
  wire csa_tree_add_12_51_groupi_n_2665, csa_tree_add_12_51_groupi_n_2666, csa_tree_add_12_51_groupi_n_2667, csa_tree_add_12_51_groupi_n_2668, csa_tree_add_12_51_groupi_n_2669, csa_tree_add_12_51_groupi_n_2670, csa_tree_add_12_51_groupi_n_2671, csa_tree_add_12_51_groupi_n_2672;
  wire csa_tree_add_12_51_groupi_n_2673, csa_tree_add_12_51_groupi_n_2674, csa_tree_add_12_51_groupi_n_2675, csa_tree_add_12_51_groupi_n_2676, csa_tree_add_12_51_groupi_n_2677, csa_tree_add_12_51_groupi_n_2678, csa_tree_add_12_51_groupi_n_2679, csa_tree_add_12_51_groupi_n_2680;
  wire csa_tree_add_12_51_groupi_n_2681, csa_tree_add_12_51_groupi_n_2682, csa_tree_add_12_51_groupi_n_2683, csa_tree_add_12_51_groupi_n_2684, csa_tree_add_12_51_groupi_n_2685, csa_tree_add_12_51_groupi_n_2686, csa_tree_add_12_51_groupi_n_2687, csa_tree_add_12_51_groupi_n_2688;
  wire csa_tree_add_12_51_groupi_n_2689, csa_tree_add_12_51_groupi_n_2690, csa_tree_add_12_51_groupi_n_2691, csa_tree_add_12_51_groupi_n_2692, csa_tree_add_12_51_groupi_n_2693, csa_tree_add_12_51_groupi_n_2694, csa_tree_add_12_51_groupi_n_2695, csa_tree_add_12_51_groupi_n_2696;
  wire csa_tree_add_12_51_groupi_n_2697, csa_tree_add_12_51_groupi_n_2698, csa_tree_add_12_51_groupi_n_2699, csa_tree_add_12_51_groupi_n_2700, csa_tree_add_12_51_groupi_n_2701, csa_tree_add_12_51_groupi_n_2702, csa_tree_add_12_51_groupi_n_2703, csa_tree_add_12_51_groupi_n_2704;
  wire csa_tree_add_12_51_groupi_n_2705, csa_tree_add_12_51_groupi_n_2706, csa_tree_add_12_51_groupi_n_2707, csa_tree_add_12_51_groupi_n_2708, csa_tree_add_12_51_groupi_n_2709, csa_tree_add_12_51_groupi_n_2710, csa_tree_add_12_51_groupi_n_2711, csa_tree_add_12_51_groupi_n_2712;
  wire csa_tree_add_12_51_groupi_n_2713, csa_tree_add_12_51_groupi_n_2714, csa_tree_add_12_51_groupi_n_2715, csa_tree_add_12_51_groupi_n_2716, csa_tree_add_12_51_groupi_n_2717, csa_tree_add_12_51_groupi_n_2718, csa_tree_add_12_51_groupi_n_2719, csa_tree_add_12_51_groupi_n_2720;
  wire csa_tree_add_12_51_groupi_n_2721, csa_tree_add_12_51_groupi_n_2722, csa_tree_add_12_51_groupi_n_2723, csa_tree_add_12_51_groupi_n_2724, csa_tree_add_12_51_groupi_n_2725, csa_tree_add_12_51_groupi_n_2726, csa_tree_add_12_51_groupi_n_2727, csa_tree_add_12_51_groupi_n_2728;
  wire csa_tree_add_12_51_groupi_n_2729, csa_tree_add_12_51_groupi_n_2730, csa_tree_add_12_51_groupi_n_2731, csa_tree_add_12_51_groupi_n_2732, csa_tree_add_12_51_groupi_n_2733, csa_tree_add_12_51_groupi_n_2734, csa_tree_add_12_51_groupi_n_2735, csa_tree_add_12_51_groupi_n_2736;
  wire csa_tree_add_12_51_groupi_n_2737, csa_tree_add_12_51_groupi_n_2738, csa_tree_add_12_51_groupi_n_2739, csa_tree_add_12_51_groupi_n_2740, csa_tree_add_12_51_groupi_n_2741, csa_tree_add_12_51_groupi_n_2742, csa_tree_add_12_51_groupi_n_2743, csa_tree_add_12_51_groupi_n_2744;
  wire csa_tree_add_12_51_groupi_n_2745, csa_tree_add_12_51_groupi_n_2746, csa_tree_add_12_51_groupi_n_2747, csa_tree_add_12_51_groupi_n_2748, csa_tree_add_12_51_groupi_n_2749, csa_tree_add_12_51_groupi_n_2750, csa_tree_add_12_51_groupi_n_2751, csa_tree_add_12_51_groupi_n_2752;
  wire csa_tree_add_12_51_groupi_n_2753, csa_tree_add_12_51_groupi_n_2754, csa_tree_add_12_51_groupi_n_2755, csa_tree_add_12_51_groupi_n_2756, csa_tree_add_12_51_groupi_n_2757, csa_tree_add_12_51_groupi_n_2758, csa_tree_add_12_51_groupi_n_2759, csa_tree_add_12_51_groupi_n_2760;
  wire csa_tree_add_12_51_groupi_n_2761, csa_tree_add_12_51_groupi_n_2762, csa_tree_add_12_51_groupi_n_2763, csa_tree_add_12_51_groupi_n_2764, csa_tree_add_12_51_groupi_n_2765, csa_tree_add_12_51_groupi_n_2766, csa_tree_add_12_51_groupi_n_2767, csa_tree_add_12_51_groupi_n_2768;
  wire csa_tree_add_12_51_groupi_n_2769, csa_tree_add_12_51_groupi_n_2770, csa_tree_add_12_51_groupi_n_2771, csa_tree_add_12_51_groupi_n_2772, csa_tree_add_12_51_groupi_n_2773, csa_tree_add_12_51_groupi_n_2774, csa_tree_add_12_51_groupi_n_2775, csa_tree_add_12_51_groupi_n_2776;
  wire csa_tree_add_12_51_groupi_n_2777, csa_tree_add_12_51_groupi_n_2778, csa_tree_add_12_51_groupi_n_2779, csa_tree_add_12_51_groupi_n_2780, csa_tree_add_12_51_groupi_n_2781, csa_tree_add_12_51_groupi_n_2782, csa_tree_add_12_51_groupi_n_2783, csa_tree_add_12_51_groupi_n_2784;
  wire csa_tree_add_12_51_groupi_n_2785, csa_tree_add_12_51_groupi_n_2786, csa_tree_add_12_51_groupi_n_2787, csa_tree_add_12_51_groupi_n_2788, csa_tree_add_12_51_groupi_n_2789, csa_tree_add_12_51_groupi_n_2790, csa_tree_add_12_51_groupi_n_2791, csa_tree_add_12_51_groupi_n_2792;
  wire csa_tree_add_12_51_groupi_n_2793, csa_tree_add_12_51_groupi_n_2794, csa_tree_add_12_51_groupi_n_2795, csa_tree_add_12_51_groupi_n_2796, csa_tree_add_12_51_groupi_n_2797, csa_tree_add_12_51_groupi_n_2798, csa_tree_add_12_51_groupi_n_2799, csa_tree_add_12_51_groupi_n_2800;
  wire csa_tree_add_12_51_groupi_n_2801, csa_tree_add_12_51_groupi_n_2802, csa_tree_add_12_51_groupi_n_2803, csa_tree_add_12_51_groupi_n_2804, csa_tree_add_12_51_groupi_n_2805, csa_tree_add_12_51_groupi_n_2806, csa_tree_add_12_51_groupi_n_2807, csa_tree_add_12_51_groupi_n_2808;
  wire csa_tree_add_12_51_groupi_n_2809, csa_tree_add_12_51_groupi_n_2810, csa_tree_add_12_51_groupi_n_2811, csa_tree_add_12_51_groupi_n_2812, csa_tree_add_12_51_groupi_n_2813, csa_tree_add_12_51_groupi_n_2814, csa_tree_add_12_51_groupi_n_2815, csa_tree_add_12_51_groupi_n_2816;
  wire csa_tree_add_12_51_groupi_n_2817, csa_tree_add_12_51_groupi_n_2818, csa_tree_add_12_51_groupi_n_2819, csa_tree_add_12_51_groupi_n_2820, csa_tree_add_12_51_groupi_n_2821, csa_tree_add_12_51_groupi_n_2822, csa_tree_add_12_51_groupi_n_2823, csa_tree_add_12_51_groupi_n_2824;
  wire csa_tree_add_12_51_groupi_n_2825, csa_tree_add_12_51_groupi_n_2826, csa_tree_add_12_51_groupi_n_2827, csa_tree_add_12_51_groupi_n_2828, csa_tree_add_12_51_groupi_n_2829, csa_tree_add_12_51_groupi_n_2830, csa_tree_add_12_51_groupi_n_2831, csa_tree_add_12_51_groupi_n_2832;
  wire csa_tree_add_12_51_groupi_n_2833, csa_tree_add_12_51_groupi_n_2834, csa_tree_add_12_51_groupi_n_2835, csa_tree_add_12_51_groupi_n_2836, csa_tree_add_12_51_groupi_n_2837, csa_tree_add_12_51_groupi_n_2838, csa_tree_add_12_51_groupi_n_2839, csa_tree_add_12_51_groupi_n_2840;
  wire csa_tree_add_12_51_groupi_n_2841, csa_tree_add_12_51_groupi_n_2842, csa_tree_add_12_51_groupi_n_2843, csa_tree_add_12_51_groupi_n_2844, csa_tree_add_12_51_groupi_n_2845, csa_tree_add_12_51_groupi_n_2846, csa_tree_add_12_51_groupi_n_2847, csa_tree_add_12_51_groupi_n_2848;
  wire csa_tree_add_12_51_groupi_n_2849, csa_tree_add_12_51_groupi_n_2850, csa_tree_add_12_51_groupi_n_2851, csa_tree_add_12_51_groupi_n_2852, csa_tree_add_12_51_groupi_n_2853, csa_tree_add_12_51_groupi_n_2854, csa_tree_add_12_51_groupi_n_2855, csa_tree_add_12_51_groupi_n_2856;
  wire csa_tree_add_12_51_groupi_n_2857, csa_tree_add_12_51_groupi_n_2858, csa_tree_add_12_51_groupi_n_2859, csa_tree_add_12_51_groupi_n_2860, csa_tree_add_12_51_groupi_n_2861, csa_tree_add_12_51_groupi_n_2862, csa_tree_add_12_51_groupi_n_2863, csa_tree_add_12_51_groupi_n_2864;
  wire csa_tree_add_12_51_groupi_n_2865, csa_tree_add_12_51_groupi_n_2866, csa_tree_add_12_51_groupi_n_2867, csa_tree_add_12_51_groupi_n_2868, csa_tree_add_12_51_groupi_n_2869, csa_tree_add_12_51_groupi_n_2870, csa_tree_add_12_51_groupi_n_2871, csa_tree_add_12_51_groupi_n_2872;
  wire csa_tree_add_12_51_groupi_n_2873, csa_tree_add_12_51_groupi_n_2874, csa_tree_add_12_51_groupi_n_2875, csa_tree_add_12_51_groupi_n_2876, csa_tree_add_12_51_groupi_n_2877, csa_tree_add_12_51_groupi_n_2878, csa_tree_add_12_51_groupi_n_2879, csa_tree_add_12_51_groupi_n_2880;
  wire csa_tree_add_12_51_groupi_n_2881, csa_tree_add_12_51_groupi_n_2882, csa_tree_add_12_51_groupi_n_2883, csa_tree_add_12_51_groupi_n_2884, csa_tree_add_12_51_groupi_n_2885, csa_tree_add_12_51_groupi_n_2886, csa_tree_add_12_51_groupi_n_2887, csa_tree_add_12_51_groupi_n_2888;
  wire csa_tree_add_12_51_groupi_n_2889, csa_tree_add_12_51_groupi_n_2890, csa_tree_add_12_51_groupi_n_2891, csa_tree_add_12_51_groupi_n_2892, csa_tree_add_12_51_groupi_n_2893, csa_tree_add_12_51_groupi_n_2894, csa_tree_add_12_51_groupi_n_2895, csa_tree_add_12_51_groupi_n_2896;
  wire csa_tree_add_12_51_groupi_n_2897, csa_tree_add_12_51_groupi_n_2898, csa_tree_add_12_51_groupi_n_2899, csa_tree_add_12_51_groupi_n_2900, csa_tree_add_12_51_groupi_n_2901, csa_tree_add_12_51_groupi_n_2902, csa_tree_add_12_51_groupi_n_2903, csa_tree_add_12_51_groupi_n_2904;
  wire csa_tree_add_12_51_groupi_n_2905, csa_tree_add_12_51_groupi_n_2906, csa_tree_add_12_51_groupi_n_2907, csa_tree_add_12_51_groupi_n_2908, csa_tree_add_12_51_groupi_n_2909, csa_tree_add_12_51_groupi_n_2910, csa_tree_add_12_51_groupi_n_2911, csa_tree_add_12_51_groupi_n_2912;
  wire csa_tree_add_12_51_groupi_n_2913, csa_tree_add_12_51_groupi_n_2914, csa_tree_add_12_51_groupi_n_2915, csa_tree_add_12_51_groupi_n_2916, csa_tree_add_12_51_groupi_n_2917, csa_tree_add_12_51_groupi_n_2918, csa_tree_add_12_51_groupi_n_2919, csa_tree_add_12_51_groupi_n_2920;
  wire csa_tree_add_12_51_groupi_n_2921, csa_tree_add_12_51_groupi_n_2922, csa_tree_add_12_51_groupi_n_2923, csa_tree_add_12_51_groupi_n_2924, csa_tree_add_12_51_groupi_n_2925, csa_tree_add_12_51_groupi_n_2926, csa_tree_add_12_51_groupi_n_2927, csa_tree_add_12_51_groupi_n_2928;
  wire csa_tree_add_12_51_groupi_n_2929, csa_tree_add_12_51_groupi_n_2930, csa_tree_add_12_51_groupi_n_2931, csa_tree_add_12_51_groupi_n_2932, csa_tree_add_12_51_groupi_n_2933, csa_tree_add_12_51_groupi_n_2934, csa_tree_add_12_51_groupi_n_2935, csa_tree_add_12_51_groupi_n_2936;
  wire csa_tree_add_12_51_groupi_n_2937, csa_tree_add_12_51_groupi_n_2938, csa_tree_add_12_51_groupi_n_2939, csa_tree_add_12_51_groupi_n_2940, csa_tree_add_12_51_groupi_n_2941, csa_tree_add_12_51_groupi_n_2942, csa_tree_add_12_51_groupi_n_2943, csa_tree_add_12_51_groupi_n_2944;
  wire csa_tree_add_12_51_groupi_n_2945, csa_tree_add_12_51_groupi_n_2946, csa_tree_add_12_51_groupi_n_2947, csa_tree_add_12_51_groupi_n_2948, csa_tree_add_12_51_groupi_n_2949, csa_tree_add_12_51_groupi_n_2950, csa_tree_add_12_51_groupi_n_2951, csa_tree_add_12_51_groupi_n_2952;
  wire csa_tree_add_12_51_groupi_n_2953, csa_tree_add_12_51_groupi_n_2954, csa_tree_add_12_51_groupi_n_2955, csa_tree_add_12_51_groupi_n_2956, csa_tree_add_12_51_groupi_n_2957, csa_tree_add_12_51_groupi_n_2958, csa_tree_add_12_51_groupi_n_2959, csa_tree_add_12_51_groupi_n_2960;
  wire csa_tree_add_12_51_groupi_n_2961, csa_tree_add_12_51_groupi_n_2962, csa_tree_add_12_51_groupi_n_2963, csa_tree_add_12_51_groupi_n_2964, csa_tree_add_12_51_groupi_n_2965, csa_tree_add_12_51_groupi_n_2966, csa_tree_add_12_51_groupi_n_2967, csa_tree_add_12_51_groupi_n_2968;
  wire csa_tree_add_12_51_groupi_n_2969, csa_tree_add_12_51_groupi_n_2970, csa_tree_add_12_51_groupi_n_2971, csa_tree_add_12_51_groupi_n_2972, csa_tree_add_12_51_groupi_n_2973, csa_tree_add_12_51_groupi_n_2974, csa_tree_add_12_51_groupi_n_2975, csa_tree_add_12_51_groupi_n_2976;
  wire csa_tree_add_12_51_groupi_n_2977, csa_tree_add_12_51_groupi_n_2978, csa_tree_add_12_51_groupi_n_2979, csa_tree_add_12_51_groupi_n_2980, csa_tree_add_12_51_groupi_n_2981, csa_tree_add_12_51_groupi_n_2982, csa_tree_add_12_51_groupi_n_2983, csa_tree_add_12_51_groupi_n_2984;
  wire csa_tree_add_12_51_groupi_n_2985, csa_tree_add_12_51_groupi_n_2986, csa_tree_add_12_51_groupi_n_2987, csa_tree_add_12_51_groupi_n_2988, csa_tree_add_12_51_groupi_n_2989, csa_tree_add_12_51_groupi_n_2990, csa_tree_add_12_51_groupi_n_2991, csa_tree_add_12_51_groupi_n_2992;
  wire csa_tree_add_12_51_groupi_n_2993, csa_tree_add_12_51_groupi_n_2994, csa_tree_add_12_51_groupi_n_2995, csa_tree_add_12_51_groupi_n_2996, csa_tree_add_12_51_groupi_n_2997, csa_tree_add_12_51_groupi_n_2998, csa_tree_add_12_51_groupi_n_2999, csa_tree_add_12_51_groupi_n_3000;
  wire csa_tree_add_12_51_groupi_n_3001, csa_tree_add_12_51_groupi_n_3002, csa_tree_add_12_51_groupi_n_3003, csa_tree_add_12_51_groupi_n_3004, csa_tree_add_12_51_groupi_n_3005, csa_tree_add_12_51_groupi_n_3006, csa_tree_add_12_51_groupi_n_3007, csa_tree_add_12_51_groupi_n_3008;
  wire csa_tree_add_12_51_groupi_n_3009, csa_tree_add_12_51_groupi_n_3010, csa_tree_add_12_51_groupi_n_3011, csa_tree_add_12_51_groupi_n_3012, csa_tree_add_12_51_groupi_n_3013, csa_tree_add_12_51_groupi_n_3014, csa_tree_add_12_51_groupi_n_3015, csa_tree_add_12_51_groupi_n_3016;
  wire csa_tree_add_12_51_groupi_n_3017, csa_tree_add_12_51_groupi_n_3018, csa_tree_add_12_51_groupi_n_3019, csa_tree_add_12_51_groupi_n_3020, csa_tree_add_12_51_groupi_n_3021, csa_tree_add_12_51_groupi_n_3022, csa_tree_add_12_51_groupi_n_3023, csa_tree_add_12_51_groupi_n_3024;
  wire csa_tree_add_12_51_groupi_n_3025, csa_tree_add_12_51_groupi_n_3026, csa_tree_add_12_51_groupi_n_3027, csa_tree_add_12_51_groupi_n_3028, csa_tree_add_12_51_groupi_n_3029, csa_tree_add_12_51_groupi_n_3030, csa_tree_add_12_51_groupi_n_3031, csa_tree_add_12_51_groupi_n_3032;
  wire csa_tree_add_12_51_groupi_n_3033, csa_tree_add_12_51_groupi_n_3034, csa_tree_add_12_51_groupi_n_3035, csa_tree_add_12_51_groupi_n_3036, csa_tree_add_12_51_groupi_n_3037, csa_tree_add_12_51_groupi_n_3038, csa_tree_add_12_51_groupi_n_3039, csa_tree_add_12_51_groupi_n_3040;
  wire csa_tree_add_12_51_groupi_n_3041, csa_tree_add_12_51_groupi_n_3042, csa_tree_add_12_51_groupi_n_3043, csa_tree_add_12_51_groupi_n_3044, csa_tree_add_12_51_groupi_n_3045, csa_tree_add_12_51_groupi_n_3046, csa_tree_add_12_51_groupi_n_3047, csa_tree_add_12_51_groupi_n_3048;
  wire csa_tree_add_12_51_groupi_n_3049, csa_tree_add_12_51_groupi_n_3050, csa_tree_add_12_51_groupi_n_3051, csa_tree_add_12_51_groupi_n_3052, csa_tree_add_12_51_groupi_n_3053, csa_tree_add_12_51_groupi_n_3054, csa_tree_add_12_51_groupi_n_3055, csa_tree_add_12_51_groupi_n_3056;
  wire csa_tree_add_12_51_groupi_n_3057, csa_tree_add_12_51_groupi_n_3058, csa_tree_add_12_51_groupi_n_3059, csa_tree_add_12_51_groupi_n_3060, csa_tree_add_12_51_groupi_n_3061, csa_tree_add_12_51_groupi_n_3062, csa_tree_add_12_51_groupi_n_3063, csa_tree_add_12_51_groupi_n_3064;
  wire csa_tree_add_12_51_groupi_n_3065, csa_tree_add_12_51_groupi_n_3066, csa_tree_add_12_51_groupi_n_3067, csa_tree_add_12_51_groupi_n_3068, csa_tree_add_12_51_groupi_n_3069, csa_tree_add_12_51_groupi_n_3070, csa_tree_add_12_51_groupi_n_3071, csa_tree_add_12_51_groupi_n_3072;
  wire csa_tree_add_12_51_groupi_n_3073, csa_tree_add_12_51_groupi_n_3074, csa_tree_add_12_51_groupi_n_3075, csa_tree_add_12_51_groupi_n_3076, csa_tree_add_12_51_groupi_n_3077, csa_tree_add_12_51_groupi_n_3078, csa_tree_add_12_51_groupi_n_3079, csa_tree_add_12_51_groupi_n_3080;
  wire csa_tree_add_12_51_groupi_n_3081, csa_tree_add_12_51_groupi_n_3082, csa_tree_add_12_51_groupi_n_3083, csa_tree_add_12_51_groupi_n_3084, csa_tree_add_12_51_groupi_n_3085, csa_tree_add_12_51_groupi_n_3086, csa_tree_add_12_51_groupi_n_3087, csa_tree_add_12_51_groupi_n_3088;
  wire csa_tree_add_12_51_groupi_n_3089, csa_tree_add_12_51_groupi_n_3090, csa_tree_add_12_51_groupi_n_3091, csa_tree_add_12_51_groupi_n_3092, csa_tree_add_12_51_groupi_n_3093, csa_tree_add_12_51_groupi_n_3094, csa_tree_add_12_51_groupi_n_3095, csa_tree_add_12_51_groupi_n_3096;
  wire csa_tree_add_12_51_groupi_n_3097, csa_tree_add_12_51_groupi_n_3098, csa_tree_add_12_51_groupi_n_3099, csa_tree_add_12_51_groupi_n_3100, csa_tree_add_12_51_groupi_n_3101, csa_tree_add_12_51_groupi_n_3102, csa_tree_add_12_51_groupi_n_3103, csa_tree_add_12_51_groupi_n_3104;
  wire csa_tree_add_12_51_groupi_n_3105, csa_tree_add_12_51_groupi_n_3106, csa_tree_add_12_51_groupi_n_3107, csa_tree_add_12_51_groupi_n_3108, csa_tree_add_12_51_groupi_n_3109, csa_tree_add_12_51_groupi_n_3110, csa_tree_add_12_51_groupi_n_3111, csa_tree_add_12_51_groupi_n_3112;
  wire csa_tree_add_12_51_groupi_n_3113, csa_tree_add_12_51_groupi_n_3114, csa_tree_add_12_51_groupi_n_3115, csa_tree_add_12_51_groupi_n_3116, csa_tree_add_12_51_groupi_n_3117, csa_tree_add_12_51_groupi_n_3118, csa_tree_add_12_51_groupi_n_3119, csa_tree_add_12_51_groupi_n_3120;
  wire csa_tree_add_12_51_groupi_n_3121, csa_tree_add_12_51_groupi_n_3122, csa_tree_add_12_51_groupi_n_3123, csa_tree_add_12_51_groupi_n_3124, csa_tree_add_12_51_groupi_n_3125, csa_tree_add_12_51_groupi_n_3126, csa_tree_add_12_51_groupi_n_3127, csa_tree_add_12_51_groupi_n_3128;
  wire csa_tree_add_12_51_groupi_n_3129, csa_tree_add_12_51_groupi_n_3130, csa_tree_add_12_51_groupi_n_3131, csa_tree_add_12_51_groupi_n_3132, csa_tree_add_12_51_groupi_n_3133, csa_tree_add_12_51_groupi_n_3134, csa_tree_add_12_51_groupi_n_3135, csa_tree_add_12_51_groupi_n_3136;
  wire csa_tree_add_12_51_groupi_n_3137, csa_tree_add_12_51_groupi_n_3138, csa_tree_add_12_51_groupi_n_3139, csa_tree_add_12_51_groupi_n_3140, csa_tree_add_12_51_groupi_n_3141, csa_tree_add_12_51_groupi_n_3142, csa_tree_add_12_51_groupi_n_3143, csa_tree_add_12_51_groupi_n_3144;
  wire csa_tree_add_12_51_groupi_n_3145, csa_tree_add_12_51_groupi_n_3146, csa_tree_add_12_51_groupi_n_3147, csa_tree_add_12_51_groupi_n_3148, csa_tree_add_12_51_groupi_n_3149, csa_tree_add_12_51_groupi_n_3150, csa_tree_add_12_51_groupi_n_3151, csa_tree_add_12_51_groupi_n_3152;
  wire csa_tree_add_12_51_groupi_n_3153, csa_tree_add_12_51_groupi_n_3154, csa_tree_add_12_51_groupi_n_3155, csa_tree_add_12_51_groupi_n_3156, csa_tree_add_12_51_groupi_n_3157, csa_tree_add_12_51_groupi_n_3158, csa_tree_add_12_51_groupi_n_3159, csa_tree_add_12_51_groupi_n_3160;
  wire csa_tree_add_12_51_groupi_n_3161, csa_tree_add_12_51_groupi_n_3162, csa_tree_add_12_51_groupi_n_3163, csa_tree_add_12_51_groupi_n_3164, csa_tree_add_12_51_groupi_n_3165, csa_tree_add_12_51_groupi_n_3166, csa_tree_add_12_51_groupi_n_3167, csa_tree_add_12_51_groupi_n_3168;
  wire csa_tree_add_12_51_groupi_n_3169, csa_tree_add_12_51_groupi_n_3170, csa_tree_add_12_51_groupi_n_3171, csa_tree_add_12_51_groupi_n_3172, csa_tree_add_12_51_groupi_n_3173, csa_tree_add_12_51_groupi_n_3174, csa_tree_add_12_51_groupi_n_3175, csa_tree_add_12_51_groupi_n_3176;
  wire csa_tree_add_12_51_groupi_n_3177, csa_tree_add_12_51_groupi_n_3178, csa_tree_add_12_51_groupi_n_3179, csa_tree_add_12_51_groupi_n_3180, csa_tree_add_12_51_groupi_n_3181, csa_tree_add_12_51_groupi_n_3182, csa_tree_add_12_51_groupi_n_3183, csa_tree_add_12_51_groupi_n_3184;
  wire csa_tree_add_12_51_groupi_n_3185, csa_tree_add_12_51_groupi_n_3186, csa_tree_add_12_51_groupi_n_3187, csa_tree_add_12_51_groupi_n_3188, csa_tree_add_12_51_groupi_n_3189, csa_tree_add_12_51_groupi_n_3190, csa_tree_add_12_51_groupi_n_3191, csa_tree_add_12_51_groupi_n_3192;
  wire csa_tree_add_12_51_groupi_n_3193, csa_tree_add_12_51_groupi_n_3194, csa_tree_add_12_51_groupi_n_3195, csa_tree_add_12_51_groupi_n_3196, csa_tree_add_12_51_groupi_n_3197, csa_tree_add_12_51_groupi_n_3198, csa_tree_add_12_51_groupi_n_3199, csa_tree_add_12_51_groupi_n_3200;
  wire csa_tree_add_12_51_groupi_n_3201, csa_tree_add_12_51_groupi_n_3202, csa_tree_add_12_51_groupi_n_3203, csa_tree_add_12_51_groupi_n_3204, csa_tree_add_12_51_groupi_n_3205, csa_tree_add_12_51_groupi_n_3206, csa_tree_add_12_51_groupi_n_3207, csa_tree_add_12_51_groupi_n_3208;
  wire csa_tree_add_12_51_groupi_n_3209, csa_tree_add_12_51_groupi_n_3210, csa_tree_add_12_51_groupi_n_3211, csa_tree_add_12_51_groupi_n_3212, csa_tree_add_12_51_groupi_n_3213, csa_tree_add_12_51_groupi_n_3214, csa_tree_add_12_51_groupi_n_3215, csa_tree_add_12_51_groupi_n_3216;
  wire csa_tree_add_12_51_groupi_n_3217, csa_tree_add_12_51_groupi_n_3218, csa_tree_add_12_51_groupi_n_3219, csa_tree_add_12_51_groupi_n_3220, csa_tree_add_12_51_groupi_n_3221, csa_tree_add_12_51_groupi_n_3222, csa_tree_add_12_51_groupi_n_3223, csa_tree_add_12_51_groupi_n_3224;
  wire csa_tree_add_12_51_groupi_n_3225, csa_tree_add_12_51_groupi_n_3226, csa_tree_add_12_51_groupi_n_3227, csa_tree_add_12_51_groupi_n_3228, csa_tree_add_12_51_groupi_n_3229, csa_tree_add_12_51_groupi_n_3230, csa_tree_add_12_51_groupi_n_3231, csa_tree_add_12_51_groupi_n_3232;
  wire csa_tree_add_12_51_groupi_n_3233, csa_tree_add_12_51_groupi_n_3234, csa_tree_add_12_51_groupi_n_3235, csa_tree_add_12_51_groupi_n_3236, csa_tree_add_12_51_groupi_n_3237, csa_tree_add_12_51_groupi_n_3238, csa_tree_add_12_51_groupi_n_3239, csa_tree_add_12_51_groupi_n_3240;
  wire csa_tree_add_12_51_groupi_n_3241, csa_tree_add_12_51_groupi_n_3242, csa_tree_add_12_51_groupi_n_3243, csa_tree_add_12_51_groupi_n_3244, csa_tree_add_12_51_groupi_n_3245, csa_tree_add_12_51_groupi_n_3246, csa_tree_add_12_51_groupi_n_3247, csa_tree_add_12_51_groupi_n_3248;
  wire csa_tree_add_12_51_groupi_n_3249, csa_tree_add_12_51_groupi_n_3250, csa_tree_add_12_51_groupi_n_3251, csa_tree_add_12_51_groupi_n_3252, csa_tree_add_12_51_groupi_n_3253, csa_tree_add_12_51_groupi_n_3254, csa_tree_add_12_51_groupi_n_3255, csa_tree_add_12_51_groupi_n_3256;
  wire csa_tree_add_12_51_groupi_n_3257, csa_tree_add_12_51_groupi_n_3258, csa_tree_add_12_51_groupi_n_3259, csa_tree_add_12_51_groupi_n_3260, csa_tree_add_12_51_groupi_n_3261, csa_tree_add_12_51_groupi_n_3262, csa_tree_add_12_51_groupi_n_3263, csa_tree_add_12_51_groupi_n_3264;
  wire csa_tree_add_12_51_groupi_n_3265, csa_tree_add_12_51_groupi_n_3266, csa_tree_add_12_51_groupi_n_3267, csa_tree_add_12_51_groupi_n_3268, csa_tree_add_12_51_groupi_n_3269, csa_tree_add_12_51_groupi_n_3270, csa_tree_add_12_51_groupi_n_3271, csa_tree_add_12_51_groupi_n_3272;
  wire csa_tree_add_12_51_groupi_n_3273, csa_tree_add_12_51_groupi_n_3274, csa_tree_add_12_51_groupi_n_3275, csa_tree_add_12_51_groupi_n_3276, csa_tree_add_12_51_groupi_n_3277, csa_tree_add_12_51_groupi_n_3278, csa_tree_add_12_51_groupi_n_3279, csa_tree_add_12_51_groupi_n_3280;
  wire csa_tree_add_12_51_groupi_n_3281, csa_tree_add_12_51_groupi_n_3282, csa_tree_add_12_51_groupi_n_3283, csa_tree_add_12_51_groupi_n_3284, csa_tree_add_12_51_groupi_n_3285, csa_tree_add_12_51_groupi_n_3286, csa_tree_add_12_51_groupi_n_3287, csa_tree_add_12_51_groupi_n_3288;
  wire csa_tree_add_12_51_groupi_n_3289, csa_tree_add_12_51_groupi_n_3290, csa_tree_add_12_51_groupi_n_3291, csa_tree_add_12_51_groupi_n_3292, csa_tree_add_12_51_groupi_n_3293, csa_tree_add_12_51_groupi_n_3294, csa_tree_add_12_51_groupi_n_3295, csa_tree_add_12_51_groupi_n_3296;
  wire csa_tree_add_12_51_groupi_n_3297, csa_tree_add_12_51_groupi_n_3298, csa_tree_add_12_51_groupi_n_3299, csa_tree_add_12_51_groupi_n_3300, csa_tree_add_12_51_groupi_n_3301, csa_tree_add_12_51_groupi_n_3302, csa_tree_add_12_51_groupi_n_3303, csa_tree_add_12_51_groupi_n_3304;
  wire csa_tree_add_12_51_groupi_n_3305, csa_tree_add_12_51_groupi_n_3306, csa_tree_add_12_51_groupi_n_3307, csa_tree_add_12_51_groupi_n_3308, csa_tree_add_12_51_groupi_n_3309, csa_tree_add_12_51_groupi_n_3310, csa_tree_add_12_51_groupi_n_3311, csa_tree_add_12_51_groupi_n_3312;
  wire csa_tree_add_12_51_groupi_n_3313, csa_tree_add_12_51_groupi_n_3314, csa_tree_add_12_51_groupi_n_3315, csa_tree_add_12_51_groupi_n_3316, csa_tree_add_12_51_groupi_n_3317, csa_tree_add_12_51_groupi_n_3318, csa_tree_add_12_51_groupi_n_3319, csa_tree_add_12_51_groupi_n_3320;
  wire csa_tree_add_12_51_groupi_n_3321, csa_tree_add_12_51_groupi_n_3322, csa_tree_add_12_51_groupi_n_3323, csa_tree_add_12_51_groupi_n_3324, csa_tree_add_12_51_groupi_n_3325, csa_tree_add_12_51_groupi_n_3326, csa_tree_add_12_51_groupi_n_3327, csa_tree_add_12_51_groupi_n_3328;
  wire csa_tree_add_12_51_groupi_n_3329, csa_tree_add_12_51_groupi_n_3330, csa_tree_add_12_51_groupi_n_3331, csa_tree_add_12_51_groupi_n_3332, csa_tree_add_12_51_groupi_n_3333, csa_tree_add_12_51_groupi_n_3334, csa_tree_add_12_51_groupi_n_3335, csa_tree_add_12_51_groupi_n_3336;
  wire csa_tree_add_12_51_groupi_n_3337, csa_tree_add_12_51_groupi_n_3338, csa_tree_add_12_51_groupi_n_3339, csa_tree_add_12_51_groupi_n_3340, csa_tree_add_12_51_groupi_n_3341, csa_tree_add_12_51_groupi_n_3342, csa_tree_add_12_51_groupi_n_3343, csa_tree_add_12_51_groupi_n_3344;
  wire csa_tree_add_12_51_groupi_n_3345, csa_tree_add_12_51_groupi_n_3346, csa_tree_add_12_51_groupi_n_3347, csa_tree_add_12_51_groupi_n_3348, csa_tree_add_12_51_groupi_n_3349, csa_tree_add_12_51_groupi_n_3350, csa_tree_add_12_51_groupi_n_3351, csa_tree_add_12_51_groupi_n_3352;
  wire csa_tree_add_12_51_groupi_n_3353, csa_tree_add_12_51_groupi_n_3354, csa_tree_add_12_51_groupi_n_3355, csa_tree_add_12_51_groupi_n_3356, csa_tree_add_12_51_groupi_n_3357, csa_tree_add_12_51_groupi_n_3358, csa_tree_add_12_51_groupi_n_3359, csa_tree_add_12_51_groupi_n_3360;
  wire csa_tree_add_12_51_groupi_n_3361, csa_tree_add_12_51_groupi_n_3362, csa_tree_add_12_51_groupi_n_3363, csa_tree_add_12_51_groupi_n_3364, csa_tree_add_12_51_groupi_n_3365, csa_tree_add_12_51_groupi_n_3366, csa_tree_add_12_51_groupi_n_3367, csa_tree_add_12_51_groupi_n_3368;
  wire csa_tree_add_12_51_groupi_n_3369, csa_tree_add_12_51_groupi_n_3370, csa_tree_add_12_51_groupi_n_3371, csa_tree_add_12_51_groupi_n_3372, csa_tree_add_12_51_groupi_n_3373, csa_tree_add_12_51_groupi_n_3374, csa_tree_add_12_51_groupi_n_3375, csa_tree_add_12_51_groupi_n_3376;
  wire csa_tree_add_12_51_groupi_n_3377, csa_tree_add_12_51_groupi_n_3378, csa_tree_add_12_51_groupi_n_3379, csa_tree_add_12_51_groupi_n_3380, csa_tree_add_12_51_groupi_n_3381, csa_tree_add_12_51_groupi_n_3382, csa_tree_add_12_51_groupi_n_3383, csa_tree_add_12_51_groupi_n_3384;
  wire csa_tree_add_12_51_groupi_n_3385, csa_tree_add_12_51_groupi_n_3386, csa_tree_add_12_51_groupi_n_3387, csa_tree_add_12_51_groupi_n_3388, csa_tree_add_12_51_groupi_n_3389, csa_tree_add_12_51_groupi_n_3390, csa_tree_add_12_51_groupi_n_3391, csa_tree_add_12_51_groupi_n_3392;
  wire csa_tree_add_12_51_groupi_n_3393, csa_tree_add_12_51_groupi_n_3394, csa_tree_add_12_51_groupi_n_3395, csa_tree_add_12_51_groupi_n_3396, csa_tree_add_12_51_groupi_n_3397, csa_tree_add_12_51_groupi_n_3398, csa_tree_add_12_51_groupi_n_3399, csa_tree_add_12_51_groupi_n_3400;
  wire csa_tree_add_12_51_groupi_n_3401, csa_tree_add_12_51_groupi_n_3402, csa_tree_add_12_51_groupi_n_3403, csa_tree_add_12_51_groupi_n_3404, csa_tree_add_12_51_groupi_n_3405, csa_tree_add_12_51_groupi_n_3406, csa_tree_add_12_51_groupi_n_3407, csa_tree_add_12_51_groupi_n_3408;
  wire csa_tree_add_12_51_groupi_n_3409, csa_tree_add_12_51_groupi_n_3410, csa_tree_add_12_51_groupi_n_3411, csa_tree_add_12_51_groupi_n_3412, csa_tree_add_12_51_groupi_n_3413, csa_tree_add_12_51_groupi_n_3414, csa_tree_add_12_51_groupi_n_3415, csa_tree_add_12_51_groupi_n_3416;
  wire csa_tree_add_12_51_groupi_n_3417, csa_tree_add_12_51_groupi_n_3418, csa_tree_add_12_51_groupi_n_3419, csa_tree_add_12_51_groupi_n_3420, csa_tree_add_12_51_groupi_n_3421, csa_tree_add_12_51_groupi_n_3422, csa_tree_add_12_51_groupi_n_3423, csa_tree_add_12_51_groupi_n_3424;
  wire csa_tree_add_12_51_groupi_n_3425, csa_tree_add_12_51_groupi_n_3426, csa_tree_add_12_51_groupi_n_3427, csa_tree_add_12_51_groupi_n_3428, csa_tree_add_12_51_groupi_n_3429, csa_tree_add_12_51_groupi_n_3430, csa_tree_add_12_51_groupi_n_3431, csa_tree_add_12_51_groupi_n_3432;
  wire csa_tree_add_12_51_groupi_n_3433, csa_tree_add_12_51_groupi_n_3434, csa_tree_add_12_51_groupi_n_3435, csa_tree_add_12_51_groupi_n_3436, csa_tree_add_12_51_groupi_n_3437, csa_tree_add_12_51_groupi_n_3438, csa_tree_add_12_51_groupi_n_3439, csa_tree_add_12_51_groupi_n_3440;
  wire csa_tree_add_12_51_groupi_n_3441, csa_tree_add_12_51_groupi_n_3442, csa_tree_add_12_51_groupi_n_3443, csa_tree_add_12_51_groupi_n_3444, csa_tree_add_12_51_groupi_n_3445, csa_tree_add_12_51_groupi_n_3446, csa_tree_add_12_51_groupi_n_3447, csa_tree_add_12_51_groupi_n_3448;
  wire csa_tree_add_12_51_groupi_n_3449, csa_tree_add_12_51_groupi_n_3450, csa_tree_add_12_51_groupi_n_3451, csa_tree_add_12_51_groupi_n_3452, csa_tree_add_12_51_groupi_n_3453, csa_tree_add_12_51_groupi_n_3454, csa_tree_add_12_51_groupi_n_3455, csa_tree_add_12_51_groupi_n_3456;
  wire csa_tree_add_12_51_groupi_n_3457, csa_tree_add_12_51_groupi_n_3458, csa_tree_add_12_51_groupi_n_3459, csa_tree_add_12_51_groupi_n_3460, csa_tree_add_12_51_groupi_n_3461, csa_tree_add_12_51_groupi_n_3462, csa_tree_add_12_51_groupi_n_3463, csa_tree_add_12_51_groupi_n_3464;
  wire csa_tree_add_12_51_groupi_n_3465, csa_tree_add_12_51_groupi_n_3466, csa_tree_add_12_51_groupi_n_3467, csa_tree_add_12_51_groupi_n_3468, csa_tree_add_12_51_groupi_n_3469, csa_tree_add_12_51_groupi_n_3470, csa_tree_add_12_51_groupi_n_3471, csa_tree_add_12_51_groupi_n_3472;
  wire csa_tree_add_12_51_groupi_n_3473, csa_tree_add_12_51_groupi_n_3474, csa_tree_add_12_51_groupi_n_3475, csa_tree_add_12_51_groupi_n_3476, csa_tree_add_12_51_groupi_n_3477, csa_tree_add_12_51_groupi_n_3478, csa_tree_add_12_51_groupi_n_3479, csa_tree_add_12_51_groupi_n_3480;
  wire csa_tree_add_12_51_groupi_n_3481, csa_tree_add_12_51_groupi_n_3482, csa_tree_add_12_51_groupi_n_3483, csa_tree_add_12_51_groupi_n_3484, csa_tree_add_12_51_groupi_n_3485, csa_tree_add_12_51_groupi_n_3486, csa_tree_add_12_51_groupi_n_3487, csa_tree_add_12_51_groupi_n_3488;
  wire csa_tree_add_12_51_groupi_n_3489, csa_tree_add_12_51_groupi_n_3490, csa_tree_add_12_51_groupi_n_3491, csa_tree_add_12_51_groupi_n_3492, csa_tree_add_12_51_groupi_n_3493, csa_tree_add_12_51_groupi_n_3494, csa_tree_add_12_51_groupi_n_3495, csa_tree_add_12_51_groupi_n_3496;
  wire csa_tree_add_12_51_groupi_n_3497, csa_tree_add_12_51_groupi_n_3498, csa_tree_add_12_51_groupi_n_3499, csa_tree_add_12_51_groupi_n_3500, csa_tree_add_12_51_groupi_n_3501, csa_tree_add_12_51_groupi_n_3502, csa_tree_add_12_51_groupi_n_3503, csa_tree_add_12_51_groupi_n_3504;
  wire csa_tree_add_12_51_groupi_n_3505, csa_tree_add_12_51_groupi_n_3506, csa_tree_add_12_51_groupi_n_3507, csa_tree_add_12_51_groupi_n_3508, csa_tree_add_12_51_groupi_n_3509, csa_tree_add_12_51_groupi_n_3510, csa_tree_add_12_51_groupi_n_3511, csa_tree_add_12_51_groupi_n_3512;
  wire csa_tree_add_12_51_groupi_n_3513, csa_tree_add_12_51_groupi_n_3514, csa_tree_add_12_51_groupi_n_3515, csa_tree_add_12_51_groupi_n_3516, csa_tree_add_12_51_groupi_n_3517, csa_tree_add_12_51_groupi_n_3518, csa_tree_add_12_51_groupi_n_3519, csa_tree_add_12_51_groupi_n_3520;
  wire csa_tree_add_12_51_groupi_n_3521, csa_tree_add_12_51_groupi_n_3522, csa_tree_add_12_51_groupi_n_3523, csa_tree_add_12_51_groupi_n_3524, csa_tree_add_12_51_groupi_n_3525, csa_tree_add_12_51_groupi_n_3526, csa_tree_add_12_51_groupi_n_3527, csa_tree_add_12_51_groupi_n_3528;
  wire csa_tree_add_12_51_groupi_n_3529, csa_tree_add_12_51_groupi_n_3530, csa_tree_add_12_51_groupi_n_3531, csa_tree_add_12_51_groupi_n_3532, csa_tree_add_12_51_groupi_n_3533, csa_tree_add_12_51_groupi_n_3534, csa_tree_add_12_51_groupi_n_3535, csa_tree_add_12_51_groupi_n_3536;
  wire csa_tree_add_12_51_groupi_n_3537, csa_tree_add_12_51_groupi_n_3538, csa_tree_add_12_51_groupi_n_3539, csa_tree_add_12_51_groupi_n_3540, csa_tree_add_12_51_groupi_n_3541, csa_tree_add_12_51_groupi_n_3542, csa_tree_add_12_51_groupi_n_3543, csa_tree_add_12_51_groupi_n_3544;
  wire csa_tree_add_12_51_groupi_n_3545, csa_tree_add_12_51_groupi_n_3546, csa_tree_add_12_51_groupi_n_3547, csa_tree_add_12_51_groupi_n_3548, csa_tree_add_12_51_groupi_n_3549, csa_tree_add_12_51_groupi_n_3550, csa_tree_add_12_51_groupi_n_3551, csa_tree_add_12_51_groupi_n_3552;
  wire csa_tree_add_12_51_groupi_n_3553, csa_tree_add_12_51_groupi_n_3554, csa_tree_add_12_51_groupi_n_3555, csa_tree_add_12_51_groupi_n_3556, csa_tree_add_12_51_groupi_n_3557, csa_tree_add_12_51_groupi_n_3558, csa_tree_add_12_51_groupi_n_3559, csa_tree_add_12_51_groupi_n_3560;
  wire csa_tree_add_12_51_groupi_n_3561, csa_tree_add_12_51_groupi_n_3562, csa_tree_add_12_51_groupi_n_3563, csa_tree_add_12_51_groupi_n_3564, csa_tree_add_12_51_groupi_n_3565, csa_tree_add_12_51_groupi_n_3566, csa_tree_add_12_51_groupi_n_3567, csa_tree_add_12_51_groupi_n_3568;
  wire csa_tree_add_12_51_groupi_n_3569, csa_tree_add_12_51_groupi_n_3570, csa_tree_add_12_51_groupi_n_3571, csa_tree_add_12_51_groupi_n_3572, csa_tree_add_12_51_groupi_n_3573, csa_tree_add_12_51_groupi_n_3574, csa_tree_add_12_51_groupi_n_3575, csa_tree_add_12_51_groupi_n_3576;
  wire csa_tree_add_12_51_groupi_n_3577, csa_tree_add_12_51_groupi_n_3578, csa_tree_add_12_51_groupi_n_3579, csa_tree_add_12_51_groupi_n_3580, csa_tree_add_12_51_groupi_n_3581, csa_tree_add_12_51_groupi_n_3582, csa_tree_add_12_51_groupi_n_3583, csa_tree_add_12_51_groupi_n_3584;
  wire csa_tree_add_12_51_groupi_n_3585, csa_tree_add_12_51_groupi_n_3586, csa_tree_add_12_51_groupi_n_3587, csa_tree_add_12_51_groupi_n_3588, csa_tree_add_12_51_groupi_n_3589, csa_tree_add_12_51_groupi_n_3590, csa_tree_add_12_51_groupi_n_3591, csa_tree_add_12_51_groupi_n_3592;
  wire csa_tree_add_12_51_groupi_n_3593, csa_tree_add_12_51_groupi_n_3594, csa_tree_add_12_51_groupi_n_3595, csa_tree_add_12_51_groupi_n_3596, csa_tree_add_12_51_groupi_n_3597, csa_tree_add_12_51_groupi_n_3598, csa_tree_add_12_51_groupi_n_3599, csa_tree_add_12_51_groupi_n_3600;
  wire csa_tree_add_12_51_groupi_n_3601, csa_tree_add_12_51_groupi_n_3602, csa_tree_add_12_51_groupi_n_3603, csa_tree_add_12_51_groupi_n_3604, csa_tree_add_12_51_groupi_n_3605, csa_tree_add_12_51_groupi_n_3606, csa_tree_add_12_51_groupi_n_3607, csa_tree_add_12_51_groupi_n_3608;
  wire csa_tree_add_12_51_groupi_n_3609, csa_tree_add_12_51_groupi_n_3610, csa_tree_add_12_51_groupi_n_3611, csa_tree_add_12_51_groupi_n_3612, csa_tree_add_12_51_groupi_n_3613, csa_tree_add_12_51_groupi_n_3614, csa_tree_add_12_51_groupi_n_3615, csa_tree_add_12_51_groupi_n_3616;
  wire csa_tree_add_12_51_groupi_n_3617, csa_tree_add_12_51_groupi_n_3618, csa_tree_add_12_51_groupi_n_3619, csa_tree_add_12_51_groupi_n_3620, csa_tree_add_12_51_groupi_n_3621, csa_tree_add_12_51_groupi_n_3622, csa_tree_add_12_51_groupi_n_3623, csa_tree_add_12_51_groupi_n_3624;
  wire csa_tree_add_12_51_groupi_n_3625, csa_tree_add_12_51_groupi_n_3626, csa_tree_add_12_51_groupi_n_3627, csa_tree_add_12_51_groupi_n_3628, csa_tree_add_12_51_groupi_n_3629, csa_tree_add_12_51_groupi_n_3630, csa_tree_add_12_51_groupi_n_3631, csa_tree_add_12_51_groupi_n_3632;
  wire csa_tree_add_12_51_groupi_n_3633, csa_tree_add_12_51_groupi_n_3634, csa_tree_add_12_51_groupi_n_3635, csa_tree_add_12_51_groupi_n_3636, csa_tree_add_12_51_groupi_n_3637, csa_tree_add_12_51_groupi_n_3638, csa_tree_add_12_51_groupi_n_3639, csa_tree_add_12_51_groupi_n_3640;
  wire csa_tree_add_12_51_groupi_n_3641, csa_tree_add_12_51_groupi_n_3642, csa_tree_add_12_51_groupi_n_3643, csa_tree_add_12_51_groupi_n_3644, csa_tree_add_12_51_groupi_n_3645, csa_tree_add_12_51_groupi_n_3646, csa_tree_add_12_51_groupi_n_3647, csa_tree_add_12_51_groupi_n_3648;
  wire csa_tree_add_12_51_groupi_n_3649, csa_tree_add_12_51_groupi_n_3650, csa_tree_add_12_51_groupi_n_3651, csa_tree_add_12_51_groupi_n_3652, csa_tree_add_12_51_groupi_n_3653, csa_tree_add_12_51_groupi_n_3654, csa_tree_add_12_51_groupi_n_3655, csa_tree_add_12_51_groupi_n_3656;
  wire csa_tree_add_12_51_groupi_n_3657, csa_tree_add_12_51_groupi_n_3658, csa_tree_add_12_51_groupi_n_3659, csa_tree_add_12_51_groupi_n_3660, csa_tree_add_12_51_groupi_n_3661, csa_tree_add_12_51_groupi_n_3662, csa_tree_add_12_51_groupi_n_3663, csa_tree_add_12_51_groupi_n_3664;
  wire csa_tree_add_12_51_groupi_n_3665, csa_tree_add_12_51_groupi_n_3666, csa_tree_add_12_51_groupi_n_3667, csa_tree_add_12_51_groupi_n_3668, csa_tree_add_12_51_groupi_n_3669, csa_tree_add_12_51_groupi_n_3670, csa_tree_add_12_51_groupi_n_3671, csa_tree_add_12_51_groupi_n_3672;
  wire csa_tree_add_12_51_groupi_n_3673, csa_tree_add_12_51_groupi_n_3674, csa_tree_add_12_51_groupi_n_3675, csa_tree_add_12_51_groupi_n_3676, csa_tree_add_12_51_groupi_n_3677, csa_tree_add_12_51_groupi_n_3678, csa_tree_add_12_51_groupi_n_3679, csa_tree_add_12_51_groupi_n_3680;
  wire csa_tree_add_12_51_groupi_n_3681, csa_tree_add_12_51_groupi_n_3682, csa_tree_add_12_51_groupi_n_3683, csa_tree_add_12_51_groupi_n_3684, csa_tree_add_12_51_groupi_n_3685, csa_tree_add_12_51_groupi_n_3686, csa_tree_add_12_51_groupi_n_3687, csa_tree_add_12_51_groupi_n_3688;
  wire csa_tree_add_12_51_groupi_n_3689, csa_tree_add_12_51_groupi_n_3690, csa_tree_add_12_51_groupi_n_3691, csa_tree_add_12_51_groupi_n_3692, csa_tree_add_12_51_groupi_n_3693, csa_tree_add_12_51_groupi_n_3694, csa_tree_add_12_51_groupi_n_3695, csa_tree_add_12_51_groupi_n_3696;
  wire csa_tree_add_12_51_groupi_n_3697, csa_tree_add_12_51_groupi_n_3698, csa_tree_add_12_51_groupi_n_3699, csa_tree_add_12_51_groupi_n_3700, csa_tree_add_12_51_groupi_n_3701, csa_tree_add_12_51_groupi_n_3702, csa_tree_add_12_51_groupi_n_3703, csa_tree_add_12_51_groupi_n_3704;
  wire csa_tree_add_12_51_groupi_n_3705, csa_tree_add_12_51_groupi_n_3706, csa_tree_add_12_51_groupi_n_3707, csa_tree_add_12_51_groupi_n_3708, csa_tree_add_12_51_groupi_n_3709, csa_tree_add_12_51_groupi_n_3710, csa_tree_add_12_51_groupi_n_3711, csa_tree_add_12_51_groupi_n_3712;
  wire csa_tree_add_12_51_groupi_n_3713, csa_tree_add_12_51_groupi_n_3714, csa_tree_add_12_51_groupi_n_3715, csa_tree_add_12_51_groupi_n_3716, csa_tree_add_12_51_groupi_n_3717, csa_tree_add_12_51_groupi_n_3718, csa_tree_add_12_51_groupi_n_3719, csa_tree_add_12_51_groupi_n_3720;
  wire csa_tree_add_12_51_groupi_n_3721, csa_tree_add_12_51_groupi_n_3722, csa_tree_add_12_51_groupi_n_3723, csa_tree_add_12_51_groupi_n_3724, csa_tree_add_12_51_groupi_n_3725, csa_tree_add_12_51_groupi_n_3726, csa_tree_add_12_51_groupi_n_3727, csa_tree_add_12_51_groupi_n_3728;
  wire csa_tree_add_12_51_groupi_n_3729, csa_tree_add_12_51_groupi_n_3730, csa_tree_add_12_51_groupi_n_3731, csa_tree_add_12_51_groupi_n_3732, csa_tree_add_12_51_groupi_n_3733, csa_tree_add_12_51_groupi_n_3734, csa_tree_add_12_51_groupi_n_3735, csa_tree_add_12_51_groupi_n_3736;
  wire csa_tree_add_12_51_groupi_n_3737, csa_tree_add_12_51_groupi_n_3738, csa_tree_add_12_51_groupi_n_3739, csa_tree_add_12_51_groupi_n_3740, csa_tree_add_12_51_groupi_n_3741, csa_tree_add_12_51_groupi_n_3742, csa_tree_add_12_51_groupi_n_3743, csa_tree_add_12_51_groupi_n_3744;
  wire csa_tree_add_12_51_groupi_n_3745, csa_tree_add_12_51_groupi_n_3746, csa_tree_add_12_51_groupi_n_3747, csa_tree_add_12_51_groupi_n_3748, csa_tree_add_12_51_groupi_n_3749, csa_tree_add_12_51_groupi_n_3750, csa_tree_add_12_51_groupi_n_3751, csa_tree_add_12_51_groupi_n_3752;
  wire csa_tree_add_12_51_groupi_n_3753, csa_tree_add_12_51_groupi_n_3754, csa_tree_add_12_51_groupi_n_3755, csa_tree_add_12_51_groupi_n_3756, csa_tree_add_12_51_groupi_n_3757, csa_tree_add_12_51_groupi_n_3758, csa_tree_add_12_51_groupi_n_3759, csa_tree_add_12_51_groupi_n_3760;
  wire csa_tree_add_12_51_groupi_n_3761, csa_tree_add_12_51_groupi_n_3762, csa_tree_add_12_51_groupi_n_3763, csa_tree_add_12_51_groupi_n_3764, csa_tree_add_12_51_groupi_n_3765, csa_tree_add_12_51_groupi_n_3766, csa_tree_add_12_51_groupi_n_3767, csa_tree_add_12_51_groupi_n_3768;
  wire csa_tree_add_12_51_groupi_n_3769, csa_tree_add_12_51_groupi_n_3770, csa_tree_add_12_51_groupi_n_3771, csa_tree_add_12_51_groupi_n_3772, csa_tree_add_12_51_groupi_n_3773, csa_tree_add_12_51_groupi_n_3774, csa_tree_add_12_51_groupi_n_3775, csa_tree_add_12_51_groupi_n_3776;
  wire csa_tree_add_12_51_groupi_n_3777, csa_tree_add_12_51_groupi_n_3778, csa_tree_add_12_51_groupi_n_3779, csa_tree_add_12_51_groupi_n_3780, csa_tree_add_12_51_groupi_n_3781, csa_tree_add_12_51_groupi_n_3782, csa_tree_add_12_51_groupi_n_3783, csa_tree_add_12_51_groupi_n_3784;
  wire csa_tree_add_12_51_groupi_n_3785, csa_tree_add_12_51_groupi_n_3786, csa_tree_add_12_51_groupi_n_3787, csa_tree_add_12_51_groupi_n_3788, csa_tree_add_12_51_groupi_n_3789, csa_tree_add_12_51_groupi_n_3790, csa_tree_add_12_51_groupi_n_3791, csa_tree_add_12_51_groupi_n_3792;
  wire csa_tree_add_12_51_groupi_n_3793, csa_tree_add_12_51_groupi_n_3794, csa_tree_add_12_51_groupi_n_3795, csa_tree_add_12_51_groupi_n_3796, csa_tree_add_12_51_groupi_n_3797, csa_tree_add_12_51_groupi_n_3798, csa_tree_add_12_51_groupi_n_3799, csa_tree_add_12_51_groupi_n_3800;
  wire csa_tree_add_12_51_groupi_n_3801, csa_tree_add_12_51_groupi_n_3802, csa_tree_add_12_51_groupi_n_3803, csa_tree_add_12_51_groupi_n_3804, csa_tree_add_12_51_groupi_n_3805, csa_tree_add_12_51_groupi_n_3806, csa_tree_add_12_51_groupi_n_3807, csa_tree_add_12_51_groupi_n_3808;
  wire csa_tree_add_12_51_groupi_n_3809, csa_tree_add_12_51_groupi_n_3810, csa_tree_add_12_51_groupi_n_3811, csa_tree_add_12_51_groupi_n_3812, csa_tree_add_12_51_groupi_n_3813, csa_tree_add_12_51_groupi_n_3814, csa_tree_add_12_51_groupi_n_3815, csa_tree_add_12_51_groupi_n_3816;
  wire csa_tree_add_12_51_groupi_n_3817, csa_tree_add_12_51_groupi_n_3818, csa_tree_add_12_51_groupi_n_3819, csa_tree_add_12_51_groupi_n_3820, csa_tree_add_12_51_groupi_n_3821, csa_tree_add_12_51_groupi_n_3822, csa_tree_add_12_51_groupi_n_3823, csa_tree_add_12_51_groupi_n_3824;
  wire csa_tree_add_12_51_groupi_n_3825, csa_tree_add_12_51_groupi_n_3826, csa_tree_add_12_51_groupi_n_3827, csa_tree_add_12_51_groupi_n_3828, csa_tree_add_12_51_groupi_n_3829, csa_tree_add_12_51_groupi_n_3830, csa_tree_add_12_51_groupi_n_3831, csa_tree_add_12_51_groupi_n_3832;
  wire csa_tree_add_12_51_groupi_n_3833, csa_tree_add_12_51_groupi_n_3834, csa_tree_add_12_51_groupi_n_3835, csa_tree_add_12_51_groupi_n_3836, csa_tree_add_12_51_groupi_n_3837, csa_tree_add_12_51_groupi_n_3838, csa_tree_add_12_51_groupi_n_3839, csa_tree_add_12_51_groupi_n_3840;
  wire csa_tree_add_12_51_groupi_n_3841, csa_tree_add_12_51_groupi_n_3842, csa_tree_add_12_51_groupi_n_3843, csa_tree_add_12_51_groupi_n_3844, csa_tree_add_12_51_groupi_n_3845, csa_tree_add_12_51_groupi_n_3846, csa_tree_add_12_51_groupi_n_3847, csa_tree_add_12_51_groupi_n_3848;
  wire csa_tree_add_12_51_groupi_n_3849, csa_tree_add_12_51_groupi_n_3850, csa_tree_add_12_51_groupi_n_3851, csa_tree_add_12_51_groupi_n_3852, csa_tree_add_12_51_groupi_n_3853, csa_tree_add_12_51_groupi_n_3854, csa_tree_add_12_51_groupi_n_3855, csa_tree_add_12_51_groupi_n_3856;
  wire csa_tree_add_12_51_groupi_n_3857, csa_tree_add_12_51_groupi_n_3858, csa_tree_add_12_51_groupi_n_3859, csa_tree_add_12_51_groupi_n_3860, csa_tree_add_12_51_groupi_n_3861, csa_tree_add_12_51_groupi_n_3862, csa_tree_add_12_51_groupi_n_3863, csa_tree_add_12_51_groupi_n_3864;
  wire csa_tree_add_12_51_groupi_n_3865, csa_tree_add_12_51_groupi_n_3866, csa_tree_add_12_51_groupi_n_3867, csa_tree_add_12_51_groupi_n_3868, csa_tree_add_12_51_groupi_n_3869, csa_tree_add_12_51_groupi_n_3870, csa_tree_add_12_51_groupi_n_3871, csa_tree_add_12_51_groupi_n_3872;
  wire csa_tree_add_12_51_groupi_n_3873, csa_tree_add_12_51_groupi_n_3874, csa_tree_add_12_51_groupi_n_3875, csa_tree_add_12_51_groupi_n_3876, csa_tree_add_12_51_groupi_n_3877, csa_tree_add_12_51_groupi_n_3878, csa_tree_add_12_51_groupi_n_3879, csa_tree_add_12_51_groupi_n_3880;
  wire csa_tree_add_12_51_groupi_n_3881, csa_tree_add_12_51_groupi_n_3882, csa_tree_add_12_51_groupi_n_3883, csa_tree_add_12_51_groupi_n_3884, csa_tree_add_12_51_groupi_n_3885, csa_tree_add_12_51_groupi_n_3886, csa_tree_add_12_51_groupi_n_3887, csa_tree_add_12_51_groupi_n_3888;
  wire csa_tree_add_12_51_groupi_n_3889, csa_tree_add_12_51_groupi_n_3890, csa_tree_add_12_51_groupi_n_3891, csa_tree_add_12_51_groupi_n_3892, csa_tree_add_12_51_groupi_n_3893, csa_tree_add_12_51_groupi_n_3894, csa_tree_add_12_51_groupi_n_3895, csa_tree_add_12_51_groupi_n_3896;
  wire csa_tree_add_12_51_groupi_n_3897, csa_tree_add_12_51_groupi_n_3898, csa_tree_add_12_51_groupi_n_3899, csa_tree_add_12_51_groupi_n_3900, csa_tree_add_12_51_groupi_n_3901, csa_tree_add_12_51_groupi_n_3902, csa_tree_add_12_51_groupi_n_3903, csa_tree_add_12_51_groupi_n_3904;
  wire csa_tree_add_12_51_groupi_n_3905, csa_tree_add_12_51_groupi_n_3906, csa_tree_add_12_51_groupi_n_3907, csa_tree_add_12_51_groupi_n_3908, csa_tree_add_12_51_groupi_n_3909, csa_tree_add_12_51_groupi_n_3910, csa_tree_add_12_51_groupi_n_3911, csa_tree_add_12_51_groupi_n_3912;
  wire csa_tree_add_12_51_groupi_n_3913, csa_tree_add_12_51_groupi_n_3914, csa_tree_add_12_51_groupi_n_3915, csa_tree_add_12_51_groupi_n_3916, csa_tree_add_12_51_groupi_n_3917, csa_tree_add_12_51_groupi_n_3918, csa_tree_add_12_51_groupi_n_3919, csa_tree_add_12_51_groupi_n_3920;
  wire csa_tree_add_12_51_groupi_n_3921, csa_tree_add_12_51_groupi_n_3922, csa_tree_add_12_51_groupi_n_3923, csa_tree_add_12_51_groupi_n_3924, csa_tree_add_12_51_groupi_n_3925, csa_tree_add_12_51_groupi_n_3926, csa_tree_add_12_51_groupi_n_3927, csa_tree_add_12_51_groupi_n_3928;
  wire csa_tree_add_12_51_groupi_n_3929, csa_tree_add_12_51_groupi_n_3930, csa_tree_add_12_51_groupi_n_3931, csa_tree_add_12_51_groupi_n_3932, csa_tree_add_12_51_groupi_n_3933, csa_tree_add_12_51_groupi_n_3934, csa_tree_add_12_51_groupi_n_3935, csa_tree_add_12_51_groupi_n_3936;
  wire csa_tree_add_12_51_groupi_n_3937, csa_tree_add_12_51_groupi_n_3938, csa_tree_add_12_51_groupi_n_3939, csa_tree_add_12_51_groupi_n_3940, csa_tree_add_12_51_groupi_n_3941, csa_tree_add_12_51_groupi_n_3942, csa_tree_add_12_51_groupi_n_3943, csa_tree_add_12_51_groupi_n_3944;
  wire csa_tree_add_12_51_groupi_n_3945, csa_tree_add_12_51_groupi_n_3946, csa_tree_add_12_51_groupi_n_3947, csa_tree_add_12_51_groupi_n_3948, csa_tree_add_12_51_groupi_n_3949, csa_tree_add_12_51_groupi_n_3950, csa_tree_add_12_51_groupi_n_3951, csa_tree_add_12_51_groupi_n_3952;
  wire csa_tree_add_12_51_groupi_n_3953, csa_tree_add_12_51_groupi_n_3954, csa_tree_add_12_51_groupi_n_3955, csa_tree_add_12_51_groupi_n_3956, csa_tree_add_12_51_groupi_n_3957, csa_tree_add_12_51_groupi_n_3958, csa_tree_add_12_51_groupi_n_3959, csa_tree_add_12_51_groupi_n_3960;
  wire csa_tree_add_12_51_groupi_n_3961, csa_tree_add_12_51_groupi_n_3962, csa_tree_add_12_51_groupi_n_3963, csa_tree_add_12_51_groupi_n_3964, csa_tree_add_12_51_groupi_n_3965, csa_tree_add_12_51_groupi_n_3966, csa_tree_add_12_51_groupi_n_3967, csa_tree_add_12_51_groupi_n_3968;
  wire csa_tree_add_12_51_groupi_n_3969, csa_tree_add_12_51_groupi_n_3970, csa_tree_add_12_51_groupi_n_3971, csa_tree_add_12_51_groupi_n_3972, csa_tree_add_12_51_groupi_n_3973, csa_tree_add_12_51_groupi_n_3974, csa_tree_add_12_51_groupi_n_3975, csa_tree_add_12_51_groupi_n_3976;
  wire csa_tree_add_12_51_groupi_n_3977, csa_tree_add_12_51_groupi_n_3978, csa_tree_add_12_51_groupi_n_3979, csa_tree_add_12_51_groupi_n_3980, csa_tree_add_12_51_groupi_n_3981, csa_tree_add_12_51_groupi_n_3982, csa_tree_add_12_51_groupi_n_3983, csa_tree_add_12_51_groupi_n_3984;
  wire csa_tree_add_12_51_groupi_n_3985, csa_tree_add_12_51_groupi_n_3986, csa_tree_add_12_51_groupi_n_3987, csa_tree_add_12_51_groupi_n_3988, csa_tree_add_12_51_groupi_n_3989, csa_tree_add_12_51_groupi_n_3990, csa_tree_add_12_51_groupi_n_3991, csa_tree_add_12_51_groupi_n_3992;
  wire csa_tree_add_12_51_groupi_n_3993, csa_tree_add_12_51_groupi_n_3994, csa_tree_add_12_51_groupi_n_3995, csa_tree_add_12_51_groupi_n_3996, csa_tree_add_12_51_groupi_n_3997, csa_tree_add_12_51_groupi_n_3998, csa_tree_add_12_51_groupi_n_3999, csa_tree_add_12_51_groupi_n_4000;
  wire csa_tree_add_12_51_groupi_n_4001, csa_tree_add_12_51_groupi_n_4002, csa_tree_add_12_51_groupi_n_4003, csa_tree_add_12_51_groupi_n_4004, csa_tree_add_12_51_groupi_n_4005, csa_tree_add_12_51_groupi_n_4006, csa_tree_add_12_51_groupi_n_4007, csa_tree_add_12_51_groupi_n_4008;
  wire csa_tree_add_12_51_groupi_n_4009, csa_tree_add_12_51_groupi_n_4010, csa_tree_add_12_51_groupi_n_4011, csa_tree_add_12_51_groupi_n_4012, csa_tree_add_12_51_groupi_n_4013, csa_tree_add_12_51_groupi_n_4014, csa_tree_add_12_51_groupi_n_4015, csa_tree_add_12_51_groupi_n_4016;
  wire csa_tree_add_12_51_groupi_n_4017, csa_tree_add_12_51_groupi_n_4018, csa_tree_add_12_51_groupi_n_4019, csa_tree_add_12_51_groupi_n_4020, csa_tree_add_12_51_groupi_n_4021, csa_tree_add_12_51_groupi_n_4022, csa_tree_add_12_51_groupi_n_4023, csa_tree_add_12_51_groupi_n_4024;
  wire csa_tree_add_12_51_groupi_n_4025, csa_tree_add_12_51_groupi_n_4026, csa_tree_add_12_51_groupi_n_4027, csa_tree_add_12_51_groupi_n_4028, csa_tree_add_12_51_groupi_n_4029, csa_tree_add_12_51_groupi_n_4030, csa_tree_add_12_51_groupi_n_4031, csa_tree_add_12_51_groupi_n_4032;
  wire csa_tree_add_12_51_groupi_n_4033, csa_tree_add_12_51_groupi_n_4034, csa_tree_add_12_51_groupi_n_4035, csa_tree_add_12_51_groupi_n_4036, csa_tree_add_12_51_groupi_n_4037, csa_tree_add_12_51_groupi_n_4038, csa_tree_add_12_51_groupi_n_4039, csa_tree_add_12_51_groupi_n_4040;
  wire csa_tree_add_12_51_groupi_n_4041, csa_tree_add_12_51_groupi_n_4042, csa_tree_add_12_51_groupi_n_4043, csa_tree_add_12_51_groupi_n_4044, csa_tree_add_12_51_groupi_n_4045, csa_tree_add_12_51_groupi_n_4046, csa_tree_add_12_51_groupi_n_4047, csa_tree_add_12_51_groupi_n_4048;
  wire csa_tree_add_12_51_groupi_n_4049, csa_tree_add_12_51_groupi_n_4050, csa_tree_add_12_51_groupi_n_4051, csa_tree_add_12_51_groupi_n_4052, csa_tree_add_12_51_groupi_n_4053, csa_tree_add_12_51_groupi_n_4054, csa_tree_add_12_51_groupi_n_4055, csa_tree_add_12_51_groupi_n_4056;
  wire csa_tree_add_12_51_groupi_n_4057, csa_tree_add_12_51_groupi_n_4058, csa_tree_add_12_51_groupi_n_4059, csa_tree_add_12_51_groupi_n_4060, csa_tree_add_12_51_groupi_n_4061, csa_tree_add_12_51_groupi_n_4062, csa_tree_add_12_51_groupi_n_4063, csa_tree_add_12_51_groupi_n_4064;
  wire csa_tree_add_12_51_groupi_n_4065, csa_tree_add_12_51_groupi_n_4066, csa_tree_add_12_51_groupi_n_4067, csa_tree_add_12_51_groupi_n_4068, csa_tree_add_12_51_groupi_n_4069, csa_tree_add_12_51_groupi_n_4070, csa_tree_add_12_51_groupi_n_4071, csa_tree_add_12_51_groupi_n_4072;
  wire csa_tree_add_12_51_groupi_n_4073, csa_tree_add_12_51_groupi_n_4074, csa_tree_add_12_51_groupi_n_4075, csa_tree_add_12_51_groupi_n_4076, csa_tree_add_12_51_groupi_n_4077, csa_tree_add_12_51_groupi_n_4078, csa_tree_add_12_51_groupi_n_4079, csa_tree_add_12_51_groupi_n_4080;
  wire csa_tree_add_12_51_groupi_n_4081, csa_tree_add_12_51_groupi_n_4082, csa_tree_add_12_51_groupi_n_4083, csa_tree_add_12_51_groupi_n_4084, csa_tree_add_12_51_groupi_n_4085, csa_tree_add_12_51_groupi_n_4086, csa_tree_add_12_51_groupi_n_4087, csa_tree_add_12_51_groupi_n_4088;
  wire csa_tree_add_12_51_groupi_n_4089, csa_tree_add_12_51_groupi_n_4090, csa_tree_add_12_51_groupi_n_4091, csa_tree_add_12_51_groupi_n_4092, csa_tree_add_12_51_groupi_n_4093, csa_tree_add_12_51_groupi_n_4094, csa_tree_add_12_51_groupi_n_4095, csa_tree_add_12_51_groupi_n_4096;
  wire csa_tree_add_12_51_groupi_n_4097, csa_tree_add_12_51_groupi_n_4098, csa_tree_add_12_51_groupi_n_4099, csa_tree_add_12_51_groupi_n_4100, csa_tree_add_12_51_groupi_n_4101, csa_tree_add_12_51_groupi_n_4102, csa_tree_add_12_51_groupi_n_4103, csa_tree_add_12_51_groupi_n_4104;
  wire csa_tree_add_12_51_groupi_n_4105, csa_tree_add_12_51_groupi_n_4106, csa_tree_add_12_51_groupi_n_4107, csa_tree_add_12_51_groupi_n_4108, csa_tree_add_12_51_groupi_n_4109, csa_tree_add_12_51_groupi_n_4110, csa_tree_add_12_51_groupi_n_4111, csa_tree_add_12_51_groupi_n_4112;
  wire csa_tree_add_12_51_groupi_n_4113, csa_tree_add_12_51_groupi_n_4114, csa_tree_add_12_51_groupi_n_4115, csa_tree_add_12_51_groupi_n_4116, csa_tree_add_12_51_groupi_n_4117, csa_tree_add_12_51_groupi_n_4118, csa_tree_add_12_51_groupi_n_4119, csa_tree_add_12_51_groupi_n_4120;
  wire csa_tree_add_12_51_groupi_n_4121, csa_tree_add_12_51_groupi_n_4122, csa_tree_add_12_51_groupi_n_4123, csa_tree_add_12_51_groupi_n_4124, csa_tree_add_12_51_groupi_n_4125, csa_tree_add_12_51_groupi_n_4126, csa_tree_add_12_51_groupi_n_4127, csa_tree_add_12_51_groupi_n_4128;
  wire csa_tree_add_12_51_groupi_n_4129, csa_tree_add_12_51_groupi_n_4130, csa_tree_add_12_51_groupi_n_4131, csa_tree_add_12_51_groupi_n_4132, csa_tree_add_12_51_groupi_n_4133, csa_tree_add_12_51_groupi_n_4134, csa_tree_add_12_51_groupi_n_4135, csa_tree_add_12_51_groupi_n_4136;
  wire csa_tree_add_12_51_groupi_n_4137, csa_tree_add_12_51_groupi_n_4138, csa_tree_add_12_51_groupi_n_4139, csa_tree_add_12_51_groupi_n_4140, csa_tree_add_12_51_groupi_n_4141, csa_tree_add_12_51_groupi_n_4142, csa_tree_add_12_51_groupi_n_4143, csa_tree_add_12_51_groupi_n_4144;
  wire csa_tree_add_12_51_groupi_n_4145, csa_tree_add_12_51_groupi_n_4146, csa_tree_add_12_51_groupi_n_4147, csa_tree_add_12_51_groupi_n_4148, csa_tree_add_12_51_groupi_n_4149, csa_tree_add_12_51_groupi_n_4150, csa_tree_add_12_51_groupi_n_4151, csa_tree_add_12_51_groupi_n_4152;
  wire csa_tree_add_12_51_groupi_n_4153, csa_tree_add_12_51_groupi_n_4154, csa_tree_add_12_51_groupi_n_4155, csa_tree_add_12_51_groupi_n_4156, csa_tree_add_12_51_groupi_n_4157, csa_tree_add_12_51_groupi_n_4158, csa_tree_add_12_51_groupi_n_4159, csa_tree_add_12_51_groupi_n_4160;
  wire csa_tree_add_12_51_groupi_n_4161, csa_tree_add_12_51_groupi_n_4162, csa_tree_add_12_51_groupi_n_4163, csa_tree_add_12_51_groupi_n_4164, csa_tree_add_12_51_groupi_n_4165, csa_tree_add_12_51_groupi_n_4166, csa_tree_add_12_51_groupi_n_4167, csa_tree_add_12_51_groupi_n_4168;
  wire csa_tree_add_12_51_groupi_n_4169, csa_tree_add_12_51_groupi_n_4170, csa_tree_add_12_51_groupi_n_4171, csa_tree_add_12_51_groupi_n_4172, csa_tree_add_12_51_groupi_n_4173, csa_tree_add_12_51_groupi_n_4174, csa_tree_add_12_51_groupi_n_4175, csa_tree_add_12_51_groupi_n_4176;
  wire csa_tree_add_12_51_groupi_n_4177, csa_tree_add_12_51_groupi_n_4178, csa_tree_add_12_51_groupi_n_4179, csa_tree_add_12_51_groupi_n_4180, csa_tree_add_12_51_groupi_n_4181, csa_tree_add_12_51_groupi_n_4182, csa_tree_add_12_51_groupi_n_4183, csa_tree_add_12_51_groupi_n_4184;
  wire csa_tree_add_12_51_groupi_n_4185, csa_tree_add_12_51_groupi_n_4186, csa_tree_add_12_51_groupi_n_4187, csa_tree_add_12_51_groupi_n_4188, csa_tree_add_12_51_groupi_n_4189, csa_tree_add_12_51_groupi_n_4190, csa_tree_add_12_51_groupi_n_4191, csa_tree_add_12_51_groupi_n_4192;
  wire csa_tree_add_12_51_groupi_n_4193, csa_tree_add_12_51_groupi_n_4194, csa_tree_add_12_51_groupi_n_4195, csa_tree_add_12_51_groupi_n_4196, csa_tree_add_12_51_groupi_n_4197, csa_tree_add_12_51_groupi_n_4198, csa_tree_add_12_51_groupi_n_4199, csa_tree_add_12_51_groupi_n_4200;
  wire csa_tree_add_12_51_groupi_n_4201, csa_tree_add_12_51_groupi_n_4202, csa_tree_add_12_51_groupi_n_4203, csa_tree_add_12_51_groupi_n_4204, csa_tree_add_12_51_groupi_n_4205, csa_tree_add_12_51_groupi_n_4206, csa_tree_add_12_51_groupi_n_4207, csa_tree_add_12_51_groupi_n_4208;
  wire csa_tree_add_12_51_groupi_n_4209, csa_tree_add_12_51_groupi_n_4210, csa_tree_add_12_51_groupi_n_4211, csa_tree_add_12_51_groupi_n_4212, csa_tree_add_12_51_groupi_n_4213, csa_tree_add_12_51_groupi_n_4214, csa_tree_add_12_51_groupi_n_4215, csa_tree_add_12_51_groupi_n_4216;
  wire csa_tree_add_12_51_groupi_n_4217, csa_tree_add_12_51_groupi_n_4218, csa_tree_add_12_51_groupi_n_4219, csa_tree_add_12_51_groupi_n_4220, csa_tree_add_12_51_groupi_n_4221, csa_tree_add_12_51_groupi_n_4222, csa_tree_add_12_51_groupi_n_4223, csa_tree_add_12_51_groupi_n_4224;
  wire csa_tree_add_12_51_groupi_n_4225, csa_tree_add_12_51_groupi_n_4226, csa_tree_add_12_51_groupi_n_4227, csa_tree_add_12_51_groupi_n_4228, csa_tree_add_12_51_groupi_n_4229, csa_tree_add_12_51_groupi_n_4230, csa_tree_add_12_51_groupi_n_4231, csa_tree_add_12_51_groupi_n_4232;
  wire csa_tree_add_12_51_groupi_n_4233, csa_tree_add_12_51_groupi_n_4234, csa_tree_add_12_51_groupi_n_4235, csa_tree_add_12_51_groupi_n_4236, csa_tree_add_12_51_groupi_n_4237, csa_tree_add_12_51_groupi_n_4238, csa_tree_add_12_51_groupi_n_4239, csa_tree_add_12_51_groupi_n_4240;
  wire csa_tree_add_12_51_groupi_n_4241, csa_tree_add_12_51_groupi_n_4242, csa_tree_add_12_51_groupi_n_4243, csa_tree_add_12_51_groupi_n_4244, csa_tree_add_12_51_groupi_n_4245, csa_tree_add_12_51_groupi_n_4246, csa_tree_add_12_51_groupi_n_4247, csa_tree_add_12_51_groupi_n_4248;
  wire csa_tree_add_12_51_groupi_n_4249, csa_tree_add_12_51_groupi_n_4250, csa_tree_add_12_51_groupi_n_4251, csa_tree_add_12_51_groupi_n_4252, csa_tree_add_12_51_groupi_n_4253, csa_tree_add_12_51_groupi_n_4254, csa_tree_add_12_51_groupi_n_4255, csa_tree_add_12_51_groupi_n_4256;
  wire csa_tree_add_12_51_groupi_n_4257, csa_tree_add_12_51_groupi_n_4258, csa_tree_add_12_51_groupi_n_4259, csa_tree_add_12_51_groupi_n_4260, csa_tree_add_12_51_groupi_n_4261, csa_tree_add_12_51_groupi_n_4262, csa_tree_add_12_51_groupi_n_4263, csa_tree_add_12_51_groupi_n_4264;
  wire csa_tree_add_12_51_groupi_n_4265, csa_tree_add_12_51_groupi_n_4266, csa_tree_add_12_51_groupi_n_4267, csa_tree_add_12_51_groupi_n_4268, csa_tree_add_12_51_groupi_n_4269, csa_tree_add_12_51_groupi_n_4270, csa_tree_add_12_51_groupi_n_4271, csa_tree_add_12_51_groupi_n_4272;
  wire csa_tree_add_12_51_groupi_n_4273, csa_tree_add_12_51_groupi_n_4274, csa_tree_add_12_51_groupi_n_4275, csa_tree_add_12_51_groupi_n_4276, csa_tree_add_12_51_groupi_n_4277, csa_tree_add_12_51_groupi_n_4278, csa_tree_add_12_51_groupi_n_4279, csa_tree_add_12_51_groupi_n_4280;
  wire csa_tree_add_12_51_groupi_n_4281, csa_tree_add_12_51_groupi_n_4282, csa_tree_add_12_51_groupi_n_4283, csa_tree_add_12_51_groupi_n_4284, csa_tree_add_12_51_groupi_n_4285, csa_tree_add_12_51_groupi_n_4286, csa_tree_add_12_51_groupi_n_4287, csa_tree_add_12_51_groupi_n_4288;
  wire csa_tree_add_12_51_groupi_n_4289, csa_tree_add_12_51_groupi_n_4290, csa_tree_add_12_51_groupi_n_4291, csa_tree_add_12_51_groupi_n_4292, csa_tree_add_12_51_groupi_n_4293, csa_tree_add_12_51_groupi_n_4294, csa_tree_add_12_51_groupi_n_4295, csa_tree_add_12_51_groupi_n_4296;
  wire csa_tree_add_12_51_groupi_n_4297, csa_tree_add_12_51_groupi_n_4298, csa_tree_add_12_51_groupi_n_4299, csa_tree_add_12_51_groupi_n_4300, csa_tree_add_12_51_groupi_n_4301, csa_tree_add_12_51_groupi_n_4302, csa_tree_add_12_51_groupi_n_4303, csa_tree_add_12_51_groupi_n_4304;
  wire csa_tree_add_12_51_groupi_n_4305, csa_tree_add_12_51_groupi_n_4306, csa_tree_add_12_51_groupi_n_4307, csa_tree_add_12_51_groupi_n_4308, csa_tree_add_12_51_groupi_n_4309, csa_tree_add_12_51_groupi_n_4310, csa_tree_add_12_51_groupi_n_4311, csa_tree_add_12_51_groupi_n_4312;
  wire csa_tree_add_12_51_groupi_n_4313, csa_tree_add_12_51_groupi_n_4314, csa_tree_add_12_51_groupi_n_4315, csa_tree_add_12_51_groupi_n_4316, csa_tree_add_12_51_groupi_n_4317, csa_tree_add_12_51_groupi_n_4318, csa_tree_add_12_51_groupi_n_4319, csa_tree_add_12_51_groupi_n_4320;
  wire csa_tree_add_12_51_groupi_n_4321, csa_tree_add_12_51_groupi_n_4322, csa_tree_add_12_51_groupi_n_4323, csa_tree_add_12_51_groupi_n_4324, csa_tree_add_12_51_groupi_n_4325, csa_tree_add_12_51_groupi_n_4326, csa_tree_add_12_51_groupi_n_4327, csa_tree_add_12_51_groupi_n_4328;
  wire csa_tree_add_12_51_groupi_n_4329, csa_tree_add_12_51_groupi_n_4330, csa_tree_add_12_51_groupi_n_4331, csa_tree_add_12_51_groupi_n_4332, csa_tree_add_12_51_groupi_n_4333, csa_tree_add_12_51_groupi_n_4334, csa_tree_add_12_51_groupi_n_4335, csa_tree_add_12_51_groupi_n_4336;
  wire csa_tree_add_12_51_groupi_n_4337, csa_tree_add_12_51_groupi_n_4338, csa_tree_add_12_51_groupi_n_4339, csa_tree_add_12_51_groupi_n_4340, csa_tree_add_12_51_groupi_n_4341, csa_tree_add_12_51_groupi_n_4342, csa_tree_add_12_51_groupi_n_4343, csa_tree_add_12_51_groupi_n_4344;
  wire csa_tree_add_12_51_groupi_n_4345, csa_tree_add_12_51_groupi_n_4346, csa_tree_add_12_51_groupi_n_4347, csa_tree_add_12_51_groupi_n_4348, csa_tree_add_12_51_groupi_n_4349, csa_tree_add_12_51_groupi_n_4350, csa_tree_add_12_51_groupi_n_4351, csa_tree_add_12_51_groupi_n_4352;
  wire csa_tree_add_12_51_groupi_n_4353, csa_tree_add_12_51_groupi_n_4354, csa_tree_add_12_51_groupi_n_4355, csa_tree_add_12_51_groupi_n_4356, csa_tree_add_12_51_groupi_n_4357, csa_tree_add_12_51_groupi_n_4358, csa_tree_add_12_51_groupi_n_4359, csa_tree_add_12_51_groupi_n_4360;
  wire csa_tree_add_12_51_groupi_n_4361, csa_tree_add_12_51_groupi_n_4362, csa_tree_add_12_51_groupi_n_4363, csa_tree_add_12_51_groupi_n_4364, csa_tree_add_12_51_groupi_n_4365, csa_tree_add_12_51_groupi_n_4366, csa_tree_add_12_51_groupi_n_4367, csa_tree_add_12_51_groupi_n_4368;
  wire csa_tree_add_12_51_groupi_n_4369, csa_tree_add_12_51_groupi_n_4370, csa_tree_add_12_51_groupi_n_4371, csa_tree_add_12_51_groupi_n_4372, csa_tree_add_12_51_groupi_n_4373, csa_tree_add_12_51_groupi_n_4374, csa_tree_add_12_51_groupi_n_4375, csa_tree_add_12_51_groupi_n_4376;
  wire csa_tree_add_12_51_groupi_n_4377, csa_tree_add_12_51_groupi_n_4378, csa_tree_add_12_51_groupi_n_4379, csa_tree_add_12_51_groupi_n_4380, csa_tree_add_12_51_groupi_n_4381, csa_tree_add_12_51_groupi_n_4382, csa_tree_add_12_51_groupi_n_4383, csa_tree_add_12_51_groupi_n_4384;
  wire csa_tree_add_12_51_groupi_n_4385, csa_tree_add_12_51_groupi_n_4386, csa_tree_add_12_51_groupi_n_4387, csa_tree_add_12_51_groupi_n_4388, csa_tree_add_12_51_groupi_n_4389, csa_tree_add_12_51_groupi_n_4390, csa_tree_add_12_51_groupi_n_4391, csa_tree_add_12_51_groupi_n_4392;
  wire csa_tree_add_12_51_groupi_n_4393, csa_tree_add_12_51_groupi_n_4394, csa_tree_add_12_51_groupi_n_4395, csa_tree_add_12_51_groupi_n_4396, csa_tree_add_12_51_groupi_n_4397, csa_tree_add_12_51_groupi_n_4398, csa_tree_add_12_51_groupi_n_4399, csa_tree_add_12_51_groupi_n_4400;
  wire csa_tree_add_12_51_groupi_n_4401, csa_tree_add_12_51_groupi_n_4402, csa_tree_add_12_51_groupi_n_4403, csa_tree_add_12_51_groupi_n_4404, csa_tree_add_12_51_groupi_n_4405, csa_tree_add_12_51_groupi_n_4406, csa_tree_add_12_51_groupi_n_4407, csa_tree_add_12_51_groupi_n_4408;
  wire csa_tree_add_12_51_groupi_n_4409, csa_tree_add_12_51_groupi_n_4410, csa_tree_add_12_51_groupi_n_4411, csa_tree_add_12_51_groupi_n_4412, csa_tree_add_12_51_groupi_n_4413, csa_tree_add_12_51_groupi_n_4414, csa_tree_add_12_51_groupi_n_4415, csa_tree_add_12_51_groupi_n_4416;
  wire csa_tree_add_12_51_groupi_n_4417, csa_tree_add_12_51_groupi_n_4418, csa_tree_add_12_51_groupi_n_4419, csa_tree_add_12_51_groupi_n_4420, csa_tree_add_12_51_groupi_n_4421, csa_tree_add_12_51_groupi_n_4422, csa_tree_add_12_51_groupi_n_4423, csa_tree_add_12_51_groupi_n_4424;
  wire csa_tree_add_12_51_groupi_n_4425, csa_tree_add_12_51_groupi_n_4426, csa_tree_add_12_51_groupi_n_4427, csa_tree_add_12_51_groupi_n_4428, csa_tree_add_12_51_groupi_n_4429, csa_tree_add_12_51_groupi_n_4430, csa_tree_add_12_51_groupi_n_4431, csa_tree_add_12_51_groupi_n_4432;
  wire csa_tree_add_12_51_groupi_n_4433, csa_tree_add_12_51_groupi_n_4434, csa_tree_add_12_51_groupi_n_4435, csa_tree_add_12_51_groupi_n_4436, csa_tree_add_12_51_groupi_n_4437, csa_tree_add_12_51_groupi_n_4438, csa_tree_add_12_51_groupi_n_4439, csa_tree_add_12_51_groupi_n_4440;
  wire csa_tree_add_12_51_groupi_n_4441, csa_tree_add_12_51_groupi_n_4442, csa_tree_add_12_51_groupi_n_4443, csa_tree_add_12_51_groupi_n_4444, csa_tree_add_12_51_groupi_n_4445, csa_tree_add_12_51_groupi_n_4446, csa_tree_add_12_51_groupi_n_4447, csa_tree_add_12_51_groupi_n_4448;
  wire csa_tree_add_12_51_groupi_n_4449, csa_tree_add_12_51_groupi_n_4450, csa_tree_add_12_51_groupi_n_4451, csa_tree_add_12_51_groupi_n_4452, csa_tree_add_12_51_groupi_n_4453, csa_tree_add_12_51_groupi_n_4454, csa_tree_add_12_51_groupi_n_4455, csa_tree_add_12_51_groupi_n_4456;
  wire csa_tree_add_12_51_groupi_n_4457, csa_tree_add_12_51_groupi_n_4458, csa_tree_add_12_51_groupi_n_4459, csa_tree_add_12_51_groupi_n_4460, csa_tree_add_12_51_groupi_n_4461, csa_tree_add_12_51_groupi_n_4462, csa_tree_add_12_51_groupi_n_4463, csa_tree_add_12_51_groupi_n_4464;
  wire csa_tree_add_12_51_groupi_n_4465, csa_tree_add_12_51_groupi_n_4466, csa_tree_add_12_51_groupi_n_4467, csa_tree_add_12_51_groupi_n_4468, csa_tree_add_12_51_groupi_n_4469, csa_tree_add_12_51_groupi_n_4470, csa_tree_add_12_51_groupi_n_4471, csa_tree_add_12_51_groupi_n_4472;
  wire csa_tree_add_12_51_groupi_n_4473, csa_tree_add_12_51_groupi_n_4474, csa_tree_add_12_51_groupi_n_4475, csa_tree_add_12_51_groupi_n_4476, csa_tree_add_12_51_groupi_n_4477, csa_tree_add_12_51_groupi_n_4478, csa_tree_add_12_51_groupi_n_4479, csa_tree_add_12_51_groupi_n_4480;
  wire csa_tree_add_12_51_groupi_n_4481, csa_tree_add_12_51_groupi_n_4482, csa_tree_add_12_51_groupi_n_4483, csa_tree_add_12_51_groupi_n_4484, csa_tree_add_12_51_groupi_n_4485, csa_tree_add_12_51_groupi_n_4486, csa_tree_add_12_51_groupi_n_4487, csa_tree_add_12_51_groupi_n_4488;
  wire csa_tree_add_12_51_groupi_n_4489, csa_tree_add_12_51_groupi_n_4490, csa_tree_add_12_51_groupi_n_4491, csa_tree_add_12_51_groupi_n_4492, csa_tree_add_12_51_groupi_n_4493, csa_tree_add_12_51_groupi_n_4494, csa_tree_add_12_51_groupi_n_4495, csa_tree_add_12_51_groupi_n_4496;
  wire csa_tree_add_12_51_groupi_n_4497, csa_tree_add_12_51_groupi_n_4498, csa_tree_add_12_51_groupi_n_4499, csa_tree_add_12_51_groupi_n_4500, csa_tree_add_12_51_groupi_n_4501, csa_tree_add_12_51_groupi_n_4502, csa_tree_add_12_51_groupi_n_4503, csa_tree_add_12_51_groupi_n_4504;
  wire csa_tree_add_12_51_groupi_n_4505, csa_tree_add_12_51_groupi_n_4506, csa_tree_add_12_51_groupi_n_4507, csa_tree_add_12_51_groupi_n_4508, csa_tree_add_12_51_groupi_n_4509, csa_tree_add_12_51_groupi_n_4510, csa_tree_add_12_51_groupi_n_4511, csa_tree_add_12_51_groupi_n_4512;
  wire csa_tree_add_12_51_groupi_n_4513, csa_tree_add_12_51_groupi_n_4514, csa_tree_add_12_51_groupi_n_4515, csa_tree_add_12_51_groupi_n_4516, csa_tree_add_12_51_groupi_n_4517, csa_tree_add_12_51_groupi_n_4518, csa_tree_add_12_51_groupi_n_4519, csa_tree_add_12_51_groupi_n_4520;
  wire csa_tree_add_12_51_groupi_n_4521, csa_tree_add_12_51_groupi_n_4522, csa_tree_add_12_51_groupi_n_4523, csa_tree_add_12_51_groupi_n_4524, csa_tree_add_12_51_groupi_n_4525, csa_tree_add_12_51_groupi_n_4526, csa_tree_add_12_51_groupi_n_4527, csa_tree_add_12_51_groupi_n_4528;
  wire csa_tree_add_12_51_groupi_n_4529, csa_tree_add_12_51_groupi_n_4530, csa_tree_add_12_51_groupi_n_4531, csa_tree_add_12_51_groupi_n_4532, csa_tree_add_12_51_groupi_n_4533, csa_tree_add_12_51_groupi_n_4534, csa_tree_add_12_51_groupi_n_4535, csa_tree_add_12_51_groupi_n_4536;
  wire csa_tree_add_12_51_groupi_n_4537, csa_tree_add_12_51_groupi_n_4538, csa_tree_add_12_51_groupi_n_4539, csa_tree_add_12_51_groupi_n_4540, csa_tree_add_12_51_groupi_n_4541, csa_tree_add_12_51_groupi_n_4542, csa_tree_add_12_51_groupi_n_4543, csa_tree_add_12_51_groupi_n_4544;
  wire csa_tree_add_12_51_groupi_n_4545, csa_tree_add_12_51_groupi_n_4546, csa_tree_add_12_51_groupi_n_4547, csa_tree_add_12_51_groupi_n_4548, csa_tree_add_12_51_groupi_n_4549, csa_tree_add_12_51_groupi_n_4550, csa_tree_add_12_51_groupi_n_4551, csa_tree_add_12_51_groupi_n_4552;
  wire csa_tree_add_12_51_groupi_n_4553, csa_tree_add_12_51_groupi_n_4554, csa_tree_add_12_51_groupi_n_4555, csa_tree_add_12_51_groupi_n_4556, csa_tree_add_12_51_groupi_n_4557, csa_tree_add_12_51_groupi_n_4558, csa_tree_add_12_51_groupi_n_4559, csa_tree_add_12_51_groupi_n_4560;
  wire csa_tree_add_12_51_groupi_n_4561, csa_tree_add_12_51_groupi_n_4562, csa_tree_add_12_51_groupi_n_4563, csa_tree_add_12_51_groupi_n_4564, csa_tree_add_12_51_groupi_n_4565, csa_tree_add_12_51_groupi_n_4566, csa_tree_add_12_51_groupi_n_4567, csa_tree_add_12_51_groupi_n_4568;
  wire csa_tree_add_12_51_groupi_n_4569, csa_tree_add_12_51_groupi_n_4570, csa_tree_add_12_51_groupi_n_4571, csa_tree_add_12_51_groupi_n_4572, csa_tree_add_12_51_groupi_n_4573, csa_tree_add_12_51_groupi_n_4574, csa_tree_add_12_51_groupi_n_4575, csa_tree_add_12_51_groupi_n_4576;
  wire csa_tree_add_12_51_groupi_n_4577, csa_tree_add_12_51_groupi_n_4578, csa_tree_add_12_51_groupi_n_4579, csa_tree_add_12_51_groupi_n_4580, csa_tree_add_12_51_groupi_n_4581, csa_tree_add_12_51_groupi_n_4582, csa_tree_add_12_51_groupi_n_4583, csa_tree_add_12_51_groupi_n_4584;
  wire csa_tree_add_12_51_groupi_n_4585, csa_tree_add_12_51_groupi_n_4586, csa_tree_add_12_51_groupi_n_4587, csa_tree_add_12_51_groupi_n_4588, csa_tree_add_12_51_groupi_n_4589, csa_tree_add_12_51_groupi_n_4590, csa_tree_add_12_51_groupi_n_4591, csa_tree_add_12_51_groupi_n_4592;
  wire csa_tree_add_12_51_groupi_n_4593, csa_tree_add_12_51_groupi_n_4594, csa_tree_add_12_51_groupi_n_4595, csa_tree_add_12_51_groupi_n_4596, csa_tree_add_12_51_groupi_n_4597, csa_tree_add_12_51_groupi_n_4598, csa_tree_add_12_51_groupi_n_4599, csa_tree_add_12_51_groupi_n_4600;
  wire csa_tree_add_12_51_groupi_n_4601, csa_tree_add_12_51_groupi_n_4602, csa_tree_add_12_51_groupi_n_4603, csa_tree_add_12_51_groupi_n_4604, csa_tree_add_12_51_groupi_n_4605, csa_tree_add_12_51_groupi_n_4606, csa_tree_add_12_51_groupi_n_4607, csa_tree_add_12_51_groupi_n_4608;
  wire csa_tree_add_12_51_groupi_n_4609, csa_tree_add_12_51_groupi_n_4610, csa_tree_add_12_51_groupi_n_4611, csa_tree_add_12_51_groupi_n_4612, csa_tree_add_12_51_groupi_n_4613, csa_tree_add_12_51_groupi_n_4614, csa_tree_add_12_51_groupi_n_4615, csa_tree_add_12_51_groupi_n_4616;
  wire csa_tree_add_12_51_groupi_n_4617, csa_tree_add_12_51_groupi_n_4618, csa_tree_add_12_51_groupi_n_4619, csa_tree_add_12_51_groupi_n_4620, csa_tree_add_12_51_groupi_n_4621, csa_tree_add_12_51_groupi_n_4622, csa_tree_add_12_51_groupi_n_4623, csa_tree_add_12_51_groupi_n_4624;
  wire csa_tree_add_12_51_groupi_n_4625, csa_tree_add_12_51_groupi_n_4626, csa_tree_add_12_51_groupi_n_4627, csa_tree_add_12_51_groupi_n_4628, csa_tree_add_12_51_groupi_n_4629, csa_tree_add_12_51_groupi_n_4630, csa_tree_add_12_51_groupi_n_4631, csa_tree_add_12_51_groupi_n_4632;
  wire csa_tree_add_12_51_groupi_n_4633, csa_tree_add_12_51_groupi_n_4634, csa_tree_add_12_51_groupi_n_4635, csa_tree_add_12_51_groupi_n_4636, csa_tree_add_12_51_groupi_n_4637, csa_tree_add_12_51_groupi_n_4638, csa_tree_add_12_51_groupi_n_4639, csa_tree_add_12_51_groupi_n_4640;
  wire csa_tree_add_12_51_groupi_n_4641, csa_tree_add_12_51_groupi_n_4642, csa_tree_add_12_51_groupi_n_4643, csa_tree_add_12_51_groupi_n_4644, csa_tree_add_12_51_groupi_n_4645, csa_tree_add_12_51_groupi_n_4646, csa_tree_add_12_51_groupi_n_4647, csa_tree_add_12_51_groupi_n_4648;
  wire csa_tree_add_12_51_groupi_n_4649, csa_tree_add_12_51_groupi_n_4650, csa_tree_add_12_51_groupi_n_4651, csa_tree_add_12_51_groupi_n_4652, csa_tree_add_12_51_groupi_n_4653, csa_tree_add_12_51_groupi_n_4655, csa_tree_add_12_51_groupi_n_4656, csa_tree_add_12_51_groupi_n_4657;
  wire csa_tree_add_12_51_groupi_n_4658, csa_tree_add_12_51_groupi_n_4659, csa_tree_add_12_51_groupi_n_4660, csa_tree_add_12_51_groupi_n_4661, csa_tree_add_12_51_groupi_n_4662, csa_tree_add_12_51_groupi_n_4663, csa_tree_add_12_51_groupi_n_4664, csa_tree_add_12_51_groupi_n_4665;
  wire csa_tree_add_12_51_groupi_n_4666, csa_tree_add_12_51_groupi_n_4667, csa_tree_add_12_51_groupi_n_4668, csa_tree_add_12_51_groupi_n_4669, csa_tree_add_12_51_groupi_n_4670, csa_tree_add_12_51_groupi_n_4671, csa_tree_add_12_51_groupi_n_4672, csa_tree_add_12_51_groupi_n_4673;
  wire csa_tree_add_12_51_groupi_n_4674, csa_tree_add_12_51_groupi_n_4675, csa_tree_add_12_51_groupi_n_4676, csa_tree_add_12_51_groupi_n_4677, csa_tree_add_12_51_groupi_n_4678, csa_tree_add_12_51_groupi_n_4679, csa_tree_add_12_51_groupi_n_4680, csa_tree_add_12_51_groupi_n_4681;
  wire csa_tree_add_12_51_groupi_n_4682, csa_tree_add_12_51_groupi_n_4683, csa_tree_add_12_51_groupi_n_4684, csa_tree_add_12_51_groupi_n_4685, csa_tree_add_12_51_groupi_n_4686, csa_tree_add_12_51_groupi_n_4687, csa_tree_add_12_51_groupi_n_4688, csa_tree_add_12_51_groupi_n_4689;
  wire csa_tree_add_12_51_groupi_n_4690, csa_tree_add_12_51_groupi_n_4691, csa_tree_add_12_51_groupi_n_4692, csa_tree_add_12_51_groupi_n_4693, csa_tree_add_12_51_groupi_n_4694, csa_tree_add_12_51_groupi_n_4695, csa_tree_add_12_51_groupi_n_4696, csa_tree_add_12_51_groupi_n_4697;
  wire csa_tree_add_12_51_groupi_n_4698, csa_tree_add_12_51_groupi_n_4699, csa_tree_add_12_51_groupi_n_4700, csa_tree_add_12_51_groupi_n_4701, csa_tree_add_12_51_groupi_n_4702, csa_tree_add_12_51_groupi_n_4703, csa_tree_add_12_51_groupi_n_4704, csa_tree_add_12_51_groupi_n_4705;
  wire csa_tree_add_12_51_groupi_n_4706, csa_tree_add_12_51_groupi_n_4707, csa_tree_add_12_51_groupi_n_4708, csa_tree_add_12_51_groupi_n_4709, csa_tree_add_12_51_groupi_n_4710, csa_tree_add_12_51_groupi_n_4711, csa_tree_add_12_51_groupi_n_4712, csa_tree_add_12_51_groupi_n_4713;
  wire csa_tree_add_12_51_groupi_n_4714, csa_tree_add_12_51_groupi_n_4715, csa_tree_add_12_51_groupi_n_4716, csa_tree_add_12_51_groupi_n_4717, csa_tree_add_12_51_groupi_n_4718, csa_tree_add_12_51_groupi_n_4719, csa_tree_add_12_51_groupi_n_4720, csa_tree_add_12_51_groupi_n_4721;
  wire csa_tree_add_12_51_groupi_n_4722, csa_tree_add_12_51_groupi_n_4723, csa_tree_add_12_51_groupi_n_4724, csa_tree_add_12_51_groupi_n_4725, csa_tree_add_12_51_groupi_n_4726, csa_tree_add_12_51_groupi_n_4727, csa_tree_add_12_51_groupi_n_4728, csa_tree_add_12_51_groupi_n_4729;
  wire csa_tree_add_12_51_groupi_n_4730, csa_tree_add_12_51_groupi_n_4731, csa_tree_add_12_51_groupi_n_4732, csa_tree_add_12_51_groupi_n_4733, csa_tree_add_12_51_groupi_n_4734, csa_tree_add_12_51_groupi_n_4735, csa_tree_add_12_51_groupi_n_4736, csa_tree_add_12_51_groupi_n_4737;
  wire csa_tree_add_12_51_groupi_n_4738, csa_tree_add_12_51_groupi_n_4739, csa_tree_add_12_51_groupi_n_4740, csa_tree_add_12_51_groupi_n_4741, csa_tree_add_12_51_groupi_n_4742, csa_tree_add_12_51_groupi_n_4743, csa_tree_add_12_51_groupi_n_4744, csa_tree_add_12_51_groupi_n_4745;
  wire csa_tree_add_12_51_groupi_n_4746, csa_tree_add_12_51_groupi_n_4747, csa_tree_add_12_51_groupi_n_4748, csa_tree_add_12_51_groupi_n_4749, csa_tree_add_12_51_groupi_n_4750, csa_tree_add_12_51_groupi_n_4751, csa_tree_add_12_51_groupi_n_4752, csa_tree_add_12_51_groupi_n_4753;
  wire csa_tree_add_12_51_groupi_n_4754, csa_tree_add_12_51_groupi_n_4755, csa_tree_add_12_51_groupi_n_4756, csa_tree_add_12_51_groupi_n_4757, csa_tree_add_12_51_groupi_n_4758, csa_tree_add_12_51_groupi_n_4759, csa_tree_add_12_51_groupi_n_4760, csa_tree_add_12_51_groupi_n_4761;
  wire csa_tree_add_12_51_groupi_n_4762, csa_tree_add_12_51_groupi_n_4763, csa_tree_add_12_51_groupi_n_4764, csa_tree_add_12_51_groupi_n_4765, csa_tree_add_12_51_groupi_n_4766, csa_tree_add_12_51_groupi_n_4767, csa_tree_add_12_51_groupi_n_4768, csa_tree_add_12_51_groupi_n_4769;
  wire csa_tree_add_12_51_groupi_n_4770, csa_tree_add_12_51_groupi_n_4771, csa_tree_add_12_51_groupi_n_4772, csa_tree_add_12_51_groupi_n_4773, csa_tree_add_12_51_groupi_n_4774, csa_tree_add_12_51_groupi_n_4775, csa_tree_add_12_51_groupi_n_4776, csa_tree_add_12_51_groupi_n_4777;
  wire csa_tree_add_12_51_groupi_n_4778, csa_tree_add_12_51_groupi_n_4779, csa_tree_add_12_51_groupi_n_4780, csa_tree_add_12_51_groupi_n_4781, csa_tree_add_12_51_groupi_n_4782, csa_tree_add_12_51_groupi_n_4783, csa_tree_add_12_51_groupi_n_4784, csa_tree_add_12_51_groupi_n_4785;
  wire csa_tree_add_12_51_groupi_n_4786, csa_tree_add_12_51_groupi_n_4787, csa_tree_add_12_51_groupi_n_4788, csa_tree_add_12_51_groupi_n_4789, csa_tree_add_12_51_groupi_n_4790, csa_tree_add_12_51_groupi_n_4791, csa_tree_add_12_51_groupi_n_4792, csa_tree_add_12_51_groupi_n_4793;
  wire csa_tree_add_12_51_groupi_n_4794, csa_tree_add_12_51_groupi_n_4795, csa_tree_add_12_51_groupi_n_4796, csa_tree_add_12_51_groupi_n_4797, csa_tree_add_12_51_groupi_n_4798, csa_tree_add_12_51_groupi_n_4799, csa_tree_add_12_51_groupi_n_4800, csa_tree_add_12_51_groupi_n_4801;
  wire csa_tree_add_12_51_groupi_n_4802, csa_tree_add_12_51_groupi_n_4803, csa_tree_add_12_51_groupi_n_4804, csa_tree_add_12_51_groupi_n_4805, csa_tree_add_12_51_groupi_n_4806, csa_tree_add_12_51_groupi_n_4807, csa_tree_add_12_51_groupi_n_4808, csa_tree_add_12_51_groupi_n_4809;
  wire csa_tree_add_12_51_groupi_n_4810, csa_tree_add_12_51_groupi_n_4811, csa_tree_add_12_51_groupi_n_4812, csa_tree_add_12_51_groupi_n_4813, csa_tree_add_12_51_groupi_n_4814, csa_tree_add_12_51_groupi_n_4815, csa_tree_add_12_51_groupi_n_4816, csa_tree_add_12_51_groupi_n_4817;
  wire csa_tree_add_12_51_groupi_n_4818, csa_tree_add_12_51_groupi_n_4819, csa_tree_add_12_51_groupi_n_4820, csa_tree_add_12_51_groupi_n_4821, csa_tree_add_12_51_groupi_n_4822, csa_tree_add_12_51_groupi_n_4823, csa_tree_add_12_51_groupi_n_4824, csa_tree_add_12_51_groupi_n_4825;
  wire csa_tree_add_12_51_groupi_n_4826, csa_tree_add_12_51_groupi_n_4827, csa_tree_add_12_51_groupi_n_4828, csa_tree_add_12_51_groupi_n_4829, csa_tree_add_12_51_groupi_n_4830, csa_tree_add_12_51_groupi_n_4831, csa_tree_add_12_51_groupi_n_4832, csa_tree_add_12_51_groupi_n_4833;
  wire csa_tree_add_12_51_groupi_n_4834, csa_tree_add_12_51_groupi_n_4835, csa_tree_add_12_51_groupi_n_4836, csa_tree_add_12_51_groupi_n_4837, csa_tree_add_12_51_groupi_n_4838, csa_tree_add_12_51_groupi_n_4839, csa_tree_add_12_51_groupi_n_4840, csa_tree_add_12_51_groupi_n_4841;
  wire csa_tree_add_12_51_groupi_n_4842, csa_tree_add_12_51_groupi_n_4843, csa_tree_add_12_51_groupi_n_4844, csa_tree_add_12_51_groupi_n_4845, csa_tree_add_12_51_groupi_n_4846, csa_tree_add_12_51_groupi_n_4847, csa_tree_add_12_51_groupi_n_4848, csa_tree_add_12_51_groupi_n_4849;
  wire csa_tree_add_12_51_groupi_n_4850, csa_tree_add_12_51_groupi_n_4851, csa_tree_add_12_51_groupi_n_4852, csa_tree_add_12_51_groupi_n_4853, csa_tree_add_12_51_groupi_n_4854, csa_tree_add_12_51_groupi_n_4855, csa_tree_add_12_51_groupi_n_4856, csa_tree_add_12_51_groupi_n_4857;
  wire csa_tree_add_12_51_groupi_n_4858, csa_tree_add_12_51_groupi_n_4859, csa_tree_add_12_51_groupi_n_4860, csa_tree_add_12_51_groupi_n_4861, csa_tree_add_12_51_groupi_n_4862, csa_tree_add_12_51_groupi_n_4863, csa_tree_add_12_51_groupi_n_4864, csa_tree_add_12_51_groupi_n_4865;
  wire csa_tree_add_12_51_groupi_n_4866, csa_tree_add_12_51_groupi_n_4867, csa_tree_add_12_51_groupi_n_4868, csa_tree_add_12_51_groupi_n_4869, csa_tree_add_12_51_groupi_n_4870, csa_tree_add_12_51_groupi_n_4871, csa_tree_add_12_51_groupi_n_4872, csa_tree_add_12_51_groupi_n_4873;
  wire csa_tree_add_12_51_groupi_n_4874, csa_tree_add_12_51_groupi_n_4875, csa_tree_add_12_51_groupi_n_4876, csa_tree_add_12_51_groupi_n_4877, csa_tree_add_12_51_groupi_n_4878, csa_tree_add_12_51_groupi_n_4879, csa_tree_add_12_51_groupi_n_4880, csa_tree_add_12_51_groupi_n_4881;
  wire csa_tree_add_12_51_groupi_n_4882, csa_tree_add_12_51_groupi_n_4883, csa_tree_add_12_51_groupi_n_4884, csa_tree_add_12_51_groupi_n_4885, csa_tree_add_12_51_groupi_n_4886, csa_tree_add_12_51_groupi_n_4887, csa_tree_add_12_51_groupi_n_4888, csa_tree_add_12_51_groupi_n_4889;
  wire csa_tree_add_12_51_groupi_n_4890, csa_tree_add_12_51_groupi_n_4891, csa_tree_add_12_51_groupi_n_4892, csa_tree_add_12_51_groupi_n_4893, csa_tree_add_12_51_groupi_n_4894, csa_tree_add_12_51_groupi_n_4895, csa_tree_add_12_51_groupi_n_4896, csa_tree_add_12_51_groupi_n_4897;
  wire csa_tree_add_12_51_groupi_n_4898, csa_tree_add_12_51_groupi_n_4899, csa_tree_add_12_51_groupi_n_4900, csa_tree_add_12_51_groupi_n_4901, csa_tree_add_12_51_groupi_n_4902, csa_tree_add_12_51_groupi_n_4903, csa_tree_add_12_51_groupi_n_4904, csa_tree_add_12_51_groupi_n_4905;
  wire csa_tree_add_12_51_groupi_n_4906, csa_tree_add_12_51_groupi_n_4907, csa_tree_add_12_51_groupi_n_4908, csa_tree_add_12_51_groupi_n_4909, csa_tree_add_12_51_groupi_n_4910, csa_tree_add_12_51_groupi_n_4911, csa_tree_add_12_51_groupi_n_4912, csa_tree_add_12_51_groupi_n_4913;
  wire csa_tree_add_12_51_groupi_n_4914, csa_tree_add_12_51_groupi_n_4915, csa_tree_add_12_51_groupi_n_4916, csa_tree_add_12_51_groupi_n_4917, csa_tree_add_12_51_groupi_n_4918, csa_tree_add_12_51_groupi_n_4919, csa_tree_add_12_51_groupi_n_4920, csa_tree_add_12_51_groupi_n_4921;
  wire csa_tree_add_12_51_groupi_n_4922, csa_tree_add_12_51_groupi_n_4923, csa_tree_add_12_51_groupi_n_4924, csa_tree_add_12_51_groupi_n_4925, csa_tree_add_12_51_groupi_n_4926, csa_tree_add_12_51_groupi_n_4927, csa_tree_add_12_51_groupi_n_4928, csa_tree_add_12_51_groupi_n_4929;
  wire csa_tree_add_12_51_groupi_n_4930, csa_tree_add_12_51_groupi_n_4931, csa_tree_add_12_51_groupi_n_4932, csa_tree_add_12_51_groupi_n_4933, csa_tree_add_12_51_groupi_n_4934, csa_tree_add_12_51_groupi_n_4935, csa_tree_add_12_51_groupi_n_4936, csa_tree_add_12_51_groupi_n_4937;
  wire csa_tree_add_12_51_groupi_n_4938, csa_tree_add_12_51_groupi_n_4939, csa_tree_add_12_51_groupi_n_4940, csa_tree_add_12_51_groupi_n_4941, csa_tree_add_12_51_groupi_n_4942, csa_tree_add_12_51_groupi_n_4943, csa_tree_add_12_51_groupi_n_4944, csa_tree_add_12_51_groupi_n_4945;
  wire csa_tree_add_12_51_groupi_n_4946, csa_tree_add_12_51_groupi_n_4947, csa_tree_add_12_51_groupi_n_4948, csa_tree_add_12_51_groupi_n_4949, csa_tree_add_12_51_groupi_n_4950, csa_tree_add_12_51_groupi_n_4951, csa_tree_add_12_51_groupi_n_4952, csa_tree_add_12_51_groupi_n_4953;
  wire csa_tree_add_12_51_groupi_n_4954, csa_tree_add_12_51_groupi_n_4955, csa_tree_add_12_51_groupi_n_4956, csa_tree_add_12_51_groupi_n_4957, csa_tree_add_12_51_groupi_n_4958, csa_tree_add_12_51_groupi_n_4959, csa_tree_add_12_51_groupi_n_4960, csa_tree_add_12_51_groupi_n_4961;
  wire csa_tree_add_12_51_groupi_n_4962, csa_tree_add_12_51_groupi_n_4963, csa_tree_add_12_51_groupi_n_4964, csa_tree_add_12_51_groupi_n_4965, csa_tree_add_12_51_groupi_n_4966, csa_tree_add_12_51_groupi_n_4967, csa_tree_add_12_51_groupi_n_4968, csa_tree_add_12_51_groupi_n_4969;
  wire csa_tree_add_12_51_groupi_n_4970, csa_tree_add_12_51_groupi_n_4971, csa_tree_add_12_51_groupi_n_4972, csa_tree_add_12_51_groupi_n_4973, csa_tree_add_12_51_groupi_n_4974, csa_tree_add_12_51_groupi_n_4975, csa_tree_add_12_51_groupi_n_4976, csa_tree_add_12_51_groupi_n_4977;
  wire csa_tree_add_12_51_groupi_n_4978, csa_tree_add_12_51_groupi_n_4979, csa_tree_add_12_51_groupi_n_4980, csa_tree_add_12_51_groupi_n_4981, csa_tree_add_12_51_groupi_n_4982, csa_tree_add_12_51_groupi_n_4983, csa_tree_add_12_51_groupi_n_4984, csa_tree_add_12_51_groupi_n_4985;
  wire csa_tree_add_12_51_groupi_n_4986, csa_tree_add_12_51_groupi_n_4987, csa_tree_add_12_51_groupi_n_4988, csa_tree_add_12_51_groupi_n_4989, csa_tree_add_12_51_groupi_n_4990, csa_tree_add_12_51_groupi_n_4991, csa_tree_add_12_51_groupi_n_4992, csa_tree_add_12_51_groupi_n_4993;
  wire csa_tree_add_12_51_groupi_n_4994, csa_tree_add_12_51_groupi_n_4995, csa_tree_add_12_51_groupi_n_4996, csa_tree_add_12_51_groupi_n_4997, csa_tree_add_12_51_groupi_n_4998, csa_tree_add_12_51_groupi_n_5000, csa_tree_add_12_51_groupi_n_5001, csa_tree_add_12_51_groupi_n_5002;
  wire csa_tree_add_12_51_groupi_n_5003, csa_tree_add_12_51_groupi_n_5004, csa_tree_add_12_51_groupi_n_5005, csa_tree_add_12_51_groupi_n_5006, csa_tree_add_12_51_groupi_n_5007, csa_tree_add_12_51_groupi_n_5008, csa_tree_add_12_51_groupi_n_5009, csa_tree_add_12_51_groupi_n_5010;
  wire csa_tree_add_12_51_groupi_n_5011, csa_tree_add_12_51_groupi_n_5012, csa_tree_add_12_51_groupi_n_5013, csa_tree_add_12_51_groupi_n_5014, csa_tree_add_12_51_groupi_n_5015, csa_tree_add_12_51_groupi_n_5016, csa_tree_add_12_51_groupi_n_5017, csa_tree_add_12_51_groupi_n_5018;
  wire csa_tree_add_12_51_groupi_n_5019, csa_tree_add_12_51_groupi_n_5020, csa_tree_add_12_51_groupi_n_5021, csa_tree_add_12_51_groupi_n_5022, csa_tree_add_12_51_groupi_n_5023, csa_tree_add_12_51_groupi_n_5024, csa_tree_add_12_51_groupi_n_5025, csa_tree_add_12_51_groupi_n_5026;
  wire csa_tree_add_12_51_groupi_n_5027, csa_tree_add_12_51_groupi_n_5028, csa_tree_add_12_51_groupi_n_5029, csa_tree_add_12_51_groupi_n_5030, csa_tree_add_12_51_groupi_n_5031, csa_tree_add_12_51_groupi_n_5032, csa_tree_add_12_51_groupi_n_5033, csa_tree_add_12_51_groupi_n_5034;
  wire csa_tree_add_12_51_groupi_n_5035, csa_tree_add_12_51_groupi_n_5036, csa_tree_add_12_51_groupi_n_5037, csa_tree_add_12_51_groupi_n_5038, csa_tree_add_12_51_groupi_n_5039, csa_tree_add_12_51_groupi_n_5040, csa_tree_add_12_51_groupi_n_5041, csa_tree_add_12_51_groupi_n_5042;
  wire csa_tree_add_12_51_groupi_n_5043, csa_tree_add_12_51_groupi_n_5044, csa_tree_add_12_51_groupi_n_5045, csa_tree_add_12_51_groupi_n_5046, csa_tree_add_12_51_groupi_n_5047, csa_tree_add_12_51_groupi_n_5048, csa_tree_add_12_51_groupi_n_5049, csa_tree_add_12_51_groupi_n_5050;
  wire csa_tree_add_12_51_groupi_n_5051, csa_tree_add_12_51_groupi_n_5052, csa_tree_add_12_51_groupi_n_5053, csa_tree_add_12_51_groupi_n_5054, csa_tree_add_12_51_groupi_n_5055, csa_tree_add_12_51_groupi_n_5056, csa_tree_add_12_51_groupi_n_5057, csa_tree_add_12_51_groupi_n_5058;
  wire csa_tree_add_12_51_groupi_n_5059, csa_tree_add_12_51_groupi_n_5060, csa_tree_add_12_51_groupi_n_5061, csa_tree_add_12_51_groupi_n_5062, csa_tree_add_12_51_groupi_n_5063, csa_tree_add_12_51_groupi_n_5064, csa_tree_add_12_51_groupi_n_5065, csa_tree_add_12_51_groupi_n_5066;
  wire csa_tree_add_12_51_groupi_n_5067, csa_tree_add_12_51_groupi_n_5068, csa_tree_add_12_51_groupi_n_5069, csa_tree_add_12_51_groupi_n_5070, csa_tree_add_12_51_groupi_n_5071, csa_tree_add_12_51_groupi_n_5072, csa_tree_add_12_51_groupi_n_5073, csa_tree_add_12_51_groupi_n_5074;
  wire csa_tree_add_12_51_groupi_n_5075, csa_tree_add_12_51_groupi_n_5076, csa_tree_add_12_51_groupi_n_5077, csa_tree_add_12_51_groupi_n_5078, csa_tree_add_12_51_groupi_n_5079, csa_tree_add_12_51_groupi_n_5080, csa_tree_add_12_51_groupi_n_5081, csa_tree_add_12_51_groupi_n_5082;
  wire csa_tree_add_12_51_groupi_n_5083, csa_tree_add_12_51_groupi_n_5084, csa_tree_add_12_51_groupi_n_5085, csa_tree_add_12_51_groupi_n_5086, csa_tree_add_12_51_groupi_n_5087, csa_tree_add_12_51_groupi_n_5088, csa_tree_add_12_51_groupi_n_5089, csa_tree_add_12_51_groupi_n_5090;
  wire csa_tree_add_12_51_groupi_n_5091, csa_tree_add_12_51_groupi_n_5092, csa_tree_add_12_51_groupi_n_5093, csa_tree_add_12_51_groupi_n_5094, csa_tree_add_12_51_groupi_n_5095, csa_tree_add_12_51_groupi_n_5096, csa_tree_add_12_51_groupi_n_5097, csa_tree_add_12_51_groupi_n_5098;
  wire csa_tree_add_12_51_groupi_n_5099, csa_tree_add_12_51_groupi_n_5100, csa_tree_add_12_51_groupi_n_5101, csa_tree_add_12_51_groupi_n_5102, csa_tree_add_12_51_groupi_n_5103, csa_tree_add_12_51_groupi_n_5104, csa_tree_add_12_51_groupi_n_5105, csa_tree_add_12_51_groupi_n_5106;
  wire csa_tree_add_12_51_groupi_n_5107, csa_tree_add_12_51_groupi_n_5108, csa_tree_add_12_51_groupi_n_5109, csa_tree_add_12_51_groupi_n_5110, csa_tree_add_12_51_groupi_n_5111, csa_tree_add_12_51_groupi_n_5112, csa_tree_add_12_51_groupi_n_5113, csa_tree_add_12_51_groupi_n_5114;
  wire csa_tree_add_12_51_groupi_n_5115, csa_tree_add_12_51_groupi_n_5116, csa_tree_add_12_51_groupi_n_5117, csa_tree_add_12_51_groupi_n_5118, csa_tree_add_12_51_groupi_n_5119, csa_tree_add_12_51_groupi_n_5120, csa_tree_add_12_51_groupi_n_5121, csa_tree_add_12_51_groupi_n_5122;
  wire csa_tree_add_12_51_groupi_n_5123, csa_tree_add_12_51_groupi_n_5124, csa_tree_add_12_51_groupi_n_5125, csa_tree_add_12_51_groupi_n_5126, csa_tree_add_12_51_groupi_n_5127, csa_tree_add_12_51_groupi_n_5128, csa_tree_add_12_51_groupi_n_5129, csa_tree_add_12_51_groupi_n_5130;
  wire csa_tree_add_12_51_groupi_n_5131, csa_tree_add_12_51_groupi_n_5132, csa_tree_add_12_51_groupi_n_5133, csa_tree_add_12_51_groupi_n_5134, csa_tree_add_12_51_groupi_n_5135, csa_tree_add_12_51_groupi_n_5136, csa_tree_add_12_51_groupi_n_5137, csa_tree_add_12_51_groupi_n_5138;
  wire csa_tree_add_12_51_groupi_n_5139, csa_tree_add_12_51_groupi_n_5140, csa_tree_add_12_51_groupi_n_5141, csa_tree_add_12_51_groupi_n_5142, csa_tree_add_12_51_groupi_n_5143, csa_tree_add_12_51_groupi_n_5144, csa_tree_add_12_51_groupi_n_5145, csa_tree_add_12_51_groupi_n_5146;
  wire csa_tree_add_12_51_groupi_n_5147, csa_tree_add_12_51_groupi_n_5148, csa_tree_add_12_51_groupi_n_5149, csa_tree_add_12_51_groupi_n_5150, csa_tree_add_12_51_groupi_n_5151, csa_tree_add_12_51_groupi_n_5152, csa_tree_add_12_51_groupi_n_5153, csa_tree_add_12_51_groupi_n_5154;
  wire csa_tree_add_12_51_groupi_n_5155, csa_tree_add_12_51_groupi_n_5156, csa_tree_add_12_51_groupi_n_5157, csa_tree_add_12_51_groupi_n_5159, csa_tree_add_12_51_groupi_n_5160, csa_tree_add_12_51_groupi_n_5161, csa_tree_add_12_51_groupi_n_5162, csa_tree_add_12_51_groupi_n_5163;
  wire csa_tree_add_12_51_groupi_n_5164, csa_tree_add_12_51_groupi_n_5165, csa_tree_add_12_51_groupi_n_5166, csa_tree_add_12_51_groupi_n_5167, csa_tree_add_12_51_groupi_n_5168, csa_tree_add_12_51_groupi_n_5169, csa_tree_add_12_51_groupi_n_5170, csa_tree_add_12_51_groupi_n_5171;
  wire csa_tree_add_12_51_groupi_n_5172, csa_tree_add_12_51_groupi_n_5173, csa_tree_add_12_51_groupi_n_5174, csa_tree_add_12_51_groupi_n_5175, csa_tree_add_12_51_groupi_n_5176, csa_tree_add_12_51_groupi_n_5177, csa_tree_add_12_51_groupi_n_5178, csa_tree_add_12_51_groupi_n_5179;
  wire csa_tree_add_12_51_groupi_n_5180, csa_tree_add_12_51_groupi_n_5181, csa_tree_add_12_51_groupi_n_5182, csa_tree_add_12_51_groupi_n_5183, csa_tree_add_12_51_groupi_n_5184, csa_tree_add_12_51_groupi_n_5185, csa_tree_add_12_51_groupi_n_5186, csa_tree_add_12_51_groupi_n_5187;
  wire csa_tree_add_12_51_groupi_n_5188, csa_tree_add_12_51_groupi_n_5189, csa_tree_add_12_51_groupi_n_5190, csa_tree_add_12_51_groupi_n_5191, csa_tree_add_12_51_groupi_n_5192, csa_tree_add_12_51_groupi_n_5193, csa_tree_add_12_51_groupi_n_5194, csa_tree_add_12_51_groupi_n_5195;
  wire csa_tree_add_12_51_groupi_n_5196, csa_tree_add_12_51_groupi_n_5197, csa_tree_add_12_51_groupi_n_5198, csa_tree_add_12_51_groupi_n_5199, csa_tree_add_12_51_groupi_n_5200, csa_tree_add_12_51_groupi_n_5201, csa_tree_add_12_51_groupi_n_5202, csa_tree_add_12_51_groupi_n_5203;
  wire csa_tree_add_12_51_groupi_n_5204, csa_tree_add_12_51_groupi_n_5205, csa_tree_add_12_51_groupi_n_5206, csa_tree_add_12_51_groupi_n_5207, csa_tree_add_12_51_groupi_n_5208, csa_tree_add_12_51_groupi_n_5209, csa_tree_add_12_51_groupi_n_5210, csa_tree_add_12_51_groupi_n_5211;
  wire csa_tree_add_12_51_groupi_n_5212, csa_tree_add_12_51_groupi_n_5213, csa_tree_add_12_51_groupi_n_5214, csa_tree_add_12_51_groupi_n_5215, csa_tree_add_12_51_groupi_n_5216, csa_tree_add_12_51_groupi_n_5217, csa_tree_add_12_51_groupi_n_5218, csa_tree_add_12_51_groupi_n_5219;
  wire csa_tree_add_12_51_groupi_n_5220, csa_tree_add_12_51_groupi_n_5221, csa_tree_add_12_51_groupi_n_5222, csa_tree_add_12_51_groupi_n_5223, csa_tree_add_12_51_groupi_n_5224, csa_tree_add_12_51_groupi_n_5225, csa_tree_add_12_51_groupi_n_5226, csa_tree_add_12_51_groupi_n_5227;
  wire csa_tree_add_12_51_groupi_n_5228, csa_tree_add_12_51_groupi_n_5229, csa_tree_add_12_51_groupi_n_5230, csa_tree_add_12_51_groupi_n_5231, csa_tree_add_12_51_groupi_n_5233, csa_tree_add_12_51_groupi_n_5234, csa_tree_add_12_51_groupi_n_5235, csa_tree_add_12_51_groupi_n_5236;
  wire csa_tree_add_12_51_groupi_n_5237, csa_tree_add_12_51_groupi_n_5238, csa_tree_add_12_51_groupi_n_5239, csa_tree_add_12_51_groupi_n_5240, csa_tree_add_12_51_groupi_n_5241, csa_tree_add_12_51_groupi_n_5242, csa_tree_add_12_51_groupi_n_5243, csa_tree_add_12_51_groupi_n_5244;
  wire csa_tree_add_12_51_groupi_n_5245, csa_tree_add_12_51_groupi_n_5246, csa_tree_add_12_51_groupi_n_5247, csa_tree_add_12_51_groupi_n_5248, csa_tree_add_12_51_groupi_n_5249, csa_tree_add_12_51_groupi_n_5250, csa_tree_add_12_51_groupi_n_5251, csa_tree_add_12_51_groupi_n_5252;
  wire csa_tree_add_12_51_groupi_n_5253, csa_tree_add_12_51_groupi_n_5254, csa_tree_add_12_51_groupi_n_5255, csa_tree_add_12_51_groupi_n_5256, csa_tree_add_12_51_groupi_n_5257, csa_tree_add_12_51_groupi_n_5258, csa_tree_add_12_51_groupi_n_5259, csa_tree_add_12_51_groupi_n_5260;
  wire csa_tree_add_12_51_groupi_n_5261, csa_tree_add_12_51_groupi_n_5262, csa_tree_add_12_51_groupi_n_5263, csa_tree_add_12_51_groupi_n_5264, csa_tree_add_12_51_groupi_n_5265, csa_tree_add_12_51_groupi_n_5266, csa_tree_add_12_51_groupi_n_5267, csa_tree_add_12_51_groupi_n_5268;
  wire csa_tree_add_12_51_groupi_n_5269, csa_tree_add_12_51_groupi_n_5270, csa_tree_add_12_51_groupi_n_5271, csa_tree_add_12_51_groupi_n_5272, csa_tree_add_12_51_groupi_n_5273, csa_tree_add_12_51_groupi_n_5274, csa_tree_add_12_51_groupi_n_5275, csa_tree_add_12_51_groupi_n_5276;
  wire csa_tree_add_12_51_groupi_n_5277, csa_tree_add_12_51_groupi_n_5278, csa_tree_add_12_51_groupi_n_5279, csa_tree_add_12_51_groupi_n_5280, csa_tree_add_12_51_groupi_n_5281, csa_tree_add_12_51_groupi_n_5282, csa_tree_add_12_51_groupi_n_5283, csa_tree_add_12_51_groupi_n_5284;
  wire csa_tree_add_12_51_groupi_n_5285, csa_tree_add_12_51_groupi_n_5286, csa_tree_add_12_51_groupi_n_5287, csa_tree_add_12_51_groupi_n_5288, csa_tree_add_12_51_groupi_n_5289, csa_tree_add_12_51_groupi_n_5290, csa_tree_add_12_51_groupi_n_5291, csa_tree_add_12_51_groupi_n_5292;
  wire csa_tree_add_12_51_groupi_n_5293, csa_tree_add_12_51_groupi_n_5294, csa_tree_add_12_51_groupi_n_5295, csa_tree_add_12_51_groupi_n_5296, csa_tree_add_12_51_groupi_n_5297, csa_tree_add_12_51_groupi_n_5298, csa_tree_add_12_51_groupi_n_5299, csa_tree_add_12_51_groupi_n_5300;
  wire csa_tree_add_12_51_groupi_n_5301, csa_tree_add_12_51_groupi_n_5302, csa_tree_add_12_51_groupi_n_5303, csa_tree_add_12_51_groupi_n_5304, csa_tree_add_12_51_groupi_n_5305, csa_tree_add_12_51_groupi_n_5306, csa_tree_add_12_51_groupi_n_5307, csa_tree_add_12_51_groupi_n_5308;
  wire csa_tree_add_12_51_groupi_n_5309, csa_tree_add_12_51_groupi_n_5310, csa_tree_add_12_51_groupi_n_5311, csa_tree_add_12_51_groupi_n_5312, csa_tree_add_12_51_groupi_n_5313, csa_tree_add_12_51_groupi_n_5314, csa_tree_add_12_51_groupi_n_5315, csa_tree_add_12_51_groupi_n_5316;
  wire csa_tree_add_12_51_groupi_n_5317, csa_tree_add_12_51_groupi_n_5318, csa_tree_add_12_51_groupi_n_5319, csa_tree_add_12_51_groupi_n_5320, csa_tree_add_12_51_groupi_n_5321, csa_tree_add_12_51_groupi_n_5322, csa_tree_add_12_51_groupi_n_5323, csa_tree_add_12_51_groupi_n_5324;
  wire csa_tree_add_12_51_groupi_n_5325, csa_tree_add_12_51_groupi_n_5326, csa_tree_add_12_51_groupi_n_5327, csa_tree_add_12_51_groupi_n_5328, csa_tree_add_12_51_groupi_n_5329, csa_tree_add_12_51_groupi_n_5330, csa_tree_add_12_51_groupi_n_5331, csa_tree_add_12_51_groupi_n_5332;
  wire csa_tree_add_12_51_groupi_n_5333, csa_tree_add_12_51_groupi_n_5334, csa_tree_add_12_51_groupi_n_5335, csa_tree_add_12_51_groupi_n_5336, csa_tree_add_12_51_groupi_n_5337, csa_tree_add_12_51_groupi_n_5338, csa_tree_add_12_51_groupi_n_5339, csa_tree_add_12_51_groupi_n_5340;
  wire csa_tree_add_12_51_groupi_n_5341, csa_tree_add_12_51_groupi_n_5342, csa_tree_add_12_51_groupi_n_5343, csa_tree_add_12_51_groupi_n_5344, csa_tree_add_12_51_groupi_n_5345, csa_tree_add_12_51_groupi_n_5346, csa_tree_add_12_51_groupi_n_5347, csa_tree_add_12_51_groupi_n_5348;
  wire csa_tree_add_12_51_groupi_n_5349, csa_tree_add_12_51_groupi_n_5350, csa_tree_add_12_51_groupi_n_5351, csa_tree_add_12_51_groupi_n_5352, csa_tree_add_12_51_groupi_n_5353, csa_tree_add_12_51_groupi_n_5354, csa_tree_add_12_51_groupi_n_5355, csa_tree_add_12_51_groupi_n_5356;
  wire csa_tree_add_12_51_groupi_n_5357, csa_tree_add_12_51_groupi_n_5358, csa_tree_add_12_51_groupi_n_5359, csa_tree_add_12_51_groupi_n_5360, csa_tree_add_12_51_groupi_n_5361, csa_tree_add_12_51_groupi_n_5362, csa_tree_add_12_51_groupi_n_5363, csa_tree_add_12_51_groupi_n_5364;
  wire csa_tree_add_12_51_groupi_n_5365, csa_tree_add_12_51_groupi_n_5366, csa_tree_add_12_51_groupi_n_5367, csa_tree_add_12_51_groupi_n_5368, csa_tree_add_12_51_groupi_n_5369, csa_tree_add_12_51_groupi_n_5370, csa_tree_add_12_51_groupi_n_5371, csa_tree_add_12_51_groupi_n_5372;
  wire csa_tree_add_12_51_groupi_n_5373, csa_tree_add_12_51_groupi_n_5374, csa_tree_add_12_51_groupi_n_5375, csa_tree_add_12_51_groupi_n_5376, csa_tree_add_12_51_groupi_n_5377, csa_tree_add_12_51_groupi_n_5378, csa_tree_add_12_51_groupi_n_5379, csa_tree_add_12_51_groupi_n_5380;
  wire csa_tree_add_12_51_groupi_n_5381, csa_tree_add_12_51_groupi_n_5382, csa_tree_add_12_51_groupi_n_5383, csa_tree_add_12_51_groupi_n_5384, csa_tree_add_12_51_groupi_n_5385, csa_tree_add_12_51_groupi_n_5386, csa_tree_add_12_51_groupi_n_5387, csa_tree_add_12_51_groupi_n_5388;
  wire csa_tree_add_12_51_groupi_n_5389, csa_tree_add_12_51_groupi_n_5390, csa_tree_add_12_51_groupi_n_5391, csa_tree_add_12_51_groupi_n_5392, csa_tree_add_12_51_groupi_n_5393, csa_tree_add_12_51_groupi_n_5394, csa_tree_add_12_51_groupi_n_5395, csa_tree_add_12_51_groupi_n_5396;
  wire csa_tree_add_12_51_groupi_n_5397, csa_tree_add_12_51_groupi_n_5398, csa_tree_add_12_51_groupi_n_5399, csa_tree_add_12_51_groupi_n_5400, csa_tree_add_12_51_groupi_n_5401, csa_tree_add_12_51_groupi_n_5402, csa_tree_add_12_51_groupi_n_5403, csa_tree_add_12_51_groupi_n_5404;
  wire csa_tree_add_12_51_groupi_n_5405, csa_tree_add_12_51_groupi_n_5406, csa_tree_add_12_51_groupi_n_5407, csa_tree_add_12_51_groupi_n_5408, csa_tree_add_12_51_groupi_n_5409, csa_tree_add_12_51_groupi_n_5410, csa_tree_add_12_51_groupi_n_5411, csa_tree_add_12_51_groupi_n_5412;
  wire csa_tree_add_12_51_groupi_n_5413, csa_tree_add_12_51_groupi_n_5414, csa_tree_add_12_51_groupi_n_5415, csa_tree_add_12_51_groupi_n_5416, csa_tree_add_12_51_groupi_n_5417, csa_tree_add_12_51_groupi_n_5418, csa_tree_add_12_51_groupi_n_5419, csa_tree_add_12_51_groupi_n_5420;
  wire csa_tree_add_12_51_groupi_n_5421, csa_tree_add_12_51_groupi_n_5422, csa_tree_add_12_51_groupi_n_5423, csa_tree_add_12_51_groupi_n_5424, csa_tree_add_12_51_groupi_n_5425, csa_tree_add_12_51_groupi_n_5426, csa_tree_add_12_51_groupi_n_5427, csa_tree_add_12_51_groupi_n_5428;
  wire csa_tree_add_12_51_groupi_n_5429, csa_tree_add_12_51_groupi_n_5430, csa_tree_add_12_51_groupi_n_5431, csa_tree_add_12_51_groupi_n_5432, csa_tree_add_12_51_groupi_n_5433, csa_tree_add_12_51_groupi_n_5434, csa_tree_add_12_51_groupi_n_5435, csa_tree_add_12_51_groupi_n_5436;
  wire csa_tree_add_12_51_groupi_n_5437, csa_tree_add_12_51_groupi_n_5438, csa_tree_add_12_51_groupi_n_5439, csa_tree_add_12_51_groupi_n_5440, csa_tree_add_12_51_groupi_n_5441, csa_tree_add_12_51_groupi_n_5442, csa_tree_add_12_51_groupi_n_5443, csa_tree_add_12_51_groupi_n_5444;
  wire csa_tree_add_12_51_groupi_n_5445, csa_tree_add_12_51_groupi_n_5446, csa_tree_add_12_51_groupi_n_5447, csa_tree_add_12_51_groupi_n_5448, csa_tree_add_12_51_groupi_n_5449, csa_tree_add_12_51_groupi_n_5450, csa_tree_add_12_51_groupi_n_5451, csa_tree_add_12_51_groupi_n_5452;
  wire csa_tree_add_12_51_groupi_n_5453, csa_tree_add_12_51_groupi_n_5454, csa_tree_add_12_51_groupi_n_5455, csa_tree_add_12_51_groupi_n_5456, csa_tree_add_12_51_groupi_n_5457, csa_tree_add_12_51_groupi_n_5458, csa_tree_add_12_51_groupi_n_5459, csa_tree_add_12_51_groupi_n_5460;
  wire csa_tree_add_12_51_groupi_n_5461, csa_tree_add_12_51_groupi_n_5462, csa_tree_add_12_51_groupi_n_5463, csa_tree_add_12_51_groupi_n_5464, csa_tree_add_12_51_groupi_n_5465, csa_tree_add_12_51_groupi_n_5466, csa_tree_add_12_51_groupi_n_5467, csa_tree_add_12_51_groupi_n_5468;
  wire csa_tree_add_12_51_groupi_n_5469, csa_tree_add_12_51_groupi_n_5470, csa_tree_add_12_51_groupi_n_5471, csa_tree_add_12_51_groupi_n_5472, csa_tree_add_12_51_groupi_n_5473, csa_tree_add_12_51_groupi_n_5474, csa_tree_add_12_51_groupi_n_5475, csa_tree_add_12_51_groupi_n_5476;
  wire csa_tree_add_12_51_groupi_n_5477, csa_tree_add_12_51_groupi_n_5478, csa_tree_add_12_51_groupi_n_5479, csa_tree_add_12_51_groupi_n_5480, csa_tree_add_12_51_groupi_n_5481, csa_tree_add_12_51_groupi_n_5483, csa_tree_add_12_51_groupi_n_5484, csa_tree_add_12_51_groupi_n_5485;
  wire csa_tree_add_12_51_groupi_n_5486, csa_tree_add_12_51_groupi_n_5487, csa_tree_add_12_51_groupi_n_5488, csa_tree_add_12_51_groupi_n_5489, csa_tree_add_12_51_groupi_n_5490, csa_tree_add_12_51_groupi_n_5491, csa_tree_add_12_51_groupi_n_5492, csa_tree_add_12_51_groupi_n_5493;
  wire csa_tree_add_12_51_groupi_n_5494, csa_tree_add_12_51_groupi_n_5495, csa_tree_add_12_51_groupi_n_5496, csa_tree_add_12_51_groupi_n_5497, csa_tree_add_12_51_groupi_n_5498, csa_tree_add_12_51_groupi_n_5499, csa_tree_add_12_51_groupi_n_5500, csa_tree_add_12_51_groupi_n_5501;
  wire csa_tree_add_12_51_groupi_n_5502, csa_tree_add_12_51_groupi_n_5503, csa_tree_add_12_51_groupi_n_5504, csa_tree_add_12_51_groupi_n_5505, csa_tree_add_12_51_groupi_n_5506, csa_tree_add_12_51_groupi_n_5507, csa_tree_add_12_51_groupi_n_5508, csa_tree_add_12_51_groupi_n_5509;
  wire csa_tree_add_12_51_groupi_n_5510, csa_tree_add_12_51_groupi_n_5511, csa_tree_add_12_51_groupi_n_5512, csa_tree_add_12_51_groupi_n_5513, csa_tree_add_12_51_groupi_n_5514, csa_tree_add_12_51_groupi_n_5515, csa_tree_add_12_51_groupi_n_5516, csa_tree_add_12_51_groupi_n_5517;
  wire csa_tree_add_12_51_groupi_n_5518, csa_tree_add_12_51_groupi_n_5519, csa_tree_add_12_51_groupi_n_5520, csa_tree_add_12_51_groupi_n_5521, csa_tree_add_12_51_groupi_n_5522, csa_tree_add_12_51_groupi_n_5523, csa_tree_add_12_51_groupi_n_5524, csa_tree_add_12_51_groupi_n_5525;
  wire csa_tree_add_12_51_groupi_n_5526, csa_tree_add_12_51_groupi_n_5527, csa_tree_add_12_51_groupi_n_5528, csa_tree_add_12_51_groupi_n_5529, csa_tree_add_12_51_groupi_n_5530, csa_tree_add_12_51_groupi_n_5531, csa_tree_add_12_51_groupi_n_5532, csa_tree_add_12_51_groupi_n_5533;
  wire csa_tree_add_12_51_groupi_n_5534, csa_tree_add_12_51_groupi_n_5535, csa_tree_add_12_51_groupi_n_5536, csa_tree_add_12_51_groupi_n_5537, csa_tree_add_12_51_groupi_n_5538, csa_tree_add_12_51_groupi_n_5539, csa_tree_add_12_51_groupi_n_5540, csa_tree_add_12_51_groupi_n_5541;
  wire csa_tree_add_12_51_groupi_n_5542, csa_tree_add_12_51_groupi_n_5543, csa_tree_add_12_51_groupi_n_5544, csa_tree_add_12_51_groupi_n_5545, csa_tree_add_12_51_groupi_n_5546, csa_tree_add_12_51_groupi_n_5547, csa_tree_add_12_51_groupi_n_5548, csa_tree_add_12_51_groupi_n_5549;
  wire csa_tree_add_12_51_groupi_n_5550, csa_tree_add_12_51_groupi_n_5551, csa_tree_add_12_51_groupi_n_5552, csa_tree_add_12_51_groupi_n_5553, csa_tree_add_12_51_groupi_n_5554, csa_tree_add_12_51_groupi_n_5555, csa_tree_add_12_51_groupi_n_5556, csa_tree_add_12_51_groupi_n_5557;
  wire csa_tree_add_12_51_groupi_n_5558, csa_tree_add_12_51_groupi_n_5559, csa_tree_add_12_51_groupi_n_5560, csa_tree_add_12_51_groupi_n_5561, csa_tree_add_12_51_groupi_n_5562, csa_tree_add_12_51_groupi_n_5563, csa_tree_add_12_51_groupi_n_5564, csa_tree_add_12_51_groupi_n_5565;
  wire csa_tree_add_12_51_groupi_n_5566, csa_tree_add_12_51_groupi_n_5567, csa_tree_add_12_51_groupi_n_5568, csa_tree_add_12_51_groupi_n_5569, csa_tree_add_12_51_groupi_n_5570, csa_tree_add_12_51_groupi_n_5571, csa_tree_add_12_51_groupi_n_5572, csa_tree_add_12_51_groupi_n_5573;
  wire csa_tree_add_12_51_groupi_n_5574, csa_tree_add_12_51_groupi_n_5575, csa_tree_add_12_51_groupi_n_5576, csa_tree_add_12_51_groupi_n_5577, csa_tree_add_12_51_groupi_n_5578, csa_tree_add_12_51_groupi_n_5579, csa_tree_add_12_51_groupi_n_5580, csa_tree_add_12_51_groupi_n_5581;
  wire csa_tree_add_12_51_groupi_n_5582, csa_tree_add_12_51_groupi_n_5583, csa_tree_add_12_51_groupi_n_5584, csa_tree_add_12_51_groupi_n_5585, csa_tree_add_12_51_groupi_n_5586, csa_tree_add_12_51_groupi_n_5587, csa_tree_add_12_51_groupi_n_5588, csa_tree_add_12_51_groupi_n_5589;
  wire csa_tree_add_12_51_groupi_n_5590, csa_tree_add_12_51_groupi_n_5591, csa_tree_add_12_51_groupi_n_5592, csa_tree_add_12_51_groupi_n_5593, csa_tree_add_12_51_groupi_n_5594, csa_tree_add_12_51_groupi_n_5595, csa_tree_add_12_51_groupi_n_5596, csa_tree_add_12_51_groupi_n_5597;
  wire csa_tree_add_12_51_groupi_n_5598, csa_tree_add_12_51_groupi_n_5599, csa_tree_add_12_51_groupi_n_5600, csa_tree_add_12_51_groupi_n_5601, csa_tree_add_12_51_groupi_n_5602, csa_tree_add_12_51_groupi_n_5603, csa_tree_add_12_51_groupi_n_5604, csa_tree_add_12_51_groupi_n_5605;
  wire csa_tree_add_12_51_groupi_n_5606, csa_tree_add_12_51_groupi_n_5607, csa_tree_add_12_51_groupi_n_5608, csa_tree_add_12_51_groupi_n_5609, csa_tree_add_12_51_groupi_n_5610, csa_tree_add_12_51_groupi_n_5611, csa_tree_add_12_51_groupi_n_5612, csa_tree_add_12_51_groupi_n_5613;
  wire csa_tree_add_12_51_groupi_n_5614, csa_tree_add_12_51_groupi_n_5615, csa_tree_add_12_51_groupi_n_5616, csa_tree_add_12_51_groupi_n_5617, csa_tree_add_12_51_groupi_n_5618, csa_tree_add_12_51_groupi_n_5619, csa_tree_add_12_51_groupi_n_5620, csa_tree_add_12_51_groupi_n_5621;
  wire csa_tree_add_12_51_groupi_n_5622, csa_tree_add_12_51_groupi_n_5623, csa_tree_add_12_51_groupi_n_5624, csa_tree_add_12_51_groupi_n_5625, csa_tree_add_12_51_groupi_n_5626, csa_tree_add_12_51_groupi_n_5627, csa_tree_add_12_51_groupi_n_5628, csa_tree_add_12_51_groupi_n_5629;
  wire csa_tree_add_12_51_groupi_n_5630, csa_tree_add_12_51_groupi_n_5631, csa_tree_add_12_51_groupi_n_5632, csa_tree_add_12_51_groupi_n_5633, csa_tree_add_12_51_groupi_n_5634, csa_tree_add_12_51_groupi_n_5635, csa_tree_add_12_51_groupi_n_5636, csa_tree_add_12_51_groupi_n_5637;
  wire csa_tree_add_12_51_groupi_n_5638, csa_tree_add_12_51_groupi_n_5639, csa_tree_add_12_51_groupi_n_5640, csa_tree_add_12_51_groupi_n_5641, csa_tree_add_12_51_groupi_n_5642, csa_tree_add_12_51_groupi_n_5643, csa_tree_add_12_51_groupi_n_5644, csa_tree_add_12_51_groupi_n_5645;
  wire csa_tree_add_12_51_groupi_n_5646, csa_tree_add_12_51_groupi_n_5647, csa_tree_add_12_51_groupi_n_5648, csa_tree_add_12_51_groupi_n_5649, csa_tree_add_12_51_groupi_n_5650, csa_tree_add_12_51_groupi_n_5651, csa_tree_add_12_51_groupi_n_5652, csa_tree_add_12_51_groupi_n_5653;
  wire csa_tree_add_12_51_groupi_n_5654, csa_tree_add_12_51_groupi_n_5655, csa_tree_add_12_51_groupi_n_5656, csa_tree_add_12_51_groupi_n_5657, csa_tree_add_12_51_groupi_n_5658, csa_tree_add_12_51_groupi_n_5659, csa_tree_add_12_51_groupi_n_5660, csa_tree_add_12_51_groupi_n_5661;
  wire csa_tree_add_12_51_groupi_n_5662, csa_tree_add_12_51_groupi_n_5663, csa_tree_add_12_51_groupi_n_5664, csa_tree_add_12_51_groupi_n_5665, csa_tree_add_12_51_groupi_n_5666, csa_tree_add_12_51_groupi_n_5667, csa_tree_add_12_51_groupi_n_5668, csa_tree_add_12_51_groupi_n_5669;
  wire csa_tree_add_12_51_groupi_n_5670, csa_tree_add_12_51_groupi_n_5671, csa_tree_add_12_51_groupi_n_5672, csa_tree_add_12_51_groupi_n_5673, csa_tree_add_12_51_groupi_n_5674, csa_tree_add_12_51_groupi_n_5675, csa_tree_add_12_51_groupi_n_5676, csa_tree_add_12_51_groupi_n_5677;
  wire csa_tree_add_12_51_groupi_n_5678, csa_tree_add_12_51_groupi_n_5679, csa_tree_add_12_51_groupi_n_5680, csa_tree_add_12_51_groupi_n_5681, csa_tree_add_12_51_groupi_n_5682, csa_tree_add_12_51_groupi_n_5683, csa_tree_add_12_51_groupi_n_5684, csa_tree_add_12_51_groupi_n_5685;
  wire csa_tree_add_12_51_groupi_n_5686, csa_tree_add_12_51_groupi_n_5687, csa_tree_add_12_51_groupi_n_5688, csa_tree_add_12_51_groupi_n_5689, csa_tree_add_12_51_groupi_n_5690, csa_tree_add_12_51_groupi_n_5691, csa_tree_add_12_51_groupi_n_5692, csa_tree_add_12_51_groupi_n_5693;
  wire csa_tree_add_12_51_groupi_n_5694, csa_tree_add_12_51_groupi_n_5695, csa_tree_add_12_51_groupi_n_5696, csa_tree_add_12_51_groupi_n_5697, csa_tree_add_12_51_groupi_n_5698, csa_tree_add_12_51_groupi_n_5699, csa_tree_add_12_51_groupi_n_5700, csa_tree_add_12_51_groupi_n_5701;
  wire csa_tree_add_12_51_groupi_n_5702, csa_tree_add_12_51_groupi_n_5703, csa_tree_add_12_51_groupi_n_5704, csa_tree_add_12_51_groupi_n_5705, csa_tree_add_12_51_groupi_n_5706, csa_tree_add_12_51_groupi_n_5707, csa_tree_add_12_51_groupi_n_5708, csa_tree_add_12_51_groupi_n_5709;
  wire csa_tree_add_12_51_groupi_n_5710, csa_tree_add_12_51_groupi_n_5711, csa_tree_add_12_51_groupi_n_5712, csa_tree_add_12_51_groupi_n_5713, csa_tree_add_12_51_groupi_n_5714, csa_tree_add_12_51_groupi_n_5715, csa_tree_add_12_51_groupi_n_5716, csa_tree_add_12_51_groupi_n_5717;
  wire csa_tree_add_12_51_groupi_n_5718, csa_tree_add_12_51_groupi_n_5719, csa_tree_add_12_51_groupi_n_5720, csa_tree_add_12_51_groupi_n_5721, csa_tree_add_12_51_groupi_n_5722, csa_tree_add_12_51_groupi_n_5723, csa_tree_add_12_51_groupi_n_5724, csa_tree_add_12_51_groupi_n_5725;
  wire csa_tree_add_12_51_groupi_n_5726, csa_tree_add_12_51_groupi_n_5727, csa_tree_add_12_51_groupi_n_5728, csa_tree_add_12_51_groupi_n_5729, csa_tree_add_12_51_groupi_n_5731, csa_tree_add_12_51_groupi_n_5732, csa_tree_add_12_51_groupi_n_5733, csa_tree_add_12_51_groupi_n_5734;
  wire csa_tree_add_12_51_groupi_n_5735, csa_tree_add_12_51_groupi_n_5736, csa_tree_add_12_51_groupi_n_5737, csa_tree_add_12_51_groupi_n_5738, csa_tree_add_12_51_groupi_n_5739, csa_tree_add_12_51_groupi_n_5740, csa_tree_add_12_51_groupi_n_5741, csa_tree_add_12_51_groupi_n_5742;
  wire csa_tree_add_12_51_groupi_n_5743, csa_tree_add_12_51_groupi_n_5744, csa_tree_add_12_51_groupi_n_5745, csa_tree_add_12_51_groupi_n_5746, csa_tree_add_12_51_groupi_n_5747, csa_tree_add_12_51_groupi_n_5748, csa_tree_add_12_51_groupi_n_5749, csa_tree_add_12_51_groupi_n_5750;
  wire csa_tree_add_12_51_groupi_n_5751, csa_tree_add_12_51_groupi_n_5752, csa_tree_add_12_51_groupi_n_5753, csa_tree_add_12_51_groupi_n_5754, csa_tree_add_12_51_groupi_n_5755, csa_tree_add_12_51_groupi_n_5756, csa_tree_add_12_51_groupi_n_5757, csa_tree_add_12_51_groupi_n_5758;
  wire csa_tree_add_12_51_groupi_n_5759, csa_tree_add_12_51_groupi_n_5760, csa_tree_add_12_51_groupi_n_5761, csa_tree_add_12_51_groupi_n_5762, csa_tree_add_12_51_groupi_n_5763, csa_tree_add_12_51_groupi_n_5764, csa_tree_add_12_51_groupi_n_5765, csa_tree_add_12_51_groupi_n_5766;
  wire csa_tree_add_12_51_groupi_n_5767, csa_tree_add_12_51_groupi_n_5768, csa_tree_add_12_51_groupi_n_5769, csa_tree_add_12_51_groupi_n_5770, csa_tree_add_12_51_groupi_n_5771, csa_tree_add_12_51_groupi_n_5772, csa_tree_add_12_51_groupi_n_5773, csa_tree_add_12_51_groupi_n_5774;
  wire csa_tree_add_12_51_groupi_n_5775, csa_tree_add_12_51_groupi_n_5776, csa_tree_add_12_51_groupi_n_5777, csa_tree_add_12_51_groupi_n_5778, csa_tree_add_12_51_groupi_n_5779, csa_tree_add_12_51_groupi_n_5780, csa_tree_add_12_51_groupi_n_5781, csa_tree_add_12_51_groupi_n_5782;
  wire csa_tree_add_12_51_groupi_n_5783, csa_tree_add_12_51_groupi_n_5784, csa_tree_add_12_51_groupi_n_5785, csa_tree_add_12_51_groupi_n_5786, csa_tree_add_12_51_groupi_n_5787, csa_tree_add_12_51_groupi_n_5788, csa_tree_add_12_51_groupi_n_5789, csa_tree_add_12_51_groupi_n_5790;
  wire csa_tree_add_12_51_groupi_n_5791, csa_tree_add_12_51_groupi_n_5792, csa_tree_add_12_51_groupi_n_5793, csa_tree_add_12_51_groupi_n_5794, csa_tree_add_12_51_groupi_n_5795, csa_tree_add_12_51_groupi_n_5796, csa_tree_add_12_51_groupi_n_5797, csa_tree_add_12_51_groupi_n_5798;
  wire csa_tree_add_12_51_groupi_n_5799, csa_tree_add_12_51_groupi_n_5800, csa_tree_add_12_51_groupi_n_5801, csa_tree_add_12_51_groupi_n_5802, csa_tree_add_12_51_groupi_n_5803, csa_tree_add_12_51_groupi_n_5804, csa_tree_add_12_51_groupi_n_5805, csa_tree_add_12_51_groupi_n_5806;
  wire csa_tree_add_12_51_groupi_n_5807, csa_tree_add_12_51_groupi_n_5808, csa_tree_add_12_51_groupi_n_5809, csa_tree_add_12_51_groupi_n_5810, csa_tree_add_12_51_groupi_n_5811, csa_tree_add_12_51_groupi_n_5812, csa_tree_add_12_51_groupi_n_5813, csa_tree_add_12_51_groupi_n_5814;
  wire csa_tree_add_12_51_groupi_n_5815, csa_tree_add_12_51_groupi_n_5816, csa_tree_add_12_51_groupi_n_5817, csa_tree_add_12_51_groupi_n_5818, csa_tree_add_12_51_groupi_n_5819, csa_tree_add_12_51_groupi_n_5820, csa_tree_add_12_51_groupi_n_5821, csa_tree_add_12_51_groupi_n_5822;
  wire csa_tree_add_12_51_groupi_n_5823, csa_tree_add_12_51_groupi_n_5824, csa_tree_add_12_51_groupi_n_5825, csa_tree_add_12_51_groupi_n_5826, csa_tree_add_12_51_groupi_n_5827, csa_tree_add_12_51_groupi_n_5828, csa_tree_add_12_51_groupi_n_5829, csa_tree_add_12_51_groupi_n_5830;
  wire csa_tree_add_12_51_groupi_n_5831, csa_tree_add_12_51_groupi_n_5832, csa_tree_add_12_51_groupi_n_5833, csa_tree_add_12_51_groupi_n_5834, csa_tree_add_12_51_groupi_n_5835, csa_tree_add_12_51_groupi_n_5836, csa_tree_add_12_51_groupi_n_5837, csa_tree_add_12_51_groupi_n_5838;
  wire csa_tree_add_12_51_groupi_n_5839, csa_tree_add_12_51_groupi_n_5840, csa_tree_add_12_51_groupi_n_5841, csa_tree_add_12_51_groupi_n_5842, csa_tree_add_12_51_groupi_n_5843, csa_tree_add_12_51_groupi_n_5844, csa_tree_add_12_51_groupi_n_5845, csa_tree_add_12_51_groupi_n_5846;
  wire csa_tree_add_12_51_groupi_n_5847, csa_tree_add_12_51_groupi_n_5848, csa_tree_add_12_51_groupi_n_5849, csa_tree_add_12_51_groupi_n_5850, csa_tree_add_12_51_groupi_n_5851, csa_tree_add_12_51_groupi_n_5852, csa_tree_add_12_51_groupi_n_5853, csa_tree_add_12_51_groupi_n_5854;
  wire csa_tree_add_12_51_groupi_n_5855, csa_tree_add_12_51_groupi_n_5856, csa_tree_add_12_51_groupi_n_5857, csa_tree_add_12_51_groupi_n_5858, csa_tree_add_12_51_groupi_n_5859, csa_tree_add_12_51_groupi_n_5860, csa_tree_add_12_51_groupi_n_5861, csa_tree_add_12_51_groupi_n_5862;
  wire csa_tree_add_12_51_groupi_n_5863, csa_tree_add_12_51_groupi_n_5864, csa_tree_add_12_51_groupi_n_5865, csa_tree_add_12_51_groupi_n_5866, csa_tree_add_12_51_groupi_n_5867, csa_tree_add_12_51_groupi_n_5868, csa_tree_add_12_51_groupi_n_5869, csa_tree_add_12_51_groupi_n_5870;
  wire csa_tree_add_12_51_groupi_n_5871, csa_tree_add_12_51_groupi_n_5872, csa_tree_add_12_51_groupi_n_5873, csa_tree_add_12_51_groupi_n_5874, csa_tree_add_12_51_groupi_n_5875, csa_tree_add_12_51_groupi_n_5876, csa_tree_add_12_51_groupi_n_5877, csa_tree_add_12_51_groupi_n_5878;
  wire csa_tree_add_12_51_groupi_n_5879, csa_tree_add_12_51_groupi_n_5880, csa_tree_add_12_51_groupi_n_5881, csa_tree_add_12_51_groupi_n_5882, csa_tree_add_12_51_groupi_n_5883, csa_tree_add_12_51_groupi_n_5884, csa_tree_add_12_51_groupi_n_5885, csa_tree_add_12_51_groupi_n_5886;
  wire csa_tree_add_12_51_groupi_n_5887, csa_tree_add_12_51_groupi_n_5888, csa_tree_add_12_51_groupi_n_5889, csa_tree_add_12_51_groupi_n_5890, csa_tree_add_12_51_groupi_n_5891, csa_tree_add_12_51_groupi_n_5892, csa_tree_add_12_51_groupi_n_5893, csa_tree_add_12_51_groupi_n_5894;
  wire csa_tree_add_12_51_groupi_n_5895, csa_tree_add_12_51_groupi_n_5896, csa_tree_add_12_51_groupi_n_5897, csa_tree_add_12_51_groupi_n_5898, csa_tree_add_12_51_groupi_n_5900, csa_tree_add_12_51_groupi_n_5901, csa_tree_add_12_51_groupi_n_5902, csa_tree_add_12_51_groupi_n_5903;
  wire csa_tree_add_12_51_groupi_n_5904, csa_tree_add_12_51_groupi_n_5905, csa_tree_add_12_51_groupi_n_5906, csa_tree_add_12_51_groupi_n_5907, csa_tree_add_12_51_groupi_n_5908, csa_tree_add_12_51_groupi_n_5909, csa_tree_add_12_51_groupi_n_5910, csa_tree_add_12_51_groupi_n_5911;
  wire csa_tree_add_12_51_groupi_n_5912, csa_tree_add_12_51_groupi_n_5913, csa_tree_add_12_51_groupi_n_5914, csa_tree_add_12_51_groupi_n_5915, csa_tree_add_12_51_groupi_n_5916, csa_tree_add_12_51_groupi_n_5917, csa_tree_add_12_51_groupi_n_5918, csa_tree_add_12_51_groupi_n_5919;
  wire csa_tree_add_12_51_groupi_n_5920, csa_tree_add_12_51_groupi_n_5921, csa_tree_add_12_51_groupi_n_5922, csa_tree_add_12_51_groupi_n_5923, csa_tree_add_12_51_groupi_n_5924, csa_tree_add_12_51_groupi_n_5925, csa_tree_add_12_51_groupi_n_5926, csa_tree_add_12_51_groupi_n_5927;
  wire csa_tree_add_12_51_groupi_n_5928, csa_tree_add_12_51_groupi_n_5929, csa_tree_add_12_51_groupi_n_5930, csa_tree_add_12_51_groupi_n_5931, csa_tree_add_12_51_groupi_n_5932, csa_tree_add_12_51_groupi_n_5933, csa_tree_add_12_51_groupi_n_5934, csa_tree_add_12_51_groupi_n_5935;
  wire csa_tree_add_12_51_groupi_n_5936, csa_tree_add_12_51_groupi_n_5937, csa_tree_add_12_51_groupi_n_5938, csa_tree_add_12_51_groupi_n_5939, csa_tree_add_12_51_groupi_n_5940, csa_tree_add_12_51_groupi_n_5941, csa_tree_add_12_51_groupi_n_5942, csa_tree_add_12_51_groupi_n_5943;
  wire csa_tree_add_12_51_groupi_n_5944, csa_tree_add_12_51_groupi_n_5945, csa_tree_add_12_51_groupi_n_5946, csa_tree_add_12_51_groupi_n_5947, csa_tree_add_12_51_groupi_n_5948, csa_tree_add_12_51_groupi_n_5949, csa_tree_add_12_51_groupi_n_5950, csa_tree_add_12_51_groupi_n_5951;
  wire csa_tree_add_12_51_groupi_n_5952, csa_tree_add_12_51_groupi_n_5953, csa_tree_add_12_51_groupi_n_5954, csa_tree_add_12_51_groupi_n_5955, csa_tree_add_12_51_groupi_n_5956, csa_tree_add_12_51_groupi_n_5957, csa_tree_add_12_51_groupi_n_5958, csa_tree_add_12_51_groupi_n_5959;
  wire csa_tree_add_12_51_groupi_n_5960, csa_tree_add_12_51_groupi_n_5961, csa_tree_add_12_51_groupi_n_5962, csa_tree_add_12_51_groupi_n_5963, csa_tree_add_12_51_groupi_n_5964, csa_tree_add_12_51_groupi_n_5965, csa_tree_add_12_51_groupi_n_5966, csa_tree_add_12_51_groupi_n_5967;
  wire csa_tree_add_12_51_groupi_n_5968, csa_tree_add_12_51_groupi_n_5969, csa_tree_add_12_51_groupi_n_5970, csa_tree_add_12_51_groupi_n_5971, csa_tree_add_12_51_groupi_n_5972, csa_tree_add_12_51_groupi_n_5973, csa_tree_add_12_51_groupi_n_5974, csa_tree_add_12_51_groupi_n_5975;
  wire csa_tree_add_12_51_groupi_n_5976, csa_tree_add_12_51_groupi_n_5977, csa_tree_add_12_51_groupi_n_5978, csa_tree_add_12_51_groupi_n_5979, csa_tree_add_12_51_groupi_n_5980, csa_tree_add_12_51_groupi_n_5981, csa_tree_add_12_51_groupi_n_5982, csa_tree_add_12_51_groupi_n_5983;
  wire csa_tree_add_12_51_groupi_n_5984, csa_tree_add_12_51_groupi_n_5985, csa_tree_add_12_51_groupi_n_5986, csa_tree_add_12_51_groupi_n_5987, csa_tree_add_12_51_groupi_n_5988, csa_tree_add_12_51_groupi_n_5989, csa_tree_add_12_51_groupi_n_5990, csa_tree_add_12_51_groupi_n_5991;
  wire csa_tree_add_12_51_groupi_n_5992, csa_tree_add_12_51_groupi_n_5993, csa_tree_add_12_51_groupi_n_5994, csa_tree_add_12_51_groupi_n_5995, csa_tree_add_12_51_groupi_n_5996, csa_tree_add_12_51_groupi_n_5997, csa_tree_add_12_51_groupi_n_5998, csa_tree_add_12_51_groupi_n_5999;
  wire csa_tree_add_12_51_groupi_n_6000, csa_tree_add_12_51_groupi_n_6001, csa_tree_add_12_51_groupi_n_6002, csa_tree_add_12_51_groupi_n_6003, csa_tree_add_12_51_groupi_n_6004, csa_tree_add_12_51_groupi_n_6005, csa_tree_add_12_51_groupi_n_6006, csa_tree_add_12_51_groupi_n_6007;
  wire csa_tree_add_12_51_groupi_n_6008, csa_tree_add_12_51_groupi_n_6009, csa_tree_add_12_51_groupi_n_6010, csa_tree_add_12_51_groupi_n_6011, csa_tree_add_12_51_groupi_n_6012, csa_tree_add_12_51_groupi_n_6013, csa_tree_add_12_51_groupi_n_6014, csa_tree_add_12_51_groupi_n_6015;
  wire csa_tree_add_12_51_groupi_n_6016, csa_tree_add_12_51_groupi_n_6017, csa_tree_add_12_51_groupi_n_6018, csa_tree_add_12_51_groupi_n_6019, csa_tree_add_12_51_groupi_n_6020, csa_tree_add_12_51_groupi_n_6021, csa_tree_add_12_51_groupi_n_6022, csa_tree_add_12_51_groupi_n_6023;
  wire csa_tree_add_12_51_groupi_n_6024, csa_tree_add_12_51_groupi_n_6025, csa_tree_add_12_51_groupi_n_6026, csa_tree_add_12_51_groupi_n_6027, csa_tree_add_12_51_groupi_n_6028, csa_tree_add_12_51_groupi_n_6029, csa_tree_add_12_51_groupi_n_6030, csa_tree_add_12_51_groupi_n_6031;
  wire csa_tree_add_12_51_groupi_n_6032, csa_tree_add_12_51_groupi_n_6033, csa_tree_add_12_51_groupi_n_6034, csa_tree_add_12_51_groupi_n_6035, csa_tree_add_12_51_groupi_n_6036, csa_tree_add_12_51_groupi_n_6037, csa_tree_add_12_51_groupi_n_6038, csa_tree_add_12_51_groupi_n_6039;
  wire csa_tree_add_12_51_groupi_n_6040, csa_tree_add_12_51_groupi_n_6041, csa_tree_add_12_51_groupi_n_6042, csa_tree_add_12_51_groupi_n_6043, csa_tree_add_12_51_groupi_n_6044, csa_tree_add_12_51_groupi_n_6045, csa_tree_add_12_51_groupi_n_6046, csa_tree_add_12_51_groupi_n_6047;
  wire csa_tree_add_12_51_groupi_n_6048, csa_tree_add_12_51_groupi_n_6049, csa_tree_add_12_51_groupi_n_6050, csa_tree_add_12_51_groupi_n_6051, csa_tree_add_12_51_groupi_n_6052, csa_tree_add_12_51_groupi_n_6053, csa_tree_add_12_51_groupi_n_6054, csa_tree_add_12_51_groupi_n_6055;
  wire csa_tree_add_12_51_groupi_n_6056, csa_tree_add_12_51_groupi_n_6057, csa_tree_add_12_51_groupi_n_6058, csa_tree_add_12_51_groupi_n_6059, csa_tree_add_12_51_groupi_n_6060, csa_tree_add_12_51_groupi_n_6061, csa_tree_add_12_51_groupi_n_6062, csa_tree_add_12_51_groupi_n_6063;
  wire csa_tree_add_12_51_groupi_n_6064, csa_tree_add_12_51_groupi_n_6065, csa_tree_add_12_51_groupi_n_6066, csa_tree_add_12_51_groupi_n_6067, csa_tree_add_12_51_groupi_n_6068, csa_tree_add_12_51_groupi_n_6069, csa_tree_add_12_51_groupi_n_6070, csa_tree_add_12_51_groupi_n_6071;
  wire csa_tree_add_12_51_groupi_n_6072, csa_tree_add_12_51_groupi_n_6073, csa_tree_add_12_51_groupi_n_6074, csa_tree_add_12_51_groupi_n_6075, csa_tree_add_12_51_groupi_n_6076, csa_tree_add_12_51_groupi_n_6077, csa_tree_add_12_51_groupi_n_6078, csa_tree_add_12_51_groupi_n_6079;
  wire csa_tree_add_12_51_groupi_n_6080, csa_tree_add_12_51_groupi_n_6081, csa_tree_add_12_51_groupi_n_6082, csa_tree_add_12_51_groupi_n_6083, csa_tree_add_12_51_groupi_n_6084, csa_tree_add_12_51_groupi_n_6085, csa_tree_add_12_51_groupi_n_6086, csa_tree_add_12_51_groupi_n_6087;
  wire csa_tree_add_12_51_groupi_n_6088, csa_tree_add_12_51_groupi_n_6089, csa_tree_add_12_51_groupi_n_6090, csa_tree_add_12_51_groupi_n_6091, csa_tree_add_12_51_groupi_n_6092, csa_tree_add_12_51_groupi_n_6093, csa_tree_add_12_51_groupi_n_6094, csa_tree_add_12_51_groupi_n_6095;
  wire csa_tree_add_12_51_groupi_n_6096, csa_tree_add_12_51_groupi_n_6097, csa_tree_add_12_51_groupi_n_6098, csa_tree_add_12_51_groupi_n_6099, csa_tree_add_12_51_groupi_n_6100, csa_tree_add_12_51_groupi_n_6101, csa_tree_add_12_51_groupi_n_6102, csa_tree_add_12_51_groupi_n_6103;
  wire csa_tree_add_12_51_groupi_n_6104, csa_tree_add_12_51_groupi_n_6105, csa_tree_add_12_51_groupi_n_6106, csa_tree_add_12_51_groupi_n_6107, csa_tree_add_12_51_groupi_n_6108, csa_tree_add_12_51_groupi_n_6109, csa_tree_add_12_51_groupi_n_6110, csa_tree_add_12_51_groupi_n_6111;
  wire csa_tree_add_12_51_groupi_n_6112, csa_tree_add_12_51_groupi_n_6113, csa_tree_add_12_51_groupi_n_6114, csa_tree_add_12_51_groupi_n_6115, csa_tree_add_12_51_groupi_n_6116, csa_tree_add_12_51_groupi_n_6117, csa_tree_add_12_51_groupi_n_6118, csa_tree_add_12_51_groupi_n_6119;
  wire csa_tree_add_12_51_groupi_n_6120, csa_tree_add_12_51_groupi_n_6121, csa_tree_add_12_51_groupi_n_6122, csa_tree_add_12_51_groupi_n_6123, csa_tree_add_12_51_groupi_n_6124, csa_tree_add_12_51_groupi_n_6125, csa_tree_add_12_51_groupi_n_6126, csa_tree_add_12_51_groupi_n_6127;
  wire csa_tree_add_12_51_groupi_n_6128, csa_tree_add_12_51_groupi_n_6129, csa_tree_add_12_51_groupi_n_6130, csa_tree_add_12_51_groupi_n_6131, csa_tree_add_12_51_groupi_n_6132, csa_tree_add_12_51_groupi_n_6133, csa_tree_add_12_51_groupi_n_6134, csa_tree_add_12_51_groupi_n_6135;
  wire csa_tree_add_12_51_groupi_n_6136, csa_tree_add_12_51_groupi_n_6137, csa_tree_add_12_51_groupi_n_6138, csa_tree_add_12_51_groupi_n_6139, csa_tree_add_12_51_groupi_n_6140, csa_tree_add_12_51_groupi_n_6141, csa_tree_add_12_51_groupi_n_6142, csa_tree_add_12_51_groupi_n_6143;
  wire csa_tree_add_12_51_groupi_n_6144, csa_tree_add_12_51_groupi_n_6145, csa_tree_add_12_51_groupi_n_6146, csa_tree_add_12_51_groupi_n_6147, csa_tree_add_12_51_groupi_n_6148, csa_tree_add_12_51_groupi_n_6149, csa_tree_add_12_51_groupi_n_6150, csa_tree_add_12_51_groupi_n_6151;
  wire csa_tree_add_12_51_groupi_n_6152, csa_tree_add_12_51_groupi_n_6153, csa_tree_add_12_51_groupi_n_6154, csa_tree_add_12_51_groupi_n_6155, csa_tree_add_12_51_groupi_n_6156, csa_tree_add_12_51_groupi_n_6157, csa_tree_add_12_51_groupi_n_6158, csa_tree_add_12_51_groupi_n_6159;
  wire csa_tree_add_12_51_groupi_n_6160, csa_tree_add_12_51_groupi_n_6161, csa_tree_add_12_51_groupi_n_6162, csa_tree_add_12_51_groupi_n_6163, csa_tree_add_12_51_groupi_n_6164, csa_tree_add_12_51_groupi_n_6165, csa_tree_add_12_51_groupi_n_6166, csa_tree_add_12_51_groupi_n_6167;
  wire csa_tree_add_12_51_groupi_n_6168, csa_tree_add_12_51_groupi_n_6169, csa_tree_add_12_51_groupi_n_6170, csa_tree_add_12_51_groupi_n_6171, csa_tree_add_12_51_groupi_n_6172, csa_tree_add_12_51_groupi_n_6173, csa_tree_add_12_51_groupi_n_6174, csa_tree_add_12_51_groupi_n_6175;
  wire csa_tree_add_12_51_groupi_n_6176, csa_tree_add_12_51_groupi_n_6178, csa_tree_add_12_51_groupi_n_6179, csa_tree_add_12_51_groupi_n_6180, csa_tree_add_12_51_groupi_n_6181, csa_tree_add_12_51_groupi_n_6182, csa_tree_add_12_51_groupi_n_6183, csa_tree_add_12_51_groupi_n_6184;
  wire csa_tree_add_12_51_groupi_n_6185, csa_tree_add_12_51_groupi_n_6186, csa_tree_add_12_51_groupi_n_6187, csa_tree_add_12_51_groupi_n_6188, csa_tree_add_12_51_groupi_n_6189, csa_tree_add_12_51_groupi_n_6190, csa_tree_add_12_51_groupi_n_6191, csa_tree_add_12_51_groupi_n_6192;
  wire csa_tree_add_12_51_groupi_n_6193, csa_tree_add_12_51_groupi_n_6194, csa_tree_add_12_51_groupi_n_6195, csa_tree_add_12_51_groupi_n_6196, csa_tree_add_12_51_groupi_n_6197, csa_tree_add_12_51_groupi_n_6198, csa_tree_add_12_51_groupi_n_6199, csa_tree_add_12_51_groupi_n_6200;
  wire csa_tree_add_12_51_groupi_n_6201, csa_tree_add_12_51_groupi_n_6202, csa_tree_add_12_51_groupi_n_6203, csa_tree_add_12_51_groupi_n_6204, csa_tree_add_12_51_groupi_n_6205, csa_tree_add_12_51_groupi_n_6206, csa_tree_add_12_51_groupi_n_6207, csa_tree_add_12_51_groupi_n_6208;
  wire csa_tree_add_12_51_groupi_n_6209, csa_tree_add_12_51_groupi_n_6210, csa_tree_add_12_51_groupi_n_6211, csa_tree_add_12_51_groupi_n_6212, csa_tree_add_12_51_groupi_n_6213, csa_tree_add_12_51_groupi_n_6214, csa_tree_add_12_51_groupi_n_6215, csa_tree_add_12_51_groupi_n_6216;
  wire csa_tree_add_12_51_groupi_n_6217, csa_tree_add_12_51_groupi_n_6218, csa_tree_add_12_51_groupi_n_6219, csa_tree_add_12_51_groupi_n_6220, csa_tree_add_12_51_groupi_n_6221, csa_tree_add_12_51_groupi_n_6222, csa_tree_add_12_51_groupi_n_6223, csa_tree_add_12_51_groupi_n_6224;
  wire csa_tree_add_12_51_groupi_n_6225, csa_tree_add_12_51_groupi_n_6226, csa_tree_add_12_51_groupi_n_6227, csa_tree_add_12_51_groupi_n_6228, csa_tree_add_12_51_groupi_n_6229, csa_tree_add_12_51_groupi_n_6230, csa_tree_add_12_51_groupi_n_6231, csa_tree_add_12_51_groupi_n_6232;
  wire csa_tree_add_12_51_groupi_n_6233, csa_tree_add_12_51_groupi_n_6234, csa_tree_add_12_51_groupi_n_6235, csa_tree_add_12_51_groupi_n_6236, csa_tree_add_12_51_groupi_n_6237, csa_tree_add_12_51_groupi_n_6238, csa_tree_add_12_51_groupi_n_6239, csa_tree_add_12_51_groupi_n_6240;
  wire csa_tree_add_12_51_groupi_n_6241, csa_tree_add_12_51_groupi_n_6242, csa_tree_add_12_51_groupi_n_6243, csa_tree_add_12_51_groupi_n_6244, csa_tree_add_12_51_groupi_n_6245, csa_tree_add_12_51_groupi_n_6246, csa_tree_add_12_51_groupi_n_6247, csa_tree_add_12_51_groupi_n_6248;
  wire csa_tree_add_12_51_groupi_n_6249, csa_tree_add_12_51_groupi_n_6250, csa_tree_add_12_51_groupi_n_6251, csa_tree_add_12_51_groupi_n_6252, csa_tree_add_12_51_groupi_n_6253, csa_tree_add_12_51_groupi_n_6254, csa_tree_add_12_51_groupi_n_6255, csa_tree_add_12_51_groupi_n_6256;
  wire csa_tree_add_12_51_groupi_n_6257, csa_tree_add_12_51_groupi_n_6258, csa_tree_add_12_51_groupi_n_6259, csa_tree_add_12_51_groupi_n_6260, csa_tree_add_12_51_groupi_n_6261, csa_tree_add_12_51_groupi_n_6262, csa_tree_add_12_51_groupi_n_6263, csa_tree_add_12_51_groupi_n_6264;
  wire csa_tree_add_12_51_groupi_n_6265, csa_tree_add_12_51_groupi_n_6266, csa_tree_add_12_51_groupi_n_6267, csa_tree_add_12_51_groupi_n_6268, csa_tree_add_12_51_groupi_n_6269, csa_tree_add_12_51_groupi_n_6270, csa_tree_add_12_51_groupi_n_6271, csa_tree_add_12_51_groupi_n_6273;
  wire csa_tree_add_12_51_groupi_n_6274, csa_tree_add_12_51_groupi_n_6275, csa_tree_add_12_51_groupi_n_6276, csa_tree_add_12_51_groupi_n_6277, csa_tree_add_12_51_groupi_n_6278, csa_tree_add_12_51_groupi_n_6279, csa_tree_add_12_51_groupi_n_6280, csa_tree_add_12_51_groupi_n_6281;
  wire csa_tree_add_12_51_groupi_n_6282, csa_tree_add_12_51_groupi_n_6283, csa_tree_add_12_51_groupi_n_6284, csa_tree_add_12_51_groupi_n_6285, csa_tree_add_12_51_groupi_n_6286, csa_tree_add_12_51_groupi_n_6287, csa_tree_add_12_51_groupi_n_6288, csa_tree_add_12_51_groupi_n_6289;
  wire csa_tree_add_12_51_groupi_n_6290, csa_tree_add_12_51_groupi_n_6291, csa_tree_add_12_51_groupi_n_6292, csa_tree_add_12_51_groupi_n_6293, csa_tree_add_12_51_groupi_n_6294, csa_tree_add_12_51_groupi_n_6295, csa_tree_add_12_51_groupi_n_6296, csa_tree_add_12_51_groupi_n_6297;
  wire csa_tree_add_12_51_groupi_n_6298, csa_tree_add_12_51_groupi_n_6299, csa_tree_add_12_51_groupi_n_6300, csa_tree_add_12_51_groupi_n_6301, csa_tree_add_12_51_groupi_n_6302, csa_tree_add_12_51_groupi_n_6303, csa_tree_add_12_51_groupi_n_6304, csa_tree_add_12_51_groupi_n_6305;
  wire csa_tree_add_12_51_groupi_n_6306, csa_tree_add_12_51_groupi_n_6307, csa_tree_add_12_51_groupi_n_6308, csa_tree_add_12_51_groupi_n_6309, csa_tree_add_12_51_groupi_n_6310, csa_tree_add_12_51_groupi_n_6311, csa_tree_add_12_51_groupi_n_6312, csa_tree_add_12_51_groupi_n_6313;
  wire csa_tree_add_12_51_groupi_n_6314, csa_tree_add_12_51_groupi_n_6315, csa_tree_add_12_51_groupi_n_6316, csa_tree_add_12_51_groupi_n_6317, csa_tree_add_12_51_groupi_n_6318, csa_tree_add_12_51_groupi_n_6319, csa_tree_add_12_51_groupi_n_6320, csa_tree_add_12_51_groupi_n_6321;
  wire csa_tree_add_12_51_groupi_n_6322, csa_tree_add_12_51_groupi_n_6323, csa_tree_add_12_51_groupi_n_6324, csa_tree_add_12_51_groupi_n_6325, csa_tree_add_12_51_groupi_n_6326, csa_tree_add_12_51_groupi_n_6327, csa_tree_add_12_51_groupi_n_6328, csa_tree_add_12_51_groupi_n_6329;
  wire csa_tree_add_12_51_groupi_n_6330, csa_tree_add_12_51_groupi_n_6331, csa_tree_add_12_51_groupi_n_6332, csa_tree_add_12_51_groupi_n_6333, csa_tree_add_12_51_groupi_n_6334, csa_tree_add_12_51_groupi_n_6335, csa_tree_add_12_51_groupi_n_6336, csa_tree_add_12_51_groupi_n_6337;
  wire csa_tree_add_12_51_groupi_n_6338, csa_tree_add_12_51_groupi_n_6339, csa_tree_add_12_51_groupi_n_6340, csa_tree_add_12_51_groupi_n_6341, csa_tree_add_12_51_groupi_n_6342, csa_tree_add_12_51_groupi_n_6343, csa_tree_add_12_51_groupi_n_6344, csa_tree_add_12_51_groupi_n_6345;
  wire csa_tree_add_12_51_groupi_n_6346, csa_tree_add_12_51_groupi_n_6347, csa_tree_add_12_51_groupi_n_6348, csa_tree_add_12_51_groupi_n_6349, csa_tree_add_12_51_groupi_n_6350, csa_tree_add_12_51_groupi_n_6351, csa_tree_add_12_51_groupi_n_6352, csa_tree_add_12_51_groupi_n_6353;
  wire csa_tree_add_12_51_groupi_n_6354, csa_tree_add_12_51_groupi_n_6355, csa_tree_add_12_51_groupi_n_6356, csa_tree_add_12_51_groupi_n_6357, csa_tree_add_12_51_groupi_n_6358, csa_tree_add_12_51_groupi_n_6359, csa_tree_add_12_51_groupi_n_6360, csa_tree_add_12_51_groupi_n_6361;
  wire csa_tree_add_12_51_groupi_n_6362, csa_tree_add_12_51_groupi_n_6363, csa_tree_add_12_51_groupi_n_6364, csa_tree_add_12_51_groupi_n_6365, csa_tree_add_12_51_groupi_n_6366, csa_tree_add_12_51_groupi_n_6367, csa_tree_add_12_51_groupi_n_6368, csa_tree_add_12_51_groupi_n_6369;
  wire csa_tree_add_12_51_groupi_n_6370, csa_tree_add_12_51_groupi_n_6371, csa_tree_add_12_51_groupi_n_6372, csa_tree_add_12_51_groupi_n_6373, csa_tree_add_12_51_groupi_n_6374, csa_tree_add_12_51_groupi_n_6375, csa_tree_add_12_51_groupi_n_6376, csa_tree_add_12_51_groupi_n_6377;
  wire csa_tree_add_12_51_groupi_n_6378, csa_tree_add_12_51_groupi_n_6379, csa_tree_add_12_51_groupi_n_6380, csa_tree_add_12_51_groupi_n_6381, csa_tree_add_12_51_groupi_n_6382, csa_tree_add_12_51_groupi_n_6383, csa_tree_add_12_51_groupi_n_6384, csa_tree_add_12_51_groupi_n_6385;
  wire csa_tree_add_12_51_groupi_n_6386, csa_tree_add_12_51_groupi_n_6387, csa_tree_add_12_51_groupi_n_6388, csa_tree_add_12_51_groupi_n_6389, csa_tree_add_12_51_groupi_n_6390, csa_tree_add_12_51_groupi_n_6391, csa_tree_add_12_51_groupi_n_6392, csa_tree_add_12_51_groupi_n_6393;
  wire csa_tree_add_12_51_groupi_n_6394, csa_tree_add_12_51_groupi_n_6395, csa_tree_add_12_51_groupi_n_6396, csa_tree_add_12_51_groupi_n_6397, csa_tree_add_12_51_groupi_n_6398, csa_tree_add_12_51_groupi_n_6399, csa_tree_add_12_51_groupi_n_6400, csa_tree_add_12_51_groupi_n_6401;
  wire csa_tree_add_12_51_groupi_n_6402, csa_tree_add_12_51_groupi_n_6403, csa_tree_add_12_51_groupi_n_6404, csa_tree_add_12_51_groupi_n_6405, csa_tree_add_12_51_groupi_n_6406, csa_tree_add_12_51_groupi_n_6407, csa_tree_add_12_51_groupi_n_6408, csa_tree_add_12_51_groupi_n_6409;
  wire csa_tree_add_12_51_groupi_n_6410, csa_tree_add_12_51_groupi_n_6411, csa_tree_add_12_51_groupi_n_6412, csa_tree_add_12_51_groupi_n_6413, csa_tree_add_12_51_groupi_n_6414, csa_tree_add_12_51_groupi_n_6415, csa_tree_add_12_51_groupi_n_6416, csa_tree_add_12_51_groupi_n_6417;
  wire csa_tree_add_12_51_groupi_n_6418, csa_tree_add_12_51_groupi_n_6419, csa_tree_add_12_51_groupi_n_6420, csa_tree_add_12_51_groupi_n_6421, csa_tree_add_12_51_groupi_n_6422, csa_tree_add_12_51_groupi_n_6423, csa_tree_add_12_51_groupi_n_6424, csa_tree_add_12_51_groupi_n_6425;
  wire csa_tree_add_12_51_groupi_n_6426, csa_tree_add_12_51_groupi_n_6427, csa_tree_add_12_51_groupi_n_6428, csa_tree_add_12_51_groupi_n_6429, csa_tree_add_12_51_groupi_n_6430, csa_tree_add_12_51_groupi_n_6431, csa_tree_add_12_51_groupi_n_6432, csa_tree_add_12_51_groupi_n_6433;
  wire csa_tree_add_12_51_groupi_n_6434, csa_tree_add_12_51_groupi_n_6435, csa_tree_add_12_51_groupi_n_6436, csa_tree_add_12_51_groupi_n_6437, csa_tree_add_12_51_groupi_n_6438, csa_tree_add_12_51_groupi_n_6439, csa_tree_add_12_51_groupi_n_6440, csa_tree_add_12_51_groupi_n_6442;
  wire csa_tree_add_12_51_groupi_n_6443, csa_tree_add_12_51_groupi_n_6444, csa_tree_add_12_51_groupi_n_6445, csa_tree_add_12_51_groupi_n_6446, csa_tree_add_12_51_groupi_n_6447, csa_tree_add_12_51_groupi_n_6448, csa_tree_add_12_51_groupi_n_6449, csa_tree_add_12_51_groupi_n_6450;
  wire csa_tree_add_12_51_groupi_n_6451, csa_tree_add_12_51_groupi_n_6452, csa_tree_add_12_51_groupi_n_6453, csa_tree_add_12_51_groupi_n_6454, csa_tree_add_12_51_groupi_n_6455, csa_tree_add_12_51_groupi_n_6456, csa_tree_add_12_51_groupi_n_6457, csa_tree_add_12_51_groupi_n_6458;
  wire csa_tree_add_12_51_groupi_n_6459, csa_tree_add_12_51_groupi_n_6460, csa_tree_add_12_51_groupi_n_6461, csa_tree_add_12_51_groupi_n_6462, csa_tree_add_12_51_groupi_n_6463, csa_tree_add_12_51_groupi_n_6464, csa_tree_add_12_51_groupi_n_6465, csa_tree_add_12_51_groupi_n_6466;
  wire csa_tree_add_12_51_groupi_n_6467, csa_tree_add_12_51_groupi_n_6468, csa_tree_add_12_51_groupi_n_6469, csa_tree_add_12_51_groupi_n_6470, csa_tree_add_12_51_groupi_n_6471, csa_tree_add_12_51_groupi_n_6472, csa_tree_add_12_51_groupi_n_6473, csa_tree_add_12_51_groupi_n_6474;
  wire csa_tree_add_12_51_groupi_n_6475, csa_tree_add_12_51_groupi_n_6476, csa_tree_add_12_51_groupi_n_6477, csa_tree_add_12_51_groupi_n_6478, csa_tree_add_12_51_groupi_n_6479, csa_tree_add_12_51_groupi_n_6480, csa_tree_add_12_51_groupi_n_6481, csa_tree_add_12_51_groupi_n_6482;
  wire csa_tree_add_12_51_groupi_n_6483, csa_tree_add_12_51_groupi_n_6484, csa_tree_add_12_51_groupi_n_6485, csa_tree_add_12_51_groupi_n_6486, csa_tree_add_12_51_groupi_n_6487, csa_tree_add_12_51_groupi_n_6488, csa_tree_add_12_51_groupi_n_6489, csa_tree_add_12_51_groupi_n_6490;
  wire csa_tree_add_12_51_groupi_n_6491, csa_tree_add_12_51_groupi_n_6492, csa_tree_add_12_51_groupi_n_6493, csa_tree_add_12_51_groupi_n_6494, csa_tree_add_12_51_groupi_n_6495, csa_tree_add_12_51_groupi_n_6496, csa_tree_add_12_51_groupi_n_6497, csa_tree_add_12_51_groupi_n_6498;
  wire csa_tree_add_12_51_groupi_n_6499, csa_tree_add_12_51_groupi_n_6500, csa_tree_add_12_51_groupi_n_6501, csa_tree_add_12_51_groupi_n_6502, csa_tree_add_12_51_groupi_n_6503, csa_tree_add_12_51_groupi_n_6504, csa_tree_add_12_51_groupi_n_6505, csa_tree_add_12_51_groupi_n_6506;
  wire csa_tree_add_12_51_groupi_n_6507, csa_tree_add_12_51_groupi_n_6508, csa_tree_add_12_51_groupi_n_6509, csa_tree_add_12_51_groupi_n_6510, csa_tree_add_12_51_groupi_n_6511, csa_tree_add_12_51_groupi_n_6512, csa_tree_add_12_51_groupi_n_6513, csa_tree_add_12_51_groupi_n_6514;
  wire csa_tree_add_12_51_groupi_n_6515, csa_tree_add_12_51_groupi_n_6516, csa_tree_add_12_51_groupi_n_6517, csa_tree_add_12_51_groupi_n_6518, csa_tree_add_12_51_groupi_n_6519, csa_tree_add_12_51_groupi_n_6520, csa_tree_add_12_51_groupi_n_6521, csa_tree_add_12_51_groupi_n_6522;
  wire csa_tree_add_12_51_groupi_n_6523, csa_tree_add_12_51_groupi_n_6524, csa_tree_add_12_51_groupi_n_6525, csa_tree_add_12_51_groupi_n_6526, csa_tree_add_12_51_groupi_n_6527, csa_tree_add_12_51_groupi_n_6528, csa_tree_add_12_51_groupi_n_6529, csa_tree_add_12_51_groupi_n_6530;
  wire csa_tree_add_12_51_groupi_n_6531, csa_tree_add_12_51_groupi_n_6532, csa_tree_add_12_51_groupi_n_6533, csa_tree_add_12_51_groupi_n_6534, csa_tree_add_12_51_groupi_n_6535, csa_tree_add_12_51_groupi_n_6536, csa_tree_add_12_51_groupi_n_6537, csa_tree_add_12_51_groupi_n_6538;
  wire csa_tree_add_12_51_groupi_n_6539, csa_tree_add_12_51_groupi_n_6540, csa_tree_add_12_51_groupi_n_6541, csa_tree_add_12_51_groupi_n_6542, csa_tree_add_12_51_groupi_n_6543, csa_tree_add_12_51_groupi_n_6544, csa_tree_add_12_51_groupi_n_6545, csa_tree_add_12_51_groupi_n_6546;
  wire csa_tree_add_12_51_groupi_n_6547, csa_tree_add_12_51_groupi_n_6548, csa_tree_add_12_51_groupi_n_6549, csa_tree_add_12_51_groupi_n_6550, csa_tree_add_12_51_groupi_n_6551, csa_tree_add_12_51_groupi_n_6552, csa_tree_add_12_51_groupi_n_6553, csa_tree_add_12_51_groupi_n_6554;
  wire csa_tree_add_12_51_groupi_n_6555, csa_tree_add_12_51_groupi_n_6556, csa_tree_add_12_51_groupi_n_6557, csa_tree_add_12_51_groupi_n_6558, csa_tree_add_12_51_groupi_n_6559, csa_tree_add_12_51_groupi_n_6560, csa_tree_add_12_51_groupi_n_6561, csa_tree_add_12_51_groupi_n_6562;
  wire csa_tree_add_12_51_groupi_n_6563, csa_tree_add_12_51_groupi_n_6564, csa_tree_add_12_51_groupi_n_6565, csa_tree_add_12_51_groupi_n_6566, csa_tree_add_12_51_groupi_n_6567, csa_tree_add_12_51_groupi_n_6568, csa_tree_add_12_51_groupi_n_6569, csa_tree_add_12_51_groupi_n_6570;
  wire csa_tree_add_12_51_groupi_n_6571, csa_tree_add_12_51_groupi_n_6572, csa_tree_add_12_51_groupi_n_6573, csa_tree_add_12_51_groupi_n_6574, csa_tree_add_12_51_groupi_n_6575, csa_tree_add_12_51_groupi_n_6576, csa_tree_add_12_51_groupi_n_6577, csa_tree_add_12_51_groupi_n_6578;
  wire csa_tree_add_12_51_groupi_n_6579, csa_tree_add_12_51_groupi_n_6580, csa_tree_add_12_51_groupi_n_6581, csa_tree_add_12_51_groupi_n_6582, csa_tree_add_12_51_groupi_n_6583, csa_tree_add_12_51_groupi_n_6584, csa_tree_add_12_51_groupi_n_6585, csa_tree_add_12_51_groupi_n_6586;
  wire csa_tree_add_12_51_groupi_n_6587, csa_tree_add_12_51_groupi_n_6588, csa_tree_add_12_51_groupi_n_6589, csa_tree_add_12_51_groupi_n_6590, csa_tree_add_12_51_groupi_n_6591, csa_tree_add_12_51_groupi_n_6592, csa_tree_add_12_51_groupi_n_6593, csa_tree_add_12_51_groupi_n_6594;
  wire csa_tree_add_12_51_groupi_n_6595, csa_tree_add_12_51_groupi_n_6596, csa_tree_add_12_51_groupi_n_6597, csa_tree_add_12_51_groupi_n_6598, csa_tree_add_12_51_groupi_n_6599, csa_tree_add_12_51_groupi_n_6600, csa_tree_add_12_51_groupi_n_6601, csa_tree_add_12_51_groupi_n_6602;
  wire csa_tree_add_12_51_groupi_n_6603, csa_tree_add_12_51_groupi_n_6604, csa_tree_add_12_51_groupi_n_6605, csa_tree_add_12_51_groupi_n_6606, csa_tree_add_12_51_groupi_n_6607, csa_tree_add_12_51_groupi_n_6608, csa_tree_add_12_51_groupi_n_6609, csa_tree_add_12_51_groupi_n_6610;
  wire csa_tree_add_12_51_groupi_n_6611, csa_tree_add_12_51_groupi_n_6612, csa_tree_add_12_51_groupi_n_6613, csa_tree_add_12_51_groupi_n_6614, csa_tree_add_12_51_groupi_n_6615, csa_tree_add_12_51_groupi_n_6616, csa_tree_add_12_51_groupi_n_6617, csa_tree_add_12_51_groupi_n_6618;
  wire csa_tree_add_12_51_groupi_n_6619, csa_tree_add_12_51_groupi_n_6621, csa_tree_add_12_51_groupi_n_6622, csa_tree_add_12_51_groupi_n_6623, csa_tree_add_12_51_groupi_n_6624, csa_tree_add_12_51_groupi_n_6625, csa_tree_add_12_51_groupi_n_6626, csa_tree_add_12_51_groupi_n_6627;
  wire csa_tree_add_12_51_groupi_n_6628, csa_tree_add_12_51_groupi_n_6629, csa_tree_add_12_51_groupi_n_6630, csa_tree_add_12_51_groupi_n_6631, csa_tree_add_12_51_groupi_n_6632, csa_tree_add_12_51_groupi_n_6633, csa_tree_add_12_51_groupi_n_6634, csa_tree_add_12_51_groupi_n_6635;
  wire csa_tree_add_12_51_groupi_n_6636, csa_tree_add_12_51_groupi_n_6637, csa_tree_add_12_51_groupi_n_6638, csa_tree_add_12_51_groupi_n_6639, csa_tree_add_12_51_groupi_n_6640, csa_tree_add_12_51_groupi_n_6641, csa_tree_add_12_51_groupi_n_6642, csa_tree_add_12_51_groupi_n_6643;
  wire csa_tree_add_12_51_groupi_n_6644, csa_tree_add_12_51_groupi_n_6645, csa_tree_add_12_51_groupi_n_6646, csa_tree_add_12_51_groupi_n_6647, csa_tree_add_12_51_groupi_n_6648, csa_tree_add_12_51_groupi_n_6649, csa_tree_add_12_51_groupi_n_6650, csa_tree_add_12_51_groupi_n_6651;
  wire csa_tree_add_12_51_groupi_n_6652, csa_tree_add_12_51_groupi_n_6653, csa_tree_add_12_51_groupi_n_6654, csa_tree_add_12_51_groupi_n_6655, csa_tree_add_12_51_groupi_n_6656, csa_tree_add_12_51_groupi_n_6657, csa_tree_add_12_51_groupi_n_6658, csa_tree_add_12_51_groupi_n_6659;
  wire csa_tree_add_12_51_groupi_n_6660, csa_tree_add_12_51_groupi_n_6661, csa_tree_add_12_51_groupi_n_6662, csa_tree_add_12_51_groupi_n_6663, csa_tree_add_12_51_groupi_n_6664, csa_tree_add_12_51_groupi_n_6665, csa_tree_add_12_51_groupi_n_6666, csa_tree_add_12_51_groupi_n_6667;
  wire csa_tree_add_12_51_groupi_n_6668, csa_tree_add_12_51_groupi_n_6669, csa_tree_add_12_51_groupi_n_6670, csa_tree_add_12_51_groupi_n_6671, csa_tree_add_12_51_groupi_n_6672, csa_tree_add_12_51_groupi_n_6673, csa_tree_add_12_51_groupi_n_6674, csa_tree_add_12_51_groupi_n_6675;
  wire csa_tree_add_12_51_groupi_n_6676, csa_tree_add_12_51_groupi_n_6677, csa_tree_add_12_51_groupi_n_6678, csa_tree_add_12_51_groupi_n_6679, csa_tree_add_12_51_groupi_n_6680, csa_tree_add_12_51_groupi_n_6681, csa_tree_add_12_51_groupi_n_6682, csa_tree_add_12_51_groupi_n_6683;
  wire csa_tree_add_12_51_groupi_n_6684, csa_tree_add_12_51_groupi_n_6685, csa_tree_add_12_51_groupi_n_6686, csa_tree_add_12_51_groupi_n_6687, csa_tree_add_12_51_groupi_n_6688, csa_tree_add_12_51_groupi_n_6689, csa_tree_add_12_51_groupi_n_6690, csa_tree_add_12_51_groupi_n_6691;
  wire csa_tree_add_12_51_groupi_n_6692, csa_tree_add_12_51_groupi_n_6693, csa_tree_add_12_51_groupi_n_6694, csa_tree_add_12_51_groupi_n_6695, csa_tree_add_12_51_groupi_n_6696, csa_tree_add_12_51_groupi_n_6697, csa_tree_add_12_51_groupi_n_6698, csa_tree_add_12_51_groupi_n_6699;
  wire csa_tree_add_12_51_groupi_n_6700, csa_tree_add_12_51_groupi_n_6701, csa_tree_add_12_51_groupi_n_6702, csa_tree_add_12_51_groupi_n_6703, csa_tree_add_12_51_groupi_n_6704, csa_tree_add_12_51_groupi_n_6705, csa_tree_add_12_51_groupi_n_6706, csa_tree_add_12_51_groupi_n_6707;
  wire csa_tree_add_12_51_groupi_n_6708, csa_tree_add_12_51_groupi_n_6709, csa_tree_add_12_51_groupi_n_6710, csa_tree_add_12_51_groupi_n_6711, csa_tree_add_12_51_groupi_n_6712, csa_tree_add_12_51_groupi_n_6713, csa_tree_add_12_51_groupi_n_6714, csa_tree_add_12_51_groupi_n_6715;
  wire csa_tree_add_12_51_groupi_n_6716, csa_tree_add_12_51_groupi_n_6717, csa_tree_add_12_51_groupi_n_6718, csa_tree_add_12_51_groupi_n_6719, csa_tree_add_12_51_groupi_n_6720, csa_tree_add_12_51_groupi_n_6721, csa_tree_add_12_51_groupi_n_6722, csa_tree_add_12_51_groupi_n_6723;
  wire csa_tree_add_12_51_groupi_n_6724, csa_tree_add_12_51_groupi_n_6725, csa_tree_add_12_51_groupi_n_6726, csa_tree_add_12_51_groupi_n_6727, csa_tree_add_12_51_groupi_n_6728, csa_tree_add_12_51_groupi_n_6729, csa_tree_add_12_51_groupi_n_6730, csa_tree_add_12_51_groupi_n_6731;
  wire csa_tree_add_12_51_groupi_n_6732, csa_tree_add_12_51_groupi_n_6733, csa_tree_add_12_51_groupi_n_6734, csa_tree_add_12_51_groupi_n_6735, csa_tree_add_12_51_groupi_n_6736, csa_tree_add_12_51_groupi_n_6737, csa_tree_add_12_51_groupi_n_6739, csa_tree_add_12_51_groupi_n_6740;
  wire csa_tree_add_12_51_groupi_n_6741, csa_tree_add_12_51_groupi_n_6742, csa_tree_add_12_51_groupi_n_6743, csa_tree_add_12_51_groupi_n_6744, csa_tree_add_12_51_groupi_n_6745, csa_tree_add_12_51_groupi_n_6746, csa_tree_add_12_51_groupi_n_6747, csa_tree_add_12_51_groupi_n_6748;
  wire csa_tree_add_12_51_groupi_n_6749, csa_tree_add_12_51_groupi_n_6750, csa_tree_add_12_51_groupi_n_6751, csa_tree_add_12_51_groupi_n_6752, csa_tree_add_12_51_groupi_n_6753, csa_tree_add_12_51_groupi_n_6754, csa_tree_add_12_51_groupi_n_6755, csa_tree_add_12_51_groupi_n_6756;
  wire csa_tree_add_12_51_groupi_n_6757, csa_tree_add_12_51_groupi_n_6758, csa_tree_add_12_51_groupi_n_6759, csa_tree_add_12_51_groupi_n_6760, csa_tree_add_12_51_groupi_n_6761, csa_tree_add_12_51_groupi_n_6762, csa_tree_add_12_51_groupi_n_6763, csa_tree_add_12_51_groupi_n_6764;
  wire csa_tree_add_12_51_groupi_n_6765, csa_tree_add_12_51_groupi_n_6766, csa_tree_add_12_51_groupi_n_6767, csa_tree_add_12_51_groupi_n_6768, csa_tree_add_12_51_groupi_n_6769, csa_tree_add_12_51_groupi_n_6770, csa_tree_add_12_51_groupi_n_6771, csa_tree_add_12_51_groupi_n_6772;
  wire csa_tree_add_12_51_groupi_n_6773, csa_tree_add_12_51_groupi_n_6774, csa_tree_add_12_51_groupi_n_6775, csa_tree_add_12_51_groupi_n_6776, csa_tree_add_12_51_groupi_n_6777, csa_tree_add_12_51_groupi_n_6778, csa_tree_add_12_51_groupi_n_6779, csa_tree_add_12_51_groupi_n_6780;
  wire csa_tree_add_12_51_groupi_n_6781, csa_tree_add_12_51_groupi_n_6782, csa_tree_add_12_51_groupi_n_6783, csa_tree_add_12_51_groupi_n_6784, csa_tree_add_12_51_groupi_n_6785, csa_tree_add_12_51_groupi_n_6786, csa_tree_add_12_51_groupi_n_6787, csa_tree_add_12_51_groupi_n_6788;
  wire csa_tree_add_12_51_groupi_n_6789, csa_tree_add_12_51_groupi_n_6790, csa_tree_add_12_51_groupi_n_6791, csa_tree_add_12_51_groupi_n_6792, csa_tree_add_12_51_groupi_n_6793, csa_tree_add_12_51_groupi_n_6794, csa_tree_add_12_51_groupi_n_6795, csa_tree_add_12_51_groupi_n_6796;
  wire csa_tree_add_12_51_groupi_n_6797, csa_tree_add_12_51_groupi_n_6798, csa_tree_add_12_51_groupi_n_6799, csa_tree_add_12_51_groupi_n_6800, csa_tree_add_12_51_groupi_n_6801, csa_tree_add_12_51_groupi_n_6802, csa_tree_add_12_51_groupi_n_6803, csa_tree_add_12_51_groupi_n_6804;
  wire csa_tree_add_12_51_groupi_n_6805, csa_tree_add_12_51_groupi_n_6806, csa_tree_add_12_51_groupi_n_6807, csa_tree_add_12_51_groupi_n_6808, csa_tree_add_12_51_groupi_n_6809, csa_tree_add_12_51_groupi_n_6810, csa_tree_add_12_51_groupi_n_6811, csa_tree_add_12_51_groupi_n_6812;
  wire csa_tree_add_12_51_groupi_n_6813, csa_tree_add_12_51_groupi_n_6814, csa_tree_add_12_51_groupi_n_6815, csa_tree_add_12_51_groupi_n_6816, csa_tree_add_12_51_groupi_n_6817, csa_tree_add_12_51_groupi_n_6818, csa_tree_add_12_51_groupi_n_6819, csa_tree_add_12_51_groupi_n_6820;
  wire csa_tree_add_12_51_groupi_n_6821, csa_tree_add_12_51_groupi_n_6822, csa_tree_add_12_51_groupi_n_6823, csa_tree_add_12_51_groupi_n_6824, csa_tree_add_12_51_groupi_n_6825, csa_tree_add_12_51_groupi_n_6826, csa_tree_add_12_51_groupi_n_6827, csa_tree_add_12_51_groupi_n_6828;
  wire csa_tree_add_12_51_groupi_n_6829, csa_tree_add_12_51_groupi_n_6830, csa_tree_add_12_51_groupi_n_6831, csa_tree_add_12_51_groupi_n_6832, csa_tree_add_12_51_groupi_n_6833, csa_tree_add_12_51_groupi_n_6834, csa_tree_add_12_51_groupi_n_6835, csa_tree_add_12_51_groupi_n_6836;
  wire csa_tree_add_12_51_groupi_n_6837, csa_tree_add_12_51_groupi_n_6838, csa_tree_add_12_51_groupi_n_6839, csa_tree_add_12_51_groupi_n_6840, csa_tree_add_12_51_groupi_n_6841, csa_tree_add_12_51_groupi_n_6842, csa_tree_add_12_51_groupi_n_6843, csa_tree_add_12_51_groupi_n_6844;
  wire csa_tree_add_12_51_groupi_n_6845, csa_tree_add_12_51_groupi_n_6846, csa_tree_add_12_51_groupi_n_6847, csa_tree_add_12_51_groupi_n_6848, csa_tree_add_12_51_groupi_n_6849, csa_tree_add_12_51_groupi_n_6850, csa_tree_add_12_51_groupi_n_6851, csa_tree_add_12_51_groupi_n_6852;
  wire csa_tree_add_12_51_groupi_n_6854, csa_tree_add_12_51_groupi_n_6855, csa_tree_add_12_51_groupi_n_6856, csa_tree_add_12_51_groupi_n_6857, csa_tree_add_12_51_groupi_n_6858, csa_tree_add_12_51_groupi_n_6859, csa_tree_add_12_51_groupi_n_6860, csa_tree_add_12_51_groupi_n_6861;
  wire csa_tree_add_12_51_groupi_n_6862, csa_tree_add_12_51_groupi_n_6863, csa_tree_add_12_51_groupi_n_6864, csa_tree_add_12_51_groupi_n_6865, csa_tree_add_12_51_groupi_n_6866, csa_tree_add_12_51_groupi_n_6867, csa_tree_add_12_51_groupi_n_6868, csa_tree_add_12_51_groupi_n_6869;
  wire csa_tree_add_12_51_groupi_n_6870, csa_tree_add_12_51_groupi_n_6871, csa_tree_add_12_51_groupi_n_6872, csa_tree_add_12_51_groupi_n_6873, csa_tree_add_12_51_groupi_n_6874, csa_tree_add_12_51_groupi_n_6875, csa_tree_add_12_51_groupi_n_6876, csa_tree_add_12_51_groupi_n_6877;
  wire csa_tree_add_12_51_groupi_n_6878, csa_tree_add_12_51_groupi_n_6879, csa_tree_add_12_51_groupi_n_6880, csa_tree_add_12_51_groupi_n_6881, csa_tree_add_12_51_groupi_n_6882, csa_tree_add_12_51_groupi_n_6883, csa_tree_add_12_51_groupi_n_6884, csa_tree_add_12_51_groupi_n_6885;
  wire csa_tree_add_12_51_groupi_n_6886, csa_tree_add_12_51_groupi_n_6887, csa_tree_add_12_51_groupi_n_6888, csa_tree_add_12_51_groupi_n_6889, csa_tree_add_12_51_groupi_n_6890, csa_tree_add_12_51_groupi_n_6891, csa_tree_add_12_51_groupi_n_6892, csa_tree_add_12_51_groupi_n_6893;
  wire csa_tree_add_12_51_groupi_n_6894, csa_tree_add_12_51_groupi_n_6895, csa_tree_add_12_51_groupi_n_6896, csa_tree_add_12_51_groupi_n_6897, csa_tree_add_12_51_groupi_n_6898, csa_tree_add_12_51_groupi_n_6899, csa_tree_add_12_51_groupi_n_6900, csa_tree_add_12_51_groupi_n_6901;
  wire csa_tree_add_12_51_groupi_n_6902, csa_tree_add_12_51_groupi_n_6903, csa_tree_add_12_51_groupi_n_6904, csa_tree_add_12_51_groupi_n_6905, csa_tree_add_12_51_groupi_n_6906, csa_tree_add_12_51_groupi_n_6907, csa_tree_add_12_51_groupi_n_6908, csa_tree_add_12_51_groupi_n_6909;
  wire csa_tree_add_12_51_groupi_n_6910, csa_tree_add_12_51_groupi_n_6911, csa_tree_add_12_51_groupi_n_6912, csa_tree_add_12_51_groupi_n_6913, csa_tree_add_12_51_groupi_n_6914, csa_tree_add_12_51_groupi_n_6915, csa_tree_add_12_51_groupi_n_6916, csa_tree_add_12_51_groupi_n_6917;
  wire csa_tree_add_12_51_groupi_n_6918, csa_tree_add_12_51_groupi_n_6919, csa_tree_add_12_51_groupi_n_6920, csa_tree_add_12_51_groupi_n_6921, csa_tree_add_12_51_groupi_n_6922, csa_tree_add_12_51_groupi_n_6923, csa_tree_add_12_51_groupi_n_6924, csa_tree_add_12_51_groupi_n_6925;
  wire csa_tree_add_12_51_groupi_n_6926, csa_tree_add_12_51_groupi_n_6927, csa_tree_add_12_51_groupi_n_6928, csa_tree_add_12_51_groupi_n_6929, csa_tree_add_12_51_groupi_n_6930, csa_tree_add_12_51_groupi_n_6931, csa_tree_add_12_51_groupi_n_6932, csa_tree_add_12_51_groupi_n_6934;
  wire csa_tree_add_12_51_groupi_n_6935, csa_tree_add_12_51_groupi_n_6936, csa_tree_add_12_51_groupi_n_6937, csa_tree_add_12_51_groupi_n_6938, csa_tree_add_12_51_groupi_n_6939, csa_tree_add_12_51_groupi_n_6940, csa_tree_add_12_51_groupi_n_6941, csa_tree_add_12_51_groupi_n_6942;
  wire csa_tree_add_12_51_groupi_n_6943, csa_tree_add_12_51_groupi_n_6944, csa_tree_add_12_51_groupi_n_6945, csa_tree_add_12_51_groupi_n_6946, csa_tree_add_12_51_groupi_n_6947, csa_tree_add_12_51_groupi_n_6948, csa_tree_add_12_51_groupi_n_6949, csa_tree_add_12_51_groupi_n_6950;
  wire csa_tree_add_12_51_groupi_n_6951, csa_tree_add_12_51_groupi_n_6952, csa_tree_add_12_51_groupi_n_6953, csa_tree_add_12_51_groupi_n_6954, csa_tree_add_12_51_groupi_n_6955, csa_tree_add_12_51_groupi_n_6956, csa_tree_add_12_51_groupi_n_6957, csa_tree_add_12_51_groupi_n_6958;
  wire csa_tree_add_12_51_groupi_n_6959, csa_tree_add_12_51_groupi_n_6960, csa_tree_add_12_51_groupi_n_6961, csa_tree_add_12_51_groupi_n_6962, csa_tree_add_12_51_groupi_n_6963, csa_tree_add_12_51_groupi_n_6964, csa_tree_add_12_51_groupi_n_6965, csa_tree_add_12_51_groupi_n_6966;
  wire csa_tree_add_12_51_groupi_n_6967, csa_tree_add_12_51_groupi_n_6968, csa_tree_add_12_51_groupi_n_6969, csa_tree_add_12_51_groupi_n_6970, csa_tree_add_12_51_groupi_n_6971, csa_tree_add_12_51_groupi_n_6972, csa_tree_add_12_51_groupi_n_6973, csa_tree_add_12_51_groupi_n_6974;
  wire csa_tree_add_12_51_groupi_n_6975, csa_tree_add_12_51_groupi_n_6976, csa_tree_add_12_51_groupi_n_6977, csa_tree_add_12_51_groupi_n_6978, csa_tree_add_12_51_groupi_n_6979, csa_tree_add_12_51_groupi_n_6980, csa_tree_add_12_51_groupi_n_6981, csa_tree_add_12_51_groupi_n_6982;
  wire csa_tree_add_12_51_groupi_n_6983, csa_tree_add_12_51_groupi_n_6984, csa_tree_add_12_51_groupi_n_6985, csa_tree_add_12_51_groupi_n_6986, csa_tree_add_12_51_groupi_n_6987, csa_tree_add_12_51_groupi_n_6988, csa_tree_add_12_51_groupi_n_6989, csa_tree_add_12_51_groupi_n_6990;
  wire csa_tree_add_12_51_groupi_n_6991, csa_tree_add_12_51_groupi_n_6992, csa_tree_add_12_51_groupi_n_6993, csa_tree_add_12_51_groupi_n_6994, csa_tree_add_12_51_groupi_n_6995, csa_tree_add_12_51_groupi_n_6996, csa_tree_add_12_51_groupi_n_6997, csa_tree_add_12_51_groupi_n_6998;
  wire csa_tree_add_12_51_groupi_n_6999, csa_tree_add_12_51_groupi_n_7000, csa_tree_add_12_51_groupi_n_7001, csa_tree_add_12_51_groupi_n_7002, csa_tree_add_12_51_groupi_n_7003, csa_tree_add_12_51_groupi_n_7005, csa_tree_add_12_51_groupi_n_7006, csa_tree_add_12_51_groupi_n_7007;
  wire csa_tree_add_12_51_groupi_n_7008, csa_tree_add_12_51_groupi_n_7009, csa_tree_add_12_51_groupi_n_7010, csa_tree_add_12_51_groupi_n_7011, csa_tree_add_12_51_groupi_n_7012, csa_tree_add_12_51_groupi_n_7013, csa_tree_add_12_51_groupi_n_7014, csa_tree_add_12_51_groupi_n_7015;
  wire csa_tree_add_12_51_groupi_n_7016, csa_tree_add_12_51_groupi_n_7017, csa_tree_add_12_51_groupi_n_7018, csa_tree_add_12_51_groupi_n_7019, csa_tree_add_12_51_groupi_n_7020, csa_tree_add_12_51_groupi_n_7021, csa_tree_add_12_51_groupi_n_7022, csa_tree_add_12_51_groupi_n_7023;
  wire csa_tree_add_12_51_groupi_n_7024, csa_tree_add_12_51_groupi_n_7025, csa_tree_add_12_51_groupi_n_7026, csa_tree_add_12_51_groupi_n_7027, csa_tree_add_12_51_groupi_n_7028, csa_tree_add_12_51_groupi_n_7029, csa_tree_add_12_51_groupi_n_7030, csa_tree_add_12_51_groupi_n_7031;
  wire csa_tree_add_12_51_groupi_n_7032, csa_tree_add_12_51_groupi_n_7033, csa_tree_add_12_51_groupi_n_7034, csa_tree_add_12_51_groupi_n_7035, csa_tree_add_12_51_groupi_n_7036, csa_tree_add_12_51_groupi_n_7037, csa_tree_add_12_51_groupi_n_7038, csa_tree_add_12_51_groupi_n_7039;
  wire csa_tree_add_12_51_groupi_n_7040, csa_tree_add_12_51_groupi_n_7041, csa_tree_add_12_51_groupi_n_7042, csa_tree_add_12_51_groupi_n_7043, csa_tree_add_12_51_groupi_n_7044, csa_tree_add_12_51_groupi_n_7045, csa_tree_add_12_51_groupi_n_7046, csa_tree_add_12_51_groupi_n_7047;
  wire csa_tree_add_12_51_groupi_n_7048, csa_tree_add_12_51_groupi_n_7049, csa_tree_add_12_51_groupi_n_7050, csa_tree_add_12_51_groupi_n_7051, csa_tree_add_12_51_groupi_n_7052, csa_tree_add_12_51_groupi_n_7053, csa_tree_add_12_51_groupi_n_7054, csa_tree_add_12_51_groupi_n_7055;
  wire csa_tree_add_12_51_groupi_n_7056, csa_tree_add_12_51_groupi_n_7058, csa_tree_add_12_51_groupi_n_7059, csa_tree_add_12_51_groupi_n_7060, csa_tree_add_12_51_groupi_n_7061, csa_tree_add_12_51_groupi_n_7062, csa_tree_add_12_51_groupi_n_7063, csa_tree_add_12_51_groupi_n_7064;
  wire csa_tree_add_12_51_groupi_n_7065, csa_tree_add_12_51_groupi_n_7066, csa_tree_add_12_51_groupi_n_7067, csa_tree_add_12_51_groupi_n_7068, csa_tree_add_12_51_groupi_n_7069, csa_tree_add_12_51_groupi_n_7070, csa_tree_add_12_51_groupi_n_7071, csa_tree_add_12_51_groupi_n_7072;
  wire csa_tree_add_12_51_groupi_n_7073, csa_tree_add_12_51_groupi_n_7074, csa_tree_add_12_51_groupi_n_7075, csa_tree_add_12_51_groupi_n_7076, csa_tree_add_12_51_groupi_n_7077, csa_tree_add_12_51_groupi_n_7078, csa_tree_add_12_51_groupi_n_7079, csa_tree_add_12_51_groupi_n_7080;
  wire csa_tree_add_12_51_groupi_n_7081, csa_tree_add_12_51_groupi_n_7082, csa_tree_add_12_51_groupi_n_7083, csa_tree_add_12_51_groupi_n_7084, csa_tree_add_12_51_groupi_n_7085, csa_tree_add_12_51_groupi_n_7086, csa_tree_add_12_51_groupi_n_7087, csa_tree_add_12_51_groupi_n_7088;
  wire csa_tree_add_12_51_groupi_n_7089, csa_tree_add_12_51_groupi_n_7090, csa_tree_add_12_51_groupi_n_7091, csa_tree_add_12_51_groupi_n_7092, csa_tree_add_12_51_groupi_n_7093, csa_tree_add_12_51_groupi_n_7094, csa_tree_add_12_51_groupi_n_7095, csa_tree_add_12_51_groupi_n_7096;
  wire csa_tree_add_12_51_groupi_n_7097, csa_tree_add_12_51_groupi_n_7098, csa_tree_add_12_51_groupi_n_7099, csa_tree_add_12_51_groupi_n_7101, csa_tree_add_12_51_groupi_n_7102, csa_tree_add_12_51_groupi_n_7103, csa_tree_add_12_51_groupi_n_7104, csa_tree_add_12_51_groupi_n_7105;
  wire csa_tree_add_12_51_groupi_n_7106, csa_tree_add_12_51_groupi_n_7107, csa_tree_add_12_51_groupi_n_7108, csa_tree_add_12_51_groupi_n_7109, csa_tree_add_12_51_groupi_n_7110, csa_tree_add_12_51_groupi_n_7111, csa_tree_add_12_51_groupi_n_7112, csa_tree_add_12_51_groupi_n_7113;
  wire csa_tree_add_12_51_groupi_n_7114, csa_tree_add_12_51_groupi_n_7115, csa_tree_add_12_51_groupi_n_7116, csa_tree_add_12_51_groupi_n_7117, csa_tree_add_12_51_groupi_n_7118, csa_tree_add_12_51_groupi_n_7119, csa_tree_add_12_51_groupi_n_7120, csa_tree_add_12_51_groupi_n_7121;
  wire csa_tree_add_12_51_groupi_n_7122, csa_tree_add_12_51_groupi_n_7123, csa_tree_add_12_51_groupi_n_7124, csa_tree_add_12_51_groupi_n_7125, csa_tree_add_12_51_groupi_n_7126, csa_tree_add_12_51_groupi_n_7128, csa_tree_add_12_51_groupi_n_7129, csa_tree_add_12_51_groupi_n_7131;
  wire csa_tree_add_12_51_groupi_n_7132, csa_tree_add_12_51_groupi_n_7134, csa_tree_add_12_51_groupi_n_7135, csa_tree_add_12_51_groupi_n_7137, csa_tree_add_12_51_groupi_n_7138, csa_tree_add_12_51_groupi_n_7140, csa_tree_add_12_51_groupi_n_7141, csa_tree_add_12_51_groupi_n_7143;
  wire csa_tree_add_12_51_groupi_n_7144, csa_tree_add_12_51_groupi_n_7146, csa_tree_add_12_51_groupi_n_7147, csa_tree_add_12_51_groupi_n_7149, csa_tree_add_12_51_groupi_n_7150, csa_tree_add_12_51_groupi_n_7152, csa_tree_add_12_51_groupi_n_7153, csa_tree_add_12_51_groupi_n_7155;
  wire csa_tree_add_12_51_groupi_n_7156, csa_tree_add_12_51_groupi_n_7158, csa_tree_add_12_51_groupi_n_7159, csa_tree_add_12_51_groupi_n_7161, csa_tree_add_12_51_groupi_n_7162, csa_tree_add_12_51_groupi_n_7163, csa_tree_add_12_51_groupi_n_7165, csa_tree_add_12_51_groupi_n_7166;
  wire csa_tree_add_12_51_groupi_n_7168, csa_tree_add_12_51_groupi_n_7169, csa_tree_add_12_51_groupi_n_7170, csa_tree_add_12_51_groupi_n_7172, csa_tree_add_12_51_groupi_n_7173, csa_tree_add_12_51_groupi_n_7175, sub_11_21_n_0, sub_11_21_n_1;
  wire sub_11_21_n_2, sub_11_21_n_3, sub_11_21_n_4, sub_11_21_n_5, sub_11_21_n_6, sub_11_21_n_7, sub_11_21_n_8, sub_11_21_n_9;
  wire sub_11_21_n_10, sub_11_21_n_11, sub_11_21_n_12, sub_11_21_n_13, sub_11_21_n_14, sub_11_21_n_15, sub_11_21_n_16, sub_11_21_n_17;
  wire sub_11_21_n_18, sub_11_21_n_19, sub_11_21_n_20, sub_11_21_n_21, sub_11_21_n_22, sub_11_21_n_23, sub_11_21_n_24, sub_11_21_n_25;
  wire sub_11_21_n_26, sub_11_21_n_27, sub_11_21_n_28, sub_11_21_n_29, sub_11_21_n_30, sub_11_21_n_31, sub_11_21_n_32, sub_11_21_n_33;
  wire sub_11_21_n_34, sub_11_21_n_35, sub_11_21_n_36, sub_11_21_n_37, sub_11_21_n_38, sub_11_21_n_39, sub_11_21_n_40, sub_11_21_n_41;
  wire sub_11_21_n_42, sub_11_21_n_43, sub_11_21_n_44, sub_11_21_n_45, sub_11_21_n_46, sub_11_21_n_47, sub_11_21_n_48, sub_11_21_n_49;
  wire sub_11_21_n_50, sub_11_21_n_51, sub_11_21_n_52, sub_11_21_n_53, sub_11_21_n_54, sub_11_21_n_55, sub_11_21_n_56, sub_11_21_n_57;
  wire sub_11_21_n_58, sub_11_21_n_59, sub_11_21_n_60, sub_11_21_n_61, sub_11_21_n_62, sub_11_21_n_63, sub_11_21_n_64, sub_11_21_n_65;
  wire sub_11_21_n_66, sub_11_21_n_67, sub_11_21_n_68, sub_11_21_n_69, sub_11_21_n_70, sub_11_21_n_71, sub_11_21_n_72, sub_11_21_n_73;
  wire sub_11_21_n_74, sub_11_21_n_75, sub_11_21_n_76, sub_11_21_n_77, sub_11_21_n_78, sub_11_21_n_79, sub_11_21_n_80, sub_11_21_n_81;
  wire sub_11_21_n_82, sub_11_21_n_83, sub_11_21_n_84, sub_11_21_n_85, sub_11_21_n_86, sub_11_21_n_87, sub_11_21_n_88, sub_11_21_n_89;
  wire sub_11_21_n_90, sub_11_21_n_91, sub_11_21_n_92, sub_11_21_n_93, sub_11_21_n_94, sub_11_21_n_95, sub_11_21_n_96, sub_11_21_n_98;
  wire sub_11_21_n_100, sub_11_21_n_102, sub_11_21_n_103, sub_11_21_n_105, sub_11_21_n_106, sub_11_21_n_108, sub_11_21_n_109, sub_11_21_n_111;
  wire sub_11_21_n_112, sub_11_21_n_114, sub_11_21_n_115, sub_11_21_n_117, sub_11_21_n_118, sub_11_21_n_120, sub_11_21_n_121, sub_11_21_n_123;
  wire sub_11_21_n_124, sub_11_21_n_126, sub_11_21_n_127, sub_11_21_n_129, sub_11_21_n_130, sub_11_21_n_132, sub_11_21_n_133, sub_11_21_n_135;
  wire sub_11_21_n_136, sub_11_21_n_138, sub_11_21_n_139, sub_11_21_n_141;
  or add_10_21_g333__2398(out1[16] ,add_10_21_n_30 ,add_10_21_n_93);
  xnor add_10_21_g334__5107(out1[15] ,add_10_21_n_92 ,add_10_21_n_40);
  and add_10_21_g335__6260(add_10_21_n_93 ,add_10_21_n_16 ,add_10_21_n_92);
  or add_10_21_g336__4319(add_10_21_n_92 ,add_10_21_n_25 ,add_10_21_n_90);
  xnor add_10_21_g337__8428(out1[14] ,add_10_21_n_89 ,add_10_21_n_39);
  and add_10_21_g338__5526(add_10_21_n_90 ,add_10_21_n_10 ,add_10_21_n_89);
  or add_10_21_g339__6783(add_10_21_n_89 ,add_10_21_n_21 ,add_10_21_n_87);
  xnor add_10_21_g340__3680(out1[13] ,add_10_21_n_86 ,add_10_21_n_38);
  and add_10_21_g341__1617(add_10_21_n_87 ,add_10_21_n_17 ,add_10_21_n_86);
  or add_10_21_g342__2802(add_10_21_n_86 ,add_10_21_n_11 ,add_10_21_n_84);
  xnor add_10_21_g343__1705(out1[12] ,add_10_21_n_83 ,add_10_21_n_37);
  and add_10_21_g344__5122(add_10_21_n_84 ,add_10_21_n_13 ,add_10_21_n_83);
  or add_10_21_g345__8246(add_10_21_n_83 ,add_10_21_n_9 ,add_10_21_n_81);
  xnor add_10_21_g346__7098(out1[11] ,add_10_21_n_80 ,add_10_21_n_36);
  and add_10_21_g347__6131(add_10_21_n_81 ,add_10_21_n_23 ,add_10_21_n_80);
  or add_10_21_g348__1881(add_10_21_n_80 ,add_10_21_n_33 ,add_10_21_n_78);
  xnor add_10_21_g349__5115(out1[10] ,add_10_21_n_77 ,add_10_21_n_43);
  and add_10_21_g350__7482(add_10_21_n_78 ,add_10_21_n_3 ,add_10_21_n_77);
  or add_10_21_g351__4733(add_10_21_n_77 ,add_10_21_n_22 ,add_10_21_n_75);
  xnor add_10_21_g352__6161(out1[9] ,add_10_21_n_74 ,add_10_21_n_49);
  and add_10_21_g353__9315(add_10_21_n_75 ,add_10_21_n_20 ,add_10_21_n_74);
  or add_10_21_g354__9945(add_10_21_n_74 ,add_10_21_n_29 ,add_10_21_n_72);
  xnor add_10_21_g355__2883(out1[8] ,add_10_21_n_71 ,add_10_21_n_48);
  and add_10_21_g356__2346(add_10_21_n_72 ,add_10_21_n_12 ,add_10_21_n_71);
  or add_10_21_g357__1666(add_10_21_n_71 ,add_10_21_n_18 ,add_10_21_n_69);
  xnor add_10_21_g358__7410(out1[7] ,add_10_21_n_68 ,add_10_21_n_47);
  and add_10_21_g359__6417(add_10_21_n_69 ,add_10_21_n_26 ,add_10_21_n_68);
  or add_10_21_g360__5477(add_10_21_n_68 ,add_10_21_n_7 ,add_10_21_n_66);
  xnor add_10_21_g361__2398(out1[6] ,add_10_21_n_65 ,add_10_21_n_46);
  and add_10_21_g362__5107(add_10_21_n_66 ,add_10_21_n_19 ,add_10_21_n_65);
  or add_10_21_g363__6260(add_10_21_n_65 ,add_10_21_n_4 ,add_10_21_n_63);
  xnor add_10_21_g364__4319(out1[5] ,add_10_21_n_62 ,add_10_21_n_45);
  and add_10_21_g365__8428(add_10_21_n_63 ,add_10_21_n_31 ,add_10_21_n_62);
  or add_10_21_g366__5526(add_10_21_n_62 ,add_10_21_n_32 ,add_10_21_n_60);
  xnor add_10_21_g367__6783(out1[4] ,add_10_21_n_59 ,add_10_21_n_44);
  and add_10_21_g368__3680(add_10_21_n_60 ,add_10_21_n_27 ,add_10_21_n_59);
  or add_10_21_g369__1617(add_10_21_n_59 ,add_10_21_n_28 ,add_10_21_n_57);
  xnor add_10_21_g370__2802(out1[3] ,add_10_21_n_56 ,add_10_21_n_35);
  and add_10_21_g371__1705(add_10_21_n_57 ,add_10_21_n_8 ,add_10_21_n_56);
  or add_10_21_g372__5122(add_10_21_n_56 ,add_10_21_n_6 ,add_10_21_n_54);
  xnor add_10_21_g373__8246(out1[2] ,add_10_21_n_52 ,add_10_21_n_42);
  and add_10_21_g374__7098(add_10_21_n_54 ,add_10_21_n_24 ,add_10_21_n_52);
  xor add_10_21_g375__6131(out1[1] ,add_10_21_n_34 ,add_10_21_n_41);
  or add_10_21_g376__1881(add_10_21_n_52 ,add_10_21_n_5 ,add_10_21_n_50);
  and add_10_21_g377__5115(add_10_21_n_51 ,add_10_21_n_34 ,add_10_21_n_14);
  nor add_10_21_g378__7482(add_10_21_n_50 ,add_10_21_n_34 ,add_10_21_n_15);
  xnor add_10_21_g379__4733(add_10_21_n_49 ,in1[9] ,in2[9]);
  xnor add_10_21_g380__6161(add_10_21_n_48 ,in1[8] ,in2[8]);
  xnor add_10_21_g381__9315(add_10_21_n_47 ,in1[7] ,in2[7]);
  xnor add_10_21_g382__9945(add_10_21_n_46 ,in1[6] ,in2[6]);
  xnor add_10_21_g383__2883(add_10_21_n_45 ,in1[5] ,in2[5]);
  xnor add_10_21_g384__2346(add_10_21_n_44 ,in1[4] ,in2[4]);
  xnor add_10_21_g385__1666(add_10_21_n_43 ,in1[10] ,in2[10]);
  xnor add_10_21_g386__7410(add_10_21_n_42 ,in1[2] ,in2[2]);
  xnor add_10_21_g387__6417(add_10_21_n_41 ,in1[1] ,in2[1]);
  xnor add_10_21_g388__5477(add_10_21_n_40 ,in1[15] ,in2[15]);
  xnor add_10_21_g389__2398(add_10_21_n_39 ,in1[14] ,in2[14]);
  xnor add_10_21_g390__5107(add_10_21_n_38 ,in1[13] ,in2[13]);
  xnor add_10_21_g391__6260(add_10_21_n_37 ,in1[12] ,in2[12]);
  xnor add_10_21_g392__4319(add_10_21_n_36 ,in1[11] ,in2[11]);
  xnor add_10_21_g393__8428(add_10_21_n_35 ,in1[3] ,in2[3]);
  and add_10_21_g394__5526(add_10_21_n_33 ,in1[10] ,in2[10]);
  and add_10_21_g395__6783(add_10_21_n_32 ,in1[4] ,in2[4]);
  or add_10_21_g396__3680(add_10_21_n_31 ,in1[5] ,in2[5]);
  and add_10_21_g397__1617(add_10_21_n_30 ,in1[15] ,in2[15]);
  and add_10_21_g398__2802(add_10_21_n_29 ,in1[8] ,in2[8]);
  and add_10_21_g399__1705(add_10_21_n_28 ,in1[3] ,in2[3]);
  or add_10_21_g400__5122(add_10_21_n_27 ,in1[4] ,in2[4]);
  or add_10_21_g401__8246(add_10_21_n_26 ,in1[7] ,in2[7]);
  and add_10_21_g402__7098(add_10_21_n_25 ,in1[14] ,in2[14]);
  or add_10_21_g403__6131(add_10_21_n_24 ,in1[2] ,in2[2]);
  or add_10_21_g404__1881(add_10_21_n_23 ,in1[11] ,in2[11]);
  and add_10_21_g405__5115(add_10_21_n_22 ,in1[9] ,in2[9]);
  and add_10_21_g406__7482(add_10_21_n_21 ,in1[13] ,in2[13]);
  or add_10_21_g407__4733(add_10_21_n_20 ,in1[9] ,in2[9]);
  or add_10_21_g408__6161(add_10_21_n_19 ,in1[6] ,in2[6]);
  or add_10_21_g409__9315(add_10_21_n_34 ,add_10_21_n_2 ,add_10_21_n_1);
  and add_10_21_g410__9945(add_10_21_n_18 ,in1[7] ,in2[7]);
  or add_10_21_g411__2883(add_10_21_n_17 ,in1[13] ,in2[13]);
  or add_10_21_g412__2346(add_10_21_n_16 ,in1[15] ,in2[15]);
  nor add_10_21_g413__1666(add_10_21_n_15 ,in1[1] ,in2[1]);
  or add_10_21_g414__7410(add_10_21_n_14 ,in1[0] ,in2[0]);
  or add_10_21_g415__6417(add_10_21_n_13 ,in1[12] ,in2[12]);
  or add_10_21_g416__5477(add_10_21_n_12 ,in1[8] ,in2[8]);
  and add_10_21_g417__2398(add_10_21_n_11 ,in1[12] ,in2[12]);
  or add_10_21_g418__5107(add_10_21_n_10 ,in1[14] ,in2[14]);
  and add_10_21_g419__6260(add_10_21_n_9 ,in1[11] ,in2[11]);
  or add_10_21_g420__4319(add_10_21_n_8 ,in1[3] ,in2[3]);
  and add_10_21_g421__8428(add_10_21_n_7 ,in1[6] ,in2[6]);
  and add_10_21_g422__5526(add_10_21_n_6 ,in1[2] ,in2[2]);
  and add_10_21_g423__6783(add_10_21_n_5 ,in1[1] ,in2[1]);
  and add_10_21_g424__3680(add_10_21_n_4 ,in1[5] ,in2[5]);
  or add_10_21_g425__1617(add_10_21_n_3 ,in1[10] ,in2[10]);
  not add_10_21_g426(add_10_21_n_2 ,in1[0]);
  not add_10_21_g427(add_10_21_n_1 ,in2[0]);
  buf add_10_21_drc_bufs(out1[0] ,add_10_21_n_51);
  xnor csa_tree_add_12_51_groupi_g14586__2802(out3[33] ,csa_tree_add_12_51_groupi_n_4774 ,csa_tree_add_12_51_groupi_n_7175);
  or csa_tree_add_12_51_groupi_g14587__1705(csa_tree_add_12_51_groupi_n_7175 ,csa_tree_add_12_51_groupi_n_5292 ,csa_tree_add_12_51_groupi_n_7173);
  xnor csa_tree_add_12_51_groupi_g14588__5122(out3[32] ,csa_tree_add_12_51_groupi_n_7172 ,csa_tree_add_12_51_groupi_n_5326);
  nor csa_tree_add_12_51_groupi_g14589__8246(csa_tree_add_12_51_groupi_n_7173 ,csa_tree_add_12_51_groupi_n_5291 ,csa_tree_add_12_51_groupi_n_7172);
  and csa_tree_add_12_51_groupi_g14590__7098(csa_tree_add_12_51_groupi_n_7172 ,csa_tree_add_12_51_groupi_n_6984 ,csa_tree_add_12_51_groupi_n_7170);
  xnor csa_tree_add_12_51_groupi_g14591__6131(out3[31] ,csa_tree_add_12_51_groupi_n_7168 ,csa_tree_add_12_51_groupi_n_6995);
  or csa_tree_add_12_51_groupi_g14592__1881(csa_tree_add_12_51_groupi_n_7170 ,csa_tree_add_12_51_groupi_n_6986 ,csa_tree_add_12_51_groupi_n_7169);
  not csa_tree_add_12_51_groupi_g14593(csa_tree_add_12_51_groupi_n_7169 ,csa_tree_add_12_51_groupi_n_7168);
  or csa_tree_add_12_51_groupi_g14594__5115(csa_tree_add_12_51_groupi_n_7168 ,csa_tree_add_12_51_groupi_n_7045 ,csa_tree_add_12_51_groupi_n_7166);
  xnor csa_tree_add_12_51_groupi_g14595__7482(out3[30] ,csa_tree_add_12_51_groupi_n_7165 ,csa_tree_add_12_51_groupi_n_7055);
  nor csa_tree_add_12_51_groupi_g14596__4733(csa_tree_add_12_51_groupi_n_7166 ,csa_tree_add_12_51_groupi_n_7052 ,csa_tree_add_12_51_groupi_n_7165);
  and csa_tree_add_12_51_groupi_g14597__6161(csa_tree_add_12_51_groupi_n_7165 ,csa_tree_add_12_51_groupi_n_7087 ,csa_tree_add_12_51_groupi_n_7163);
  xnor csa_tree_add_12_51_groupi_g14598__9315(out3[29] ,csa_tree_add_12_51_groupi_n_7161 ,csa_tree_add_12_51_groupi_n_7096);
  or csa_tree_add_12_51_groupi_g14599__9945(csa_tree_add_12_51_groupi_n_7163 ,csa_tree_add_12_51_groupi_n_7162 ,csa_tree_add_12_51_groupi_n_7094);
  not csa_tree_add_12_51_groupi_g14600(csa_tree_add_12_51_groupi_n_7162 ,csa_tree_add_12_51_groupi_n_7161);
  or csa_tree_add_12_51_groupi_g14601__2883(csa_tree_add_12_51_groupi_n_7161 ,csa_tree_add_12_51_groupi_n_7159 ,csa_tree_add_12_51_groupi_n_7092);
  xnor csa_tree_add_12_51_groupi_g14602__2346(out3[28] ,csa_tree_add_12_51_groupi_n_7158 ,csa_tree_add_12_51_groupi_n_7099);
  and csa_tree_add_12_51_groupi_g14603__1666(csa_tree_add_12_51_groupi_n_7159 ,csa_tree_add_12_51_groupi_n_7093 ,csa_tree_add_12_51_groupi_n_7158);
  or csa_tree_add_12_51_groupi_g14604__7410(csa_tree_add_12_51_groupi_n_7158 ,csa_tree_add_12_51_groupi_n_7156 ,csa_tree_add_12_51_groupi_n_7114);
  xnor csa_tree_add_12_51_groupi_g14605__6417(out3[27] ,csa_tree_add_12_51_groupi_n_7155 ,csa_tree_add_12_51_groupi_n_7125);
  and csa_tree_add_12_51_groupi_g14606__5477(csa_tree_add_12_51_groupi_n_7156 ,csa_tree_add_12_51_groupi_n_7111 ,csa_tree_add_12_51_groupi_n_7155);
  or csa_tree_add_12_51_groupi_g14607__2398(csa_tree_add_12_51_groupi_n_7155 ,csa_tree_add_12_51_groupi_n_7153 ,csa_tree_add_12_51_groupi_n_7113);
  xnor csa_tree_add_12_51_groupi_g14608__5107(out3[26] ,csa_tree_add_12_51_groupi_n_7152 ,csa_tree_add_12_51_groupi_n_7124);
  and csa_tree_add_12_51_groupi_g14609__6260(csa_tree_add_12_51_groupi_n_7153 ,csa_tree_add_12_51_groupi_n_7115 ,csa_tree_add_12_51_groupi_n_7152);
  or csa_tree_add_12_51_groupi_g14610__4319(csa_tree_add_12_51_groupi_n_7152 ,csa_tree_add_12_51_groupi_n_7106 ,csa_tree_add_12_51_groupi_n_7150);
  xnor csa_tree_add_12_51_groupi_g14611__8428(out3[25] ,csa_tree_add_12_51_groupi_n_7149 ,csa_tree_add_12_51_groupi_n_7123);
  and csa_tree_add_12_51_groupi_g14612__5526(csa_tree_add_12_51_groupi_n_7150 ,csa_tree_add_12_51_groupi_n_7109 ,csa_tree_add_12_51_groupi_n_7149);
  or csa_tree_add_12_51_groupi_g14613__6783(csa_tree_add_12_51_groupi_n_7149 ,csa_tree_add_12_51_groupi_n_7147 ,csa_tree_add_12_51_groupi_n_7105);
  xnor csa_tree_add_12_51_groupi_g14614__3680(out3[24] ,csa_tree_add_12_51_groupi_n_7146 ,csa_tree_add_12_51_groupi_n_7122);
  and csa_tree_add_12_51_groupi_g14615__1617(csa_tree_add_12_51_groupi_n_7147 ,csa_tree_add_12_51_groupi_n_7108 ,csa_tree_add_12_51_groupi_n_7146);
  or csa_tree_add_12_51_groupi_g14616__2802(csa_tree_add_12_51_groupi_n_7146 ,csa_tree_add_12_51_groupi_n_7144 ,csa_tree_add_12_51_groupi_n_7101);
  xnor csa_tree_add_12_51_groupi_g14617__1705(out3[23] ,csa_tree_add_12_51_groupi_n_7143 ,csa_tree_add_12_51_groupi_n_7121);
  and csa_tree_add_12_51_groupi_g14618__5122(csa_tree_add_12_51_groupi_n_7144 ,csa_tree_add_12_51_groupi_n_7143 ,csa_tree_add_12_51_groupi_n_7102);
  or csa_tree_add_12_51_groupi_g14619__8246(csa_tree_add_12_51_groupi_n_7143 ,csa_tree_add_12_51_groupi_n_7107 ,csa_tree_add_12_51_groupi_n_7141);
  xnor csa_tree_add_12_51_groupi_g14620__7098(out3[22] ,csa_tree_add_12_51_groupi_n_7140 ,csa_tree_add_12_51_groupi_n_7120);
  and csa_tree_add_12_51_groupi_g14621__6131(csa_tree_add_12_51_groupi_n_7141 ,csa_tree_add_12_51_groupi_n_7140 ,csa_tree_add_12_51_groupi_n_7103);
  or csa_tree_add_12_51_groupi_g14622__1881(csa_tree_add_12_51_groupi_n_7140 ,csa_tree_add_12_51_groupi_n_7138 ,csa_tree_add_12_51_groupi_n_7104);
  xnor csa_tree_add_12_51_groupi_g14623__5115(out3[21] ,csa_tree_add_12_51_groupi_n_7137 ,csa_tree_add_12_51_groupi_n_7119);
  and csa_tree_add_12_51_groupi_g14624__7482(csa_tree_add_12_51_groupi_n_7138 ,csa_tree_add_12_51_groupi_n_7137 ,csa_tree_add_12_51_groupi_n_7110);
  or csa_tree_add_12_51_groupi_g14625__4733(csa_tree_add_12_51_groupi_n_7137 ,csa_tree_add_12_51_groupi_n_7095 ,csa_tree_add_12_51_groupi_n_7135);
  xnor csa_tree_add_12_51_groupi_g14626__6161(out3[20] ,csa_tree_add_12_51_groupi_n_7134 ,csa_tree_add_12_51_groupi_n_7097);
  and csa_tree_add_12_51_groupi_g14627__9315(csa_tree_add_12_51_groupi_n_7135 ,csa_tree_add_12_51_groupi_n_7134 ,csa_tree_add_12_51_groupi_n_7088);
  or csa_tree_add_12_51_groupi_g14628__9945(csa_tree_add_12_51_groupi_n_7134 ,csa_tree_add_12_51_groupi_n_7132 ,csa_tree_add_12_51_groupi_n_7112);
  xnor csa_tree_add_12_51_groupi_g14629__2883(out3[19] ,csa_tree_add_12_51_groupi_n_7131 ,csa_tree_add_12_51_groupi_n_7118);
  and csa_tree_add_12_51_groupi_g14630__2346(csa_tree_add_12_51_groupi_n_7132 ,csa_tree_add_12_51_groupi_n_7116 ,csa_tree_add_12_51_groupi_n_7131);
  or csa_tree_add_12_51_groupi_g14631__1666(csa_tree_add_12_51_groupi_n_7131 ,csa_tree_add_12_51_groupi_n_7091 ,csa_tree_add_12_51_groupi_n_7129);
  xnor csa_tree_add_12_51_groupi_g14632__7410(out3[18] ,csa_tree_add_12_51_groupi_n_7128 ,csa_tree_add_12_51_groupi_n_7098);
  and csa_tree_add_12_51_groupi_g14633__6417(csa_tree_add_12_51_groupi_n_7129 ,csa_tree_add_12_51_groupi_n_7128 ,csa_tree_add_12_51_groupi_n_7090);
  or csa_tree_add_12_51_groupi_g14634__5477(csa_tree_add_12_51_groupi_n_7128 ,csa_tree_add_12_51_groupi_n_7126 ,csa_tree_add_12_51_groupi_n_7065);
  xnor csa_tree_add_12_51_groupi_g14635__2398(out3[17] ,csa_tree_add_12_51_groupi_n_7117 ,csa_tree_add_12_51_groupi_n_7076);
  nor csa_tree_add_12_51_groupi_g14636__5107(csa_tree_add_12_51_groupi_n_7126 ,csa_tree_add_12_51_groupi_n_7117 ,csa_tree_add_12_51_groupi_n_7066);
  xnor csa_tree_add_12_51_groupi_g14637__6260(csa_tree_add_12_51_groupi_n_7125 ,csa_tree_add_12_51_groupi_n_7084 ,csa_tree_add_12_51_groupi_n_7067);
  xnor csa_tree_add_12_51_groupi_g14638__4319(csa_tree_add_12_51_groupi_n_7124 ,csa_tree_add_12_51_groupi_n_7054 ,csa_tree_add_12_51_groupi_n_7080);
  xnor csa_tree_add_12_51_groupi_g14639__8428(csa_tree_add_12_51_groupi_n_7123 ,csa_tree_add_12_51_groupi_n_7072 ,csa_tree_add_12_51_groupi_n_7083);
  xnor csa_tree_add_12_51_groupi_g14640__5526(csa_tree_add_12_51_groupi_n_7122 ,csa_tree_add_12_51_groupi_n_7082 ,csa_tree_add_12_51_groupi_n_7071);
  xnor csa_tree_add_12_51_groupi_g14641__6783(csa_tree_add_12_51_groupi_n_7121 ,csa_tree_add_12_51_groupi_n_7070 ,csa_tree_add_12_51_groupi_n_7077);
  xnor csa_tree_add_12_51_groupi_g14642__3680(csa_tree_add_12_51_groupi_n_7120 ,csa_tree_add_12_51_groupi_n_7081 ,csa_tree_add_12_51_groupi_n_7058);
  xnor csa_tree_add_12_51_groupi_g14643__1617(csa_tree_add_12_51_groupi_n_7119 ,csa_tree_add_12_51_groupi_n_7061 ,csa_tree_add_12_51_groupi_n_7078);
  xnor csa_tree_add_12_51_groupi_g14644__2802(csa_tree_add_12_51_groupi_n_7118 ,csa_tree_add_12_51_groupi_n_7086 ,csa_tree_add_12_51_groupi_n_7069);
  or csa_tree_add_12_51_groupi_g14645__1705(csa_tree_add_12_51_groupi_n_7116 ,csa_tree_add_12_51_groupi_n_7068 ,csa_tree_add_12_51_groupi_n_7085);
  or csa_tree_add_12_51_groupi_g14646__5122(csa_tree_add_12_51_groupi_n_7115 ,csa_tree_add_12_51_groupi_n_7079 ,csa_tree_add_12_51_groupi_n_7053);
  and csa_tree_add_12_51_groupi_g14647__8246(csa_tree_add_12_51_groupi_n_7114 ,csa_tree_add_12_51_groupi_n_7084 ,csa_tree_add_12_51_groupi_n_7067);
  nor csa_tree_add_12_51_groupi_g14648__7098(csa_tree_add_12_51_groupi_n_7113 ,csa_tree_add_12_51_groupi_n_7080 ,csa_tree_add_12_51_groupi_n_7054);
  nor csa_tree_add_12_51_groupi_g14649__6131(csa_tree_add_12_51_groupi_n_7112 ,csa_tree_add_12_51_groupi_n_7069 ,csa_tree_add_12_51_groupi_n_7086);
  or csa_tree_add_12_51_groupi_g14650__1881(csa_tree_add_12_51_groupi_n_7111 ,csa_tree_add_12_51_groupi_n_7084 ,csa_tree_add_12_51_groupi_n_7067);
  or csa_tree_add_12_51_groupi_g14651__5115(csa_tree_add_12_51_groupi_n_7110 ,csa_tree_add_12_51_groupi_n_7061 ,csa_tree_add_12_51_groupi_n_7078);
  or csa_tree_add_12_51_groupi_g14652__7482(csa_tree_add_12_51_groupi_n_7109 ,csa_tree_add_12_51_groupi_n_7072 ,csa_tree_add_12_51_groupi_n_7083);
  or csa_tree_add_12_51_groupi_g14653__4733(csa_tree_add_12_51_groupi_n_7108 ,csa_tree_add_12_51_groupi_n_7082 ,csa_tree_add_12_51_groupi_n_7071);
  and csa_tree_add_12_51_groupi_g14654__6161(csa_tree_add_12_51_groupi_n_7107 ,csa_tree_add_12_51_groupi_n_7081 ,csa_tree_add_12_51_groupi_n_7058);
  and csa_tree_add_12_51_groupi_g14655__9315(csa_tree_add_12_51_groupi_n_7117 ,csa_tree_add_12_51_groupi_n_7089 ,csa_tree_add_12_51_groupi_n_7042);
  and csa_tree_add_12_51_groupi_g14656__9945(csa_tree_add_12_51_groupi_n_7106 ,csa_tree_add_12_51_groupi_n_7072 ,csa_tree_add_12_51_groupi_n_7083);
  and csa_tree_add_12_51_groupi_g14657__2883(csa_tree_add_12_51_groupi_n_7105 ,csa_tree_add_12_51_groupi_n_7082 ,csa_tree_add_12_51_groupi_n_7071);
  and csa_tree_add_12_51_groupi_g14658__2346(csa_tree_add_12_51_groupi_n_7104 ,csa_tree_add_12_51_groupi_n_7061 ,csa_tree_add_12_51_groupi_n_7078);
  or csa_tree_add_12_51_groupi_g14659__1666(csa_tree_add_12_51_groupi_n_7103 ,csa_tree_add_12_51_groupi_n_7081 ,csa_tree_add_12_51_groupi_n_7058);
  or csa_tree_add_12_51_groupi_g14660__7410(csa_tree_add_12_51_groupi_n_7102 ,csa_tree_add_12_51_groupi_n_7070 ,csa_tree_add_12_51_groupi_n_7077);
  and csa_tree_add_12_51_groupi_g14661__6417(csa_tree_add_12_51_groupi_n_7101 ,csa_tree_add_12_51_groupi_n_7070 ,csa_tree_add_12_51_groupi_n_7077);
  xnor csa_tree_add_12_51_groupi_g14662__5477(out3[16] ,csa_tree_add_12_51_groupi_n_7075 ,csa_tree_add_12_51_groupi_n_7056);
  xnor csa_tree_add_12_51_groupi_g14663__2398(csa_tree_add_12_51_groupi_n_7099 ,csa_tree_add_12_51_groupi_n_7074 ,csa_tree_add_12_51_groupi_n_7041);
  xnor csa_tree_add_12_51_groupi_g14664__5107(csa_tree_add_12_51_groupi_n_7098 ,csa_tree_add_12_51_groupi_n_7023 ,csa_tree_add_12_51_groupi_n_7059);
  xnor csa_tree_add_12_51_groupi_g14665__6260(csa_tree_add_12_51_groupi_n_7097 ,csa_tree_add_12_51_groupi_n_7062 ,csa_tree_add_12_51_groupi_n_7060);
  xnor csa_tree_add_12_51_groupi_g14666__4319(csa_tree_add_12_51_groupi_n_7096 ,csa_tree_add_12_51_groupi_n_7006 ,csa_tree_add_12_51_groupi_n_7064);
  and csa_tree_add_12_51_groupi_g14667__8428(csa_tree_add_12_51_groupi_n_7095 ,csa_tree_add_12_51_groupi_n_7062 ,csa_tree_add_12_51_groupi_n_7060);
  nor csa_tree_add_12_51_groupi_g14668__5526(csa_tree_add_12_51_groupi_n_7094 ,csa_tree_add_12_51_groupi_n_7006 ,csa_tree_add_12_51_groupi_n_7064);
  or csa_tree_add_12_51_groupi_g14669__6783(csa_tree_add_12_51_groupi_n_7093 ,csa_tree_add_12_51_groupi_n_7040 ,csa_tree_add_12_51_groupi_n_7073);
  nor csa_tree_add_12_51_groupi_g14670__3680(csa_tree_add_12_51_groupi_n_7092 ,csa_tree_add_12_51_groupi_n_7041 ,csa_tree_add_12_51_groupi_n_7074);
  and csa_tree_add_12_51_groupi_g14671__1617(csa_tree_add_12_51_groupi_n_7091 ,csa_tree_add_12_51_groupi_n_7023 ,csa_tree_add_12_51_groupi_n_7059);
  or csa_tree_add_12_51_groupi_g14672__2802(csa_tree_add_12_51_groupi_n_7090 ,csa_tree_add_12_51_groupi_n_7023 ,csa_tree_add_12_51_groupi_n_7059);
  or csa_tree_add_12_51_groupi_g14673__1705(csa_tree_add_12_51_groupi_n_7089 ,csa_tree_add_12_51_groupi_n_7043 ,csa_tree_add_12_51_groupi_n_7075);
  or csa_tree_add_12_51_groupi_g14674__5122(csa_tree_add_12_51_groupi_n_7088 ,csa_tree_add_12_51_groupi_n_7062 ,csa_tree_add_12_51_groupi_n_7060);
  or csa_tree_add_12_51_groupi_g14675__8246(csa_tree_add_12_51_groupi_n_7087 ,csa_tree_add_12_51_groupi_n_7005 ,csa_tree_add_12_51_groupi_n_7063);
  not csa_tree_add_12_51_groupi_g14676(csa_tree_add_12_51_groupi_n_7086 ,csa_tree_add_12_51_groupi_n_7085);
  not csa_tree_add_12_51_groupi_g14677(csa_tree_add_12_51_groupi_n_7080 ,csa_tree_add_12_51_groupi_n_7079);
  xnor csa_tree_add_12_51_groupi_g14678__7098(csa_tree_add_12_51_groupi_n_7076 ,csa_tree_add_12_51_groupi_n_7038 ,csa_tree_add_12_51_groupi_n_6990);
  xnor csa_tree_add_12_51_groupi_g14679__6131(csa_tree_add_12_51_groupi_n_7085 ,csa_tree_add_12_51_groupi_n_6991 ,csa_tree_add_12_51_groupi_n_7033);
  xnor csa_tree_add_12_51_groupi_g14680__1881(csa_tree_add_12_51_groupi_n_7084 ,csa_tree_add_12_51_groupi_n_6959 ,csa_tree_add_12_51_groupi_n_7031);
  xnor csa_tree_add_12_51_groupi_g14681__5115(csa_tree_add_12_51_groupi_n_7083 ,csa_tree_add_12_51_groupi_n_6958 ,csa_tree_add_12_51_groupi_n_7034);
  xnor csa_tree_add_12_51_groupi_g14682__7482(csa_tree_add_12_51_groupi_n_7082 ,csa_tree_add_12_51_groupi_n_7024 ,csa_tree_add_12_51_groupi_n_7030);
  xnor csa_tree_add_12_51_groupi_g14683__4733(csa_tree_add_12_51_groupi_n_7081 ,csa_tree_add_12_51_groupi_n_6943 ,csa_tree_add_12_51_groupi_n_7029);
  xnor csa_tree_add_12_51_groupi_g14684__6161(csa_tree_add_12_51_groupi_n_7079 ,csa_tree_add_12_51_groupi_n_6972 ,csa_tree_add_12_51_groupi_n_16);
  xnor csa_tree_add_12_51_groupi_g14685__9315(csa_tree_add_12_51_groupi_n_7078 ,csa_tree_add_12_51_groupi_n_7027 ,csa_tree_add_12_51_groupi_n_7028);
  xnor csa_tree_add_12_51_groupi_g14686__9945(csa_tree_add_12_51_groupi_n_7077 ,csa_tree_add_12_51_groupi_n_7009 ,csa_tree_add_12_51_groupi_n_7032);
  not csa_tree_add_12_51_groupi_g14687(csa_tree_add_12_51_groupi_n_7073 ,csa_tree_add_12_51_groupi_n_7074);
  not csa_tree_add_12_51_groupi_g14688(csa_tree_add_12_51_groupi_n_7068 ,csa_tree_add_12_51_groupi_n_7069);
  and csa_tree_add_12_51_groupi_g14689__2883(csa_tree_add_12_51_groupi_n_7066 ,csa_tree_add_12_51_groupi_n_7039 ,csa_tree_add_12_51_groupi_n_6990);
  nor csa_tree_add_12_51_groupi_g14690__2346(csa_tree_add_12_51_groupi_n_7065 ,csa_tree_add_12_51_groupi_n_7039 ,csa_tree_add_12_51_groupi_n_6990);
  and csa_tree_add_12_51_groupi_g14691__1666(csa_tree_add_12_51_groupi_n_7075 ,csa_tree_add_12_51_groupi_n_7044 ,csa_tree_add_12_51_groupi_n_6963);
  and csa_tree_add_12_51_groupi_g14692__7410(csa_tree_add_12_51_groupi_n_7074 ,csa_tree_add_12_51_groupi_n_7048 ,csa_tree_add_12_51_groupi_n_7018);
  or csa_tree_add_12_51_groupi_g14693__6417(csa_tree_add_12_51_groupi_n_7072 ,csa_tree_add_12_51_groupi_n_7047 ,csa_tree_add_12_51_groupi_n_7020);
  or csa_tree_add_12_51_groupi_g14694__5477(csa_tree_add_12_51_groupi_n_7071 ,csa_tree_add_12_51_groupi_n_6998 ,csa_tree_add_12_51_groupi_n_7051);
  or csa_tree_add_12_51_groupi_g14695__2398(csa_tree_add_12_51_groupi_n_7070 ,csa_tree_add_12_51_groupi_n_7017 ,csa_tree_add_12_51_groupi_n_7050);
  and csa_tree_add_12_51_groupi_g14696__5107(csa_tree_add_12_51_groupi_n_7069 ,csa_tree_add_12_51_groupi_n_7049 ,csa_tree_add_12_51_groupi_n_7014);
  or csa_tree_add_12_51_groupi_g14697__6260(csa_tree_add_12_51_groupi_n_7067 ,csa_tree_add_12_51_groupi_n_7046 ,csa_tree_add_12_51_groupi_n_7012);
  not csa_tree_add_12_51_groupi_g14698(csa_tree_add_12_51_groupi_n_7063 ,csa_tree_add_12_51_groupi_n_7064);
  xnor csa_tree_add_12_51_groupi_g14699__4319(out3[15] ,csa_tree_add_12_51_groupi_n_7025 ,csa_tree_add_12_51_groupi_n_6994);
  xnor csa_tree_add_12_51_groupi_g14700__8428(csa_tree_add_12_51_groupi_n_7056 ,csa_tree_add_12_51_groupi_n_7008 ,csa_tree_add_12_51_groupi_n_6922);
  xnor csa_tree_add_12_51_groupi_g14701__5526(csa_tree_add_12_51_groupi_n_7055 ,csa_tree_add_12_51_groupi_n_6938 ,csa_tree_add_12_51_groupi_n_7022);
  xnor csa_tree_add_12_51_groupi_g14702__6783(csa_tree_add_12_51_groupi_n_7064 ,csa_tree_add_12_51_groupi_n_6918 ,csa_tree_add_12_51_groupi_n_6996);
  xnor csa_tree_add_12_51_groupi_g14703__3680(csa_tree_add_12_51_groupi_n_7062 ,csa_tree_add_12_51_groupi_n_7010 ,csa_tree_add_12_51_groupi_n_6993);
  or csa_tree_add_12_51_groupi_g14704__1617(csa_tree_add_12_51_groupi_n_7061 ,csa_tree_add_12_51_groupi_n_6965 ,csa_tree_add_12_51_groupi_n_7036);
  or csa_tree_add_12_51_groupi_g14705__2802(csa_tree_add_12_51_groupi_n_7060 ,csa_tree_add_12_51_groupi_n_7035 ,csa_tree_add_12_51_groupi_n_6999);
  xnor csa_tree_add_12_51_groupi_g14706__1705(csa_tree_add_12_51_groupi_n_7059 ,csa_tree_add_12_51_groupi_n_6967 ,csa_tree_add_12_51_groupi_n_6997);
  or csa_tree_add_12_51_groupi_g14707__5122(csa_tree_add_12_51_groupi_n_7058 ,csa_tree_add_12_51_groupi_n_7037 ,csa_tree_add_12_51_groupi_n_7001);
  not csa_tree_add_12_51_groupi_g14708(csa_tree_add_12_51_groupi_n_7053 ,csa_tree_add_12_51_groupi_n_7054);
  and csa_tree_add_12_51_groupi_g14709__8246(csa_tree_add_12_51_groupi_n_7052 ,csa_tree_add_12_51_groupi_n_6939 ,csa_tree_add_12_51_groupi_n_7022);
  and csa_tree_add_12_51_groupi_g14710__7098(csa_tree_add_12_51_groupi_n_7051 ,csa_tree_add_12_51_groupi_n_7003 ,csa_tree_add_12_51_groupi_n_7009);
  nor csa_tree_add_12_51_groupi_g14711__6131(csa_tree_add_12_51_groupi_n_7050 ,csa_tree_add_12_51_groupi_n_7016 ,csa_tree_add_12_51_groupi_n_6943);
  or csa_tree_add_12_51_groupi_g14712__1881(csa_tree_add_12_51_groupi_n_7049 ,csa_tree_add_12_51_groupi_n_6940 ,csa_tree_add_12_51_groupi_n_7011);
  or csa_tree_add_12_51_groupi_g14713__5115(csa_tree_add_12_51_groupi_n_7048 ,csa_tree_add_12_51_groupi_n_6959 ,csa_tree_add_12_51_groupi_n_7015);
  and csa_tree_add_12_51_groupi_g14714__7482(csa_tree_add_12_51_groupi_n_7047 ,csa_tree_add_12_51_groupi_n_7021 ,csa_tree_add_12_51_groupi_n_7024);
  nor csa_tree_add_12_51_groupi_g14715__4733(csa_tree_add_12_51_groupi_n_7046 ,csa_tree_add_12_51_groupi_n_7013 ,csa_tree_add_12_51_groupi_n_6992);
  nor csa_tree_add_12_51_groupi_g14716__6161(csa_tree_add_12_51_groupi_n_7045 ,csa_tree_add_12_51_groupi_n_6939 ,csa_tree_add_12_51_groupi_n_7022);
  or csa_tree_add_12_51_groupi_g14717__9315(csa_tree_add_12_51_groupi_n_7044 ,csa_tree_add_12_51_groupi_n_6988 ,csa_tree_add_12_51_groupi_n_7026);
  nor csa_tree_add_12_51_groupi_g14718__9945(csa_tree_add_12_51_groupi_n_7043 ,csa_tree_add_12_51_groupi_n_7007 ,csa_tree_add_12_51_groupi_n_6922);
  or csa_tree_add_12_51_groupi_g14719__2883(csa_tree_add_12_51_groupi_n_7042 ,csa_tree_add_12_51_groupi_n_7008 ,csa_tree_add_12_51_groupi_n_6921);
  and csa_tree_add_12_51_groupi_g14720__2346(csa_tree_add_12_51_groupi_n_7054 ,csa_tree_add_12_51_groupi_n_6980 ,csa_tree_add_12_51_groupi_n_7019);
  not csa_tree_add_12_51_groupi_g14721(csa_tree_add_12_51_groupi_n_7041 ,csa_tree_add_12_51_groupi_n_7040);
  not csa_tree_add_12_51_groupi_g14722(csa_tree_add_12_51_groupi_n_7039 ,csa_tree_add_12_51_groupi_n_7038);
  nor csa_tree_add_12_51_groupi_g14723__1666(csa_tree_add_12_51_groupi_n_7037 ,csa_tree_add_12_51_groupi_n_7027 ,csa_tree_add_12_51_groupi_n_7002);
  nor csa_tree_add_12_51_groupi_g14724__7410(csa_tree_add_12_51_groupi_n_7036 ,csa_tree_add_12_51_groupi_n_6966 ,csa_tree_add_12_51_groupi_n_7010);
  nor csa_tree_add_12_51_groupi_g14725__6417(csa_tree_add_12_51_groupi_n_7035 ,csa_tree_add_12_51_groupi_n_6991 ,csa_tree_add_12_51_groupi_n_7000);
  xnor csa_tree_add_12_51_groupi_g14727__5477(csa_tree_add_12_51_groupi_n_7034 ,csa_tree_add_12_51_groupi_n_6978 ,csa_tree_add_12_51_groupi_n_6920);
  xnor csa_tree_add_12_51_groupi_g14728__2398(csa_tree_add_12_51_groupi_n_7033 ,csa_tree_add_12_51_groupi_n_6894 ,csa_tree_add_12_51_groupi_n_6973);
  xnor csa_tree_add_12_51_groupi_g14729__5107(csa_tree_add_12_51_groupi_n_7032 ,csa_tree_add_12_51_groupi_n_6989 ,csa_tree_add_12_51_groupi_n_6900);
  xnor csa_tree_add_12_51_groupi_g14730__6260(csa_tree_add_12_51_groupi_n_7031 ,csa_tree_add_12_51_groupi_n_6969 ,csa_tree_add_12_51_groupi_n_6818);
  xnor csa_tree_add_12_51_groupi_g14731__4319(csa_tree_add_12_51_groupi_n_7030 ,csa_tree_add_12_51_groupi_n_6971 ,csa_tree_add_12_51_groupi_n_6937);
  xnor csa_tree_add_12_51_groupi_g14732__8428(csa_tree_add_12_51_groupi_n_7029 ,csa_tree_add_12_51_groupi_n_6882 ,csa_tree_add_12_51_groupi_n_6977);
  xnor csa_tree_add_12_51_groupi_g14733__5526(csa_tree_add_12_51_groupi_n_7028 ,csa_tree_add_12_51_groupi_n_6895 ,csa_tree_add_12_51_groupi_n_6975);
  xnor csa_tree_add_12_51_groupi_g14734__6783(csa_tree_add_12_51_groupi_n_7040 ,csa_tree_add_12_51_groupi_n_6923 ,csa_tree_add_12_51_groupi_n_6962);
  xnor csa_tree_add_12_51_groupi_g14735__3680(csa_tree_add_12_51_groupi_n_7038 ,csa_tree_add_12_51_groupi_n_6941 ,csa_tree_add_12_51_groupi_n_6961);
  not csa_tree_add_12_51_groupi_g14736(csa_tree_add_12_51_groupi_n_7026 ,csa_tree_add_12_51_groupi_n_7025);
  or csa_tree_add_12_51_groupi_g14737__1617(csa_tree_add_12_51_groupi_n_7021 ,csa_tree_add_12_51_groupi_n_2354 ,csa_tree_add_12_51_groupi_n_6970);
  nor csa_tree_add_12_51_groupi_g14738__2802(csa_tree_add_12_51_groupi_n_7020 ,csa_tree_add_12_51_groupi_n_2151 ,csa_tree_add_12_51_groupi_n_6971);
  or csa_tree_add_12_51_groupi_g14739__1705(csa_tree_add_12_51_groupi_n_7019 ,csa_tree_add_12_51_groupi_n_6979 ,csa_tree_add_12_51_groupi_n_6978);
  or csa_tree_add_12_51_groupi_g14740__5122(csa_tree_add_12_51_groupi_n_7018 ,csa_tree_add_12_51_groupi_n_6968 ,csa_tree_add_12_51_groupi_n_6818);
  nor csa_tree_add_12_51_groupi_g14741__8246(csa_tree_add_12_51_groupi_n_7017 ,csa_tree_add_12_51_groupi_n_6883 ,csa_tree_add_12_51_groupi_n_6977);
  and csa_tree_add_12_51_groupi_g14742__7098(csa_tree_add_12_51_groupi_n_7016 ,csa_tree_add_12_51_groupi_n_6883 ,csa_tree_add_12_51_groupi_n_6977);
  nor csa_tree_add_12_51_groupi_g14743__6131(csa_tree_add_12_51_groupi_n_7015 ,csa_tree_add_12_51_groupi_n_6969 ,csa_tree_add_12_51_groupi_n_6817);
  or csa_tree_add_12_51_groupi_g14744__1881(csa_tree_add_12_51_groupi_n_7014 ,csa_tree_add_12_51_groupi_n_6884 ,csa_tree_add_12_51_groupi_n_6967);
  and csa_tree_add_12_51_groupi_g14745__5115(csa_tree_add_12_51_groupi_n_7013 ,csa_tree_add_12_51_groupi_n_6749 ,csa_tree_add_12_51_groupi_n_6972);
  nor csa_tree_add_12_51_groupi_g14746__7482(csa_tree_add_12_51_groupi_n_7012 ,csa_tree_add_12_51_groupi_n_6749 ,csa_tree_add_12_51_groupi_n_6972);
  and csa_tree_add_12_51_groupi_g14747__4733(csa_tree_add_12_51_groupi_n_7011 ,csa_tree_add_12_51_groupi_n_6884 ,csa_tree_add_12_51_groupi_n_6967);
  and csa_tree_add_12_51_groupi_g14748__6161(csa_tree_add_12_51_groupi_n_7027 ,csa_tree_add_12_51_groupi_n_6944 ,csa_tree_add_12_51_groupi_n_6983);
  or csa_tree_add_12_51_groupi_g14749__9315(csa_tree_add_12_51_groupi_n_7025 ,csa_tree_add_12_51_groupi_n_6912 ,csa_tree_add_12_51_groupi_n_6985);
  or csa_tree_add_12_51_groupi_g14750__9945(csa_tree_add_12_51_groupi_n_7024 ,csa_tree_add_12_51_groupi_n_6953 ,csa_tree_add_12_51_groupi_n_6981);
  or csa_tree_add_12_51_groupi_g14751__2883(csa_tree_add_12_51_groupi_n_7023 ,csa_tree_add_12_51_groupi_n_6987 ,csa_tree_add_12_51_groupi_n_6952);
  and csa_tree_add_12_51_groupi_g14752__2346(csa_tree_add_12_51_groupi_n_7022 ,csa_tree_add_12_51_groupi_n_6946 ,csa_tree_add_12_51_groupi_n_6982);
  not csa_tree_add_12_51_groupi_g14753(csa_tree_add_12_51_groupi_n_7007 ,csa_tree_add_12_51_groupi_n_7008);
  not csa_tree_add_12_51_groupi_g14754(csa_tree_add_12_51_groupi_n_7006 ,csa_tree_add_12_51_groupi_n_7005);
  xnor csa_tree_add_12_51_groupi_g14755__1666(out3[14] ,csa_tree_add_12_51_groupi_n_6960 ,csa_tree_add_12_51_groupi_n_6928);
  or csa_tree_add_12_51_groupi_g14756__7410(csa_tree_add_12_51_groupi_n_7003 ,csa_tree_add_12_51_groupi_n_6989 ,csa_tree_add_12_51_groupi_n_6900);
  and csa_tree_add_12_51_groupi_g14757__6417(csa_tree_add_12_51_groupi_n_7002 ,csa_tree_add_12_51_groupi_n_6895 ,csa_tree_add_12_51_groupi_n_6976);
  nor csa_tree_add_12_51_groupi_g14758__5477(csa_tree_add_12_51_groupi_n_7001 ,csa_tree_add_12_51_groupi_n_6895 ,csa_tree_add_12_51_groupi_n_6976);
  and csa_tree_add_12_51_groupi_g14759__2398(csa_tree_add_12_51_groupi_n_7000 ,csa_tree_add_12_51_groupi_n_6894 ,csa_tree_add_12_51_groupi_n_6974);
  nor csa_tree_add_12_51_groupi_g14760__5107(csa_tree_add_12_51_groupi_n_6999 ,csa_tree_add_12_51_groupi_n_6894 ,csa_tree_add_12_51_groupi_n_6974);
  and csa_tree_add_12_51_groupi_g14761__6260(csa_tree_add_12_51_groupi_n_6998 ,csa_tree_add_12_51_groupi_n_6989 ,csa_tree_add_12_51_groupi_n_6900);
  xor csa_tree_add_12_51_groupi_g14762__4319(csa_tree_add_12_51_groupi_n_6997 ,csa_tree_add_12_51_groupi_n_6884 ,csa_tree_add_12_51_groupi_n_6940);
  xnor csa_tree_add_12_51_groupi_g14763__8428(csa_tree_add_12_51_groupi_n_6996 ,csa_tree_add_12_51_groupi_n_6942 ,csa_tree_add_12_51_groupi_n_6748);
  xnor csa_tree_add_12_51_groupi_g14764__5526(csa_tree_add_12_51_groupi_n_6995 ,csa_tree_add_12_51_groupi_n_5186 ,csa_tree_add_12_51_groupi_n_6956);
  xnor csa_tree_add_12_51_groupi_g14765__6783(csa_tree_add_12_51_groupi_n_6994 ,csa_tree_add_12_51_groupi_n_6807 ,csa_tree_add_12_51_groupi_n_6936);
  xnor csa_tree_add_12_51_groupi_g14766__3680(csa_tree_add_12_51_groupi_n_6993 ,csa_tree_add_12_51_groupi_n_6934 ,csa_tree_add_12_51_groupi_n_6811);
  xnor csa_tree_add_12_51_groupi_g14767__1617(csa_tree_add_12_51_groupi_n_7010 ,csa_tree_add_12_51_groupi_n_6899 ,csa_tree_add_12_51_groupi_n_6926);
  xnor csa_tree_add_12_51_groupi_g14768__2802(csa_tree_add_12_51_groupi_n_7009 ,csa_tree_add_12_51_groupi_n_6901 ,csa_tree_add_12_51_groupi_n_6927);
  xnor csa_tree_add_12_51_groupi_g14769__1705(csa_tree_add_12_51_groupi_n_7008 ,csa_tree_add_12_51_groupi_n_6903 ,csa_tree_add_12_51_groupi_n_6929);
  and csa_tree_add_12_51_groupi_g14770__5122(csa_tree_add_12_51_groupi_n_7005 ,csa_tree_add_12_51_groupi_n_6964 ,csa_tree_add_12_51_groupi_n_6931);
  nor csa_tree_add_12_51_groupi_g14771__8246(csa_tree_add_12_51_groupi_n_6988 ,csa_tree_add_12_51_groupi_n_6807 ,csa_tree_add_12_51_groupi_n_6936);
  and csa_tree_add_12_51_groupi_g14772__7098(csa_tree_add_12_51_groupi_n_6987 ,csa_tree_add_12_51_groupi_n_6941 ,csa_tree_add_12_51_groupi_n_6947);
  nor csa_tree_add_12_51_groupi_g14773__6131(csa_tree_add_12_51_groupi_n_6986 ,csa_tree_add_12_51_groupi_n_5186 ,csa_tree_add_12_51_groupi_n_6956);
  and csa_tree_add_12_51_groupi_g14774__1881(csa_tree_add_12_51_groupi_n_6985 ,csa_tree_add_12_51_groupi_n_6960 ,csa_tree_add_12_51_groupi_n_6911);
  or csa_tree_add_12_51_groupi_g14775__5115(csa_tree_add_12_51_groupi_n_6984 ,csa_tree_add_12_51_groupi_n_5185 ,csa_tree_add_12_51_groupi_n_6955);
  or csa_tree_add_12_51_groupi_g14776__7482(csa_tree_add_12_51_groupi_n_6983 ,csa_tree_add_12_51_groupi_n_6886 ,csa_tree_add_12_51_groupi_n_6948);
  or csa_tree_add_12_51_groupi_g14777__4733(csa_tree_add_12_51_groupi_n_6982 ,csa_tree_add_12_51_groupi_n_6942 ,csa_tree_add_12_51_groupi_n_6945);
  nor csa_tree_add_12_51_groupi_g14778__6161(csa_tree_add_12_51_groupi_n_6981 ,csa_tree_add_12_51_groupi_n_6950 ,csa_tree_add_12_51_groupi_n_6885);
  or csa_tree_add_12_51_groupi_g14779__9315(csa_tree_add_12_51_groupi_n_6980 ,csa_tree_add_12_51_groupi_n_6958 ,csa_tree_add_12_51_groupi_n_6919);
  nor csa_tree_add_12_51_groupi_g14780__9945(csa_tree_add_12_51_groupi_n_6979 ,csa_tree_add_12_51_groupi_n_6957 ,csa_tree_add_12_51_groupi_n_6920);
  and csa_tree_add_12_51_groupi_g14781__2883(csa_tree_add_12_51_groupi_n_6992 ,csa_tree_add_12_51_groupi_n_6930 ,csa_tree_add_12_51_groupi_n_6872);
  and csa_tree_add_12_51_groupi_g14782__2346(csa_tree_add_12_51_groupi_n_6991 ,csa_tree_add_12_51_groupi_n_6954 ,csa_tree_add_12_51_groupi_n_6873);
  and csa_tree_add_12_51_groupi_g14783__1666(csa_tree_add_12_51_groupi_n_6990 ,csa_tree_add_12_51_groupi_n_6949 ,csa_tree_add_12_51_groupi_n_6908);
  or csa_tree_add_12_51_groupi_g14784__7410(csa_tree_add_12_51_groupi_n_6989 ,csa_tree_add_12_51_groupi_n_6951 ,csa_tree_add_12_51_groupi_n_6877);
  not csa_tree_add_12_51_groupi_g14785(csa_tree_add_12_51_groupi_n_6976 ,csa_tree_add_12_51_groupi_n_6975);
  not csa_tree_add_12_51_groupi_g14786(csa_tree_add_12_51_groupi_n_6974 ,csa_tree_add_12_51_groupi_n_6973);
  not csa_tree_add_12_51_groupi_g14787(csa_tree_add_12_51_groupi_n_6971 ,csa_tree_add_12_51_groupi_n_6970);
  not csa_tree_add_12_51_groupi_g14788(csa_tree_add_12_51_groupi_n_6969 ,csa_tree_add_12_51_groupi_n_6968);
  and csa_tree_add_12_51_groupi_g14789__6417(csa_tree_add_12_51_groupi_n_6966 ,csa_tree_add_12_51_groupi_n_6934 ,csa_tree_add_12_51_groupi_n_6812);
  nor csa_tree_add_12_51_groupi_g14790__5477(csa_tree_add_12_51_groupi_n_6965 ,csa_tree_add_12_51_groupi_n_6934 ,csa_tree_add_12_51_groupi_n_6812);
  or csa_tree_add_12_51_groupi_g14791__2398(csa_tree_add_12_51_groupi_n_6964 ,csa_tree_add_12_51_groupi_n_6923 ,csa_tree_add_12_51_groupi_n_6932);
  or csa_tree_add_12_51_groupi_g14792__5107(csa_tree_add_12_51_groupi_n_6963 ,csa_tree_add_12_51_groupi_n_6806 ,csa_tree_add_12_51_groupi_n_6935);
  xnor csa_tree_add_12_51_groupi_g14793__6260(csa_tree_add_12_51_groupi_n_6962 ,csa_tree_add_12_51_groupi_n_6820 ,csa_tree_add_12_51_groupi_n_6897);
  xnor csa_tree_add_12_51_groupi_g14794__4319(csa_tree_add_12_51_groupi_n_6961 ,csa_tree_add_12_51_groupi_n_6916 ,csa_tree_add_12_51_groupi_n_6859);
  xnor csa_tree_add_12_51_groupi_g14795__8428(csa_tree_add_12_51_groupi_n_6978 ,csa_tree_add_12_51_groupi_n_6924 ,csa_tree_add_12_51_groupi_n_6893);
  xnor csa_tree_add_12_51_groupi_g14796__5526(csa_tree_add_12_51_groupi_n_6977 ,csa_tree_add_12_51_groupi_n_6902 ,csa_tree_add_12_51_groupi_n_6892);
  xnor csa_tree_add_12_51_groupi_g14797__6783(csa_tree_add_12_51_groupi_n_6975 ,csa_tree_add_12_51_groupi_n_6846 ,csa_tree_add_12_51_groupi_n_6887);
  xnor csa_tree_add_12_51_groupi_g14798__3680(csa_tree_add_12_51_groupi_n_6973 ,csa_tree_add_12_51_groupi_n_6863 ,csa_tree_add_12_51_groupi_n_6888);
  xnor csa_tree_add_12_51_groupi_g14799__1617(csa_tree_add_12_51_groupi_n_6972 ,csa_tree_add_12_51_groupi_n_6867 ,csa_tree_add_12_51_groupi_n_6891);
  xnor csa_tree_add_12_51_groupi_g14800__2802(csa_tree_add_12_51_groupi_n_6970 ,csa_tree_add_12_51_groupi_n_6821 ,csa_tree_add_12_51_groupi_n_6889);
  xnor csa_tree_add_12_51_groupi_g14801__1705(csa_tree_add_12_51_groupi_n_6968 ,csa_tree_add_12_51_groupi_n_6726 ,csa_tree_add_12_51_groupi_n_17);
  xnor csa_tree_add_12_51_groupi_g14802__5122(csa_tree_add_12_51_groupi_n_6967 ,csa_tree_add_12_51_groupi_n_6904 ,csa_tree_add_12_51_groupi_n_6890);
  not csa_tree_add_12_51_groupi_g14803(csa_tree_add_12_51_groupi_n_6958 ,csa_tree_add_12_51_groupi_n_6957);
  not csa_tree_add_12_51_groupi_g14804(csa_tree_add_12_51_groupi_n_6955 ,csa_tree_add_12_51_groupi_n_6956);
  or csa_tree_add_12_51_groupi_g14805__8246(csa_tree_add_12_51_groupi_n_6954 ,csa_tree_add_12_51_groupi_n_6904 ,csa_tree_add_12_51_groupi_n_6874);
  and csa_tree_add_12_51_groupi_g14806__7098(csa_tree_add_12_51_groupi_n_6953 ,csa_tree_add_12_51_groupi_n_6901 ,csa_tree_add_12_51_groupi_n_6784);
  and csa_tree_add_12_51_groupi_g14807__6131(csa_tree_add_12_51_groupi_n_6952 ,csa_tree_add_12_51_groupi_n_6916 ,csa_tree_add_12_51_groupi_n_6859);
  nor csa_tree_add_12_51_groupi_g14808__1881(csa_tree_add_12_51_groupi_n_6951 ,csa_tree_add_12_51_groupi_n_6878 ,csa_tree_add_12_51_groupi_n_6902);
  nor csa_tree_add_12_51_groupi_g14809__5115(csa_tree_add_12_51_groupi_n_6950 ,csa_tree_add_12_51_groupi_n_6901 ,csa_tree_add_12_51_groupi_n_6784);
  or csa_tree_add_12_51_groupi_g14810__7482(csa_tree_add_12_51_groupi_n_6949 ,csa_tree_add_12_51_groupi_n_6909 ,csa_tree_add_12_51_groupi_n_6903);
  nor csa_tree_add_12_51_groupi_g14811__4733(csa_tree_add_12_51_groupi_n_6948 ,csa_tree_add_12_51_groupi_n_6899 ,csa_tree_add_12_51_groupi_n_6781);
  or csa_tree_add_12_51_groupi_g14812__6161(csa_tree_add_12_51_groupi_n_6947 ,csa_tree_add_12_51_groupi_n_6916 ,csa_tree_add_12_51_groupi_n_6859);
  or csa_tree_add_12_51_groupi_g14813__9315(csa_tree_add_12_51_groupi_n_6946 ,csa_tree_add_12_51_groupi_n_6748 ,csa_tree_add_12_51_groupi_n_6917);
  nor csa_tree_add_12_51_groupi_g14814__9945(csa_tree_add_12_51_groupi_n_6945 ,csa_tree_add_12_51_groupi_n_6747 ,csa_tree_add_12_51_groupi_n_6918);
  or csa_tree_add_12_51_groupi_g14815__2883(csa_tree_add_12_51_groupi_n_6944 ,csa_tree_add_12_51_groupi_n_6898 ,csa_tree_add_12_51_groupi_n_6780);
  or csa_tree_add_12_51_groupi_g14816__2346(csa_tree_add_12_51_groupi_n_6960 ,csa_tree_add_12_51_groupi_n_6833 ,csa_tree_add_12_51_groupi_n_6910);
  and csa_tree_add_12_51_groupi_g14817__1666(csa_tree_add_12_51_groupi_n_6959 ,csa_tree_add_12_51_groupi_n_6915 ,csa_tree_add_12_51_groupi_n_6869);
  or csa_tree_add_12_51_groupi_g14818__7410(csa_tree_add_12_51_groupi_n_6957 ,csa_tree_add_12_51_groupi_n_6875 ,csa_tree_add_12_51_groupi_n_6905);
  or csa_tree_add_12_51_groupi_g14819__6417(csa_tree_add_12_51_groupi_n_6956 ,csa_tree_add_12_51_groupi_n_6764 ,csa_tree_add_12_51_groupi_n_6913);
  not csa_tree_add_12_51_groupi_g14820(csa_tree_add_12_51_groupi_n_6939 ,csa_tree_add_12_51_groupi_n_6938);
  not csa_tree_add_12_51_groupi_g14822(csa_tree_add_12_51_groupi_n_6935 ,csa_tree_add_12_51_groupi_n_6936);
  xnor csa_tree_add_12_51_groupi_g14823__5477(out3[13] ,csa_tree_add_12_51_groupi_n_6866 ,csa_tree_add_12_51_groupi_n_6850);
  nor csa_tree_add_12_51_groupi_g14824__2398(csa_tree_add_12_51_groupi_n_6932 ,csa_tree_add_12_51_groupi_n_6820 ,csa_tree_add_12_51_groupi_n_6896);
  or csa_tree_add_12_51_groupi_g14825__5107(csa_tree_add_12_51_groupi_n_6931 ,csa_tree_add_12_51_groupi_n_6819 ,csa_tree_add_12_51_groupi_n_6897);
  or csa_tree_add_12_51_groupi_g14826__6260(csa_tree_add_12_51_groupi_n_6930 ,csa_tree_add_12_51_groupi_n_6925 ,csa_tree_add_12_51_groupi_n_6868);
  xnor csa_tree_add_12_51_groupi_g14827__4319(csa_tree_add_12_51_groupi_n_6929 ,csa_tree_add_12_51_groupi_n_6862 ,csa_tree_add_12_51_groupi_n_6786);
  xnor csa_tree_add_12_51_groupi_g14828__8428(csa_tree_add_12_51_groupi_n_6928 ,csa_tree_add_12_51_groupi_n_6860 ,csa_tree_add_12_51_groupi_n_6787);
  xor csa_tree_add_12_51_groupi_g14829__5526(csa_tree_add_12_51_groupi_n_6927 ,csa_tree_add_12_51_groupi_n_6885 ,csa_tree_add_12_51_groupi_n_6784);
  xnor csa_tree_add_12_51_groupi_g14830__6783(csa_tree_add_12_51_groupi_n_6926 ,csa_tree_add_12_51_groupi_n_6886 ,csa_tree_add_12_51_groupi_n_6781);
  and csa_tree_add_12_51_groupi_g14831__3680(csa_tree_add_12_51_groupi_n_6943 ,csa_tree_add_12_51_groupi_n_6914 ,csa_tree_add_12_51_groupi_n_6854);
  xnor csa_tree_add_12_51_groupi_g14832__1617(csa_tree_add_12_51_groupi_n_6942 ,csa_tree_add_12_51_groupi_n_5024 ,csa_tree_add_12_51_groupi_n_6851);
  xnor csa_tree_add_12_51_groupi_g14833__2802(csa_tree_add_12_51_groupi_n_6941 ,csa_tree_add_12_51_groupi_n_6864 ,csa_tree_add_12_51_groupi_n_6849);
  and csa_tree_add_12_51_groupi_g14834__1705(csa_tree_add_12_51_groupi_n_6940 ,csa_tree_add_12_51_groupi_n_6907 ,csa_tree_add_12_51_groupi_n_6827);
  xnor csa_tree_add_12_51_groupi_g14835__5122(csa_tree_add_12_51_groupi_n_6938 ,csa_tree_add_12_51_groupi_n_6865 ,csa_tree_add_12_51_groupi_n_6797);
  xnor csa_tree_add_12_51_groupi_g14836__8246(csa_tree_add_12_51_groupi_n_6937 ,csa_tree_add_12_51_groupi_n_6759 ,csa_tree_add_12_51_groupi_n_6848);
  xnor csa_tree_add_12_51_groupi_g14837__7098(csa_tree_add_12_51_groupi_n_6936 ,csa_tree_add_12_51_groupi_n_6822 ,csa_tree_add_12_51_groupi_n_6852);
  and csa_tree_add_12_51_groupi_g14838__6131(csa_tree_add_12_51_groupi_n_6934 ,csa_tree_add_12_51_groupi_n_6906 ,csa_tree_add_12_51_groupi_n_6857);
  not csa_tree_add_12_51_groupi_g14839(csa_tree_add_12_51_groupi_n_6925 ,csa_tree_add_12_51_groupi_n_6924);
  not csa_tree_add_12_51_groupi_g14840(csa_tree_add_12_51_groupi_n_6921 ,csa_tree_add_12_51_groupi_n_6922);
  not csa_tree_add_12_51_groupi_g14841(csa_tree_add_12_51_groupi_n_6919 ,csa_tree_add_12_51_groupi_n_6920);
  not csa_tree_add_12_51_groupi_g14842(csa_tree_add_12_51_groupi_n_6917 ,csa_tree_add_12_51_groupi_n_6918);
  or csa_tree_add_12_51_groupi_g14843__1881(csa_tree_add_12_51_groupi_n_6915 ,csa_tree_add_12_51_groupi_n_6870 ,csa_tree_add_12_51_groupi_n_6867);
  or csa_tree_add_12_51_groupi_g14844__5115(csa_tree_add_12_51_groupi_n_6914 ,csa_tree_add_12_51_groupi_n_6846 ,csa_tree_add_12_51_groupi_n_6855);
  and csa_tree_add_12_51_groupi_g14845__7482(csa_tree_add_12_51_groupi_n_6913 ,csa_tree_add_12_51_groupi_n_6778 ,csa_tree_add_12_51_groupi_n_6865);
  and csa_tree_add_12_51_groupi_g14846__4733(csa_tree_add_12_51_groupi_n_6912 ,csa_tree_add_12_51_groupi_n_6860 ,csa_tree_add_12_51_groupi_n_6787);
  or csa_tree_add_12_51_groupi_g14847__6161(csa_tree_add_12_51_groupi_n_6911 ,csa_tree_add_12_51_groupi_n_6860 ,csa_tree_add_12_51_groupi_n_6787);
  and csa_tree_add_12_51_groupi_g14848__9315(csa_tree_add_12_51_groupi_n_6910 ,csa_tree_add_12_51_groupi_n_6866 ,csa_tree_add_12_51_groupi_n_6832);
  nor csa_tree_add_12_51_groupi_g14849__9945(csa_tree_add_12_51_groupi_n_6909 ,csa_tree_add_12_51_groupi_n_6862 ,csa_tree_add_12_51_groupi_n_6786);
  or csa_tree_add_12_51_groupi_g14850__2883(csa_tree_add_12_51_groupi_n_6908 ,csa_tree_add_12_51_groupi_n_6861 ,csa_tree_add_12_51_groupi_n_6785);
  or csa_tree_add_12_51_groupi_g14851__2346(csa_tree_add_12_51_groupi_n_6907 ,csa_tree_add_12_51_groupi_n_6864 ,csa_tree_add_12_51_groupi_n_6826);
  or csa_tree_add_12_51_groupi_g14852__1666(csa_tree_add_12_51_groupi_n_6906 ,csa_tree_add_12_51_groupi_n_6863 ,csa_tree_add_12_51_groupi_n_6858);
  nor csa_tree_add_12_51_groupi_g14853__7410(csa_tree_add_12_51_groupi_n_6905 ,csa_tree_add_12_51_groupi_n_6876 ,csa_tree_add_12_51_groupi_n_6821);
  or csa_tree_add_12_51_groupi_g14854__6417(csa_tree_add_12_51_groupi_n_6924 ,csa_tree_add_12_51_groupi_n_6823 ,csa_tree_add_12_51_groupi_n_6880);
  and csa_tree_add_12_51_groupi_g14855__5477(csa_tree_add_12_51_groupi_n_6923 ,csa_tree_add_12_51_groupi_n_6829 ,csa_tree_add_12_51_groupi_n_6856);
  or csa_tree_add_12_51_groupi_g14856__2398(csa_tree_add_12_51_groupi_n_6922 ,csa_tree_add_12_51_groupi_n_6839 ,csa_tree_add_12_51_groupi_n_6879);
  xnor csa_tree_add_12_51_groupi_g14857__5107(csa_tree_add_12_51_groupi_n_6920 ,csa_tree_add_12_51_groupi_n_6634 ,csa_tree_add_12_51_groupi_n_6794);
  or csa_tree_add_12_51_groupi_g14858__6260(csa_tree_add_12_51_groupi_n_6918 ,csa_tree_add_12_51_groupi_n_6831 ,csa_tree_add_12_51_groupi_n_6881);
  or csa_tree_add_12_51_groupi_g14859__4319(csa_tree_add_12_51_groupi_n_6916 ,csa_tree_add_12_51_groupi_n_6871 ,csa_tree_add_12_51_groupi_n_6825);
  not csa_tree_add_12_51_groupi_g14860(csa_tree_add_12_51_groupi_n_6898 ,csa_tree_add_12_51_groupi_n_6899);
  not csa_tree_add_12_51_groupi_g14861(csa_tree_add_12_51_groupi_n_6896 ,csa_tree_add_12_51_groupi_n_6897);
  xnor csa_tree_add_12_51_groupi_g14862__8428(csa_tree_add_12_51_groupi_n_6893 ,csa_tree_add_12_51_groupi_n_6816 ,csa_tree_add_12_51_groupi_n_6720);
  xnor csa_tree_add_12_51_groupi_g14863__5526(csa_tree_add_12_51_groupi_n_6892 ,csa_tree_add_12_51_groupi_n_6715 ,csa_tree_add_12_51_groupi_n_6810);
  xnor csa_tree_add_12_51_groupi_g14865__6783(csa_tree_add_12_51_groupi_n_6891 ,csa_tree_add_12_51_groupi_n_6789 ,csa_tree_add_12_51_groupi_n_6843);
  xnor csa_tree_add_12_51_groupi_g14866__3680(csa_tree_add_12_51_groupi_n_6890 ,csa_tree_add_12_51_groupi_n_6746 ,csa_tree_add_12_51_groupi_n_6845);
  xnor csa_tree_add_12_51_groupi_g14867__1617(csa_tree_add_12_51_groupi_n_6889 ,csa_tree_add_12_51_groupi_n_6841 ,csa_tree_add_12_51_groupi_n_6713);
  xnor csa_tree_add_12_51_groupi_g14868__2802(csa_tree_add_12_51_groupi_n_6888 ,csa_tree_add_12_51_groupi_n_6809 ,csa_tree_add_12_51_groupi_n_6690);
  xnor csa_tree_add_12_51_groupi_g14869__1705(csa_tree_add_12_51_groupi_n_6887 ,csa_tree_add_12_51_groupi_n_6744 ,csa_tree_add_12_51_groupi_n_6814);
  xnor csa_tree_add_12_51_groupi_g14870__5122(csa_tree_add_12_51_groupi_n_6904 ,csa_tree_add_12_51_groupi_n_6762 ,csa_tree_add_12_51_groupi_n_6799);
  xnor csa_tree_add_12_51_groupi_g14871__8246(csa_tree_add_12_51_groupi_n_6903 ,csa_tree_add_12_51_groupi_n_6753 ,csa_tree_add_12_51_groupi_n_6793);
  xnor csa_tree_add_12_51_groupi_g14872__7098(csa_tree_add_12_51_groupi_n_6902 ,csa_tree_add_12_51_groupi_n_6760 ,csa_tree_add_12_51_groupi_n_6796);
  xnor csa_tree_add_12_51_groupi_g14873__6131(csa_tree_add_12_51_groupi_n_6901 ,csa_tree_add_12_51_groupi_n_6465 ,csa_tree_add_12_51_groupi_n_6802);
  xnor csa_tree_add_12_51_groupi_g14874__1881(csa_tree_add_12_51_groupi_n_6900 ,csa_tree_add_12_51_groupi_n_6442 ,csa_tree_add_12_51_groupi_n_15);
  xnor csa_tree_add_12_51_groupi_g14875__5115(csa_tree_add_12_51_groupi_n_6899 ,csa_tree_add_12_51_groupi_n_6463 ,csa_tree_add_12_51_groupi_n_6801);
  xnor csa_tree_add_12_51_groupi_g14876__7482(csa_tree_add_12_51_groupi_n_6897 ,csa_tree_add_12_51_groupi_n_6779 ,csa_tree_add_12_51_groupi_n_6798);
  xnor csa_tree_add_12_51_groupi_g14877__4733(csa_tree_add_12_51_groupi_n_6895 ,csa_tree_add_12_51_groupi_n_6758 ,csa_tree_add_12_51_groupi_n_6800);
  xnor csa_tree_add_12_51_groupi_g14878__6161(csa_tree_add_12_51_groupi_n_6894 ,csa_tree_add_12_51_groupi_n_6761 ,csa_tree_add_12_51_groupi_n_6795);
  not csa_tree_add_12_51_groupi_g14879(csa_tree_add_12_51_groupi_n_6883 ,csa_tree_add_12_51_groupi_n_6882);
  nor csa_tree_add_12_51_groupi_g14880__9315(csa_tree_add_12_51_groupi_n_6881 ,csa_tree_add_12_51_groupi_n_6730 ,csa_tree_add_12_51_groupi_n_6830);
  and csa_tree_add_12_51_groupi_g14881__9945(csa_tree_add_12_51_groupi_n_6880 ,csa_tree_add_12_51_groupi_n_6759 ,csa_tree_add_12_51_groupi_n_6834);
  and csa_tree_add_12_51_groupi_g14882__2883(csa_tree_add_12_51_groupi_n_6879 ,csa_tree_add_12_51_groupi_n_6838 ,csa_tree_add_12_51_groupi_n_6822);
  nor csa_tree_add_12_51_groupi_g14883__2346(csa_tree_add_12_51_groupi_n_6878 ,csa_tree_add_12_51_groupi_n_6715 ,csa_tree_add_12_51_groupi_n_6810);
  and csa_tree_add_12_51_groupi_g14884__1666(csa_tree_add_12_51_groupi_n_6877 ,csa_tree_add_12_51_groupi_n_6715 ,csa_tree_add_12_51_groupi_n_6810);
  and csa_tree_add_12_51_groupi_g14885__7410(csa_tree_add_12_51_groupi_n_6876 ,csa_tree_add_12_51_groupi_n_6841 ,csa_tree_add_12_51_groupi_n_6714);
  nor csa_tree_add_12_51_groupi_g14886__6417(csa_tree_add_12_51_groupi_n_6875 ,csa_tree_add_12_51_groupi_n_6841 ,csa_tree_add_12_51_groupi_n_6714);
  nor csa_tree_add_12_51_groupi_g14887__5477(csa_tree_add_12_51_groupi_n_6874 ,csa_tree_add_12_51_groupi_n_6746 ,csa_tree_add_12_51_groupi_n_6845);
  or csa_tree_add_12_51_groupi_g14888__2398(csa_tree_add_12_51_groupi_n_6873 ,csa_tree_add_12_51_groupi_n_6745 ,csa_tree_add_12_51_groupi_n_6844);
  or csa_tree_add_12_51_groupi_g14889__5107(csa_tree_add_12_51_groupi_n_6872 ,csa_tree_add_12_51_groupi_n_6816 ,csa_tree_add_12_51_groupi_n_6719);
  nor csa_tree_add_12_51_groupi_g14890__6260(csa_tree_add_12_51_groupi_n_6871 ,csa_tree_add_12_51_groupi_n_6729 ,csa_tree_add_12_51_groupi_n_6824);
  nor csa_tree_add_12_51_groupi_g14891__4319(csa_tree_add_12_51_groupi_n_6870 ,csa_tree_add_12_51_groupi_n_6789 ,csa_tree_add_12_51_groupi_n_6843);
  or csa_tree_add_12_51_groupi_g14892__8428(csa_tree_add_12_51_groupi_n_6869 ,csa_tree_add_12_51_groupi_n_6788 ,csa_tree_add_12_51_groupi_n_6842);
  nor csa_tree_add_12_51_groupi_g14893__5526(csa_tree_add_12_51_groupi_n_6868 ,csa_tree_add_12_51_groupi_n_6815 ,csa_tree_add_12_51_groupi_n_6720);
  and csa_tree_add_12_51_groupi_g14894__6783(csa_tree_add_12_51_groupi_n_6886 ,csa_tree_add_12_51_groupi_n_6772 ,csa_tree_add_12_51_groupi_n_6835);
  and csa_tree_add_12_51_groupi_g14895__3680(csa_tree_add_12_51_groupi_n_6885 ,csa_tree_add_12_51_groupi_n_6840 ,csa_tree_add_12_51_groupi_n_6776);
  and csa_tree_add_12_51_groupi_g14896__1617(csa_tree_add_12_51_groupi_n_6884 ,csa_tree_add_12_51_groupi_n_6527 ,csa_tree_add_12_51_groupi_n_6837);
  or csa_tree_add_12_51_groupi_g14897__2802(csa_tree_add_12_51_groupi_n_6882 ,csa_tree_add_12_51_groupi_n_6836 ,csa_tree_add_12_51_groupi_n_6739);
  not csa_tree_add_12_51_groupi_g14898(csa_tree_add_12_51_groupi_n_6861 ,csa_tree_add_12_51_groupi_n_6862);
  nor csa_tree_add_12_51_groupi_g14899__1705(csa_tree_add_12_51_groupi_n_6858 ,csa_tree_add_12_51_groupi_n_6809 ,csa_tree_add_12_51_groupi_n_6689);
  or csa_tree_add_12_51_groupi_g14900__5122(csa_tree_add_12_51_groupi_n_6857 ,csa_tree_add_12_51_groupi_n_6808 ,csa_tree_add_12_51_groupi_n_6690);
  or csa_tree_add_12_51_groupi_g14901__8246(csa_tree_add_12_51_groupi_n_6856 ,csa_tree_add_12_51_groupi_n_6828 ,csa_tree_add_12_51_groupi_n_6847);
  nor csa_tree_add_12_51_groupi_g14902__7098(csa_tree_add_12_51_groupi_n_6855 ,csa_tree_add_12_51_groupi_n_6744 ,csa_tree_add_12_51_groupi_n_6813);
  or csa_tree_add_12_51_groupi_g14903__6131(csa_tree_add_12_51_groupi_n_6854 ,csa_tree_add_12_51_groupi_n_6743 ,csa_tree_add_12_51_groupi_n_6814);
  xnor csa_tree_add_12_51_groupi_g14904__1881(out3[12] ,csa_tree_add_12_51_groupi_n_6757 ,csa_tree_add_12_51_groupi_n_6737);
  xnor csa_tree_add_12_51_groupi_g14905__5115(csa_tree_add_12_51_groupi_n_6852 ,csa_tree_add_12_51_groupi_n_6754 ,csa_tree_add_12_51_groupi_n_6716);
  xnor csa_tree_add_12_51_groupi_g14906__7482(csa_tree_add_12_51_groupi_n_6851 ,csa_tree_add_12_51_groupi_n_6692 ,csa_tree_add_12_51_groupi_n_6790);
  xnor csa_tree_add_12_51_groupi_g14907__4733(csa_tree_add_12_51_groupi_n_6850 ,csa_tree_add_12_51_groupi_n_6750 ,csa_tree_add_12_51_groupi_n_6668);
  xnor csa_tree_add_12_51_groupi_g14908__6161(csa_tree_add_12_51_groupi_n_6849 ,csa_tree_add_12_51_groupi_n_6453 ,csa_tree_add_12_51_groupi_n_6783);
  xnor csa_tree_add_12_51_groupi_g14909__9315(csa_tree_add_12_51_groupi_n_6848 ,csa_tree_add_12_51_groupi_n_6752 ,csa_tree_add_12_51_groupi_n_6394);
  xnor csa_tree_add_12_51_groupi_g14910__9945(csa_tree_add_12_51_groupi_n_6867 ,csa_tree_add_12_51_groupi_n_6698 ,csa_tree_add_12_51_groupi_n_6735);
  or csa_tree_add_12_51_groupi_g14911__2883(csa_tree_add_12_51_groupi_n_6866 ,csa_tree_add_12_51_groupi_n_6803 ,csa_tree_add_12_51_groupi_n_6680);
  or csa_tree_add_12_51_groupi_g14912__2346(csa_tree_add_12_51_groupi_n_6865 ,csa_tree_add_12_51_groupi_n_6766 ,csa_tree_add_12_51_groupi_n_6805);
  xnor csa_tree_add_12_51_groupi_g14913__1666(csa_tree_add_12_51_groupi_n_6864 ,csa_tree_add_12_51_groupi_n_6695 ,csa_tree_add_12_51_groupi_n_6736);
  and csa_tree_add_12_51_groupi_g14914__7410(csa_tree_add_12_51_groupi_n_6863 ,csa_tree_add_12_51_groupi_n_6804 ,csa_tree_add_12_51_groupi_n_6742);
  xnor csa_tree_add_12_51_groupi_g14915__6417(csa_tree_add_12_51_groupi_n_6862 ,csa_tree_add_12_51_groupi_n_6552 ,csa_tree_add_12_51_groupi_n_6734);
  xnor csa_tree_add_12_51_groupi_g14916__5477(csa_tree_add_12_51_groupi_n_6860 ,csa_tree_add_12_51_groupi_n_6694 ,csa_tree_add_12_51_groupi_n_6733);
  xnor csa_tree_add_12_51_groupi_g14917__2398(csa_tree_add_12_51_groupi_n_6859 ,csa_tree_add_12_51_groupi_n_6791 ,csa_tree_add_12_51_groupi_n_6603);
  not csa_tree_add_12_51_groupi_g14919(csa_tree_add_12_51_groupi_n_6844 ,csa_tree_add_12_51_groupi_n_6845);
  not csa_tree_add_12_51_groupi_g14920(csa_tree_add_12_51_groupi_n_6842 ,csa_tree_add_12_51_groupi_n_6843);
  or csa_tree_add_12_51_groupi_g14921__5107(csa_tree_add_12_51_groupi_n_6840 ,csa_tree_add_12_51_groupi_n_6777 ,csa_tree_add_12_51_groupi_n_6760);
  and csa_tree_add_12_51_groupi_g14922__6260(csa_tree_add_12_51_groupi_n_6839 ,csa_tree_add_12_51_groupi_n_6754 ,csa_tree_add_12_51_groupi_n_6716);
  or csa_tree_add_12_51_groupi_g14923__4319(csa_tree_add_12_51_groupi_n_6838 ,csa_tree_add_12_51_groupi_n_6754 ,csa_tree_add_12_51_groupi_n_6716);
  or csa_tree_add_12_51_groupi_g14924__8428(csa_tree_add_12_51_groupi_n_6837 ,csa_tree_add_12_51_groupi_n_6526 ,csa_tree_add_12_51_groupi_n_6792);
  and csa_tree_add_12_51_groupi_g14925__5526(csa_tree_add_12_51_groupi_n_6836 ,csa_tree_add_12_51_groupi_n_6758 ,csa_tree_add_12_51_groupi_n_6763);
  or csa_tree_add_12_51_groupi_g14926__6783(csa_tree_add_12_51_groupi_n_6835 ,csa_tree_add_12_51_groupi_n_6771 ,csa_tree_add_12_51_groupi_n_6761);
  or csa_tree_add_12_51_groupi_g14927__3680(csa_tree_add_12_51_groupi_n_6834 ,csa_tree_add_12_51_groupi_n_6752 ,csa_tree_add_12_51_groupi_n_6393);
  and csa_tree_add_12_51_groupi_g14928__1617(csa_tree_add_12_51_groupi_n_6833 ,csa_tree_add_12_51_groupi_n_6750 ,csa_tree_add_12_51_groupi_n_6668);
  or csa_tree_add_12_51_groupi_g14929__2802(csa_tree_add_12_51_groupi_n_6832 ,csa_tree_add_12_51_groupi_n_6750 ,csa_tree_add_12_51_groupi_n_6668);
  and csa_tree_add_12_51_groupi_g14930__1705(csa_tree_add_12_51_groupi_n_6831 ,csa_tree_add_12_51_groupi_n_6688 ,csa_tree_add_12_51_groupi_n_6779);
  nor csa_tree_add_12_51_groupi_g14931__5122(csa_tree_add_12_51_groupi_n_6830 ,csa_tree_add_12_51_groupi_n_6688 ,csa_tree_add_12_51_groupi_n_6779);
  or csa_tree_add_12_51_groupi_g14932__8246(csa_tree_add_12_51_groupi_n_6829 ,csa_tree_add_12_51_groupi_n_6726 ,csa_tree_add_12_51_groupi_n_6755);
  nor csa_tree_add_12_51_groupi_g14933__7098(csa_tree_add_12_51_groupi_n_6828 ,csa_tree_add_12_51_groupi_n_6725 ,csa_tree_add_12_51_groupi_n_6756);
  or csa_tree_add_12_51_groupi_g14934__6131(csa_tree_add_12_51_groupi_n_6827 ,csa_tree_add_12_51_groupi_n_6453 ,csa_tree_add_12_51_groupi_n_6782);
  nor csa_tree_add_12_51_groupi_g14935__1881(csa_tree_add_12_51_groupi_n_6826 ,csa_tree_add_12_51_groupi_n_6452 ,csa_tree_add_12_51_groupi_n_6783);
  nor csa_tree_add_12_51_groupi_g14936__5115(csa_tree_add_12_51_groupi_n_6825 ,csa_tree_add_12_51_groupi_n_6554 ,csa_tree_add_12_51_groupi_n_6753);
  and csa_tree_add_12_51_groupi_g14937__7482(csa_tree_add_12_51_groupi_n_6824 ,csa_tree_add_12_51_groupi_n_6554 ,csa_tree_add_12_51_groupi_n_6753);
  nor csa_tree_add_12_51_groupi_g14938__4733(csa_tree_add_12_51_groupi_n_6823 ,csa_tree_add_12_51_groupi_n_6751 ,csa_tree_add_12_51_groupi_n_6394);
  and csa_tree_add_12_51_groupi_g14939__6161(csa_tree_add_12_51_groupi_n_6847 ,csa_tree_add_12_51_groupi_n_6702 ,csa_tree_add_12_51_groupi_n_6767);
  and csa_tree_add_12_51_groupi_g14940__9315(csa_tree_add_12_51_groupi_n_6846 ,csa_tree_add_12_51_groupi_n_6582 ,csa_tree_add_12_51_groupi_n_6775);
  or csa_tree_add_12_51_groupi_g14941__9945(csa_tree_add_12_51_groupi_n_6845 ,csa_tree_add_12_51_groupi_n_6686 ,csa_tree_add_12_51_groupi_n_6765);
  or csa_tree_add_12_51_groupi_g14942__2883(csa_tree_add_12_51_groupi_n_6843 ,csa_tree_add_12_51_groupi_n_6700 ,csa_tree_add_12_51_groupi_n_6768);
  and csa_tree_add_12_51_groupi_g14943__2346(csa_tree_add_12_51_groupi_n_6841 ,csa_tree_add_12_51_groupi_n_6576 ,csa_tree_add_12_51_groupi_n_6774);
  not csa_tree_add_12_51_groupi_g14944(csa_tree_add_12_51_groupi_n_6819 ,csa_tree_add_12_51_groupi_n_6820);
  not csa_tree_add_12_51_groupi_g14945(csa_tree_add_12_51_groupi_n_6817 ,csa_tree_add_12_51_groupi_n_6818);
  not csa_tree_add_12_51_groupi_g14946(csa_tree_add_12_51_groupi_n_6815 ,csa_tree_add_12_51_groupi_n_6816);
  not csa_tree_add_12_51_groupi_g14947(csa_tree_add_12_51_groupi_n_6813 ,csa_tree_add_12_51_groupi_n_6814);
  not csa_tree_add_12_51_groupi_g14948(csa_tree_add_12_51_groupi_n_6812 ,csa_tree_add_12_51_groupi_n_6811);
  not csa_tree_add_12_51_groupi_g14949(csa_tree_add_12_51_groupi_n_6808 ,csa_tree_add_12_51_groupi_n_6809);
  not csa_tree_add_12_51_groupi_g14950(csa_tree_add_12_51_groupi_n_6806 ,csa_tree_add_12_51_groupi_n_6807);
  and csa_tree_add_12_51_groupi_g14951__1666(csa_tree_add_12_51_groupi_n_6805 ,csa_tree_add_12_51_groupi_n_6769 ,csa_tree_add_12_51_groupi_n_6790);
  or csa_tree_add_12_51_groupi_g14952__7410(csa_tree_add_12_51_groupi_n_6804 ,csa_tree_add_12_51_groupi_n_6762 ,csa_tree_add_12_51_groupi_n_6741);
  and csa_tree_add_12_51_groupi_g14953__6417(csa_tree_add_12_51_groupi_n_6803 ,csa_tree_add_12_51_groupi_n_6678 ,csa_tree_add_12_51_groupi_n_6757);
  xnor csa_tree_add_12_51_groupi_g14954__5477(csa_tree_add_12_51_groupi_n_6802 ,csa_tree_add_12_51_groupi_n_6631 ,csa_tree_add_12_51_groupi_n_6696);
  xnor csa_tree_add_12_51_groupi_g14955__2398(csa_tree_add_12_51_groupi_n_6801 ,csa_tree_add_12_51_groupi_n_6633 ,csa_tree_add_12_51_groupi_n_6697);
  xnor csa_tree_add_12_51_groupi_g14957__5107(csa_tree_add_12_51_groupi_n_6800 ,csa_tree_add_12_51_groupi_n_6539 ,csa_tree_add_12_51_groupi_n_6727);
  xnor csa_tree_add_12_51_groupi_g14958__6260(csa_tree_add_12_51_groupi_n_6799 ,csa_tree_add_12_51_groupi_n_6548 ,csa_tree_add_12_51_groupi_n_6718);
  xnor csa_tree_add_12_51_groupi_g14959__4319(csa_tree_add_12_51_groupi_n_6798 ,csa_tree_add_12_51_groupi_n_6730 ,csa_tree_add_12_51_groupi_n_6688);
  xnor csa_tree_add_12_51_groupi_g14960__8428(csa_tree_add_12_51_groupi_n_6797 ,csa_tree_add_12_51_groupi_n_5022 ,csa_tree_add_12_51_groupi_n_6724);
  xnor csa_tree_add_12_51_groupi_g14961__5526(csa_tree_add_12_51_groupi_n_6796 ,csa_tree_add_12_51_groupi_n_6556 ,csa_tree_add_12_51_groupi_n_6712);
  xnor csa_tree_add_12_51_groupi_g14962__6783(csa_tree_add_12_51_groupi_n_6795 ,csa_tree_add_12_51_groupi_n_6536 ,csa_tree_add_12_51_groupi_n_6722);
  xnor csa_tree_add_12_51_groupi_g14963__3680(csa_tree_add_12_51_groupi_n_6794 ,csa_tree_add_12_51_groupi_n_6538 ,csa_tree_add_12_51_groupi_n_6728);
  xnor csa_tree_add_12_51_groupi_g14964__1617(csa_tree_add_12_51_groupi_n_6793 ,csa_tree_add_12_51_groupi_n_6729 ,csa_tree_add_12_51_groupi_n_6554);
  xnor csa_tree_add_12_51_groupi_g14965__2802(csa_tree_add_12_51_groupi_n_6822 ,csa_tree_add_12_51_groupi_n_6636 ,csa_tree_add_12_51_groupi_n_6675);
  and csa_tree_add_12_51_groupi_g14966__1705(csa_tree_add_12_51_groupi_n_6821 ,csa_tree_add_12_51_groupi_n_6687 ,csa_tree_add_12_51_groupi_n_6773);
  xnor csa_tree_add_12_51_groupi_g14967__5122(csa_tree_add_12_51_groupi_n_6820 ,csa_tree_add_12_51_groupi_n_5056 ,csa_tree_add_12_51_groupi_n_6670);
  xnor csa_tree_add_12_51_groupi_g14968__8246(csa_tree_add_12_51_groupi_n_6818 ,csa_tree_add_12_51_groupi_n_6600 ,csa_tree_add_12_51_groupi_n_6672);
  xnor csa_tree_add_12_51_groupi_g14969__7098(csa_tree_add_12_51_groupi_n_6816 ,csa_tree_add_12_51_groupi_n_6546 ,csa_tree_add_12_51_groupi_n_6673);
  and csa_tree_add_12_51_groupi_g14970__6131(csa_tree_add_12_51_groupi_n_6814 ,csa_tree_add_12_51_groupi_n_6682 ,csa_tree_add_12_51_groupi_n_6770);
  xnor csa_tree_add_12_51_groupi_g14971__1881(csa_tree_add_12_51_groupi_n_6811 ,csa_tree_add_12_51_groupi_n_6731 ,csa_tree_add_12_51_groupi_n_6610);
  xnor csa_tree_add_12_51_groupi_g14972__5115(csa_tree_add_12_51_groupi_n_6810 ,csa_tree_add_12_51_groupi_n_6550 ,csa_tree_add_12_51_groupi_n_6671);
  xnor csa_tree_add_12_51_groupi_g14973__7482(csa_tree_add_12_51_groupi_n_6809 ,csa_tree_add_12_51_groupi_n_6559 ,csa_tree_add_12_51_groupi_n_6674);
  or csa_tree_add_12_51_groupi_g14974__4733(csa_tree_add_12_51_groupi_n_6807 ,csa_tree_add_12_51_groupi_n_6677 ,csa_tree_add_12_51_groupi_n_6740);
  not csa_tree_add_12_51_groupi_g14975(csa_tree_add_12_51_groupi_n_6792 ,csa_tree_add_12_51_groupi_n_6791);
  not csa_tree_add_12_51_groupi_g14976(csa_tree_add_12_51_groupi_n_6789 ,csa_tree_add_12_51_groupi_n_6788);
  not csa_tree_add_12_51_groupi_g14977(csa_tree_add_12_51_groupi_n_6785 ,csa_tree_add_12_51_groupi_n_6786);
  not csa_tree_add_12_51_groupi_g14978(csa_tree_add_12_51_groupi_n_6782 ,csa_tree_add_12_51_groupi_n_6783);
  not csa_tree_add_12_51_groupi_g14979(csa_tree_add_12_51_groupi_n_6780 ,csa_tree_add_12_51_groupi_n_6781);
  or csa_tree_add_12_51_groupi_g14980__6161(csa_tree_add_12_51_groupi_n_6778 ,csa_tree_add_12_51_groupi_n_6723 ,csa_tree_add_12_51_groupi_n_5021);
  nor csa_tree_add_12_51_groupi_g14981__9315(csa_tree_add_12_51_groupi_n_6777 ,csa_tree_add_12_51_groupi_n_6556 ,csa_tree_add_12_51_groupi_n_6712);
  or csa_tree_add_12_51_groupi_g14982__9945(csa_tree_add_12_51_groupi_n_6776 ,csa_tree_add_12_51_groupi_n_6555 ,csa_tree_add_12_51_groupi_n_6711);
  or csa_tree_add_12_51_groupi_g14983__2883(csa_tree_add_12_51_groupi_n_6775 ,csa_tree_add_12_51_groupi_n_6581 ,csa_tree_add_12_51_groupi_n_6732);
  or csa_tree_add_12_51_groupi_g14984__2346(csa_tree_add_12_51_groupi_n_6774 ,csa_tree_add_12_51_groupi_n_6573 ,csa_tree_add_12_51_groupi_n_6693);
  or csa_tree_add_12_51_groupi_g14985__1666(csa_tree_add_12_51_groupi_n_6773 ,csa_tree_add_12_51_groupi_n_6684 ,csa_tree_add_12_51_groupi_n_6696);
  or csa_tree_add_12_51_groupi_g14986__7410(csa_tree_add_12_51_groupi_n_6772 ,csa_tree_add_12_51_groupi_n_6535 ,csa_tree_add_12_51_groupi_n_6721);
  nor csa_tree_add_12_51_groupi_g14987__6417(csa_tree_add_12_51_groupi_n_6771 ,csa_tree_add_12_51_groupi_n_6536 ,csa_tree_add_12_51_groupi_n_6722);
  or csa_tree_add_12_51_groupi_g14988__5477(csa_tree_add_12_51_groupi_n_6770 ,csa_tree_add_12_51_groupi_n_6681 ,csa_tree_add_12_51_groupi_n_6697);
  or csa_tree_add_12_51_groupi_g14989__2398(csa_tree_add_12_51_groupi_n_6769 ,csa_tree_add_12_51_groupi_n_5023 ,csa_tree_add_12_51_groupi_n_6692);
  and csa_tree_add_12_51_groupi_g14990__5107(csa_tree_add_12_51_groupi_n_6768 ,csa_tree_add_12_51_groupi_n_6728 ,csa_tree_add_12_51_groupi_n_6699);
  or csa_tree_add_12_51_groupi_g14991__6260(csa_tree_add_12_51_groupi_n_6767 ,csa_tree_add_12_51_groupi_n_6698 ,csa_tree_add_12_51_groupi_n_6707);
  nor csa_tree_add_12_51_groupi_g14992__4319(csa_tree_add_12_51_groupi_n_6766 ,csa_tree_add_12_51_groupi_n_5024 ,csa_tree_add_12_51_groupi_n_6691);
  and csa_tree_add_12_51_groupi_g14993__8428(csa_tree_add_12_51_groupi_n_6765 ,csa_tree_add_12_51_groupi_n_6695 ,csa_tree_add_12_51_groupi_n_6685);
  nor csa_tree_add_12_51_groupi_g14994__5526(csa_tree_add_12_51_groupi_n_6764 ,csa_tree_add_12_51_groupi_n_6724 ,csa_tree_add_12_51_groupi_n_5022);
  or csa_tree_add_12_51_groupi_g14995__6783(csa_tree_add_12_51_groupi_n_6763 ,csa_tree_add_12_51_groupi_n_6540 ,csa_tree_add_12_51_groupi_n_6727);
  or csa_tree_add_12_51_groupi_g14996__3680(csa_tree_add_12_51_groupi_n_6791 ,csa_tree_add_12_51_groupi_n_6622 ,csa_tree_add_12_51_groupi_n_6683);
  or csa_tree_add_12_51_groupi_g14997__1617(csa_tree_add_12_51_groupi_n_6790 ,csa_tree_add_12_51_groupi_n_6648 ,csa_tree_add_12_51_groupi_n_6703);
  and csa_tree_add_12_51_groupi_g14998__2802(csa_tree_add_12_51_groupi_n_6788 ,csa_tree_add_12_51_groupi_n_6651 ,csa_tree_add_12_51_groupi_n_6708);
  or csa_tree_add_12_51_groupi_g14999__1705(csa_tree_add_12_51_groupi_n_6787 ,csa_tree_add_12_51_groupi_n_6642 ,csa_tree_add_12_51_groupi_n_6706);
  or csa_tree_add_12_51_groupi_g15000__5122(csa_tree_add_12_51_groupi_n_6786 ,csa_tree_add_12_51_groupi_n_6705 ,csa_tree_add_12_51_groupi_n_6645);
  or csa_tree_add_12_51_groupi_g15001__8246(csa_tree_add_12_51_groupi_n_6784 ,csa_tree_add_12_51_groupi_n_6649 ,csa_tree_add_12_51_groupi_n_6709);
  or csa_tree_add_12_51_groupi_g15002__7098(csa_tree_add_12_51_groupi_n_6783 ,csa_tree_add_12_51_groupi_n_6667 ,csa_tree_add_12_51_groupi_n_6701);
  or csa_tree_add_12_51_groupi_g15003__6131(csa_tree_add_12_51_groupi_n_6781 ,csa_tree_add_12_51_groupi_n_6656 ,csa_tree_add_12_51_groupi_n_6704);
  or csa_tree_add_12_51_groupi_g15004__1881(csa_tree_add_12_51_groupi_n_6779 ,csa_tree_add_12_51_groupi_n_6639 ,csa_tree_add_12_51_groupi_n_6710);
  not csa_tree_add_12_51_groupi_g15005(csa_tree_add_12_51_groupi_n_6755 ,csa_tree_add_12_51_groupi_n_6756);
  not csa_tree_add_12_51_groupi_g15006(csa_tree_add_12_51_groupi_n_6751 ,csa_tree_add_12_51_groupi_n_6752);
  not csa_tree_add_12_51_groupi_g15008(csa_tree_add_12_51_groupi_n_6747 ,csa_tree_add_12_51_groupi_n_6748);
  not csa_tree_add_12_51_groupi_g15009(csa_tree_add_12_51_groupi_n_6745 ,csa_tree_add_12_51_groupi_n_6746);
  not csa_tree_add_12_51_groupi_g15010(csa_tree_add_12_51_groupi_n_6744 ,csa_tree_add_12_51_groupi_n_6743);
  or csa_tree_add_12_51_groupi_g15011__5115(csa_tree_add_12_51_groupi_n_6742 ,csa_tree_add_12_51_groupi_n_6547 ,csa_tree_add_12_51_groupi_n_6717);
  nor csa_tree_add_12_51_groupi_g15012__7482(csa_tree_add_12_51_groupi_n_6741 ,csa_tree_add_12_51_groupi_n_6548 ,csa_tree_add_12_51_groupi_n_6718);
  and csa_tree_add_12_51_groupi_g15013__4733(csa_tree_add_12_51_groupi_n_6740 ,csa_tree_add_12_51_groupi_n_6694 ,csa_tree_add_12_51_groupi_n_6676);
  and csa_tree_add_12_51_groupi_g15014__6161(csa_tree_add_12_51_groupi_n_6739 ,csa_tree_add_12_51_groupi_n_6540 ,csa_tree_add_12_51_groupi_n_6727);
  xnor csa_tree_add_12_51_groupi_g15015__9315(out3[11] ,csa_tree_add_12_51_groupi_n_6637 ,csa_tree_add_12_51_groupi_n_6606);
  xnor csa_tree_add_12_51_groupi_g15016__9945(csa_tree_add_12_51_groupi_n_6737 ,csa_tree_add_12_51_groupi_n_6423 ,csa_tree_add_12_51_groupi_n_6635);
  xnor csa_tree_add_12_51_groupi_g15017__2883(csa_tree_add_12_51_groupi_n_6736 ,csa_tree_add_12_51_groupi_n_6627 ,csa_tree_add_12_51_groupi_n_6534);
  xnor csa_tree_add_12_51_groupi_g15018__2346(csa_tree_add_12_51_groupi_n_6735 ,csa_tree_add_12_51_groupi_n_6629 ,csa_tree_add_12_51_groupi_n_6594);
  xnor csa_tree_add_12_51_groupi_g15019__1666(csa_tree_add_12_51_groupi_n_6734 ,csa_tree_add_12_51_groupi_n_6557 ,csa_tree_add_12_51_groupi_n_6669);
  xnor csa_tree_add_12_51_groupi_g15020__7410(csa_tree_add_12_51_groupi_n_6733 ,csa_tree_add_12_51_groupi_n_6541 ,csa_tree_add_12_51_groupi_n_6625);
  xnor csa_tree_add_12_51_groupi_g15021__6417(csa_tree_add_12_51_groupi_n_6762 ,csa_tree_add_12_51_groupi_n_6599 ,csa_tree_add_12_51_groupi_n_6612);
  xnor csa_tree_add_12_51_groupi_g15022__5477(csa_tree_add_12_51_groupi_n_6761 ,csa_tree_add_12_51_groupi_n_6466 ,csa_tree_add_12_51_groupi_n_6602);
  xnor csa_tree_add_12_51_groupi_g15023__2398(csa_tree_add_12_51_groupi_n_6760 ,csa_tree_add_12_51_groupi_n_6467 ,csa_tree_add_12_51_groupi_n_6614);
  xnor csa_tree_add_12_51_groupi_g15024__5107(csa_tree_add_12_51_groupi_n_6759 ,csa_tree_add_12_51_groupi_n_6598 ,csa_tree_add_12_51_groupi_n_6604);
  xnor csa_tree_add_12_51_groupi_g15025__6260(csa_tree_add_12_51_groupi_n_6758 ,csa_tree_add_12_51_groupi_n_6601 ,csa_tree_add_12_51_groupi_n_6613);
  or csa_tree_add_12_51_groupi_g15026__4319(csa_tree_add_12_51_groupi_n_6757 ,csa_tree_add_12_51_groupi_n_6679 ,csa_tree_add_12_51_groupi_n_6528);
  xnor csa_tree_add_12_51_groupi_g15027__8428(csa_tree_add_12_51_groupi_n_6756 ,csa_tree_add_12_51_groupi_n_6514 ,csa_tree_add_12_51_groupi_n_6608);
  xnor csa_tree_add_12_51_groupi_g15028__5526(csa_tree_add_12_51_groupi_n_6754 ,csa_tree_add_12_51_groupi_n_6511 ,csa_tree_add_12_51_groupi_n_6616);
  xnor csa_tree_add_12_51_groupi_g15029__6783(csa_tree_add_12_51_groupi_n_6753 ,csa_tree_add_12_51_groupi_n_6542 ,csa_tree_add_12_51_groupi_n_6607);
  xnor csa_tree_add_12_51_groupi_g15030__3680(csa_tree_add_12_51_groupi_n_6752 ,csa_tree_add_12_51_groupi_n_6510 ,csa_tree_add_12_51_groupi_n_6618);
  xnor csa_tree_add_12_51_groupi_g15031__1617(csa_tree_add_12_51_groupi_n_6750 ,csa_tree_add_12_51_groupi_n_6549 ,csa_tree_add_12_51_groupi_n_6617);
  xnor csa_tree_add_12_51_groupi_g15032__2802(csa_tree_add_12_51_groupi_n_6749 ,csa_tree_add_12_51_groupi_n_6470 ,csa_tree_add_12_51_groupi_n_6605);
  xnor csa_tree_add_12_51_groupi_g15033__1705(csa_tree_add_12_51_groupi_n_6748 ,csa_tree_add_12_51_groupi_n_6471 ,csa_tree_add_12_51_groupi_n_6611);
  xnor csa_tree_add_12_51_groupi_g15034__5122(csa_tree_add_12_51_groupi_n_6746 ,csa_tree_add_12_51_groupi_n_6516 ,csa_tree_add_12_51_groupi_n_6615);
  xnor csa_tree_add_12_51_groupi_g15035__8246(csa_tree_add_12_51_groupi_n_6743 ,csa_tree_add_12_51_groupi_n_6500 ,csa_tree_add_12_51_groupi_n_6609);
  not csa_tree_add_12_51_groupi_g15036(csa_tree_add_12_51_groupi_n_6732 ,csa_tree_add_12_51_groupi_n_6731);
  not csa_tree_add_12_51_groupi_g15037(csa_tree_add_12_51_groupi_n_6725 ,csa_tree_add_12_51_groupi_n_6726);
  not csa_tree_add_12_51_groupi_g15038(csa_tree_add_12_51_groupi_n_6723 ,csa_tree_add_12_51_groupi_n_6724);
  not csa_tree_add_12_51_groupi_g15039(csa_tree_add_12_51_groupi_n_6721 ,csa_tree_add_12_51_groupi_n_6722);
  not csa_tree_add_12_51_groupi_g15040(csa_tree_add_12_51_groupi_n_6719 ,csa_tree_add_12_51_groupi_n_6720);
  not csa_tree_add_12_51_groupi_g15041(csa_tree_add_12_51_groupi_n_6717 ,csa_tree_add_12_51_groupi_n_6718);
  not csa_tree_add_12_51_groupi_g15042(csa_tree_add_12_51_groupi_n_6714 ,csa_tree_add_12_51_groupi_n_6713);
  not csa_tree_add_12_51_groupi_g15043(csa_tree_add_12_51_groupi_n_6711 ,csa_tree_add_12_51_groupi_n_6712);
  and csa_tree_add_12_51_groupi_g15044__7098(csa_tree_add_12_51_groupi_n_6710 ,csa_tree_add_12_51_groupi_n_6638 ,csa_tree_add_12_51_groupi_n_6600);
  nor csa_tree_add_12_51_groupi_g15045__6131(csa_tree_add_12_51_groupi_n_6709 ,csa_tree_add_12_51_groupi_n_6558 ,csa_tree_add_12_51_groupi_n_6665);
  or csa_tree_add_12_51_groupi_g15046__1881(csa_tree_add_12_51_groupi_n_6708 ,csa_tree_add_12_51_groupi_n_6664 ,csa_tree_add_12_51_groupi_n_6472);
  nor csa_tree_add_12_51_groupi_g15047__5115(csa_tree_add_12_51_groupi_n_6707 ,csa_tree_add_12_51_groupi_n_6629 ,csa_tree_add_12_51_groupi_n_6594);
  nor csa_tree_add_12_51_groupi_g15048__7482(csa_tree_add_12_51_groupi_n_6706 ,csa_tree_add_12_51_groupi_n_6429 ,csa_tree_add_12_51_groupi_n_6641);
  and csa_tree_add_12_51_groupi_g15049__4733(csa_tree_add_12_51_groupi_n_6705 ,csa_tree_add_12_51_groupi_n_6636 ,csa_tree_add_12_51_groupi_n_6646);
  and csa_tree_add_12_51_groupi_g15050__6161(csa_tree_add_12_51_groupi_n_6704 ,csa_tree_add_12_51_groupi_n_6559 ,csa_tree_add_12_51_groupi_n_6655);
  nor csa_tree_add_12_51_groupi_g15051__9315(csa_tree_add_12_51_groupi_n_6703 ,csa_tree_add_12_51_groupi_n_6562 ,csa_tree_add_12_51_groupi_n_6647);
  or csa_tree_add_12_51_groupi_g15052__9945(csa_tree_add_12_51_groupi_n_6702 ,csa_tree_add_12_51_groupi_n_6628 ,csa_tree_add_12_51_groupi_n_6593);
  and csa_tree_add_12_51_groupi_g15053__2883(csa_tree_add_12_51_groupi_n_6701 ,csa_tree_add_12_51_groupi_n_6650 ,csa_tree_add_12_51_groupi_n_6669);
  and csa_tree_add_12_51_groupi_g15054__2346(csa_tree_add_12_51_groupi_n_6700 ,csa_tree_add_12_51_groupi_n_6538 ,csa_tree_add_12_51_groupi_n_6634);
  or csa_tree_add_12_51_groupi_g15055__1666(csa_tree_add_12_51_groupi_n_6699 ,csa_tree_add_12_51_groupi_n_6538 ,csa_tree_add_12_51_groupi_n_6634);
  or csa_tree_add_12_51_groupi_g15056__7410(csa_tree_add_12_51_groupi_n_6731 ,csa_tree_add_12_51_groupi_n_6661 ,csa_tree_add_12_51_groupi_n_6575);
  and csa_tree_add_12_51_groupi_g15057__6417(csa_tree_add_12_51_groupi_n_6730 ,csa_tree_add_12_51_groupi_n_6574 ,csa_tree_add_12_51_groupi_n_6658);
  and csa_tree_add_12_51_groupi_g15058__5477(csa_tree_add_12_51_groupi_n_6729 ,csa_tree_add_12_51_groupi_n_6591 ,csa_tree_add_12_51_groupi_n_6666);
  or csa_tree_add_12_51_groupi_g15059__2398(csa_tree_add_12_51_groupi_n_6728 ,csa_tree_add_12_51_groupi_n_6588 ,csa_tree_add_12_51_groupi_n_6663);
  or csa_tree_add_12_51_groupi_g15060__5107(csa_tree_add_12_51_groupi_n_6727 ,csa_tree_add_12_51_groupi_n_6483 ,csa_tree_add_12_51_groupi_n_6657);
  and csa_tree_add_12_51_groupi_g15061__6260(csa_tree_add_12_51_groupi_n_6726 ,csa_tree_add_12_51_groupi_n_6571 ,csa_tree_add_12_51_groupi_n_6653);
  and csa_tree_add_12_51_groupi_g15062__4319(csa_tree_add_12_51_groupi_n_6724 ,csa_tree_add_12_51_groupi_n_6568 ,csa_tree_add_12_51_groupi_n_6660);
  or csa_tree_add_12_51_groupi_g15063__8428(csa_tree_add_12_51_groupi_n_6722 ,csa_tree_add_12_51_groupi_n_6570 ,csa_tree_add_12_51_groupi_n_6654);
  or csa_tree_add_12_51_groupi_g15064__5526(csa_tree_add_12_51_groupi_n_6720 ,csa_tree_add_12_51_groupi_n_6578 ,csa_tree_add_12_51_groupi_n_6659);
  or csa_tree_add_12_51_groupi_g15065__6783(csa_tree_add_12_51_groupi_n_6718 ,csa_tree_add_12_51_groupi_n_6564 ,csa_tree_add_12_51_groupi_n_6644);
  or csa_tree_add_12_51_groupi_g15066__3680(csa_tree_add_12_51_groupi_n_6716 ,csa_tree_add_12_51_groupi_n_6566 ,csa_tree_add_12_51_groupi_n_6643);
  or csa_tree_add_12_51_groupi_g15067__1617(csa_tree_add_12_51_groupi_n_6715 ,csa_tree_add_12_51_groupi_n_6586 ,csa_tree_add_12_51_groupi_n_6662);
  or csa_tree_add_12_51_groupi_g15068__2802(csa_tree_add_12_51_groupi_n_6713 ,csa_tree_add_12_51_groupi_n_6525 ,csa_tree_add_12_51_groupi_n_6652);
  or csa_tree_add_12_51_groupi_g15069__1705(csa_tree_add_12_51_groupi_n_6712 ,csa_tree_add_12_51_groupi_n_6592 ,csa_tree_add_12_51_groupi_n_6640);
  not csa_tree_add_12_51_groupi_g15071(csa_tree_add_12_51_groupi_n_6691 ,csa_tree_add_12_51_groupi_n_6692);
  not csa_tree_add_12_51_groupi_g15072(csa_tree_add_12_51_groupi_n_6690 ,csa_tree_add_12_51_groupi_n_6689);
  or csa_tree_add_12_51_groupi_g15073__5122(csa_tree_add_12_51_groupi_n_6687 ,csa_tree_add_12_51_groupi_n_6465 ,csa_tree_add_12_51_groupi_n_6630);
  nor csa_tree_add_12_51_groupi_g15074__8246(csa_tree_add_12_51_groupi_n_6686 ,csa_tree_add_12_51_groupi_n_6627 ,csa_tree_add_12_51_groupi_n_6533);
  or csa_tree_add_12_51_groupi_g15075__7098(csa_tree_add_12_51_groupi_n_6685 ,csa_tree_add_12_51_groupi_n_6626 ,csa_tree_add_12_51_groupi_n_6534);
  nor csa_tree_add_12_51_groupi_g15076__6131(csa_tree_add_12_51_groupi_n_6684 ,csa_tree_add_12_51_groupi_n_6464 ,csa_tree_add_12_51_groupi_n_6631);
  nor csa_tree_add_12_51_groupi_g15077__1881(csa_tree_add_12_51_groupi_n_6683 ,csa_tree_add_12_51_groupi_n_6621 ,csa_tree_add_12_51_groupi_n_6400);
  or csa_tree_add_12_51_groupi_g15078__5115(csa_tree_add_12_51_groupi_n_6682 ,csa_tree_add_12_51_groupi_n_6463 ,csa_tree_add_12_51_groupi_n_6632);
  nor csa_tree_add_12_51_groupi_g15079__7482(csa_tree_add_12_51_groupi_n_6681 ,csa_tree_add_12_51_groupi_n_6462 ,csa_tree_add_12_51_groupi_n_6633);
  and csa_tree_add_12_51_groupi_g15080__4733(csa_tree_add_12_51_groupi_n_6680 ,csa_tree_add_12_51_groupi_n_6423 ,csa_tree_add_12_51_groupi_n_6635);
  and csa_tree_add_12_51_groupi_g15081__6161(csa_tree_add_12_51_groupi_n_6679 ,csa_tree_add_12_51_groupi_n_6522 ,csa_tree_add_12_51_groupi_n_6637);
  or csa_tree_add_12_51_groupi_g15082__9315(csa_tree_add_12_51_groupi_n_6678 ,csa_tree_add_12_51_groupi_n_6423 ,csa_tree_add_12_51_groupi_n_6635);
  and csa_tree_add_12_51_groupi_g15083__9945(csa_tree_add_12_51_groupi_n_6677 ,csa_tree_add_12_51_groupi_n_6541 ,csa_tree_add_12_51_groupi_n_6625);
  or csa_tree_add_12_51_groupi_g15084__2883(csa_tree_add_12_51_groupi_n_6676 ,csa_tree_add_12_51_groupi_n_6541 ,csa_tree_add_12_51_groupi_n_6625);
  xnor csa_tree_add_12_51_groupi_g15085__2346(csa_tree_add_12_51_groupi_n_6675 ,csa_tree_add_12_51_groupi_n_6504 ,csa_tree_add_12_51_groupi_n_6597);
  xnor csa_tree_add_12_51_groupi_g15086__1666(csa_tree_add_12_51_groupi_n_6674 ,csa_tree_add_12_51_groupi_n_6537 ,csa_tree_add_12_51_groupi_n_6509);
  xnor csa_tree_add_12_51_groupi_g15087__7410(csa_tree_add_12_51_groupi_n_6673 ,csa_tree_add_12_51_groupi_n_6544 ,csa_tree_add_12_51_groupi_n_6472);
  xnor csa_tree_add_12_51_groupi_g15088__6417(csa_tree_add_12_51_groupi_n_6672 ,csa_tree_add_12_51_groupi_n_6596 ,csa_tree_add_12_51_groupi_n_5177);
  xnor csa_tree_add_12_51_groupi_g15089__5477(csa_tree_add_12_51_groupi_n_6671 ,csa_tree_add_12_51_groupi_n_6495 ,csa_tree_add_12_51_groupi_n_6558);
  xnor csa_tree_add_12_51_groupi_g15090__2398(csa_tree_add_12_51_groupi_n_6670 ,csa_tree_add_12_51_groupi_n_6562 ,csa_tree_add_12_51_groupi_n_6553);
  xnor csa_tree_add_12_51_groupi_g15091__5107(csa_tree_add_12_51_groupi_n_6698 ,csa_tree_add_12_51_groupi_n_5028 ,csa_tree_add_12_51_groupi_n_6517);
  xnor csa_tree_add_12_51_groupi_g15092__6260(csa_tree_add_12_51_groupi_n_6697 ,csa_tree_add_12_51_groupi_n_6561 ,csa_tree_add_12_51_groupi_n_6521);
  xnor csa_tree_add_12_51_groupi_g15093__4319(csa_tree_add_12_51_groupi_n_6696 ,csa_tree_add_12_51_groupi_n_6444 ,csa_tree_add_12_51_groupi_n_6519);
  xnor csa_tree_add_12_51_groupi_g15094__8428(csa_tree_add_12_51_groupi_n_6695 ,csa_tree_add_12_51_groupi_n_6448 ,csa_tree_add_12_51_groupi_n_6520);
  xnor csa_tree_add_12_51_groupi_g15095__5526(csa_tree_add_12_51_groupi_n_6694 ,csa_tree_add_12_51_groupi_n_6445 ,csa_tree_add_12_51_groupi_n_6518);
  and csa_tree_add_12_51_groupi_g15096__6783(csa_tree_add_12_51_groupi_n_6693 ,csa_tree_add_12_51_groupi_n_6623 ,csa_tree_add_12_51_groupi_n_6585);
  or csa_tree_add_12_51_groupi_g15097__3680(csa_tree_add_12_51_groupi_n_6692 ,csa_tree_add_12_51_groupi_n_4802 ,csa_tree_add_12_51_groupi_n_6624);
  or csa_tree_add_12_51_groupi_g15098__1617(csa_tree_add_12_51_groupi_n_6689 ,csa_tree_add_12_51_groupi_n_6530 ,csa_tree_add_12_51_groupi_n_6619);
  xnor csa_tree_add_12_51_groupi_g15099__2802(csa_tree_add_12_51_groupi_n_6688 ,csa_tree_add_12_51_groupi_n_6560 ,csa_tree_add_12_51_groupi_n_4824);
  and csa_tree_add_12_51_groupi_g15100__1705(csa_tree_add_12_51_groupi_n_6667 ,csa_tree_add_12_51_groupi_n_6552 ,csa_tree_add_12_51_groupi_n_6557);
  or csa_tree_add_12_51_groupi_g15101__5122(csa_tree_add_12_51_groupi_n_6666 ,csa_tree_add_12_51_groupi_n_6512 ,csa_tree_add_12_51_groupi_n_6590);
  and csa_tree_add_12_51_groupi_g15102__8246(csa_tree_add_12_51_groupi_n_6665 ,csa_tree_add_12_51_groupi_n_6551 ,csa_tree_add_12_51_groupi_n_6495);
  nor csa_tree_add_12_51_groupi_g15103__7098(csa_tree_add_12_51_groupi_n_6664 ,csa_tree_add_12_51_groupi_n_6546 ,csa_tree_add_12_51_groupi_n_6544);
  and csa_tree_add_12_51_groupi_g15104__6131(csa_tree_add_12_51_groupi_n_6663 ,csa_tree_add_12_51_groupi_n_6510 ,csa_tree_add_12_51_groupi_n_6587);
  and csa_tree_add_12_51_groupi_g15105__1881(csa_tree_add_12_51_groupi_n_6662 ,csa_tree_add_12_51_groupi_n_6584 ,csa_tree_add_12_51_groupi_n_6601);
  nor csa_tree_add_12_51_groupi_g15106__5115(csa_tree_add_12_51_groupi_n_6661 ,csa_tree_add_12_51_groupi_n_6580 ,csa_tree_add_12_51_groupi_n_6466);
  or csa_tree_add_12_51_groupi_g15107__7482(csa_tree_add_12_51_groupi_n_6660 ,csa_tree_add_12_51_groupi_n_6471 ,csa_tree_add_12_51_groupi_n_6579);
  and csa_tree_add_12_51_groupi_g15108__4733(csa_tree_add_12_51_groupi_n_6659 ,csa_tree_add_12_51_groupi_n_6598 ,csa_tree_add_12_51_groupi_n_6577);
  or csa_tree_add_12_51_groupi_g15109__6161(csa_tree_add_12_51_groupi_n_6658 ,csa_tree_add_12_51_groupi_n_6515 ,csa_tree_add_12_51_groupi_n_6572);
  nor csa_tree_add_12_51_groupi_g15110__9315(csa_tree_add_12_51_groupi_n_6657 ,csa_tree_add_12_51_groupi_n_6482 ,csa_tree_add_12_51_groupi_n_6561);
  and csa_tree_add_12_51_groupi_g15111__9945(csa_tree_add_12_51_groupi_n_6656 ,csa_tree_add_12_51_groupi_n_6537 ,csa_tree_add_12_51_groupi_n_6509);
  or csa_tree_add_12_51_groupi_g15112__2883(csa_tree_add_12_51_groupi_n_6655 ,csa_tree_add_12_51_groupi_n_6537 ,csa_tree_add_12_51_groupi_n_6509);
  and csa_tree_add_12_51_groupi_g15113__2346(csa_tree_add_12_51_groupi_n_6654 ,csa_tree_add_12_51_groupi_n_6516 ,csa_tree_add_12_51_groupi_n_6569);
  or csa_tree_add_12_51_groupi_g15114__1666(csa_tree_add_12_51_groupi_n_6653 ,csa_tree_add_12_51_groupi_n_6470 ,csa_tree_add_12_51_groupi_n_6567);
  and csa_tree_add_12_51_groupi_g15115__7410(csa_tree_add_12_51_groupi_n_6652 ,csa_tree_add_12_51_groupi_n_6524 ,csa_tree_add_12_51_groupi_n_6428);
  or csa_tree_add_12_51_groupi_g15116__6417(csa_tree_add_12_51_groupi_n_6651 ,csa_tree_add_12_51_groupi_n_6545 ,csa_tree_add_12_51_groupi_n_6543);
  or csa_tree_add_12_51_groupi_g15117__5477(csa_tree_add_12_51_groupi_n_6650 ,csa_tree_add_12_51_groupi_n_6552 ,csa_tree_add_12_51_groupi_n_6557);
  nor csa_tree_add_12_51_groupi_g15118__2398(csa_tree_add_12_51_groupi_n_6649 ,csa_tree_add_12_51_groupi_n_6551 ,csa_tree_add_12_51_groupi_n_6495);
  nor csa_tree_add_12_51_groupi_g15119__5107(csa_tree_add_12_51_groupi_n_6648 ,csa_tree_add_12_51_groupi_n_6553 ,csa_tree_add_12_51_groupi_n_5057);
  and csa_tree_add_12_51_groupi_g15120__6260(csa_tree_add_12_51_groupi_n_6647 ,csa_tree_add_12_51_groupi_n_6553 ,csa_tree_add_12_51_groupi_n_5057);
  or csa_tree_add_12_51_groupi_g15121__4319(csa_tree_add_12_51_groupi_n_6646 ,csa_tree_add_12_51_groupi_n_6504 ,csa_tree_add_12_51_groupi_n_6597);
  and csa_tree_add_12_51_groupi_g15122__8428(csa_tree_add_12_51_groupi_n_6645 ,csa_tree_add_12_51_groupi_n_6504 ,csa_tree_add_12_51_groupi_n_6597);
  nor csa_tree_add_12_51_groupi_g15123__5526(csa_tree_add_12_51_groupi_n_6644 ,csa_tree_add_12_51_groupi_n_6563 ,csa_tree_add_12_51_groupi_n_6427);
  nor csa_tree_add_12_51_groupi_g15124__6783(csa_tree_add_12_51_groupi_n_6643 ,csa_tree_add_12_51_groupi_n_6430 ,csa_tree_add_12_51_groupi_n_6583);
  and csa_tree_add_12_51_groupi_g15125__3680(csa_tree_add_12_51_groupi_n_6642 ,csa_tree_add_12_51_groupi_n_6492 ,csa_tree_add_12_51_groupi_n_6549);
  nor csa_tree_add_12_51_groupi_g15126__1617(csa_tree_add_12_51_groupi_n_6641 ,csa_tree_add_12_51_groupi_n_6492 ,csa_tree_add_12_51_groupi_n_6549);
  nor csa_tree_add_12_51_groupi_g15127__2802(csa_tree_add_12_51_groupi_n_6640 ,csa_tree_add_12_51_groupi_n_6469 ,csa_tree_add_12_51_groupi_n_6532);
  nor csa_tree_add_12_51_groupi_g15128__1705(csa_tree_add_12_51_groupi_n_6639 ,csa_tree_add_12_51_groupi_n_6595 ,csa_tree_add_12_51_groupi_n_5177);
  or csa_tree_add_12_51_groupi_g15129__5122(csa_tree_add_12_51_groupi_n_6638 ,csa_tree_add_12_51_groupi_n_6596 ,csa_tree_add_12_51_groupi_n_5176);
  or csa_tree_add_12_51_groupi_g15130__8246(csa_tree_add_12_51_groupi_n_6669 ,csa_tree_add_12_51_groupi_n_6478 ,csa_tree_add_12_51_groupi_n_6565);
  or csa_tree_add_12_51_groupi_g15131__7098(csa_tree_add_12_51_groupi_n_6668 ,csa_tree_add_12_51_groupi_n_6487 ,csa_tree_add_12_51_groupi_n_6531);
  not csa_tree_add_12_51_groupi_g15132(csa_tree_add_12_51_groupi_n_6632 ,csa_tree_add_12_51_groupi_n_6633);
  not csa_tree_add_12_51_groupi_g15133(csa_tree_add_12_51_groupi_n_6630 ,csa_tree_add_12_51_groupi_n_6631);
  not csa_tree_add_12_51_groupi_g15134(csa_tree_add_12_51_groupi_n_6628 ,csa_tree_add_12_51_groupi_n_6629);
  not csa_tree_add_12_51_groupi_g15135(csa_tree_add_12_51_groupi_n_6626 ,csa_tree_add_12_51_groupi_n_6627);
  and csa_tree_add_12_51_groupi_g15136__6131(csa_tree_add_12_51_groupi_n_6624 ,csa_tree_add_12_51_groupi_n_6560 ,csa_tree_add_12_51_groupi_n_4804);
  or csa_tree_add_12_51_groupi_g15137__1881(csa_tree_add_12_51_groupi_n_6623 ,csa_tree_add_12_51_groupi_n_6468 ,csa_tree_add_12_51_groupi_n_6589);
  nor csa_tree_add_12_51_groupi_g15138__5115(csa_tree_add_12_51_groupi_n_6622 ,csa_tree_add_12_51_groupi_n_6542 ,csa_tree_add_12_51_groupi_n_6446);
  and csa_tree_add_12_51_groupi_g15139__7482(csa_tree_add_12_51_groupi_n_6621 ,csa_tree_add_12_51_groupi_n_6542 ,csa_tree_add_12_51_groupi_n_6446);
  xnor csa_tree_add_12_51_groupi_g15140__4733(out3[10] ,csa_tree_add_12_51_groupi_n_6513 ,csa_tree_add_12_51_groupi_n_6436);
  and csa_tree_add_12_51_groupi_g15141__6161(csa_tree_add_12_51_groupi_n_6619 ,csa_tree_add_12_51_groupi_n_6529 ,csa_tree_add_12_51_groupi_n_6599);
  xnor csa_tree_add_12_51_groupi_g15142__9315(csa_tree_add_12_51_groupi_n_6618 ,csa_tree_add_12_51_groupi_n_6503 ,csa_tree_add_12_51_groupi_n_6306);
  xor csa_tree_add_12_51_groupi_g15143__9945(csa_tree_add_12_51_groupi_n_6617 ,csa_tree_add_12_51_groupi_n_6429 ,csa_tree_add_12_51_groupi_n_6492);
  xnor csa_tree_add_12_51_groupi_g15144__2883(csa_tree_add_12_51_groupi_n_6616 ,csa_tree_add_12_51_groupi_n_6497 ,csa_tree_add_12_51_groupi_n_6494);
  xnor csa_tree_add_12_51_groupi_g15145__2346(csa_tree_add_12_51_groupi_n_6615 ,csa_tree_add_12_51_groupi_n_6501 ,csa_tree_add_12_51_groupi_n_6309);
  xnor csa_tree_add_12_51_groupi_g15146__1666(csa_tree_add_12_51_groupi_n_6614 ,csa_tree_add_12_51_groupi_n_6099 ,csa_tree_add_12_51_groupi_n_6499);
  xnor csa_tree_add_12_51_groupi_g15147__7410(csa_tree_add_12_51_groupi_n_6613 ,csa_tree_add_12_51_groupi_n_6460 ,csa_tree_add_12_51_groupi_n_6491);
  xnor csa_tree_add_12_51_groupi_g15148__6417(csa_tree_add_12_51_groupi_n_6612 ,csa_tree_add_12_51_groupi_n_6490 ,csa_tree_add_12_51_groupi_n_6397);
  xnor csa_tree_add_12_51_groupi_g15149__5477(csa_tree_add_12_51_groupi_n_6611 ,csa_tree_add_12_51_groupi_n_6451 ,csa_tree_add_12_51_groupi_n_6450);
  xnor csa_tree_add_12_51_groupi_g15150__2398(csa_tree_add_12_51_groupi_n_6610 ,csa_tree_add_12_51_groupi_n_6458 ,csa_tree_add_12_51_groupi_n_6459);
  xnor csa_tree_add_12_51_groupi_g15151__5107(csa_tree_add_12_51_groupi_n_6609 ,csa_tree_add_12_51_groupi_n_6469 ,csa_tree_add_12_51_groupi_n_6299);
  xnor csa_tree_add_12_51_groupi_g15152__6260(csa_tree_add_12_51_groupi_n_6608 ,csa_tree_add_12_51_groupi_n_6508 ,csa_tree_add_12_51_groupi_n_6506);
  xnor csa_tree_add_12_51_groupi_g15153__4319(csa_tree_add_12_51_groupi_n_6607 ,csa_tree_add_12_51_groupi_n_6446 ,csa_tree_add_12_51_groupi_n_6400);
  xnor csa_tree_add_12_51_groupi_g15154__8428(csa_tree_add_12_51_groupi_n_6606 ,csa_tree_add_12_51_groupi_n_6461 ,csa_tree_add_12_51_groupi_n_6246);
  xnor csa_tree_add_12_51_groupi_g15155__5526(csa_tree_add_12_51_groupi_n_6605 ,csa_tree_add_12_51_groupi_n_6456 ,csa_tree_add_12_51_groupi_n_6457);
  xnor csa_tree_add_12_51_groupi_g15156__6783(csa_tree_add_12_51_groupi_n_6604 ,csa_tree_add_12_51_groupi_n_6502 ,csa_tree_add_12_51_groupi_n_6488);
  xnor csa_tree_add_12_51_groupi_g15157__3680(csa_tree_add_12_51_groupi_n_6603 ,csa_tree_add_12_51_groupi_n_6454 ,csa_tree_add_12_51_groupi_n_6455);
  xnor csa_tree_add_12_51_groupi_g15158__1617(csa_tree_add_12_51_groupi_n_6602 ,csa_tree_add_12_51_groupi_n_6208 ,csa_tree_add_12_51_groupi_n_6449);
  or csa_tree_add_12_51_groupi_g15159__2802(csa_tree_add_12_51_groupi_n_6637 ,csa_tree_add_12_51_groupi_n_6388 ,csa_tree_add_12_51_groupi_n_6523);
  xnor csa_tree_add_12_51_groupi_g15160__1705(csa_tree_add_12_51_groupi_n_6636 ,csa_tree_add_12_51_groupi_n_6399 ,csa_tree_add_12_51_groupi_n_6433);
  xnor csa_tree_add_12_51_groupi_g15161__5122(csa_tree_add_12_51_groupi_n_6635 ,csa_tree_add_12_51_groupi_n_6398 ,csa_tree_add_12_51_groupi_n_6437);
  xnor csa_tree_add_12_51_groupi_g15162__8246(csa_tree_add_12_51_groupi_n_6634 ,csa_tree_add_12_51_groupi_n_6307 ,csa_tree_add_12_51_groupi_n_6438);
  xnor csa_tree_add_12_51_groupi_g15163__7098(csa_tree_add_12_51_groupi_n_6633 ,csa_tree_add_12_51_groupi_n_6310 ,csa_tree_add_12_51_groupi_n_6432);
  xnor csa_tree_add_12_51_groupi_g15164__6131(csa_tree_add_12_51_groupi_n_6631 ,csa_tree_add_12_51_groupi_n_6315 ,csa_tree_add_12_51_groupi_n_6434);
  xnor csa_tree_add_12_51_groupi_g15165__1881(csa_tree_add_12_51_groupi_n_6629 ,csa_tree_add_12_51_groupi_n_6290 ,csa_tree_add_12_51_groupi_n_6440);
  xnor csa_tree_add_12_51_groupi_g15166__5115(csa_tree_add_12_51_groupi_n_6627 ,csa_tree_add_12_51_groupi_n_6289 ,csa_tree_add_12_51_groupi_n_6439);
  xnor csa_tree_add_12_51_groupi_g15167__7482(csa_tree_add_12_51_groupi_n_6625 ,csa_tree_add_12_51_groupi_n_6304 ,csa_tree_add_12_51_groupi_n_6435);
  not csa_tree_add_12_51_groupi_g15168(csa_tree_add_12_51_groupi_n_6595 ,csa_tree_add_12_51_groupi_n_6596);
  not csa_tree_add_12_51_groupi_g15169(csa_tree_add_12_51_groupi_n_6593 ,csa_tree_add_12_51_groupi_n_6594);
  and csa_tree_add_12_51_groupi_g15170__4733(csa_tree_add_12_51_groupi_n_6592 ,csa_tree_add_12_51_groupi_n_6500 ,csa_tree_add_12_51_groupi_n_6299);
  or csa_tree_add_12_51_groupi_g15171__6161(csa_tree_add_12_51_groupi_n_6591 ,csa_tree_add_12_51_groupi_n_6496 ,csa_tree_add_12_51_groupi_n_6493);
  nor csa_tree_add_12_51_groupi_g15172__9315(csa_tree_add_12_51_groupi_n_6590 ,csa_tree_add_12_51_groupi_n_6497 ,csa_tree_add_12_51_groupi_n_6494);
  nor csa_tree_add_12_51_groupi_g15173__9945(csa_tree_add_12_51_groupi_n_6589 ,csa_tree_add_12_51_groupi_n_6098 ,csa_tree_add_12_51_groupi_n_6499);
  and csa_tree_add_12_51_groupi_g15174__2883(csa_tree_add_12_51_groupi_n_6588 ,csa_tree_add_12_51_groupi_n_6503 ,csa_tree_add_12_51_groupi_n_6306);
  or csa_tree_add_12_51_groupi_g15175__2346(csa_tree_add_12_51_groupi_n_6587 ,csa_tree_add_12_51_groupi_n_6503 ,csa_tree_add_12_51_groupi_n_6306);
  and csa_tree_add_12_51_groupi_g15176__1666(csa_tree_add_12_51_groupi_n_6586 ,csa_tree_add_12_51_groupi_n_6460 ,csa_tree_add_12_51_groupi_n_6491);
  or csa_tree_add_12_51_groupi_g15177__7410(csa_tree_add_12_51_groupi_n_6585 ,csa_tree_add_12_51_groupi_n_6099 ,csa_tree_add_12_51_groupi_n_6498);
  or csa_tree_add_12_51_groupi_g15178__6417(csa_tree_add_12_51_groupi_n_6584 ,csa_tree_add_12_51_groupi_n_6460 ,csa_tree_add_12_51_groupi_n_6491);
  nor csa_tree_add_12_51_groupi_g15179__5477(csa_tree_add_12_51_groupi_n_6583 ,csa_tree_add_12_51_groupi_n_6293 ,csa_tree_add_12_51_groupi_n_6445);
  or csa_tree_add_12_51_groupi_g15180__2398(csa_tree_add_12_51_groupi_n_6582 ,csa_tree_add_12_51_groupi_n_6459 ,csa_tree_add_12_51_groupi_n_6458);
  and csa_tree_add_12_51_groupi_g15181__5107(csa_tree_add_12_51_groupi_n_6581 ,csa_tree_add_12_51_groupi_n_6459 ,csa_tree_add_12_51_groupi_n_6458);
  nor csa_tree_add_12_51_groupi_g15182__6260(csa_tree_add_12_51_groupi_n_6580 ,csa_tree_add_12_51_groupi_n_6208 ,csa_tree_add_12_51_groupi_n_6449);
  and csa_tree_add_12_51_groupi_g15183__4319(csa_tree_add_12_51_groupi_n_6579 ,csa_tree_add_12_51_groupi_n_6450 ,csa_tree_add_12_51_groupi_n_6451);
  and csa_tree_add_12_51_groupi_g15184__8428(csa_tree_add_12_51_groupi_n_6578 ,csa_tree_add_12_51_groupi_n_6502 ,csa_tree_add_12_51_groupi_n_6488);
  or csa_tree_add_12_51_groupi_g15185__5526(csa_tree_add_12_51_groupi_n_6577 ,csa_tree_add_12_51_groupi_n_6502 ,csa_tree_add_12_51_groupi_n_6488);
  or csa_tree_add_12_51_groupi_g15186__6783(csa_tree_add_12_51_groupi_n_6576 ,csa_tree_add_12_51_groupi_n_6442 ,csa_tree_add_12_51_groupi_n_6447);
  and csa_tree_add_12_51_groupi_g15187__3680(csa_tree_add_12_51_groupi_n_6575 ,csa_tree_add_12_51_groupi_n_6208 ,csa_tree_add_12_51_groupi_n_6449);
  or csa_tree_add_12_51_groupi_g15188__1617(csa_tree_add_12_51_groupi_n_6574 ,csa_tree_add_12_51_groupi_n_6507 ,csa_tree_add_12_51_groupi_n_6505);
  and csa_tree_add_12_51_groupi_g15189__2802(csa_tree_add_12_51_groupi_n_6573 ,csa_tree_add_12_51_groupi_n_6442 ,csa_tree_add_12_51_groupi_n_6447);
  nor csa_tree_add_12_51_groupi_g15190__1705(csa_tree_add_12_51_groupi_n_6572 ,csa_tree_add_12_51_groupi_n_6508 ,csa_tree_add_12_51_groupi_n_6506);
  or csa_tree_add_12_51_groupi_g15191__5122(csa_tree_add_12_51_groupi_n_6571 ,csa_tree_add_12_51_groupi_n_6457 ,csa_tree_add_12_51_groupi_n_6456);
  and csa_tree_add_12_51_groupi_g15192__8246(csa_tree_add_12_51_groupi_n_6570 ,csa_tree_add_12_51_groupi_n_6501 ,csa_tree_add_12_51_groupi_n_6309);
  or csa_tree_add_12_51_groupi_g15193__7098(csa_tree_add_12_51_groupi_n_6569 ,csa_tree_add_12_51_groupi_n_6501 ,csa_tree_add_12_51_groupi_n_6309);
  or csa_tree_add_12_51_groupi_g15194__6131(csa_tree_add_12_51_groupi_n_6568 ,csa_tree_add_12_51_groupi_n_6450 ,csa_tree_add_12_51_groupi_n_6451);
  and csa_tree_add_12_51_groupi_g15195__1881(csa_tree_add_12_51_groupi_n_6567 ,csa_tree_add_12_51_groupi_n_6457 ,csa_tree_add_12_51_groupi_n_6456);
  and csa_tree_add_12_51_groupi_g15196__5115(csa_tree_add_12_51_groupi_n_6566 ,csa_tree_add_12_51_groupi_n_6293 ,csa_tree_add_12_51_groupi_n_6445);
  nor csa_tree_add_12_51_groupi_g15197__7482(csa_tree_add_12_51_groupi_n_6565 ,csa_tree_add_12_51_groupi_n_6479 ,csa_tree_add_12_51_groupi_n_6254);
  and csa_tree_add_12_51_groupi_g15198__4733(csa_tree_add_12_51_groupi_n_6564 ,csa_tree_add_12_51_groupi_n_6296 ,csa_tree_add_12_51_groupi_n_6448);
  nor csa_tree_add_12_51_groupi_g15199__6161(csa_tree_add_12_51_groupi_n_6563 ,csa_tree_add_12_51_groupi_n_6296 ,csa_tree_add_12_51_groupi_n_6448);
  or csa_tree_add_12_51_groupi_g15200__9315(csa_tree_add_12_51_groupi_n_6601 ,csa_tree_add_12_51_groupi_n_6415 ,csa_tree_add_12_51_groupi_n_6485);
  or csa_tree_add_12_51_groupi_g15201__9945(csa_tree_add_12_51_groupi_n_6600 ,csa_tree_add_12_51_groupi_n_6405 ,csa_tree_add_12_51_groupi_n_6476);
  or csa_tree_add_12_51_groupi_g15202__2883(csa_tree_add_12_51_groupi_n_6599 ,csa_tree_add_12_51_groupi_n_6411 ,csa_tree_add_12_51_groupi_n_6481);
  or csa_tree_add_12_51_groupi_g15203__2346(csa_tree_add_12_51_groupi_n_6598 ,csa_tree_add_12_51_groupi_n_6416 ,csa_tree_add_12_51_groupi_n_6484);
  or csa_tree_add_12_51_groupi_g15204__1666(csa_tree_add_12_51_groupi_n_6597 ,csa_tree_add_12_51_groupi_n_6419 ,csa_tree_add_12_51_groupi_n_6486);
  or csa_tree_add_12_51_groupi_g15205__7410(csa_tree_add_12_51_groupi_n_6596 ,csa_tree_add_12_51_groupi_n_6421 ,csa_tree_add_12_51_groupi_n_6475);
  or csa_tree_add_12_51_groupi_g15206__6417(csa_tree_add_12_51_groupi_n_6594 ,csa_tree_add_12_51_groupi_n_6409 ,csa_tree_add_12_51_groupi_n_6480);
  not csa_tree_add_12_51_groupi_g15207(csa_tree_add_12_51_groupi_n_6555 ,csa_tree_add_12_51_groupi_n_6556);
  not csa_tree_add_12_51_groupi_g15208(csa_tree_add_12_51_groupi_n_6551 ,csa_tree_add_12_51_groupi_n_6550);
  not csa_tree_add_12_51_groupi_g15209(csa_tree_add_12_51_groupi_n_6548 ,csa_tree_add_12_51_groupi_n_6547);
  not csa_tree_add_12_51_groupi_g15210(csa_tree_add_12_51_groupi_n_6545 ,csa_tree_add_12_51_groupi_n_6546);
  not csa_tree_add_12_51_groupi_g15211(csa_tree_add_12_51_groupi_n_6543 ,csa_tree_add_12_51_groupi_n_6544);
  not csa_tree_add_12_51_groupi_g15212(csa_tree_add_12_51_groupi_n_6540 ,csa_tree_add_12_51_groupi_n_6539);
  not csa_tree_add_12_51_groupi_g15213(csa_tree_add_12_51_groupi_n_6535 ,csa_tree_add_12_51_groupi_n_6536);
  not csa_tree_add_12_51_groupi_g15214(csa_tree_add_12_51_groupi_n_6533 ,csa_tree_add_12_51_groupi_n_6534);
  nor csa_tree_add_12_51_groupi_g15215__5477(csa_tree_add_12_51_groupi_n_6532 ,csa_tree_add_12_51_groupi_n_6500 ,csa_tree_add_12_51_groupi_n_6299);
  nor csa_tree_add_12_51_groupi_g15216__2398(csa_tree_add_12_51_groupi_n_6531 ,csa_tree_add_12_51_groupi_n_6477 ,csa_tree_add_12_51_groupi_n_6253);
  nor csa_tree_add_12_51_groupi_g15217__5107(csa_tree_add_12_51_groupi_n_6530 ,csa_tree_add_12_51_groupi_n_6489 ,csa_tree_add_12_51_groupi_n_6397);
  or csa_tree_add_12_51_groupi_g15218__6260(csa_tree_add_12_51_groupi_n_6529 ,csa_tree_add_12_51_groupi_n_6490 ,csa_tree_add_12_51_groupi_n_6396);
  and csa_tree_add_12_51_groupi_g15219__4319(csa_tree_add_12_51_groupi_n_6528 ,csa_tree_add_12_51_groupi_n_6461 ,csa_tree_add_12_51_groupi_n_6246);
  or csa_tree_add_12_51_groupi_g15220__8428(csa_tree_add_12_51_groupi_n_6527 ,csa_tree_add_12_51_groupi_n_6455 ,csa_tree_add_12_51_groupi_n_6454);
  and csa_tree_add_12_51_groupi_g15221__5526(csa_tree_add_12_51_groupi_n_6526 ,csa_tree_add_12_51_groupi_n_6455 ,csa_tree_add_12_51_groupi_n_6454);
  nor csa_tree_add_12_51_groupi_g15222__6783(csa_tree_add_12_51_groupi_n_6525 ,csa_tree_add_12_51_groupi_n_6444 ,csa_tree_add_12_51_groupi_n_6424);
  or csa_tree_add_12_51_groupi_g15223__3680(csa_tree_add_12_51_groupi_n_6524 ,csa_tree_add_12_51_groupi_n_6443 ,csa_tree_add_12_51_groupi_n_6425);
  and csa_tree_add_12_51_groupi_g15224__1617(csa_tree_add_12_51_groupi_n_6523 ,csa_tree_add_12_51_groupi_n_6387 ,csa_tree_add_12_51_groupi_n_6513);
  or csa_tree_add_12_51_groupi_g15225__2802(csa_tree_add_12_51_groupi_n_6522 ,csa_tree_add_12_51_groupi_n_6461 ,csa_tree_add_12_51_groupi_n_6246);
  xnor csa_tree_add_12_51_groupi_g15226__1705(csa_tree_add_12_51_groupi_n_6521 ,csa_tree_add_12_51_groupi_n_6426 ,csa_tree_add_12_51_groupi_n_6395);
  xor csa_tree_add_12_51_groupi_g15227__5122(csa_tree_add_12_51_groupi_n_6520 ,csa_tree_add_12_51_groupi_n_6296 ,csa_tree_add_12_51_groupi_n_6427);
  xnor csa_tree_add_12_51_groupi_g15228__8246(csa_tree_add_12_51_groupi_n_6519 ,csa_tree_add_12_51_groupi_n_6428 ,csa_tree_add_12_51_groupi_n_6425);
  xor csa_tree_add_12_51_groupi_g15229__7098(csa_tree_add_12_51_groupi_n_6518 ,csa_tree_add_12_51_groupi_n_6293 ,csa_tree_add_12_51_groupi_n_6430);
  xnor csa_tree_add_12_51_groupi_g15230__6131(csa_tree_add_12_51_groupi_n_6517 ,csa_tree_add_12_51_groupi_n_6431 ,csa_tree_add_12_51_groupi_n_6368);
  xnor csa_tree_add_12_51_groupi_g15231__1881(csa_tree_add_12_51_groupi_n_6562 ,csa_tree_add_12_51_groupi_n_6378 ,in3[14]);
  xnor csa_tree_add_12_51_groupi_g15232__5115(csa_tree_add_12_51_groupi_n_6561 ,csa_tree_add_12_51_groupi_n_6211 ,csa_tree_add_12_51_groupi_n_6377);
  xnor csa_tree_add_12_51_groupi_g15233__7482(csa_tree_add_12_51_groupi_n_6560 ,csa_tree_add_12_51_groupi_n_6384 ,in4[14]);
  xnor csa_tree_add_12_51_groupi_g15234__4733(csa_tree_add_12_51_groupi_n_6559 ,csa_tree_add_12_51_groupi_n_6382 ,in3[5]);
  xnor csa_tree_add_12_51_groupi_g15235__6161(csa_tree_add_12_51_groupi_n_6558 ,csa_tree_add_12_51_groupi_n_6372 ,in3[8]);
  xnor csa_tree_add_12_51_groupi_g15236__9315(csa_tree_add_12_51_groupi_n_6557 ,csa_tree_add_12_51_groupi_n_6402 ,in3[2]);
  xnor csa_tree_add_12_51_groupi_g15237__9945(csa_tree_add_12_51_groupi_n_6556 ,csa_tree_add_12_51_groupi_n_6385 ,in4[8]);
  xnor csa_tree_add_12_51_groupi_g15238__2883(csa_tree_add_12_51_groupi_n_6554 ,csa_tree_add_12_51_groupi_n_104 ,csa_tree_add_12_51_groupi_n_6403);
  xnor csa_tree_add_12_51_groupi_g15239__2346(csa_tree_add_12_51_groupi_n_6553 ,csa_tree_add_12_51_groupi_n_6381 ,in2[14]);
  xnor csa_tree_add_12_51_groupi_g15240__1666(csa_tree_add_12_51_groupi_n_6552 ,csa_tree_add_12_51_groupi_n_6401 ,in4[2]);
  xnor csa_tree_add_12_51_groupi_g15241__7410(csa_tree_add_12_51_groupi_n_6550 ,csa_tree_add_12_51_groupi_n_6379 ,in2[8]);
  xnor csa_tree_add_12_51_groupi_g15242__6417(csa_tree_add_12_51_groupi_n_6549 ,csa_tree_add_12_51_groupi_n_6303 ,csa_tree_add_12_51_groupi_n_14);
  xnor csa_tree_add_12_51_groupi_g15243__5477(csa_tree_add_12_51_groupi_n_6547 ,csa_tree_add_12_51_groupi_n_6207 ,csa_tree_add_12_51_groupi_n_6376);
  xnor csa_tree_add_12_51_groupi_g15244__2398(csa_tree_add_12_51_groupi_n_6546 ,csa_tree_add_12_51_groupi_n_6374 ,in4[11]);
  xnor csa_tree_add_12_51_groupi_g15245__5107(csa_tree_add_12_51_groupi_n_6544 ,csa_tree_add_12_51_groupi_n_6373 ,in2[11]);
  xnor csa_tree_add_12_51_groupi_g15246__6260(csa_tree_add_12_51_groupi_n_6542 ,csa_tree_add_12_51_groupi_n_6294 ,csa_tree_add_12_51_groupi_n_6370);
  or csa_tree_add_12_51_groupi_g15247__4319(csa_tree_add_12_51_groupi_n_6541 ,csa_tree_add_12_51_groupi_n_6390 ,csa_tree_add_12_51_groupi_n_6474);
  xnor csa_tree_add_12_51_groupi_g15248__8428(csa_tree_add_12_51_groupi_n_6539 ,csa_tree_add_12_51_groupi_n_6209 ,csa_tree_add_12_51_groupi_n_6375);
  xnor csa_tree_add_12_51_groupi_g15249__5526(csa_tree_add_12_51_groupi_n_6538 ,csa_tree_add_12_51_groupi_n_6371 ,in3[11]);
  xnor csa_tree_add_12_51_groupi_g15250__6783(csa_tree_add_12_51_groupi_n_6537 ,csa_tree_add_12_51_groupi_n_6383 ,in2[5]);
  xnor csa_tree_add_12_51_groupi_g15251__3680(csa_tree_add_12_51_groupi_n_6536 ,csa_tree_add_12_51_groupi_n_6380 ,in4[5]);
  or csa_tree_add_12_51_groupi_g15252__1617(csa_tree_add_12_51_groupi_n_6534 ,csa_tree_add_12_51_groupi_n_6407 ,csa_tree_add_12_51_groupi_n_6473);
  not csa_tree_add_12_51_groupi_g15253(csa_tree_add_12_51_groupi_n_6515 ,csa_tree_add_12_51_groupi_n_6514);
  not csa_tree_add_12_51_groupi_g15254(csa_tree_add_12_51_groupi_n_6512 ,csa_tree_add_12_51_groupi_n_6511);
  not csa_tree_add_12_51_groupi_g15255(csa_tree_add_12_51_groupi_n_6507 ,csa_tree_add_12_51_groupi_n_6508);
  not csa_tree_add_12_51_groupi_g15256(csa_tree_add_12_51_groupi_n_6505 ,csa_tree_add_12_51_groupi_n_6506);
  not csa_tree_add_12_51_groupi_g15257(csa_tree_add_12_51_groupi_n_6498 ,csa_tree_add_12_51_groupi_n_6499);
  not csa_tree_add_12_51_groupi_g15258(csa_tree_add_12_51_groupi_n_6496 ,csa_tree_add_12_51_groupi_n_6497);
  not csa_tree_add_12_51_groupi_g15259(csa_tree_add_12_51_groupi_n_6493 ,csa_tree_add_12_51_groupi_n_6494);
  not csa_tree_add_12_51_groupi_g15260(csa_tree_add_12_51_groupi_n_6489 ,csa_tree_add_12_51_groupi_n_6490);
  and csa_tree_add_12_51_groupi_g15261__2802(csa_tree_add_12_51_groupi_n_6487 ,csa_tree_add_12_51_groupi_n_6398 ,csa_tree_add_12_51_groupi_n_6302);
  nor csa_tree_add_12_51_groupi_g15262__1705(csa_tree_add_12_51_groupi_n_6486 ,csa_tree_add_12_51_groupi_n_6418 ,csa_tree_add_12_51_groupi_n_6214);
  nor csa_tree_add_12_51_groupi_g15263__5122(csa_tree_add_12_51_groupi_n_6485 ,csa_tree_add_12_51_groupi_n_6312 ,csa_tree_add_12_51_groupi_n_6414);
  and csa_tree_add_12_51_groupi_g15264__8246(csa_tree_add_12_51_groupi_n_6484 ,csa_tree_add_12_51_groupi_n_6315 ,csa_tree_add_12_51_groupi_n_6413);
  and csa_tree_add_12_51_groupi_g15265__7098(csa_tree_add_12_51_groupi_n_6483 ,csa_tree_add_12_51_groupi_n_6426 ,csa_tree_add_12_51_groupi_n_6395);
  nor csa_tree_add_12_51_groupi_g15266__6131(csa_tree_add_12_51_groupi_n_6482 ,csa_tree_add_12_51_groupi_n_6426 ,csa_tree_add_12_51_groupi_n_6395);
  nor csa_tree_add_12_51_groupi_g15267__1881(csa_tree_add_12_51_groupi_n_6481 ,csa_tree_add_12_51_groupi_n_6410 ,csa_tree_add_12_51_groupi_n_6252);
  nor csa_tree_add_12_51_groupi_g15268__5115(csa_tree_add_12_51_groupi_n_6480 ,csa_tree_add_12_51_groupi_n_6408 ,csa_tree_add_12_51_groupi_n_6369);
  nor csa_tree_add_12_51_groupi_g15269__7482(csa_tree_add_12_51_groupi_n_6479 ,csa_tree_add_12_51_groupi_n_6288 ,csa_tree_add_12_51_groupi_n_6399);
  and csa_tree_add_12_51_groupi_g15270__4733(csa_tree_add_12_51_groupi_n_6478 ,csa_tree_add_12_51_groupi_n_6288 ,csa_tree_add_12_51_groupi_n_6399);
  nor csa_tree_add_12_51_groupi_g15271__6161(csa_tree_add_12_51_groupi_n_6477 ,csa_tree_add_12_51_groupi_n_6398 ,csa_tree_add_12_51_groupi_n_6302);
  and csa_tree_add_12_51_groupi_g15272__9315(csa_tree_add_12_51_groupi_n_6476 ,csa_tree_add_12_51_groupi_n_6431 ,csa_tree_add_12_51_groupi_n_6406);
  nor csa_tree_add_12_51_groupi_g15273__9945(csa_tree_add_12_51_groupi_n_6475 ,csa_tree_add_12_51_groupi_n_6314 ,csa_tree_add_12_51_groupi_n_6420);
  nor csa_tree_add_12_51_groupi_g15274__2883(csa_tree_add_12_51_groupi_n_6474 ,csa_tree_add_12_51_groupi_n_6389 ,csa_tree_add_12_51_groupi_n_6251);
  nor csa_tree_add_12_51_groupi_g15275__2346(csa_tree_add_12_51_groupi_n_6473 ,csa_tree_add_12_51_groupi_n_6257 ,csa_tree_add_12_51_groupi_n_6412);
  xnor csa_tree_add_12_51_groupi_g15276__1666(csa_tree_add_12_51_groupi_n_6516 ,csa_tree_add_12_51_groupi_n_6338 ,in2[5]);
  xnor csa_tree_add_12_51_groupi_g15277__7410(csa_tree_add_12_51_groupi_n_6514 ,csa_tree_add_12_51_groupi_n_6336 ,in3[14]);
  or csa_tree_add_12_51_groupi_g15278__6417(csa_tree_add_12_51_groupi_n_6513 ,csa_tree_add_12_51_groupi_n_6392 ,csa_tree_add_12_51_groupi_n_6185);
  xnor csa_tree_add_12_51_groupi_g15279__5477(csa_tree_add_12_51_groupi_n_6511 ,csa_tree_add_12_51_groupi_n_6343 ,in2[2]);
  xnor csa_tree_add_12_51_groupi_g15280__2398(csa_tree_add_12_51_groupi_n_6510 ,csa_tree_add_12_51_groupi_n_6339 ,in3[11]);
  or csa_tree_add_12_51_groupi_g15281__5107(csa_tree_add_12_51_groupi_n_6509 ,csa_tree_add_12_51_groupi_n_6386 ,csa_tree_add_12_51_groupi_n_6360);
  xnor csa_tree_add_12_51_groupi_g15282__6260(csa_tree_add_12_51_groupi_n_6508 ,csa_tree_add_12_51_groupi_n_6334 ,in4[14]);
  xnor csa_tree_add_12_51_groupi_g15283__4319(csa_tree_add_12_51_groupi_n_6506 ,csa_tree_add_12_51_groupi_n_6335 ,in2[14]);
  xnor csa_tree_add_12_51_groupi_g15284__8428(csa_tree_add_12_51_groupi_n_6504 ,csa_tree_add_12_51_groupi_n_6344 ,in3[2]);
  xnor csa_tree_add_12_51_groupi_g15285__5526(csa_tree_add_12_51_groupi_n_6503 ,csa_tree_add_12_51_groupi_n_6341 ,in4[11]);
  xnor csa_tree_add_12_51_groupi_g15286__6783(csa_tree_add_12_51_groupi_n_6502 ,csa_tree_add_12_51_groupi_n_6333 ,in2[11]);
  xnor csa_tree_add_12_51_groupi_g15287__3680(csa_tree_add_12_51_groupi_n_6501 ,csa_tree_add_12_51_groupi_n_6337 ,in4[5]);
  or csa_tree_add_12_51_groupi_g15288__1617(csa_tree_add_12_51_groupi_n_6500 ,csa_tree_add_12_51_groupi_n_6422 ,csa_tree_add_12_51_groupi_n_6356);
  xnor csa_tree_add_12_51_groupi_g15289__2802(csa_tree_add_12_51_groupi_n_6499 ,csa_tree_add_12_51_groupi_n_6104 ,csa_tree_add_12_51_groupi_n_6259);
  xnor csa_tree_add_12_51_groupi_g15290__1705(csa_tree_add_12_51_groupi_n_6497 ,csa_tree_add_12_51_groupi_n_6342 ,in4[2]);
  and csa_tree_add_12_51_groupi_g15291__5122(csa_tree_add_12_51_groupi_n_6495 ,csa_tree_add_12_51_groupi_n_6361 ,csa_tree_add_12_51_groupi_n_6417);
  or csa_tree_add_12_51_groupi_g15292__8246(csa_tree_add_12_51_groupi_n_6494 ,csa_tree_add_12_51_groupi_n_6404 ,csa_tree_add_12_51_groupi_n_6349);
  xnor csa_tree_add_12_51_groupi_g15293__7098(csa_tree_add_12_51_groupi_n_6492 ,csa_tree_add_12_51_groupi_n_6109 ,csa_tree_add_12_51_groupi_n_6261);
  xnor csa_tree_add_12_51_groupi_g15294__6131(csa_tree_add_12_51_groupi_n_6491 ,csa_tree_add_12_51_groupi_n_6332 ,in3[8]);
  xnor csa_tree_add_12_51_groupi_g15295__1881(csa_tree_add_12_51_groupi_n_6490 ,csa_tree_add_12_51_groupi_n_6340 ,in3[5]);
  or csa_tree_add_12_51_groupi_g15296__5115(csa_tree_add_12_51_groupi_n_6488 ,csa_tree_add_12_51_groupi_n_6353 ,csa_tree_add_12_51_groupi_n_6391);
  not csa_tree_add_12_51_groupi_g15297(csa_tree_add_12_51_groupi_n_6468 ,csa_tree_add_12_51_groupi_n_6467);
  not csa_tree_add_12_51_groupi_g15298(csa_tree_add_12_51_groupi_n_6464 ,csa_tree_add_12_51_groupi_n_6465);
  not csa_tree_add_12_51_groupi_g15299(csa_tree_add_12_51_groupi_n_6462 ,csa_tree_add_12_51_groupi_n_6463);
  not csa_tree_add_12_51_groupi_g15300(csa_tree_add_12_51_groupi_n_6452 ,csa_tree_add_12_51_groupi_n_6453);
  not csa_tree_add_12_51_groupi_g15301(csa_tree_add_12_51_groupi_n_6443 ,csa_tree_add_12_51_groupi_n_6444);
  xnor csa_tree_add_12_51_groupi_g15302__7482(out3[9] ,csa_tree_add_12_51_groupi_n_6313 ,csa_tree_add_12_51_groupi_n_6267);
  xnor csa_tree_add_12_51_groupi_g15303__4733(csa_tree_add_12_51_groupi_n_6440 ,csa_tree_add_12_51_groupi_n_6314 ,csa_tree_add_12_51_groupi_n_6292);
  xnor csa_tree_add_12_51_groupi_g15304__6161(csa_tree_add_12_51_groupi_n_6439 ,csa_tree_add_12_51_groupi_n_6297 ,csa_tree_add_12_51_groupi_n_6252);
  xnor csa_tree_add_12_51_groupi_g15305__9315(csa_tree_add_12_51_groupi_n_6438 ,csa_tree_add_12_51_groupi_n_6369 ,csa_tree_add_12_51_groupi_n_6245);
  xor csa_tree_add_12_51_groupi_g15306__9945(csa_tree_add_12_51_groupi_n_6437 ,csa_tree_add_12_51_groupi_n_6253 ,csa_tree_add_12_51_groupi_n_6302);
  xnor csa_tree_add_12_51_groupi_g15307__2883(csa_tree_add_12_51_groupi_n_6436 ,csa_tree_add_12_51_groupi_n_6169 ,csa_tree_add_12_51_groupi_n_6301);
  xnor csa_tree_add_12_51_groupi_g15308__2346(csa_tree_add_12_51_groupi_n_6435 ,csa_tree_add_12_51_groupi_n_6214 ,csa_tree_add_12_51_groupi_n_6295);
  xnor csa_tree_add_12_51_groupi_g15309__1666(csa_tree_add_12_51_groupi_n_6434 ,csa_tree_add_12_51_groupi_n_6300 ,csa_tree_add_12_51_groupi_n_6298);
  xor csa_tree_add_12_51_groupi_g15310__7410(csa_tree_add_12_51_groupi_n_6433 ,csa_tree_add_12_51_groupi_n_6288 ,csa_tree_add_12_51_groupi_n_6254);
  xnor csa_tree_add_12_51_groupi_g15311__6417(csa_tree_add_12_51_groupi_n_6432 ,csa_tree_add_12_51_groupi_n_6312 ,csa_tree_add_12_51_groupi_n_6287);
  xnor csa_tree_add_12_51_groupi_g15312__5477(csa_tree_add_12_51_groupi_n_6472 ,csa_tree_add_12_51_groupi_n_6122 ,csa_tree_add_12_51_groupi_n_6264);
  xnor csa_tree_add_12_51_groupi_g15313__2398(csa_tree_add_12_51_groupi_n_6471 ,csa_tree_add_12_51_groupi_n_6321 ,in3[14]);
  xnor csa_tree_add_12_51_groupi_g15314__5107(csa_tree_add_12_51_groupi_n_6470 ,csa_tree_add_12_51_groupi_n_6317 ,in3[11]);
  xnor csa_tree_add_12_51_groupi_g15315__6260(csa_tree_add_12_51_groupi_n_6469 ,csa_tree_add_12_51_groupi_n_1924 ,csa_tree_add_12_51_groupi_n_6330);
  xnor csa_tree_add_12_51_groupi_g15316__4319(csa_tree_add_12_51_groupi_n_6467 ,csa_tree_add_12_51_groupi_n_6248 ,csa_tree_add_12_51_groupi_n_6260);
  xnor csa_tree_add_12_51_groupi_g15317__8428(csa_tree_add_12_51_groupi_n_6466 ,csa_tree_add_12_51_groupi_n_6250 ,csa_tree_add_12_51_groupi_n_6268);
  xnor csa_tree_add_12_51_groupi_g15318__5526(csa_tree_add_12_51_groupi_n_6465 ,csa_tree_add_12_51_groupi_n_6322 ,in4[8]);
  xnor csa_tree_add_12_51_groupi_g15319__6783(csa_tree_add_12_51_groupi_n_6463 ,csa_tree_add_12_51_groupi_n_6324 ,in3[5]);
  xnor csa_tree_add_12_51_groupi_g15320__3680(csa_tree_add_12_51_groupi_n_6461 ,csa_tree_add_12_51_groupi_n_6215 ,csa_tree_add_12_51_groupi_n_6265);
  xnor csa_tree_add_12_51_groupi_g15321__1617(csa_tree_add_12_51_groupi_n_6460 ,csa_tree_add_12_51_groupi_n_6331 ,in4[8]);
  xnor csa_tree_add_12_51_groupi_g15322__2802(csa_tree_add_12_51_groupi_n_6459 ,csa_tree_add_12_51_groupi_n_6320 ,in4[5]);
  xnor csa_tree_add_12_51_groupi_g15323__1705(csa_tree_add_12_51_groupi_n_6458 ,csa_tree_add_12_51_groupi_n_6319 ,in2[5]);
  xnor csa_tree_add_12_51_groupi_g15324__5122(csa_tree_add_12_51_groupi_n_6457 ,csa_tree_add_12_51_groupi_n_6316 ,in4[11]);
  xnor csa_tree_add_12_51_groupi_g15325__8246(csa_tree_add_12_51_groupi_n_6456 ,csa_tree_add_12_51_groupi_n_6329 ,in2[11]);
  xnor csa_tree_add_12_51_groupi_g15326__7098(csa_tree_add_12_51_groupi_n_6455 ,csa_tree_add_12_51_groupi_n_6345 ,in4[2]);
  xnor csa_tree_add_12_51_groupi_g15327__6131(csa_tree_add_12_51_groupi_n_6454 ,csa_tree_add_12_51_groupi_n_6328 ,in2[2]);
  xnor csa_tree_add_12_51_groupi_g15328__1881(csa_tree_add_12_51_groupi_n_6453 ,csa_tree_add_12_51_groupi_n_6327 ,in3[2]);
  xnor csa_tree_add_12_51_groupi_g15329__5115(csa_tree_add_12_51_groupi_n_6451 ,csa_tree_add_12_51_groupi_n_6326 ,in2[14]);
  xnor csa_tree_add_12_51_groupi_g15330__7482(csa_tree_add_12_51_groupi_n_6450 ,csa_tree_add_12_51_groupi_n_6323 ,in4[14]);
  xnor csa_tree_add_12_51_groupi_g15331__4733(csa_tree_add_12_51_groupi_n_6449 ,csa_tree_add_12_51_groupi_n_6118 ,csa_tree_add_12_51_groupi_n_6262);
  xnor csa_tree_add_12_51_groupi_g15332__6161(csa_tree_add_12_51_groupi_n_6448 ,csa_tree_add_12_51_groupi_n_6213 ,csa_tree_add_12_51_groupi_n_6269);
  xnor csa_tree_add_12_51_groupi_g15333__9315(csa_tree_add_12_51_groupi_n_6447 ,csa_tree_add_12_51_groupi_n_6318 ,in3[8]);
  xnor csa_tree_add_12_51_groupi_g15334__9945(csa_tree_add_12_51_groupi_n_6446 ,csa_tree_add_12_51_groupi_n_6090 ,csa_tree_add_12_51_groupi_n_6266);
  xnor csa_tree_add_12_51_groupi_g15335__2883(csa_tree_add_12_51_groupi_n_6445 ,csa_tree_add_12_51_groupi_n_6212 ,csa_tree_add_12_51_groupi_n_6263);
  xnor csa_tree_add_12_51_groupi_g15336__2346(csa_tree_add_12_51_groupi_n_6444 ,csa_tree_add_12_51_groupi_n_6210 ,csa_tree_add_12_51_groupi_n_6270);
  xnor csa_tree_add_12_51_groupi_g15337__1666(csa_tree_add_12_51_groupi_n_6442 ,csa_tree_add_12_51_groupi_n_6325 ,in2[8]);
  not csa_tree_add_12_51_groupi_g15338(csa_tree_add_12_51_groupi_n_6425 ,csa_tree_add_12_51_groupi_n_6424);
  nor csa_tree_add_12_51_groupi_g15339__7410(csa_tree_add_12_51_groupi_n_6422 ,csa_tree_add_12_51_groupi_n_6258 ,csa_tree_add_12_51_groupi_n_6355);
  nor csa_tree_add_12_51_groupi_g15340__6417(csa_tree_add_12_51_groupi_n_6421 ,csa_tree_add_12_51_groupi_n_6292 ,csa_tree_add_12_51_groupi_n_6291);
  and csa_tree_add_12_51_groupi_g15341__5477(csa_tree_add_12_51_groupi_n_6420 ,csa_tree_add_12_51_groupi_n_6292 ,csa_tree_add_12_51_groupi_n_6291);
  nor csa_tree_add_12_51_groupi_g15342__2398(csa_tree_add_12_51_groupi_n_6419 ,csa_tree_add_12_51_groupi_n_6295 ,csa_tree_add_12_51_groupi_n_6305);
  and csa_tree_add_12_51_groupi_g15343__5107(csa_tree_add_12_51_groupi_n_6418 ,csa_tree_add_12_51_groupi_n_6295 ,csa_tree_add_12_51_groupi_n_6305);
  or csa_tree_add_12_51_groupi_g15344__6260(csa_tree_add_12_51_groupi_n_6417 ,csa_tree_add_12_51_groupi_n_6362 ,csa_tree_add_12_51_groupi_n_6247);
  and csa_tree_add_12_51_groupi_g15345__4319(csa_tree_add_12_51_groupi_n_6416 ,csa_tree_add_12_51_groupi_n_6300 ,csa_tree_add_12_51_groupi_n_6298);
  nor csa_tree_add_12_51_groupi_g15346__8428(csa_tree_add_12_51_groupi_n_6415 ,csa_tree_add_12_51_groupi_n_6287 ,csa_tree_add_12_51_groupi_n_6311);
  and csa_tree_add_12_51_groupi_g15347__5526(csa_tree_add_12_51_groupi_n_6414 ,csa_tree_add_12_51_groupi_n_6287 ,csa_tree_add_12_51_groupi_n_6311);
  or csa_tree_add_12_51_groupi_g15348__6783(csa_tree_add_12_51_groupi_n_6413 ,csa_tree_add_12_51_groupi_n_6300 ,csa_tree_add_12_51_groupi_n_6298);
  and csa_tree_add_12_51_groupi_g15349__3680(csa_tree_add_12_51_groupi_n_6412 ,csa_tree_add_12_51_groupi_n_6107 ,csa_tree_add_12_51_groupi_n_6294);
  and csa_tree_add_12_51_groupi_g15350__1617(csa_tree_add_12_51_groupi_n_6411 ,csa_tree_add_12_51_groupi_n_6297 ,csa_tree_add_12_51_groupi_n_6289);
  nor csa_tree_add_12_51_groupi_g15351__2802(csa_tree_add_12_51_groupi_n_6410 ,csa_tree_add_12_51_groupi_n_6297 ,csa_tree_add_12_51_groupi_n_6289);
  nor csa_tree_add_12_51_groupi_g15352__1705(csa_tree_add_12_51_groupi_n_6409 ,csa_tree_add_12_51_groupi_n_6245 ,csa_tree_add_12_51_groupi_n_6308);
  and csa_tree_add_12_51_groupi_g15353__5122(csa_tree_add_12_51_groupi_n_6408 ,csa_tree_add_12_51_groupi_n_6245 ,csa_tree_add_12_51_groupi_n_6308);
  nor csa_tree_add_12_51_groupi_g15354__8246(csa_tree_add_12_51_groupi_n_6407 ,csa_tree_add_12_51_groupi_n_6107 ,csa_tree_add_12_51_groupi_n_6294);
  or csa_tree_add_12_51_groupi_g15355__7098(csa_tree_add_12_51_groupi_n_6406 ,csa_tree_add_12_51_groupi_n_5027 ,csa_tree_add_12_51_groupi_n_6368);
  nor csa_tree_add_12_51_groupi_g15356__6131(csa_tree_add_12_51_groupi_n_6405 ,csa_tree_add_12_51_groupi_n_5028 ,csa_tree_add_12_51_groupi_n_6367);
  nor csa_tree_add_12_51_groupi_g15357__1881(csa_tree_add_12_51_groupi_n_6404 ,csa_tree_add_12_51_groupi_n_6172 ,csa_tree_add_12_51_groupi_n_6348);
  nor csa_tree_add_12_51_groupi_g15358__5115(csa_tree_add_12_51_groupi_n_6403 ,csa_tree_add_12_51_groupi_n_3476 ,csa_tree_add_12_51_groupi_n_6275);
  nor csa_tree_add_12_51_groupi_g15359__7482(csa_tree_add_12_51_groupi_n_6402 ,csa_tree_add_12_51_groupi_n_3475 ,csa_tree_add_12_51_groupi_n_6273);
  nor csa_tree_add_12_51_groupi_g15360__4733(csa_tree_add_12_51_groupi_n_6401 ,csa_tree_add_12_51_groupi_n_3479 ,csa_tree_add_12_51_groupi_n_6274);
  or csa_tree_add_12_51_groupi_g15361__6161(csa_tree_add_12_51_groupi_n_6431 ,csa_tree_add_12_51_groupi_n_6227 ,csa_tree_add_12_51_groupi_n_6354);
  and csa_tree_add_12_51_groupi_g15362__9315(csa_tree_add_12_51_groupi_n_6430 ,csa_tree_add_12_51_groupi_n_6230 ,csa_tree_add_12_51_groupi_n_6365);
  and csa_tree_add_12_51_groupi_g15363__9945(csa_tree_add_12_51_groupi_n_6429 ,csa_tree_add_12_51_groupi_n_6233 ,csa_tree_add_12_51_groupi_n_6346);
  or csa_tree_add_12_51_groupi_g15364__2883(csa_tree_add_12_51_groupi_n_6428 ,csa_tree_add_12_51_groupi_n_6235 ,csa_tree_add_12_51_groupi_n_6350);
  and csa_tree_add_12_51_groupi_g15365__2346(csa_tree_add_12_51_groupi_n_6427 ,csa_tree_add_12_51_groupi_n_6239 ,csa_tree_add_12_51_groupi_n_6352);
  or csa_tree_add_12_51_groupi_g15366__1666(csa_tree_add_12_51_groupi_n_6426 ,csa_tree_add_12_51_groupi_n_6242 ,csa_tree_add_12_51_groupi_n_6358);
  and csa_tree_add_12_51_groupi_g15367__7410(csa_tree_add_12_51_groupi_n_6424 ,csa_tree_add_12_51_groupi_n_6351 ,csa_tree_add_12_51_groupi_n_6236);
  or csa_tree_add_12_51_groupi_g15368__6417(csa_tree_add_12_51_groupi_n_6423 ,csa_tree_add_12_51_groupi_n_6347 ,csa_tree_add_12_51_groupi_n_6244);
  not csa_tree_add_12_51_groupi_g15369(csa_tree_add_12_51_groupi_n_6396 ,csa_tree_add_12_51_groupi_n_6397);
  not csa_tree_add_12_51_groupi_g15370(csa_tree_add_12_51_groupi_n_6393 ,csa_tree_add_12_51_groupi_n_6394);
  and csa_tree_add_12_51_groupi_g15371__5477(csa_tree_add_12_51_groupi_n_6392 ,csa_tree_add_12_51_groupi_n_6313 ,csa_tree_add_12_51_groupi_n_6186);
  nor csa_tree_add_12_51_groupi_g15372__2398(csa_tree_add_12_51_groupi_n_6391 ,csa_tree_add_12_51_groupi_n_6170 ,csa_tree_add_12_51_groupi_n_6366);
  and csa_tree_add_12_51_groupi_g15373__5107(csa_tree_add_12_51_groupi_n_6390 ,csa_tree_add_12_51_groupi_n_6063 ,csa_tree_add_12_51_groupi_n_6303);
  nor csa_tree_add_12_51_groupi_g15374__6260(csa_tree_add_12_51_groupi_n_6389 ,csa_tree_add_12_51_groupi_n_6063 ,csa_tree_add_12_51_groupi_n_6303);
  and csa_tree_add_12_51_groupi_g15375__4319(csa_tree_add_12_51_groupi_n_6388 ,csa_tree_add_12_51_groupi_n_6169 ,csa_tree_add_12_51_groupi_n_6301);
  or csa_tree_add_12_51_groupi_g15376__8428(csa_tree_add_12_51_groupi_n_6387 ,csa_tree_add_12_51_groupi_n_6169 ,csa_tree_add_12_51_groupi_n_6301);
  nor csa_tree_add_12_51_groupi_g15377__5526(csa_tree_add_12_51_groupi_n_6386 ,csa_tree_add_12_51_groupi_n_6256 ,csa_tree_add_12_51_groupi_n_6359);
  nor csa_tree_add_12_51_groupi_g15378__6783(csa_tree_add_12_51_groupi_n_6385 ,csa_tree_add_12_51_groupi_n_4074 ,csa_tree_add_12_51_groupi_n_6286);
  nor csa_tree_add_12_51_groupi_g15379__3680(csa_tree_add_12_51_groupi_n_6384 ,csa_tree_add_12_51_groupi_n_4083 ,csa_tree_add_12_51_groupi_n_6271);
  nor csa_tree_add_12_51_groupi_g15380__1617(csa_tree_add_12_51_groupi_n_6383 ,csa_tree_add_12_51_groupi_n_4080 ,csa_tree_add_12_51_groupi_n_6280);
  nor csa_tree_add_12_51_groupi_g15381__2802(csa_tree_add_12_51_groupi_n_6382 ,csa_tree_add_12_51_groupi_n_4078 ,csa_tree_add_12_51_groupi_n_6285);
  or csa_tree_add_12_51_groupi_g15382__1705(csa_tree_add_12_51_groupi_n_6381 ,csa_tree_add_12_51_groupi_n_4077 ,csa_tree_add_12_51_groupi_n_6284);
  nor csa_tree_add_12_51_groupi_g15383__5122(csa_tree_add_12_51_groupi_n_6380 ,csa_tree_add_12_51_groupi_n_4079 ,csa_tree_add_12_51_groupi_n_6279);
  nor csa_tree_add_12_51_groupi_g15384__8246(csa_tree_add_12_51_groupi_n_6379 ,csa_tree_add_12_51_groupi_n_4076 ,csa_tree_add_12_51_groupi_n_6283);
  or csa_tree_add_12_51_groupi_g15385__7098(csa_tree_add_12_51_groupi_n_6378 ,csa_tree_add_12_51_groupi_n_4072 ,csa_tree_add_12_51_groupi_n_6278);
  xnor csa_tree_add_12_51_groupi_g15386__6131(csa_tree_add_12_51_groupi_n_6377 ,csa_tree_add_12_51_groupi_n_6258 ,csa_tree_add_12_51_groupi_n_6106);
  xnor csa_tree_add_12_51_groupi_g15387__1881(csa_tree_add_12_51_groupi_n_6376 ,csa_tree_add_12_51_groupi_n_6255 ,csa_tree_add_12_51_groupi_n_6061);
  xnor csa_tree_add_12_51_groupi_g15388__5115(csa_tree_add_12_51_groupi_n_6375 ,csa_tree_add_12_51_groupi_n_6247 ,csa_tree_add_12_51_groupi_n_6058);
  nor csa_tree_add_12_51_groupi_g15389__7482(csa_tree_add_12_51_groupi_n_6374 ,csa_tree_add_12_51_groupi_n_4086 ,csa_tree_add_12_51_groupi_n_6277);
  nor csa_tree_add_12_51_groupi_g15390__4733(csa_tree_add_12_51_groupi_n_6373 ,csa_tree_add_12_51_groupi_n_4084 ,csa_tree_add_12_51_groupi_n_6276);
  or csa_tree_add_12_51_groupi_g15391__6161(csa_tree_add_12_51_groupi_n_6372 ,csa_tree_add_12_51_groupi_n_4075 ,csa_tree_add_12_51_groupi_n_6282);
  nor csa_tree_add_12_51_groupi_g15392__9315(csa_tree_add_12_51_groupi_n_6371 ,csa_tree_add_12_51_groupi_n_4085 ,csa_tree_add_12_51_groupi_n_6281);
  xnor csa_tree_add_12_51_groupi_g15393__9945(csa_tree_add_12_51_groupi_n_6370 ,csa_tree_add_12_51_groupi_n_6257 ,csa_tree_add_12_51_groupi_n_6107);
  and csa_tree_add_12_51_groupi_g15395__2883(csa_tree_add_12_51_groupi_n_6400 ,csa_tree_add_12_51_groupi_n_6194 ,csa_tree_add_12_51_groupi_n_6363);
  xnor csa_tree_add_12_51_groupi_g15396__2346(csa_tree_add_12_51_groupi_n_6399 ,csa_tree_add_12_51_groupi_n_6111 ,csa_tree_add_12_51_groupi_n_6176);
  xnor csa_tree_add_12_51_groupi_g15397__1666(csa_tree_add_12_51_groupi_n_6398 ,csa_tree_add_12_51_groupi_n_6115 ,csa_tree_add_12_51_groupi_n_6175);
  and csa_tree_add_12_51_groupi_g15398__7410(csa_tree_add_12_51_groupi_n_6397 ,csa_tree_add_12_51_groupi_n_6364 ,csa_tree_add_12_51_groupi_n_6221);
  or csa_tree_add_12_51_groupi_g15399__6417(csa_tree_add_12_51_groupi_n_6395 ,csa_tree_add_12_51_groupi_n_6224 ,csa_tree_add_12_51_groupi_n_6357);
  xnor csa_tree_add_12_51_groupi_g15400__5477(csa_tree_add_12_51_groupi_n_6394 ,csa_tree_add_12_51_groupi_n_6064 ,csa_tree_add_12_51_groupi_n_6174);
  not csa_tree_add_12_51_groupi_g15401(csa_tree_add_12_51_groupi_n_6367 ,csa_tree_add_12_51_groupi_n_6368);
  and csa_tree_add_12_51_groupi_g15402__2398(csa_tree_add_12_51_groupi_n_6366 ,csa_tree_add_12_51_groupi_n_6091 ,csa_tree_add_12_51_groupi_n_6210);
  or csa_tree_add_12_51_groupi_g15403__5107(csa_tree_add_12_51_groupi_n_6365 ,csa_tree_add_12_51_groupi_n_6125 ,csa_tree_add_12_51_groupi_n_6243);
  or csa_tree_add_12_51_groupi_g15404__6260(csa_tree_add_12_51_groupi_n_6364 ,csa_tree_add_12_51_groupi_n_6213 ,csa_tree_add_12_51_groupi_n_6222);
  or csa_tree_add_12_51_groupi_g15405__4319(csa_tree_add_12_51_groupi_n_6363 ,csa_tree_add_12_51_groupi_n_6066 ,csa_tree_add_12_51_groupi_n_6193);
  and csa_tree_add_12_51_groupi_g15406__8428(csa_tree_add_12_51_groupi_n_6362 ,csa_tree_add_12_51_groupi_n_6058 ,csa_tree_add_12_51_groupi_n_6209);
  or csa_tree_add_12_51_groupi_g15407__5526(csa_tree_add_12_51_groupi_n_6361 ,csa_tree_add_12_51_groupi_n_6058 ,csa_tree_add_12_51_groupi_n_6209);
  nor csa_tree_add_12_51_groupi_g15408__6783(csa_tree_add_12_51_groupi_n_6360 ,csa_tree_add_12_51_groupi_n_6207 ,csa_tree_add_12_51_groupi_n_6062);
  and csa_tree_add_12_51_groupi_g15409__3680(csa_tree_add_12_51_groupi_n_6359 ,csa_tree_add_12_51_groupi_n_6207 ,csa_tree_add_12_51_groupi_n_6062);
  nor csa_tree_add_12_51_groupi_g15410__1617(csa_tree_add_12_51_groupi_n_6358 ,csa_tree_add_12_51_groupi_n_6123 ,csa_tree_add_12_51_groupi_n_6241);
  and csa_tree_add_12_51_groupi_g15411__2802(csa_tree_add_12_51_groupi_n_6357 ,csa_tree_add_12_51_groupi_n_6250 ,csa_tree_add_12_51_groupi_n_6223);
  nor csa_tree_add_12_51_groupi_g15412__1705(csa_tree_add_12_51_groupi_n_6356 ,csa_tree_add_12_51_groupi_n_6106 ,csa_tree_add_12_51_groupi_n_6211);
  and csa_tree_add_12_51_groupi_g15413__5122(csa_tree_add_12_51_groupi_n_6355 ,csa_tree_add_12_51_groupi_n_6106 ,csa_tree_add_12_51_groupi_n_6211);
  and csa_tree_add_12_51_groupi_g15414__8246(csa_tree_add_12_51_groupi_n_6354 ,csa_tree_add_12_51_groupi_n_6122 ,csa_tree_add_12_51_groupi_n_6226);
  nor csa_tree_add_12_51_groupi_g15415__7098(csa_tree_add_12_51_groupi_n_6353 ,csa_tree_add_12_51_groupi_n_6091 ,csa_tree_add_12_51_groupi_n_6210);
  or csa_tree_add_12_51_groupi_g15416__6131(csa_tree_add_12_51_groupi_n_6352 ,csa_tree_add_12_51_groupi_n_6238 ,csa_tree_add_12_51_groupi_n_6173);
  or csa_tree_add_12_51_groupi_g15417__1881(csa_tree_add_12_51_groupi_n_6351 ,csa_tree_add_12_51_groupi_n_6249 ,csa_tree_add_12_51_groupi_n_6237);
  nor csa_tree_add_12_51_groupi_g15418__5115(csa_tree_add_12_51_groupi_n_6350 ,csa_tree_add_12_51_groupi_n_6124 ,csa_tree_add_12_51_groupi_n_6234);
  and csa_tree_add_12_51_groupi_g15419__7482(csa_tree_add_12_51_groupi_n_6349 ,csa_tree_add_12_51_groupi_n_6120 ,csa_tree_add_12_51_groupi_n_6212);
  nor csa_tree_add_12_51_groupi_g15420__4733(csa_tree_add_12_51_groupi_n_6348 ,csa_tree_add_12_51_groupi_n_6120 ,csa_tree_add_12_51_groupi_n_6212);
  and csa_tree_add_12_51_groupi_g15421__6161(csa_tree_add_12_51_groupi_n_6347 ,csa_tree_add_12_51_groupi_n_6231 ,csa_tree_add_12_51_groupi_n_6215);
  or csa_tree_add_12_51_groupi_g15422__9315(csa_tree_add_12_51_groupi_n_6346 ,csa_tree_add_12_51_groupi_n_6067 ,csa_tree_add_12_51_groupi_n_6232);
  or csa_tree_add_12_51_groupi_g15423__9945(csa_tree_add_12_51_groupi_n_6345 ,csa_tree_add_12_51_groupi_n_2877 ,csa_tree_add_12_51_groupi_n_6198);
  nor csa_tree_add_12_51_groupi_g15424__2883(csa_tree_add_12_51_groupi_n_6344 ,csa_tree_add_12_51_groupi_n_3467 ,csa_tree_add_12_51_groupi_n_6199);
  nor csa_tree_add_12_51_groupi_g15425__2346(csa_tree_add_12_51_groupi_n_6343 ,csa_tree_add_12_51_groupi_n_3468 ,csa_tree_add_12_51_groupi_n_6200);
  nor csa_tree_add_12_51_groupi_g15426__1666(csa_tree_add_12_51_groupi_n_6342 ,csa_tree_add_12_51_groupi_n_3453 ,csa_tree_add_12_51_groupi_n_6201);
  nor csa_tree_add_12_51_groupi_g15427__7410(csa_tree_add_12_51_groupi_n_6341 ,csa_tree_add_12_51_groupi_n_3931 ,csa_tree_add_12_51_groupi_n_6203);
  nor csa_tree_add_12_51_groupi_g15428__6417(csa_tree_add_12_51_groupi_n_6340 ,csa_tree_add_12_51_groupi_n_3943 ,csa_tree_add_12_51_groupi_n_6228);
  nor csa_tree_add_12_51_groupi_g15429__5477(csa_tree_add_12_51_groupi_n_6339 ,csa_tree_add_12_51_groupi_n_3937 ,csa_tree_add_12_51_groupi_n_6240);
  nor csa_tree_add_12_51_groupi_g15430__2398(csa_tree_add_12_51_groupi_n_6338 ,csa_tree_add_12_51_groupi_n_3934 ,csa_tree_add_12_51_groupi_n_6204);
  nor csa_tree_add_12_51_groupi_g15431__5107(csa_tree_add_12_51_groupi_n_6337 ,csa_tree_add_12_51_groupi_n_4070 ,csa_tree_add_12_51_groupi_n_6219);
  nor csa_tree_add_12_51_groupi_g15432__6260(csa_tree_add_12_51_groupi_n_6336 ,csa_tree_add_12_51_groupi_n_3936 ,csa_tree_add_12_51_groupi_n_6191);
  nor csa_tree_add_12_51_groupi_g15433__4319(csa_tree_add_12_51_groupi_n_6335 ,csa_tree_add_12_51_groupi_n_3947 ,csa_tree_add_12_51_groupi_n_6216);
  nor csa_tree_add_12_51_groupi_g15434__8428(csa_tree_add_12_51_groupi_n_6334 ,csa_tree_add_12_51_groupi_n_4105 ,csa_tree_add_12_51_groupi_n_6220);
  nor csa_tree_add_12_51_groupi_g15435__5526(csa_tree_add_12_51_groupi_n_6333 ,csa_tree_add_12_51_groupi_n_3930 ,csa_tree_add_12_51_groupi_n_6202);
  nor csa_tree_add_12_51_groupi_g15436__6783(csa_tree_add_12_51_groupi_n_6332 ,csa_tree_add_12_51_groupi_n_3932 ,csa_tree_add_12_51_groupi_n_6195);
  nor csa_tree_add_12_51_groupi_g15437__3680(csa_tree_add_12_51_groupi_n_6331 ,csa_tree_add_12_51_groupi_n_3941 ,csa_tree_add_12_51_groupi_n_6217);
  nor csa_tree_add_12_51_groupi_g15438__1617(csa_tree_add_12_51_groupi_n_6330 ,csa_tree_add_12_51_groupi_n_3939 ,csa_tree_add_12_51_groupi_n_6218);
  or csa_tree_add_12_51_groupi_g15439__2802(csa_tree_add_12_51_groupi_n_6329 ,csa_tree_add_12_51_groupi_n_3752 ,csa_tree_add_12_51_groupi_n_6178);
  or csa_tree_add_12_51_groupi_g15440__1705(csa_tree_add_12_51_groupi_n_6328 ,csa_tree_add_12_51_groupi_n_2875 ,csa_tree_add_12_51_groupi_n_6197);
  or csa_tree_add_12_51_groupi_g15441__5122(csa_tree_add_12_51_groupi_n_6327 ,csa_tree_add_12_51_groupi_n_2878 ,csa_tree_add_12_51_groupi_n_6196);
  or csa_tree_add_12_51_groupi_g15442__8246(csa_tree_add_12_51_groupi_n_6326 ,csa_tree_add_12_51_groupi_n_3754 ,csa_tree_add_12_51_groupi_n_6192);
  or csa_tree_add_12_51_groupi_g15443__7098(csa_tree_add_12_51_groupi_n_6325 ,csa_tree_add_12_51_groupi_n_3749 ,csa_tree_add_12_51_groupi_n_6205);
  or csa_tree_add_12_51_groupi_g15444__6131(csa_tree_add_12_51_groupi_n_6324 ,csa_tree_add_12_51_groupi_n_3750 ,csa_tree_add_12_51_groupi_n_6190);
  or csa_tree_add_12_51_groupi_g15445__1881(csa_tree_add_12_51_groupi_n_6323 ,csa_tree_add_12_51_groupi_n_3746 ,csa_tree_add_12_51_groupi_n_6188);
  or csa_tree_add_12_51_groupi_g15446__5115(csa_tree_add_12_51_groupi_n_6322 ,csa_tree_add_12_51_groupi_n_3739 ,csa_tree_add_12_51_groupi_n_6189);
  or csa_tree_add_12_51_groupi_g15447__7482(csa_tree_add_12_51_groupi_n_6321 ,csa_tree_add_12_51_groupi_n_3757 ,csa_tree_add_12_51_groupi_n_6184);
  or csa_tree_add_12_51_groupi_g15448__4733(csa_tree_add_12_51_groupi_n_6320 ,csa_tree_add_12_51_groupi_n_3738 ,csa_tree_add_12_51_groupi_n_6183);
  or csa_tree_add_12_51_groupi_g15449__6161(csa_tree_add_12_51_groupi_n_6319 ,csa_tree_add_12_51_groupi_n_3759 ,csa_tree_add_12_51_groupi_n_6182);
  or csa_tree_add_12_51_groupi_g15450__9315(csa_tree_add_12_51_groupi_n_6318 ,csa_tree_add_12_51_groupi_n_3747 ,csa_tree_add_12_51_groupi_n_6181);
  or csa_tree_add_12_51_groupi_g15451__9945(csa_tree_add_12_51_groupi_n_6317 ,csa_tree_add_12_51_groupi_n_3761 ,csa_tree_add_12_51_groupi_n_6180);
  or csa_tree_add_12_51_groupi_g15452__2883(csa_tree_add_12_51_groupi_n_6316 ,csa_tree_add_12_51_groupi_n_3748 ,csa_tree_add_12_51_groupi_n_6179);
  and csa_tree_add_12_51_groupi_g15453__2346(csa_tree_add_12_51_groupi_n_6369 ,csa_tree_add_12_51_groupi_n_6146 ,csa_tree_add_12_51_groupi_n_6225);
  or csa_tree_add_12_51_groupi_g15454__1666(csa_tree_add_12_51_groupi_n_6368 ,csa_tree_add_12_51_groupi_n_5033 ,csa_tree_add_12_51_groupi_n_6229);
  not csa_tree_add_12_51_groupi_g15455(csa_tree_add_12_51_groupi_n_6311 ,csa_tree_add_12_51_groupi_n_6310);
  not csa_tree_add_12_51_groupi_g15456(csa_tree_add_12_51_groupi_n_6308 ,csa_tree_add_12_51_groupi_n_6307);
  not csa_tree_add_12_51_groupi_g15457(csa_tree_add_12_51_groupi_n_6305 ,csa_tree_add_12_51_groupi_n_6304);
  not csa_tree_add_12_51_groupi_g15458(csa_tree_add_12_51_groupi_n_6291 ,csa_tree_add_12_51_groupi_n_6290);
  nor csa_tree_add_12_51_groupi_g15459__7410(csa_tree_add_12_51_groupi_n_6286 ,csa_tree_add_12_51_groupi_n_1890 ,csa_tree_add_12_51_groupi_n_989);
  nor csa_tree_add_12_51_groupi_g15460__6417(csa_tree_add_12_51_groupi_n_6285 ,csa_tree_add_12_51_groupi_n_1872 ,csa_tree_add_12_51_groupi_n_992);
  nor csa_tree_add_12_51_groupi_g15461__5477(csa_tree_add_12_51_groupi_n_6284 ,csa_tree_add_12_51_groupi_n_1881 ,csa_tree_add_12_51_groupi_n_179);
  nor csa_tree_add_12_51_groupi_g15462__2398(csa_tree_add_12_51_groupi_n_6283 ,csa_tree_add_12_51_groupi_n_1878 ,csa_tree_add_12_51_groupi_n_989);
  nor csa_tree_add_12_51_groupi_g15463__5107(csa_tree_add_12_51_groupi_n_6282 ,csa_tree_add_12_51_groupi_n_1884 ,csa_tree_add_12_51_groupi_n_990);
  nor csa_tree_add_12_51_groupi_g15464__6260(csa_tree_add_12_51_groupi_n_6281 ,csa_tree_add_12_51_groupi_n_1875 ,csa_tree_add_12_51_groupi_n_993);
  nor csa_tree_add_12_51_groupi_g15465__4319(csa_tree_add_12_51_groupi_n_6280 ,csa_tree_add_12_51_groupi_n_1866 ,csa_tree_add_12_51_groupi_n_960);
  nor csa_tree_add_12_51_groupi_g15466__8428(csa_tree_add_12_51_groupi_n_6279 ,csa_tree_add_12_51_groupi_n_1863 ,csa_tree_add_12_51_groupi_n_959);
  nor csa_tree_add_12_51_groupi_g15467__5526(csa_tree_add_12_51_groupi_n_6278 ,csa_tree_add_12_51_groupi_n_1854 ,csa_tree_add_12_51_groupi_n_990);
  nor csa_tree_add_12_51_groupi_g15468__6783(csa_tree_add_12_51_groupi_n_6277 ,csa_tree_add_12_51_groupi_n_1887 ,csa_tree_add_12_51_groupi_n_959);
  nor csa_tree_add_12_51_groupi_g15469__3680(csa_tree_add_12_51_groupi_n_6276 ,csa_tree_add_12_51_groupi_n_1848 ,csa_tree_add_12_51_groupi_n_993);
  nor csa_tree_add_12_51_groupi_g15470__1617(csa_tree_add_12_51_groupi_n_6275 ,csa_tree_add_12_51_groupi_n_1857 ,csa_tree_add_12_51_groupi_n_992);
  nor csa_tree_add_12_51_groupi_g15471__2802(csa_tree_add_12_51_groupi_n_6274 ,csa_tree_add_12_51_groupi_n_1851 ,csa_tree_add_12_51_groupi_n_1962);
  nor csa_tree_add_12_51_groupi_g15472__1705(csa_tree_add_12_51_groupi_n_6273 ,csa_tree_add_12_51_groupi_n_1860 ,csa_tree_add_12_51_groupi_n_960);
  xnor csa_tree_add_12_51_groupi_g15473__5122(out3[8] ,csa_tree_add_12_51_groupi_n_6171 ,csa_tree_add_12_51_groupi_n_6069);
  nor csa_tree_add_12_51_groupi_g15474__8246(csa_tree_add_12_51_groupi_n_6271 ,csa_tree_add_12_51_groupi_n_1869 ,csa_tree_add_12_51_groupi_n_179);
  xnor csa_tree_add_12_51_groupi_g15475__7098(csa_tree_add_12_51_groupi_n_6270 ,csa_tree_add_12_51_groupi_n_6170 ,csa_tree_add_12_51_groupi_n_6091);
  xnor csa_tree_add_12_51_groupi_g15476__6131(csa_tree_add_12_51_groupi_n_6269 ,csa_tree_add_12_51_groupi_n_6060 ,csa_tree_add_12_51_groupi_n_6101);
  xnor csa_tree_add_12_51_groupi_g15477__1881(csa_tree_add_12_51_groupi_n_6268 ,csa_tree_add_12_51_groupi_n_6097 ,csa_tree_add_12_51_groupi_n_6168);
  xnor csa_tree_add_12_51_groupi_g15478__5115(csa_tree_add_12_51_groupi_n_6267 ,csa_tree_add_12_51_groupi_n_6112 ,csa_tree_add_12_51_groupi_n_5844);
  xnor csa_tree_add_12_51_groupi_g15479__7482(csa_tree_add_12_51_groupi_n_6266 ,csa_tree_add_12_51_groupi_n_6103 ,csa_tree_add_12_51_groupi_n_6173);
  xnor csa_tree_add_12_51_groupi_g15480__4733(csa_tree_add_12_51_groupi_n_6265 ,csa_tree_add_12_51_groupi_n_6113 ,csa_tree_add_12_51_groupi_n_6055);
  xnor csa_tree_add_12_51_groupi_g15481__6161(csa_tree_add_12_51_groupi_n_6264 ,csa_tree_add_12_51_groupi_n_4214 ,csa_tree_add_12_51_groupi_n_6093);
  xor csa_tree_add_12_51_groupi_g15482__9315(csa_tree_add_12_51_groupi_n_6263 ,csa_tree_add_12_51_groupi_n_6120 ,csa_tree_add_12_51_groupi_n_6172);
  xnor csa_tree_add_12_51_groupi_g15483__9945(csa_tree_add_12_51_groupi_n_6262 ,csa_tree_add_12_51_groupi_n_5917 ,csa_tree_add_12_51_groupi_n_6123);
  xnor csa_tree_add_12_51_groupi_g15484__2883(csa_tree_add_12_51_groupi_n_6261 ,csa_tree_add_12_51_groupi_n_6125 ,csa_tree_add_12_51_groupi_n_6117);
  xnor csa_tree_add_12_51_groupi_g15485__2346(csa_tree_add_12_51_groupi_n_6260 ,csa_tree_add_12_51_groupi_n_6095 ,csa_tree_add_12_51_groupi_n_6166);
  xnor csa_tree_add_12_51_groupi_g15486__1666(csa_tree_add_12_51_groupi_n_6259 ,csa_tree_add_12_51_groupi_n_5814 ,csa_tree_add_12_51_groupi_n_6124);
  xnor csa_tree_add_12_51_groupi_g15487__7410(csa_tree_add_12_51_groupi_n_6315 ,csa_tree_add_12_51_groupi_n_6135 ,in3[11]);
  xnor csa_tree_add_12_51_groupi_g15488__6417(csa_tree_add_12_51_groupi_n_6314 ,csa_tree_add_12_51_groupi_n_1930 ,csa_tree_add_12_51_groupi_n_6134);
  or csa_tree_add_12_51_groupi_g15489__5477(csa_tree_add_12_51_groupi_n_6313 ,csa_tree_add_12_51_groupi_n_6002 ,csa_tree_add_12_51_groupi_n_6187);
  xnor csa_tree_add_12_51_groupi_g15490__2398(csa_tree_add_12_51_groupi_n_6312 ,csa_tree_add_12_51_groupi_n_1953 ,csa_tree_add_12_51_groupi_n_6136);
  xnor csa_tree_add_12_51_groupi_g15491__5107(csa_tree_add_12_51_groupi_n_6310 ,csa_tree_add_12_51_groupi_n_6126 ,in2[8]);
  xnor csa_tree_add_12_51_groupi_g15492__6260(csa_tree_add_12_51_groupi_n_6309 ,csa_tree_add_12_51_groupi_n_5909 ,csa_tree_add_12_51_groupi_n_6074);
  xnor csa_tree_add_12_51_groupi_g15493__4319(csa_tree_add_12_51_groupi_n_6307 ,csa_tree_add_12_51_groupi_n_6121 ,csa_tree_add_12_51_groupi_n_5072);
  xnor csa_tree_add_12_51_groupi_g15494__8428(csa_tree_add_12_51_groupi_n_6306 ,csa_tree_add_12_51_groupi_n_5912 ,csa_tree_add_12_51_groupi_n_6077);
  xnor csa_tree_add_12_51_groupi_g15495__5526(csa_tree_add_12_51_groupi_n_6304 ,csa_tree_add_12_51_groupi_n_6133 ,in3[2]);
  xnor csa_tree_add_12_51_groupi_g15496__6783(csa_tree_add_12_51_groupi_n_6303 ,csa_tree_add_12_51_groupi_n_6025 ,csa_tree_add_12_51_groupi_n_6070);
  xnor csa_tree_add_12_51_groupi_g15497__3680(csa_tree_add_12_51_groupi_n_6302 ,csa_tree_add_12_51_groupi_n_5908 ,csa_tree_add_12_51_groupi_n_6071);
  xnor csa_tree_add_12_51_groupi_g15498__1617(csa_tree_add_12_51_groupi_n_6301 ,csa_tree_add_12_51_groupi_n_6028 ,csa_tree_add_12_51_groupi_n_6072);
  xnor csa_tree_add_12_51_groupi_g15499__2802(csa_tree_add_12_51_groupi_n_6300 ,csa_tree_add_12_51_groupi_n_6128 ,in2[11]);
  xnor csa_tree_add_12_51_groupi_g15500__1705(csa_tree_add_12_51_groupi_n_6299 ,csa_tree_add_12_51_groupi_n_5885 ,csa_tree_add_12_51_groupi_n_6076);
  xnor csa_tree_add_12_51_groupi_g15501__5122(csa_tree_add_12_51_groupi_n_6298 ,csa_tree_add_12_51_groupi_n_6137 ,in4[11]);
  xnor csa_tree_add_12_51_groupi_g15502__8246(csa_tree_add_12_51_groupi_n_6297 ,csa_tree_add_12_51_groupi_n_6131 ,in2[5]);
  xnor csa_tree_add_12_51_groupi_g15503__7098(csa_tree_add_12_51_groupi_n_6296 ,csa_tree_add_12_51_groupi_n_6129 ,in4[5]);
  xnor csa_tree_add_12_51_groupi_g15504__6131(csa_tree_add_12_51_groupi_n_6295 ,csa_tree_add_12_51_groupi_n_110 ,csa_tree_add_12_51_groupi_n_6140);
  xnor csa_tree_add_12_51_groupi_g15505__1881(csa_tree_add_12_51_groupi_n_6294 ,csa_tree_add_12_51_groupi_n_6027 ,csa_tree_add_12_51_groupi_n_6073);
  xnor csa_tree_add_12_51_groupi_g15506__5115(csa_tree_add_12_51_groupi_n_6293 ,csa_tree_add_12_51_groupi_n_6138 ,in4[2]);
  xnor csa_tree_add_12_51_groupi_g15507__7482(csa_tree_add_12_51_groupi_n_6292 ,csa_tree_add_12_51_groupi_n_1901 ,csa_tree_add_12_51_groupi_n_6139);
  xnor csa_tree_add_12_51_groupi_g15508__4733(csa_tree_add_12_51_groupi_n_6290 ,csa_tree_add_12_51_groupi_n_6132 ,in2[14]);
  xnor csa_tree_add_12_51_groupi_g15509__6161(csa_tree_add_12_51_groupi_n_6289 ,csa_tree_add_12_51_groupi_n_6130 ,in3[5]);
  xnor csa_tree_add_12_51_groupi_g15510__9315(csa_tree_add_12_51_groupi_n_6288 ,csa_tree_add_12_51_groupi_n_5923 ,csa_tree_add_12_51_groupi_n_6075);
  xnor csa_tree_add_12_51_groupi_g15511__9945(csa_tree_add_12_51_groupi_n_6287 ,csa_tree_add_12_51_groupi_n_1957 ,csa_tree_add_12_51_groupi_n_6127);
  not csa_tree_add_12_51_groupi_g15512(csa_tree_add_12_51_groupi_n_6256 ,csa_tree_add_12_51_groupi_n_6255);
  not csa_tree_add_12_51_groupi_g15513(csa_tree_add_12_51_groupi_n_6249 ,csa_tree_add_12_51_groupi_n_6248);
  and csa_tree_add_12_51_groupi_g15514__2883(csa_tree_add_12_51_groupi_n_6244 ,csa_tree_add_12_51_groupi_n_6113 ,csa_tree_add_12_51_groupi_n_6055);
  nor csa_tree_add_12_51_groupi_g15515__2346(csa_tree_add_12_51_groupi_n_6243 ,csa_tree_add_12_51_groupi_n_6109 ,csa_tree_add_12_51_groupi_n_6116);
  nor csa_tree_add_12_51_groupi_g15516__1666(csa_tree_add_12_51_groupi_n_6242 ,csa_tree_add_12_51_groupi_n_6119 ,csa_tree_add_12_51_groupi_n_5917);
  and csa_tree_add_12_51_groupi_g15517__7410(csa_tree_add_12_51_groupi_n_6241 ,csa_tree_add_12_51_groupi_n_6119 ,csa_tree_add_12_51_groupi_n_5917);
  or csa_tree_add_12_51_groupi_g15518__6417(csa_tree_add_12_51_groupi_n_6240 ,csa_tree_add_12_51_groupi_n_3582 ,csa_tree_add_12_51_groupi_n_6085);
  or csa_tree_add_12_51_groupi_g15519__5477(csa_tree_add_12_51_groupi_n_6239 ,csa_tree_add_12_51_groupi_n_6102 ,csa_tree_add_12_51_groupi_n_6089);
  nor csa_tree_add_12_51_groupi_g15520__2398(csa_tree_add_12_51_groupi_n_6238 ,csa_tree_add_12_51_groupi_n_6103 ,csa_tree_add_12_51_groupi_n_6090);
  nor csa_tree_add_12_51_groupi_g15521__5107(csa_tree_add_12_51_groupi_n_6237 ,csa_tree_add_12_51_groupi_n_6095 ,csa_tree_add_12_51_groupi_n_6166);
  or csa_tree_add_12_51_groupi_g15522__6260(csa_tree_add_12_51_groupi_n_6236 ,csa_tree_add_12_51_groupi_n_6094 ,csa_tree_add_12_51_groupi_n_6165);
  nor csa_tree_add_12_51_groupi_g15523__4319(csa_tree_add_12_51_groupi_n_6235 ,csa_tree_add_12_51_groupi_n_6105 ,csa_tree_add_12_51_groupi_n_5814);
  and csa_tree_add_12_51_groupi_g15524__8428(csa_tree_add_12_51_groupi_n_6234 ,csa_tree_add_12_51_groupi_n_6105 ,csa_tree_add_12_51_groupi_n_5814);
  or csa_tree_add_12_51_groupi_g15525__5526(csa_tree_add_12_51_groupi_n_6233 ,csa_tree_add_12_51_groupi_n_5916 ,csa_tree_add_12_51_groupi_n_6114);
  nor csa_tree_add_12_51_groupi_g15526__6783(csa_tree_add_12_51_groupi_n_6232 ,csa_tree_add_12_51_groupi_n_5915 ,csa_tree_add_12_51_groupi_n_6115);
  or csa_tree_add_12_51_groupi_g15527__3680(csa_tree_add_12_51_groupi_n_6231 ,csa_tree_add_12_51_groupi_n_6113 ,csa_tree_add_12_51_groupi_n_6055);
  or csa_tree_add_12_51_groupi_g15528__1617(csa_tree_add_12_51_groupi_n_6230 ,csa_tree_add_12_51_groupi_n_6108 ,csa_tree_add_12_51_groupi_n_6117);
  and csa_tree_add_12_51_groupi_g15529__2802(csa_tree_add_12_51_groupi_n_6229 ,csa_tree_add_12_51_groupi_n_6121 ,csa_tree_add_12_51_groupi_n_5032);
  or csa_tree_add_12_51_groupi_g15530__1705(csa_tree_add_12_51_groupi_n_6228 ,csa_tree_add_12_51_groupi_n_3630 ,csa_tree_add_12_51_groupi_n_6086);
  nor csa_tree_add_12_51_groupi_g15531__5122(csa_tree_add_12_51_groupi_n_6227 ,csa_tree_add_12_51_groupi_n_4214 ,csa_tree_add_12_51_groupi_n_6092);
  or csa_tree_add_12_51_groupi_g15532__8246(csa_tree_add_12_51_groupi_n_6226 ,csa_tree_add_12_51_groupi_n_4213 ,csa_tree_add_12_51_groupi_n_6093);
  or csa_tree_add_12_51_groupi_g15533__7098(csa_tree_add_12_51_groupi_n_6225 ,csa_tree_add_12_51_groupi_n_6145 ,csa_tree_add_12_51_groupi_n_6065);
  nor csa_tree_add_12_51_groupi_g15534__6131(csa_tree_add_12_51_groupi_n_6224 ,csa_tree_add_12_51_groupi_n_6096 ,csa_tree_add_12_51_groupi_n_6168);
  or csa_tree_add_12_51_groupi_g15535__1881(csa_tree_add_12_51_groupi_n_6223 ,csa_tree_add_12_51_groupi_n_6097 ,csa_tree_add_12_51_groupi_n_6167);
  nor csa_tree_add_12_51_groupi_g15536__5115(csa_tree_add_12_51_groupi_n_6222 ,csa_tree_add_12_51_groupi_n_6060 ,csa_tree_add_12_51_groupi_n_6100);
  or csa_tree_add_12_51_groupi_g15537__7482(csa_tree_add_12_51_groupi_n_6221 ,csa_tree_add_12_51_groupi_n_6059 ,csa_tree_add_12_51_groupi_n_6101);
  or csa_tree_add_12_51_groupi_g15538__4733(csa_tree_add_12_51_groupi_n_6220 ,csa_tree_add_12_51_groupi_n_3415 ,csa_tree_add_12_51_groupi_n_6083);
  or csa_tree_add_12_51_groupi_g15539__6161(csa_tree_add_12_51_groupi_n_6219 ,csa_tree_add_12_51_groupi_n_3412 ,csa_tree_add_12_51_groupi_n_6082);
  or csa_tree_add_12_51_groupi_g15540__9315(csa_tree_add_12_51_groupi_n_6218 ,csa_tree_add_12_51_groupi_n_3723 ,csa_tree_add_12_51_groupi_n_6157);
  or csa_tree_add_12_51_groupi_g15541__9945(csa_tree_add_12_51_groupi_n_6217 ,csa_tree_add_12_51_groupi_n_3668 ,csa_tree_add_12_51_groupi_n_6078);
  or csa_tree_add_12_51_groupi_g15542__2883(csa_tree_add_12_51_groupi_n_6216 ,csa_tree_add_12_51_groupi_n_3595 ,csa_tree_add_12_51_groupi_n_6087);
  and csa_tree_add_12_51_groupi_g15543__2346(csa_tree_add_12_51_groupi_n_6258 ,csa_tree_add_12_51_groupi_n_6036 ,csa_tree_add_12_51_groupi_n_6160);
  and csa_tree_add_12_51_groupi_g15544__1666(csa_tree_add_12_51_groupi_n_6257 ,csa_tree_add_12_51_groupi_n_6041 ,csa_tree_add_12_51_groupi_n_6154);
  or csa_tree_add_12_51_groupi_g15545__7410(csa_tree_add_12_51_groupi_n_6255 ,csa_tree_add_12_51_groupi_n_6143 ,csa_tree_add_12_51_groupi_n_6022);
  and csa_tree_add_12_51_groupi_g15546__6417(csa_tree_add_12_51_groupi_n_6254 ,csa_tree_add_12_51_groupi_n_6035 ,csa_tree_add_12_51_groupi_n_6151);
  and csa_tree_add_12_51_groupi_g15547__5477(csa_tree_add_12_51_groupi_n_6253 ,csa_tree_add_12_51_groupi_n_6150 ,csa_tree_add_12_51_groupi_n_6031);
  and csa_tree_add_12_51_groupi_g15548__2398(csa_tree_add_12_51_groupi_n_6252 ,csa_tree_add_12_51_groupi_n_6037 ,csa_tree_add_12_51_groupi_n_6153);
  and csa_tree_add_12_51_groupi_g15549__5107(csa_tree_add_12_51_groupi_n_6251 ,csa_tree_add_12_51_groupi_n_6052 ,csa_tree_add_12_51_groupi_n_6159);
  or csa_tree_add_12_51_groupi_g15550__6260(csa_tree_add_12_51_groupi_n_6250 ,csa_tree_add_12_51_groupi_n_6050 ,csa_tree_add_12_51_groupi_n_6158);
  or csa_tree_add_12_51_groupi_g15551__4319(csa_tree_add_12_51_groupi_n_6248 ,csa_tree_add_12_51_groupi_n_6047 ,csa_tree_add_12_51_groupi_n_6156);
  and csa_tree_add_12_51_groupi_g15552__8428(csa_tree_add_12_51_groupi_n_6247 ,csa_tree_add_12_51_groupi_n_6000 ,csa_tree_add_12_51_groupi_n_6144);
  or csa_tree_add_12_51_groupi_g15553__5526(csa_tree_add_12_51_groupi_n_6246 ,csa_tree_add_12_51_groupi_n_6149 ,csa_tree_add_12_51_groupi_n_6029);
  and csa_tree_add_12_51_groupi_g15554__6783(csa_tree_add_12_51_groupi_n_6245 ,csa_tree_add_12_51_groupi_n_6045 ,csa_tree_add_12_51_groupi_n_6155);
  nor csa_tree_add_12_51_groupi_g15555__3680(csa_tree_add_12_51_groupi_n_6205 ,csa_tree_add_12_51_groupi_n_1614 ,csa_tree_add_12_51_groupi_n_2181);
  or csa_tree_add_12_51_groupi_g15556__1617(csa_tree_add_12_51_groupi_n_6204 ,csa_tree_add_12_51_groupi_n_3633 ,csa_tree_add_12_51_groupi_n_6081);
  or csa_tree_add_12_51_groupi_g15557__2802(csa_tree_add_12_51_groupi_n_6203 ,csa_tree_add_12_51_groupi_n_3703 ,csa_tree_add_12_51_groupi_n_6080);
  or csa_tree_add_12_51_groupi_g15558__1705(csa_tree_add_12_51_groupi_n_6202 ,csa_tree_add_12_51_groupi_n_3675 ,csa_tree_add_12_51_groupi_n_6079);
  or csa_tree_add_12_51_groupi_g15559__5122(csa_tree_add_12_51_groupi_n_6201 ,csa_tree_add_12_51_groupi_n_3190 ,csa_tree_add_12_51_groupi_n_6142);
  or csa_tree_add_12_51_groupi_g15560__8246(csa_tree_add_12_51_groupi_n_6200 ,csa_tree_add_12_51_groupi_n_3180 ,csa_tree_add_12_51_groupi_n_6147);
  or csa_tree_add_12_51_groupi_g15561__7098(csa_tree_add_12_51_groupi_n_6199 ,csa_tree_add_12_51_groupi_n_3196 ,csa_tree_add_12_51_groupi_n_6148);
  nor csa_tree_add_12_51_groupi_g15562__6131(csa_tree_add_12_51_groupi_n_6198 ,csa_tree_add_12_51_groupi_n_1581 ,csa_tree_add_12_51_groupi_n_2177);
  nor csa_tree_add_12_51_groupi_g15563__1881(csa_tree_add_12_51_groupi_n_6197 ,csa_tree_add_12_51_groupi_n_1590 ,csa_tree_add_12_51_groupi_n_2183);
  nor csa_tree_add_12_51_groupi_g15564__5115(csa_tree_add_12_51_groupi_n_6196 ,csa_tree_add_12_51_groupi_n_1602 ,csa_tree_add_12_51_groupi_n_2178);
  or csa_tree_add_12_51_groupi_g15565__7482(csa_tree_add_12_51_groupi_n_6195 ,csa_tree_add_12_51_groupi_n_3672 ,csa_tree_add_12_51_groupi_n_6084);
  or csa_tree_add_12_51_groupi_g15566__4733(csa_tree_add_12_51_groupi_n_6194 ,csa_tree_add_12_51_groupi_n_5874 ,csa_tree_add_12_51_groupi_n_6110);
  nor csa_tree_add_12_51_groupi_g15567__6161(csa_tree_add_12_51_groupi_n_6193 ,csa_tree_add_12_51_groupi_n_5873 ,csa_tree_add_12_51_groupi_n_6111);
  nor csa_tree_add_12_51_groupi_g15568__9315(csa_tree_add_12_51_groupi_n_6192 ,csa_tree_add_12_51_groupi_n_1620 ,csa_tree_add_12_51_groupi_n_2183);
  or csa_tree_add_12_51_groupi_g15569__9945(csa_tree_add_12_51_groupi_n_6191 ,csa_tree_add_12_51_groupi_n_3711 ,csa_tree_add_12_51_groupi_n_6088);
  nor csa_tree_add_12_51_groupi_g15570__2883(csa_tree_add_12_51_groupi_n_6190 ,csa_tree_add_12_51_groupi_n_1608 ,csa_tree_add_12_51_groupi_n_2184);
  nor csa_tree_add_12_51_groupi_g15571__2346(csa_tree_add_12_51_groupi_n_6189 ,csa_tree_add_12_51_groupi_n_1689 ,csa_tree_add_12_51_groupi_n_2184);
  nor csa_tree_add_12_51_groupi_g15572__1666(csa_tree_add_12_51_groupi_n_6188 ,csa_tree_add_12_51_groupi_n_1596 ,csa_tree_add_12_51_groupi_n_2180);
  and csa_tree_add_12_51_groupi_g15573__7410(csa_tree_add_12_51_groupi_n_6187 ,csa_tree_add_12_51_groupi_n_6171 ,csa_tree_add_12_51_groupi_n_6001);
  or csa_tree_add_12_51_groupi_g15574__6417(csa_tree_add_12_51_groupi_n_6186 ,csa_tree_add_12_51_groupi_n_6112 ,csa_tree_add_12_51_groupi_n_5844);
  and csa_tree_add_12_51_groupi_g15575__5477(csa_tree_add_12_51_groupi_n_6185 ,csa_tree_add_12_51_groupi_n_6112 ,csa_tree_add_12_51_groupi_n_5844);
  nor csa_tree_add_12_51_groupi_g15576__2398(csa_tree_add_12_51_groupi_n_6184 ,csa_tree_add_12_51_groupi_n_1650 ,csa_tree_add_12_51_groupi_n_2155);
  nor csa_tree_add_12_51_groupi_g15577__5107(csa_tree_add_12_51_groupi_n_6183 ,csa_tree_add_12_51_groupi_n_1632 ,csa_tree_add_12_51_groupi_n_6164);
  nor csa_tree_add_12_51_groupi_g15578__6260(csa_tree_add_12_51_groupi_n_6182 ,csa_tree_add_12_51_groupi_n_1671 ,csa_tree_add_12_51_groupi_n_2177);
  nor csa_tree_add_12_51_groupi_g15579__4319(csa_tree_add_12_51_groupi_n_6181 ,csa_tree_add_12_51_groupi_n_1644 ,csa_tree_add_12_51_groupi_n_2178);
  nor csa_tree_add_12_51_groupi_g15580__8428(csa_tree_add_12_51_groupi_n_6180 ,csa_tree_add_12_51_groupi_n_1638 ,csa_tree_add_12_51_groupi_n_2155);
  nor csa_tree_add_12_51_groupi_g15581__5526(csa_tree_add_12_51_groupi_n_6179 ,csa_tree_add_12_51_groupi_n_1659 ,csa_tree_add_12_51_groupi_n_2181);
  nor csa_tree_add_12_51_groupi_g15582__6783(csa_tree_add_12_51_groupi_n_6178 ,csa_tree_add_12_51_groupi_n_1626 ,csa_tree_add_12_51_groupi_n_2180);
  xnor csa_tree_add_12_51_groupi_g15583__3680(out3[7] ,csa_tree_add_12_51_groupi_n_5884 ,csa_tree_add_12_51_groupi_n_5996);
  xnor csa_tree_add_12_51_groupi_g15584__1617(csa_tree_add_12_51_groupi_n_6176 ,csa_tree_add_12_51_groupi_n_5874 ,csa_tree_add_12_51_groupi_n_6066);
  xnor csa_tree_add_12_51_groupi_g15585__2802(csa_tree_add_12_51_groupi_n_6175 ,csa_tree_add_12_51_groupi_n_6067 ,csa_tree_add_12_51_groupi_n_5916);
  xnor csa_tree_add_12_51_groupi_g15586__1705(csa_tree_add_12_51_groupi_n_6174 ,csa_tree_add_12_51_groupi_n_6057 ,csa_tree_add_12_51_groupi_n_5094);
  xnor csa_tree_add_12_51_groupi_g15587__5122(csa_tree_add_12_51_groupi_n_6215 ,csa_tree_add_12_51_groupi_n_5931 ,csa_tree_add_12_51_groupi_n_5997);
  and csa_tree_add_12_51_groupi_g15588__8246(csa_tree_add_12_51_groupi_n_6214 ,csa_tree_add_12_51_groupi_n_6004 ,csa_tree_add_12_51_groupi_n_6152);
  xnor csa_tree_add_12_51_groupi_g15589__7098(csa_tree_add_12_51_groupi_n_6213 ,csa_tree_add_12_51_groupi_n_5919 ,csa_tree_add_12_51_groupi_n_5993);
  xnor csa_tree_add_12_51_groupi_g15590__6131(csa_tree_add_12_51_groupi_n_6212 ,csa_tree_add_12_51_groupi_n_5933 ,csa_tree_add_12_51_groupi_n_5992);
  xnor csa_tree_add_12_51_groupi_g15591__1881(csa_tree_add_12_51_groupi_n_6211 ,csa_tree_add_12_51_groupi_n_5918 ,csa_tree_add_12_51_groupi_n_5995);
  xnor csa_tree_add_12_51_groupi_g15592__5115(csa_tree_add_12_51_groupi_n_6210 ,csa_tree_add_12_51_groupi_n_4921 ,csa_tree_add_12_51_groupi_n_5998);
  xnor csa_tree_add_12_51_groupi_g15593__7482(csa_tree_add_12_51_groupi_n_6209 ,csa_tree_add_12_51_groupi_n_5946 ,csa_tree_add_12_51_groupi_n_5999);
  xnor csa_tree_add_12_51_groupi_g15594__4733(csa_tree_add_12_51_groupi_n_6208 ,csa_tree_add_12_51_groupi_n_5929 ,csa_tree_add_12_51_groupi_n_5994);
  xnor csa_tree_add_12_51_groupi_g15595__6161(csa_tree_add_12_51_groupi_n_6207 ,csa_tree_add_12_51_groupi_n_5851 ,csa_tree_add_12_51_groupi_n_13);
  or csa_tree_add_12_51_groupi_g15596(csa_tree_add_12_51_groupi_n_6206 ,csa_tree_add_12_51_groupi_n_1904 ,csa_tree_add_12_51_groupi_n_6141);
  not csa_tree_add_12_51_groupi_g15597(csa_tree_add_12_51_groupi_n_6168 ,csa_tree_add_12_51_groupi_n_6167);
  not csa_tree_add_12_51_groupi_g15598(csa_tree_add_12_51_groupi_n_6165 ,csa_tree_add_12_51_groupi_n_6166);
  not csa_tree_add_12_51_groupi_g15599(csa_tree_add_12_51_groupi_n_6164 ,csa_tree_add_12_51_groupi_n_6163);
  not csa_tree_add_12_51_groupi_g15600(csa_tree_add_12_51_groupi_n_6162 ,csa_tree_add_12_51_groupi_n_1904);
  not csa_tree_add_12_51_groupi_g15602(csa_tree_add_12_51_groupi_n_6161 ,csa_tree_add_12_51_groupi_n_6163);
  or csa_tree_add_12_51_groupi_g15603(csa_tree_add_12_51_groupi_n_6160 ,csa_tree_add_12_51_groupi_n_6053 ,csa_tree_add_12_51_groupi_n_5853);
  or csa_tree_add_12_51_groupi_g15604(csa_tree_add_12_51_groupi_n_6159 ,csa_tree_add_12_51_groupi_n_6051 ,csa_tree_add_12_51_groupi_n_5991);
  nor csa_tree_add_12_51_groupi_g15605(csa_tree_add_12_51_groupi_n_6158 ,csa_tree_add_12_51_groupi_n_5947 ,csa_tree_add_12_51_groupi_n_6049);
  nor csa_tree_add_12_51_groupi_g15606(csa_tree_add_12_51_groupi_n_6157 ,csa_tree_add_12_51_groupi_n_1613 ,csa_tree_add_12_51_groupi_n_1013);
  and csa_tree_add_12_51_groupi_g15607(csa_tree_add_12_51_groupi_n_6156 ,csa_tree_add_12_51_groupi_n_6046 ,csa_tree_add_12_51_groupi_n_5885);
  or csa_tree_add_12_51_groupi_g15608(csa_tree_add_12_51_groupi_n_6155 ,csa_tree_add_12_51_groupi_n_5944 ,csa_tree_add_12_51_groupi_n_6044);
  or csa_tree_add_12_51_groupi_g15609(csa_tree_add_12_51_groupi_n_6154 ,csa_tree_add_12_51_groupi_n_5945 ,csa_tree_add_12_51_groupi_n_6040);
  or csa_tree_add_12_51_groupi_g15610(csa_tree_add_12_51_groupi_n_6153 ,csa_tree_add_12_51_groupi_n_6027 ,csa_tree_add_12_51_groupi_n_6038);
  or csa_tree_add_12_51_groupi_g15611(csa_tree_add_12_51_groupi_n_6152 ,csa_tree_add_12_51_groupi_n_6003 ,csa_tree_add_12_51_groupi_n_6026);
  or csa_tree_add_12_51_groupi_g15612(csa_tree_add_12_51_groupi_n_6151 ,csa_tree_add_12_51_groupi_n_5881 ,csa_tree_add_12_51_groupi_n_6034);
  or csa_tree_add_12_51_groupi_g15613(csa_tree_add_12_51_groupi_n_6150 ,csa_tree_add_12_51_groupi_n_6033 ,csa_tree_add_12_51_groupi_n_5886);
  and csa_tree_add_12_51_groupi_g15614(csa_tree_add_12_51_groupi_n_6149 ,csa_tree_add_12_51_groupi_n_6030 ,csa_tree_add_12_51_groupi_n_6028);
  nor csa_tree_add_12_51_groupi_g15615(csa_tree_add_12_51_groupi_n_6148 ,csa_tree_add_12_51_groupi_n_1601 ,csa_tree_add_12_51_groupi_n_1016);
  nor csa_tree_add_12_51_groupi_g15616(csa_tree_add_12_51_groupi_n_6147 ,csa_tree_add_12_51_groupi_n_1589 ,csa_tree_add_12_51_groupi_n_163);
  or csa_tree_add_12_51_groupi_g15617(csa_tree_add_12_51_groupi_n_6146 ,csa_tree_add_12_51_groupi_n_6056 ,csa_tree_add_12_51_groupi_n_5094);
  nor csa_tree_add_12_51_groupi_g15618(csa_tree_add_12_51_groupi_n_6145 ,csa_tree_add_12_51_groupi_n_6057 ,csa_tree_add_12_51_groupi_n_5093);
  or csa_tree_add_12_51_groupi_g15619(csa_tree_add_12_51_groupi_n_6144 ,csa_tree_add_12_51_groupi_n_5889 ,csa_tree_add_12_51_groupi_n_6042);
  nor csa_tree_add_12_51_groupi_g15620(csa_tree_add_12_51_groupi_n_6143 ,csa_tree_add_12_51_groupi_n_6023 ,csa_tree_add_12_51_groupi_n_5883);
  nor csa_tree_add_12_51_groupi_g15621(csa_tree_add_12_51_groupi_n_6142 ,csa_tree_add_12_51_groupi_n_1580 ,csa_tree_add_12_51_groupi_n_1013);
  nor csa_tree_add_12_51_groupi_g15622(csa_tree_add_12_51_groupi_n_6141 ,in1[15] ,csa_tree_add_12_51_groupi_n_6068);
  nor csa_tree_add_12_51_groupi_g15623(csa_tree_add_12_51_groupi_n_6140 ,csa_tree_add_12_51_groupi_n_3466 ,csa_tree_add_12_51_groupi_n_6007);
  nor csa_tree_add_12_51_groupi_g15624(csa_tree_add_12_51_groupi_n_6139 ,csa_tree_add_12_51_groupi_n_3918 ,csa_tree_add_12_51_groupi_n_6016);
  nor csa_tree_add_12_51_groupi_g15625(csa_tree_add_12_51_groupi_n_6138 ,csa_tree_add_12_51_groupi_n_3465 ,csa_tree_add_12_51_groupi_n_6005);
  nor csa_tree_add_12_51_groupi_g15626(csa_tree_add_12_51_groupi_n_6137 ,csa_tree_add_12_51_groupi_n_3842 ,csa_tree_add_12_51_groupi_n_6009);
  nor csa_tree_add_12_51_groupi_g15627(csa_tree_add_12_51_groupi_n_6136 ,csa_tree_add_12_51_groupi_n_3869 ,csa_tree_add_12_51_groupi_n_6011);
  nor csa_tree_add_12_51_groupi_g15628(csa_tree_add_12_51_groupi_n_6135 ,csa_tree_add_12_51_groupi_n_3870 ,csa_tree_add_12_51_groupi_n_6010);
  nor csa_tree_add_12_51_groupi_g15629(csa_tree_add_12_51_groupi_n_6134 ,csa_tree_add_12_51_groupi_n_3855 ,csa_tree_add_12_51_groupi_n_6012);
  nor csa_tree_add_12_51_groupi_g15630(csa_tree_add_12_51_groupi_n_6133 ,csa_tree_add_12_51_groupi_n_3452 ,csa_tree_add_12_51_groupi_n_6006);
  nor csa_tree_add_12_51_groupi_g15631(csa_tree_add_12_51_groupi_n_6132 ,csa_tree_add_12_51_groupi_n_3891 ,csa_tree_add_12_51_groupi_n_6015);
  nor csa_tree_add_12_51_groupi_g15632(csa_tree_add_12_51_groupi_n_6131 ,csa_tree_add_12_51_groupi_n_4042 ,csa_tree_add_12_51_groupi_n_6019);
  nor csa_tree_add_12_51_groupi_g15633(csa_tree_add_12_51_groupi_n_6130 ,csa_tree_add_12_51_groupi_n_4041 ,csa_tree_add_12_51_groupi_n_6020);
  nor csa_tree_add_12_51_groupi_g15634(csa_tree_add_12_51_groupi_n_6129 ,csa_tree_add_12_51_groupi_n_4039 ,csa_tree_add_12_51_groupi_n_6018);
  nor csa_tree_add_12_51_groupi_g15635(csa_tree_add_12_51_groupi_n_6128 ,csa_tree_add_12_51_groupi_n_4061 ,csa_tree_add_12_51_groupi_n_6017);
  nor csa_tree_add_12_51_groupi_g15636(csa_tree_add_12_51_groupi_n_6127 ,csa_tree_add_12_51_groupi_n_3904 ,csa_tree_add_12_51_groupi_n_6014);
  nor csa_tree_add_12_51_groupi_g15637(csa_tree_add_12_51_groupi_n_6126 ,csa_tree_add_12_51_groupi_n_3907 ,csa_tree_add_12_51_groupi_n_6013);
  and csa_tree_add_12_51_groupi_g15638(csa_tree_add_12_51_groupi_n_6173 ,csa_tree_add_12_51_groupi_n_6039 ,csa_tree_add_12_51_groupi_n_5964);
  and csa_tree_add_12_51_groupi_g15639(csa_tree_add_12_51_groupi_n_6172 ,csa_tree_add_12_51_groupi_n_6054 ,csa_tree_add_12_51_groupi_n_5969);
  or csa_tree_add_12_51_groupi_g15640(csa_tree_add_12_51_groupi_n_6171 ,csa_tree_add_12_51_groupi_n_5966 ,csa_tree_add_12_51_groupi_n_6032);
  and csa_tree_add_12_51_groupi_g15641(csa_tree_add_12_51_groupi_n_6170 ,csa_tree_add_12_51_groupi_n_5867 ,csa_tree_add_12_51_groupi_n_6008);
  or csa_tree_add_12_51_groupi_g15642(csa_tree_add_12_51_groupi_n_6169 ,csa_tree_add_12_51_groupi_n_5869 ,csa_tree_add_12_51_groupi_n_6048);
  or csa_tree_add_12_51_groupi_g15643(csa_tree_add_12_51_groupi_n_6167 ,csa_tree_add_12_51_groupi_n_6021 ,csa_tree_add_12_51_groupi_n_5980);
  or csa_tree_add_12_51_groupi_g15644(csa_tree_add_12_51_groupi_n_6166 ,csa_tree_add_12_51_groupi_n_5973 ,csa_tree_add_12_51_groupi_n_6043);
  and csa_tree_add_12_51_groupi_g15645(csa_tree_add_12_51_groupi_n_6163 ,in1[15] ,csa_tree_add_12_51_groupi_n_6068);
  not csa_tree_add_12_51_groupi_g15646(csa_tree_add_12_51_groupi_n_6119 ,csa_tree_add_12_51_groupi_n_6118);
  not csa_tree_add_12_51_groupi_g15647(csa_tree_add_12_51_groupi_n_6117 ,csa_tree_add_12_51_groupi_n_6116);
  not csa_tree_add_12_51_groupi_g15648(csa_tree_add_12_51_groupi_n_6114 ,csa_tree_add_12_51_groupi_n_6115);
  not csa_tree_add_12_51_groupi_g15649(csa_tree_add_12_51_groupi_n_6110 ,csa_tree_add_12_51_groupi_n_6111);
  not csa_tree_add_12_51_groupi_g15650(csa_tree_add_12_51_groupi_n_6108 ,csa_tree_add_12_51_groupi_n_6109);
  not csa_tree_add_12_51_groupi_g15651(csa_tree_add_12_51_groupi_n_6105 ,csa_tree_add_12_51_groupi_n_6104);
  not csa_tree_add_12_51_groupi_g15652(csa_tree_add_12_51_groupi_n_6102 ,csa_tree_add_12_51_groupi_n_6103);
  not csa_tree_add_12_51_groupi_g15653(csa_tree_add_12_51_groupi_n_6100 ,csa_tree_add_12_51_groupi_n_6101);
  not csa_tree_add_12_51_groupi_g15654(csa_tree_add_12_51_groupi_n_6098 ,csa_tree_add_12_51_groupi_n_6099);
  not csa_tree_add_12_51_groupi_g15655(csa_tree_add_12_51_groupi_n_6097 ,csa_tree_add_12_51_groupi_n_6096);
  not csa_tree_add_12_51_groupi_g15656(csa_tree_add_12_51_groupi_n_6094 ,csa_tree_add_12_51_groupi_n_6095);
  not csa_tree_add_12_51_groupi_g15657(csa_tree_add_12_51_groupi_n_6093 ,csa_tree_add_12_51_groupi_n_6092);
  not csa_tree_add_12_51_groupi_g15658(csa_tree_add_12_51_groupi_n_6089 ,csa_tree_add_12_51_groupi_n_6090);
  nor csa_tree_add_12_51_groupi_g15659(csa_tree_add_12_51_groupi_n_6088 ,csa_tree_add_12_51_groupi_n_1649 ,csa_tree_add_12_51_groupi_n_1014);
  nor csa_tree_add_12_51_groupi_g15660(csa_tree_add_12_51_groupi_n_6087 ,csa_tree_add_12_51_groupi_n_1619 ,csa_tree_add_12_51_groupi_n_1017);
  nor csa_tree_add_12_51_groupi_g15661(csa_tree_add_12_51_groupi_n_6086 ,csa_tree_add_12_51_groupi_n_1607 ,csa_tree_add_12_51_groupi_n_861);
  nor csa_tree_add_12_51_groupi_g15662(csa_tree_add_12_51_groupi_n_6085 ,csa_tree_add_12_51_groupi_n_1637 ,csa_tree_add_12_51_groupi_n_860);
  nor csa_tree_add_12_51_groupi_g15663(csa_tree_add_12_51_groupi_n_6084 ,csa_tree_add_12_51_groupi_n_1643 ,csa_tree_add_12_51_groupi_n_1014);
  nor csa_tree_add_12_51_groupi_g15664(csa_tree_add_12_51_groupi_n_6083 ,csa_tree_add_12_51_groupi_n_1595 ,csa_tree_add_12_51_groupi_n_860);
  nor csa_tree_add_12_51_groupi_g15665(csa_tree_add_12_51_groupi_n_6082 ,csa_tree_add_12_51_groupi_n_1631 ,csa_tree_add_12_51_groupi_n_1017);
  nor csa_tree_add_12_51_groupi_g15666(csa_tree_add_12_51_groupi_n_6081 ,csa_tree_add_12_51_groupi_n_1670 ,csa_tree_add_12_51_groupi_n_1016);
  nor csa_tree_add_12_51_groupi_g15667(csa_tree_add_12_51_groupi_n_6080 ,csa_tree_add_12_51_groupi_n_1658 ,csa_tree_add_12_51_groupi_n_2001);
  nor csa_tree_add_12_51_groupi_g15668(csa_tree_add_12_51_groupi_n_6079 ,csa_tree_add_12_51_groupi_n_1625 ,csa_tree_add_12_51_groupi_n_861);
  nor csa_tree_add_12_51_groupi_g15669(csa_tree_add_12_51_groupi_n_6078 ,csa_tree_add_12_51_groupi_n_1688 ,csa_tree_add_12_51_groupi_n_163);
  xnor csa_tree_add_12_51_groupi_g15670(csa_tree_add_12_51_groupi_n_6077 ,csa_tree_add_12_51_groupi_n_5944 ,csa_tree_add_12_51_groupi_n_5914);
  xnor csa_tree_add_12_51_groupi_g15671(csa_tree_add_12_51_groupi_n_6076 ,csa_tree_add_12_51_groupi_n_5920 ,csa_tree_add_12_51_groupi_n_5921);
  xnor csa_tree_add_12_51_groupi_g15672(csa_tree_add_12_51_groupi_n_6075 ,csa_tree_add_12_51_groupi_n_5945 ,csa_tree_add_12_51_groupi_n_5925);
  xnor csa_tree_add_12_51_groupi_g15673(csa_tree_add_12_51_groupi_n_6074 ,csa_tree_add_12_51_groupi_n_5947 ,csa_tree_add_12_51_groupi_n_5940);
  xnor csa_tree_add_12_51_groupi_g15674(csa_tree_add_12_51_groupi_n_6073 ,csa_tree_add_12_51_groupi_n_5935 ,csa_tree_add_12_51_groupi_n_5876);
  xnor csa_tree_add_12_51_groupi_g15675(csa_tree_add_12_51_groupi_n_6072 ,csa_tree_add_12_51_groupi_n_5927 ,csa_tree_add_12_51_groupi_n_5880);
  xnor csa_tree_add_12_51_groupi_g15676(csa_tree_add_12_51_groupi_n_6071 ,csa_tree_add_12_51_groupi_n_5991 ,csa_tree_add_12_51_groupi_n_5939);
  xnor csa_tree_add_12_51_groupi_g15677(csa_tree_add_12_51_groupi_n_6070 ,csa_tree_add_12_51_groupi_n_5846 ,csa_tree_add_12_51_groupi_n_5937);
  xnor csa_tree_add_12_51_groupi_g15678(csa_tree_add_12_51_groupi_n_6069 ,csa_tree_add_12_51_groupi_n_5843 ,csa_tree_add_12_51_groupi_n_5926);
  xnor csa_tree_add_12_51_groupi_g15679(csa_tree_add_12_51_groupi_n_6125 ,csa_tree_add_12_51_groupi_n_106 ,csa_tree_add_12_51_groupi_n_5953);
  xnor csa_tree_add_12_51_groupi_g15680(csa_tree_add_12_51_groupi_n_6124 ,csa_tree_add_12_51_groupi_n_1920 ,csa_tree_add_12_51_groupi_n_5958);
  xnor csa_tree_add_12_51_groupi_g15681(csa_tree_add_12_51_groupi_n_6123 ,csa_tree_add_12_51_groupi_n_115 ,csa_tree_add_12_51_groupi_n_5962);
  xnor csa_tree_add_12_51_groupi_g15682(csa_tree_add_12_51_groupi_n_6122 ,csa_tree_add_12_51_groupi_n_5952 ,in2[14]);
  xnor csa_tree_add_12_51_groupi_g15683(csa_tree_add_12_51_groupi_n_6121 ,csa_tree_add_12_51_groupi_n_5949 ,in3[14]);
  xnor csa_tree_add_12_51_groupi_g15684(csa_tree_add_12_51_groupi_n_6120 ,csa_tree_add_12_51_groupi_n_5743 ,csa_tree_add_12_51_groupi_n_5896);
  xnor csa_tree_add_12_51_groupi_g15685(csa_tree_add_12_51_groupi_n_6118 ,csa_tree_add_12_51_groupi_n_5948 ,in4[8]);
  xnor csa_tree_add_12_51_groupi_g15686(csa_tree_add_12_51_groupi_n_6116 ,csa_tree_add_12_51_groupi_n_5961 ,in2[2]);
  xnor csa_tree_add_12_51_groupi_g15687(csa_tree_add_12_51_groupi_n_6115 ,csa_tree_add_12_51_groupi_n_5854 ,csa_tree_add_12_51_groupi_n_5893);
  xnor csa_tree_add_12_51_groupi_g15688(csa_tree_add_12_51_groupi_n_6113 ,csa_tree_add_12_51_groupi_n_5752 ,csa_tree_add_12_51_groupi_n_5894);
  xnor csa_tree_add_12_51_groupi_g15689(csa_tree_add_12_51_groupi_n_6112 ,csa_tree_add_12_51_groupi_n_5943 ,csa_tree_add_12_51_groupi_n_5898);
  xnor csa_tree_add_12_51_groupi_g15690(csa_tree_add_12_51_groupi_n_6111 ,csa_tree_add_12_51_groupi_n_5850 ,csa_tree_add_12_51_groupi_n_5895);
  xnor csa_tree_add_12_51_groupi_g15691(csa_tree_add_12_51_groupi_n_6109 ,csa_tree_add_12_51_groupi_n_5960 ,in4[2]);
  xnor csa_tree_add_12_51_groupi_g15692(csa_tree_add_12_51_groupi_n_6107 ,csa_tree_add_12_51_groupi_n_1933 ,csa_tree_add_12_51_groupi_n_5959);
  xnor csa_tree_add_12_51_groupi_g15693(csa_tree_add_12_51_groupi_n_6106 ,csa_tree_add_12_51_groupi_n_5746 ,csa_tree_add_12_51_groupi_n_5897);
  xnor csa_tree_add_12_51_groupi_g15694(csa_tree_add_12_51_groupi_n_6104 ,csa_tree_add_12_51_groupi_n_5957 ,in4[11]);
  xnor csa_tree_add_12_51_groupi_g15695(csa_tree_add_12_51_groupi_n_6103 ,csa_tree_add_12_51_groupi_n_5955 ,in2[5]);
  xnor csa_tree_add_12_51_groupi_g15696(csa_tree_add_12_51_groupi_n_6101 ,csa_tree_add_12_51_groupi_n_5761 ,csa_tree_add_12_51_groupi_n_5891);
  xnor csa_tree_add_12_51_groupi_g15697(csa_tree_add_12_51_groupi_n_6099 ,csa_tree_add_12_51_groupi_n_5941 ,csa_tree_add_12_51_groupi_n_5890);
  xnor csa_tree_add_12_51_groupi_g15698(csa_tree_add_12_51_groupi_n_6096 ,csa_tree_add_12_51_groupi_n_96 ,csa_tree_add_12_51_groupi_n_5950);
  xnor csa_tree_add_12_51_groupi_g15699(csa_tree_add_12_51_groupi_n_6095 ,csa_tree_add_12_51_groupi_n_5954 ,in3[11]);
  xnor csa_tree_add_12_51_groupi_g15700(csa_tree_add_12_51_groupi_n_6092 ,csa_tree_add_12_51_groupi_n_1901 ,csa_tree_add_12_51_groupi_n_5951);
  xnor csa_tree_add_12_51_groupi_g15701(csa_tree_add_12_51_groupi_n_6091 ,csa_tree_add_12_51_groupi_n_5739 ,csa_tree_add_12_51_groupi_n_5892);
  xnor csa_tree_add_12_51_groupi_g15702(csa_tree_add_12_51_groupi_n_6090 ,csa_tree_add_12_51_groupi_n_5956 ,in3[5]);
  not csa_tree_add_12_51_groupi_g15703(csa_tree_add_12_51_groupi_n_6065 ,csa_tree_add_12_51_groupi_n_6064);
  not csa_tree_add_12_51_groupi_g15705(csa_tree_add_12_51_groupi_n_6062 ,csa_tree_add_12_51_groupi_n_6061);
  not csa_tree_add_12_51_groupi_g15706(csa_tree_add_12_51_groupi_n_6059 ,csa_tree_add_12_51_groupi_n_6060);
  not csa_tree_add_12_51_groupi_g15707(csa_tree_add_12_51_groupi_n_6056 ,csa_tree_add_12_51_groupi_n_6057);
  or csa_tree_add_12_51_groupi_g15708(csa_tree_add_12_51_groupi_n_6054 ,csa_tree_add_12_51_groupi_n_5970 ,csa_tree_add_12_51_groupi_n_5716);
  nor csa_tree_add_12_51_groupi_g15709(csa_tree_add_12_51_groupi_n_6053 ,csa_tree_add_12_51_groupi_n_5707 ,csa_tree_add_12_51_groupi_n_5929);
  or csa_tree_add_12_51_groupi_g15710(csa_tree_add_12_51_groupi_n_6052 ,csa_tree_add_12_51_groupi_n_5939 ,csa_tree_add_12_51_groupi_n_5907);
  nor csa_tree_add_12_51_groupi_g15711(csa_tree_add_12_51_groupi_n_6051 ,csa_tree_add_12_51_groupi_n_5938 ,csa_tree_add_12_51_groupi_n_5908);
  nor csa_tree_add_12_51_groupi_g15712(csa_tree_add_12_51_groupi_n_6050 ,csa_tree_add_12_51_groupi_n_5940 ,csa_tree_add_12_51_groupi_n_5910);
  and csa_tree_add_12_51_groupi_g15713(csa_tree_add_12_51_groupi_n_6049 ,csa_tree_add_12_51_groupi_n_5940 ,csa_tree_add_12_51_groupi_n_5910);
  and csa_tree_add_12_51_groupi_g15714(csa_tree_add_12_51_groupi_n_6048 ,csa_tree_add_12_51_groupi_n_5868 ,csa_tree_add_12_51_groupi_n_5943);
  and csa_tree_add_12_51_groupi_g15715(csa_tree_add_12_51_groupi_n_6047 ,csa_tree_add_12_51_groupi_n_5920 ,csa_tree_add_12_51_groupi_n_5921);
  or csa_tree_add_12_51_groupi_g15716(csa_tree_add_12_51_groupi_n_6046 ,csa_tree_add_12_51_groupi_n_5920 ,csa_tree_add_12_51_groupi_n_5921);
  or csa_tree_add_12_51_groupi_g15717(csa_tree_add_12_51_groupi_n_6045 ,csa_tree_add_12_51_groupi_n_5911 ,csa_tree_add_12_51_groupi_n_5914);
  nor csa_tree_add_12_51_groupi_g15718(csa_tree_add_12_51_groupi_n_6044 ,csa_tree_add_12_51_groupi_n_5912 ,csa_tree_add_12_51_groupi_n_5913);
  and csa_tree_add_12_51_groupi_g15719(csa_tree_add_12_51_groupi_n_6043 ,csa_tree_add_12_51_groupi_n_5946 ,csa_tree_add_12_51_groupi_n_5974);
  and csa_tree_add_12_51_groupi_g15720(csa_tree_add_12_51_groupi_n_6042 ,csa_tree_add_12_51_groupi_n_5877 ,csa_tree_add_12_51_groupi_n_5918);
  or csa_tree_add_12_51_groupi_g15721(csa_tree_add_12_51_groupi_n_6041 ,csa_tree_add_12_51_groupi_n_5922 ,csa_tree_add_12_51_groupi_n_5925);
  nor csa_tree_add_12_51_groupi_g15722(csa_tree_add_12_51_groupi_n_6040 ,csa_tree_add_12_51_groupi_n_5923 ,csa_tree_add_12_51_groupi_n_5924);
  or csa_tree_add_12_51_groupi_g15723(csa_tree_add_12_51_groupi_n_6039 ,csa_tree_add_12_51_groupi_n_5815 ,csa_tree_add_12_51_groupi_n_5965);
  nor csa_tree_add_12_51_groupi_g15724(csa_tree_add_12_51_groupi_n_6038 ,csa_tree_add_12_51_groupi_n_5935 ,csa_tree_add_12_51_groupi_n_5876);
  or csa_tree_add_12_51_groupi_g15725(csa_tree_add_12_51_groupi_n_6037 ,csa_tree_add_12_51_groupi_n_5934 ,csa_tree_add_12_51_groupi_n_5875);
  or csa_tree_add_12_51_groupi_g15726(csa_tree_add_12_51_groupi_n_6036 ,csa_tree_add_12_51_groupi_n_5708 ,csa_tree_add_12_51_groupi_n_5928);
  or csa_tree_add_12_51_groupi_g15727(csa_tree_add_12_51_groupi_n_6035 ,csa_tree_add_12_51_groupi_n_5750 ,csa_tree_add_12_51_groupi_n_5932);
  nor csa_tree_add_12_51_groupi_g15728(csa_tree_add_12_51_groupi_n_6034 ,csa_tree_add_12_51_groupi_n_5749 ,csa_tree_add_12_51_groupi_n_5933);
  nor csa_tree_add_12_51_groupi_g15729(csa_tree_add_12_51_groupi_n_6033 ,csa_tree_add_12_51_groupi_n_5753 ,csa_tree_add_12_51_groupi_n_5931);
  and csa_tree_add_12_51_groupi_g15730(csa_tree_add_12_51_groupi_n_6032 ,csa_tree_add_12_51_groupi_n_5884 ,csa_tree_add_12_51_groupi_n_5967);
  or csa_tree_add_12_51_groupi_g15731(csa_tree_add_12_51_groupi_n_6031 ,csa_tree_add_12_51_groupi_n_5754 ,csa_tree_add_12_51_groupi_n_5930);
  or csa_tree_add_12_51_groupi_g15732(csa_tree_add_12_51_groupi_n_6030 ,csa_tree_add_12_51_groupi_n_5927 ,csa_tree_add_12_51_groupi_n_5880);
  and csa_tree_add_12_51_groupi_g15733(csa_tree_add_12_51_groupi_n_6029 ,csa_tree_add_12_51_groupi_n_5927 ,csa_tree_add_12_51_groupi_n_5880);
  or csa_tree_add_12_51_groupi_g15734(csa_tree_add_12_51_groupi_n_6068 ,csa_tree_add_12_51_groupi_n_2441 ,csa_tree_add_12_51_groupi_n_5979);
  and csa_tree_add_12_51_groupi_g15735(csa_tree_add_12_51_groupi_n_6067 ,csa_tree_add_12_51_groupi_n_5856 ,csa_tree_add_12_51_groupi_n_5968);
  and csa_tree_add_12_51_groupi_g15736(csa_tree_add_12_51_groupi_n_6066 ,csa_tree_add_12_51_groupi_n_5864 ,csa_tree_add_12_51_groupi_n_5976);
  or csa_tree_add_12_51_groupi_g15737(csa_tree_add_12_51_groupi_n_6064 ,csa_tree_add_12_51_groupi_n_5871 ,csa_tree_add_12_51_groupi_n_5972);
  or csa_tree_add_12_51_groupi_g15738(csa_tree_add_12_51_groupi_n_6063 ,csa_tree_add_12_51_groupi_n_5963 ,csa_tree_add_12_51_groupi_n_5859);
  or csa_tree_add_12_51_groupi_g15739(csa_tree_add_12_51_groupi_n_6061 ,csa_tree_add_12_51_groupi_n_5839 ,csa_tree_add_12_51_groupi_n_5981);
  or csa_tree_add_12_51_groupi_g15740(csa_tree_add_12_51_groupi_n_6060 ,csa_tree_add_12_51_groupi_n_5982 ,csa_tree_add_12_51_groupi_n_5837);
  and csa_tree_add_12_51_groupi_g15741(csa_tree_add_12_51_groupi_n_6058 ,csa_tree_add_12_51_groupi_n_5863 ,csa_tree_add_12_51_groupi_n_5975);
  or csa_tree_add_12_51_groupi_g15742(csa_tree_add_12_51_groupi_n_6057 ,csa_tree_add_12_51_groupi_n_5866 ,csa_tree_add_12_51_groupi_n_5978);
  or csa_tree_add_12_51_groupi_g15743(csa_tree_add_12_51_groupi_n_6055 ,csa_tree_add_12_51_groupi_n_5971 ,csa_tree_add_12_51_groupi_n_5855);
  not csa_tree_add_12_51_groupi_g15744(csa_tree_add_12_51_groupi_n_6026 ,csa_tree_add_12_51_groupi_n_6025);
  and csa_tree_add_12_51_groupi_g15745(csa_tree_add_12_51_groupi_n_6023 ,csa_tree_add_12_51_groupi_n_5760 ,csa_tree_add_12_51_groupi_n_5919);
  nor csa_tree_add_12_51_groupi_g15746(csa_tree_add_12_51_groupi_n_6022 ,csa_tree_add_12_51_groupi_n_5760 ,csa_tree_add_12_51_groupi_n_5919);
  nor csa_tree_add_12_51_groupi_g15747(csa_tree_add_12_51_groupi_n_6021 ,csa_tree_add_12_51_groupi_n_5977 ,csa_tree_add_12_51_groupi_n_5888);
  or csa_tree_add_12_51_groupi_g15748(csa_tree_add_12_51_groupi_n_6020 ,csa_tree_add_12_51_groupi_n_3384 ,csa_tree_add_12_51_groupi_n_5990);
  or csa_tree_add_12_51_groupi_g15749(csa_tree_add_12_51_groupi_n_6019 ,csa_tree_add_12_51_groupi_n_3312 ,csa_tree_add_12_51_groupi_n_5904);
  or csa_tree_add_12_51_groupi_g15750(csa_tree_add_12_51_groupi_n_6018 ,csa_tree_add_12_51_groupi_n_3323 ,csa_tree_add_12_51_groupi_n_5903);
  or csa_tree_add_12_51_groupi_g15751(csa_tree_add_12_51_groupi_n_6017 ,csa_tree_add_12_51_groupi_n_3259 ,csa_tree_add_12_51_groupi_n_5906);
  or csa_tree_add_12_51_groupi_g15752(csa_tree_add_12_51_groupi_n_6016 ,csa_tree_add_12_51_groupi_n_3725 ,csa_tree_add_12_51_groupi_n_5986);
  or csa_tree_add_12_51_groupi_g15753(csa_tree_add_12_51_groupi_n_6015 ,csa_tree_add_12_51_groupi_n_3624 ,csa_tree_add_12_51_groupi_n_5987);
  or csa_tree_add_12_51_groupi_g15754(csa_tree_add_12_51_groupi_n_6014 ,csa_tree_add_12_51_groupi_n_3658 ,csa_tree_add_12_51_groupi_n_5988);
  or csa_tree_add_12_51_groupi_g15755(csa_tree_add_12_51_groupi_n_6013 ,csa_tree_add_12_51_groupi_n_3688 ,csa_tree_add_12_51_groupi_n_5989);
  or csa_tree_add_12_51_groupi_g15756(csa_tree_add_12_51_groupi_n_6012 ,csa_tree_add_12_51_groupi_n_3709 ,csa_tree_add_12_51_groupi_n_5900);
  or csa_tree_add_12_51_groupi_g15757(csa_tree_add_12_51_groupi_n_6011 ,csa_tree_add_12_51_groupi_n_3641 ,csa_tree_add_12_51_groupi_n_5902);
  or csa_tree_add_12_51_groupi_g15758(csa_tree_add_12_51_groupi_n_6010 ,csa_tree_add_12_51_groupi_n_3715 ,csa_tree_add_12_51_groupi_n_5905);
  or csa_tree_add_12_51_groupi_g15759(csa_tree_add_12_51_groupi_n_6009 ,csa_tree_add_12_51_groupi_n_3679 ,csa_tree_add_12_51_groupi_n_5901);
  or csa_tree_add_12_51_groupi_g15760(csa_tree_add_12_51_groupi_n_6008 ,csa_tree_add_12_51_groupi_n_5942 ,csa_tree_add_12_51_groupi_n_5870);
  or csa_tree_add_12_51_groupi_g15761(csa_tree_add_12_51_groupi_n_6007 ,csa_tree_add_12_51_groupi_n_3041 ,csa_tree_add_12_51_groupi_n_5983);
  or csa_tree_add_12_51_groupi_g15762(csa_tree_add_12_51_groupi_n_6006 ,csa_tree_add_12_51_groupi_n_3080 ,csa_tree_add_12_51_groupi_n_5984);
  or csa_tree_add_12_51_groupi_g15763(csa_tree_add_12_51_groupi_n_6005 ,csa_tree_add_12_51_groupi_n_3140 ,csa_tree_add_12_51_groupi_n_5985);
  or csa_tree_add_12_51_groupi_g15764(csa_tree_add_12_51_groupi_n_6004 ,csa_tree_add_12_51_groupi_n_5845 ,csa_tree_add_12_51_groupi_n_5936);
  nor csa_tree_add_12_51_groupi_g15765(csa_tree_add_12_51_groupi_n_6003 ,csa_tree_add_12_51_groupi_n_5846 ,csa_tree_add_12_51_groupi_n_5937);
  and csa_tree_add_12_51_groupi_g15766(csa_tree_add_12_51_groupi_n_6002 ,csa_tree_add_12_51_groupi_n_5843 ,csa_tree_add_12_51_groupi_n_5926);
  or csa_tree_add_12_51_groupi_g15767(csa_tree_add_12_51_groupi_n_6001 ,csa_tree_add_12_51_groupi_n_5843 ,csa_tree_add_12_51_groupi_n_5926);
  or csa_tree_add_12_51_groupi_g15768(csa_tree_add_12_51_groupi_n_6000 ,csa_tree_add_12_51_groupi_n_5877 ,csa_tree_add_12_51_groupi_n_5918);
  xnor csa_tree_add_12_51_groupi_g15769(csa_tree_add_12_51_groupi_n_5999 ,csa_tree_add_12_51_groupi_n_5765 ,csa_tree_add_12_51_groupi_n_5848);
  xnor csa_tree_add_12_51_groupi_g15770(csa_tree_add_12_51_groupi_n_5998 ,csa_tree_add_12_51_groupi_n_5887 ,csa_tree_add_12_51_groupi_n_5812);
  xnor csa_tree_add_12_51_groupi_g15771(csa_tree_add_12_51_groupi_n_5997 ,csa_tree_add_12_51_groupi_n_5886 ,csa_tree_add_12_51_groupi_n_5754);
  xnor csa_tree_add_12_51_groupi_g15773(csa_tree_add_12_51_groupi_n_5996 ,csa_tree_add_12_51_groupi_n_5538 ,csa_tree_add_12_51_groupi_n_5852);
  xnor csa_tree_add_12_51_groupi_g15774(csa_tree_add_12_51_groupi_n_5995 ,csa_tree_add_12_51_groupi_n_5889 ,csa_tree_add_12_51_groupi_n_5877);
  xnor csa_tree_add_12_51_groupi_g15775(csa_tree_add_12_51_groupi_n_5994 ,csa_tree_add_12_51_groupi_n_5853 ,csa_tree_add_12_51_groupi_n_5708);
  xnor csa_tree_add_12_51_groupi_g15776(csa_tree_add_12_51_groupi_n_5993 ,csa_tree_add_12_51_groupi_n_5883 ,csa_tree_add_12_51_groupi_n_5760);
  xnor csa_tree_add_12_51_groupi_g15777(csa_tree_add_12_51_groupi_n_5992 ,csa_tree_add_12_51_groupi_n_5881 ,csa_tree_add_12_51_groupi_n_5750);
  xnor csa_tree_add_12_51_groupi_g15778(csa_tree_add_12_51_groupi_n_6028 ,csa_tree_add_12_51_groupi_n_5766 ,csa_tree_add_12_51_groupi_n_5820);
  xnor csa_tree_add_12_51_groupi_g15779(csa_tree_add_12_51_groupi_n_6027 ,csa_tree_add_12_51_groupi_n_5757 ,csa_tree_add_12_51_groupi_n_5821);
  xnor csa_tree_add_12_51_groupi_g15780(csa_tree_add_12_51_groupi_n_6025 ,csa_tree_add_12_51_groupi_n_5879 ,csa_tree_add_12_51_groupi_n_5819);
  xnor csa_tree_add_12_51_groupi_g15781(csa_tree_add_12_51_groupi_n_6024 ,csa_tree_add_12_51_groupi_n_5882 ,csa_tree_add_12_51_groupi_n_2568);
  nor csa_tree_add_12_51_groupi_g15782(csa_tree_add_12_51_groupi_n_5990 ,csa_tree_add_12_51_groupi_n_1607 ,csa_tree_add_12_51_groupi_n_806);
  nor csa_tree_add_12_51_groupi_g15783(csa_tree_add_12_51_groupi_n_5989 ,csa_tree_add_12_51_groupi_n_1613 ,csa_tree_add_12_51_groupi_n_809);
  nor csa_tree_add_12_51_groupi_g15784(csa_tree_add_12_51_groupi_n_5988 ,csa_tree_add_12_51_groupi_n_1688 ,csa_tree_add_12_51_groupi_n_177);
  nor csa_tree_add_12_51_groupi_g15785(csa_tree_add_12_51_groupi_n_5987 ,csa_tree_add_12_51_groupi_n_1619 ,csa_tree_add_12_51_groupi_n_806);
  nor csa_tree_add_12_51_groupi_g15786(csa_tree_add_12_51_groupi_n_5986 ,csa_tree_add_12_51_groupi_n_1595 ,csa_tree_add_12_51_groupi_n_807);
  nor csa_tree_add_12_51_groupi_g15787(csa_tree_add_12_51_groupi_n_5985 ,csa_tree_add_12_51_groupi_n_1580 ,csa_tree_add_12_51_groupi_n_810);
  nor csa_tree_add_12_51_groupi_g15788(csa_tree_add_12_51_groupi_n_5984 ,csa_tree_add_12_51_groupi_n_1601 ,csa_tree_add_12_51_groupi_n_909);
  nor csa_tree_add_12_51_groupi_g15789(csa_tree_add_12_51_groupi_n_5983 ,csa_tree_add_12_51_groupi_n_1589 ,csa_tree_add_12_51_groupi_n_908);
  nor csa_tree_add_12_51_groupi_g15790(csa_tree_add_12_51_groupi_n_5982 ,csa_tree_add_12_51_groupi_n_5714 ,csa_tree_add_12_51_groupi_n_5838);
  nor csa_tree_add_12_51_groupi_g15791(csa_tree_add_12_51_groupi_n_5981 ,csa_tree_add_12_51_groupi_n_0 ,csa_tree_add_12_51_groupi_n_5840);
  nor csa_tree_add_12_51_groupi_g15792(csa_tree_add_12_51_groupi_n_5980 ,csa_tree_add_12_51_groupi_n_5756 ,csa_tree_add_12_51_groupi_n_5851);
  nor csa_tree_add_12_51_groupi_g15793(csa_tree_add_12_51_groupi_n_5979 ,csa_tree_add_12_51_groupi_n_2440 ,csa_tree_add_12_51_groupi_n_5882);
  nor csa_tree_add_12_51_groupi_g15794(csa_tree_add_12_51_groupi_n_5978 ,csa_tree_add_12_51_groupi_n_5769 ,csa_tree_add_12_51_groupi_n_5865);
  and csa_tree_add_12_51_groupi_g15795(csa_tree_add_12_51_groupi_n_5977 ,csa_tree_add_12_51_groupi_n_5756 ,csa_tree_add_12_51_groupi_n_5851);
  or csa_tree_add_12_51_groupi_g15796(csa_tree_add_12_51_groupi_n_5976 ,csa_tree_add_12_51_groupi_n_5862 ,csa_tree_add_12_51_groupi_n_5818);
  or csa_tree_add_12_51_groupi_g15797(csa_tree_add_12_51_groupi_n_5975 ,csa_tree_add_12_51_groupi_n_5771 ,csa_tree_add_12_51_groupi_n_5861);
  or csa_tree_add_12_51_groupi_g15798(csa_tree_add_12_51_groupi_n_5974 ,csa_tree_add_12_51_groupi_n_5765 ,csa_tree_add_12_51_groupi_n_5847);
  nor csa_tree_add_12_51_groupi_g15799(csa_tree_add_12_51_groupi_n_5973 ,csa_tree_add_12_51_groupi_n_5764 ,csa_tree_add_12_51_groupi_n_5848);
  and csa_tree_add_12_51_groupi_g15800(csa_tree_add_12_51_groupi_n_5972 ,csa_tree_add_12_51_groupi_n_5887 ,csa_tree_add_12_51_groupi_n_5860);
  nor csa_tree_add_12_51_groupi_g15801(csa_tree_add_12_51_groupi_n_5971 ,csa_tree_add_12_51_groupi_n_5712 ,csa_tree_add_12_51_groupi_n_5872);
  nor csa_tree_add_12_51_groupi_g15802(csa_tree_add_12_51_groupi_n_5970 ,csa_tree_add_12_51_groupi_n_5573 ,csa_tree_add_12_51_groupi_n_5879);
  or csa_tree_add_12_51_groupi_g15803(csa_tree_add_12_51_groupi_n_5969 ,csa_tree_add_12_51_groupi_n_5574 ,csa_tree_add_12_51_groupi_n_5878);
  or csa_tree_add_12_51_groupi_g15804(csa_tree_add_12_51_groupi_n_5968 ,csa_tree_add_12_51_groupi_n_5770 ,csa_tree_add_12_51_groupi_n_5857);
  or csa_tree_add_12_51_groupi_g15805(csa_tree_add_12_51_groupi_n_5967 ,csa_tree_add_12_51_groupi_n_5538 ,csa_tree_add_12_51_groupi_n_5852);
  and csa_tree_add_12_51_groupi_g15806(csa_tree_add_12_51_groupi_n_5966 ,csa_tree_add_12_51_groupi_n_5538 ,csa_tree_add_12_51_groupi_n_5852);
  nor csa_tree_add_12_51_groupi_g15807(csa_tree_add_12_51_groupi_n_5965 ,csa_tree_add_12_51_groupi_n_5850 ,csa_tree_add_12_51_groupi_n_5762);
  or csa_tree_add_12_51_groupi_g15808(csa_tree_add_12_51_groupi_n_5964 ,csa_tree_add_12_51_groupi_n_5849 ,csa_tree_add_12_51_groupi_n_5763);
  and csa_tree_add_12_51_groupi_g15809(csa_tree_add_12_51_groupi_n_5963 ,csa_tree_add_12_51_groupi_n_5858 ,csa_tree_add_12_51_groupi_n_5854);
  nor csa_tree_add_12_51_groupi_g15810(csa_tree_add_12_51_groupi_n_5962 ,csa_tree_add_12_51_groupi_n_3902 ,csa_tree_add_12_51_groupi_n_5835);
  nor csa_tree_add_12_51_groupi_g15811(csa_tree_add_12_51_groupi_n_5961 ,csa_tree_add_12_51_groupi_n_3439 ,csa_tree_add_12_51_groupi_n_5823);
  nor csa_tree_add_12_51_groupi_g15812(csa_tree_add_12_51_groupi_n_5960 ,csa_tree_add_12_51_groupi_n_3463 ,csa_tree_add_12_51_groupi_n_5824);
  nor csa_tree_add_12_51_groupi_g15813(csa_tree_add_12_51_groupi_n_5959 ,csa_tree_add_12_51_groupi_n_3853 ,csa_tree_add_12_51_groupi_n_5827);
  nor csa_tree_add_12_51_groupi_g15814(csa_tree_add_12_51_groupi_n_5958 ,csa_tree_add_12_51_groupi_n_3832 ,csa_tree_add_12_51_groupi_n_5841);
  nor csa_tree_add_12_51_groupi_g15815(csa_tree_add_12_51_groupi_n_5957 ,csa_tree_add_12_51_groupi_n_3834 ,csa_tree_add_12_51_groupi_n_5826);
  nor csa_tree_add_12_51_groupi_g15816(csa_tree_add_12_51_groupi_n_5956 ,csa_tree_add_12_51_groupi_n_3893 ,csa_tree_add_12_51_groupi_n_5832);
  nor csa_tree_add_12_51_groupi_g15817(csa_tree_add_12_51_groupi_n_5955 ,csa_tree_add_12_51_groupi_n_3856 ,csa_tree_add_12_51_groupi_n_5828);
  nor csa_tree_add_12_51_groupi_g15818(csa_tree_add_12_51_groupi_n_5954 ,csa_tree_add_12_51_groupi_n_3859 ,csa_tree_add_12_51_groupi_n_5829);
  nor csa_tree_add_12_51_groupi_g15819(csa_tree_add_12_51_groupi_n_5953 ,csa_tree_add_12_51_groupi_n_3462 ,csa_tree_add_12_51_groupi_n_5822);
  nor csa_tree_add_12_51_groupi_g15820(csa_tree_add_12_51_groupi_n_5952 ,csa_tree_add_12_51_groupi_n_3906 ,csa_tree_add_12_51_groupi_n_5833);
  nor csa_tree_add_12_51_groupi_g15821(csa_tree_add_12_51_groupi_n_5951 ,csa_tree_add_12_51_groupi_n_3914 ,csa_tree_add_12_51_groupi_n_5834);
  nor csa_tree_add_12_51_groupi_g15822(csa_tree_add_12_51_groupi_n_5950 ,csa_tree_add_12_51_groupi_n_3878 ,csa_tree_add_12_51_groupi_n_5830);
  nor csa_tree_add_12_51_groupi_g15823(csa_tree_add_12_51_groupi_n_5949 ,csa_tree_add_12_51_groupi_n_3868 ,csa_tree_add_12_51_groupi_n_5831);
  nor csa_tree_add_12_51_groupi_g15824(csa_tree_add_12_51_groupi_n_5948 ,csa_tree_add_12_51_groupi_n_4110 ,csa_tree_add_12_51_groupi_n_5836);
  and csa_tree_add_12_51_groupi_g15825(csa_tree_add_12_51_groupi_n_5991 ,csa_tree_add_12_51_groupi_n_5825 ,csa_tree_add_12_51_groupi_n_5652);
  not csa_tree_add_12_51_groupi_g15826(csa_tree_add_12_51_groupi_n_5942 ,csa_tree_add_12_51_groupi_n_5941);
  not csa_tree_add_12_51_groupi_g15827(csa_tree_add_12_51_groupi_n_5939 ,csa_tree_add_12_51_groupi_n_5938);
  not csa_tree_add_12_51_groupi_g15828(csa_tree_add_12_51_groupi_n_5936 ,csa_tree_add_12_51_groupi_n_5937);
  not csa_tree_add_12_51_groupi_g15829(csa_tree_add_12_51_groupi_n_5934 ,csa_tree_add_12_51_groupi_n_5935);
  not csa_tree_add_12_51_groupi_g15830(csa_tree_add_12_51_groupi_n_5932 ,csa_tree_add_12_51_groupi_n_5933);
  not csa_tree_add_12_51_groupi_g15831(csa_tree_add_12_51_groupi_n_5930 ,csa_tree_add_12_51_groupi_n_5931);
  not csa_tree_add_12_51_groupi_g15832(csa_tree_add_12_51_groupi_n_5928 ,csa_tree_add_12_51_groupi_n_5929);
  not csa_tree_add_12_51_groupi_g15833(csa_tree_add_12_51_groupi_n_5925 ,csa_tree_add_12_51_groupi_n_5924);
  not csa_tree_add_12_51_groupi_g15834(csa_tree_add_12_51_groupi_n_5923 ,csa_tree_add_12_51_groupi_n_5922);
  not csa_tree_add_12_51_groupi_g15835(csa_tree_add_12_51_groupi_n_5916 ,csa_tree_add_12_51_groupi_n_5915);
  not csa_tree_add_12_51_groupi_g15836(csa_tree_add_12_51_groupi_n_5914 ,csa_tree_add_12_51_groupi_n_5913);
  not csa_tree_add_12_51_groupi_g15837(csa_tree_add_12_51_groupi_n_5912 ,csa_tree_add_12_51_groupi_n_5911);
  not csa_tree_add_12_51_groupi_g15838(csa_tree_add_12_51_groupi_n_5910 ,csa_tree_add_12_51_groupi_n_5909);
  not csa_tree_add_12_51_groupi_g15839(csa_tree_add_12_51_groupi_n_5908 ,csa_tree_add_12_51_groupi_n_5907);
  nor csa_tree_add_12_51_groupi_g15840(csa_tree_add_12_51_groupi_n_5906 ,csa_tree_add_12_51_groupi_n_1625 ,csa_tree_add_12_51_groupi_n_807);
  nor csa_tree_add_12_51_groupi_g15841(csa_tree_add_12_51_groupi_n_5905 ,csa_tree_add_12_51_groupi_n_1637 ,csa_tree_add_12_51_groupi_n_908);
  nor csa_tree_add_12_51_groupi_g15842(csa_tree_add_12_51_groupi_n_5904 ,csa_tree_add_12_51_groupi_n_1670 ,csa_tree_add_12_51_groupi_n_810);
  nor csa_tree_add_12_51_groupi_g15843(csa_tree_add_12_51_groupi_n_5903 ,csa_tree_add_12_51_groupi_n_1631 ,csa_tree_add_12_51_groupi_n_809);
  nor csa_tree_add_12_51_groupi_g15844(csa_tree_add_12_51_groupi_n_5902 ,csa_tree_add_12_51_groupi_n_1643 ,csa_tree_add_12_51_groupi_n_1998);
  nor csa_tree_add_12_51_groupi_g15845(csa_tree_add_12_51_groupi_n_5901 ,csa_tree_add_12_51_groupi_n_1658 ,csa_tree_add_12_51_groupi_n_909);
  nor csa_tree_add_12_51_groupi_g15846(csa_tree_add_12_51_groupi_n_5900 ,csa_tree_add_12_51_groupi_n_1649 ,csa_tree_add_12_51_groupi_n_177);
  xnor csa_tree_add_12_51_groupi_g15847(out3[6] ,csa_tree_add_12_51_groupi_n_5711 ,csa_tree_add_12_51_groupi_n_5718);
  xnor csa_tree_add_12_51_groupi_g15848(csa_tree_add_12_51_groupi_n_5898 ,csa_tree_add_12_51_groupi_n_5758 ,csa_tree_add_12_51_groupi_n_5813);
  xnor csa_tree_add_12_51_groupi_g15849(csa_tree_add_12_51_groupi_n_5897 ,csa_tree_add_12_51_groupi_n_5771 ,csa_tree_add_12_51_groupi_n_5745);
  xnor csa_tree_add_12_51_groupi_g15850(csa_tree_add_12_51_groupi_n_5896 ,csa_tree_add_12_51_groupi_n_5818 ,csa_tree_add_12_51_groupi_n_5741);
  xnor csa_tree_add_12_51_groupi_g15851(csa_tree_add_12_51_groupi_n_5895 ,csa_tree_add_12_51_groupi_n_5815 ,csa_tree_add_12_51_groupi_n_5763);
  xnor csa_tree_add_12_51_groupi_g15852(csa_tree_add_12_51_groupi_n_5894 ,csa_tree_add_12_51_groupi_n_5768 ,csa_tree_add_12_51_groupi_n_5770);
  xnor csa_tree_add_12_51_groupi_g15853(csa_tree_add_12_51_groupi_n_5893 ,csa_tree_add_12_51_groupi_n_5759 ,csa_tree_add_12_51_groupi_n_5709);
  xnor csa_tree_add_12_51_groupi_g15854(csa_tree_add_12_51_groupi_n_5892 ,csa_tree_add_12_51_groupi_n_5769 ,csa_tree_add_12_51_groupi_n_5738);
  xnor csa_tree_add_12_51_groupi_g15855(csa_tree_add_12_51_groupi_n_5891 ,csa_tree_add_12_51_groupi_n_0 ,csa_tree_add_12_51_groupi_n_5571);
  xnor csa_tree_add_12_51_groupi_g15856(csa_tree_add_12_51_groupi_n_5890 ,csa_tree_add_12_51_groupi_n_5706 ,csa_tree_add_12_51_groupi_n_5748);
  xnor csa_tree_add_12_51_groupi_g15857(csa_tree_add_12_51_groupi_n_5947 ,csa_tree_add_12_51_groupi_n_1944 ,csa_tree_add_12_51_groupi_n_5784);
  xnor csa_tree_add_12_51_groupi_g15858(csa_tree_add_12_51_groupi_n_5946 ,csa_tree_add_12_51_groupi_n_5774 ,in3[11]);
  xnor csa_tree_add_12_51_groupi_g15859(csa_tree_add_12_51_groupi_n_5945 ,csa_tree_add_12_51_groupi_n_1894 ,csa_tree_add_12_51_groupi_n_5780);
  xnor csa_tree_add_12_51_groupi_g15860(csa_tree_add_12_51_groupi_n_5944 ,csa_tree_add_12_51_groupi_n_108 ,csa_tree_add_12_51_groupi_n_5773);
  xnor csa_tree_add_12_51_groupi_g15861(csa_tree_add_12_51_groupi_n_5943 ,csa_tree_add_12_51_groupi_n_5542 ,csa_tree_add_12_51_groupi_n_5721);
  xnor csa_tree_add_12_51_groupi_g15862(csa_tree_add_12_51_groupi_n_5941 ,csa_tree_add_12_51_groupi_n_5565 ,csa_tree_add_12_51_groupi_n_5725);
  xnor csa_tree_add_12_51_groupi_g15863(csa_tree_add_12_51_groupi_n_5940 ,csa_tree_add_12_51_groupi_n_1949 ,csa_tree_add_12_51_groupi_n_5786);
  xnor csa_tree_add_12_51_groupi_g15864(csa_tree_add_12_51_groupi_n_5938 ,csa_tree_add_12_51_groupi_n_5781 ,in4[2]);
  xnor csa_tree_add_12_51_groupi_g15865(csa_tree_add_12_51_groupi_n_5937 ,csa_tree_add_12_51_groupi_n_5588 ,csa_tree_add_12_51_groupi_n_5724);
  xnor csa_tree_add_12_51_groupi_g15866(csa_tree_add_12_51_groupi_n_5935 ,csa_tree_add_12_51_groupi_n_5562 ,csa_tree_add_12_51_groupi_n_5722);
  xnor csa_tree_add_12_51_groupi_g15867(csa_tree_add_12_51_groupi_n_5933 ,csa_tree_add_12_51_groupi_n_5677 ,csa_tree_add_12_51_groupi_n_5723);
  xnor csa_tree_add_12_51_groupi_g15868(csa_tree_add_12_51_groupi_n_5931 ,csa_tree_add_12_51_groupi_n_5816 ,csa_tree_add_12_51_groupi_n_5720);
  xnor csa_tree_add_12_51_groupi_g15869(csa_tree_add_12_51_groupi_n_5929 ,csa_tree_add_12_51_groupi_n_5590 ,csa_tree_add_12_51_groupi_n_5726);
  xnor csa_tree_add_12_51_groupi_g15870(csa_tree_add_12_51_groupi_n_5927 ,csa_tree_add_12_51_groupi_n_5596 ,csa_tree_add_12_51_groupi_n_5719);
  xnor csa_tree_add_12_51_groupi_g15871(csa_tree_add_12_51_groupi_n_5926 ,csa_tree_add_12_51_groupi_n_5713 ,csa_tree_add_12_51_groupi_n_5717);
  xnor csa_tree_add_12_51_groupi_g15872(csa_tree_add_12_51_groupi_n_5924 ,csa_tree_add_12_51_groupi_n_5776 ,in2[5]);
  xnor csa_tree_add_12_51_groupi_g15873(csa_tree_add_12_51_groupi_n_5922 ,csa_tree_add_12_51_groupi_n_5775 ,csa_tree_add_12_51_groupi_n_1932);
  xnor csa_tree_add_12_51_groupi_g15874(csa_tree_add_12_51_groupi_n_5921 ,csa_tree_add_12_51_groupi_n_5778 ,in2[11]);
  xnor csa_tree_add_12_51_groupi_g15875(csa_tree_add_12_51_groupi_n_5920 ,csa_tree_add_12_51_groupi_n_5779 ,in4[11]);
  xnor csa_tree_add_12_51_groupi_g15876(csa_tree_add_12_51_groupi_n_5919 ,csa_tree_add_12_51_groupi_n_5710 ,csa_tree_add_12_51_groupi_n_5727);
  xnor csa_tree_add_12_51_groupi_g15877(csa_tree_add_12_51_groupi_n_5918 ,csa_tree_add_12_51_groupi_n_5678 ,csa_tree_add_12_51_groupi_n_5729);
  xnor csa_tree_add_12_51_groupi_g15878(csa_tree_add_12_51_groupi_n_5917 ,csa_tree_add_12_51_groupi_n_5564 ,csa_tree_add_12_51_groupi_n_5728);
  xnor csa_tree_add_12_51_groupi_g15879(csa_tree_add_12_51_groupi_n_5915 ,csa_tree_add_12_51_groupi_n_5783 ,in3[2]);
  xnor csa_tree_add_12_51_groupi_g15880(csa_tree_add_12_51_groupi_n_5913 ,csa_tree_add_12_51_groupi_n_5772 ,in2[14]);
  xnor csa_tree_add_12_51_groupi_g15881(csa_tree_add_12_51_groupi_n_5911 ,csa_tree_add_12_51_groupi_n_5777 ,csa_tree_add_12_51_groupi_n_2366);
  xnor csa_tree_add_12_51_groupi_g15882(csa_tree_add_12_51_groupi_n_5909 ,csa_tree_add_12_51_groupi_n_5785 ,in4[8]);
  xnor csa_tree_add_12_51_groupi_g15883(csa_tree_add_12_51_groupi_n_5907 ,csa_tree_add_12_51_groupi_n_118 ,csa_tree_add_12_51_groupi_n_5782);
  not csa_tree_add_12_51_groupi_g15885(csa_tree_add_12_51_groupi_n_5878 ,csa_tree_add_12_51_groupi_n_5879);
  not csa_tree_add_12_51_groupi_g15886(csa_tree_add_12_51_groupi_n_5875 ,csa_tree_add_12_51_groupi_n_5876);
  not csa_tree_add_12_51_groupi_g15887(csa_tree_add_12_51_groupi_n_5874 ,csa_tree_add_12_51_groupi_n_5873);
  nor csa_tree_add_12_51_groupi_g15888(csa_tree_add_12_51_groupi_n_5872 ,csa_tree_add_12_51_groupi_n_5575 ,csa_tree_add_12_51_groupi_n_5766);
  nor csa_tree_add_12_51_groupi_g15889(csa_tree_add_12_51_groupi_n_5871 ,csa_tree_add_12_51_groupi_n_4921 ,csa_tree_add_12_51_groupi_n_5811);
  nor csa_tree_add_12_51_groupi_g15890(csa_tree_add_12_51_groupi_n_5870 ,csa_tree_add_12_51_groupi_n_5706 ,csa_tree_add_12_51_groupi_n_5747);
  and csa_tree_add_12_51_groupi_g15891(csa_tree_add_12_51_groupi_n_5869 ,csa_tree_add_12_51_groupi_n_5758 ,csa_tree_add_12_51_groupi_n_5813);
  or csa_tree_add_12_51_groupi_g15892(csa_tree_add_12_51_groupi_n_5868 ,csa_tree_add_12_51_groupi_n_5758 ,csa_tree_add_12_51_groupi_n_5813);
  or csa_tree_add_12_51_groupi_g15893(csa_tree_add_12_51_groupi_n_5867 ,csa_tree_add_12_51_groupi_n_5705 ,csa_tree_add_12_51_groupi_n_5748);
  and csa_tree_add_12_51_groupi_g15894(csa_tree_add_12_51_groupi_n_5866 ,csa_tree_add_12_51_groupi_n_5739 ,csa_tree_add_12_51_groupi_n_5738);
  nor csa_tree_add_12_51_groupi_g15895(csa_tree_add_12_51_groupi_n_5865 ,csa_tree_add_12_51_groupi_n_5739 ,csa_tree_add_12_51_groupi_n_5738);
  or csa_tree_add_12_51_groupi_g15896(csa_tree_add_12_51_groupi_n_5864 ,csa_tree_add_12_51_groupi_n_5741 ,csa_tree_add_12_51_groupi_n_5742);
  or csa_tree_add_12_51_groupi_g15897(csa_tree_add_12_51_groupi_n_5863 ,csa_tree_add_12_51_groupi_n_5744 ,csa_tree_add_12_51_groupi_n_4);
  nor csa_tree_add_12_51_groupi_g15898(csa_tree_add_12_51_groupi_n_5862 ,csa_tree_add_12_51_groupi_n_5740 ,csa_tree_add_12_51_groupi_n_5743);
  nor csa_tree_add_12_51_groupi_g15899(csa_tree_add_12_51_groupi_n_5861 ,csa_tree_add_12_51_groupi_n_5745 ,csa_tree_add_12_51_groupi_n_5746);
  or csa_tree_add_12_51_groupi_g15900(csa_tree_add_12_51_groupi_n_5860 ,csa_tree_add_12_51_groupi_n_4920 ,csa_tree_add_12_51_groupi_n_5812);
  and csa_tree_add_12_51_groupi_g15901(csa_tree_add_12_51_groupi_n_5859 ,csa_tree_add_12_51_groupi_n_5759 ,csa_tree_add_12_51_groupi_n_5709);
  or csa_tree_add_12_51_groupi_g15902(csa_tree_add_12_51_groupi_n_5858 ,csa_tree_add_12_51_groupi_n_5759 ,csa_tree_add_12_51_groupi_n_5709);
  nor csa_tree_add_12_51_groupi_g15903(csa_tree_add_12_51_groupi_n_5857 ,csa_tree_add_12_51_groupi_n_5752 ,csa_tree_add_12_51_groupi_n_5767);
  or csa_tree_add_12_51_groupi_g15904(csa_tree_add_12_51_groupi_n_5856 ,csa_tree_add_12_51_groupi_n_5751 ,csa_tree_add_12_51_groupi_n_5768);
  and csa_tree_add_12_51_groupi_g15905(csa_tree_add_12_51_groupi_n_5855 ,csa_tree_add_12_51_groupi_n_5575 ,csa_tree_add_12_51_groupi_n_5766);
  and csa_tree_add_12_51_groupi_g15906(csa_tree_add_12_51_groupi_n_5889 ,csa_tree_add_12_51_groupi_n_5700 ,csa_tree_add_12_51_groupi_n_5808);
  and csa_tree_add_12_51_groupi_g15907(csa_tree_add_12_51_groupi_n_5888 ,csa_tree_add_12_51_groupi_n_5804 ,csa_tree_add_12_51_groupi_n_5694);
  or csa_tree_add_12_51_groupi_g15908(csa_tree_add_12_51_groupi_n_5887 ,csa_tree_add_12_51_groupi_n_5686 ,csa_tree_add_12_51_groupi_n_5810);
  and csa_tree_add_12_51_groupi_g15909(csa_tree_add_12_51_groupi_n_5886 ,csa_tree_add_12_51_groupi_n_5695 ,csa_tree_add_12_51_groupi_n_5791);
  or csa_tree_add_12_51_groupi_g15910(csa_tree_add_12_51_groupi_n_5885 ,csa_tree_add_12_51_groupi_n_5693 ,csa_tree_add_12_51_groupi_n_5801);
  or csa_tree_add_12_51_groupi_g15911(csa_tree_add_12_51_groupi_n_5884 ,csa_tree_add_12_51_groupi_n_5649 ,csa_tree_add_12_51_groupi_n_5794);
  and csa_tree_add_12_51_groupi_g15912(csa_tree_add_12_51_groupi_n_5883 ,csa_tree_add_12_51_groupi_n_5675 ,csa_tree_add_12_51_groupi_n_5795);
  and csa_tree_add_12_51_groupi_g15913(csa_tree_add_12_51_groupi_n_5882 ,csa_tree_add_12_51_groupi_n_2436 ,csa_tree_add_12_51_groupi_n_5793);
  and csa_tree_add_12_51_groupi_g15914(csa_tree_add_12_51_groupi_n_5881 ,csa_tree_add_12_51_groupi_n_5704 ,csa_tree_add_12_51_groupi_n_5789);
  or csa_tree_add_12_51_groupi_g15915(csa_tree_add_12_51_groupi_n_5880 ,csa_tree_add_12_51_groupi_n_5792 ,csa_tree_add_12_51_groupi_n_5698);
  or csa_tree_add_12_51_groupi_g15916(csa_tree_add_12_51_groupi_n_5879 ,csa_tree_add_12_51_groupi_n_5683 ,csa_tree_add_12_51_groupi_n_5788);
  and csa_tree_add_12_51_groupi_g15917(csa_tree_add_12_51_groupi_n_5877 ,csa_tree_add_12_51_groupi_n_5689 ,csa_tree_add_12_51_groupi_n_5809);
  or csa_tree_add_12_51_groupi_g15918(csa_tree_add_12_51_groupi_n_5876 ,csa_tree_add_12_51_groupi_n_5684 ,csa_tree_add_12_51_groupi_n_5790);
  or csa_tree_add_12_51_groupi_g15919(csa_tree_add_12_51_groupi_n_5873 ,csa_tree_add_12_51_groupi_n_5787 ,csa_tree_add_12_51_groupi_n_5679);
  not csa_tree_add_12_51_groupi_g15920(csa_tree_add_12_51_groupi_n_5849 ,csa_tree_add_12_51_groupi_n_5850);
  not csa_tree_add_12_51_groupi_g15921(csa_tree_add_12_51_groupi_n_5847 ,csa_tree_add_12_51_groupi_n_5848);
  not csa_tree_add_12_51_groupi_g15922(csa_tree_add_12_51_groupi_n_5845 ,csa_tree_add_12_51_groupi_n_5846);
  or csa_tree_add_12_51_groupi_g15923(csa_tree_add_12_51_groupi_n_5841 ,csa_tree_add_12_51_groupi_n_3727 ,csa_tree_add_12_51_groupi_n_5731);
  nor csa_tree_add_12_51_groupi_g15924(csa_tree_add_12_51_groupi_n_5840 ,csa_tree_add_12_51_groupi_n_5761 ,csa_tree_add_12_51_groupi_n_5571);
  and csa_tree_add_12_51_groupi_g15925(csa_tree_add_12_51_groupi_n_5839 ,csa_tree_add_12_51_groupi_n_5761 ,csa_tree_add_12_51_groupi_n_5571);
  and csa_tree_add_12_51_groupi_g15926(csa_tree_add_12_51_groupi_n_5838 ,csa_tree_add_12_51_groupi_n_5587 ,csa_tree_add_12_51_groupi_n_5757);
  nor csa_tree_add_12_51_groupi_g15927(csa_tree_add_12_51_groupi_n_5837 ,csa_tree_add_12_51_groupi_n_5587 ,csa_tree_add_12_51_groupi_n_5757);
  or csa_tree_add_12_51_groupi_g15928(csa_tree_add_12_51_groupi_n_5836 ,csa_tree_add_12_51_groupi_n_3363 ,csa_tree_add_12_51_groupi_n_5800);
  or csa_tree_add_12_51_groupi_g15929(csa_tree_add_12_51_groupi_n_5835 ,csa_tree_add_12_51_groupi_n_3648 ,csa_tree_add_12_51_groupi_n_5802);
  or csa_tree_add_12_51_groupi_g15930(csa_tree_add_12_51_groupi_n_5834 ,csa_tree_add_12_51_groupi_n_3713 ,csa_tree_add_12_51_groupi_n_5803);
  or csa_tree_add_12_51_groupi_g15931(csa_tree_add_12_51_groupi_n_5833 ,csa_tree_add_12_51_groupi_n_3653 ,csa_tree_add_12_51_groupi_n_5805);
  or csa_tree_add_12_51_groupi_g15932(csa_tree_add_12_51_groupi_n_5832 ,csa_tree_add_12_51_groupi_n_3731 ,csa_tree_add_12_51_groupi_n_5806);
  or csa_tree_add_12_51_groupi_g15933(csa_tree_add_12_51_groupi_n_5831 ,csa_tree_add_12_51_groupi_n_3585 ,csa_tree_add_12_51_groupi_n_5736);
  or csa_tree_add_12_51_groupi_g15934(csa_tree_add_12_51_groupi_n_5830 ,csa_tree_add_12_51_groupi_n_3608 ,csa_tree_add_12_51_groupi_n_5737);
  or csa_tree_add_12_51_groupi_g15935(csa_tree_add_12_51_groupi_n_5829 ,csa_tree_add_12_51_groupi_n_3698 ,csa_tree_add_12_51_groupi_n_5735);
  or csa_tree_add_12_51_groupi_g15936(csa_tree_add_12_51_groupi_n_5828 ,csa_tree_add_12_51_groupi_n_3618 ,csa_tree_add_12_51_groupi_n_5734);
  or csa_tree_add_12_51_groupi_g15937(csa_tree_add_12_51_groupi_n_5827 ,csa_tree_add_12_51_groupi_n_3599 ,csa_tree_add_12_51_groupi_n_5733);
  or csa_tree_add_12_51_groupi_g15938(csa_tree_add_12_51_groupi_n_5826 ,csa_tree_add_12_51_groupi_n_3693 ,csa_tree_add_12_51_groupi_n_5732);
  or csa_tree_add_12_51_groupi_g15939(csa_tree_add_12_51_groupi_n_5825 ,csa_tree_add_12_51_groupi_n_5653 ,csa_tree_add_12_51_groupi_n_5817);
  or csa_tree_add_12_51_groupi_g15940(csa_tree_add_12_51_groupi_n_5824 ,csa_tree_add_12_51_groupi_n_3124 ,csa_tree_add_12_51_groupi_n_5797);
  or csa_tree_add_12_51_groupi_g15941(csa_tree_add_12_51_groupi_n_5823 ,csa_tree_add_12_51_groupi_n_3164 ,csa_tree_add_12_51_groupi_n_5798);
  or csa_tree_add_12_51_groupi_g15942(csa_tree_add_12_51_groupi_n_5822 ,csa_tree_add_12_51_groupi_n_3074 ,csa_tree_add_12_51_groupi_n_5799);
  xnor csa_tree_add_12_51_groupi_g15943(csa_tree_add_12_51_groupi_n_5821 ,csa_tree_add_12_51_groupi_n_5714 ,csa_tree_add_12_51_groupi_n_5587);
  xor csa_tree_add_12_51_groupi_g15944(csa_tree_add_12_51_groupi_n_5820 ,csa_tree_add_12_51_groupi_n_5575 ,csa_tree_add_12_51_groupi_n_5712);
  xnor csa_tree_add_12_51_groupi_g15945(csa_tree_add_12_51_groupi_n_5819 ,csa_tree_add_12_51_groupi_n_5716 ,csa_tree_add_12_51_groupi_n_5574);
  xnor csa_tree_add_12_51_groupi_g15946(csa_tree_add_12_51_groupi_n_5854 ,csa_tree_add_12_51_groupi_n_5580 ,csa_tree_add_12_51_groupi_n_5644);
  and csa_tree_add_12_51_groupi_g15947(csa_tree_add_12_51_groupi_n_5853 ,csa_tree_add_12_51_groupi_n_5670 ,csa_tree_add_12_51_groupi_n_5796);
  xnor csa_tree_add_12_51_groupi_g15948(csa_tree_add_12_51_groupi_n_5852 ,csa_tree_add_12_51_groupi_n_5428 ,csa_tree_add_12_51_groupi_n_5647);
  xnor csa_tree_add_12_51_groupi_g15949(csa_tree_add_12_51_groupi_n_5851 ,csa_tree_add_12_51_groupi_n_5576 ,csa_tree_add_12_51_groupi_n_5643);
  xnor csa_tree_add_12_51_groupi_g15950(csa_tree_add_12_51_groupi_n_5850 ,csa_tree_add_12_51_groupi_n_5581 ,csa_tree_add_12_51_groupi_n_5642);
  xnor csa_tree_add_12_51_groupi_g15951(csa_tree_add_12_51_groupi_n_5848 ,csa_tree_add_12_51_groupi_n_4841 ,csa_tree_add_12_51_groupi_n_5648);
  xnor csa_tree_add_12_51_groupi_g15952(csa_tree_add_12_51_groupi_n_5846 ,csa_tree_add_12_51_groupi_n_5429 ,csa_tree_add_12_51_groupi_n_5646);
  or csa_tree_add_12_51_groupi_g15953(csa_tree_add_12_51_groupi_n_5844 ,csa_tree_add_12_51_groupi_n_5807 ,csa_tree_add_12_51_groupi_n_5651);
  xnor csa_tree_add_12_51_groupi_g15954(csa_tree_add_12_51_groupi_n_5843 ,csa_tree_add_12_51_groupi_n_5379 ,csa_tree_add_12_51_groupi_n_5645);
  xnor csa_tree_add_12_51_groupi_g15955(csa_tree_add_12_51_groupi_n_5842 ,csa_tree_add_12_51_groupi_n_5715 ,csa_tree_add_12_51_groupi_n_2564);
  not csa_tree_add_12_51_groupi_g15956(csa_tree_add_12_51_groupi_n_5817 ,csa_tree_add_12_51_groupi_n_5816);
  not csa_tree_add_12_51_groupi_g15957(csa_tree_add_12_51_groupi_n_5811 ,csa_tree_add_12_51_groupi_n_5812);
  nor csa_tree_add_12_51_groupi_g15958(csa_tree_add_12_51_groupi_n_5810 ,csa_tree_add_12_51_groupi_n_5595 ,csa_tree_add_12_51_groupi_n_5703);
  or csa_tree_add_12_51_groupi_g15959(csa_tree_add_12_51_groupi_n_5809 ,csa_tree_add_12_51_groupi_n_5591 ,csa_tree_add_12_51_groupi_n_5701);
  or csa_tree_add_12_51_groupi_g15960(csa_tree_add_12_51_groupi_n_5808 ,csa_tree_add_12_51_groupi_n_5592 ,csa_tree_add_12_51_groupi_n_5699);
  and csa_tree_add_12_51_groupi_g15961(csa_tree_add_12_51_groupi_n_5807 ,csa_tree_add_12_51_groupi_n_5650 ,csa_tree_add_12_51_groupi_n_5713);
  nor csa_tree_add_12_51_groupi_g15962(csa_tree_add_12_51_groupi_n_5806 ,csa_tree_add_12_51_groupi_n_1871 ,csa_tree_add_12_51_groupi_n_794);
  nor csa_tree_add_12_51_groupi_g15963(csa_tree_add_12_51_groupi_n_5805 ,csa_tree_add_12_51_groupi_n_1880 ,csa_tree_add_12_51_groupi_n_797);
  or csa_tree_add_12_51_groupi_g15964(csa_tree_add_12_51_groupi_n_5804 ,csa_tree_add_12_51_groupi_n_5696 ,csa_tree_add_12_51_groupi_n_5710);
  nor csa_tree_add_12_51_groupi_g15965(csa_tree_add_12_51_groupi_n_5803 ,csa_tree_add_12_51_groupi_n_1868 ,csa_tree_add_12_51_groupi_n_159);
  nor csa_tree_add_12_51_groupi_g15966(csa_tree_add_12_51_groupi_n_5802 ,csa_tree_add_12_51_groupi_n_1877 ,csa_tree_add_12_51_groupi_n_794);
  nor csa_tree_add_12_51_groupi_g15967(csa_tree_add_12_51_groupi_n_5801 ,csa_tree_add_12_51_groupi_n_5678 ,csa_tree_add_12_51_groupi_n_5690);
  nor csa_tree_add_12_51_groupi_g15968(csa_tree_add_12_51_groupi_n_5800 ,csa_tree_add_12_51_groupi_n_1889 ,csa_tree_add_12_51_groupi_n_795);
  nor csa_tree_add_12_51_groupi_g15969(csa_tree_add_12_51_groupi_n_5799 ,csa_tree_add_12_51_groupi_n_1859 ,csa_tree_add_12_51_groupi_n_798);
  nor csa_tree_add_12_51_groupi_g15970(csa_tree_add_12_51_groupi_n_5798 ,csa_tree_add_12_51_groupi_n_1856 ,csa_tree_add_12_51_groupi_n_843);
  nor csa_tree_add_12_51_groupi_g15971(csa_tree_add_12_51_groupi_n_5797 ,csa_tree_add_12_51_groupi_n_1850 ,csa_tree_add_12_51_groupi_n_842);
  or csa_tree_add_12_51_groupi_g15972(csa_tree_add_12_51_groupi_n_5796 ,csa_tree_add_12_51_groupi_n_5539 ,csa_tree_add_12_51_groupi_n_5669);
  or csa_tree_add_12_51_groupi_g15973(csa_tree_add_12_51_groupi_n_5795 ,csa_tree_add_12_51_groupi_n_5594 ,csa_tree_add_12_51_groupi_n_5674);
  and csa_tree_add_12_51_groupi_g15974(csa_tree_add_12_51_groupi_n_5794 ,csa_tree_add_12_51_groupi_n_5711 ,csa_tree_add_12_51_groupi_n_5702);
  or csa_tree_add_12_51_groupi_g15975(csa_tree_add_12_51_groupi_n_5793 ,csa_tree_add_12_51_groupi_n_2431 ,csa_tree_add_12_51_groupi_n_5715);
  and csa_tree_add_12_51_groupi_g15976(csa_tree_add_12_51_groupi_n_5792 ,csa_tree_add_12_51_groupi_n_5542 ,csa_tree_add_12_51_groupi_n_5691);
  or csa_tree_add_12_51_groupi_g15977(csa_tree_add_12_51_groupi_n_5791 ,csa_tree_add_12_51_groupi_n_5597 ,csa_tree_add_12_51_groupi_n_5697);
  nor csa_tree_add_12_51_groupi_g15978(csa_tree_add_12_51_groupi_n_5790 ,csa_tree_add_12_51_groupi_n_5543 ,csa_tree_add_12_51_groupi_n_5687);
  or csa_tree_add_12_51_groupi_g15979(csa_tree_add_12_51_groupi_n_5789 ,csa_tree_add_12_51_groupi_n_5589 ,csa_tree_add_12_51_groupi_n_5685);
  nor csa_tree_add_12_51_groupi_g15980(csa_tree_add_12_51_groupi_n_5788 ,csa_tree_add_12_51_groupi_n_5682 ,csa_tree_add_12_51_groupi_n_5540);
  and csa_tree_add_12_51_groupi_g15981(csa_tree_add_12_51_groupi_n_5787 ,csa_tree_add_12_51_groupi_n_5677 ,csa_tree_add_12_51_groupi_n_5680);
  nor csa_tree_add_12_51_groupi_g15982(csa_tree_add_12_51_groupi_n_5786 ,csa_tree_add_12_51_groupi_n_4101 ,csa_tree_add_12_51_groupi_n_5666);
  nor csa_tree_add_12_51_groupi_g15983(csa_tree_add_12_51_groupi_n_5785 ,csa_tree_add_12_51_groupi_n_4035 ,csa_tree_add_12_51_groupi_n_5668);
  nor csa_tree_add_12_51_groupi_g15984(csa_tree_add_12_51_groupi_n_5784 ,csa_tree_add_12_51_groupi_n_4036 ,csa_tree_add_12_51_groupi_n_5667);
  nor csa_tree_add_12_51_groupi_g15985(csa_tree_add_12_51_groupi_n_5783 ,csa_tree_add_12_51_groupi_n_3460 ,csa_tree_add_12_51_groupi_n_5654);
  nor csa_tree_add_12_51_groupi_g15986(csa_tree_add_12_51_groupi_n_5782 ,csa_tree_add_12_51_groupi_n_3473 ,csa_tree_add_12_51_groupi_n_5655);
  nor csa_tree_add_12_51_groupi_g15987(csa_tree_add_12_51_groupi_n_5781 ,csa_tree_add_12_51_groupi_n_3472 ,csa_tree_add_12_51_groupi_n_5656);
  nor csa_tree_add_12_51_groupi_g15988(csa_tree_add_12_51_groupi_n_5780 ,csa_tree_add_12_51_groupi_n_3888 ,csa_tree_add_12_51_groupi_n_5663);
  nor csa_tree_add_12_51_groupi_g15989(csa_tree_add_12_51_groupi_n_5779 ,csa_tree_add_12_51_groupi_n_3844 ,csa_tree_add_12_51_groupi_n_5658);
  nor csa_tree_add_12_51_groupi_g15990(csa_tree_add_12_51_groupi_n_5778 ,csa_tree_add_12_51_groupi_n_3831 ,csa_tree_add_12_51_groupi_n_5657);
  nor csa_tree_add_12_51_groupi_g15991(csa_tree_add_12_51_groupi_n_5777 ,csa_tree_add_12_51_groupi_n_3916 ,csa_tree_add_12_51_groupi_n_5665);
  nor csa_tree_add_12_51_groupi_g15992(csa_tree_add_12_51_groupi_n_5776 ,csa_tree_add_12_51_groupi_n_3851 ,csa_tree_add_12_51_groupi_n_5659);
  nor csa_tree_add_12_51_groupi_g15993(csa_tree_add_12_51_groupi_n_5775 ,csa_tree_add_12_51_groupi_n_3852 ,csa_tree_add_12_51_groupi_n_5660);
  nor csa_tree_add_12_51_groupi_g15994(csa_tree_add_12_51_groupi_n_5774 ,csa_tree_add_12_51_groupi_n_3857 ,csa_tree_add_12_51_groupi_n_5661);
  nor csa_tree_add_12_51_groupi_g15995(csa_tree_add_12_51_groupi_n_5773 ,csa_tree_add_12_51_groupi_n_3866 ,csa_tree_add_12_51_groupi_n_5662);
  nor csa_tree_add_12_51_groupi_g15996(csa_tree_add_12_51_groupi_n_5772 ,csa_tree_add_12_51_groupi_n_3910 ,csa_tree_add_12_51_groupi_n_5664);
  and csa_tree_add_12_51_groupi_g15997(csa_tree_add_12_51_groupi_n_5818 ,csa_tree_add_12_51_groupi_n_5623 ,csa_tree_add_12_51_groupi_n_5673);
  or csa_tree_add_12_51_groupi_g15998(csa_tree_add_12_51_groupi_n_5816 ,csa_tree_add_12_51_groupi_n_5626 ,csa_tree_add_12_51_groupi_n_5692);
  and csa_tree_add_12_51_groupi_g15999(csa_tree_add_12_51_groupi_n_5815 ,csa_tree_add_12_51_groupi_n_5688 ,csa_tree_add_12_51_groupi_n_5627);
  and csa_tree_add_12_51_groupi_g16000(csa_tree_add_12_51_groupi_n_5814 ,csa_tree_add_12_51_groupi_n_5621 ,csa_tree_add_12_51_groupi_n_5671);
  or csa_tree_add_12_51_groupi_g16001(csa_tree_add_12_51_groupi_n_5813 ,csa_tree_add_12_51_groupi_n_5630 ,csa_tree_add_12_51_groupi_n_5681);
  or csa_tree_add_12_51_groupi_g16002(csa_tree_add_12_51_groupi_n_5812 ,csa_tree_add_12_51_groupi_n_4801 ,csa_tree_add_12_51_groupi_n_5672);
  not csa_tree_add_12_51_groupi_g16003(csa_tree_add_12_51_groupi_n_5768 ,csa_tree_add_12_51_groupi_n_5767);
  not csa_tree_add_12_51_groupi_g16004(csa_tree_add_12_51_groupi_n_5764 ,csa_tree_add_12_51_groupi_n_5765);
  not csa_tree_add_12_51_groupi_g16005(csa_tree_add_12_51_groupi_n_5763 ,csa_tree_add_12_51_groupi_n_5762);
  not csa_tree_add_12_51_groupi_g16006(csa_tree_add_12_51_groupi_n_5756 ,csa_tree_add_12_51_groupi_n_5755);
  not csa_tree_add_12_51_groupi_g16007(csa_tree_add_12_51_groupi_n_5754 ,csa_tree_add_12_51_groupi_n_5753);
  not csa_tree_add_12_51_groupi_g16008(csa_tree_add_12_51_groupi_n_5752 ,csa_tree_add_12_51_groupi_n_5751);
  not csa_tree_add_12_51_groupi_g16009(csa_tree_add_12_51_groupi_n_5750 ,csa_tree_add_12_51_groupi_n_5749);
  not csa_tree_add_12_51_groupi_g16010(csa_tree_add_12_51_groupi_n_5747 ,csa_tree_add_12_51_groupi_n_5748);
  not csa_tree_add_12_51_groupi_g16011(csa_tree_add_12_51_groupi_n_5746 ,csa_tree_add_12_51_groupi_n_4);
  not csa_tree_add_12_51_groupi_g16012(csa_tree_add_12_51_groupi_n_5744 ,csa_tree_add_12_51_groupi_n_5745);
  not csa_tree_add_12_51_groupi_g16013(csa_tree_add_12_51_groupi_n_5742 ,csa_tree_add_12_51_groupi_n_5743);
  not csa_tree_add_12_51_groupi_g16014(csa_tree_add_12_51_groupi_n_5741 ,csa_tree_add_12_51_groupi_n_5740);
  nor csa_tree_add_12_51_groupi_g16015(csa_tree_add_12_51_groupi_n_5737 ,csa_tree_add_12_51_groupi_n_1883 ,csa_tree_add_12_51_groupi_n_795);
  nor csa_tree_add_12_51_groupi_g16016(csa_tree_add_12_51_groupi_n_5736 ,csa_tree_add_12_51_groupi_n_1853 ,csa_tree_add_12_51_groupi_n_842);
  nor csa_tree_add_12_51_groupi_g16017(csa_tree_add_12_51_groupi_n_5735 ,csa_tree_add_12_51_groupi_n_1874 ,csa_tree_add_12_51_groupi_n_798);
  nor csa_tree_add_12_51_groupi_g16018(csa_tree_add_12_51_groupi_n_5734 ,csa_tree_add_12_51_groupi_n_1865 ,csa_tree_add_12_51_groupi_n_797);
  nor csa_tree_add_12_51_groupi_g16019(csa_tree_add_12_51_groupi_n_5733 ,csa_tree_add_12_51_groupi_n_1862 ,csa_tree_add_12_51_groupi_n_1986);
  nor csa_tree_add_12_51_groupi_g16020(csa_tree_add_12_51_groupi_n_5732 ,csa_tree_add_12_51_groupi_n_1886 ,csa_tree_add_12_51_groupi_n_843);
  nor csa_tree_add_12_51_groupi_g16021(csa_tree_add_12_51_groupi_n_5731 ,csa_tree_add_12_51_groupi_n_1847 ,csa_tree_add_12_51_groupi_n_159);
  xnor csa_tree_add_12_51_groupi_g16022(out3[5] ,csa_tree_add_12_51_groupi_n_5479 ,csa_tree_add_12_51_groupi_n_5551);
  xnor csa_tree_add_12_51_groupi_g16023(csa_tree_add_12_51_groupi_n_5729 ,csa_tree_add_12_51_groupi_n_5572 ,csa_tree_add_12_51_groupi_n_5473);
  xnor csa_tree_add_12_51_groupi_g16024(csa_tree_add_12_51_groupi_n_5728 ,csa_tree_add_12_51_groupi_n_5592 ,csa_tree_add_12_51_groupi_n_5408);
  xnor csa_tree_add_12_51_groupi_g16025(csa_tree_add_12_51_groupi_n_5727 ,csa_tree_add_12_51_groupi_n_5583 ,csa_tree_add_12_51_groupi_n_5349);
  xnor csa_tree_add_12_51_groupi_g16026(csa_tree_add_12_51_groupi_n_5726 ,csa_tree_add_12_51_groupi_n_5503 ,csa_tree_add_12_51_groupi_n_5641);
  xnor csa_tree_add_12_51_groupi_g16027(csa_tree_add_12_51_groupi_n_5725 ,csa_tree_add_12_51_groupi_n_4586 ,csa_tree_add_12_51_groupi_n_5595);
  xnor csa_tree_add_12_51_groupi_g16028(csa_tree_add_12_51_groupi_n_5724 ,csa_tree_add_12_51_groupi_n_5568 ,csa_tree_add_12_51_groupi_n_5533);
  xnor csa_tree_add_12_51_groupi_g16029(csa_tree_add_12_51_groupi_n_5723 ,csa_tree_add_12_51_groupi_n_5475 ,csa_tree_add_12_51_groupi_n_5586);
  xnor csa_tree_add_12_51_groupi_g16030(csa_tree_add_12_51_groupi_n_5722 ,csa_tree_add_12_51_groupi_n_5537 ,csa_tree_add_12_51_groupi_n_5594);
  xnor csa_tree_add_12_51_groupi_g16031(csa_tree_add_12_51_groupi_n_5721 ,csa_tree_add_12_51_groupi_n_5406 ,csa_tree_add_12_51_groupi_n_5579);
  xnor csa_tree_add_12_51_groupi_g16032(csa_tree_add_12_51_groupi_n_5720 ,csa_tree_add_12_51_groupi_n_5378 ,csa_tree_add_12_51_groupi_n_5585);
  xnor csa_tree_add_12_51_groupi_g16033(csa_tree_add_12_51_groupi_n_5719 ,csa_tree_add_12_51_groupi_n_5570 ,csa_tree_add_12_51_groupi_n_5531);
  xnor csa_tree_add_12_51_groupi_g16034(csa_tree_add_12_51_groupi_n_5718 ,csa_tree_add_12_51_groupi_n_5577 ,csa_tree_add_12_51_groupi_n_5376);
  xnor csa_tree_add_12_51_groupi_g16035(csa_tree_add_12_51_groupi_n_5717 ,csa_tree_add_12_51_groupi_n_5578 ,csa_tree_add_12_51_groupi_n_5474);
  xnor csa_tree_add_12_51_groupi_g16036(csa_tree_add_12_51_groupi_n_5771 ,csa_tree_add_12_51_groupi_n_1896 ,csa_tree_add_12_51_groupi_n_5607);
  xnor csa_tree_add_12_51_groupi_g16037(csa_tree_add_12_51_groupi_n_5770 ,csa_tree_add_12_51_groupi_n_102 ,csa_tree_add_12_51_groupi_n_5600);
  xnor csa_tree_add_12_51_groupi_g16038(csa_tree_add_12_51_groupi_n_5769 ,csa_tree_add_12_51_groupi_n_1955 ,csa_tree_add_12_51_groupi_n_5612);
  xnor csa_tree_add_12_51_groupi_g16040(csa_tree_add_12_51_groupi_n_5767 ,csa_tree_add_12_51_groupi_n_5385 ,csa_tree_add_12_51_groupi_n_5549);
  xnor csa_tree_add_12_51_groupi_g16041(csa_tree_add_12_51_groupi_n_5766 ,csa_tree_add_12_51_groupi_n_5501 ,csa_tree_add_12_51_groupi_n_5550);
  xnor csa_tree_add_12_51_groupi_g16042(csa_tree_add_12_51_groupi_n_5765 ,csa_tree_add_12_51_groupi_n_5409 ,csa_tree_add_12_51_groupi_n_5552);
  xnor csa_tree_add_12_51_groupi_g16043(csa_tree_add_12_51_groupi_n_5762 ,csa_tree_add_12_51_groupi_n_5424 ,csa_tree_add_12_51_groupi_n_5547);
  xnor csa_tree_add_12_51_groupi_g16044(csa_tree_add_12_51_groupi_n_5761 ,csa_tree_add_12_51_groupi_n_5601 ,in4[8]);
  xnor csa_tree_add_12_51_groupi_g16045(csa_tree_add_12_51_groupi_n_5760 ,csa_tree_add_12_51_groupi_n_1923 ,csa_tree_add_12_51_groupi_n_5606);
  xnor csa_tree_add_12_51_groupi_g16046(csa_tree_add_12_51_groupi_n_5759 ,csa_tree_add_12_51_groupi_n_5417 ,csa_tree_add_12_51_groupi_n_5548);
  xnor csa_tree_add_12_51_groupi_g16047(csa_tree_add_12_51_groupi_n_5758 ,csa_tree_add_12_51_groupi_n_5427 ,csa_tree_add_12_51_groupi_n_5545);
  xnor csa_tree_add_12_51_groupi_g16048(csa_tree_add_12_51_groupi_n_5757 ,csa_tree_add_12_51_groupi_n_5414 ,csa_tree_add_12_51_groupi_n_5544);
  xnor csa_tree_add_12_51_groupi_g16049(csa_tree_add_12_51_groupi_n_5755 ,csa_tree_add_12_51_groupi_n_5418 ,csa_tree_add_12_51_groupi_n_5546);
  xnor csa_tree_add_12_51_groupi_g16050(csa_tree_add_12_51_groupi_n_5753 ,csa_tree_add_12_51_groupi_n_5602 ,in4[2]);
  xnor csa_tree_add_12_51_groupi_g16051(csa_tree_add_12_51_groupi_n_5751 ,csa_tree_add_12_51_groupi_n_1941 ,csa_tree_add_12_51_groupi_n_5604);
  xnor csa_tree_add_12_51_groupi_g16052(csa_tree_add_12_51_groupi_n_5749 ,csa_tree_add_12_51_groupi_n_5603 ,in3[5]);
  xnor csa_tree_add_12_51_groupi_g16053(csa_tree_add_12_51_groupi_n_5748 ,csa_tree_add_12_51_groupi_n_5593 ,csa_tree_add_12_51_groupi_n_4819);
  xnor csa_tree_add_12_51_groupi_g16055(csa_tree_add_12_51_groupi_n_5745 ,csa_tree_add_12_51_groupi_n_5609 ,in4[11]);
  xnor csa_tree_add_12_51_groupi_g16056(csa_tree_add_12_51_groupi_n_5743 ,csa_tree_add_12_51_groupi_n_5610 ,in2[5]);
  xnor csa_tree_add_12_51_groupi_g16057(csa_tree_add_12_51_groupi_n_5740 ,csa_tree_add_12_51_groupi_n_5611 ,in4[5]);
  xnor csa_tree_add_12_51_groupi_g16058(csa_tree_add_12_51_groupi_n_5739 ,csa_tree_add_12_51_groupi_n_5599 ,in4[14]);
  xnor csa_tree_add_12_51_groupi_g16059(csa_tree_add_12_51_groupi_n_5738 ,csa_tree_add_12_51_groupi_n_5598 ,in2[14]);
  not csa_tree_add_12_51_groupi_g16060(csa_tree_add_12_51_groupi_n_5708 ,csa_tree_add_12_51_groupi_n_5707);
  not csa_tree_add_12_51_groupi_g16061(csa_tree_add_12_51_groupi_n_5705 ,csa_tree_add_12_51_groupi_n_5706);
  or csa_tree_add_12_51_groupi_g16062(csa_tree_add_12_51_groupi_n_5704 ,csa_tree_add_12_51_groupi_n_5567 ,csa_tree_add_12_51_groupi_n_5532);
  and csa_tree_add_12_51_groupi_g16063(csa_tree_add_12_51_groupi_n_5703 ,csa_tree_add_12_51_groupi_n_5566 ,csa_tree_add_12_51_groupi_n_4586);
  or csa_tree_add_12_51_groupi_g16064(csa_tree_add_12_51_groupi_n_5702 ,csa_tree_add_12_51_groupi_n_5577 ,csa_tree_add_12_51_groupi_n_5376);
  nor csa_tree_add_12_51_groupi_g16065(csa_tree_add_12_51_groupi_n_5701 ,csa_tree_add_12_51_groupi_n_5503 ,csa_tree_add_12_51_groupi_n_5641);
  or csa_tree_add_12_51_groupi_g16066(csa_tree_add_12_51_groupi_n_5700 ,csa_tree_add_12_51_groupi_n_5563 ,csa_tree_add_12_51_groupi_n_5407);
  nor csa_tree_add_12_51_groupi_g16067(csa_tree_add_12_51_groupi_n_5699 ,csa_tree_add_12_51_groupi_n_5564 ,csa_tree_add_12_51_groupi_n_5408);
  and csa_tree_add_12_51_groupi_g16068(csa_tree_add_12_51_groupi_n_5698 ,csa_tree_add_12_51_groupi_n_5406 ,csa_tree_add_12_51_groupi_n_5579);
  nor csa_tree_add_12_51_groupi_g16069(csa_tree_add_12_51_groupi_n_5697 ,csa_tree_add_12_51_groupi_n_5570 ,csa_tree_add_12_51_groupi_n_5531);
  nor csa_tree_add_12_51_groupi_g16070(csa_tree_add_12_51_groupi_n_5696 ,csa_tree_add_12_51_groupi_n_5583 ,csa_tree_add_12_51_groupi_n_5349);
  or csa_tree_add_12_51_groupi_g16071(csa_tree_add_12_51_groupi_n_5695 ,csa_tree_add_12_51_groupi_n_5569 ,csa_tree_add_12_51_groupi_n_5530);
  or csa_tree_add_12_51_groupi_g16072(csa_tree_add_12_51_groupi_n_5694 ,csa_tree_add_12_51_groupi_n_5582 ,csa_tree_add_12_51_groupi_n_5348);
  and csa_tree_add_12_51_groupi_g16073(csa_tree_add_12_51_groupi_n_5693 ,csa_tree_add_12_51_groupi_n_5572 ,csa_tree_add_12_51_groupi_n_5473);
  nor csa_tree_add_12_51_groupi_g16074(csa_tree_add_12_51_groupi_n_5692 ,csa_tree_add_12_51_groupi_n_5431 ,csa_tree_add_12_51_groupi_n_5625);
  or csa_tree_add_12_51_groupi_g16075(csa_tree_add_12_51_groupi_n_5691 ,csa_tree_add_12_51_groupi_n_5406 ,csa_tree_add_12_51_groupi_n_5579);
  nor csa_tree_add_12_51_groupi_g16076(csa_tree_add_12_51_groupi_n_5690 ,csa_tree_add_12_51_groupi_n_5572 ,csa_tree_add_12_51_groupi_n_5473);
  or csa_tree_add_12_51_groupi_g16077(csa_tree_add_12_51_groupi_n_5689 ,csa_tree_add_12_51_groupi_n_5502 ,csa_tree_add_12_51_groupi_n_5640);
  or csa_tree_add_12_51_groupi_g16078(csa_tree_add_12_51_groupi_n_5688 ,csa_tree_add_12_51_groupi_n_5381 ,csa_tree_add_12_51_groupi_n_5628);
  nor csa_tree_add_12_51_groupi_g16079(csa_tree_add_12_51_groupi_n_5687 ,csa_tree_add_12_51_groupi_n_5420 ,csa_tree_add_12_51_groupi_n_5581);
  nor csa_tree_add_12_51_groupi_g16080(csa_tree_add_12_51_groupi_n_5686 ,csa_tree_add_12_51_groupi_n_5566 ,csa_tree_add_12_51_groupi_n_4586);
  nor csa_tree_add_12_51_groupi_g16081(csa_tree_add_12_51_groupi_n_5685 ,csa_tree_add_12_51_groupi_n_5568 ,csa_tree_add_12_51_groupi_n_5533);
  and csa_tree_add_12_51_groupi_g16082(csa_tree_add_12_51_groupi_n_5684 ,csa_tree_add_12_51_groupi_n_5420 ,csa_tree_add_12_51_groupi_n_5581);
  and csa_tree_add_12_51_groupi_g16083(csa_tree_add_12_51_groupi_n_5683 ,csa_tree_add_12_51_groupi_n_5415 ,csa_tree_add_12_51_groupi_n_5580);
  nor csa_tree_add_12_51_groupi_g16084(csa_tree_add_12_51_groupi_n_5682 ,csa_tree_add_12_51_groupi_n_5415 ,csa_tree_add_12_51_groupi_n_5580);
  and csa_tree_add_12_51_groupi_g16085(csa_tree_add_12_51_groupi_n_5681 ,csa_tree_add_12_51_groupi_n_5379 ,csa_tree_add_12_51_groupi_n_5629);
  or csa_tree_add_12_51_groupi_g16086(csa_tree_add_12_51_groupi_n_5680 ,csa_tree_add_12_51_groupi_n_5475 ,csa_tree_add_12_51_groupi_n_5586);
  and csa_tree_add_12_51_groupi_g16087(csa_tree_add_12_51_groupi_n_5679 ,csa_tree_add_12_51_groupi_n_5475 ,csa_tree_add_12_51_groupi_n_5586);
  and csa_tree_add_12_51_groupi_g16088(csa_tree_add_12_51_groupi_n_5716 ,csa_tree_add_12_51_groupi_n_5528 ,csa_tree_add_12_51_groupi_n_5639);
  and csa_tree_add_12_51_groupi_g16089(csa_tree_add_12_51_groupi_n_5715 ,csa_tree_add_12_51_groupi_n_2434 ,csa_tree_add_12_51_groupi_n_5633);
  and csa_tree_add_12_51_groupi_g16090(csa_tree_add_12_51_groupi_n_5714 ,csa_tree_add_12_51_groupi_n_5517 ,csa_tree_add_12_51_groupi_n_5634);
  or csa_tree_add_12_51_groupi_g16091(csa_tree_add_12_51_groupi_n_5713 ,csa_tree_add_12_51_groupi_n_5520 ,csa_tree_add_12_51_groupi_n_5635);
  and csa_tree_add_12_51_groupi_g16092(csa_tree_add_12_51_groupi_n_5712 ,csa_tree_add_12_51_groupi_n_5518 ,csa_tree_add_12_51_groupi_n_5637);
  or csa_tree_add_12_51_groupi_g16093(csa_tree_add_12_51_groupi_n_5711 ,csa_tree_add_12_51_groupi_n_5624 ,csa_tree_add_12_51_groupi_n_5529);
  and csa_tree_add_12_51_groupi_g16094(csa_tree_add_12_51_groupi_n_5710 ,csa_tree_add_12_51_groupi_n_5514 ,csa_tree_add_12_51_groupi_n_5632);
  or csa_tree_add_12_51_groupi_g16095(csa_tree_add_12_51_groupi_n_5709 ,csa_tree_add_12_51_groupi_n_5631 ,csa_tree_add_12_51_groupi_n_5512);
  or csa_tree_add_12_51_groupi_g16096(csa_tree_add_12_51_groupi_n_5707 ,csa_tree_add_12_51_groupi_n_5526 ,csa_tree_add_12_51_groupi_n_5638);
  or csa_tree_add_12_51_groupi_g16097(csa_tree_add_12_51_groupi_n_5706 ,csa_tree_add_12_51_groupi_n_5522 ,csa_tree_add_12_51_groupi_n_5636);
  or csa_tree_add_12_51_groupi_g16098(csa_tree_add_12_51_groupi_n_5675 ,csa_tree_add_12_51_groupi_n_5561 ,csa_tree_add_12_51_groupi_n_5537);
  nor csa_tree_add_12_51_groupi_g16099(csa_tree_add_12_51_groupi_n_5674 ,csa_tree_add_12_51_groupi_n_5562 ,csa_tree_add_12_51_groupi_n_5536);
  or csa_tree_add_12_51_groupi_g16100(csa_tree_add_12_51_groupi_n_5673 ,csa_tree_add_12_51_groupi_n_5622 ,csa_tree_add_12_51_groupi_n_5430);
  and csa_tree_add_12_51_groupi_g16101(csa_tree_add_12_51_groupi_n_5672 ,csa_tree_add_12_51_groupi_n_5593 ,csa_tree_add_12_51_groupi_n_4800);
  or csa_tree_add_12_51_groupi_g16102(csa_tree_add_12_51_groupi_n_5671 ,csa_tree_add_12_51_groupi_n_5620 ,csa_tree_add_12_51_groupi_n_5510);
  or csa_tree_add_12_51_groupi_g16103(csa_tree_add_12_51_groupi_n_5670 ,csa_tree_add_12_51_groupi_n_5506 ,csa_tree_add_12_51_groupi_n_5576);
  and csa_tree_add_12_51_groupi_g16104(csa_tree_add_12_51_groupi_n_5669 ,csa_tree_add_12_51_groupi_n_5506 ,csa_tree_add_12_51_groupi_n_5576);
  or csa_tree_add_12_51_groupi_g16105(csa_tree_add_12_51_groupi_n_5668 ,csa_tree_add_12_51_groupi_n_3361 ,csa_tree_add_12_51_groupi_n_5614);
  or csa_tree_add_12_51_groupi_g16106(csa_tree_add_12_51_groupi_n_5667 ,csa_tree_add_12_51_groupi_n_3306 ,csa_tree_add_12_51_groupi_n_5560);
  or csa_tree_add_12_51_groupi_g16107(csa_tree_add_12_51_groupi_n_5666 ,csa_tree_add_12_51_groupi_n_3070 ,csa_tree_add_12_51_groupi_n_5615);
  or csa_tree_add_12_51_groupi_g16108(csa_tree_add_12_51_groupi_n_5665 ,csa_tree_add_12_51_groupi_n_3701 ,csa_tree_add_12_51_groupi_n_5613);
  or csa_tree_add_12_51_groupi_g16109(csa_tree_add_12_51_groupi_n_5664 ,csa_tree_add_12_51_groupi_n_3702 ,csa_tree_add_12_51_groupi_n_5619);
  or csa_tree_add_12_51_groupi_g16110(csa_tree_add_12_51_groupi_n_5663 ,csa_tree_add_12_51_groupi_n_3736 ,csa_tree_add_12_51_groupi_n_5553);
  or csa_tree_add_12_51_groupi_g16111(csa_tree_add_12_51_groupi_n_5662 ,csa_tree_add_12_51_groupi_n_3612 ,csa_tree_add_12_51_groupi_n_5559);
  or csa_tree_add_12_51_groupi_g16112(csa_tree_add_12_51_groupi_n_5661 ,csa_tree_add_12_51_groupi_n_3607 ,csa_tree_add_12_51_groupi_n_5558);
  or csa_tree_add_12_51_groupi_g16113(csa_tree_add_12_51_groupi_n_5660 ,csa_tree_add_12_51_groupi_n_3597 ,csa_tree_add_12_51_groupi_n_5557);
  or csa_tree_add_12_51_groupi_g16114(csa_tree_add_12_51_groupi_n_5659 ,csa_tree_add_12_51_groupi_n_3596 ,csa_tree_add_12_51_groupi_n_5556);
  or csa_tree_add_12_51_groupi_g16115(csa_tree_add_12_51_groupi_n_5658 ,csa_tree_add_12_51_groupi_n_3684 ,csa_tree_add_12_51_groupi_n_5555);
  or csa_tree_add_12_51_groupi_g16116(csa_tree_add_12_51_groupi_n_5657 ,csa_tree_add_12_51_groupi_n_3591 ,csa_tree_add_12_51_groupi_n_5554);
  or csa_tree_add_12_51_groupi_g16117(csa_tree_add_12_51_groupi_n_5656 ,csa_tree_add_12_51_groupi_n_3016 ,csa_tree_add_12_51_groupi_n_5618);
  or csa_tree_add_12_51_groupi_g16118(csa_tree_add_12_51_groupi_n_5655 ,csa_tree_add_12_51_groupi_n_3102 ,csa_tree_add_12_51_groupi_n_5617);
  or csa_tree_add_12_51_groupi_g16119(csa_tree_add_12_51_groupi_n_5654 ,csa_tree_add_12_51_groupi_n_3095 ,csa_tree_add_12_51_groupi_n_5616);
  nor csa_tree_add_12_51_groupi_g16120(csa_tree_add_12_51_groupi_n_5653 ,csa_tree_add_12_51_groupi_n_5378 ,csa_tree_add_12_51_groupi_n_5585);
  or csa_tree_add_12_51_groupi_g16121(csa_tree_add_12_51_groupi_n_5652 ,csa_tree_add_12_51_groupi_n_5377 ,csa_tree_add_12_51_groupi_n_5584);
  and csa_tree_add_12_51_groupi_g16122(csa_tree_add_12_51_groupi_n_5651 ,csa_tree_add_12_51_groupi_n_5578 ,csa_tree_add_12_51_groupi_n_5474);
  or csa_tree_add_12_51_groupi_g16123(csa_tree_add_12_51_groupi_n_5650 ,csa_tree_add_12_51_groupi_n_5578 ,csa_tree_add_12_51_groupi_n_5474);
  and csa_tree_add_12_51_groupi_g16124(csa_tree_add_12_51_groupi_n_5649 ,csa_tree_add_12_51_groupi_n_5577 ,csa_tree_add_12_51_groupi_n_5376);
  xnor csa_tree_add_12_51_groupi_g16125(csa_tree_add_12_51_groupi_n_5648 ,csa_tree_add_12_51_groupi_n_5535 ,csa_tree_add_12_51_groupi_n_5509);
  xnor csa_tree_add_12_51_groupi_g16126(csa_tree_add_12_51_groupi_n_5647 ,csa_tree_add_12_51_groupi_n_5216 ,csa_tree_add_12_51_groupi_n_5511);
  xnor csa_tree_add_12_51_groupi_g16127(csa_tree_add_12_51_groupi_n_5646 ,csa_tree_add_12_51_groupi_n_5508 ,csa_tree_add_12_51_groupi_n_5181);
  xnor csa_tree_add_12_51_groupi_g16128(csa_tree_add_12_51_groupi_n_5645 ,csa_tree_add_12_51_groupi_n_5260 ,csa_tree_add_12_51_groupi_n_5500);
  xor csa_tree_add_12_51_groupi_g16129(csa_tree_add_12_51_groupi_n_5644 ,csa_tree_add_12_51_groupi_n_5415 ,csa_tree_add_12_51_groupi_n_5540);
  xnor csa_tree_add_12_51_groupi_g16130(csa_tree_add_12_51_groupi_n_5643 ,csa_tree_add_12_51_groupi_n_5506 ,csa_tree_add_12_51_groupi_n_5539);
  xor csa_tree_add_12_51_groupi_g16131(csa_tree_add_12_51_groupi_n_5642 ,csa_tree_add_12_51_groupi_n_5420 ,csa_tree_add_12_51_groupi_n_5543);
  xnor csa_tree_add_12_51_groupi_g16132(csa_tree_add_12_51_groupi_n_5678 ,csa_tree_add_12_51_groupi_n_4668 ,csa_tree_add_12_51_groupi_n_5480);
  xnor csa_tree_add_12_51_groupi_g16133(csa_tree_add_12_51_groupi_n_5677 ,csa_tree_add_12_51_groupi_n_5505 ,csa_tree_add_12_51_groupi_n_5481);
  xnor csa_tree_add_12_51_groupi_g16134(csa_tree_add_12_51_groupi_n_5676 ,csa_tree_add_12_51_groupi_n_5541 ,csa_tree_add_12_51_groupi_n_2570);
  not csa_tree_add_12_51_groupi_g16135(csa_tree_add_12_51_groupi_n_5640 ,csa_tree_add_12_51_groupi_n_5641);
  or csa_tree_add_12_51_groupi_g16136(csa_tree_add_12_51_groupi_n_5639 ,csa_tree_add_12_51_groupi_n_5433 ,csa_tree_add_12_51_groupi_n_5527);
  nor csa_tree_add_12_51_groupi_g16137(csa_tree_add_12_51_groupi_n_5638 ,csa_tree_add_12_51_groupi_n_5432 ,csa_tree_add_12_51_groupi_n_5525);
  or csa_tree_add_12_51_groupi_g16138(csa_tree_add_12_51_groupi_n_5637 ,csa_tree_add_12_51_groupi_n_5434 ,csa_tree_add_12_51_groupi_n_5524);
  nor csa_tree_add_12_51_groupi_g16139(csa_tree_add_12_51_groupi_n_5636 ,csa_tree_add_12_51_groupi_n_5436 ,csa_tree_add_12_51_groupi_n_5521);
  and csa_tree_add_12_51_groupi_g16140(csa_tree_add_12_51_groupi_n_5635 ,csa_tree_add_12_51_groupi_n_5519 ,csa_tree_add_12_51_groupi_n_5511);
  or csa_tree_add_12_51_groupi_g16141(csa_tree_add_12_51_groupi_n_5634 ,csa_tree_add_12_51_groupi_n_5516 ,csa_tree_add_12_51_groupi_n_5478);
  or csa_tree_add_12_51_groupi_g16142(csa_tree_add_12_51_groupi_n_5633 ,csa_tree_add_12_51_groupi_n_2437 ,csa_tree_add_12_51_groupi_n_5541);
  or csa_tree_add_12_51_groupi_g16143(csa_tree_add_12_51_groupi_n_5632 ,csa_tree_add_12_51_groupi_n_5515 ,csa_tree_add_12_51_groupi_n_5435);
  and csa_tree_add_12_51_groupi_g16144(csa_tree_add_12_51_groupi_n_5631 ,csa_tree_add_12_51_groupi_n_5385 ,csa_tree_add_12_51_groupi_n_5513);
  and csa_tree_add_12_51_groupi_g16145(csa_tree_add_12_51_groupi_n_5630 ,csa_tree_add_12_51_groupi_n_5260 ,csa_tree_add_12_51_groupi_n_5500);
  or csa_tree_add_12_51_groupi_g16146(csa_tree_add_12_51_groupi_n_5629 ,csa_tree_add_12_51_groupi_n_5260 ,csa_tree_add_12_51_groupi_n_5500);
  nor csa_tree_add_12_51_groupi_g16147(csa_tree_add_12_51_groupi_n_5628 ,csa_tree_add_12_51_groupi_n_5246 ,csa_tree_add_12_51_groupi_n_5505);
  or csa_tree_add_12_51_groupi_g16148(csa_tree_add_12_51_groupi_n_5627 ,csa_tree_add_12_51_groupi_n_5247 ,csa_tree_add_12_51_groupi_n_5504);
  and csa_tree_add_12_51_groupi_g16149(csa_tree_add_12_51_groupi_n_5626 ,csa_tree_add_12_51_groupi_n_5501 ,csa_tree_add_12_51_groupi_n_5219);
  nor csa_tree_add_12_51_groupi_g16150(csa_tree_add_12_51_groupi_n_5625 ,csa_tree_add_12_51_groupi_n_5501 ,csa_tree_add_12_51_groupi_n_5219);
  and csa_tree_add_12_51_groupi_g16151(csa_tree_add_12_51_groupi_n_5624 ,csa_tree_add_12_51_groupi_n_5479 ,csa_tree_add_12_51_groupi_n_5523);
  or csa_tree_add_12_51_groupi_g16152(csa_tree_add_12_51_groupi_n_5623 ,csa_tree_add_12_51_groupi_n_5507 ,csa_tree_add_12_51_groupi_n_5180);
  nor csa_tree_add_12_51_groupi_g16153(csa_tree_add_12_51_groupi_n_5622 ,csa_tree_add_12_51_groupi_n_5508 ,csa_tree_add_12_51_groupi_n_5181);
  or csa_tree_add_12_51_groupi_g16154(csa_tree_add_12_51_groupi_n_5621 ,csa_tree_add_12_51_groupi_n_5534 ,csa_tree_add_12_51_groupi_n_4841);
  nor csa_tree_add_12_51_groupi_g16155(csa_tree_add_12_51_groupi_n_5620 ,csa_tree_add_12_51_groupi_n_5535 ,csa_tree_add_12_51_groupi_n_4840);
  nor csa_tree_add_12_51_groupi_g16156(csa_tree_add_12_51_groupi_n_5619 ,csa_tree_add_12_51_groupi_n_1655 ,csa_tree_add_12_51_groupi_n_1007);
  nor csa_tree_add_12_51_groupi_g16157(csa_tree_add_12_51_groupi_n_5618 ,csa_tree_add_12_51_groupi_n_1583 ,csa_tree_add_12_51_groupi_n_1010);
  nor csa_tree_add_12_51_groupi_g16158(csa_tree_add_12_51_groupi_n_5617 ,csa_tree_add_12_51_groupi_n_1592 ,csa_tree_add_12_51_groupi_n_161);
  nor csa_tree_add_12_51_groupi_g16159(csa_tree_add_12_51_groupi_n_5616 ,csa_tree_add_12_51_groupi_n_1604 ,csa_tree_add_12_51_groupi_n_1007);
  nor csa_tree_add_12_51_groupi_g16160(csa_tree_add_12_51_groupi_n_5615 ,csa_tree_add_12_51_groupi_n_1640 ,csa_tree_add_12_51_groupi_n_1008);
  nor csa_tree_add_12_51_groupi_g16161(csa_tree_add_12_51_groupi_n_5614 ,csa_tree_add_12_51_groupi_n_1622 ,csa_tree_add_12_51_groupi_n_1011);
  nor csa_tree_add_12_51_groupi_g16162(csa_tree_add_12_51_groupi_n_5613 ,csa_tree_add_12_51_groupi_n_1616 ,csa_tree_add_12_51_groupi_n_930);
  nor csa_tree_add_12_51_groupi_g16163(csa_tree_add_12_51_groupi_n_5612 ,csa_tree_add_12_51_groupi_n_4095 ,csa_tree_add_12_51_groupi_n_5490);
  nor csa_tree_add_12_51_groupi_g16164(csa_tree_add_12_51_groupi_n_5611 ,csa_tree_add_12_51_groupi_n_3848 ,csa_tree_add_12_51_groupi_n_5489);
  nor csa_tree_add_12_51_groupi_g16165(csa_tree_add_12_51_groupi_n_5610 ,csa_tree_add_12_51_groupi_n_3847 ,csa_tree_add_12_51_groupi_n_5488);
  nor csa_tree_add_12_51_groupi_g16166(csa_tree_add_12_51_groupi_n_5609 ,csa_tree_add_12_51_groupi_n_3837 ,csa_tree_add_12_51_groupi_n_5487);
  nor csa_tree_add_12_51_groupi_g16167(csa_tree_add_12_51_groupi_n_5608 ,csa_tree_add_12_51_groupi_n_3830 ,csa_tree_add_12_51_groupi_n_5486);
  nor csa_tree_add_12_51_groupi_g16168(csa_tree_add_12_51_groupi_n_5607 ,csa_tree_add_12_51_groupi_n_4034 ,csa_tree_add_12_51_groupi_n_5494);
  nor csa_tree_add_12_51_groupi_g16169(csa_tree_add_12_51_groupi_n_5606 ,csa_tree_add_12_51_groupi_n_4106 ,csa_tree_add_12_51_groupi_n_5497);
  nor csa_tree_add_12_51_groupi_g16170(csa_tree_add_12_51_groupi_n_5605 ,csa_tree_add_12_51_groupi_n_4108 ,csa_tree_add_12_51_groupi_n_5495);
  nor csa_tree_add_12_51_groupi_g16171(csa_tree_add_12_51_groupi_n_5604 ,csa_tree_add_12_51_groupi_n_3459 ,csa_tree_add_12_51_groupi_n_5485);
  nor csa_tree_add_12_51_groupi_g16172(csa_tree_add_12_51_groupi_n_5603 ,csa_tree_add_12_51_groupi_n_3927 ,csa_tree_add_12_51_groupi_n_5493);
  nor csa_tree_add_12_51_groupi_g16173(csa_tree_add_12_51_groupi_n_5602 ,csa_tree_add_12_51_groupi_n_3448 ,csa_tree_add_12_51_groupi_n_5483);
  nor csa_tree_add_12_51_groupi_g16174(csa_tree_add_12_51_groupi_n_5601 ,csa_tree_add_12_51_groupi_n_4068 ,csa_tree_add_12_51_groupi_n_5496);
  nor csa_tree_add_12_51_groupi_g16175(csa_tree_add_12_51_groupi_n_5600 ,csa_tree_add_12_51_groupi_n_3444 ,csa_tree_add_12_51_groupi_n_5484);
  nor csa_tree_add_12_51_groupi_g16176(csa_tree_add_12_51_groupi_n_5599 ,csa_tree_add_12_51_groupi_n_3922 ,csa_tree_add_12_51_groupi_n_5492);
  nor csa_tree_add_12_51_groupi_g16177(csa_tree_add_12_51_groupi_n_5598 ,csa_tree_add_12_51_groupi_n_3890 ,csa_tree_add_12_51_groupi_n_5491);
  or csa_tree_add_12_51_groupi_g16178(csa_tree_add_12_51_groupi_n_5641 ,csa_tree_add_12_51_groupi_n_5463 ,csa_tree_add_12_51_groupi_n_5498);
  not csa_tree_add_12_51_groupi_g16179(csa_tree_add_12_51_groupi_n_5597 ,csa_tree_add_12_51_groupi_n_5596);
  not csa_tree_add_12_51_groupi_g16180(csa_tree_add_12_51_groupi_n_5591 ,csa_tree_add_12_51_groupi_n_5590);
  not csa_tree_add_12_51_groupi_g16181(csa_tree_add_12_51_groupi_n_5589 ,csa_tree_add_12_51_groupi_n_5588);
  not csa_tree_add_12_51_groupi_g16182(csa_tree_add_12_51_groupi_n_5584 ,csa_tree_add_12_51_groupi_n_5585);
  not csa_tree_add_12_51_groupi_g16183(csa_tree_add_12_51_groupi_n_5582 ,csa_tree_add_12_51_groupi_n_5583);
  not csa_tree_add_12_51_groupi_g16184(csa_tree_add_12_51_groupi_n_5574 ,csa_tree_add_12_51_groupi_n_5573);
  not csa_tree_add_12_51_groupi_g16185(csa_tree_add_12_51_groupi_n_5569 ,csa_tree_add_12_51_groupi_n_5570);
  not csa_tree_add_12_51_groupi_g16186(csa_tree_add_12_51_groupi_n_5568 ,csa_tree_add_12_51_groupi_n_5567);
  not csa_tree_add_12_51_groupi_g16187(csa_tree_add_12_51_groupi_n_5566 ,csa_tree_add_12_51_groupi_n_5565);
  not csa_tree_add_12_51_groupi_g16188(csa_tree_add_12_51_groupi_n_5563 ,csa_tree_add_12_51_groupi_n_5564);
  not csa_tree_add_12_51_groupi_g16189(csa_tree_add_12_51_groupi_n_5562 ,csa_tree_add_12_51_groupi_n_5561);
  nor csa_tree_add_12_51_groupi_g16190(csa_tree_add_12_51_groupi_n_5560 ,csa_tree_add_12_51_groupi_n_1634 ,csa_tree_add_12_51_groupi_n_929);
  nor csa_tree_add_12_51_groupi_g16191(csa_tree_add_12_51_groupi_n_5559 ,csa_tree_add_12_51_groupi_n_1664 ,csa_tree_add_12_51_groupi_n_1008);
  nor csa_tree_add_12_51_groupi_g16192(csa_tree_add_12_51_groupi_n_5558 ,csa_tree_add_12_51_groupi_n_1610 ,csa_tree_add_12_51_groupi_n_929);
  nor csa_tree_add_12_51_groupi_g16193(csa_tree_add_12_51_groupi_n_5557 ,csa_tree_add_12_51_groupi_n_1586 ,csa_tree_add_12_51_groupi_n_1011);
  nor csa_tree_add_12_51_groupi_g16194(csa_tree_add_12_51_groupi_n_5556 ,csa_tree_add_12_51_groupi_n_1646 ,csa_tree_add_12_51_groupi_n_1010);
  nor csa_tree_add_12_51_groupi_g16195(csa_tree_add_12_51_groupi_n_5555 ,csa_tree_add_12_51_groupi_n_1598 ,csa_tree_add_12_51_groupi_n_1974);
  nor csa_tree_add_12_51_groupi_g16196(csa_tree_add_12_51_groupi_n_5554 ,csa_tree_add_12_51_groupi_n_1679 ,csa_tree_add_12_51_groupi_n_930);
  nor csa_tree_add_12_51_groupi_g16197(csa_tree_add_12_51_groupi_n_5553 ,csa_tree_add_12_51_groupi_n_1628 ,csa_tree_add_12_51_groupi_n_161);
  xnor csa_tree_add_12_51_groupi_g16198(csa_tree_add_12_51_groupi_n_5552 ,csa_tree_add_12_51_groupi_n_5436 ,csa_tree_add_12_51_groupi_n_5411);
  xnor csa_tree_add_12_51_groupi_g16199(csa_tree_add_12_51_groupi_n_5551 ,csa_tree_add_12_51_groupi_n_5148 ,csa_tree_add_12_51_groupi_n_5425);
  xor csa_tree_add_12_51_groupi_g16200(csa_tree_add_12_51_groupi_n_5550 ,csa_tree_add_12_51_groupi_n_5431 ,csa_tree_add_12_51_groupi_n_5219);
  xnor csa_tree_add_12_51_groupi_g16201(csa_tree_add_12_51_groupi_n_5549 ,csa_tree_add_12_51_groupi_n_5255 ,csa_tree_add_12_51_groupi_n_5405);
  xnor csa_tree_add_12_51_groupi_g16202(csa_tree_add_12_51_groupi_n_5548 ,csa_tree_add_12_51_groupi_n_5375 ,csa_tree_add_12_51_groupi_n_5433);
  xnor csa_tree_add_12_51_groupi_g16203(csa_tree_add_12_51_groupi_n_5547 ,csa_tree_add_12_51_groupi_n_5478 ,csa_tree_add_12_51_groupi_n_5422);
  xnor csa_tree_add_12_51_groupi_g16204(csa_tree_add_12_51_groupi_n_5546 ,csa_tree_add_12_51_groupi_n_5432 ,csa_tree_add_12_51_groupi_n_5412);
  xnor csa_tree_add_12_51_groupi_g16205(csa_tree_add_12_51_groupi_n_5545 ,csa_tree_add_12_51_groupi_n_5477 ,csa_tree_add_12_51_groupi_n_5434);
  xnor csa_tree_add_12_51_groupi_g16206(csa_tree_add_12_51_groupi_n_5544 ,csa_tree_add_12_51_groupi_n_5214 ,csa_tree_add_12_51_groupi_n_5435);
  xnor csa_tree_add_12_51_groupi_g16207(csa_tree_add_12_51_groupi_n_5596 ,csa_tree_add_12_51_groupi_n_5450 ,in2[2]);
  xnor csa_tree_add_12_51_groupi_g16208(csa_tree_add_12_51_groupi_n_5595 ,csa_tree_add_12_51_groupi_n_1898 ,csa_tree_add_12_51_groupi_n_5442);
  xnor csa_tree_add_12_51_groupi_g16209(csa_tree_add_12_51_groupi_n_5594 ,csa_tree_add_12_51_groupi_n_96 ,csa_tree_add_12_51_groupi_n_5444);
  xnor csa_tree_add_12_51_groupi_g16210(csa_tree_add_12_51_groupi_n_5593 ,csa_tree_add_12_51_groupi_n_5451 ,in3[14]);
  xnor csa_tree_add_12_51_groupi_g16211(csa_tree_add_12_51_groupi_n_5592 ,csa_tree_add_12_51_groupi_n_1947 ,csa_tree_add_12_51_groupi_n_5440);
  xnor csa_tree_add_12_51_groupi_g16212(csa_tree_add_12_51_groupi_n_5590 ,csa_tree_add_12_51_groupi_n_5438 ,in3[11]);
  xnor csa_tree_add_12_51_groupi_g16213(csa_tree_add_12_51_groupi_n_5588 ,csa_tree_add_12_51_groupi_n_5445 ,in2[5]);
  xnor csa_tree_add_12_51_groupi_g16214(csa_tree_add_12_51_groupi_n_5587 ,csa_tree_add_12_51_groupi_n_115 ,csa_tree_add_12_51_groupi_n_5446);
  xnor csa_tree_add_12_51_groupi_g16215(csa_tree_add_12_51_groupi_n_5586 ,csa_tree_add_12_51_groupi_n_5269 ,csa_tree_add_12_51_groupi_n_5394);
  xnor csa_tree_add_12_51_groupi_g16216(csa_tree_add_12_51_groupi_n_5585 ,csa_tree_add_12_51_groupi_n_5252 ,csa_tree_add_12_51_groupi_n_5392);
  xnor csa_tree_add_12_51_groupi_g16217(csa_tree_add_12_51_groupi_n_5583 ,csa_tree_add_12_51_groupi_n_5274 ,csa_tree_add_12_51_groupi_n_5395);
  xnor csa_tree_add_12_51_groupi_g16218(csa_tree_add_12_51_groupi_n_5581 ,csa_tree_add_12_51_groupi_n_5350 ,csa_tree_add_12_51_groupi_n_5393);
  xnor csa_tree_add_12_51_groupi_g16219(csa_tree_add_12_51_groupi_n_5580 ,csa_tree_add_12_51_groupi_n_5351 ,csa_tree_add_12_51_groupi_n_5389);
  xnor csa_tree_add_12_51_groupi_g16220(csa_tree_add_12_51_groupi_n_5579 ,csa_tree_add_12_51_groupi_n_5271 ,csa_tree_add_12_51_groupi_n_5390);
  xnor csa_tree_add_12_51_groupi_g16221(csa_tree_add_12_51_groupi_n_5578 ,csa_tree_add_12_51_groupi_n_5272 ,csa_tree_add_12_51_groupi_n_5391);
  xnor csa_tree_add_12_51_groupi_g16222(csa_tree_add_12_51_groupi_n_5577 ,csa_tree_add_12_51_groupi_n_5273 ,csa_tree_add_12_51_groupi_n_5388);
  xnor csa_tree_add_12_51_groupi_g16223(csa_tree_add_12_51_groupi_n_5576 ,csa_tree_add_12_51_groupi_n_5347 ,csa_tree_add_12_51_groupi_n_5387);
  xnor csa_tree_add_12_51_groupi_g16224(csa_tree_add_12_51_groupi_n_5575 ,csa_tree_add_12_51_groupi_n_5447 ,in3[2]);
  xnor csa_tree_add_12_51_groupi_g16225(csa_tree_add_12_51_groupi_n_5573 ,csa_tree_add_12_51_groupi_n_5437 ,in3[5]);
  xnor csa_tree_add_12_51_groupi_g16226(csa_tree_add_12_51_groupi_n_5572 ,csa_tree_add_12_51_groupi_n_5248 ,csa_tree_add_12_51_groupi_n_5396);
  xnor csa_tree_add_12_51_groupi_g16227(csa_tree_add_12_51_groupi_n_5571 ,csa_tree_add_12_51_groupi_n_5383 ,csa_tree_add_12_51_groupi_n_5386);
  xnor csa_tree_add_12_51_groupi_g16228(csa_tree_add_12_51_groupi_n_5570 ,csa_tree_add_12_51_groupi_n_5448 ,in4[2]);
  xnor csa_tree_add_12_51_groupi_g16229(csa_tree_add_12_51_groupi_n_5567 ,csa_tree_add_12_51_groupi_n_5449 ,csa_tree_add_12_51_groupi_n_1936);
  xnor csa_tree_add_12_51_groupi_g16230(csa_tree_add_12_51_groupi_n_5565 ,csa_tree_add_12_51_groupi_n_5443 ,in4[14]);
  xnor csa_tree_add_12_51_groupi_g16231(csa_tree_add_12_51_groupi_n_5564 ,csa_tree_add_12_51_groupi_n_5439 ,in4[11]);
  xnor csa_tree_add_12_51_groupi_g16232(csa_tree_add_12_51_groupi_n_5561 ,csa_tree_add_12_51_groupi_n_5441 ,csa_tree_add_12_51_groupi_n_1939);
  not csa_tree_add_12_51_groupi_g16233(csa_tree_add_12_51_groupi_n_5537 ,csa_tree_add_12_51_groupi_n_5536);
  not csa_tree_add_12_51_groupi_g16234(csa_tree_add_12_51_groupi_n_5534 ,csa_tree_add_12_51_groupi_n_5535);
  not csa_tree_add_12_51_groupi_g16235(csa_tree_add_12_51_groupi_n_5532 ,csa_tree_add_12_51_groupi_n_5533);
  not csa_tree_add_12_51_groupi_g16236(csa_tree_add_12_51_groupi_n_5530 ,csa_tree_add_12_51_groupi_n_5531);
  and csa_tree_add_12_51_groupi_g16237(csa_tree_add_12_51_groupi_n_5529 ,csa_tree_add_12_51_groupi_n_5148 ,csa_tree_add_12_51_groupi_n_5425);
  or csa_tree_add_12_51_groupi_g16238(csa_tree_add_12_51_groupi_n_5528 ,csa_tree_add_12_51_groupi_n_5416 ,csa_tree_add_12_51_groupi_n_5375);
  nor csa_tree_add_12_51_groupi_g16239(csa_tree_add_12_51_groupi_n_5527 ,csa_tree_add_12_51_groupi_n_5417 ,csa_tree_add_12_51_groupi_n_5374);
  nor csa_tree_add_12_51_groupi_g16240(csa_tree_add_12_51_groupi_n_5526 ,csa_tree_add_12_51_groupi_n_5419 ,csa_tree_add_12_51_groupi_n_5412);
  and csa_tree_add_12_51_groupi_g16241(csa_tree_add_12_51_groupi_n_5525 ,csa_tree_add_12_51_groupi_n_5419 ,csa_tree_add_12_51_groupi_n_5412);
  nor csa_tree_add_12_51_groupi_g16242(csa_tree_add_12_51_groupi_n_5524 ,csa_tree_add_12_51_groupi_n_5427 ,csa_tree_add_12_51_groupi_n_5476);
  or csa_tree_add_12_51_groupi_g16243(csa_tree_add_12_51_groupi_n_5523 ,csa_tree_add_12_51_groupi_n_5148 ,csa_tree_add_12_51_groupi_n_5425);
  nor csa_tree_add_12_51_groupi_g16244(csa_tree_add_12_51_groupi_n_5522 ,csa_tree_add_12_51_groupi_n_5410 ,csa_tree_add_12_51_groupi_n_5411);
  and csa_tree_add_12_51_groupi_g16245(csa_tree_add_12_51_groupi_n_5521 ,csa_tree_add_12_51_groupi_n_5410 ,csa_tree_add_12_51_groupi_n_5411);
  and csa_tree_add_12_51_groupi_g16246(csa_tree_add_12_51_groupi_n_5520 ,csa_tree_add_12_51_groupi_n_5216 ,csa_tree_add_12_51_groupi_n_5428);
  or csa_tree_add_12_51_groupi_g16247(csa_tree_add_12_51_groupi_n_5519 ,csa_tree_add_12_51_groupi_n_5216 ,csa_tree_add_12_51_groupi_n_5428);
  or csa_tree_add_12_51_groupi_g16248(csa_tree_add_12_51_groupi_n_5518 ,csa_tree_add_12_51_groupi_n_5426 ,csa_tree_add_12_51_groupi_n_5477);
  or csa_tree_add_12_51_groupi_g16249(csa_tree_add_12_51_groupi_n_5517 ,csa_tree_add_12_51_groupi_n_5422 ,csa_tree_add_12_51_groupi_n_5423);
  nor csa_tree_add_12_51_groupi_g16250(csa_tree_add_12_51_groupi_n_5516 ,csa_tree_add_12_51_groupi_n_5421 ,csa_tree_add_12_51_groupi_n_5424);
  nor csa_tree_add_12_51_groupi_g16251(csa_tree_add_12_51_groupi_n_5515 ,csa_tree_add_12_51_groupi_n_5214 ,csa_tree_add_12_51_groupi_n_5414);
  or csa_tree_add_12_51_groupi_g16252(csa_tree_add_12_51_groupi_n_5514 ,csa_tree_add_12_51_groupi_n_5213 ,csa_tree_add_12_51_groupi_n_5413);
  or csa_tree_add_12_51_groupi_g16253(csa_tree_add_12_51_groupi_n_5513 ,csa_tree_add_12_51_groupi_n_5255 ,csa_tree_add_12_51_groupi_n_5405);
  and csa_tree_add_12_51_groupi_g16254(csa_tree_add_12_51_groupi_n_5512 ,csa_tree_add_12_51_groupi_n_5255 ,csa_tree_add_12_51_groupi_n_5405);
  and csa_tree_add_12_51_groupi_g16255(csa_tree_add_12_51_groupi_n_5543 ,csa_tree_add_12_51_groupi_n_5370 ,csa_tree_add_12_51_groupi_n_5459);
  or csa_tree_add_12_51_groupi_g16256(csa_tree_add_12_51_groupi_n_5542 ,csa_tree_add_12_51_groupi_n_5369 ,csa_tree_add_12_51_groupi_n_5457);
  and csa_tree_add_12_51_groupi_g16257(csa_tree_add_12_51_groupi_n_5541 ,csa_tree_add_12_51_groupi_n_2423 ,csa_tree_add_12_51_groupi_n_5455);
  and csa_tree_add_12_51_groupi_g16258(csa_tree_add_12_51_groupi_n_5540 ,csa_tree_add_12_51_groupi_n_5372 ,csa_tree_add_12_51_groupi_n_5465);
  and csa_tree_add_12_51_groupi_g16259(csa_tree_add_12_51_groupi_n_5539 ,csa_tree_add_12_51_groupi_n_5368 ,csa_tree_add_12_51_groupi_n_5461);
  or csa_tree_add_12_51_groupi_g16260(csa_tree_add_12_51_groupi_n_5538 ,csa_tree_add_12_51_groupi_n_5356 ,csa_tree_add_12_51_groupi_n_5452);
  or csa_tree_add_12_51_groupi_g16261(csa_tree_add_12_51_groupi_n_5536 ,csa_tree_add_12_51_groupi_n_5353 ,csa_tree_add_12_51_groupi_n_5453);
  or csa_tree_add_12_51_groupi_g16262(csa_tree_add_12_51_groupi_n_5535 ,csa_tree_add_12_51_groupi_n_5362 ,csa_tree_add_12_51_groupi_n_5456);
  or csa_tree_add_12_51_groupi_g16263(csa_tree_add_12_51_groupi_n_5533 ,csa_tree_add_12_51_groupi_n_5357 ,csa_tree_add_12_51_groupi_n_5454);
  or csa_tree_add_12_51_groupi_g16264(csa_tree_add_12_51_groupi_n_5531 ,csa_tree_add_12_51_groupi_n_5363 ,csa_tree_add_12_51_groupi_n_5458);
  not csa_tree_add_12_51_groupi_g16265(csa_tree_add_12_51_groupi_n_5510 ,csa_tree_add_12_51_groupi_n_5509);
  not csa_tree_add_12_51_groupi_g16266(csa_tree_add_12_51_groupi_n_5507 ,csa_tree_add_12_51_groupi_n_5508);
  not csa_tree_add_12_51_groupi_g16267(csa_tree_add_12_51_groupi_n_5504 ,csa_tree_add_12_51_groupi_n_5505);
  not csa_tree_add_12_51_groupi_g16268(csa_tree_add_12_51_groupi_n_5502 ,csa_tree_add_12_51_groupi_n_5503);
  nor csa_tree_add_12_51_groupi_g16269(csa_tree_add_12_51_groupi_n_5498 ,csa_tree_add_12_51_groupi_n_5464 ,csa_tree_add_12_51_groupi_n_5318);
  or csa_tree_add_12_51_groupi_g16270(csa_tree_add_12_51_groupi_n_5497 ,csa_tree_add_12_51_groupi_n_3372 ,csa_tree_add_12_51_groupi_n_5470);
  or csa_tree_add_12_51_groupi_g16271(csa_tree_add_12_51_groupi_n_5496 ,csa_tree_add_12_51_groupi_n_3496 ,csa_tree_add_12_51_groupi_n_5471);
  or csa_tree_add_12_51_groupi_g16272(csa_tree_add_12_51_groupi_n_5495 ,csa_tree_add_12_51_groupi_n_3302 ,csa_tree_add_12_51_groupi_n_5400);
  or csa_tree_add_12_51_groupi_g16273(csa_tree_add_12_51_groupi_n_5494 ,csa_tree_add_12_51_groupi_n_3298 ,csa_tree_add_12_51_groupi_n_5404);
  or csa_tree_add_12_51_groupi_g16274(csa_tree_add_12_51_groupi_n_5493 ,csa_tree_add_12_51_groupi_n_3677 ,csa_tree_add_12_51_groupi_n_5469);
  or csa_tree_add_12_51_groupi_g16275(csa_tree_add_12_51_groupi_n_5492 ,csa_tree_add_12_51_groupi_n_3666 ,csa_tree_add_12_51_groupi_n_5472);
  or csa_tree_add_12_51_groupi_g16276(csa_tree_add_12_51_groupi_n_5491 ,csa_tree_add_12_51_groupi_n_3615 ,csa_tree_add_12_51_groupi_n_5397);
  or csa_tree_add_12_51_groupi_g16277(csa_tree_add_12_51_groupi_n_5490 ,csa_tree_add_12_51_groupi_n_3097 ,csa_tree_add_12_51_groupi_n_5403);
  or csa_tree_add_12_51_groupi_g16278(csa_tree_add_12_51_groupi_n_5489 ,csa_tree_add_12_51_groupi_n_3583 ,csa_tree_add_12_51_groupi_n_5402);
  or csa_tree_add_12_51_groupi_g16279(csa_tree_add_12_51_groupi_n_5488 ,csa_tree_add_12_51_groupi_n_3661 ,csa_tree_add_12_51_groupi_n_5401);
  or csa_tree_add_12_51_groupi_g16280(csa_tree_add_12_51_groupi_n_5487 ,csa_tree_add_12_51_groupi_n_3735 ,csa_tree_add_12_51_groupi_n_5399);
  or csa_tree_add_12_51_groupi_g16281(csa_tree_add_12_51_groupi_n_5486 ,csa_tree_add_12_51_groupi_n_3613 ,csa_tree_add_12_51_groupi_n_5398);
  or csa_tree_add_12_51_groupi_g16282(csa_tree_add_12_51_groupi_n_5485 ,csa_tree_add_12_51_groupi_n_3099 ,csa_tree_add_12_51_groupi_n_5466);
  or csa_tree_add_12_51_groupi_g16283(csa_tree_add_12_51_groupi_n_5484 ,csa_tree_add_12_51_groupi_n_3035 ,csa_tree_add_12_51_groupi_n_5467);
  or csa_tree_add_12_51_groupi_g16284(csa_tree_add_12_51_groupi_n_5483 ,csa_tree_add_12_51_groupi_n_3110 ,csa_tree_add_12_51_groupi_n_5468);
  xnor csa_tree_add_12_51_groupi_g16285(out3[4] ,csa_tree_add_12_51_groupi_n_5316 ,csa_tree_add_12_51_groupi_n_5322);
  xnor csa_tree_add_12_51_groupi_g16286(csa_tree_add_12_51_groupi_n_5481 ,csa_tree_add_12_51_groupi_n_5381 ,csa_tree_add_12_51_groupi_n_5247);
  xnor csa_tree_add_12_51_groupi_g16287(csa_tree_add_12_51_groupi_n_5480 ,csa_tree_add_12_51_groupi_n_4714 ,csa_tree_add_12_51_groupi_n_5380);
  xnor csa_tree_add_12_51_groupi_g16288(csa_tree_add_12_51_groupi_n_5511 ,csa_tree_add_12_51_groupi_n_5187 ,csa_tree_add_12_51_groupi_n_5321);
  or csa_tree_add_12_51_groupi_g16289(csa_tree_add_12_51_groupi_n_5509 ,csa_tree_add_12_51_groupi_n_4795 ,csa_tree_add_12_51_groupi_n_5460);
  xnor csa_tree_add_12_51_groupi_g16290(csa_tree_add_12_51_groupi_n_5508 ,csa_tree_add_12_51_groupi_n_5086 ,csa_tree_add_12_51_groupi_n_5323);
  and csa_tree_add_12_51_groupi_g16291(csa_tree_add_12_51_groupi_n_5506 ,csa_tree_add_12_51_groupi_n_5343 ,csa_tree_add_12_51_groupi_n_5462);
  xnor csa_tree_add_12_51_groupi_g16292(csa_tree_add_12_51_groupi_n_5505 ,csa_tree_add_12_51_groupi_n_5105 ,csa_tree_add_12_51_groupi_n_5324);
  xnor csa_tree_add_12_51_groupi_g16293(csa_tree_add_12_51_groupi_n_5503 ,csa_tree_add_12_51_groupi_n_4678 ,csa_tree_add_12_51_groupi_n_5325);
  xnor csa_tree_add_12_51_groupi_g16294(csa_tree_add_12_51_groupi_n_5501 ,csa_tree_add_12_51_groupi_n_5098 ,csa_tree_add_12_51_groupi_n_5320);
  xnor csa_tree_add_12_51_groupi_g16295(csa_tree_add_12_51_groupi_n_5500 ,csa_tree_add_12_51_groupi_n_5110 ,csa_tree_add_12_51_groupi_n_5319);
  xnor csa_tree_add_12_51_groupi_g16296(csa_tree_add_12_51_groupi_n_5499 ,csa_tree_add_12_51_groupi_n_5382 ,csa_tree_add_12_51_groupi_n_2567);
  not csa_tree_add_12_51_groupi_g16297(csa_tree_add_12_51_groupi_n_5477 ,csa_tree_add_12_51_groupi_n_5476);
  nor csa_tree_add_12_51_groupi_g16298(csa_tree_add_12_51_groupi_n_5472 ,csa_tree_add_12_51_groupi_n_1823 ,csa_tree_add_12_51_groupi_n_1001);
  nor csa_tree_add_12_51_groupi_g16299(csa_tree_add_12_51_groupi_n_5471 ,csa_tree_add_12_51_groupi_n_1817 ,csa_tree_add_12_51_groupi_n_1004);
  nor csa_tree_add_12_51_groupi_g16300(csa_tree_add_12_51_groupi_n_5470 ,csa_tree_add_12_51_groupi_n_1829 ,csa_tree_add_12_51_groupi_n_153);
  nor csa_tree_add_12_51_groupi_g16301(csa_tree_add_12_51_groupi_n_5469 ,csa_tree_add_12_51_groupi_n_1827 ,csa_tree_add_12_51_groupi_n_1001);
  nor csa_tree_add_12_51_groupi_g16302(csa_tree_add_12_51_groupi_n_5468 ,csa_tree_add_12_51_groupi_n_1819 ,csa_tree_add_12_51_groupi_n_1002);
  nor csa_tree_add_12_51_groupi_g16303(csa_tree_add_12_51_groupi_n_5467 ,csa_tree_add_12_51_groupi_n_1825 ,csa_tree_add_12_51_groupi_n_1005);
  nor csa_tree_add_12_51_groupi_g16304(csa_tree_add_12_51_groupi_n_5466 ,csa_tree_add_12_51_groupi_n_1821 ,csa_tree_add_12_51_groupi_n_948);
  or csa_tree_add_12_51_groupi_g16305(csa_tree_add_12_51_groupi_n_5465 ,csa_tree_add_12_51_groupi_n_5371 ,csa_tree_add_12_51_groupi_n_5154);
  nor csa_tree_add_12_51_groupi_g16306(csa_tree_add_12_51_groupi_n_5464 ,csa_tree_add_12_51_groupi_n_5261 ,csa_tree_add_12_51_groupi_n_5347);
  and csa_tree_add_12_51_groupi_g16307(csa_tree_add_12_51_groupi_n_5463 ,csa_tree_add_12_51_groupi_n_5261 ,csa_tree_add_12_51_groupi_n_5347);
  or csa_tree_add_12_51_groupi_g16308(csa_tree_add_12_51_groupi_n_5462 ,csa_tree_add_12_51_groupi_n_5384 ,csa_tree_add_12_51_groupi_n_5342);
  or csa_tree_add_12_51_groupi_g16309(csa_tree_add_12_51_groupi_n_5461 ,csa_tree_add_12_51_groupi_n_5275 ,csa_tree_add_12_51_groupi_n_5366);
  and csa_tree_add_12_51_groupi_g16310(csa_tree_add_12_51_groupi_n_5460 ,csa_tree_add_12_51_groupi_n_5380 ,csa_tree_add_12_51_groupi_n_4796);
  or csa_tree_add_12_51_groupi_g16311(csa_tree_add_12_51_groupi_n_5459 ,csa_tree_add_12_51_groupi_n_5270 ,csa_tree_add_12_51_groupi_n_5329);
  and csa_tree_add_12_51_groupi_g16312(csa_tree_add_12_51_groupi_n_5458 ,csa_tree_add_12_51_groupi_n_5271 ,csa_tree_add_12_51_groupi_n_5365);
  and csa_tree_add_12_51_groupi_g16313(csa_tree_add_12_51_groupi_n_5457 ,csa_tree_add_12_51_groupi_n_5272 ,csa_tree_add_12_51_groupi_n_5360);
  nor csa_tree_add_12_51_groupi_g16314(csa_tree_add_12_51_groupi_n_5456 ,csa_tree_add_12_51_groupi_n_2 ,csa_tree_add_12_51_groupi_n_5361);
  or csa_tree_add_12_51_groupi_g16315(csa_tree_add_12_51_groupi_n_5455 ,csa_tree_add_12_51_groupi_n_2432 ,csa_tree_add_12_51_groupi_n_5382);
  and csa_tree_add_12_51_groupi_g16316(csa_tree_add_12_51_groupi_n_5454 ,csa_tree_add_12_51_groupi_n_5351 ,csa_tree_add_12_51_groupi_n_5359);
  and csa_tree_add_12_51_groupi_g16317(csa_tree_add_12_51_groupi_n_5453 ,csa_tree_add_12_51_groupi_n_5352 ,csa_tree_add_12_51_groupi_n_5350);
  and csa_tree_add_12_51_groupi_g16318(csa_tree_add_12_51_groupi_n_5452 ,csa_tree_add_12_51_groupi_n_5273 ,csa_tree_add_12_51_groupi_n_5354);
  nor csa_tree_add_12_51_groupi_g16319(csa_tree_add_12_51_groupi_n_5451 ,csa_tree_add_12_51_groupi_n_3876 ,csa_tree_add_12_51_groupi_n_5334);
  nor csa_tree_add_12_51_groupi_g16320(csa_tree_add_12_51_groupi_n_5450 ,csa_tree_add_12_51_groupi_n_3469 ,csa_tree_add_12_51_groupi_n_5327);
  nor csa_tree_add_12_51_groupi_g16321(csa_tree_add_12_51_groupi_n_5449 ,csa_tree_add_12_51_groupi_n_3880 ,csa_tree_add_12_51_groupi_n_5335);
  nor csa_tree_add_12_51_groupi_g16322(csa_tree_add_12_51_groupi_n_5448 ,csa_tree_add_12_51_groupi_n_3445 ,csa_tree_add_12_51_groupi_n_5328);
  nor csa_tree_add_12_51_groupi_g16323(csa_tree_add_12_51_groupi_n_5447 ,csa_tree_add_12_51_groupi_n_3446 ,csa_tree_add_12_51_groupi_n_5341);
  nor csa_tree_add_12_51_groupi_g16324(csa_tree_add_12_51_groupi_n_5446 ,csa_tree_add_12_51_groupi_n_4100 ,csa_tree_add_12_51_groupi_n_5336);
  nor csa_tree_add_12_51_groupi_g16325(csa_tree_add_12_51_groupi_n_5445 ,csa_tree_add_12_51_groupi_n_3879 ,csa_tree_add_12_51_groupi_n_5333);
  nor csa_tree_add_12_51_groupi_g16326(csa_tree_add_12_51_groupi_n_5444 ,csa_tree_add_12_51_groupi_n_3865 ,csa_tree_add_12_51_groupi_n_5331);
  nor csa_tree_add_12_51_groupi_g16327(csa_tree_add_12_51_groupi_n_5443 ,csa_tree_add_12_51_groupi_n_3915 ,csa_tree_add_12_51_groupi_n_5340);
  nor csa_tree_add_12_51_groupi_g16328(csa_tree_add_12_51_groupi_n_5442 ,csa_tree_add_12_51_groupi_n_3908 ,csa_tree_add_12_51_groupi_n_5339);
  nor csa_tree_add_12_51_groupi_g16329(csa_tree_add_12_51_groupi_n_5441 ,csa_tree_add_12_51_groupi_n_3917 ,csa_tree_add_12_51_groupi_n_5337);
  nor csa_tree_add_12_51_groupi_g16330(csa_tree_add_12_51_groupi_n_5440 ,csa_tree_add_12_51_groupi_n_3841 ,csa_tree_add_12_51_groupi_n_5345);
  nor csa_tree_add_12_51_groupi_g16331(csa_tree_add_12_51_groupi_n_5439 ,csa_tree_add_12_51_groupi_n_3845 ,csa_tree_add_12_51_groupi_n_5330);
  nor csa_tree_add_12_51_groupi_g16332(csa_tree_add_12_51_groupi_n_5438 ,csa_tree_add_12_51_groupi_n_3850 ,csa_tree_add_12_51_groupi_n_5332);
  nor csa_tree_add_12_51_groupi_g16333(csa_tree_add_12_51_groupi_n_5437 ,csa_tree_add_12_51_groupi_n_3920 ,csa_tree_add_12_51_groupi_n_5338);
  or csa_tree_add_12_51_groupi_g16334(csa_tree_add_12_51_groupi_n_5479 ,csa_tree_add_12_51_groupi_n_5296 ,csa_tree_add_12_51_groupi_n_5344);
  and csa_tree_add_12_51_groupi_g16335(csa_tree_add_12_51_groupi_n_5478 ,csa_tree_add_12_51_groupi_n_5302 ,csa_tree_add_12_51_groupi_n_5355);
  or csa_tree_add_12_51_groupi_g16336(csa_tree_add_12_51_groupi_n_5476 ,csa_tree_add_12_51_groupi_n_5300 ,csa_tree_add_12_51_groupi_n_5367);
  or csa_tree_add_12_51_groupi_g16337(csa_tree_add_12_51_groupi_n_5475 ,csa_tree_add_12_51_groupi_n_5212 ,csa_tree_add_12_51_groupi_n_5373);
  or csa_tree_add_12_51_groupi_g16338(csa_tree_add_12_51_groupi_n_5474 ,csa_tree_add_12_51_groupi_n_5306 ,csa_tree_add_12_51_groupi_n_5358);
  or csa_tree_add_12_51_groupi_g16339(csa_tree_add_12_51_groupi_n_5473 ,csa_tree_add_12_51_groupi_n_5311 ,csa_tree_add_12_51_groupi_n_5364);
  not csa_tree_add_12_51_groupi_g16340(csa_tree_add_12_51_groupi_n_5430 ,csa_tree_add_12_51_groupi_n_5429);
  not csa_tree_add_12_51_groupi_g16341(csa_tree_add_12_51_groupi_n_5426 ,csa_tree_add_12_51_groupi_n_5427);
  not csa_tree_add_12_51_groupi_g16342(csa_tree_add_12_51_groupi_n_5424 ,csa_tree_add_12_51_groupi_n_5423);
  not csa_tree_add_12_51_groupi_g16343(csa_tree_add_12_51_groupi_n_5422 ,csa_tree_add_12_51_groupi_n_5421);
  not csa_tree_add_12_51_groupi_g16344(csa_tree_add_12_51_groupi_n_5419 ,csa_tree_add_12_51_groupi_n_5418);
  not csa_tree_add_12_51_groupi_g16345(csa_tree_add_12_51_groupi_n_5417 ,csa_tree_add_12_51_groupi_n_5416);
  not csa_tree_add_12_51_groupi_g16346(csa_tree_add_12_51_groupi_n_5413 ,csa_tree_add_12_51_groupi_n_5414);
  not csa_tree_add_12_51_groupi_g16347(csa_tree_add_12_51_groupi_n_5410 ,csa_tree_add_12_51_groupi_n_5409);
  not csa_tree_add_12_51_groupi_g16348(csa_tree_add_12_51_groupi_n_5407 ,csa_tree_add_12_51_groupi_n_5408);
  nor csa_tree_add_12_51_groupi_g16349(csa_tree_add_12_51_groupi_n_5404 ,csa_tree_add_12_51_groupi_n_1837 ,csa_tree_add_12_51_groupi_n_947);
  nor csa_tree_add_12_51_groupi_g16350(csa_tree_add_12_51_groupi_n_5403 ,csa_tree_add_12_51_groupi_n_1841 ,csa_tree_add_12_51_groupi_n_1002);
  nor csa_tree_add_12_51_groupi_g16351(csa_tree_add_12_51_groupi_n_5402 ,csa_tree_add_12_51_groupi_n_1835 ,csa_tree_add_12_51_groupi_n_947);
  nor csa_tree_add_12_51_groupi_g16352(csa_tree_add_12_51_groupi_n_5401 ,csa_tree_add_12_51_groupi_n_1845 ,csa_tree_add_12_51_groupi_n_1005);
  nor csa_tree_add_12_51_groupi_g16353(csa_tree_add_12_51_groupi_n_5400 ,csa_tree_add_12_51_groupi_n_1839 ,csa_tree_add_12_51_groupi_n_1004);
  nor csa_tree_add_12_51_groupi_g16354(csa_tree_add_12_51_groupi_n_5399 ,csa_tree_add_12_51_groupi_n_1843 ,csa_tree_add_12_51_groupi_n_1971);
  nor csa_tree_add_12_51_groupi_g16355(csa_tree_add_12_51_groupi_n_5398 ,csa_tree_add_12_51_groupi_n_1833 ,csa_tree_add_12_51_groupi_n_948);
  nor csa_tree_add_12_51_groupi_g16356(csa_tree_add_12_51_groupi_n_5397 ,csa_tree_add_12_51_groupi_n_1831 ,csa_tree_add_12_51_groupi_n_153);
  xnor csa_tree_add_12_51_groupi_g16357(csa_tree_add_12_51_groupi_n_5396 ,csa_tree_add_12_51_groupi_n_2 ,csa_tree_add_12_51_groupi_n_5250);
  xnor csa_tree_add_12_51_groupi_g16358(csa_tree_add_12_51_groupi_n_5395 ,csa_tree_add_12_51_groupi_n_5259 ,csa_tree_add_12_51_groupi_n_5100);
  xnor csa_tree_add_12_51_groupi_g16359(csa_tree_add_12_51_groupi_n_5394 ,csa_tree_add_12_51_groupi_n_5262 ,csa_tree_add_12_51_groupi_n_5150);
  xnor csa_tree_add_12_51_groupi_g16360(csa_tree_add_12_51_groupi_n_5393 ,csa_tree_add_12_51_groupi_n_5054 ,csa_tree_add_12_51_groupi_n_5268);
  xnor csa_tree_add_12_51_groupi_g16361(csa_tree_add_12_51_groupi_n_5392 ,csa_tree_add_12_51_groupi_n_5154 ,csa_tree_add_12_51_groupi_n_5265);
  xnor csa_tree_add_12_51_groupi_g16362(csa_tree_add_12_51_groupi_n_5391 ,csa_tree_add_12_51_groupi_n_5245 ,csa_tree_add_12_51_groupi_n_5147);
  xnor csa_tree_add_12_51_groupi_g16363(csa_tree_add_12_51_groupi_n_5390 ,csa_tree_add_12_51_groupi_n_5052 ,csa_tree_add_12_51_groupi_n_5266);
  xnor csa_tree_add_12_51_groupi_g16364(csa_tree_add_12_51_groupi_n_5389 ,csa_tree_add_12_51_groupi_n_5053 ,csa_tree_add_12_51_groupi_n_5267);
  xnor csa_tree_add_12_51_groupi_g16365(csa_tree_add_12_51_groupi_n_5388 ,csa_tree_add_12_51_groupi_n_5055 ,csa_tree_add_12_51_groupi_n_5263);
  xnor csa_tree_add_12_51_groupi_g16366(csa_tree_add_12_51_groupi_n_5387 ,csa_tree_add_12_51_groupi_n_5261 ,csa_tree_add_12_51_groupi_n_5318);
  xnor csa_tree_add_12_51_groupi_g16367(csa_tree_add_12_51_groupi_n_5386 ,csa_tree_add_12_51_groupi_n_5254 ,csa_tree_add_12_51_groupi_n_5257);
  xnor csa_tree_add_12_51_groupi_g16368(csa_tree_add_12_51_groupi_n_5436 ,csa_tree_add_12_51_groupi_n_1929 ,csa_tree_add_12_51_groupi_n_5290);
  xnor csa_tree_add_12_51_groupi_g16369(csa_tree_add_12_51_groupi_n_5435 ,csa_tree_add_12_51_groupi_n_5221 ,csa_tree_add_12_51_groupi_n_5224);
  xnor csa_tree_add_12_51_groupi_g16370(csa_tree_add_12_51_groupi_n_5434 ,csa_tree_add_12_51_groupi_n_102 ,csa_tree_add_12_51_groupi_n_5284);
  xnor csa_tree_add_12_51_groupi_g16371(csa_tree_add_12_51_groupi_n_5433 ,csa_tree_add_12_51_groupi_n_1903 ,csa_tree_add_12_51_groupi_n_5280);
  xnor csa_tree_add_12_51_groupi_g16372(csa_tree_add_12_51_groupi_n_5432 ,csa_tree_add_12_51_groupi_n_1892 ,csa_tree_add_12_51_groupi_n_5288);
  xnor csa_tree_add_12_51_groupi_g16373(csa_tree_add_12_51_groupi_n_5431 ,csa_tree_add_12_51_groupi_n_5223 ,csa_tree_add_12_51_groupi_n_5230);
  xnor csa_tree_add_12_51_groupi_g16374(csa_tree_add_12_51_groupi_n_5429 ,csa_tree_add_12_51_groupi_n_5317 ,csa_tree_add_12_51_groupi_n_5228);
  xnor csa_tree_add_12_51_groupi_g16375(csa_tree_add_12_51_groupi_n_5428 ,csa_tree_add_12_51_groupi_n_5109 ,csa_tree_add_12_51_groupi_n_5229);
  xnor csa_tree_add_12_51_groupi_g16376(csa_tree_add_12_51_groupi_n_5427 ,csa_tree_add_12_51_groupi_n_5278 ,in4[2]);
  xnor csa_tree_add_12_51_groupi_g16377(csa_tree_add_12_51_groupi_n_5425 ,csa_tree_add_12_51_groupi_n_5111 ,csa_tree_add_12_51_groupi_n_5226);
  xnor csa_tree_add_12_51_groupi_g16378(csa_tree_add_12_51_groupi_n_5423 ,csa_tree_add_12_51_groupi_n_1923 ,csa_tree_add_12_51_groupi_n_5285);
  xnor csa_tree_add_12_51_groupi_g16379(csa_tree_add_12_51_groupi_n_5421 ,csa_tree_add_12_51_groupi_n_5286 ,in4[8]);
  xnor csa_tree_add_12_51_groupi_g16380(csa_tree_add_12_51_groupi_n_5420 ,csa_tree_add_12_51_groupi_n_5283 ,in3[8]);
  xnor csa_tree_add_12_51_groupi_g16381(csa_tree_add_12_51_groupi_n_5418 ,csa_tree_add_12_51_groupi_n_5289 ,in4[11]);
  xnor csa_tree_add_12_51_groupi_g16382(csa_tree_add_12_51_groupi_n_5416 ,csa_tree_add_12_51_groupi_n_5282 ,csa_tree_add_12_51_groupi_n_1935);
  xnor csa_tree_add_12_51_groupi_g16383(csa_tree_add_12_51_groupi_n_5415 ,csa_tree_add_12_51_groupi_n_5279 ,in2[5]);
  xnor csa_tree_add_12_51_groupi_g16384(csa_tree_add_12_51_groupi_n_5414 ,csa_tree_add_12_51_groupi_n_5107 ,csa_tree_add_12_51_groupi_n_5231);
  xnor csa_tree_add_12_51_groupi_g16385(csa_tree_add_12_51_groupi_n_5412 ,csa_tree_add_12_51_groupi_n_1921 ,csa_tree_add_12_51_groupi_n_5287);
  xnor csa_tree_add_12_51_groupi_g16386(csa_tree_add_12_51_groupi_n_5411 ,csa_tree_add_12_51_groupi_n_1898 ,csa_tree_add_12_51_groupi_n_5276);
  xnor csa_tree_add_12_51_groupi_g16387(csa_tree_add_12_51_groupi_n_5409 ,csa_tree_add_12_51_groupi_n_5281 ,in4[14]);
  xnor csa_tree_add_12_51_groupi_g16388(csa_tree_add_12_51_groupi_n_5408 ,csa_tree_add_12_51_groupi_n_5112 ,csa_tree_add_12_51_groupi_n_5225);
  xnor csa_tree_add_12_51_groupi_g16389(csa_tree_add_12_51_groupi_n_5406 ,csa_tree_add_12_51_groupi_n_5277 ,in2[2]);
  xnor csa_tree_add_12_51_groupi_g16390(csa_tree_add_12_51_groupi_n_5405 ,csa_tree_add_12_51_groupi_n_5108 ,csa_tree_add_12_51_groupi_n_5227);
  not csa_tree_add_12_51_groupi_g16391(csa_tree_add_12_51_groupi_n_5384 ,csa_tree_add_12_51_groupi_n_5383);
  not csa_tree_add_12_51_groupi_g16392(csa_tree_add_12_51_groupi_n_5377 ,csa_tree_add_12_51_groupi_n_5378);
  not csa_tree_add_12_51_groupi_g16393(csa_tree_add_12_51_groupi_n_5375 ,csa_tree_add_12_51_groupi_n_5374);
  and csa_tree_add_12_51_groupi_g16394(csa_tree_add_12_51_groupi_n_5373 ,csa_tree_add_12_51_groupi_n_5211 ,csa_tree_add_12_51_groupi_n_5317);
  or csa_tree_add_12_51_groupi_g16395(csa_tree_add_12_51_groupi_n_5372 ,csa_tree_add_12_51_groupi_n_5251 ,csa_tree_add_12_51_groupi_n_5265);
  nor csa_tree_add_12_51_groupi_g16396(csa_tree_add_12_51_groupi_n_5371 ,csa_tree_add_12_51_groupi_n_5252 ,csa_tree_add_12_51_groupi_n_5264);
  or csa_tree_add_12_51_groupi_g16397(csa_tree_add_12_51_groupi_n_5370 ,csa_tree_add_12_51_groupi_n_6 ,csa_tree_add_12_51_groupi_n_5149);
  and csa_tree_add_12_51_groupi_g16398(csa_tree_add_12_51_groupi_n_5369 ,csa_tree_add_12_51_groupi_n_5245 ,csa_tree_add_12_51_groupi_n_5147);
  or csa_tree_add_12_51_groupi_g16399(csa_tree_add_12_51_groupi_n_5368 ,csa_tree_add_12_51_groupi_n_5258 ,csa_tree_add_12_51_groupi_n_5099);
  and csa_tree_add_12_51_groupi_g16400(csa_tree_add_12_51_groupi_n_5367 ,csa_tree_add_12_51_groupi_n_5110 ,csa_tree_add_12_51_groupi_n_5299);
  nor csa_tree_add_12_51_groupi_g16401(csa_tree_add_12_51_groupi_n_5366 ,csa_tree_add_12_51_groupi_n_5259 ,csa_tree_add_12_51_groupi_n_5100);
  or csa_tree_add_12_51_groupi_g16402(csa_tree_add_12_51_groupi_n_5365 ,csa_tree_add_12_51_groupi_n_5052 ,csa_tree_add_12_51_groupi_n_5266);
  nor csa_tree_add_12_51_groupi_g16403(csa_tree_add_12_51_groupi_n_5364 ,csa_tree_add_12_51_groupi_n_5220 ,csa_tree_add_12_51_groupi_n_5310);
  and csa_tree_add_12_51_groupi_g16404(csa_tree_add_12_51_groupi_n_5363 ,csa_tree_add_12_51_groupi_n_5052 ,csa_tree_add_12_51_groupi_n_5266);
  nor csa_tree_add_12_51_groupi_g16405(csa_tree_add_12_51_groupi_n_5362 ,csa_tree_add_12_51_groupi_n_5250 ,csa_tree_add_12_51_groupi_n_5249);
  and csa_tree_add_12_51_groupi_g16406(csa_tree_add_12_51_groupi_n_5361 ,csa_tree_add_12_51_groupi_n_5250 ,csa_tree_add_12_51_groupi_n_5249);
  or csa_tree_add_12_51_groupi_g16407(csa_tree_add_12_51_groupi_n_5360 ,csa_tree_add_12_51_groupi_n_5245 ,csa_tree_add_12_51_groupi_n_5147);
  or csa_tree_add_12_51_groupi_g16408(csa_tree_add_12_51_groupi_n_5359 ,csa_tree_add_12_51_groupi_n_5053 ,csa_tree_add_12_51_groupi_n_5267);
  and csa_tree_add_12_51_groupi_g16409(csa_tree_add_12_51_groupi_n_5358 ,csa_tree_add_12_51_groupi_n_5187 ,csa_tree_add_12_51_groupi_n_5305);
  and csa_tree_add_12_51_groupi_g16410(csa_tree_add_12_51_groupi_n_5357 ,csa_tree_add_12_51_groupi_n_5053 ,csa_tree_add_12_51_groupi_n_5267);
  and csa_tree_add_12_51_groupi_g16411(csa_tree_add_12_51_groupi_n_5356 ,csa_tree_add_12_51_groupi_n_5055 ,csa_tree_add_12_51_groupi_n_5263);
  or csa_tree_add_12_51_groupi_g16412(csa_tree_add_12_51_groupi_n_5355 ,csa_tree_add_12_51_groupi_n_5106 ,csa_tree_add_12_51_groupi_n_5301);
  or csa_tree_add_12_51_groupi_g16413(csa_tree_add_12_51_groupi_n_5354 ,csa_tree_add_12_51_groupi_n_5055 ,csa_tree_add_12_51_groupi_n_5263);
  and csa_tree_add_12_51_groupi_g16414(csa_tree_add_12_51_groupi_n_5353 ,csa_tree_add_12_51_groupi_n_5054 ,csa_tree_add_12_51_groupi_n_5268);
  or csa_tree_add_12_51_groupi_g16415(csa_tree_add_12_51_groupi_n_5352 ,csa_tree_add_12_51_groupi_n_5054 ,csa_tree_add_12_51_groupi_n_5268);
  or csa_tree_add_12_51_groupi_g16416(csa_tree_add_12_51_groupi_n_5385 ,csa_tree_add_12_51_groupi_n_5210 ,csa_tree_add_12_51_groupi_n_5303);
  or csa_tree_add_12_51_groupi_g16417(csa_tree_add_12_51_groupi_n_5383 ,csa_tree_add_12_51_groupi_n_5209 ,csa_tree_add_12_51_groupi_n_5313);
  and csa_tree_add_12_51_groupi_g16418(csa_tree_add_12_51_groupi_n_5382 ,csa_tree_add_12_51_groupi_n_2456 ,csa_tree_add_12_51_groupi_n_5307);
  and csa_tree_add_12_51_groupi_g16419(csa_tree_add_12_51_groupi_n_5381 ,csa_tree_add_12_51_groupi_n_5197 ,csa_tree_add_12_51_groupi_n_5308);
  or csa_tree_add_12_51_groupi_g16420(csa_tree_add_12_51_groupi_n_5380 ,csa_tree_add_12_51_groupi_n_5199 ,csa_tree_add_12_51_groupi_n_5309);
  or csa_tree_add_12_51_groupi_g16421(csa_tree_add_12_51_groupi_n_5379 ,csa_tree_add_12_51_groupi_n_5203 ,csa_tree_add_12_51_groupi_n_5312);
  or csa_tree_add_12_51_groupi_g16422(csa_tree_add_12_51_groupi_n_5378 ,csa_tree_add_12_51_groupi_n_5206 ,csa_tree_add_12_51_groupi_n_5314);
  or csa_tree_add_12_51_groupi_g16423(csa_tree_add_12_51_groupi_n_5376 ,csa_tree_add_12_51_groupi_n_5191 ,csa_tree_add_12_51_groupi_n_5315);
  or csa_tree_add_12_51_groupi_g16424(csa_tree_add_12_51_groupi_n_5374 ,csa_tree_add_12_51_groupi_n_5192 ,csa_tree_add_12_51_groupi_n_5304);
  not csa_tree_add_12_51_groupi_g16425(csa_tree_add_12_51_groupi_n_5348 ,csa_tree_add_12_51_groupi_n_5349);
  or csa_tree_add_12_51_groupi_g16426(csa_tree_add_12_51_groupi_n_5345 ,csa_tree_add_12_51_groupi_n_3714 ,csa_tree_add_12_51_groupi_n_5235);
  and csa_tree_add_12_51_groupi_g16427(csa_tree_add_12_51_groupi_n_5344 ,csa_tree_add_12_51_groupi_n_5316 ,csa_tree_add_12_51_groupi_n_5295);
  or csa_tree_add_12_51_groupi_g16428(csa_tree_add_12_51_groupi_n_5343 ,csa_tree_add_12_51_groupi_n_5253 ,csa_tree_add_12_51_groupi_n_5256);
  nor csa_tree_add_12_51_groupi_g16429(csa_tree_add_12_51_groupi_n_5342 ,csa_tree_add_12_51_groupi_n_5254 ,csa_tree_add_12_51_groupi_n_5257);
  or csa_tree_add_12_51_groupi_g16430(csa_tree_add_12_51_groupi_n_5341 ,csa_tree_add_12_51_groupi_n_3112 ,csa_tree_add_12_51_groupi_n_5298);
  or csa_tree_add_12_51_groupi_g16431(csa_tree_add_12_51_groupi_n_5340 ,csa_tree_add_12_51_groupi_n_3730 ,csa_tree_add_12_51_groupi_n_5233);
  or csa_tree_add_12_51_groupi_g16432(csa_tree_add_12_51_groupi_n_5339 ,csa_tree_add_12_51_groupi_n_3726 ,csa_tree_add_12_51_groupi_n_5244);
  or csa_tree_add_12_51_groupi_g16433(csa_tree_add_12_51_groupi_n_5338 ,csa_tree_add_12_51_groupi_n_3649 ,csa_tree_add_12_51_groupi_n_5242);
  or csa_tree_add_12_51_groupi_g16434(csa_tree_add_12_51_groupi_n_5337 ,csa_tree_add_12_51_groupi_n_3671 ,csa_tree_add_12_51_groupi_n_5243);
  or csa_tree_add_12_51_groupi_g16435(csa_tree_add_12_51_groupi_n_5336 ,csa_tree_add_12_51_groupi_n_2985 ,csa_tree_add_12_51_groupi_n_5241);
  or csa_tree_add_12_51_groupi_g16436(csa_tree_add_12_51_groupi_n_5335 ,csa_tree_add_12_51_groupi_n_3586 ,csa_tree_add_12_51_groupi_n_5236);
  or csa_tree_add_12_51_groupi_g16437(csa_tree_add_12_51_groupi_n_5334 ,csa_tree_add_12_51_groupi_n_3737 ,csa_tree_add_12_51_groupi_n_5240);
  or csa_tree_add_12_51_groupi_g16438(csa_tree_add_12_51_groupi_n_5333 ,csa_tree_add_12_51_groupi_n_3697 ,csa_tree_add_12_51_groupi_n_5239);
  or csa_tree_add_12_51_groupi_g16439(csa_tree_add_12_51_groupi_n_5332 ,csa_tree_add_12_51_groupi_n_3720 ,csa_tree_add_12_51_groupi_n_5238);
  or csa_tree_add_12_51_groupi_g16440(csa_tree_add_12_51_groupi_n_5331 ,csa_tree_add_12_51_groupi_n_3647 ,csa_tree_add_12_51_groupi_n_5237);
  or csa_tree_add_12_51_groupi_g16441(csa_tree_add_12_51_groupi_n_5330 ,csa_tree_add_12_51_groupi_n_3685 ,csa_tree_add_12_51_groupi_n_5234);
  nor csa_tree_add_12_51_groupi_g16442(csa_tree_add_12_51_groupi_n_5329 ,csa_tree_add_12_51_groupi_n_5262 ,csa_tree_add_12_51_groupi_n_5150);
  or csa_tree_add_12_51_groupi_g16443(csa_tree_add_12_51_groupi_n_5328 ,csa_tree_add_12_51_groupi_n_3155 ,csa_tree_add_12_51_groupi_n_5293);
  or csa_tree_add_12_51_groupi_g16444(csa_tree_add_12_51_groupi_n_5327 ,csa_tree_add_12_51_groupi_n_3046 ,csa_tree_add_12_51_groupi_n_5297);
  xnor csa_tree_add_12_51_groupi_g16445(csa_tree_add_12_51_groupi_n_5326 ,csa_tree_add_12_51_groupi_n_4848 ,csa_tree_add_12_51_groupi_n_5217);
  xnor csa_tree_add_12_51_groupi_g16446(csa_tree_add_12_51_groupi_n_5325 ,csa_tree_add_12_51_groupi_n_5220 ,csa_tree_add_12_51_groupi_n_5215);
  xnor csa_tree_add_12_51_groupi_g16447(csa_tree_add_12_51_groupi_n_5324 ,csa_tree_add_12_51_groupi_n_4884 ,csa_tree_add_12_51_groupi_n_5183);
  xnor csa_tree_add_12_51_groupi_g16448(csa_tree_add_12_51_groupi_n_5323 ,csa_tree_add_12_51_groupi_n_4935 ,csa_tree_add_12_51_groupi_n_5189);
  xnor csa_tree_add_12_51_groupi_g16449(csa_tree_add_12_51_groupi_n_5322 ,csa_tree_add_12_51_groupi_n_4936 ,csa_tree_add_12_51_groupi_n_5184);
  xnor csa_tree_add_12_51_groupi_g16450(csa_tree_add_12_51_groupi_n_5321 ,csa_tree_add_12_51_groupi_n_5090 ,csa_tree_add_12_51_groupi_n_5178);
  xnor csa_tree_add_12_51_groupi_g16451(csa_tree_add_12_51_groupi_n_5320 ,csa_tree_add_12_51_groupi_n_4933 ,csa_tree_add_12_51_groupi_n_5188);
  xnor csa_tree_add_12_51_groupi_g16452(csa_tree_add_12_51_groupi_n_5319 ,csa_tree_add_12_51_groupi_n_4885 ,csa_tree_add_12_51_groupi_n_5179);
  xnor csa_tree_add_12_51_groupi_g16453(csa_tree_add_12_51_groupi_n_5351 ,csa_tree_add_12_51_groupi_n_4944 ,csa_tree_add_12_51_groupi_n_5157);
  xnor csa_tree_add_12_51_groupi_g16454(csa_tree_add_12_51_groupi_n_5350 ,csa_tree_add_12_51_groupi_n_4929 ,csa_tree_add_12_51_groupi_n_5156);
  or csa_tree_add_12_51_groupi_g16455(csa_tree_add_12_51_groupi_n_5349 ,csa_tree_add_12_51_groupi_n_5204 ,csa_tree_add_12_51_groupi_n_5294);
  xnor csa_tree_add_12_51_groupi_g16456(csa_tree_add_12_51_groupi_n_5347 ,csa_tree_add_12_51_groupi_n_4490 ,csa_tree_add_12_51_groupi_n_5155);
  xnor csa_tree_add_12_51_groupi_g16457(csa_tree_add_12_51_groupi_n_5346 ,csa_tree_add_12_51_groupi_n_5222 ,csa_tree_add_12_51_groupi_n_2557);
  and csa_tree_add_12_51_groupi_g16458(csa_tree_add_12_51_groupi_n_5315 ,csa_tree_add_12_51_groupi_n_5111 ,csa_tree_add_12_51_groupi_n_5194);
  nor csa_tree_add_12_51_groupi_g16459(csa_tree_add_12_51_groupi_n_5314 ,csa_tree_add_12_51_groupi_n_5205 ,csa_tree_add_12_51_groupi_n_5223);
  and csa_tree_add_12_51_groupi_g16460(csa_tree_add_12_51_groupi_n_5313 ,csa_tree_add_12_51_groupi_n_5107 ,csa_tree_add_12_51_groupi_n_5207);
  and csa_tree_add_12_51_groupi_g16461(csa_tree_add_12_51_groupi_n_5312 ,csa_tree_add_12_51_groupi_n_5109 ,csa_tree_add_12_51_groupi_n_5202);
  nor csa_tree_add_12_51_groupi_g16462(csa_tree_add_12_51_groupi_n_5311 ,csa_tree_add_12_51_groupi_n_5215 ,csa_tree_add_12_51_groupi_n_4679);
  and csa_tree_add_12_51_groupi_g16463(csa_tree_add_12_51_groupi_n_5310 ,csa_tree_add_12_51_groupi_n_5215 ,csa_tree_add_12_51_groupi_n_4679);
  and csa_tree_add_12_51_groupi_g16464(csa_tree_add_12_51_groupi_n_5309 ,csa_tree_add_12_51_groupi_n_5112 ,csa_tree_add_12_51_groupi_n_5198);
  or csa_tree_add_12_51_groupi_g16465(csa_tree_add_12_51_groupi_n_5308 ,csa_tree_add_12_51_groupi_n_5196 ,csa_tree_add_12_51_groupi_n_5190);
  or csa_tree_add_12_51_groupi_g16466(csa_tree_add_12_51_groupi_n_5307 ,csa_tree_add_12_51_groupi_n_2458 ,csa_tree_add_12_51_groupi_n_5222);
  and csa_tree_add_12_51_groupi_g16467(csa_tree_add_12_51_groupi_n_5306 ,csa_tree_add_12_51_groupi_n_5090 ,csa_tree_add_12_51_groupi_n_5178);
  or csa_tree_add_12_51_groupi_g16468(csa_tree_add_12_51_groupi_n_5305 ,csa_tree_add_12_51_groupi_n_5090 ,csa_tree_add_12_51_groupi_n_5178);
  and csa_tree_add_12_51_groupi_g16469(csa_tree_add_12_51_groupi_n_5304 ,csa_tree_add_12_51_groupi_n_5108 ,csa_tree_add_12_51_groupi_n_5193);
  and csa_tree_add_12_51_groupi_g16470(csa_tree_add_12_51_groupi_n_5303 ,csa_tree_add_12_51_groupi_n_5208 ,csa_tree_add_12_51_groupi_n_5188);
  or csa_tree_add_12_51_groupi_g16471(csa_tree_add_12_51_groupi_n_5302 ,csa_tree_add_12_51_groupi_n_4883 ,csa_tree_add_12_51_groupi_n_5182);
  nor csa_tree_add_12_51_groupi_g16472(csa_tree_add_12_51_groupi_n_5301 ,csa_tree_add_12_51_groupi_n_4884 ,csa_tree_add_12_51_groupi_n_5183);
  and csa_tree_add_12_51_groupi_g16473(csa_tree_add_12_51_groupi_n_5300 ,csa_tree_add_12_51_groupi_n_4885 ,csa_tree_add_12_51_groupi_n_5179);
  or csa_tree_add_12_51_groupi_g16474(csa_tree_add_12_51_groupi_n_5299 ,csa_tree_add_12_51_groupi_n_4885 ,csa_tree_add_12_51_groupi_n_5179);
  nor csa_tree_add_12_51_groupi_g16475(csa_tree_add_12_51_groupi_n_5298 ,csa_tree_add_12_51_groupi_n_1605 ,csa_tree_add_12_51_groupi_n_824);
  nor csa_tree_add_12_51_groupi_g16476(csa_tree_add_12_51_groupi_n_5297 ,csa_tree_add_12_51_groupi_n_1593 ,csa_tree_add_12_51_groupi_n_827);
  and csa_tree_add_12_51_groupi_g16477(csa_tree_add_12_51_groupi_n_5296 ,csa_tree_add_12_51_groupi_n_4936 ,csa_tree_add_12_51_groupi_n_5184);
  or csa_tree_add_12_51_groupi_g16478(csa_tree_add_12_51_groupi_n_5295 ,csa_tree_add_12_51_groupi_n_4936 ,csa_tree_add_12_51_groupi_n_5184);
  and csa_tree_add_12_51_groupi_g16479(csa_tree_add_12_51_groupi_n_5294 ,csa_tree_add_12_51_groupi_n_5201 ,csa_tree_add_12_51_groupi_n_5221);
  nor csa_tree_add_12_51_groupi_g16480(csa_tree_add_12_51_groupi_n_5293 ,csa_tree_add_12_51_groupi_n_1584 ,csa_tree_add_12_51_groupi_n_181);
  nor csa_tree_add_12_51_groupi_g16481(csa_tree_add_12_51_groupi_n_5292 ,csa_tree_add_12_51_groupi_n_4848 ,csa_tree_add_12_51_groupi_n_5218);
  and csa_tree_add_12_51_groupi_g16482(csa_tree_add_12_51_groupi_n_5291 ,csa_tree_add_12_51_groupi_n_4848 ,csa_tree_add_12_51_groupi_n_5218);
  nor csa_tree_add_12_51_groupi_g16483(csa_tree_add_12_51_groupi_n_5290 ,csa_tree_add_12_51_groupi_n_3858 ,csa_tree_add_12_51_groupi_n_5164);
  nor csa_tree_add_12_51_groupi_g16484(csa_tree_add_12_51_groupi_n_5289 ,csa_tree_add_12_51_groupi_n_4064 ,csa_tree_add_12_51_groupi_n_5173);
  nor csa_tree_add_12_51_groupi_g16485(csa_tree_add_12_51_groupi_n_5288 ,csa_tree_add_12_51_groupi_n_4066 ,csa_tree_add_12_51_groupi_n_5174);
  nor csa_tree_add_12_51_groupi_g16486(csa_tree_add_12_51_groupi_n_5287 ,csa_tree_add_12_51_groupi_n_4114 ,csa_tree_add_12_51_groupi_n_5172);
  nor csa_tree_add_12_51_groupi_g16487(csa_tree_add_12_51_groupi_n_5286 ,csa_tree_add_12_51_groupi_n_3901 ,csa_tree_add_12_51_groupi_n_5168);
  nor csa_tree_add_12_51_groupi_g16488(csa_tree_add_12_51_groupi_n_5285 ,csa_tree_add_12_51_groupi_n_3900 ,csa_tree_add_12_51_groupi_n_5167);
  nor csa_tree_add_12_51_groupi_g16489(csa_tree_add_12_51_groupi_n_5284 ,csa_tree_add_12_51_groupi_n_3457 ,csa_tree_add_12_51_groupi_n_5161);
  nor csa_tree_add_12_51_groupi_g16490(csa_tree_add_12_51_groupi_n_5283 ,csa_tree_add_12_51_groupi_n_3861 ,csa_tree_add_12_51_groupi_n_5163);
  nor csa_tree_add_12_51_groupi_g16491(csa_tree_add_12_51_groupi_n_5282 ,csa_tree_add_12_51_groupi_n_3849 ,csa_tree_add_12_51_groupi_n_5165);
  nor csa_tree_add_12_51_groupi_g16492(csa_tree_add_12_51_groupi_n_5281 ,csa_tree_add_12_51_groupi_n_3905 ,csa_tree_add_12_51_groupi_n_5170);
  nor csa_tree_add_12_51_groupi_g16493(csa_tree_add_12_51_groupi_n_5280 ,csa_tree_add_12_51_groupi_n_3919 ,csa_tree_add_12_51_groupi_n_5171);
  nor csa_tree_add_12_51_groupi_g16494(csa_tree_add_12_51_groupi_n_5279 ,csa_tree_add_12_51_groupi_n_3864 ,csa_tree_add_12_51_groupi_n_5166);
  nor csa_tree_add_12_51_groupi_g16495(csa_tree_add_12_51_groupi_n_5278 ,csa_tree_add_12_51_groupi_n_3456 ,csa_tree_add_12_51_groupi_n_5162);
  nor csa_tree_add_12_51_groupi_g16496(csa_tree_add_12_51_groupi_n_5277 ,csa_tree_add_12_51_groupi_n_3442 ,csa_tree_add_12_51_groupi_n_5160);
  nor csa_tree_add_12_51_groupi_g16497(csa_tree_add_12_51_groupi_n_5276 ,csa_tree_add_12_51_groupi_n_3926 ,csa_tree_add_12_51_groupi_n_5169);
  and csa_tree_add_12_51_groupi_g16498(csa_tree_add_12_51_groupi_n_5318 ,csa_tree_add_12_51_groupi_n_4963 ,csa_tree_add_12_51_groupi_n_5159);
  or csa_tree_add_12_51_groupi_g16499(csa_tree_add_12_51_groupi_n_5317 ,csa_tree_add_12_51_groupi_n_5139 ,csa_tree_add_12_51_groupi_n_5200);
  or csa_tree_add_12_51_groupi_g16500(csa_tree_add_12_51_groupi_n_5316 ,csa_tree_add_12_51_groupi_n_5030 ,csa_tree_add_12_51_groupi_n_5195);
  not csa_tree_add_12_51_groupi_g16501(csa_tree_add_12_51_groupi_n_5275 ,csa_tree_add_12_51_groupi_n_5274);
  not csa_tree_add_12_51_groupi_g16502(csa_tree_add_12_51_groupi_n_5270 ,csa_tree_add_12_51_groupi_n_5269);
  not csa_tree_add_12_51_groupi_g16503(csa_tree_add_12_51_groupi_n_5265 ,csa_tree_add_12_51_groupi_n_5264);
  not csa_tree_add_12_51_groupi_g16504(csa_tree_add_12_51_groupi_n_5262 ,csa_tree_add_12_51_groupi_n_6);
  not csa_tree_add_12_51_groupi_g16505(csa_tree_add_12_51_groupi_n_5259 ,csa_tree_add_12_51_groupi_n_5258);
  not csa_tree_add_12_51_groupi_g16506(csa_tree_add_12_51_groupi_n_5257 ,csa_tree_add_12_51_groupi_n_5256);
  not csa_tree_add_12_51_groupi_g16507(csa_tree_add_12_51_groupi_n_5253 ,csa_tree_add_12_51_groupi_n_5254);
  not csa_tree_add_12_51_groupi_g16508(csa_tree_add_12_51_groupi_n_5251 ,csa_tree_add_12_51_groupi_n_5252);
  not csa_tree_add_12_51_groupi_g16509(csa_tree_add_12_51_groupi_n_5249 ,csa_tree_add_12_51_groupi_n_5248);
  not csa_tree_add_12_51_groupi_g16510(csa_tree_add_12_51_groupi_n_5247 ,csa_tree_add_12_51_groupi_n_5246);
  nor csa_tree_add_12_51_groupi_g16511(csa_tree_add_12_51_groupi_n_5244 ,csa_tree_add_12_51_groupi_n_1656 ,csa_tree_add_12_51_groupi_n_824);
  nor csa_tree_add_12_51_groupi_g16512(csa_tree_add_12_51_groupi_n_5243 ,csa_tree_add_12_51_groupi_n_1623 ,csa_tree_add_12_51_groupi_n_825);
  nor csa_tree_add_12_51_groupi_g16513(csa_tree_add_12_51_groupi_n_5242 ,csa_tree_add_12_51_groupi_n_1629 ,csa_tree_add_12_51_groupi_n_828);
  nor csa_tree_add_12_51_groupi_g16514(csa_tree_add_12_51_groupi_n_5241 ,csa_tree_add_12_51_groupi_n_1641 ,csa_tree_add_12_51_groupi_n_900);
  nor csa_tree_add_12_51_groupi_g16515(csa_tree_add_12_51_groupi_n_5240 ,csa_tree_add_12_51_groupi_n_1665 ,csa_tree_add_12_51_groupi_n_899);
  nor csa_tree_add_12_51_groupi_g16516(csa_tree_add_12_51_groupi_n_5239 ,csa_tree_add_12_51_groupi_n_1647 ,csa_tree_add_12_51_groupi_n_825);
  nor csa_tree_add_12_51_groupi_g16517(csa_tree_add_12_51_groupi_n_5238 ,csa_tree_add_12_51_groupi_n_1611 ,csa_tree_add_12_51_groupi_n_899);
  nor csa_tree_add_12_51_groupi_g16518(csa_tree_add_12_51_groupi_n_5237 ,csa_tree_add_12_51_groupi_n_1635 ,csa_tree_add_12_51_groupi_n_828);
  nor csa_tree_add_12_51_groupi_g16519(csa_tree_add_12_51_groupi_n_5236 ,csa_tree_add_12_51_groupi_n_1587 ,csa_tree_add_12_51_groupi_n_827);
  nor csa_tree_add_12_51_groupi_g16520(csa_tree_add_12_51_groupi_n_5235 ,csa_tree_add_12_51_groupi_n_1680 ,csa_tree_add_12_51_groupi_n_2004);
  nor csa_tree_add_12_51_groupi_g16521(csa_tree_add_12_51_groupi_n_5234 ,csa_tree_add_12_51_groupi_n_1599 ,csa_tree_add_12_51_groupi_n_900);
  nor csa_tree_add_12_51_groupi_g16522(csa_tree_add_12_51_groupi_n_5233 ,csa_tree_add_12_51_groupi_n_1617 ,csa_tree_add_12_51_groupi_n_181);
  xnor csa_tree_add_12_51_groupi_g16523(out3[3] ,csa_tree_add_12_51_groupi_n_5153 ,csa_tree_add_12_51_groupi_n_5068);
  xnor csa_tree_add_12_51_groupi_g16524(csa_tree_add_12_51_groupi_n_5231 ,csa_tree_add_12_51_groupi_n_5088 ,csa_tree_add_12_51_groupi_n_4924);
  xnor csa_tree_add_12_51_groupi_g16525(csa_tree_add_12_51_groupi_n_5230 ,csa_tree_add_12_51_groupi_n_5095 ,csa_tree_add_12_51_groupi_n_5089);
  xnor csa_tree_add_12_51_groupi_g16526(csa_tree_add_12_51_groupi_n_5229 ,csa_tree_add_12_51_groupi_n_5097 ,csa_tree_add_12_51_groupi_n_4916);
  xnor csa_tree_add_12_51_groupi_g16527(csa_tree_add_12_51_groupi_n_5228 ,csa_tree_add_12_51_groupi_n_5103 ,csa_tree_add_12_51_groupi_n_5096);
  xnor csa_tree_add_12_51_groupi_g16528(csa_tree_add_12_51_groupi_n_5227 ,csa_tree_add_12_51_groupi_n_4882 ,csa_tree_add_12_51_groupi_n_5102);
  xnor csa_tree_add_12_51_groupi_g16529(csa_tree_add_12_51_groupi_n_5226 ,csa_tree_add_12_51_groupi_n_4886 ,csa_tree_add_12_51_groupi_n_5101);
  xnor csa_tree_add_12_51_groupi_g16530(csa_tree_add_12_51_groupi_n_5225 ,csa_tree_add_12_51_groupi_n_5104 ,csa_tree_add_12_51_groupi_n_5087);
  xnor csa_tree_add_12_51_groupi_g16531(csa_tree_add_12_51_groupi_n_5224 ,csa_tree_add_12_51_groupi_n_5092 ,csa_tree_add_12_51_groupi_n_5026);
  xnor csa_tree_add_12_51_groupi_g16533(csa_tree_add_12_51_groupi_n_5274 ,csa_tree_add_12_51_groupi_n_5125 ,in3[11]);
  xnor csa_tree_add_12_51_groupi_g16534(csa_tree_add_12_51_groupi_n_5273 ,csa_tree_add_12_51_groupi_n_4939 ,csa_tree_add_12_51_groupi_n_5073);
  xnor csa_tree_add_12_51_groupi_g16535(csa_tree_add_12_51_groupi_n_5272 ,csa_tree_add_12_51_groupi_n_5124 ,in2[2]);
  xnor csa_tree_add_12_51_groupi_g16536(csa_tree_add_12_51_groupi_n_5271 ,csa_tree_add_12_51_groupi_n_5061 ,csa_tree_add_12_51_groupi_n_5074);
  xnor csa_tree_add_12_51_groupi_g16537(csa_tree_add_12_51_groupi_n_5269 ,csa_tree_add_12_51_groupi_n_5116 ,in2[8]);
  xnor csa_tree_add_12_51_groupi_g16538(csa_tree_add_12_51_groupi_n_5268 ,csa_tree_add_12_51_groupi_n_4940 ,csa_tree_add_12_51_groupi_n_5071);
  xnor csa_tree_add_12_51_groupi_g16539(csa_tree_add_12_51_groupi_n_5267 ,csa_tree_add_12_51_groupi_n_4941 ,csa_tree_add_12_51_groupi_n_5075);
  xnor csa_tree_add_12_51_groupi_g16540(csa_tree_add_12_51_groupi_n_5266 ,csa_tree_add_12_51_groupi_n_4943 ,csa_tree_add_12_51_groupi_n_5069);
  xnor csa_tree_add_12_51_groupi_g16541(csa_tree_add_12_51_groupi_n_5264 ,csa_tree_add_12_51_groupi_n_5122 ,in3[5]);
  xnor csa_tree_add_12_51_groupi_g16542(csa_tree_add_12_51_groupi_n_5263 ,csa_tree_add_12_51_groupi_n_5066 ,csa_tree_add_12_51_groupi_n_5070);
  xnor csa_tree_add_12_51_groupi_g16544(csa_tree_add_12_51_groupi_n_5261 ,csa_tree_add_12_51_groupi_n_4634 ,csa_tree_add_12_51_groupi_n_5067);
  xnor csa_tree_add_12_51_groupi_g16545(csa_tree_add_12_51_groupi_n_5260 ,csa_tree_add_12_51_groupi_n_5127 ,in3[2]);
  xnor csa_tree_add_12_51_groupi_g16546(csa_tree_add_12_51_groupi_n_5258 ,csa_tree_add_12_51_groupi_n_112 ,csa_tree_add_12_51_groupi_n_5126);
  xnor csa_tree_add_12_51_groupi_g16547(csa_tree_add_12_51_groupi_n_5256 ,csa_tree_add_12_51_groupi_n_5151 ,csa_tree_add_12_51_groupi_n_4991);
  xnor csa_tree_add_12_51_groupi_g16548(csa_tree_add_12_51_groupi_n_5255 ,csa_tree_add_12_51_groupi_n_5114 ,in4[5]);
  xnor csa_tree_add_12_51_groupi_g16549(csa_tree_add_12_51_groupi_n_5254 ,csa_tree_add_12_51_groupi_n_5118 ,in4[11]);
  xnor csa_tree_add_12_51_groupi_g16550(csa_tree_add_12_51_groupi_n_5252 ,csa_tree_add_12_51_groupi_n_5123 ,in2[5]);
  xnor csa_tree_add_12_51_groupi_g16551(csa_tree_add_12_51_groupi_n_5250 ,csa_tree_add_12_51_groupi_n_1918 ,csa_tree_add_12_51_groupi_n_5119);
  xnor csa_tree_add_12_51_groupi_g16552(csa_tree_add_12_51_groupi_n_5248 ,csa_tree_add_12_51_groupi_n_5121 ,in2[14]);
  xnor csa_tree_add_12_51_groupi_g16553(csa_tree_add_12_51_groupi_n_5246 ,csa_tree_add_12_51_groupi_n_5115 ,in3[8]);
  xnor csa_tree_add_12_51_groupi_g16554(csa_tree_add_12_51_groupi_n_5245 ,csa_tree_add_12_51_groupi_n_5113 ,in4[2]);
  not csa_tree_add_12_51_groupi_g16555(csa_tree_add_12_51_groupi_n_5218 ,csa_tree_add_12_51_groupi_n_5217);
  not csa_tree_add_12_51_groupi_g16556(csa_tree_add_12_51_groupi_n_5213 ,csa_tree_add_12_51_groupi_n_5214);
  and csa_tree_add_12_51_groupi_g16557(csa_tree_add_12_51_groupi_n_5212 ,csa_tree_add_12_51_groupi_n_5103 ,csa_tree_add_12_51_groupi_n_5096);
  or csa_tree_add_12_51_groupi_g16558(csa_tree_add_12_51_groupi_n_5211 ,csa_tree_add_12_51_groupi_n_5103 ,csa_tree_add_12_51_groupi_n_5096);
  and csa_tree_add_12_51_groupi_g16559(csa_tree_add_12_51_groupi_n_5210 ,csa_tree_add_12_51_groupi_n_5098 ,csa_tree_add_12_51_groupi_n_4933);
  and csa_tree_add_12_51_groupi_g16560(csa_tree_add_12_51_groupi_n_5209 ,csa_tree_add_12_51_groupi_n_5088 ,csa_tree_add_12_51_groupi_n_4924);
  or csa_tree_add_12_51_groupi_g16561(csa_tree_add_12_51_groupi_n_5208 ,csa_tree_add_12_51_groupi_n_5098 ,csa_tree_add_12_51_groupi_n_4933);
  or csa_tree_add_12_51_groupi_g16562(csa_tree_add_12_51_groupi_n_5207 ,csa_tree_add_12_51_groupi_n_5088 ,csa_tree_add_12_51_groupi_n_4924);
  and csa_tree_add_12_51_groupi_g16563(csa_tree_add_12_51_groupi_n_5206 ,csa_tree_add_12_51_groupi_n_5095 ,csa_tree_add_12_51_groupi_n_5089);
  nor csa_tree_add_12_51_groupi_g16564(csa_tree_add_12_51_groupi_n_5205 ,csa_tree_add_12_51_groupi_n_5095 ,csa_tree_add_12_51_groupi_n_5089);
  nor csa_tree_add_12_51_groupi_g16565(csa_tree_add_12_51_groupi_n_5204 ,csa_tree_add_12_51_groupi_n_5091 ,csa_tree_add_12_51_groupi_n_5026);
  and csa_tree_add_12_51_groupi_g16566(csa_tree_add_12_51_groupi_n_5203 ,csa_tree_add_12_51_groupi_n_5097 ,csa_tree_add_12_51_groupi_n_4916);
  or csa_tree_add_12_51_groupi_g16567(csa_tree_add_12_51_groupi_n_5202 ,csa_tree_add_12_51_groupi_n_5097 ,csa_tree_add_12_51_groupi_n_4916);
  or csa_tree_add_12_51_groupi_g16568(csa_tree_add_12_51_groupi_n_5201 ,csa_tree_add_12_51_groupi_n_5092 ,csa_tree_add_12_51_groupi_n_5025);
  and csa_tree_add_12_51_groupi_g16569(csa_tree_add_12_51_groupi_n_5200 ,csa_tree_add_12_51_groupi_n_4944 ,csa_tree_add_12_51_groupi_n_5140);
  and csa_tree_add_12_51_groupi_g16570(csa_tree_add_12_51_groupi_n_5199 ,csa_tree_add_12_51_groupi_n_5104 ,csa_tree_add_12_51_groupi_n_5087);
  or csa_tree_add_12_51_groupi_g16571(csa_tree_add_12_51_groupi_n_5198 ,csa_tree_add_12_51_groupi_n_5104 ,csa_tree_add_12_51_groupi_n_5087);
  or csa_tree_add_12_51_groupi_g16572(csa_tree_add_12_51_groupi_n_5197 ,csa_tree_add_12_51_groupi_n_5085 ,csa_tree_add_12_51_groupi_n_4934);
  nor csa_tree_add_12_51_groupi_g16573(csa_tree_add_12_51_groupi_n_5196 ,csa_tree_add_12_51_groupi_n_5086 ,csa_tree_add_12_51_groupi_n_4935);
  and csa_tree_add_12_51_groupi_g16574(csa_tree_add_12_51_groupi_n_5195 ,csa_tree_add_12_51_groupi_n_5153 ,csa_tree_add_12_51_groupi_n_5031);
  or csa_tree_add_12_51_groupi_g16575(csa_tree_add_12_51_groupi_n_5194 ,csa_tree_add_12_51_groupi_n_4886 ,csa_tree_add_12_51_groupi_n_5101);
  or csa_tree_add_12_51_groupi_g16576(csa_tree_add_12_51_groupi_n_5193 ,csa_tree_add_12_51_groupi_n_4882 ,csa_tree_add_12_51_groupi_n_5102);
  and csa_tree_add_12_51_groupi_g16577(csa_tree_add_12_51_groupi_n_5192 ,csa_tree_add_12_51_groupi_n_4882 ,csa_tree_add_12_51_groupi_n_5102);
  and csa_tree_add_12_51_groupi_g16578(csa_tree_add_12_51_groupi_n_5191 ,csa_tree_add_12_51_groupi_n_4886 ,csa_tree_add_12_51_groupi_n_5101);
  and csa_tree_add_12_51_groupi_g16579(csa_tree_add_12_51_groupi_n_5223 ,csa_tree_add_12_51_groupi_n_5049 ,csa_tree_add_12_51_groupi_n_5137);
  and csa_tree_add_12_51_groupi_g16580(csa_tree_add_12_51_groupi_n_5222 ,csa_tree_add_12_51_groupi_n_2427 ,csa_tree_add_12_51_groupi_n_5142);
  or csa_tree_add_12_51_groupi_g16581(csa_tree_add_12_51_groupi_n_5221 ,csa_tree_add_12_51_groupi_n_5014 ,csa_tree_add_12_51_groupi_n_5146);
  and csa_tree_add_12_51_groupi_g16582(csa_tree_add_12_51_groupi_n_5220 ,csa_tree_add_12_51_groupi_n_5043 ,csa_tree_add_12_51_groupi_n_5143);
  or csa_tree_add_12_51_groupi_g16583(csa_tree_add_12_51_groupi_n_5219 ,csa_tree_add_12_51_groupi_n_5006 ,csa_tree_add_12_51_groupi_n_5135);
  or csa_tree_add_12_51_groupi_g16584(csa_tree_add_12_51_groupi_n_5217 ,csa_tree_add_12_51_groupi_n_4810 ,csa_tree_add_12_51_groupi_n_5136);
  or csa_tree_add_12_51_groupi_g16585(csa_tree_add_12_51_groupi_n_5216 ,csa_tree_add_12_51_groupi_n_5045 ,csa_tree_add_12_51_groupi_n_5144);
  and csa_tree_add_12_51_groupi_g16586(csa_tree_add_12_51_groupi_n_5215 ,csa_tree_add_12_51_groupi_n_5029 ,csa_tree_add_12_51_groupi_n_5138);
  or csa_tree_add_12_51_groupi_g16587(csa_tree_add_12_51_groupi_n_5214 ,csa_tree_add_12_51_groupi_n_5039 ,csa_tree_add_12_51_groupi_n_5145);
  not csa_tree_add_12_51_groupi_g16588(csa_tree_add_12_51_groupi_n_5190 ,csa_tree_add_12_51_groupi_n_5189);
  not csa_tree_add_12_51_groupi_g16589(csa_tree_add_12_51_groupi_n_5185 ,csa_tree_add_12_51_groupi_n_5186);
  not csa_tree_add_12_51_groupi_g16590(csa_tree_add_12_51_groupi_n_5182 ,csa_tree_add_12_51_groupi_n_5183);
  not csa_tree_add_12_51_groupi_g16591(csa_tree_add_12_51_groupi_n_5180 ,csa_tree_add_12_51_groupi_n_5181);
  not csa_tree_add_12_51_groupi_g16592(csa_tree_add_12_51_groupi_n_5176 ,csa_tree_add_12_51_groupi_n_5177);
  or csa_tree_add_12_51_groupi_g16593(csa_tree_add_12_51_groupi_n_5174 ,csa_tree_add_12_51_groupi_n_3280 ,csa_tree_add_12_51_groupi_n_5080);
  or csa_tree_add_12_51_groupi_g16594(csa_tree_add_12_51_groupi_n_5173 ,csa_tree_add_12_51_groupi_n_3258 ,csa_tree_add_12_51_groupi_n_5077);
  or csa_tree_add_12_51_groupi_g16595(csa_tree_add_12_51_groupi_n_5172 ,csa_tree_add_12_51_groupi_n_3263 ,csa_tree_add_12_51_groupi_n_5076);
  or csa_tree_add_12_51_groupi_g16596(csa_tree_add_12_51_groupi_n_5171 ,csa_tree_add_12_51_groupi_n_3659 ,csa_tree_add_12_51_groupi_n_5133);
  or csa_tree_add_12_51_groupi_g16597(csa_tree_add_12_51_groupi_n_5170 ,csa_tree_add_12_51_groupi_n_3704 ,csa_tree_add_12_51_groupi_n_5134);
  or csa_tree_add_12_51_groupi_g16598(csa_tree_add_12_51_groupi_n_5169 ,csa_tree_add_12_51_groupi_n_3691 ,csa_tree_add_12_51_groupi_n_5141);
  or csa_tree_add_12_51_groupi_g16599(csa_tree_add_12_51_groupi_n_5168 ,csa_tree_add_12_51_groupi_n_3602 ,csa_tree_add_12_51_groupi_n_5084);
  or csa_tree_add_12_51_groupi_g16600(csa_tree_add_12_51_groupi_n_5167 ,csa_tree_add_12_51_groupi_n_3628 ,csa_tree_add_12_51_groupi_n_5083);
  or csa_tree_add_12_51_groupi_g16601(csa_tree_add_12_51_groupi_n_5166 ,csa_tree_add_12_51_groupi_n_3763 ,csa_tree_add_12_51_groupi_n_5082);
  or csa_tree_add_12_51_groupi_g16602(csa_tree_add_12_51_groupi_n_5165 ,csa_tree_add_12_51_groupi_n_3674 ,csa_tree_add_12_51_groupi_n_5081);
  or csa_tree_add_12_51_groupi_g16603(csa_tree_add_12_51_groupi_n_5164 ,csa_tree_add_12_51_groupi_n_3663 ,csa_tree_add_12_51_groupi_n_5079);
  or csa_tree_add_12_51_groupi_g16604(csa_tree_add_12_51_groupi_n_5163 ,csa_tree_add_12_51_groupi_n_3728 ,csa_tree_add_12_51_groupi_n_5078);
  or csa_tree_add_12_51_groupi_g16605(csa_tree_add_12_51_groupi_n_5162 ,csa_tree_add_12_51_groupi_n_3037 ,csa_tree_add_12_51_groupi_n_5130);
  or csa_tree_add_12_51_groupi_g16606(csa_tree_add_12_51_groupi_n_5161 ,csa_tree_add_12_51_groupi_n_3018 ,csa_tree_add_12_51_groupi_n_5131);
  or csa_tree_add_12_51_groupi_g16607(csa_tree_add_12_51_groupi_n_5160 ,csa_tree_add_12_51_groupi_n_3113 ,csa_tree_add_12_51_groupi_n_5129);
  or csa_tree_add_12_51_groupi_g16608(csa_tree_add_12_51_groupi_n_5159 ,csa_tree_add_12_51_groupi_n_4962 ,csa_tree_add_12_51_groupi_n_5152);
  xnor csa_tree_add_12_51_groupi_g16609(out3[2] ,csa_tree_add_12_51_groupi_n_4893 ,csa_tree_add_12_51_groupi_n_4990);
  xnor csa_tree_add_12_51_groupi_g16610(csa_tree_add_12_51_groupi_n_5157 ,csa_tree_add_12_51_groupi_n_4930 ,csa_tree_add_12_51_groupi_n_5058);
  xnor csa_tree_add_12_51_groupi_g16611(csa_tree_add_12_51_groupi_n_5156 ,csa_tree_add_12_51_groupi_n_4937 ,csa_tree_add_12_51_groupi_n_5064);
  xnor csa_tree_add_12_51_groupi_g16612(csa_tree_add_12_51_groupi_n_5155 ,csa_tree_add_12_51_groupi_n_4917 ,csa_tree_add_12_51_groupi_n_5059);
  xnor csa_tree_add_12_51_groupi_g16613(csa_tree_add_12_51_groupi_n_5189 ,csa_tree_add_12_51_groupi_n_4890 ,csa_tree_add_12_51_groupi_n_4994);
  xnor csa_tree_add_12_51_groupi_g16614(csa_tree_add_12_51_groupi_n_5188 ,csa_tree_add_12_51_groupi_n_4880 ,csa_tree_add_12_51_groupi_n_4993);
  or csa_tree_add_12_51_groupi_g16615(csa_tree_add_12_51_groupi_n_5187 ,csa_tree_add_12_51_groupi_n_5003 ,csa_tree_add_12_51_groupi_n_5128);
  xnor csa_tree_add_12_51_groupi_g16616(csa_tree_add_12_51_groupi_n_5186 ,csa_tree_add_12_51_groupi_n_5065 ,csa_tree_add_12_51_groupi_n_4823);
  xnor csa_tree_add_12_51_groupi_g16617(csa_tree_add_12_51_groupi_n_5184 ,csa_tree_add_12_51_groupi_n_4892 ,csa_tree_add_12_51_groupi_n_4997);
  xnor csa_tree_add_12_51_groupi_g16618(csa_tree_add_12_51_groupi_n_5183 ,csa_tree_add_12_51_groupi_n_4766 ,csa_tree_add_12_51_groupi_n_4992);
  or csa_tree_add_12_51_groupi_g16619(csa_tree_add_12_51_groupi_n_5181 ,csa_tree_add_12_51_groupi_n_5008 ,csa_tree_add_12_51_groupi_n_5132);
  xnor csa_tree_add_12_51_groupi_g16620(csa_tree_add_12_51_groupi_n_5179 ,csa_tree_add_12_51_groupi_n_4765 ,csa_tree_add_12_51_groupi_n_4996);
  xnor csa_tree_add_12_51_groupi_g16621(csa_tree_add_12_51_groupi_n_5178 ,csa_tree_add_12_51_groupi_n_4881 ,csa_tree_add_12_51_groupi_n_4995);
  xnor csa_tree_add_12_51_groupi_g16622(csa_tree_add_12_51_groupi_n_5177 ,csa_tree_add_12_51_groupi_n_4493 ,csa_tree_add_12_51_groupi_n_4998);
  xnor csa_tree_add_12_51_groupi_g16623(csa_tree_add_12_51_groupi_n_5175 ,csa_tree_add_12_51_groupi_n_5063 ,csa_tree_add_12_51_groupi_n_2566);
  not csa_tree_add_12_51_groupi_g16624(csa_tree_add_12_51_groupi_n_5152 ,csa_tree_add_12_51_groupi_n_5151);
  not csa_tree_add_12_51_groupi_g16625(csa_tree_add_12_51_groupi_n_5149 ,csa_tree_add_12_51_groupi_n_5150);
  and csa_tree_add_12_51_groupi_g16626(csa_tree_add_12_51_groupi_n_5146 ,csa_tree_add_12_51_groupi_n_4940 ,csa_tree_add_12_51_groupi_n_5013);
  and csa_tree_add_12_51_groupi_g16627(csa_tree_add_12_51_groupi_n_5145 ,csa_tree_add_12_51_groupi_n_5046 ,csa_tree_add_12_51_groupi_n_5064);
  and csa_tree_add_12_51_groupi_g16628(csa_tree_add_12_51_groupi_n_5144 ,csa_tree_add_12_51_groupi_n_4939 ,csa_tree_add_12_51_groupi_n_5038);
  or csa_tree_add_12_51_groupi_g16629(csa_tree_add_12_51_groupi_n_5143 ,csa_tree_add_12_51_groupi_n_5041 ,csa_tree_add_12_51_groupi_n_5060);
  or csa_tree_add_12_51_groupi_g16630(csa_tree_add_12_51_groupi_n_5142 ,csa_tree_add_12_51_groupi_n_2433 ,csa_tree_add_12_51_groupi_n_5063);
  nor csa_tree_add_12_51_groupi_g16631(csa_tree_add_12_51_groupi_n_5141 ,csa_tree_add_12_51_groupi_n_90 ,csa_tree_add_12_51_groupi_n_800);
  or csa_tree_add_12_51_groupi_g16632(csa_tree_add_12_51_groupi_n_5140 ,csa_tree_add_12_51_groupi_n_4930 ,csa_tree_add_12_51_groupi_n_5058);
  and csa_tree_add_12_51_groupi_g16633(csa_tree_add_12_51_groupi_n_5139 ,csa_tree_add_12_51_groupi_n_4930 ,csa_tree_add_12_51_groupi_n_5058);
  or csa_tree_add_12_51_groupi_g16634(csa_tree_add_12_51_groupi_n_5138 ,csa_tree_add_12_51_groupi_n_4942 ,csa_tree_add_12_51_groupi_n_5034);
  or csa_tree_add_12_51_groupi_g16635(csa_tree_add_12_51_groupi_n_5137 ,csa_tree_add_12_51_groupi_n_5048 ,csa_tree_add_12_51_groupi_n_5062);
  and csa_tree_add_12_51_groupi_g16636(csa_tree_add_12_51_groupi_n_5136 ,csa_tree_add_12_51_groupi_n_4811 ,csa_tree_add_12_51_groupi_n_5065);
  and csa_tree_add_12_51_groupi_g16637(csa_tree_add_12_51_groupi_n_5135 ,csa_tree_add_12_51_groupi_n_4943 ,csa_tree_add_12_51_groupi_n_5005);
  nor csa_tree_add_12_51_groupi_g16638(csa_tree_add_12_51_groupi_n_5134 ,csa_tree_add_12_51_groupi_n_88 ,csa_tree_add_12_51_groupi_n_803);
  nor csa_tree_add_12_51_groupi_g16639(csa_tree_add_12_51_groupi_n_5133 ,csa_tree_add_12_51_groupi_n_70 ,csa_tree_add_12_51_groupi_n_171);
  and csa_tree_add_12_51_groupi_g16640(csa_tree_add_12_51_groupi_n_5132 ,csa_tree_add_12_51_groupi_n_4941 ,csa_tree_add_12_51_groupi_n_5007);
  nor csa_tree_add_12_51_groupi_g16641(csa_tree_add_12_51_groupi_n_5131 ,csa_tree_add_12_51_groupi_n_80 ,csa_tree_add_12_51_groupi_n_800);
  nor csa_tree_add_12_51_groupi_g16642(csa_tree_add_12_51_groupi_n_5130 ,csa_tree_add_12_51_groupi_n_68 ,csa_tree_add_12_51_groupi_n_801);
  nor csa_tree_add_12_51_groupi_g16643(csa_tree_add_12_51_groupi_n_5129 ,csa_tree_add_12_51_groupi_n_74 ,csa_tree_add_12_51_groupi_n_804);
  and csa_tree_add_12_51_groupi_g16644(csa_tree_add_12_51_groupi_n_5128 ,csa_tree_add_12_51_groupi_n_5066 ,csa_tree_add_12_51_groupi_n_5002);
  nor csa_tree_add_12_51_groupi_g16645(csa_tree_add_12_51_groupi_n_5127 ,csa_tree_add_12_51_groupi_n_3449 ,csa_tree_add_12_51_groupi_n_5010);
  nor csa_tree_add_12_51_groupi_g16646(csa_tree_add_12_51_groupi_n_5126 ,csa_tree_add_12_51_groupi_n_4094 ,csa_tree_add_12_51_groupi_n_5015);
  nor csa_tree_add_12_51_groupi_g16647(csa_tree_add_12_51_groupi_n_5125 ,csa_tree_add_12_51_groupi_n_4067 ,csa_tree_add_12_51_groupi_n_5040);
  nor csa_tree_add_12_51_groupi_g16648(csa_tree_add_12_51_groupi_n_5124 ,csa_tree_add_12_51_groupi_n_3447 ,csa_tree_add_12_51_groupi_n_5012);
  nor csa_tree_add_12_51_groupi_g16649(csa_tree_add_12_51_groupi_n_5123 ,csa_tree_add_12_51_groupi_n_3881 ,csa_tree_add_12_51_groupi_n_5018);
  nor csa_tree_add_12_51_groupi_g16650(csa_tree_add_12_51_groupi_n_5122 ,csa_tree_add_12_51_groupi_n_3925 ,csa_tree_add_12_51_groupi_n_5044);
  nor csa_tree_add_12_51_groupi_g16651(csa_tree_add_12_51_groupi_n_5121 ,csa_tree_add_12_51_groupi_n_3921 ,csa_tree_add_12_51_groupi_n_5047);
  nor csa_tree_add_12_51_groupi_g16652(csa_tree_add_12_51_groupi_n_5120 ,csa_tree_add_12_51_groupi_n_3863 ,csa_tree_add_12_51_groupi_n_5017);
  nor csa_tree_add_12_51_groupi_g16653(csa_tree_add_12_51_groupi_n_5119 ,csa_tree_add_12_51_groupi_n_3886 ,csa_tree_add_12_51_groupi_n_5051);
  nor csa_tree_add_12_51_groupi_g16654(csa_tree_add_12_51_groupi_n_5118 ,csa_tree_add_12_51_groupi_n_4103 ,csa_tree_add_12_51_groupi_n_5042);
  nor csa_tree_add_12_51_groupi_g16655(csa_tree_add_12_51_groupi_n_5117 ,csa_tree_add_12_51_groupi_n_3896 ,csa_tree_add_12_51_groupi_n_5019);
  nor csa_tree_add_12_51_groupi_g16656(csa_tree_add_12_51_groupi_n_5116 ,csa_tree_add_12_51_groupi_n_3894 ,csa_tree_add_12_51_groupi_n_5000);
  nor csa_tree_add_12_51_groupi_g16657(csa_tree_add_12_51_groupi_n_5115 ,csa_tree_add_12_51_groupi_n_3854 ,csa_tree_add_12_51_groupi_n_5016);
  nor csa_tree_add_12_51_groupi_g16658(csa_tree_add_12_51_groupi_n_5114 ,csa_tree_add_12_51_groupi_n_4054 ,csa_tree_add_12_51_groupi_n_5037);
  nor csa_tree_add_12_51_groupi_g16659(csa_tree_add_12_51_groupi_n_5113 ,csa_tree_add_12_51_groupi_n_3455 ,csa_tree_add_12_51_groupi_n_5011);
  and csa_tree_add_12_51_groupi_g16660(csa_tree_add_12_51_groupi_n_5154 ,csa_tree_add_12_51_groupi_n_4976 ,csa_tree_add_12_51_groupi_n_5009);
  or csa_tree_add_12_51_groupi_g16661(csa_tree_add_12_51_groupi_n_5153 ,csa_tree_add_12_51_groupi_n_4961 ,csa_tree_add_12_51_groupi_n_5035);
  or csa_tree_add_12_51_groupi_g16662(csa_tree_add_12_51_groupi_n_5151 ,csa_tree_add_12_51_groupi_n_4970 ,csa_tree_add_12_51_groupi_n_5050);
  or csa_tree_add_12_51_groupi_g16663(csa_tree_add_12_51_groupi_n_5150 ,csa_tree_add_12_51_groupi_n_4982 ,csa_tree_add_12_51_groupi_n_5001);
  or csa_tree_add_12_51_groupi_g16664(csa_tree_add_12_51_groupi_n_5148 ,csa_tree_add_12_51_groupi_n_4912 ,csa_tree_add_12_51_groupi_n_5036);
  or csa_tree_add_12_51_groupi_g16665(csa_tree_add_12_51_groupi_n_5147 ,csa_tree_add_12_51_groupi_n_4981 ,csa_tree_add_12_51_groupi_n_5004);
  not csa_tree_add_12_51_groupi_g16666(csa_tree_add_12_51_groupi_n_5106 ,csa_tree_add_12_51_groupi_n_5105);
  not csa_tree_add_12_51_groupi_g16667(csa_tree_add_12_51_groupi_n_5099 ,csa_tree_add_12_51_groupi_n_5100);
  not csa_tree_add_12_51_groupi_g16668(csa_tree_add_12_51_groupi_n_5093 ,csa_tree_add_12_51_groupi_n_5094);
  not csa_tree_add_12_51_groupi_g16669(csa_tree_add_12_51_groupi_n_5091 ,csa_tree_add_12_51_groupi_n_5092);
  not csa_tree_add_12_51_groupi_g16670(csa_tree_add_12_51_groupi_n_5086 ,csa_tree_add_12_51_groupi_n_5085);
  nor csa_tree_add_12_51_groupi_g16671(csa_tree_add_12_51_groupi_n_5084 ,csa_tree_add_12_51_groupi_n_94 ,csa_tree_add_12_51_groupi_n_846);
  nor csa_tree_add_12_51_groupi_g16672(csa_tree_add_12_51_groupi_n_5083 ,csa_tree_add_12_51_groupi_n_84 ,csa_tree_add_12_51_groupi_n_845);
  nor csa_tree_add_12_51_groupi_g16673(csa_tree_add_12_51_groupi_n_5082 ,csa_tree_add_12_51_groupi_n_86 ,csa_tree_add_12_51_groupi_n_801);
  nor csa_tree_add_12_51_groupi_g16674(csa_tree_add_12_51_groupi_n_5081 ,csa_tree_add_12_51_groupi_n_82 ,csa_tree_add_12_51_groupi_n_845);
  nor csa_tree_add_12_51_groupi_g16675(csa_tree_add_12_51_groupi_n_5080 ,csa_tree_add_12_51_groupi_n_76 ,csa_tree_add_12_51_groupi_n_804);
  nor csa_tree_add_12_51_groupi_g16676(csa_tree_add_12_51_groupi_n_5079 ,csa_tree_add_12_51_groupi_n_72 ,csa_tree_add_12_51_groupi_n_803);
  nor csa_tree_add_12_51_groupi_g16677(csa_tree_add_12_51_groupi_n_5078 ,csa_tree_add_12_51_groupi_n_78 ,csa_tree_add_12_51_groupi_n_1989);
  nor csa_tree_add_12_51_groupi_g16678(csa_tree_add_12_51_groupi_n_5077 ,csa_tree_add_12_51_groupi_n_92 ,csa_tree_add_12_51_groupi_n_846);
  nor csa_tree_add_12_51_groupi_g16679(csa_tree_add_12_51_groupi_n_5076 ,csa_tree_add_12_51_groupi_n_66 ,csa_tree_add_12_51_groupi_n_171);
  xnor csa_tree_add_12_51_groupi_g16680(csa_tree_add_12_51_groupi_n_5075 ,csa_tree_add_12_51_groupi_n_4846 ,csa_tree_add_12_51_groupi_n_4928);
  xnor csa_tree_add_12_51_groupi_g16681(csa_tree_add_12_51_groupi_n_5074 ,csa_tree_add_12_51_groupi_n_4923 ,csa_tree_add_12_51_groupi_n_4932);
  xnor csa_tree_add_12_51_groupi_g16682(csa_tree_add_12_51_groupi_n_5073 ,csa_tree_add_12_51_groupi_n_4915 ,csa_tree_add_12_51_groupi_n_4914);
  xnor csa_tree_add_12_51_groupi_g16683(csa_tree_add_12_51_groupi_n_5072 ,csa_tree_add_12_51_groupi_n_4666 ,csa_tree_add_12_51_groupi_n_4989);
  xnor csa_tree_add_12_51_groupi_g16684(csa_tree_add_12_51_groupi_n_5071 ,csa_tree_add_12_51_groupi_n_4755 ,csa_tree_add_12_51_groupi_n_4927);
  xnor csa_tree_add_12_51_groupi_g16685(csa_tree_add_12_51_groupi_n_5070 ,csa_tree_add_12_51_groupi_n_4850 ,csa_tree_add_12_51_groupi_n_4926);
  xnor csa_tree_add_12_51_groupi_g16686(csa_tree_add_12_51_groupi_n_5069 ,csa_tree_add_12_51_groupi_n_4842 ,csa_tree_add_12_51_groupi_n_4925);
  xnor csa_tree_add_12_51_groupi_g16687(csa_tree_add_12_51_groupi_n_5068 ,csa_tree_add_12_51_groupi_n_4938 ,csa_tree_add_12_51_groupi_n_4849);
  xnor csa_tree_add_12_51_groupi_g16688(csa_tree_add_12_51_groupi_n_5067 ,csa_tree_add_12_51_groupi_n_4919 ,csa_tree_add_12_51_groupi_n_4942);
  xnor csa_tree_add_12_51_groupi_g16689(csa_tree_add_12_51_groupi_n_5112 ,csa_tree_add_12_51_groupi_n_4954 ,in3[14]);
  xnor csa_tree_add_12_51_groupi_g16690(csa_tree_add_12_51_groupi_n_5111 ,csa_tree_add_12_51_groupi_n_4758 ,csa_tree_add_12_51_groupi_n_4898);
  xnor csa_tree_add_12_51_groupi_g16691(csa_tree_add_12_51_groupi_n_5110 ,csa_tree_add_12_51_groupi_n_4773 ,csa_tree_add_12_51_groupi_n_4901);
  xnor csa_tree_add_12_51_groupi_g16692(csa_tree_add_12_51_groupi_n_5109 ,csa_tree_add_12_51_groupi_n_4957 ,in2[2]);
  xnor csa_tree_add_12_51_groupi_g16693(csa_tree_add_12_51_groupi_n_5108 ,csa_tree_add_12_51_groupi_n_4771 ,csa_tree_add_12_51_groupi_n_4899);
  xnor csa_tree_add_12_51_groupi_g16694(csa_tree_add_12_51_groupi_n_5107 ,csa_tree_add_12_51_groupi_n_4945 ,in3[11]);
  xnor csa_tree_add_12_51_groupi_g16695(csa_tree_add_12_51_groupi_n_5105 ,csa_tree_add_12_51_groupi_n_4770 ,csa_tree_add_12_51_groupi_n_4896);
  xnor csa_tree_add_12_51_groupi_g16696(csa_tree_add_12_51_groupi_n_5104 ,csa_tree_add_12_51_groupi_n_4952 ,in4[14]);
  xnor csa_tree_add_12_51_groupi_g16697(csa_tree_add_12_51_groupi_n_5103 ,csa_tree_add_12_51_groupi_n_4951 ,in2[8]);
  xnor csa_tree_add_12_51_groupi_g16698(csa_tree_add_12_51_groupi_n_5102 ,csa_tree_add_12_51_groupi_n_4891 ,csa_tree_add_12_51_groupi_n_4900);
  xnor csa_tree_add_12_51_groupi_g16699(csa_tree_add_12_51_groupi_n_5101 ,csa_tree_add_12_51_groupi_n_4855 ,csa_tree_add_12_51_groupi_n_4897);
  xnor csa_tree_add_12_51_groupi_g16700(csa_tree_add_12_51_groupi_n_5100 ,csa_tree_add_12_51_groupi_n_4772 ,csa_tree_add_12_51_groupi_n_4895);
  xnor csa_tree_add_12_51_groupi_g16701(csa_tree_add_12_51_groupi_n_5098 ,csa_tree_add_12_51_groupi_n_4950 ,in3[5]);
  xnor csa_tree_add_12_51_groupi_g16702(csa_tree_add_12_51_groupi_n_5097 ,csa_tree_add_12_51_groupi_n_4956 ,in4[2]);
  xnor csa_tree_add_12_51_groupi_g16703(csa_tree_add_12_51_groupi_n_5096 ,csa_tree_add_12_51_groupi_n_4955 ,in3[8]);
  xnor csa_tree_add_12_51_groupi_g16704(csa_tree_add_12_51_groupi_n_5095 ,csa_tree_add_12_51_groupi_n_4946 ,in4[5]);
  xnor csa_tree_add_12_51_groupi_g16705(csa_tree_add_12_51_groupi_n_5094 ,csa_tree_add_12_51_groupi_n_4498 ,csa_tree_add_12_51_groupi_n_4894);
  xnor csa_tree_add_12_51_groupi_g16706(csa_tree_add_12_51_groupi_n_5092 ,csa_tree_add_12_51_groupi_n_4949 ,in4[11]);
  xnor csa_tree_add_12_51_groupi_g16707(csa_tree_add_12_51_groupi_n_5090 ,csa_tree_add_12_51_groupi_n_4958 ,in3[2]);
  xnor csa_tree_add_12_51_groupi_g16708(csa_tree_add_12_51_groupi_n_5089 ,csa_tree_add_12_51_groupi_n_4947 ,in2[5]);
  xnor csa_tree_add_12_51_groupi_g16709(csa_tree_add_12_51_groupi_n_5088 ,csa_tree_add_12_51_groupi_n_4959 ,in2[11]);
  xnor csa_tree_add_12_51_groupi_g16710(csa_tree_add_12_51_groupi_n_5087 ,csa_tree_add_12_51_groupi_n_4953 ,in2[14]);
  xnor csa_tree_add_12_51_groupi_g16711(csa_tree_add_12_51_groupi_n_5085 ,csa_tree_add_12_51_groupi_n_4948 ,csa_tree_add_12_51_groupi_n_1939);
  not csa_tree_add_12_51_groupi_g16712(csa_tree_add_12_51_groupi_n_5062 ,csa_tree_add_12_51_groupi_n_5061);
  not csa_tree_add_12_51_groupi_g16713(csa_tree_add_12_51_groupi_n_5060 ,csa_tree_add_12_51_groupi_n_5059);
  not csa_tree_add_12_51_groupi_g16714(csa_tree_add_12_51_groupi_n_5057 ,csa_tree_add_12_51_groupi_n_5056);
  or csa_tree_add_12_51_groupi_g16715(csa_tree_add_12_51_groupi_n_5051 ,csa_tree_add_12_51_groupi_n_3690 ,csa_tree_add_12_51_groupi_n_4902);
  and csa_tree_add_12_51_groupi_g16716(csa_tree_add_12_51_groupi_n_5050 ,csa_tree_add_12_51_groupi_n_4719 ,csa_tree_add_12_51_groupi_n_4972);
  or csa_tree_add_12_51_groupi_g16717(csa_tree_add_12_51_groupi_n_5049 ,csa_tree_add_12_51_groupi_n_4922 ,csa_tree_add_12_51_groupi_n_4931);
  nor csa_tree_add_12_51_groupi_g16718(csa_tree_add_12_51_groupi_n_5048 ,csa_tree_add_12_51_groupi_n_4923 ,csa_tree_add_12_51_groupi_n_4932);
  or csa_tree_add_12_51_groupi_g16719(csa_tree_add_12_51_groupi_n_5047 ,csa_tree_add_12_51_groupi_n_3681 ,csa_tree_add_12_51_groupi_n_4986);
  or csa_tree_add_12_51_groupi_g16720(csa_tree_add_12_51_groupi_n_5046 ,csa_tree_add_12_51_groupi_n_4929 ,csa_tree_add_12_51_groupi_n_4937);
  and csa_tree_add_12_51_groupi_g16721(csa_tree_add_12_51_groupi_n_5045 ,csa_tree_add_12_51_groupi_n_4915 ,csa_tree_add_12_51_groupi_n_4914);
  or csa_tree_add_12_51_groupi_g16722(csa_tree_add_12_51_groupi_n_5044 ,csa_tree_add_12_51_groupi_n_3603 ,csa_tree_add_12_51_groupi_n_4985);
  or csa_tree_add_12_51_groupi_g16723(csa_tree_add_12_51_groupi_n_5043 ,csa_tree_add_12_51_groupi_n_9 ,csa_tree_add_12_51_groupi_n_4489);
  or csa_tree_add_12_51_groupi_g16724(csa_tree_add_12_51_groupi_n_5042 ,csa_tree_add_12_51_groupi_n_3256 ,csa_tree_add_12_51_groupi_n_4905);
  nor csa_tree_add_12_51_groupi_g16725(csa_tree_add_12_51_groupi_n_5041 ,csa_tree_add_12_51_groupi_n_4917 ,csa_tree_add_12_51_groupi_n_4490);
  or csa_tree_add_12_51_groupi_g16726(csa_tree_add_12_51_groupi_n_5040 ,csa_tree_add_12_51_groupi_n_3288 ,csa_tree_add_12_51_groupi_n_4909);
  and csa_tree_add_12_51_groupi_g16727(csa_tree_add_12_51_groupi_n_5039 ,csa_tree_add_12_51_groupi_n_4929 ,csa_tree_add_12_51_groupi_n_4937);
  or csa_tree_add_12_51_groupi_g16728(csa_tree_add_12_51_groupi_n_5038 ,csa_tree_add_12_51_groupi_n_4915 ,csa_tree_add_12_51_groupi_n_4914);
  or csa_tree_add_12_51_groupi_g16729(csa_tree_add_12_51_groupi_n_5037 ,csa_tree_add_12_51_groupi_n_3296 ,csa_tree_add_12_51_groupi_n_4907);
  and csa_tree_add_12_51_groupi_g16730(csa_tree_add_12_51_groupi_n_5036 ,csa_tree_add_12_51_groupi_n_4892 ,csa_tree_add_12_51_groupi_n_4911);
  and csa_tree_add_12_51_groupi_g16731(csa_tree_add_12_51_groupi_n_5035 ,csa_tree_add_12_51_groupi_n_4893 ,csa_tree_add_12_51_groupi_n_4960);
  nor csa_tree_add_12_51_groupi_g16732(csa_tree_add_12_51_groupi_n_5034 ,csa_tree_add_12_51_groupi_n_4918 ,csa_tree_add_12_51_groupi_n_4634);
  and csa_tree_add_12_51_groupi_g16733(csa_tree_add_12_51_groupi_n_5033 ,csa_tree_add_12_51_groupi_n_4666 ,csa_tree_add_12_51_groupi_n_4989);
  or csa_tree_add_12_51_groupi_g16734(csa_tree_add_12_51_groupi_n_5032 ,csa_tree_add_12_51_groupi_n_4666 ,csa_tree_add_12_51_groupi_n_4989);
  or csa_tree_add_12_51_groupi_g16735(csa_tree_add_12_51_groupi_n_5031 ,csa_tree_add_12_51_groupi_n_4938 ,csa_tree_add_12_51_groupi_n_4849);
  and csa_tree_add_12_51_groupi_g16736(csa_tree_add_12_51_groupi_n_5030 ,csa_tree_add_12_51_groupi_n_4938 ,csa_tree_add_12_51_groupi_n_4849);
  or csa_tree_add_12_51_groupi_g16737(csa_tree_add_12_51_groupi_n_5029 ,csa_tree_add_12_51_groupi_n_4919 ,csa_tree_add_12_51_groupi_n_4633);
  or csa_tree_add_12_51_groupi_g16738(csa_tree_add_12_51_groupi_n_5066 ,csa_tree_add_12_51_groupi_n_4865 ,csa_tree_add_12_51_groupi_n_4965);
  or csa_tree_add_12_51_groupi_g16739(csa_tree_add_12_51_groupi_n_5065 ,csa_tree_add_12_51_groupi_n_4627 ,csa_tree_add_12_51_groupi_n_4968);
  or csa_tree_add_12_51_groupi_g16740(csa_tree_add_12_51_groupi_n_5064 ,csa_tree_add_12_51_groupi_n_4856 ,csa_tree_add_12_51_groupi_n_4967);
  and csa_tree_add_12_51_groupi_g16741(csa_tree_add_12_51_groupi_n_5063 ,csa_tree_add_12_51_groupi_n_2422 ,csa_tree_add_12_51_groupi_n_4971);
  or csa_tree_add_12_51_groupi_g16742(csa_tree_add_12_51_groupi_n_5061 ,csa_tree_add_12_51_groupi_n_4871 ,csa_tree_add_12_51_groupi_n_4964);
  or csa_tree_add_12_51_groupi_g16743(csa_tree_add_12_51_groupi_n_5059 ,csa_tree_add_12_51_groupi_n_4859 ,csa_tree_add_12_51_groupi_n_4978);
  or csa_tree_add_12_51_groupi_g16744(csa_tree_add_12_51_groupi_n_5058 ,csa_tree_add_12_51_groupi_n_4864 ,csa_tree_add_12_51_groupi_n_4966);
  or csa_tree_add_12_51_groupi_g16745(csa_tree_add_12_51_groupi_n_5056 ,csa_tree_add_12_51_groupi_n_4572 ,csa_tree_add_12_51_groupi_n_4969);
  or csa_tree_add_12_51_groupi_g16746(csa_tree_add_12_51_groupi_n_5055 ,csa_tree_add_12_51_groupi_n_4866 ,csa_tree_add_12_51_groupi_n_4988);
  or csa_tree_add_12_51_groupi_g16747(csa_tree_add_12_51_groupi_n_5054 ,csa_tree_add_12_51_groupi_n_4863 ,csa_tree_add_12_51_groupi_n_4979);
  or csa_tree_add_12_51_groupi_g16748(csa_tree_add_12_51_groupi_n_5053 ,csa_tree_add_12_51_groupi_n_4861 ,csa_tree_add_12_51_groupi_n_4987);
  or csa_tree_add_12_51_groupi_g16749(csa_tree_add_12_51_groupi_n_5052 ,csa_tree_add_12_51_groupi_n_4867 ,csa_tree_add_12_51_groupi_n_4983);
  not csa_tree_add_12_51_groupi_g16750(csa_tree_add_12_51_groupi_n_5027 ,csa_tree_add_12_51_groupi_n_5028);
  not csa_tree_add_12_51_groupi_g16751(csa_tree_add_12_51_groupi_n_5025 ,csa_tree_add_12_51_groupi_n_5026);
  not csa_tree_add_12_51_groupi_g16752(csa_tree_add_12_51_groupi_n_5023 ,csa_tree_add_12_51_groupi_n_5024);
  not csa_tree_add_12_51_groupi_g16753(csa_tree_add_12_51_groupi_n_5021 ,csa_tree_add_12_51_groupi_n_5022);
  or csa_tree_add_12_51_groupi_g16754(csa_tree_add_12_51_groupi_n_5019 ,csa_tree_add_12_51_groupi_n_3695 ,csa_tree_add_12_51_groupi_n_4903);
  or csa_tree_add_12_51_groupi_g16755(csa_tree_add_12_51_groupi_n_5018 ,csa_tree_add_12_51_groupi_n_3600 ,csa_tree_add_12_51_groupi_n_4910);
  or csa_tree_add_12_51_groupi_g16756(csa_tree_add_12_51_groupi_n_5017 ,csa_tree_add_12_51_groupi_n_3592 ,csa_tree_add_12_51_groupi_n_4908);
  or csa_tree_add_12_51_groupi_g16757(csa_tree_add_12_51_groupi_n_5016 ,csa_tree_add_12_51_groupi_n_3601 ,csa_tree_add_12_51_groupi_n_4906);
  or csa_tree_add_12_51_groupi_g16758(csa_tree_add_12_51_groupi_n_5015 ,csa_tree_add_12_51_groupi_n_3073 ,csa_tree_add_12_51_groupi_n_4904);
  and csa_tree_add_12_51_groupi_g16759(csa_tree_add_12_51_groupi_n_5014 ,csa_tree_add_12_51_groupi_n_4755 ,csa_tree_add_12_51_groupi_n_4927);
  or csa_tree_add_12_51_groupi_g16760(csa_tree_add_12_51_groupi_n_5013 ,csa_tree_add_12_51_groupi_n_4755 ,csa_tree_add_12_51_groupi_n_4927);
  or csa_tree_add_12_51_groupi_g16761(csa_tree_add_12_51_groupi_n_5012 ,csa_tree_add_12_51_groupi_n_3082 ,csa_tree_add_12_51_groupi_n_4974);
  or csa_tree_add_12_51_groupi_g16762(csa_tree_add_12_51_groupi_n_5011 ,csa_tree_add_12_51_groupi_n_3052 ,csa_tree_add_12_51_groupi_n_4975);
  or csa_tree_add_12_51_groupi_g16763(csa_tree_add_12_51_groupi_n_5010 ,csa_tree_add_12_51_groupi_n_3094 ,csa_tree_add_12_51_groupi_n_4973);
  or csa_tree_add_12_51_groupi_g16764(csa_tree_add_12_51_groupi_n_5009 ,csa_tree_add_12_51_groupi_n_4728 ,csa_tree_add_12_51_groupi_n_4977);
  and csa_tree_add_12_51_groupi_g16765(csa_tree_add_12_51_groupi_n_5008 ,csa_tree_add_12_51_groupi_n_4846 ,csa_tree_add_12_51_groupi_n_4928);
  or csa_tree_add_12_51_groupi_g16766(csa_tree_add_12_51_groupi_n_5007 ,csa_tree_add_12_51_groupi_n_4846 ,csa_tree_add_12_51_groupi_n_4928);
  and csa_tree_add_12_51_groupi_g16767(csa_tree_add_12_51_groupi_n_5006 ,csa_tree_add_12_51_groupi_n_4842 ,csa_tree_add_12_51_groupi_n_4925);
  or csa_tree_add_12_51_groupi_g16768(csa_tree_add_12_51_groupi_n_5005 ,csa_tree_add_12_51_groupi_n_4842 ,csa_tree_add_12_51_groupi_n_4925);
  nor csa_tree_add_12_51_groupi_g16769(csa_tree_add_12_51_groupi_n_5004 ,csa_tree_add_12_51_groupi_n_4723 ,csa_tree_add_12_51_groupi_n_4980);
  and csa_tree_add_12_51_groupi_g16770(csa_tree_add_12_51_groupi_n_5003 ,csa_tree_add_12_51_groupi_n_4850 ,csa_tree_add_12_51_groupi_n_4926);
  or csa_tree_add_12_51_groupi_g16771(csa_tree_add_12_51_groupi_n_5002 ,csa_tree_add_12_51_groupi_n_4850 ,csa_tree_add_12_51_groupi_n_4926);
  and csa_tree_add_12_51_groupi_g16772(csa_tree_add_12_51_groupi_n_5001 ,csa_tree_add_12_51_groupi_n_4890 ,csa_tree_add_12_51_groupi_n_4984);
  or csa_tree_add_12_51_groupi_g16773(csa_tree_add_12_51_groupi_n_5000 ,csa_tree_add_12_51_groupi_n_3614 ,csa_tree_add_12_51_groupi_n_4913);
  xnor csa_tree_add_12_51_groupi_g16774(out3[1] ,csa_tree_add_12_51_groupi_n_4541 ,csa_tree_add_12_51_groupi_n_4822);
  xnor csa_tree_add_12_51_groupi_g16775(csa_tree_add_12_51_groupi_n_4998 ,csa_tree_add_12_51_groupi_n_4211 ,csa_tree_add_12_51_groupi_n_4854);
  xnor csa_tree_add_12_51_groupi_g16776(csa_tree_add_12_51_groupi_n_4997 ,csa_tree_add_12_51_groupi_n_4715 ,csa_tree_add_12_51_groupi_n_4847);
  xnor csa_tree_add_12_51_groupi_g16777(csa_tree_add_12_51_groupi_n_4996 ,csa_tree_add_12_51_groupi_n_4673 ,csa_tree_add_12_51_groupi_n_4888);
  xnor csa_tree_add_12_51_groupi_g16778(csa_tree_add_12_51_groupi_n_4995 ,csa_tree_add_12_51_groupi_n_4722 ,csa_tree_add_12_51_groupi_n_4851);
  xnor csa_tree_add_12_51_groupi_g16779(csa_tree_add_12_51_groupi_n_4994 ,csa_tree_add_12_51_groupi_n_4712 ,csa_tree_add_12_51_groupi_n_4852);
  xnor csa_tree_add_12_51_groupi_g16780(csa_tree_add_12_51_groupi_n_4993 ,csa_tree_add_12_51_groupi_n_4727 ,csa_tree_add_12_51_groupi_n_4844);
  xnor csa_tree_add_12_51_groupi_g16781(csa_tree_add_12_51_groupi_n_4992 ,csa_tree_add_12_51_groupi_n_4675 ,csa_tree_add_12_51_groupi_n_4889);
  xnor csa_tree_add_12_51_groupi_g16782(csa_tree_add_12_51_groupi_n_4991 ,csa_tree_add_12_51_groupi_n_4878 ,csa_tree_add_12_51_groupi_n_4583);
  xnor csa_tree_add_12_51_groupi_g16783(csa_tree_add_12_51_groupi_n_4990 ,csa_tree_add_12_51_groupi_n_4677 ,csa_tree_add_12_51_groupi_n_4845);
  xnor csa_tree_add_12_51_groupi_g16784(csa_tree_add_12_51_groupi_n_5028 ,csa_tree_add_12_51_groupi_n_4300 ,csa_tree_add_12_51_groupi_n_4821);
  xnor csa_tree_add_12_51_groupi_g16785(csa_tree_add_12_51_groupi_n_5026 ,csa_tree_add_12_51_groupi_n_4876 ,csa_tree_add_12_51_groupi_n_4818);
  xnor csa_tree_add_12_51_groupi_g16786(csa_tree_add_12_51_groupi_n_5024 ,csa_tree_add_12_51_groupi_n_4307 ,csa_tree_add_12_51_groupi_n_4820);
  xnor csa_tree_add_12_51_groupi_g16787(csa_tree_add_12_51_groupi_n_5022 ,csa_tree_add_12_51_groupi_n_4853 ,csa_tree_add_12_51_groupi_n_4648);
  xnor csa_tree_add_12_51_groupi_g16788(csa_tree_add_12_51_groupi_n_5020 ,csa_tree_add_12_51_groupi_n_4887 ,csa_tree_add_12_51_groupi_n_2563);
  nor csa_tree_add_12_51_groupi_g16789(csa_tree_add_12_51_groupi_n_4988 ,csa_tree_add_12_51_groupi_n_4769 ,csa_tree_add_12_51_groupi_n_4870);
  and csa_tree_add_12_51_groupi_g16790(csa_tree_add_12_51_groupi_n_4987 ,csa_tree_add_12_51_groupi_n_4771 ,csa_tree_add_12_51_groupi_n_4874);
  nor csa_tree_add_12_51_groupi_g16791(csa_tree_add_12_51_groupi_n_4986 ,csa_tree_add_12_51_groupi_n_51 ,csa_tree_add_12_51_groupi_n_1043);
  nor csa_tree_add_12_51_groupi_g16792(csa_tree_add_12_51_groupi_n_4985 ,csa_tree_add_12_51_groupi_n_60 ,csa_tree_add_12_51_groupi_n_812);
  or csa_tree_add_12_51_groupi_g16793(csa_tree_add_12_51_groupi_n_4984 ,csa_tree_add_12_51_groupi_n_4712 ,csa_tree_add_12_51_groupi_n_4852);
  and csa_tree_add_12_51_groupi_g16794(csa_tree_add_12_51_groupi_n_4983 ,csa_tree_add_12_51_groupi_n_4773 ,csa_tree_add_12_51_groupi_n_4869);
  and csa_tree_add_12_51_groupi_g16795(csa_tree_add_12_51_groupi_n_4982 ,csa_tree_add_12_51_groupi_n_4712 ,csa_tree_add_12_51_groupi_n_4852);
  and csa_tree_add_12_51_groupi_g16796(csa_tree_add_12_51_groupi_n_4981 ,csa_tree_add_12_51_groupi_n_4881 ,csa_tree_add_12_51_groupi_n_4851);
  nor csa_tree_add_12_51_groupi_g16797(csa_tree_add_12_51_groupi_n_4980 ,csa_tree_add_12_51_groupi_n_4881 ,csa_tree_add_12_51_groupi_n_4851);
  and csa_tree_add_12_51_groupi_g16798(csa_tree_add_12_51_groupi_n_4979 ,csa_tree_add_12_51_groupi_n_4770 ,csa_tree_add_12_51_groupi_n_4862);
  and csa_tree_add_12_51_groupi_g16799(csa_tree_add_12_51_groupi_n_4978 ,csa_tree_add_12_51_groupi_n_4772 ,csa_tree_add_12_51_groupi_n_4858);
  nor csa_tree_add_12_51_groupi_g16800(csa_tree_add_12_51_groupi_n_4977 ,csa_tree_add_12_51_groupi_n_4880 ,csa_tree_add_12_51_groupi_n_4844);
  or csa_tree_add_12_51_groupi_g16801(csa_tree_add_12_51_groupi_n_4976 ,csa_tree_add_12_51_groupi_n_4879 ,csa_tree_add_12_51_groupi_n_4843);
  nor csa_tree_add_12_51_groupi_g16802(csa_tree_add_12_51_groupi_n_4975 ,csa_tree_add_12_51_groupi_n_36 ,csa_tree_add_12_51_groupi_n_151);
  nor csa_tree_add_12_51_groupi_g16803(csa_tree_add_12_51_groupi_n_4974 ,csa_tree_add_12_51_groupi_n_42 ,csa_tree_add_12_51_groupi_n_1043);
  nor csa_tree_add_12_51_groupi_g16804(csa_tree_add_12_51_groupi_n_4973 ,csa_tree_add_12_51_groupi_n_27 ,csa_tree_add_12_51_groupi_n_1044);
  or csa_tree_add_12_51_groupi_g16805(csa_tree_add_12_51_groupi_n_4972 ,csa_tree_add_12_51_groupi_n_4491 ,csa_tree_add_12_51_groupi_n_4876);
  or csa_tree_add_12_51_groupi_g16806(csa_tree_add_12_51_groupi_n_4971 ,csa_tree_add_12_51_groupi_n_2419 ,csa_tree_add_12_51_groupi_n_4887);
  and csa_tree_add_12_51_groupi_g16807(csa_tree_add_12_51_groupi_n_4970 ,csa_tree_add_12_51_groupi_n_4491 ,csa_tree_add_12_51_groupi_n_4876);
  and csa_tree_add_12_51_groupi_g16808(csa_tree_add_12_51_groupi_n_4969 ,csa_tree_add_12_51_groupi_n_4571 ,csa_tree_add_12_51_groupi_n_4854);
  and csa_tree_add_12_51_groupi_g16809(csa_tree_add_12_51_groupi_n_4968 ,csa_tree_add_12_51_groupi_n_4629 ,csa_tree_add_12_51_groupi_n_4853);
  and csa_tree_add_12_51_groupi_g16810(csa_tree_add_12_51_groupi_n_4967 ,csa_tree_add_12_51_groupi_n_4889 ,csa_tree_add_12_51_groupi_n_4857);
  and csa_tree_add_12_51_groupi_g16811(csa_tree_add_12_51_groupi_n_4966 ,csa_tree_add_12_51_groupi_n_4891 ,csa_tree_add_12_51_groupi_n_4860);
  and csa_tree_add_12_51_groupi_g16812(csa_tree_add_12_51_groupi_n_4965 ,csa_tree_add_12_51_groupi_n_4855 ,csa_tree_add_12_51_groupi_n_4868);
  and csa_tree_add_12_51_groupi_g16813(csa_tree_add_12_51_groupi_n_4964 ,csa_tree_add_12_51_groupi_n_4888 ,csa_tree_add_12_51_groupi_n_4872);
  or csa_tree_add_12_51_groupi_g16814(csa_tree_add_12_51_groupi_n_4963 ,csa_tree_add_12_51_groupi_n_4877 ,csa_tree_add_12_51_groupi_n_4583);
  nor csa_tree_add_12_51_groupi_g16815(csa_tree_add_12_51_groupi_n_4962 ,csa_tree_add_12_51_groupi_n_4878 ,csa_tree_add_12_51_groupi_n_4582);
  and csa_tree_add_12_51_groupi_g16816(csa_tree_add_12_51_groupi_n_4961 ,csa_tree_add_12_51_groupi_n_4677 ,csa_tree_add_12_51_groupi_n_4845);
  or csa_tree_add_12_51_groupi_g16817(csa_tree_add_12_51_groupi_n_4960 ,csa_tree_add_12_51_groupi_n_4677 ,csa_tree_add_12_51_groupi_n_4845);
  nor csa_tree_add_12_51_groupi_g16818(csa_tree_add_12_51_groupi_n_4959 ,csa_tree_add_12_51_groupi_n_4069 ,csa_tree_add_12_51_groupi_n_4835);
  nor csa_tree_add_12_51_groupi_g16819(csa_tree_add_12_51_groupi_n_4958 ,csa_tree_add_12_51_groupi_n_3464 ,csa_tree_add_12_51_groupi_n_4826);
  nor csa_tree_add_12_51_groupi_g16820(csa_tree_add_12_51_groupi_n_4957 ,csa_tree_add_12_51_groupi_n_3438 ,csa_tree_add_12_51_groupi_n_4827);
  nor csa_tree_add_12_51_groupi_g16821(csa_tree_add_12_51_groupi_n_4956 ,csa_tree_add_12_51_groupi_n_3454 ,csa_tree_add_12_51_groupi_n_4828);
  nor csa_tree_add_12_51_groupi_g16822(csa_tree_add_12_51_groupi_n_4955 ,csa_tree_add_12_51_groupi_n_3873 ,csa_tree_add_12_51_groupi_n_4829);
  nor csa_tree_add_12_51_groupi_g16823(csa_tree_add_12_51_groupi_n_4954 ,csa_tree_add_12_51_groupi_n_3862 ,csa_tree_add_12_51_groupi_n_4830);
  nor csa_tree_add_12_51_groupi_g16824(csa_tree_add_12_51_groupi_n_4953 ,csa_tree_add_12_51_groupi_n_3895 ,csa_tree_add_12_51_groupi_n_4833);
  nor csa_tree_add_12_51_groupi_g16825(csa_tree_add_12_51_groupi_n_4952 ,csa_tree_add_12_51_groupi_n_3928 ,csa_tree_add_12_51_groupi_n_4834);
  nor csa_tree_add_12_51_groupi_g16826(csa_tree_add_12_51_groupi_n_4951 ,csa_tree_add_12_51_groupi_n_3885 ,csa_tree_add_12_51_groupi_n_4831);
  nor csa_tree_add_12_51_groupi_g16827(csa_tree_add_12_51_groupi_n_4950 ,csa_tree_add_12_51_groupi_n_4065 ,csa_tree_add_12_51_groupi_n_4873);
  nor csa_tree_add_12_51_groupi_g16828(csa_tree_add_12_51_groupi_n_4949 ,csa_tree_add_12_51_groupi_n_4104 ,csa_tree_add_12_51_groupi_n_4836);
  nor csa_tree_add_12_51_groupi_g16829(csa_tree_add_12_51_groupi_n_4948 ,csa_tree_add_12_51_groupi_n_3892 ,csa_tree_add_12_51_groupi_n_4832);
  nor csa_tree_add_12_51_groupi_g16830(csa_tree_add_12_51_groupi_n_4947 ,csa_tree_add_12_51_groupi_n_4060 ,csa_tree_add_12_51_groupi_n_4825);
  nor csa_tree_add_12_51_groupi_g16831(csa_tree_add_12_51_groupi_n_4946 ,csa_tree_add_12_51_groupi_n_4063 ,csa_tree_add_12_51_groupi_n_4838);
  nor csa_tree_add_12_51_groupi_g16832(csa_tree_add_12_51_groupi_n_4945 ,csa_tree_add_12_51_groupi_n_4057 ,csa_tree_add_12_51_groupi_n_4875);
  or csa_tree_add_12_51_groupi_g16833(csa_tree_add_12_51_groupi_n_4989 ,csa_tree_add_12_51_groupi_n_4630 ,csa_tree_add_12_51_groupi_n_4837);
  not csa_tree_add_12_51_groupi_g16834(csa_tree_add_12_51_groupi_n_4934 ,csa_tree_add_12_51_groupi_n_4935);
  not csa_tree_add_12_51_groupi_g16835(csa_tree_add_12_51_groupi_n_4931 ,csa_tree_add_12_51_groupi_n_4932);
  not csa_tree_add_12_51_groupi_g16836(csa_tree_add_12_51_groupi_n_4923 ,csa_tree_add_12_51_groupi_n_4922);
  not csa_tree_add_12_51_groupi_g16837(csa_tree_add_12_51_groupi_n_4920 ,csa_tree_add_12_51_groupi_n_4921);
  not csa_tree_add_12_51_groupi_g16838(csa_tree_add_12_51_groupi_n_4919 ,csa_tree_add_12_51_groupi_n_4918);
  not csa_tree_add_12_51_groupi_g16839(csa_tree_add_12_51_groupi_n_4917 ,csa_tree_add_12_51_groupi_n_9);
  nor csa_tree_add_12_51_groupi_g16840(csa_tree_add_12_51_groupi_n_4913 ,csa_tree_add_12_51_groupi_n_48 ,csa_tree_add_12_51_groupi_n_813);
  and csa_tree_add_12_51_groupi_g16841(csa_tree_add_12_51_groupi_n_4912 ,csa_tree_add_12_51_groupi_n_4715 ,csa_tree_add_12_51_groupi_n_4847);
  or csa_tree_add_12_51_groupi_g16842(csa_tree_add_12_51_groupi_n_4911 ,csa_tree_add_12_51_groupi_n_4715 ,csa_tree_add_12_51_groupi_n_4847);
  nor csa_tree_add_12_51_groupi_g16843(csa_tree_add_12_51_groupi_n_4910 ,csa_tree_add_12_51_groupi_n_24 ,csa_tree_add_12_51_groupi_n_840);
  nor csa_tree_add_12_51_groupi_g16844(csa_tree_add_12_51_groupi_n_4909 ,csa_tree_add_12_51_groupi_n_57 ,csa_tree_add_12_51_groupi_n_839);
  nor csa_tree_add_12_51_groupi_g16845(csa_tree_add_12_51_groupi_n_4908 ,csa_tree_add_12_51_groupi_n_21 ,csa_tree_add_12_51_groupi_n_1044);
  nor csa_tree_add_12_51_groupi_g16846(csa_tree_add_12_51_groupi_n_4907 ,csa_tree_add_12_51_groupi_n_54 ,csa_tree_add_12_51_groupi_n_839);
  nor csa_tree_add_12_51_groupi_g16847(csa_tree_add_12_51_groupi_n_4906 ,csa_tree_add_12_51_groupi_n_33 ,csa_tree_add_12_51_groupi_n_813);
  nor csa_tree_add_12_51_groupi_g16848(csa_tree_add_12_51_groupi_n_4905 ,csa_tree_add_12_51_groupi_n_63 ,csa_tree_add_12_51_groupi_n_812);
  nor csa_tree_add_12_51_groupi_g16849(csa_tree_add_12_51_groupi_n_4904 ,csa_tree_add_12_51_groupi_n_30 ,csa_tree_add_12_51_groupi_n_1983);
  nor csa_tree_add_12_51_groupi_g16850(csa_tree_add_12_51_groupi_n_4903 ,csa_tree_add_12_51_groupi_n_39 ,csa_tree_add_12_51_groupi_n_840);
  nor csa_tree_add_12_51_groupi_g16851(csa_tree_add_12_51_groupi_n_4902 ,csa_tree_add_12_51_groupi_n_45 ,csa_tree_add_12_51_groupi_n_151);
  xnor csa_tree_add_12_51_groupi_g16852(csa_tree_add_12_51_groupi_n_4901 ,csa_tree_add_12_51_groupi_n_4761 ,csa_tree_add_12_51_groupi_n_4760);
  xnor csa_tree_add_12_51_groupi_g16853(csa_tree_add_12_51_groupi_n_4900 ,csa_tree_add_12_51_groupi_n_4674 ,csa_tree_add_12_51_groupi_n_4768);
  xnor csa_tree_add_12_51_groupi_g16854(csa_tree_add_12_51_groupi_n_4899 ,csa_tree_add_12_51_groupi_n_4757 ,csa_tree_add_12_51_groupi_n_4756);
  xnor csa_tree_add_12_51_groupi_g16855(csa_tree_add_12_51_groupi_n_4898 ,csa_tree_add_12_51_groupi_n_4769 ,csa_tree_add_12_51_groupi_n_3);
  xnor csa_tree_add_12_51_groupi_g16856(csa_tree_add_12_51_groupi_n_4897 ,csa_tree_add_12_51_groupi_n_4676 ,csa_tree_add_12_51_groupi_n_4767);
  xnor csa_tree_add_12_51_groupi_g16857(csa_tree_add_12_51_groupi_n_4896 ,csa_tree_add_12_51_groupi_n_4764 ,csa_tree_add_12_51_groupi_n_4763);
  xnor csa_tree_add_12_51_groupi_g16858(csa_tree_add_12_51_groupi_n_4895 ,csa_tree_add_12_51_groupi_n_4754 ,csa_tree_add_12_51_groupi_n_4762);
  xnor csa_tree_add_12_51_groupi_g16859(csa_tree_add_12_51_groupi_n_4894 ,csa_tree_add_12_51_groupi_n_4209 ,csa_tree_add_12_51_groupi_n_4817);
  xnor csa_tree_add_12_51_groupi_g16860(csa_tree_add_12_51_groupi_n_4944 ,csa_tree_add_12_51_groupi_n_4787 ,in3[8]);
  xnor csa_tree_add_12_51_groupi_g16861(csa_tree_add_12_51_groupi_n_4943 ,csa_tree_add_12_51_groupi_n_4775 ,in3[5]);
  xnor csa_tree_add_12_51_groupi_g16862(csa_tree_add_12_51_groupi_n_4942 ,csa_tree_add_12_51_groupi_n_1929 ,csa_tree_add_12_51_groupi_n_4780);
  xnor csa_tree_add_12_51_groupi_g16863(csa_tree_add_12_51_groupi_n_4941 ,csa_tree_add_12_51_groupi_n_4784 ,in2[8]);
  xnor csa_tree_add_12_51_groupi_g16864(csa_tree_add_12_51_groupi_n_4940 ,csa_tree_add_12_51_groupi_n_4783 ,in4[11]);
  xnor csa_tree_add_12_51_groupi_g16865(csa_tree_add_12_51_groupi_n_4939 ,csa_tree_add_12_51_groupi_n_4788 ,in3[2]);
  xnor csa_tree_add_12_51_groupi_g16866(csa_tree_add_12_51_groupi_n_4938 ,csa_tree_add_12_51_groupi_n_4720 ,csa_tree_add_12_51_groupi_n_4735);
  xnor csa_tree_add_12_51_groupi_g16867(csa_tree_add_12_51_groupi_n_4937 ,csa_tree_add_12_51_groupi_n_4781 ,in3[11]);
  xnor csa_tree_add_12_51_groupi_g16868(csa_tree_add_12_51_groupi_n_4936 ,csa_tree_add_12_51_groupi_n_4575 ,csa_tree_add_12_51_groupi_n_4739);
  xnor csa_tree_add_12_51_groupi_g16869(csa_tree_add_12_51_groupi_n_4935 ,csa_tree_add_12_51_groupi_n_4593 ,csa_tree_add_12_51_groupi_n_4731);
  xnor csa_tree_add_12_51_groupi_g16870(csa_tree_add_12_51_groupi_n_4933 ,csa_tree_add_12_51_groupi_n_4594 ,csa_tree_add_12_51_groupi_n_4738);
  xnor csa_tree_add_12_51_groupi_g16871(csa_tree_add_12_51_groupi_n_4932 ,csa_tree_add_12_51_groupi_n_4778 ,in2[5]);
  xnor csa_tree_add_12_51_groupi_g16872(csa_tree_add_12_51_groupi_n_4930 ,csa_tree_add_12_51_groupi_n_4785 ,in4[8]);
  xnor csa_tree_add_12_51_groupi_g16873(csa_tree_add_12_51_groupi_n_4929 ,csa_tree_add_12_51_groupi_n_4779 ,in2[11]);
  xnor csa_tree_add_12_51_groupi_g16874(csa_tree_add_12_51_groupi_n_4928 ,csa_tree_add_12_51_groupi_n_4716 ,csa_tree_add_12_51_groupi_n_4733);
  xnor csa_tree_add_12_51_groupi_g16875(csa_tree_add_12_51_groupi_n_4927 ,csa_tree_add_12_51_groupi_n_4717 ,csa_tree_add_12_51_groupi_n_4729);
  xnor csa_tree_add_12_51_groupi_g16876(csa_tree_add_12_51_groupi_n_4926 ,csa_tree_add_12_51_groupi_n_4726 ,csa_tree_add_12_51_groupi_n_4736);
  xnor csa_tree_add_12_51_groupi_g16877(csa_tree_add_12_51_groupi_n_4925 ,csa_tree_add_12_51_groupi_n_4718 ,csa_tree_add_12_51_groupi_n_4737);
  xnor csa_tree_add_12_51_groupi_g16878(csa_tree_add_12_51_groupi_n_4924 ,csa_tree_add_12_51_groupi_n_4591 ,csa_tree_add_12_51_groupi_n_4730);
  xnor csa_tree_add_12_51_groupi_g16879(csa_tree_add_12_51_groupi_n_4922 ,csa_tree_add_12_51_groupi_n_4777 ,csa_tree_add_12_51_groupi_n_1933);
  xnor csa_tree_add_12_51_groupi_g16880(csa_tree_add_12_51_groupi_n_4921 ,csa_tree_add_12_51_groupi_n_4310 ,csa_tree_add_12_51_groupi_n_4734);
  xnor csa_tree_add_12_51_groupi_g16881(csa_tree_add_12_51_groupi_n_4918 ,csa_tree_add_12_51_groupi_n_4776 ,in2[14]);
  xnor csa_tree_add_12_51_groupi_g16883(csa_tree_add_12_51_groupi_n_4916 ,csa_tree_add_12_51_groupi_n_4592 ,csa_tree_add_12_51_groupi_n_4732);
  xnor csa_tree_add_12_51_groupi_g16884(csa_tree_add_12_51_groupi_n_4915 ,csa_tree_add_12_51_groupi_n_4789 ,in4[2]);
  xnor csa_tree_add_12_51_groupi_g16885(csa_tree_add_12_51_groupi_n_4914 ,csa_tree_add_12_51_groupi_n_4786 ,in2[2]);
  not csa_tree_add_12_51_groupi_g16886(csa_tree_add_12_51_groupi_n_4883 ,csa_tree_add_12_51_groupi_n_4884);
  not csa_tree_add_12_51_groupi_g16887(csa_tree_add_12_51_groupi_n_4879 ,csa_tree_add_12_51_groupi_n_4880);
  not csa_tree_add_12_51_groupi_g16888(csa_tree_add_12_51_groupi_n_4877 ,csa_tree_add_12_51_groupi_n_4878);
  or csa_tree_add_12_51_groupi_g16889(csa_tree_add_12_51_groupi_n_4875 ,csa_tree_add_12_51_groupi_n_3307 ,csa_tree_add_12_51_groupi_n_4746);
  or csa_tree_add_12_51_groupi_g16890(csa_tree_add_12_51_groupi_n_4874 ,csa_tree_add_12_51_groupi_n_4757 ,csa_tree_add_12_51_groupi_n_4756);
  or csa_tree_add_12_51_groupi_g16891(csa_tree_add_12_51_groupi_n_4873 ,csa_tree_add_12_51_groupi_n_3362 ,csa_tree_add_12_51_groupi_n_4751);
  or csa_tree_add_12_51_groupi_g16892(csa_tree_add_12_51_groupi_n_4872 ,csa_tree_add_12_51_groupi_n_4673 ,csa_tree_add_12_51_groupi_n_4765);
  and csa_tree_add_12_51_groupi_g16893(csa_tree_add_12_51_groupi_n_4871 ,csa_tree_add_12_51_groupi_n_4673 ,csa_tree_add_12_51_groupi_n_4765);
  and csa_tree_add_12_51_groupi_g16894(csa_tree_add_12_51_groupi_n_4870 ,csa_tree_add_12_51_groupi_n_4759 ,csa_tree_add_12_51_groupi_n_3);
  or csa_tree_add_12_51_groupi_g16895(csa_tree_add_12_51_groupi_n_4869 ,csa_tree_add_12_51_groupi_n_4761 ,csa_tree_add_12_51_groupi_n_4760);
  or csa_tree_add_12_51_groupi_g16896(csa_tree_add_12_51_groupi_n_4868 ,csa_tree_add_12_51_groupi_n_4676 ,csa_tree_add_12_51_groupi_n_4767);
  and csa_tree_add_12_51_groupi_g16897(csa_tree_add_12_51_groupi_n_4867 ,csa_tree_add_12_51_groupi_n_4761 ,csa_tree_add_12_51_groupi_n_4760);
  nor csa_tree_add_12_51_groupi_g16898(csa_tree_add_12_51_groupi_n_4866 ,csa_tree_add_12_51_groupi_n_4759 ,csa_tree_add_12_51_groupi_n_3);
  and csa_tree_add_12_51_groupi_g16899(csa_tree_add_12_51_groupi_n_4865 ,csa_tree_add_12_51_groupi_n_4676 ,csa_tree_add_12_51_groupi_n_4767);
  and csa_tree_add_12_51_groupi_g16900(csa_tree_add_12_51_groupi_n_4864 ,csa_tree_add_12_51_groupi_n_4674 ,csa_tree_add_12_51_groupi_n_4768);
  and csa_tree_add_12_51_groupi_g16901(csa_tree_add_12_51_groupi_n_4863 ,csa_tree_add_12_51_groupi_n_4764 ,csa_tree_add_12_51_groupi_n_4763);
  or csa_tree_add_12_51_groupi_g16902(csa_tree_add_12_51_groupi_n_4862 ,csa_tree_add_12_51_groupi_n_4764 ,csa_tree_add_12_51_groupi_n_4763);
  and csa_tree_add_12_51_groupi_g16903(csa_tree_add_12_51_groupi_n_4861 ,csa_tree_add_12_51_groupi_n_4757 ,csa_tree_add_12_51_groupi_n_4756);
  or csa_tree_add_12_51_groupi_g16904(csa_tree_add_12_51_groupi_n_4860 ,csa_tree_add_12_51_groupi_n_4674 ,csa_tree_add_12_51_groupi_n_4768);
  and csa_tree_add_12_51_groupi_g16905(csa_tree_add_12_51_groupi_n_4859 ,csa_tree_add_12_51_groupi_n_4754 ,csa_tree_add_12_51_groupi_n_4762);
  or csa_tree_add_12_51_groupi_g16906(csa_tree_add_12_51_groupi_n_4858 ,csa_tree_add_12_51_groupi_n_4754 ,csa_tree_add_12_51_groupi_n_4762);
  or csa_tree_add_12_51_groupi_g16907(csa_tree_add_12_51_groupi_n_4857 ,csa_tree_add_12_51_groupi_n_4675 ,csa_tree_add_12_51_groupi_n_4766);
  and csa_tree_add_12_51_groupi_g16908(csa_tree_add_12_51_groupi_n_4856 ,csa_tree_add_12_51_groupi_n_4675 ,csa_tree_add_12_51_groupi_n_4766);
  or csa_tree_add_12_51_groupi_g16909(csa_tree_add_12_51_groupi_n_4893 ,csa_tree_add_12_51_groupi_n_4622 ,csa_tree_add_12_51_groupi_n_4792);
  or csa_tree_add_12_51_groupi_g16910(csa_tree_add_12_51_groupi_n_4892 ,csa_tree_add_12_51_groupi_n_4693 ,csa_tree_add_12_51_groupi_n_4805);
  or csa_tree_add_12_51_groupi_g16911(csa_tree_add_12_51_groupi_n_4891 ,csa_tree_add_12_51_groupi_n_4700 ,csa_tree_add_12_51_groupi_n_4790);
  or csa_tree_add_12_51_groupi_g16912(csa_tree_add_12_51_groupi_n_4890 ,csa_tree_add_12_51_groupi_n_4688 ,csa_tree_add_12_51_groupi_n_4798);
  or csa_tree_add_12_51_groupi_g16913(csa_tree_add_12_51_groupi_n_4889 ,csa_tree_add_12_51_groupi_n_4613 ,csa_tree_add_12_51_groupi_n_4793);
  or csa_tree_add_12_51_groupi_g16914(csa_tree_add_12_51_groupi_n_4888 ,csa_tree_add_12_51_groupi_n_4702 ,csa_tree_add_12_51_groupi_n_4791);
  and csa_tree_add_12_51_groupi_g16915(csa_tree_add_12_51_groupi_n_4887 ,csa_tree_add_12_51_groupi_n_2428 ,csa_tree_add_12_51_groupi_n_4794);
  or csa_tree_add_12_51_groupi_g16916(csa_tree_add_12_51_groupi_n_4886 ,csa_tree_add_12_51_groupi_n_4685 ,csa_tree_add_12_51_groupi_n_4806);
  or csa_tree_add_12_51_groupi_g16917(csa_tree_add_12_51_groupi_n_4885 ,csa_tree_add_12_51_groupi_n_4699 ,csa_tree_add_12_51_groupi_n_4808);
  or csa_tree_add_12_51_groupi_g16918(csa_tree_add_12_51_groupi_n_4884 ,csa_tree_add_12_51_groupi_n_4691 ,csa_tree_add_12_51_groupi_n_4799);
  or csa_tree_add_12_51_groupi_g16919(csa_tree_add_12_51_groupi_n_4882 ,csa_tree_add_12_51_groupi_n_4689 ,csa_tree_add_12_51_groupi_n_4812);
  or csa_tree_add_12_51_groupi_g16920(csa_tree_add_12_51_groupi_n_4881 ,csa_tree_add_12_51_groupi_n_4697 ,csa_tree_add_12_51_groupi_n_4807);
  or csa_tree_add_12_51_groupi_g16921(csa_tree_add_12_51_groupi_n_4880 ,csa_tree_add_12_51_groupi_n_4706 ,csa_tree_add_12_51_groupi_n_4814);
  or csa_tree_add_12_51_groupi_g16922(csa_tree_add_12_51_groupi_n_4878 ,csa_tree_add_12_51_groupi_n_4686 ,csa_tree_add_12_51_groupi_n_4803);
  or csa_tree_add_12_51_groupi_g16923(csa_tree_add_12_51_groupi_n_4876 ,csa_tree_add_12_51_groupi_n_4698 ,csa_tree_add_12_51_groupi_n_4815);
  not csa_tree_add_12_51_groupi_g16924(csa_tree_add_12_51_groupi_n_4843 ,csa_tree_add_12_51_groupi_n_4844);
  not csa_tree_add_12_51_groupi_g16925(csa_tree_add_12_51_groupi_n_4840 ,csa_tree_add_12_51_groupi_n_4841);
  or csa_tree_add_12_51_groupi_g16926(csa_tree_add_12_51_groupi_n_4838 ,csa_tree_add_12_51_groupi_n_3294 ,csa_tree_add_12_51_groupi_n_4745);
  and csa_tree_add_12_51_groupi_g16927(csa_tree_add_12_51_groupi_n_4837 ,csa_tree_add_12_51_groupi_n_4574 ,csa_tree_add_12_51_groupi_n_4817);
  or csa_tree_add_12_51_groupi_g16928(csa_tree_add_12_51_groupi_n_4836 ,csa_tree_add_12_51_groupi_n_3266 ,csa_tree_add_12_51_groupi_n_4740);
  or csa_tree_add_12_51_groupi_g16929(csa_tree_add_12_51_groupi_n_4835 ,csa_tree_add_12_51_groupi_n_3267 ,csa_tree_add_12_51_groupi_n_4741);
  or csa_tree_add_12_51_groupi_g16930(csa_tree_add_12_51_groupi_n_4834 ,csa_tree_add_12_51_groupi_n_3708 ,csa_tree_add_12_51_groupi_n_4750);
  or csa_tree_add_12_51_groupi_g16931(csa_tree_add_12_51_groupi_n_4833 ,csa_tree_add_12_51_groupi_n_3644 ,csa_tree_add_12_51_groupi_n_4749);
  or csa_tree_add_12_51_groupi_g16932(csa_tree_add_12_51_groupi_n_4832 ,csa_tree_add_12_51_groupi_n_3716 ,csa_tree_add_12_51_groupi_n_4748);
  or csa_tree_add_12_51_groupi_g16933(csa_tree_add_12_51_groupi_n_4831 ,csa_tree_add_12_51_groupi_n_3696 ,csa_tree_add_12_51_groupi_n_4747);
  or csa_tree_add_12_51_groupi_g16934(csa_tree_add_12_51_groupi_n_4830 ,csa_tree_add_12_51_groupi_n_3643 ,csa_tree_add_12_51_groupi_n_4743);
  or csa_tree_add_12_51_groupi_g16935(csa_tree_add_12_51_groupi_n_4829 ,csa_tree_add_12_51_groupi_n_3627 ,csa_tree_add_12_51_groupi_n_4742);
  or csa_tree_add_12_51_groupi_g16936(csa_tree_add_12_51_groupi_n_4828 ,csa_tree_add_12_51_groupi_n_2979 ,csa_tree_add_12_51_groupi_n_4752);
  or csa_tree_add_12_51_groupi_g16937(csa_tree_add_12_51_groupi_n_4827 ,csa_tree_add_12_51_groupi_n_3134 ,csa_tree_add_12_51_groupi_n_4816);
  or csa_tree_add_12_51_groupi_g16938(csa_tree_add_12_51_groupi_n_4826 ,csa_tree_add_12_51_groupi_n_3004 ,csa_tree_add_12_51_groupi_n_4753);
  or csa_tree_add_12_51_groupi_g16939(csa_tree_add_12_51_groupi_n_4825 ,csa_tree_add_12_51_groupi_n_3285 ,csa_tree_add_12_51_groupi_n_4744);
  xnor csa_tree_add_12_51_groupi_g16940(csa_tree_add_12_51_groupi_n_4824 ,csa_tree_add_12_51_groupi_n_4212 ,csa_tree_add_12_51_groupi_n_4680);
  xnor csa_tree_add_12_51_groupi_g16941(csa_tree_add_12_51_groupi_n_4823 ,csa_tree_add_12_51_groupi_n_4672 ,csa_tree_add_12_51_groupi_n_4129);
  xnor csa_tree_add_12_51_groupi_g16942(csa_tree_add_12_51_groupi_n_4822 ,csa_tree_add_12_51_groupi_n_4399 ,csa_tree_add_12_51_groupi_n_4683);
  xnor csa_tree_add_12_51_groupi_g16943(csa_tree_add_12_51_groupi_n_4821 ,csa_tree_add_12_51_groupi_n_4724 ,csa_tree_add_12_51_groupi_n_3511);
  xnor csa_tree_add_12_51_groupi_g16944(csa_tree_add_12_51_groupi_n_4820 ,csa_tree_add_12_51_groupi_n_4725 ,csa_tree_add_12_51_groupi_n_3230);
  xnor csa_tree_add_12_51_groupi_g16945(csa_tree_add_12_51_groupi_n_4819 ,csa_tree_add_12_51_groupi_n_4216 ,csa_tree_add_12_51_groupi_n_4670);
  xor csa_tree_add_12_51_groupi_g16946(csa_tree_add_12_51_groupi_n_4818 ,csa_tree_add_12_51_groupi_n_4491 ,csa_tree_add_12_51_groupi_n_4719);
  or csa_tree_add_12_51_groupi_g16947(csa_tree_add_12_51_groupi_n_4855 ,csa_tree_add_12_51_groupi_n_4570 ,csa_tree_add_12_51_groupi_n_4813);
  or csa_tree_add_12_51_groupi_g16948(csa_tree_add_12_51_groupi_n_4854 ,csa_tree_add_12_51_groupi_n_4452 ,csa_tree_add_12_51_groupi_n_4809);
  or csa_tree_add_12_51_groupi_g16949(csa_tree_add_12_51_groupi_n_4853 ,csa_tree_add_12_51_groupi_n_4455 ,csa_tree_add_12_51_groupi_n_4797);
  xnor csa_tree_add_12_51_groupi_g16950(csa_tree_add_12_51_groupi_n_4852 ,csa_tree_add_12_51_groupi_n_4681 ,csa_tree_add_12_51_groupi_n_4645);
  xnor csa_tree_add_12_51_groupi_g16951(csa_tree_add_12_51_groupi_n_4851 ,csa_tree_add_12_51_groupi_n_4584 ,csa_tree_add_12_51_groupi_n_4644);
  xnor csa_tree_add_12_51_groupi_g16952(csa_tree_add_12_51_groupi_n_4850 ,csa_tree_add_12_51_groupi_n_4407 ,csa_tree_add_12_51_groupi_n_4650);
  xnor csa_tree_add_12_51_groupi_g16953(csa_tree_add_12_51_groupi_n_4849 ,csa_tree_add_12_51_groupi_n_4414 ,csa_tree_add_12_51_groupi_n_4643);
  xnor csa_tree_add_12_51_groupi_g16954(csa_tree_add_12_51_groupi_n_4848 ,csa_tree_add_12_51_groupi_n_4684 ,csa_tree_add_12_51_groupi_n_3972);
  xnor csa_tree_add_12_51_groupi_g16955(csa_tree_add_12_51_groupi_n_4847 ,csa_tree_add_12_51_groupi_n_4682 ,csa_tree_add_12_51_groupi_n_4640);
  xnor csa_tree_add_12_51_groupi_g16956(csa_tree_add_12_51_groupi_n_4846 ,csa_tree_add_12_51_groupi_n_4412 ,csa_tree_add_12_51_groupi_n_4642);
  xnor csa_tree_add_12_51_groupi_g16957(csa_tree_add_12_51_groupi_n_4845 ,csa_tree_add_12_51_groupi_n_4460 ,csa_tree_add_12_51_groupi_n_4647);
  xnor csa_tree_add_12_51_groupi_g16958(csa_tree_add_12_51_groupi_n_4844 ,csa_tree_add_12_51_groupi_n_4585 ,csa_tree_add_12_51_groupi_n_4646);
  xnor csa_tree_add_12_51_groupi_g16959(csa_tree_add_12_51_groupi_n_4842 ,csa_tree_add_12_51_groupi_n_4404 ,csa_tree_add_12_51_groupi_n_4641);
  xnor csa_tree_add_12_51_groupi_g16960(csa_tree_add_12_51_groupi_n_4841 ,csa_tree_add_12_51_groupi_n_4402 ,csa_tree_add_12_51_groupi_n_4649);
  xnor csa_tree_add_12_51_groupi_g16961(csa_tree_add_12_51_groupi_n_4839 ,csa_tree_add_12_51_groupi_n_4721 ,csa_tree_add_12_51_groupi_n_2569);
  nor csa_tree_add_12_51_groupi_g16962(csa_tree_add_12_51_groupi_n_4816 ,csa_tree_add_12_51_groupi_n_1856 ,csa_tree_add_12_51_groupi_n_1031);
  and csa_tree_add_12_51_groupi_g16963(csa_tree_add_12_51_groupi_n_4815 ,csa_tree_add_12_51_groupi_n_4707 ,csa_tree_add_12_51_groupi_n_4717);
  and csa_tree_add_12_51_groupi_g16964(csa_tree_add_12_51_groupi_n_4814 ,csa_tree_add_12_51_groupi_n_4705 ,csa_tree_add_12_51_groupi_n_4718);
  and csa_tree_add_12_51_groupi_g16965(csa_tree_add_12_51_groupi_n_4813 ,csa_tree_add_12_51_groupi_n_4569 ,csa_tree_add_12_51_groupi_n_4682);
  and csa_tree_add_12_51_groupi_g16966(csa_tree_add_12_51_groupi_n_4812 ,csa_tree_add_12_51_groupi_n_4594 ,csa_tree_add_12_51_groupi_n_4701);
  or csa_tree_add_12_51_groupi_g16967(csa_tree_add_12_51_groupi_n_4811 ,csa_tree_add_12_51_groupi_n_2352 ,csa_tree_add_12_51_groupi_n_4671);
  nor csa_tree_add_12_51_groupi_g16968(csa_tree_add_12_51_groupi_n_4810 ,csa_tree_add_12_51_groupi_n_2150 ,csa_tree_add_12_51_groupi_n_4672);
  and csa_tree_add_12_51_groupi_g16969(csa_tree_add_12_51_groupi_n_4809 ,csa_tree_add_12_51_groupi_n_4390 ,csa_tree_add_12_51_groupi_n_4724);
  and csa_tree_add_12_51_groupi_g16970(csa_tree_add_12_51_groupi_n_4808 ,csa_tree_add_12_51_groupi_n_4592 ,csa_tree_add_12_51_groupi_n_4692);
  and csa_tree_add_12_51_groupi_g16971(csa_tree_add_12_51_groupi_n_4807 ,csa_tree_add_12_51_groupi_n_4696 ,csa_tree_add_12_51_groupi_n_4726);
  nor csa_tree_add_12_51_groupi_g16972(csa_tree_add_12_51_groupi_n_4806 ,csa_tree_add_12_51_groupi_n_1 ,csa_tree_add_12_51_groupi_n_4694);
  and csa_tree_add_12_51_groupi_g16973(csa_tree_add_12_51_groupi_n_4805 ,csa_tree_add_12_51_groupi_n_4709 ,csa_tree_add_12_51_groupi_n_4720);
  or csa_tree_add_12_51_groupi_g16974(csa_tree_add_12_51_groupi_n_4804 ,csa_tree_add_12_51_groupi_n_4212 ,csa_tree_add_12_51_groupi_n_4680);
  and csa_tree_add_12_51_groupi_g16975(csa_tree_add_12_51_groupi_n_4803 ,csa_tree_add_12_51_groupi_n_4591 ,csa_tree_add_12_51_groupi_n_4711);
  and csa_tree_add_12_51_groupi_g16976(csa_tree_add_12_51_groupi_n_4802 ,csa_tree_add_12_51_groupi_n_4212 ,csa_tree_add_12_51_groupi_n_4680);
  nor csa_tree_add_12_51_groupi_g16977(csa_tree_add_12_51_groupi_n_4801 ,csa_tree_add_12_51_groupi_n_4216 ,csa_tree_add_12_51_groupi_n_4669);
  or csa_tree_add_12_51_groupi_g16978(csa_tree_add_12_51_groupi_n_4800 ,csa_tree_add_12_51_groupi_n_4215 ,csa_tree_add_12_51_groupi_n_4670);
  and csa_tree_add_12_51_groupi_g16979(csa_tree_add_12_51_groupi_n_4799 ,csa_tree_add_12_51_groupi_n_4593 ,csa_tree_add_12_51_groupi_n_4690);
  and csa_tree_add_12_51_groupi_g16980(csa_tree_add_12_51_groupi_n_4798 ,csa_tree_add_12_51_groupi_n_4687 ,csa_tree_add_12_51_groupi_n_4716);
  and csa_tree_add_12_51_groupi_g16981(csa_tree_add_12_51_groupi_n_4797 ,csa_tree_add_12_51_groupi_n_4392 ,csa_tree_add_12_51_groupi_n_4725);
  or csa_tree_add_12_51_groupi_g16982(csa_tree_add_12_51_groupi_n_4796 ,csa_tree_add_12_51_groupi_n_4667 ,csa_tree_add_12_51_groupi_n_4714);
  nor csa_tree_add_12_51_groupi_g16983(csa_tree_add_12_51_groupi_n_4795 ,csa_tree_add_12_51_groupi_n_4668 ,csa_tree_add_12_51_groupi_n_4713);
  or csa_tree_add_12_51_groupi_g16984(csa_tree_add_12_51_groupi_n_4794 ,csa_tree_add_12_51_groupi_n_2429 ,csa_tree_add_12_51_groupi_n_4721);
  and csa_tree_add_12_51_groupi_g16985(csa_tree_add_12_51_groupi_n_4793 ,csa_tree_add_12_51_groupi_n_4615 ,csa_tree_add_12_51_groupi_n_4681);
  and csa_tree_add_12_51_groupi_g16986(csa_tree_add_12_51_groupi_n_4792 ,csa_tree_add_12_51_groupi_n_4623 ,csa_tree_add_12_51_groupi_n_4683);
  nor csa_tree_add_12_51_groupi_g16987(csa_tree_add_12_51_groupi_n_4791 ,csa_tree_add_12_51_groupi_n_4507 ,csa_tree_add_12_51_groupi_n_4703);
  nor csa_tree_add_12_51_groupi_g16988(csa_tree_add_12_51_groupi_n_4790 ,csa_tree_add_12_51_groupi_n_4499 ,csa_tree_add_12_51_groupi_n_4695);
  nor csa_tree_add_12_51_groupi_g16989(csa_tree_add_12_51_groupi_n_4789 ,csa_tree_add_12_51_groupi_n_3441 ,csa_tree_add_12_51_groupi_n_4652);
  nor csa_tree_add_12_51_groupi_g16990(csa_tree_add_12_51_groupi_n_4788 ,csa_tree_add_12_51_groupi_n_3451 ,csa_tree_add_12_51_groupi_n_4653);
  nor csa_tree_add_12_51_groupi_g16991(csa_tree_add_12_51_groupi_n_4787 ,csa_tree_add_12_51_groupi_n_3882 ,csa_tree_add_12_51_groupi_n_4660);
  nor csa_tree_add_12_51_groupi_g16992(csa_tree_add_12_51_groupi_n_4786 ,csa_tree_add_12_51_groupi_n_3440 ,csa_tree_add_12_51_groupi_n_4651);
  nor csa_tree_add_12_51_groupi_g16993(csa_tree_add_12_51_groupi_n_4785 ,csa_tree_add_12_51_groupi_n_3911 ,csa_tree_add_12_51_groupi_n_4661);
  nor csa_tree_add_12_51_groupi_g16994(csa_tree_add_12_51_groupi_n_4784 ,csa_tree_add_12_51_groupi_n_3898 ,csa_tree_add_12_51_groupi_n_4662);
  nor csa_tree_add_12_51_groupi_g16995(csa_tree_add_12_51_groupi_n_4783 ,csa_tree_add_12_51_groupi_n_3839 ,csa_tree_add_12_51_groupi_n_4657);
  nor csa_tree_add_12_51_groupi_g16996(csa_tree_add_12_51_groupi_n_4782 ,csa_tree_add_12_51_groupi_n_3899 ,csa_tree_add_12_51_groupi_n_4663);
  nor csa_tree_add_12_51_groupi_g16997(csa_tree_add_12_51_groupi_n_4781 ,csa_tree_add_12_51_groupi_n_3872 ,csa_tree_add_12_51_groupi_n_4658);
  nor csa_tree_add_12_51_groupi_g16998(csa_tree_add_12_51_groupi_n_4780 ,csa_tree_add_12_51_groupi_n_4097 ,csa_tree_add_12_51_groupi_n_4659);
  nor csa_tree_add_12_51_groupi_g16999(csa_tree_add_12_51_groupi_n_4779 ,csa_tree_add_12_51_groupi_n_3838 ,csa_tree_add_12_51_groupi_n_4656);
  nor csa_tree_add_12_51_groupi_g17000(csa_tree_add_12_51_groupi_n_4778 ,csa_tree_add_12_51_groupi_n_4062 ,csa_tree_add_12_51_groupi_n_4664);
  nor csa_tree_add_12_51_groupi_g17001(csa_tree_add_12_51_groupi_n_4777 ,csa_tree_add_12_51_groupi_n_4038 ,csa_tree_add_12_51_groupi_n_4710);
  nor csa_tree_add_12_51_groupi_g17002(csa_tree_add_12_51_groupi_n_4776 ,csa_tree_add_12_51_groupi_n_4109 ,csa_tree_add_12_51_groupi_n_4708);
  nor csa_tree_add_12_51_groupi_g17003(csa_tree_add_12_51_groupi_n_4775 ,csa_tree_add_12_51_groupi_n_4037 ,csa_tree_add_12_51_groupi_n_4704);
  or csa_tree_add_12_51_groupi_g17004(csa_tree_add_12_51_groupi_n_4817 ,csa_tree_add_12_51_groupi_n_4391 ,csa_tree_add_12_51_groupi_n_4655);
  or csa_tree_add_12_51_groupi_g17005(csa_tree_add_12_51_groupi_n_4774 ,csa_tree_add_12_51_groupi_n_3973 ,csa_tree_add_12_51_groupi_n_4684);
  not csa_tree_add_12_51_groupi_g17006(csa_tree_add_12_51_groupi_n_4759 ,csa_tree_add_12_51_groupi_n_4758);
  nor csa_tree_add_12_51_groupi_g17007(csa_tree_add_12_51_groupi_n_4753 ,csa_tree_add_12_51_groupi_n_1859 ,csa_tree_add_12_51_groupi_n_1034);
  nor csa_tree_add_12_51_groupi_g17008(csa_tree_add_12_51_groupi_n_4752 ,csa_tree_add_12_51_groupi_n_1850 ,csa_tree_add_12_51_groupi_n_175);
  nor csa_tree_add_12_51_groupi_g17009(csa_tree_add_12_51_groupi_n_4751 ,csa_tree_add_12_51_groupi_n_1871 ,csa_tree_add_12_51_groupi_n_1031);
  nor csa_tree_add_12_51_groupi_g17010(csa_tree_add_12_51_groupi_n_4750 ,csa_tree_add_12_51_groupi_n_1868 ,csa_tree_add_12_51_groupi_n_1032);
  nor csa_tree_add_12_51_groupi_g17011(csa_tree_add_12_51_groupi_n_4749 ,csa_tree_add_12_51_groupi_n_1880 ,csa_tree_add_12_51_groupi_n_1035);
  nor csa_tree_add_12_51_groupi_g17012(csa_tree_add_12_51_groupi_n_4748 ,csa_tree_add_12_51_groupi_n_1889 ,csa_tree_add_12_51_groupi_n_945);
  nor csa_tree_add_12_51_groupi_g17013(csa_tree_add_12_51_groupi_n_4747 ,csa_tree_add_12_51_groupi_n_1877 ,csa_tree_add_12_51_groupi_n_944);
  nor csa_tree_add_12_51_groupi_g17014(csa_tree_add_12_51_groupi_n_4746 ,csa_tree_add_12_51_groupi_n_1874 ,csa_tree_add_12_51_groupi_n_1032);
  nor csa_tree_add_12_51_groupi_g17015(csa_tree_add_12_51_groupi_n_4745 ,csa_tree_add_12_51_groupi_n_1862 ,csa_tree_add_12_51_groupi_n_944);
  nor csa_tree_add_12_51_groupi_g17016(csa_tree_add_12_51_groupi_n_4744 ,csa_tree_add_12_51_groupi_n_1865 ,csa_tree_add_12_51_groupi_n_1035);
  nor csa_tree_add_12_51_groupi_g17017(csa_tree_add_12_51_groupi_n_4743 ,csa_tree_add_12_51_groupi_n_1853 ,csa_tree_add_12_51_groupi_n_1034);
  nor csa_tree_add_12_51_groupi_g17018(csa_tree_add_12_51_groupi_n_4742 ,csa_tree_add_12_51_groupi_n_1883 ,csa_tree_add_12_51_groupi_n_1980);
  nor csa_tree_add_12_51_groupi_g17019(csa_tree_add_12_51_groupi_n_4741 ,csa_tree_add_12_51_groupi_n_1847 ,csa_tree_add_12_51_groupi_n_945);
  nor csa_tree_add_12_51_groupi_g17020(csa_tree_add_12_51_groupi_n_4740 ,csa_tree_add_12_51_groupi_n_1886 ,csa_tree_add_12_51_groupi_n_175);
  xnor csa_tree_add_12_51_groupi_g17021(csa_tree_add_12_51_groupi_n_4739 ,csa_tree_add_12_51_groupi_n_1 ,csa_tree_add_12_51_groupi_n_4577);
  xnor csa_tree_add_12_51_groupi_g17022(csa_tree_add_12_51_groupi_n_4738 ,csa_tree_add_12_51_groupi_n_4588 ,csa_tree_add_12_51_groupi_n_4587);
  xnor csa_tree_add_12_51_groupi_g17023(csa_tree_add_12_51_groupi_n_4737 ,csa_tree_add_12_51_groupi_n_4410 ,csa_tree_add_12_51_groupi_n_4637);
  xnor csa_tree_add_12_51_groupi_g17024(csa_tree_add_12_51_groupi_n_4736 ,csa_tree_add_12_51_groupi_n_4415 ,csa_tree_add_12_51_groupi_n_4638);
  xnor csa_tree_add_12_51_groupi_g17025(csa_tree_add_12_51_groupi_n_4735 ,csa_tree_add_12_51_groupi_n_4406 ,csa_tree_add_12_51_groupi_n_4635);
  xnor csa_tree_add_12_51_groupi_g17026(csa_tree_add_12_51_groupi_n_4734 ,csa_tree_add_12_51_groupi_n_4639 ,csa_tree_add_12_51_groupi_n_3513);
  xnor csa_tree_add_12_51_groupi_g17027(csa_tree_add_12_51_groupi_n_4733 ,csa_tree_add_12_51_groupi_n_4409 ,csa_tree_add_12_51_groupi_n_4632);
  xnor csa_tree_add_12_51_groupi_g17028(csa_tree_add_12_51_groupi_n_4732 ,csa_tree_add_12_51_groupi_n_4590 ,csa_tree_add_12_51_groupi_n_4589);
  xnor csa_tree_add_12_51_groupi_g17029(csa_tree_add_12_51_groupi_n_4731 ,csa_tree_add_12_51_groupi_n_4580 ,csa_tree_add_12_51_groupi_n_4579);
  xnor csa_tree_add_12_51_groupi_g17030(csa_tree_add_12_51_groupi_n_4730 ,csa_tree_add_12_51_groupi_n_4581 ,csa_tree_add_12_51_groupi_n_4578);
  xnor csa_tree_add_12_51_groupi_g17031(csa_tree_add_12_51_groupi_n_4729 ,csa_tree_add_12_51_groupi_n_4395 ,csa_tree_add_12_51_groupi_n_4636);
  xnor csa_tree_add_12_51_groupi_g17032(csa_tree_add_12_51_groupi_n_4773 ,csa_tree_add_12_51_groupi_n_4606 ,in3[5]);
  xnor csa_tree_add_12_51_groupi_g17033(csa_tree_add_12_51_groupi_n_4772 ,csa_tree_add_12_51_groupi_n_4598 ,in3[14]);
  xnor csa_tree_add_12_51_groupi_g17034(csa_tree_add_12_51_groupi_n_4771 ,csa_tree_add_12_51_groupi_n_4599 ,in3[8]);
  xnor csa_tree_add_12_51_groupi_g17035(csa_tree_add_12_51_groupi_n_4770 ,csa_tree_add_12_51_groupi_n_4604 ,in3[11]);
  xnor csa_tree_add_12_51_groupi_g17036(csa_tree_add_12_51_groupi_n_4769 ,csa_tree_add_12_51_groupi_n_100 ,csa_tree_add_12_51_groupi_n_4601);
  xnor csa_tree_add_12_51_groupi_g17037(csa_tree_add_12_51_groupi_n_4768 ,csa_tree_add_12_51_groupi_n_4546 ,csa_tree_add_12_51_groupi_n_4550);
  xnor csa_tree_add_12_51_groupi_g17038(csa_tree_add_12_51_groupi_n_4767 ,csa_tree_add_12_51_groupi_n_4500 ,csa_tree_add_12_51_groupi_n_4551);
  xnor csa_tree_add_12_51_groupi_g17039(csa_tree_add_12_51_groupi_n_4766 ,csa_tree_add_12_51_groupi_n_4548 ,csa_tree_add_12_51_groupi_n_4549);
  xnor csa_tree_add_12_51_groupi_g17040(csa_tree_add_12_51_groupi_n_4765 ,csa_tree_add_12_51_groupi_n_4544 ,csa_tree_add_12_51_groupi_n_4553);
  xnor csa_tree_add_12_51_groupi_g17041(csa_tree_add_12_51_groupi_n_4764 ,csa_tree_add_12_51_groupi_n_4603 ,in4[11]);
  xnor csa_tree_add_12_51_groupi_g17042(csa_tree_add_12_51_groupi_n_4763 ,csa_tree_add_12_51_groupi_n_4609 ,in2[11]);
  xnor csa_tree_add_12_51_groupi_g17043(csa_tree_add_12_51_groupi_n_4762 ,csa_tree_add_12_51_groupi_n_4607 ,in2[14]);
  xnor csa_tree_add_12_51_groupi_g17044(csa_tree_add_12_51_groupi_n_4761 ,csa_tree_add_12_51_groupi_n_4597 ,in4[5]);
  xnor csa_tree_add_12_51_groupi_g17045(csa_tree_add_12_51_groupi_n_4760 ,csa_tree_add_12_51_groupi_n_4595 ,in2[5]);
  xnor csa_tree_add_12_51_groupi_g17047(csa_tree_add_12_51_groupi_n_4758 ,csa_tree_add_12_51_groupi_n_4600 ,in4[2]);
  xnor csa_tree_add_12_51_groupi_g17048(csa_tree_add_12_51_groupi_n_4757 ,csa_tree_add_12_51_groupi_n_4605 ,in4[8]);
  xnor csa_tree_add_12_51_groupi_g17049(csa_tree_add_12_51_groupi_n_4756 ,csa_tree_add_12_51_groupi_n_4608 ,in2[8]);
  xnor csa_tree_add_12_51_groupi_g17050(csa_tree_add_12_51_groupi_n_4755 ,csa_tree_add_12_51_groupi_n_4396 ,csa_tree_add_12_51_groupi_n_4552);
  xnor csa_tree_add_12_51_groupi_g17051(csa_tree_add_12_51_groupi_n_4754 ,csa_tree_add_12_51_groupi_n_4596 ,in4[14]);
  not csa_tree_add_12_51_groupi_g17052(csa_tree_add_12_51_groupi_n_4728 ,csa_tree_add_12_51_groupi_n_4727);
  not csa_tree_add_12_51_groupi_g17053(csa_tree_add_12_51_groupi_n_4723 ,csa_tree_add_12_51_groupi_n_4722);
  not csa_tree_add_12_51_groupi_g17054(csa_tree_add_12_51_groupi_n_4713 ,csa_tree_add_12_51_groupi_n_4714);
  or csa_tree_add_12_51_groupi_g17055(csa_tree_add_12_51_groupi_n_4711 ,csa_tree_add_12_51_groupi_n_4581 ,csa_tree_add_12_51_groupi_n_4578);
  or csa_tree_add_12_51_groupi_g17056(csa_tree_add_12_51_groupi_n_4710 ,csa_tree_add_12_51_groupi_n_3311 ,csa_tree_add_12_51_groupi_n_4559);
  or csa_tree_add_12_51_groupi_g17057(csa_tree_add_12_51_groupi_n_4709 ,csa_tree_add_12_51_groupi_n_4406 ,csa_tree_add_12_51_groupi_n_4635);
  or csa_tree_add_12_51_groupi_g17058(csa_tree_add_12_51_groupi_n_4708 ,csa_tree_add_12_51_groupi_n_3339 ,csa_tree_add_12_51_groupi_n_4562);
  or csa_tree_add_12_51_groupi_g17059(csa_tree_add_12_51_groupi_n_4707 ,csa_tree_add_12_51_groupi_n_4395 ,csa_tree_add_12_51_groupi_n_4636);
  and csa_tree_add_12_51_groupi_g17060(csa_tree_add_12_51_groupi_n_4706 ,csa_tree_add_12_51_groupi_n_4410 ,csa_tree_add_12_51_groupi_n_4637);
  or csa_tree_add_12_51_groupi_g17061(csa_tree_add_12_51_groupi_n_4705 ,csa_tree_add_12_51_groupi_n_4410 ,csa_tree_add_12_51_groupi_n_4637);
  or csa_tree_add_12_51_groupi_g17062(csa_tree_add_12_51_groupi_n_4704 ,csa_tree_add_12_51_groupi_n_3383 ,csa_tree_add_12_51_groupi_n_4565);
  nor csa_tree_add_12_51_groupi_g17063(csa_tree_add_12_51_groupi_n_4703 ,csa_tree_add_12_51_groupi_n_4405 ,csa_tree_add_12_51_groupi_n_4584);
  and csa_tree_add_12_51_groupi_g17064(csa_tree_add_12_51_groupi_n_4702 ,csa_tree_add_12_51_groupi_n_4405 ,csa_tree_add_12_51_groupi_n_4584);
  or csa_tree_add_12_51_groupi_g17065(csa_tree_add_12_51_groupi_n_4701 ,csa_tree_add_12_51_groupi_n_4588 ,csa_tree_add_12_51_groupi_n_4587);
  and csa_tree_add_12_51_groupi_g17066(csa_tree_add_12_51_groupi_n_4700 ,csa_tree_add_12_51_groupi_n_4411 ,csa_tree_add_12_51_groupi_n_4585);
  and csa_tree_add_12_51_groupi_g17067(csa_tree_add_12_51_groupi_n_4699 ,csa_tree_add_12_51_groupi_n_4590 ,csa_tree_add_12_51_groupi_n_4589);
  and csa_tree_add_12_51_groupi_g17068(csa_tree_add_12_51_groupi_n_4698 ,csa_tree_add_12_51_groupi_n_4395 ,csa_tree_add_12_51_groupi_n_4636);
  and csa_tree_add_12_51_groupi_g17069(csa_tree_add_12_51_groupi_n_4697 ,csa_tree_add_12_51_groupi_n_4415 ,csa_tree_add_12_51_groupi_n_4638);
  or csa_tree_add_12_51_groupi_g17070(csa_tree_add_12_51_groupi_n_4696 ,csa_tree_add_12_51_groupi_n_4415 ,csa_tree_add_12_51_groupi_n_4638);
  nor csa_tree_add_12_51_groupi_g17071(csa_tree_add_12_51_groupi_n_4695 ,csa_tree_add_12_51_groupi_n_4411 ,csa_tree_add_12_51_groupi_n_4585);
  and csa_tree_add_12_51_groupi_g17072(csa_tree_add_12_51_groupi_n_4694 ,csa_tree_add_12_51_groupi_n_4577 ,csa_tree_add_12_51_groupi_n_4576);
  and csa_tree_add_12_51_groupi_g17073(csa_tree_add_12_51_groupi_n_4693 ,csa_tree_add_12_51_groupi_n_4406 ,csa_tree_add_12_51_groupi_n_4635);
  or csa_tree_add_12_51_groupi_g17074(csa_tree_add_12_51_groupi_n_4692 ,csa_tree_add_12_51_groupi_n_4590 ,csa_tree_add_12_51_groupi_n_4589);
  and csa_tree_add_12_51_groupi_g17075(csa_tree_add_12_51_groupi_n_4691 ,csa_tree_add_12_51_groupi_n_4580 ,csa_tree_add_12_51_groupi_n_4579);
  or csa_tree_add_12_51_groupi_g17076(csa_tree_add_12_51_groupi_n_4690 ,csa_tree_add_12_51_groupi_n_4580 ,csa_tree_add_12_51_groupi_n_4579);
  and csa_tree_add_12_51_groupi_g17077(csa_tree_add_12_51_groupi_n_4689 ,csa_tree_add_12_51_groupi_n_4588 ,csa_tree_add_12_51_groupi_n_4587);
  and csa_tree_add_12_51_groupi_g17078(csa_tree_add_12_51_groupi_n_4688 ,csa_tree_add_12_51_groupi_n_4409 ,csa_tree_add_12_51_groupi_n_4632);
  or csa_tree_add_12_51_groupi_g17079(csa_tree_add_12_51_groupi_n_4687 ,csa_tree_add_12_51_groupi_n_4409 ,csa_tree_add_12_51_groupi_n_4632);
  and csa_tree_add_12_51_groupi_g17080(csa_tree_add_12_51_groupi_n_4686 ,csa_tree_add_12_51_groupi_n_4581 ,csa_tree_add_12_51_groupi_n_4578);
  nor csa_tree_add_12_51_groupi_g17081(csa_tree_add_12_51_groupi_n_4685 ,csa_tree_add_12_51_groupi_n_4577 ,csa_tree_add_12_51_groupi_n_4576);
  or csa_tree_add_12_51_groupi_g17082(csa_tree_add_12_51_groupi_n_4727 ,csa_tree_add_12_51_groupi_n_4531 ,csa_tree_add_12_51_groupi_n_4624);
  or csa_tree_add_12_51_groupi_g17083(csa_tree_add_12_51_groupi_n_4726 ,csa_tree_add_12_51_groupi_n_4526 ,csa_tree_add_12_51_groupi_n_4618);
  or csa_tree_add_12_51_groupi_g17084(csa_tree_add_12_51_groupi_n_4725 ,csa_tree_add_12_51_groupi_n_4265 ,csa_tree_add_12_51_groupi_n_4617);
  or csa_tree_add_12_51_groupi_g17085(csa_tree_add_12_51_groupi_n_4724 ,csa_tree_add_12_51_groupi_n_4267 ,csa_tree_add_12_51_groupi_n_4620);
  or csa_tree_add_12_51_groupi_g17086(csa_tree_add_12_51_groupi_n_4722 ,csa_tree_add_12_51_groupi_n_4528 ,csa_tree_add_12_51_groupi_n_4616);
  and csa_tree_add_12_51_groupi_g17087(csa_tree_add_12_51_groupi_n_4721 ,csa_tree_add_12_51_groupi_n_2459 ,csa_tree_add_12_51_groupi_n_4612);
  or csa_tree_add_12_51_groupi_g17088(csa_tree_add_12_51_groupi_n_4720 ,csa_tree_add_12_51_groupi_n_4509 ,csa_tree_add_12_51_groupi_n_4621);
  or csa_tree_add_12_51_groupi_g17089(csa_tree_add_12_51_groupi_n_4719 ,csa_tree_add_12_51_groupi_n_4532 ,csa_tree_add_12_51_groupi_n_4625);
  or csa_tree_add_12_51_groupi_g17090(csa_tree_add_12_51_groupi_n_4718 ,csa_tree_add_12_51_groupi_n_4535 ,csa_tree_add_12_51_groupi_n_4626);
  or csa_tree_add_12_51_groupi_g17091(csa_tree_add_12_51_groupi_n_4717 ,csa_tree_add_12_51_groupi_n_4520 ,csa_tree_add_12_51_groupi_n_4628);
  or csa_tree_add_12_51_groupi_g17092(csa_tree_add_12_51_groupi_n_4716 ,csa_tree_add_12_51_groupi_n_4514 ,csa_tree_add_12_51_groupi_n_4611);
  or csa_tree_add_12_51_groupi_g17093(csa_tree_add_12_51_groupi_n_4715 ,csa_tree_add_12_51_groupi_n_4521 ,csa_tree_add_12_51_groupi_n_4614);
  or csa_tree_add_12_51_groupi_g17094(csa_tree_add_12_51_groupi_n_4714 ,csa_tree_add_12_51_groupi_n_4438 ,csa_tree_add_12_51_groupi_n_4619);
  or csa_tree_add_12_51_groupi_g17095(csa_tree_add_12_51_groupi_n_4712 ,csa_tree_add_12_51_groupi_n_4518 ,csa_tree_add_12_51_groupi_n_4610);
  not csa_tree_add_12_51_groupi_g17096(csa_tree_add_12_51_groupi_n_4679 ,csa_tree_add_12_51_groupi_n_4678);
  not csa_tree_add_12_51_groupi_g17097(csa_tree_add_12_51_groupi_n_4671 ,csa_tree_add_12_51_groupi_n_4672);
  not csa_tree_add_12_51_groupi_g17098(csa_tree_add_12_51_groupi_n_4669 ,csa_tree_add_12_51_groupi_n_4670);
  not csa_tree_add_12_51_groupi_g17099(csa_tree_add_12_51_groupi_n_4667 ,csa_tree_add_12_51_groupi_n_4668);
  or csa_tree_add_12_51_groupi_g17100(csa_tree_add_12_51_groupi_n_4664 ,csa_tree_add_12_51_groupi_n_3287 ,csa_tree_add_12_51_groupi_n_4558);
  or csa_tree_add_12_51_groupi_g17101(csa_tree_add_12_51_groupi_n_4663 ,csa_tree_add_12_51_groupi_n_3656 ,csa_tree_add_12_51_groupi_n_4563);
  or csa_tree_add_12_51_groupi_g17102(csa_tree_add_12_51_groupi_n_4662 ,csa_tree_add_12_51_groupi_n_3584 ,csa_tree_add_12_51_groupi_n_4564);
  or csa_tree_add_12_51_groupi_g17103(csa_tree_add_12_51_groupi_n_4661 ,csa_tree_add_12_51_groupi_n_3665 ,csa_tree_add_12_51_groupi_n_4561);
  or csa_tree_add_12_51_groupi_g17104(csa_tree_add_12_51_groupi_n_4660 ,csa_tree_add_12_51_groupi_n_3635 ,csa_tree_add_12_51_groupi_n_4560);
  or csa_tree_add_12_51_groupi_g17105(csa_tree_add_12_51_groupi_n_4659 ,csa_tree_add_12_51_groupi_n_3091 ,csa_tree_add_12_51_groupi_n_4556);
  or csa_tree_add_12_51_groupi_g17106(csa_tree_add_12_51_groupi_n_4658 ,csa_tree_add_12_51_groupi_n_3636 ,csa_tree_add_12_51_groupi_n_4557);
  or csa_tree_add_12_51_groupi_g17107(csa_tree_add_12_51_groupi_n_4657 ,csa_tree_add_12_51_groupi_n_3587 ,csa_tree_add_12_51_groupi_n_4555);
  or csa_tree_add_12_51_groupi_g17108(csa_tree_add_12_51_groupi_n_4656 ,csa_tree_add_12_51_groupi_n_3657 ,csa_tree_add_12_51_groupi_n_4554);
  and csa_tree_add_12_51_groupi_g17109(csa_tree_add_12_51_groupi_n_4655 ,csa_tree_add_12_51_groupi_n_4393 ,csa_tree_add_12_51_groupi_n_4639);
  xnor csa_tree_add_12_51_groupi_g17110(out3[0] ,csa_tree_add_12_51_groupi_n_4138 ,csa_tree_add_12_51_groupi_n_4472);
  or csa_tree_add_12_51_groupi_g17111(csa_tree_add_12_51_groupi_n_4653 ,csa_tree_add_12_51_groupi_n_3122 ,csa_tree_add_12_51_groupi_n_4568);
  or csa_tree_add_12_51_groupi_g17112(csa_tree_add_12_51_groupi_n_4652 ,csa_tree_add_12_51_groupi_n_3093 ,csa_tree_add_12_51_groupi_n_4567);
  or csa_tree_add_12_51_groupi_g17113(csa_tree_add_12_51_groupi_n_4651 ,csa_tree_add_12_51_groupi_n_3172 ,csa_tree_add_12_51_groupi_n_4566);
  xnor csa_tree_add_12_51_groupi_g17114(csa_tree_add_12_51_groupi_n_4650 ,csa_tree_add_12_51_groupi_n_4394 ,csa_tree_add_12_51_groupi_n_4504);
  xnor csa_tree_add_12_51_groupi_g17115(csa_tree_add_12_51_groupi_n_4649 ,csa_tree_add_12_51_groupi_n_4218 ,csa_tree_add_12_51_groupi_n_4508);
  xnor csa_tree_add_12_51_groupi_g17116(csa_tree_add_12_51_groupi_n_4648 ,csa_tree_add_12_51_groupi_n_4207 ,csa_tree_add_12_51_groupi_n_4495);
  xnor csa_tree_add_12_51_groupi_g17117(csa_tree_add_12_51_groupi_n_4647 ,csa_tree_add_12_51_groupi_n_4309 ,csa_tree_add_12_51_groupi_n_4542);
  xor csa_tree_add_12_51_groupi_g17118(csa_tree_add_12_51_groupi_n_4646 ,csa_tree_add_12_51_groupi_n_4411 ,csa_tree_add_12_51_groupi_n_4499);
  xnor csa_tree_add_12_51_groupi_g17119(csa_tree_add_12_51_groupi_n_4645 ,csa_tree_add_12_51_groupi_n_4398 ,csa_tree_add_12_51_groupi_n_4488);
  xor csa_tree_add_12_51_groupi_g17120(csa_tree_add_12_51_groupi_n_4644 ,csa_tree_add_12_51_groupi_n_4405 ,csa_tree_add_12_51_groupi_n_4507);
  or csa_tree_add_12_51_groupi_g17121(csa_tree_add_12_51_groupi_n_4684 ,csa_tree_add_12_51_groupi_n_4259 ,csa_tree_add_12_51_groupi_n_4573);
  xnor csa_tree_add_12_51_groupi_g17122(csa_tree_add_12_51_groupi_n_4643 ,csa_tree_add_12_51_groupi_n_4408 ,csa_tree_add_12_51_groupi_n_4505);
  xnor csa_tree_add_12_51_groupi_g17123(csa_tree_add_12_51_groupi_n_4642 ,csa_tree_add_12_51_groupi_n_4413 ,csa_tree_add_12_51_groupi_n_4503);
  xnor csa_tree_add_12_51_groupi_g17124(csa_tree_add_12_51_groupi_n_4641 ,csa_tree_add_12_51_groupi_n_4403 ,csa_tree_add_12_51_groupi_n_4506);
  xnor csa_tree_add_12_51_groupi_g17125(csa_tree_add_12_51_groupi_n_4640 ,csa_tree_add_12_51_groupi_n_4400 ,csa_tree_add_12_51_groupi_n_4496);
  xnor csa_tree_add_12_51_groupi_g17126(csa_tree_add_12_51_groupi_n_4683 ,csa_tree_add_12_51_groupi_n_4225 ,csa_tree_add_12_51_groupi_n_4466);
  xnor csa_tree_add_12_51_groupi_g17127(csa_tree_add_12_51_groupi_n_4682 ,csa_tree_add_12_51_groupi_n_4221 ,csa_tree_add_12_51_groupi_n_4467);
  xnor csa_tree_add_12_51_groupi_g17128(csa_tree_add_12_51_groupi_n_4681 ,csa_tree_add_12_51_groupi_n_4204 ,csa_tree_add_12_51_groupi_n_4465);
  xnor csa_tree_add_12_51_groupi_g17129(csa_tree_add_12_51_groupi_n_4680 ,csa_tree_add_12_51_groupi_n_4501 ,csa_tree_add_12_51_groupi_n_4290);
  xnor csa_tree_add_12_51_groupi_g17130(csa_tree_add_12_51_groupi_n_4678 ,csa_tree_add_12_51_groupi_n_4545 ,csa_tree_add_12_51_groupi_n_4464);
  xnor csa_tree_add_12_51_groupi_g17131(csa_tree_add_12_51_groupi_n_4677 ,csa_tree_add_12_51_groupi_n_4323 ,csa_tree_add_12_51_groupi_n_4470);
  xnor csa_tree_add_12_51_groupi_g17132(csa_tree_add_12_51_groupi_n_4676 ,csa_tree_add_12_51_groupi_n_4304 ,csa_tree_add_12_51_groupi_n_4471);
  xnor csa_tree_add_12_51_groupi_g17133(csa_tree_add_12_51_groupi_n_4675 ,csa_tree_add_12_51_groupi_n_4302 ,csa_tree_add_12_51_groupi_n_4474);
  xnor csa_tree_add_12_51_groupi_g17134(csa_tree_add_12_51_groupi_n_4674 ,csa_tree_add_12_51_groupi_n_4318 ,csa_tree_add_12_51_groupi_n_4473);
  xnor csa_tree_add_12_51_groupi_g17135(csa_tree_add_12_51_groupi_n_4673 ,csa_tree_add_12_51_groupi_n_4321 ,csa_tree_add_12_51_groupi_n_4468);
  xnor csa_tree_add_12_51_groupi_g17136(csa_tree_add_12_51_groupi_n_4672 ,csa_tree_add_12_51_groupi_n_4543 ,csa_tree_add_12_51_groupi_n_4282);
  or csa_tree_add_12_51_groupi_g17137(csa_tree_add_12_51_groupi_n_4670 ,csa_tree_add_12_51_groupi_n_4479 ,csa_tree_add_12_51_groupi_n_4631);
  xnor csa_tree_add_12_51_groupi_g17138(csa_tree_add_12_51_groupi_n_4668 ,csa_tree_add_12_51_groupi_n_4228 ,csa_tree_add_12_51_groupi_n_4469);
  xnor csa_tree_add_12_51_groupi_g17139(csa_tree_add_12_51_groupi_n_4666 ,csa_tree_add_12_51_groupi_n_4502 ,csa_tree_add_12_51_groupi_n_4289);
  xnor csa_tree_add_12_51_groupi_g17140(csa_tree_add_12_51_groupi_n_4665 ,csa_tree_add_12_51_groupi_n_4547 ,csa_tree_add_12_51_groupi_n_2560);
  not csa_tree_add_12_51_groupi_g17141(csa_tree_add_12_51_groupi_n_4634 ,csa_tree_add_12_51_groupi_n_4633);
  and csa_tree_add_12_51_groupi_g17142(csa_tree_add_12_51_groupi_n_4631 ,csa_tree_add_12_51_groupi_n_4486 ,csa_tree_add_12_51_groupi_n_4508);
  nor csa_tree_add_12_51_groupi_g17143(csa_tree_add_12_51_groupi_n_4630 ,csa_tree_add_12_51_groupi_n_4209 ,csa_tree_add_12_51_groupi_n_4497);
  or csa_tree_add_12_51_groupi_g17144(csa_tree_add_12_51_groupi_n_4629 ,csa_tree_add_12_51_groupi_n_4206 ,csa_tree_add_12_51_groupi_n_4495);
  and csa_tree_add_12_51_groupi_g17145(csa_tree_add_12_51_groupi_n_4628 ,csa_tree_add_12_51_groupi_n_4538 ,csa_tree_add_12_51_groupi_n_4548);
  nor csa_tree_add_12_51_groupi_g17146(csa_tree_add_12_51_groupi_n_4627 ,csa_tree_add_12_51_groupi_n_4207 ,csa_tree_add_12_51_groupi_n_4494);
  and csa_tree_add_12_51_groupi_g17147(csa_tree_add_12_51_groupi_n_4626 ,csa_tree_add_12_51_groupi_n_4534 ,csa_tree_add_12_51_groupi_n_4544);
  nor csa_tree_add_12_51_groupi_g17148(csa_tree_add_12_51_groupi_n_4625 ,csa_tree_add_12_51_groupi_n_4416 ,csa_tree_add_12_51_groupi_n_4529);
  and csa_tree_add_12_51_groupi_g17149(csa_tree_add_12_51_groupi_n_4624 ,csa_tree_add_12_51_groupi_n_4530 ,csa_tree_add_12_51_groupi_n_4506);
  or csa_tree_add_12_51_groupi_g17150(csa_tree_add_12_51_groupi_n_4623 ,csa_tree_add_12_51_groupi_n_4399 ,csa_tree_add_12_51_groupi_n_4541);
  and csa_tree_add_12_51_groupi_g17151(csa_tree_add_12_51_groupi_n_4622 ,csa_tree_add_12_51_groupi_n_4399 ,csa_tree_add_12_51_groupi_n_4541);
  and csa_tree_add_12_51_groupi_g17152(csa_tree_add_12_51_groupi_n_4621 ,csa_tree_add_12_51_groupi_n_4510 ,csa_tree_add_12_51_groupi_n_4542);
  and csa_tree_add_12_51_groupi_g17153(csa_tree_add_12_51_groupi_n_4620 ,csa_tree_add_12_51_groupi_n_4266 ,csa_tree_add_12_51_groupi_n_4502);
  and csa_tree_add_12_51_groupi_g17154(csa_tree_add_12_51_groupi_n_4619 ,csa_tree_add_12_51_groupi_n_4440 ,csa_tree_add_12_51_groupi_n_4545);
  and csa_tree_add_12_51_groupi_g17155(csa_tree_add_12_51_groupi_n_4618 ,csa_tree_add_12_51_groupi_n_4527 ,csa_tree_add_12_51_groupi_n_4500);
  and csa_tree_add_12_51_groupi_g17156(csa_tree_add_12_51_groupi_n_4617 ,csa_tree_add_12_51_groupi_n_4268 ,csa_tree_add_12_51_groupi_n_4501);
  and csa_tree_add_12_51_groupi_g17157(csa_tree_add_12_51_groupi_n_4616 ,csa_tree_add_12_51_groupi_n_4519 ,csa_tree_add_12_51_groupi_n_4504);
  or csa_tree_add_12_51_groupi_g17158(csa_tree_add_12_51_groupi_n_4615 ,csa_tree_add_12_51_groupi_n_4398 ,csa_tree_add_12_51_groupi_n_4488);
  and csa_tree_add_12_51_groupi_g17159(csa_tree_add_12_51_groupi_n_4614 ,csa_tree_add_12_51_groupi_n_4523 ,csa_tree_add_12_51_groupi_n_4505);
  and csa_tree_add_12_51_groupi_g17160(csa_tree_add_12_51_groupi_n_4613 ,csa_tree_add_12_51_groupi_n_4398 ,csa_tree_add_12_51_groupi_n_4488);
  or csa_tree_add_12_51_groupi_g17161(csa_tree_add_12_51_groupi_n_4612 ,csa_tree_add_12_51_groupi_n_2447 ,csa_tree_add_12_51_groupi_n_4547);
  and csa_tree_add_12_51_groupi_g17162(csa_tree_add_12_51_groupi_n_4611 ,csa_tree_add_12_51_groupi_n_4516 ,csa_tree_add_12_51_groupi_n_4546);
  and csa_tree_add_12_51_groupi_g17163(csa_tree_add_12_51_groupi_n_4610 ,csa_tree_add_12_51_groupi_n_4540 ,csa_tree_add_12_51_groupi_n_4503);
  nor csa_tree_add_12_51_groupi_g17164(csa_tree_add_12_51_groupi_n_4609 ,csa_tree_add_12_51_groupi_n_3846 ,csa_tree_add_12_51_groupi_n_4481);
  nor csa_tree_add_12_51_groupi_g17165(csa_tree_add_12_51_groupi_n_4608 ,csa_tree_add_12_51_groupi_n_3912 ,csa_tree_add_12_51_groupi_n_4480);
  nor csa_tree_add_12_51_groupi_g17166(csa_tree_add_12_51_groupi_n_4607 ,csa_tree_add_12_51_groupi_n_4043 ,csa_tree_add_12_51_groupi_n_4522);
  nor csa_tree_add_12_51_groupi_g17167(csa_tree_add_12_51_groupi_n_4606 ,csa_tree_add_12_51_groupi_n_4059 ,csa_tree_add_12_51_groupi_n_4512);
  nor csa_tree_add_12_51_groupi_g17168(csa_tree_add_12_51_groupi_n_4605 ,csa_tree_add_12_51_groupi_n_3913 ,csa_tree_add_12_51_groupi_n_4475);
  nor csa_tree_add_12_51_groupi_g17169(csa_tree_add_12_51_groupi_n_4604 ,csa_tree_add_12_51_groupi_n_4098 ,csa_tree_add_12_51_groupi_n_4484);
  nor csa_tree_add_12_51_groupi_g17170(csa_tree_add_12_51_groupi_n_4603 ,csa_tree_add_12_51_groupi_n_3843 ,csa_tree_add_12_51_groupi_n_4482);
  nor csa_tree_add_12_51_groupi_g17171(csa_tree_add_12_51_groupi_n_4602 ,csa_tree_add_12_51_groupi_n_3461 ,csa_tree_add_12_51_groupi_n_4477);
  nor csa_tree_add_12_51_groupi_g17172(csa_tree_add_12_51_groupi_n_4601 ,csa_tree_add_12_51_groupi_n_3470 ,csa_tree_add_12_51_groupi_n_4476);
  nor csa_tree_add_12_51_groupi_g17173(csa_tree_add_12_51_groupi_n_4600 ,csa_tree_add_12_51_groupi_n_3458 ,csa_tree_add_12_51_groupi_n_4478);
  nor csa_tree_add_12_51_groupi_g17174(csa_tree_add_12_51_groupi_n_4599 ,csa_tree_add_12_51_groupi_n_3875 ,csa_tree_add_12_51_groupi_n_4485);
  nor csa_tree_add_12_51_groupi_g17175(csa_tree_add_12_51_groupi_n_4598 ,csa_tree_add_12_51_groupi_n_4096 ,csa_tree_add_12_51_groupi_n_4483);
  nor csa_tree_add_12_51_groupi_g17176(csa_tree_add_12_51_groupi_n_4597 ,csa_tree_add_12_51_groupi_n_4058 ,csa_tree_add_12_51_groupi_n_4533);
  nor csa_tree_add_12_51_groupi_g17177(csa_tree_add_12_51_groupi_n_4596 ,csa_tree_add_12_51_groupi_n_4111 ,csa_tree_add_12_51_groupi_n_4515);
  nor csa_tree_add_12_51_groupi_g17178(csa_tree_add_12_51_groupi_n_4595 ,csa_tree_add_12_51_groupi_n_4107 ,csa_tree_add_12_51_groupi_n_4537);
  or csa_tree_add_12_51_groupi_g17179(csa_tree_add_12_51_groupi_n_4639 ,csa_tree_add_12_51_groupi_n_4261 ,csa_tree_add_12_51_groupi_n_4511);
  or csa_tree_add_12_51_groupi_g17180(csa_tree_add_12_51_groupi_n_4638 ,csa_tree_add_12_51_groupi_n_4439 ,csa_tree_add_12_51_groupi_n_4513);
  or csa_tree_add_12_51_groupi_g17181(csa_tree_add_12_51_groupi_n_4637 ,csa_tree_add_12_51_groupi_n_4451 ,csa_tree_add_12_51_groupi_n_4536);
  or csa_tree_add_12_51_groupi_g17182(csa_tree_add_12_51_groupi_n_4636 ,csa_tree_add_12_51_groupi_n_4454 ,csa_tree_add_12_51_groupi_n_4539);
  or csa_tree_add_12_51_groupi_g17183(csa_tree_add_12_51_groupi_n_4635 ,csa_tree_add_12_51_groupi_n_4435 ,csa_tree_add_12_51_groupi_n_4525);
  and csa_tree_add_12_51_groupi_g17184(csa_tree_add_12_51_groupi_n_4633 ,csa_tree_add_12_51_groupi_n_4337 ,csa_tree_add_12_51_groupi_n_4524);
  or csa_tree_add_12_51_groupi_g17185(csa_tree_add_12_51_groupi_n_4632 ,csa_tree_add_12_51_groupi_n_4432 ,csa_tree_add_12_51_groupi_n_4517);
  not csa_tree_add_12_51_groupi_g17186(csa_tree_add_12_51_groupi_n_4582 ,csa_tree_add_12_51_groupi_n_4583);
  not csa_tree_add_12_51_groupi_g17187(csa_tree_add_12_51_groupi_n_4576 ,csa_tree_add_12_51_groupi_n_4575);
  or csa_tree_add_12_51_groupi_g17188(csa_tree_add_12_51_groupi_n_4574 ,csa_tree_add_12_51_groupi_n_4208 ,csa_tree_add_12_51_groupi_n_4498);
  and csa_tree_add_12_51_groupi_g17189(csa_tree_add_12_51_groupi_n_4573 ,csa_tree_add_12_51_groupi_n_4258 ,csa_tree_add_12_51_groupi_n_4543);
  nor csa_tree_add_12_51_groupi_g17190(csa_tree_add_12_51_groupi_n_4572 ,csa_tree_add_12_51_groupi_n_4211 ,csa_tree_add_12_51_groupi_n_4492);
  or csa_tree_add_12_51_groupi_g17191(csa_tree_add_12_51_groupi_n_4571 ,csa_tree_add_12_51_groupi_n_4210 ,csa_tree_add_12_51_groupi_n_4493);
  and csa_tree_add_12_51_groupi_g17192(csa_tree_add_12_51_groupi_n_4570 ,csa_tree_add_12_51_groupi_n_4400 ,csa_tree_add_12_51_groupi_n_4496);
  or csa_tree_add_12_51_groupi_g17193(csa_tree_add_12_51_groupi_n_4569 ,csa_tree_add_12_51_groupi_n_4400 ,csa_tree_add_12_51_groupi_n_4496);
  nor csa_tree_add_12_51_groupi_g17194(csa_tree_add_12_51_groupi_n_4568 ,csa_tree_add_12_51_groupi_n_1825 ,csa_tree_add_12_51_groupi_n_1025);
  nor csa_tree_add_12_51_groupi_g17195(csa_tree_add_12_51_groupi_n_4567 ,csa_tree_add_12_51_groupi_n_1819 ,csa_tree_add_12_51_groupi_n_1028);
  nor csa_tree_add_12_51_groupi_g17196(csa_tree_add_12_51_groupi_n_4566 ,csa_tree_add_12_51_groupi_n_1821 ,csa_tree_add_12_51_groupi_n_165);
  nor csa_tree_add_12_51_groupi_g17197(csa_tree_add_12_51_groupi_n_4565 ,csa_tree_add_12_51_groupi_n_1827 ,csa_tree_add_12_51_groupi_n_1025);
  nor csa_tree_add_12_51_groupi_g17198(csa_tree_add_12_51_groupi_n_4564 ,csa_tree_add_12_51_groupi_n_1829 ,csa_tree_add_12_51_groupi_n_1026);
  nor csa_tree_add_12_51_groupi_g17199(csa_tree_add_12_51_groupi_n_4563 ,csa_tree_add_12_51_groupi_n_1823 ,csa_tree_add_12_51_groupi_n_1029);
  nor csa_tree_add_12_51_groupi_g17200(csa_tree_add_12_51_groupi_n_4562 ,csa_tree_add_12_51_groupi_n_1831 ,csa_tree_add_12_51_groupi_n_816);
  nor csa_tree_add_12_51_groupi_g17201(csa_tree_add_12_51_groupi_n_4561 ,csa_tree_add_12_51_groupi_n_1817 ,csa_tree_add_12_51_groupi_n_815);
  nor csa_tree_add_12_51_groupi_g17202(csa_tree_add_12_51_groupi_n_4560 ,csa_tree_add_12_51_groupi_n_1839 ,csa_tree_add_12_51_groupi_n_1026);
  nor csa_tree_add_12_51_groupi_g17203(csa_tree_add_12_51_groupi_n_4559 ,csa_tree_add_12_51_groupi_n_1835 ,csa_tree_add_12_51_groupi_n_815);
  nor csa_tree_add_12_51_groupi_g17204(csa_tree_add_12_51_groupi_n_4558 ,csa_tree_add_12_51_groupi_n_1845 ,csa_tree_add_12_51_groupi_n_1029);
  nor csa_tree_add_12_51_groupi_g17205(csa_tree_add_12_51_groupi_n_4557 ,csa_tree_add_12_51_groupi_n_1837 ,csa_tree_add_12_51_groupi_n_1028);
  nor csa_tree_add_12_51_groupi_g17206(csa_tree_add_12_51_groupi_n_4556 ,csa_tree_add_12_51_groupi_n_1841 ,csa_tree_add_12_51_groupi_n_1965);
  nor csa_tree_add_12_51_groupi_g17207(csa_tree_add_12_51_groupi_n_4555 ,csa_tree_add_12_51_groupi_n_1843 ,csa_tree_add_12_51_groupi_n_816);
  nor csa_tree_add_12_51_groupi_g17208(csa_tree_add_12_51_groupi_n_4554 ,csa_tree_add_12_51_groupi_n_1833 ,csa_tree_add_12_51_groupi_n_165);
  xnor csa_tree_add_12_51_groupi_g17209(csa_tree_add_12_51_groupi_n_4553 ,csa_tree_add_12_51_groupi_n_4459 ,csa_tree_add_12_51_groupi_n_4311);
  xnor csa_tree_add_12_51_groupi_g17210(csa_tree_add_12_51_groupi_n_4552 ,csa_tree_add_12_51_groupi_n_4416 ,csa_tree_add_12_51_groupi_n_4135);
  xnor csa_tree_add_12_51_groupi_g17211(csa_tree_add_12_51_groupi_n_4551 ,csa_tree_add_12_51_groupi_n_4458 ,csa_tree_add_12_51_groupi_n_4305);
  xnor csa_tree_add_12_51_groupi_g17212(csa_tree_add_12_51_groupi_n_4550 ,csa_tree_add_12_51_groupi_n_4461 ,csa_tree_add_12_51_groupi_n_4308);
  xnor csa_tree_add_12_51_groupi_g17213(csa_tree_add_12_51_groupi_n_4549 ,csa_tree_add_12_51_groupi_n_4457 ,csa_tree_add_12_51_groupi_n_4301);
  xnor csa_tree_add_12_51_groupi_g17214(csa_tree_add_12_51_groupi_n_4594 ,csa_tree_add_12_51_groupi_n_4418 ,in3[8]);
  xnor csa_tree_add_12_51_groupi_g17215(csa_tree_add_12_51_groupi_n_4593 ,csa_tree_add_12_51_groupi_n_4420 ,in3[11]);
  xnor csa_tree_add_12_51_groupi_g17216(csa_tree_add_12_51_groupi_n_4592 ,csa_tree_add_12_51_groupi_n_4427 ,in3[5]);
  xnor csa_tree_add_12_51_groupi_g17218(csa_tree_add_12_51_groupi_n_4591 ,csa_tree_add_12_51_groupi_n_4431 ,in3[14]);
  xnor csa_tree_add_12_51_groupi_g17219(csa_tree_add_12_51_groupi_n_4590 ,csa_tree_add_12_51_groupi_n_4419 ,in4[5]);
  xnor csa_tree_add_12_51_groupi_g17220(csa_tree_add_12_51_groupi_n_4589 ,csa_tree_add_12_51_groupi_n_4417 ,in2[5]);
  xnor csa_tree_add_12_51_groupi_g17221(csa_tree_add_12_51_groupi_n_4588 ,csa_tree_add_12_51_groupi_n_4429 ,in4[8]);
  xnor csa_tree_add_12_51_groupi_g17222(csa_tree_add_12_51_groupi_n_4587 ,csa_tree_add_12_51_groupi_n_4426 ,in2[8]);
  xnor csa_tree_add_12_51_groupi_g17223(csa_tree_add_12_51_groupi_n_4586 ,csa_tree_add_12_51_groupi_n_4463 ,csa_tree_add_12_51_groupi_n_4288);
  xnor csa_tree_add_12_51_groupi_g17224(csa_tree_add_12_51_groupi_n_4585 ,csa_tree_add_12_51_groupi_n_4359 ,csa_tree_add_12_51_groupi_n_4369);
  xnor csa_tree_add_12_51_groupi_g17225(csa_tree_add_12_51_groupi_n_4584 ,csa_tree_add_12_51_groupi_n_4360 ,csa_tree_add_12_51_groupi_n_4368);
  xnor csa_tree_add_12_51_groupi_g17226(csa_tree_add_12_51_groupi_n_4583 ,csa_tree_add_12_51_groupi_n_4462 ,csa_tree_add_12_51_groupi_n_4367);
  xnor csa_tree_add_12_51_groupi_g17227(csa_tree_add_12_51_groupi_n_4581 ,csa_tree_add_12_51_groupi_n_4428 ,in4[14]);
  xnor csa_tree_add_12_51_groupi_g17228(csa_tree_add_12_51_groupi_n_4580 ,csa_tree_add_12_51_groupi_n_4425 ,in4[11]);
  xnor csa_tree_add_12_51_groupi_g17229(csa_tree_add_12_51_groupi_n_4579 ,csa_tree_add_12_51_groupi_n_4421 ,in2[11]);
  xnor csa_tree_add_12_51_groupi_g17230(csa_tree_add_12_51_groupi_n_4578 ,csa_tree_add_12_51_groupi_n_4430 ,in2[14]);
  xnor csa_tree_add_12_51_groupi_g17231(csa_tree_add_12_51_groupi_n_4577 ,csa_tree_add_12_51_groupi_n_1927 ,csa_tree_add_12_51_groupi_n_4424);
  xnor csa_tree_add_12_51_groupi_g17232(csa_tree_add_12_51_groupi_n_4575 ,csa_tree_add_12_51_groupi_n_4423 ,in2[2]);
  or csa_tree_add_12_51_groupi_g17233(csa_tree_add_12_51_groupi_n_4540 ,csa_tree_add_12_51_groupi_n_4413 ,csa_tree_add_12_51_groupi_n_4412);
  nor csa_tree_add_12_51_groupi_g17234(csa_tree_add_12_51_groupi_n_4539 ,csa_tree_add_12_51_groupi_n_4324 ,csa_tree_add_12_51_groupi_n_4453);
  or csa_tree_add_12_51_groupi_g17235(csa_tree_add_12_51_groupi_n_4538 ,csa_tree_add_12_51_groupi_n_4457 ,csa_tree_add_12_51_groupi_n_4301);
  or csa_tree_add_12_51_groupi_g17236(csa_tree_add_12_51_groupi_n_4537 ,csa_tree_add_12_51_groupi_n_3333 ,csa_tree_add_12_51_groupi_n_4373);
  and csa_tree_add_12_51_groupi_g17237(csa_tree_add_12_51_groupi_n_4536 ,csa_tree_add_12_51_groupi_n_4321 ,csa_tree_add_12_51_groupi_n_4450);
  and csa_tree_add_12_51_groupi_g17238(csa_tree_add_12_51_groupi_n_4535 ,csa_tree_add_12_51_groupi_n_4459 ,csa_tree_add_12_51_groupi_n_4311);
  or csa_tree_add_12_51_groupi_g17239(csa_tree_add_12_51_groupi_n_4534 ,csa_tree_add_12_51_groupi_n_4459 ,csa_tree_add_12_51_groupi_n_4311);
  or csa_tree_add_12_51_groupi_g17240(csa_tree_add_12_51_groupi_n_4533 ,csa_tree_add_12_51_groupi_n_3304 ,csa_tree_add_12_51_groupi_n_4374);
  nor csa_tree_add_12_51_groupi_g17241(csa_tree_add_12_51_groupi_n_4532 ,csa_tree_add_12_51_groupi_n_4135 ,csa_tree_add_12_51_groupi_n_4397);
  and csa_tree_add_12_51_groupi_g17242(csa_tree_add_12_51_groupi_n_4531 ,csa_tree_add_12_51_groupi_n_4403 ,csa_tree_add_12_51_groupi_n_4404);
  or csa_tree_add_12_51_groupi_g17243(csa_tree_add_12_51_groupi_n_4530 ,csa_tree_add_12_51_groupi_n_4403 ,csa_tree_add_12_51_groupi_n_4404);
  and csa_tree_add_12_51_groupi_g17244(csa_tree_add_12_51_groupi_n_4529 ,csa_tree_add_12_51_groupi_n_4135 ,csa_tree_add_12_51_groupi_n_4397);
  and csa_tree_add_12_51_groupi_g17245(csa_tree_add_12_51_groupi_n_4528 ,csa_tree_add_12_51_groupi_n_4394 ,csa_tree_add_12_51_groupi_n_4407);
  or csa_tree_add_12_51_groupi_g17246(csa_tree_add_12_51_groupi_n_4527 ,csa_tree_add_12_51_groupi_n_4458 ,csa_tree_add_12_51_groupi_n_4305);
  and csa_tree_add_12_51_groupi_g17247(csa_tree_add_12_51_groupi_n_4526 ,csa_tree_add_12_51_groupi_n_4458 ,csa_tree_add_12_51_groupi_n_4305);
  and csa_tree_add_12_51_groupi_g17248(csa_tree_add_12_51_groupi_n_4525 ,csa_tree_add_12_51_groupi_n_4323 ,csa_tree_add_12_51_groupi_n_4456);
  or csa_tree_add_12_51_groupi_g17249(csa_tree_add_12_51_groupi_n_4524 ,csa_tree_add_12_51_groupi_n_4338 ,csa_tree_add_12_51_groupi_n_4462);
  or csa_tree_add_12_51_groupi_g17250(csa_tree_add_12_51_groupi_n_4523 ,csa_tree_add_12_51_groupi_n_4408 ,csa_tree_add_12_51_groupi_n_4414);
  or csa_tree_add_12_51_groupi_g17251(csa_tree_add_12_51_groupi_n_4522 ,csa_tree_add_12_51_groupi_n_3335 ,csa_tree_add_12_51_groupi_n_4378);
  and csa_tree_add_12_51_groupi_g17252(csa_tree_add_12_51_groupi_n_4521 ,csa_tree_add_12_51_groupi_n_4408 ,csa_tree_add_12_51_groupi_n_4414);
  and csa_tree_add_12_51_groupi_g17253(csa_tree_add_12_51_groupi_n_4520 ,csa_tree_add_12_51_groupi_n_4457 ,csa_tree_add_12_51_groupi_n_4301);
  or csa_tree_add_12_51_groupi_g17254(csa_tree_add_12_51_groupi_n_4519 ,csa_tree_add_12_51_groupi_n_4394 ,csa_tree_add_12_51_groupi_n_4407);
  and csa_tree_add_12_51_groupi_g17255(csa_tree_add_12_51_groupi_n_4518 ,csa_tree_add_12_51_groupi_n_4413 ,csa_tree_add_12_51_groupi_n_4412);
  and csa_tree_add_12_51_groupi_g17256(csa_tree_add_12_51_groupi_n_4517 ,csa_tree_add_12_51_groupi_n_4318 ,csa_tree_add_12_51_groupi_n_4436);
  or csa_tree_add_12_51_groupi_g17257(csa_tree_add_12_51_groupi_n_4516 ,csa_tree_add_12_51_groupi_n_4461 ,csa_tree_add_12_51_groupi_n_4308);
  or csa_tree_add_12_51_groupi_g17258(csa_tree_add_12_51_groupi_n_4515 ,csa_tree_add_12_51_groupi_n_3350 ,csa_tree_add_12_51_groupi_n_4379);
  and csa_tree_add_12_51_groupi_g17259(csa_tree_add_12_51_groupi_n_4514 ,csa_tree_add_12_51_groupi_n_4461 ,csa_tree_add_12_51_groupi_n_4308);
  nor csa_tree_add_12_51_groupi_g17260(csa_tree_add_12_51_groupi_n_4513 ,csa_tree_add_12_51_groupi_n_4322 ,csa_tree_add_12_51_groupi_n_4434);
  or csa_tree_add_12_51_groupi_g17261(csa_tree_add_12_51_groupi_n_4512 ,csa_tree_add_12_51_groupi_n_3368 ,csa_tree_add_12_51_groupi_n_4381);
  and csa_tree_add_12_51_groupi_g17262(csa_tree_add_12_51_groupi_n_4511 ,csa_tree_add_12_51_groupi_n_4260 ,csa_tree_add_12_51_groupi_n_4463);
  or csa_tree_add_12_51_groupi_g17263(csa_tree_add_12_51_groupi_n_4510 ,csa_tree_add_12_51_groupi_n_4460 ,csa_tree_add_12_51_groupi_n_4309);
  and csa_tree_add_12_51_groupi_g17264(csa_tree_add_12_51_groupi_n_4509 ,csa_tree_add_12_51_groupi_n_4460 ,csa_tree_add_12_51_groupi_n_4309);
  or csa_tree_add_12_51_groupi_g17265(csa_tree_add_12_51_groupi_n_4548 ,csa_tree_add_12_51_groupi_n_4356 ,csa_tree_add_12_51_groupi_n_4449);
  and csa_tree_add_12_51_groupi_g17266(csa_tree_add_12_51_groupi_n_4547 ,csa_tree_add_12_51_groupi_n_2430 ,csa_tree_add_12_51_groupi_n_4437);
  or csa_tree_add_12_51_groupi_g17267(csa_tree_add_12_51_groupi_n_4546 ,csa_tree_add_12_51_groupi_n_4345 ,csa_tree_add_12_51_groupi_n_4433);
  or csa_tree_add_12_51_groupi_g17268(csa_tree_add_12_51_groupi_n_4545 ,csa_tree_add_12_51_groupi_n_4331 ,csa_tree_add_12_51_groupi_n_4442);
  or csa_tree_add_12_51_groupi_g17269(csa_tree_add_12_51_groupi_n_4544 ,csa_tree_add_12_51_groupi_n_4353 ,csa_tree_add_12_51_groupi_n_4448);
  or csa_tree_add_12_51_groupi_g17270(csa_tree_add_12_51_groupi_n_4543 ,csa_tree_add_12_51_groupi_n_3803 ,csa_tree_add_12_51_groupi_n_4443);
  or csa_tree_add_12_51_groupi_g17271(csa_tree_add_12_51_groupi_n_4542 ,csa_tree_add_12_51_groupi_n_4293 ,csa_tree_add_12_51_groupi_n_4441);
  or csa_tree_add_12_51_groupi_g17272(csa_tree_add_12_51_groupi_n_4541 ,csa_tree_add_12_51_groupi_n_4275 ,csa_tree_add_12_51_groupi_n_4445);
  not csa_tree_add_12_51_groupi_g17273(csa_tree_add_12_51_groupi_n_4497 ,csa_tree_add_12_51_groupi_n_4498);
  not csa_tree_add_12_51_groupi_g17274(csa_tree_add_12_51_groupi_n_4494 ,csa_tree_add_12_51_groupi_n_4495);
  not csa_tree_add_12_51_groupi_g17275(csa_tree_add_12_51_groupi_n_4492 ,csa_tree_add_12_51_groupi_n_4493);
  not csa_tree_add_12_51_groupi_g17276(csa_tree_add_12_51_groupi_n_4489 ,csa_tree_add_12_51_groupi_n_4490);
  or csa_tree_add_12_51_groupi_g17277(csa_tree_add_12_51_groupi_n_4486 ,csa_tree_add_12_51_groupi_n_4217 ,csa_tree_add_12_51_groupi_n_4402);
  or csa_tree_add_12_51_groupi_g17278(csa_tree_add_12_51_groupi_n_4485 ,csa_tree_add_12_51_groupi_n_3640 ,csa_tree_add_12_51_groupi_n_4376);
  or csa_tree_add_12_51_groupi_g17279(csa_tree_add_12_51_groupi_n_4484 ,csa_tree_add_12_51_groupi_n_3132 ,csa_tree_add_12_51_groupi_n_4375);
  or csa_tree_add_12_51_groupi_g17280(csa_tree_add_12_51_groupi_n_4483 ,csa_tree_add_12_51_groupi_n_3023 ,csa_tree_add_12_51_groupi_n_4372);
  or csa_tree_add_12_51_groupi_g17281(csa_tree_add_12_51_groupi_n_4482 ,csa_tree_add_12_51_groupi_n_3676 ,csa_tree_add_12_51_groupi_n_4370);
  or csa_tree_add_12_51_groupi_g17282(csa_tree_add_12_51_groupi_n_4481 ,csa_tree_add_12_51_groupi_n_3680 ,csa_tree_add_12_51_groupi_n_4371);
  or csa_tree_add_12_51_groupi_g17283(csa_tree_add_12_51_groupi_n_4480 ,csa_tree_add_12_51_groupi_n_3664 ,csa_tree_add_12_51_groupi_n_4380);
  nor csa_tree_add_12_51_groupi_g17284(csa_tree_add_12_51_groupi_n_4479 ,csa_tree_add_12_51_groupi_n_4218 ,csa_tree_add_12_51_groupi_n_4401);
  or csa_tree_add_12_51_groupi_g17285(csa_tree_add_12_51_groupi_n_4478 ,csa_tree_add_12_51_groupi_n_3058 ,csa_tree_add_12_51_groupi_n_4389);
  or csa_tree_add_12_51_groupi_g17286(csa_tree_add_12_51_groupi_n_4477 ,csa_tree_add_12_51_groupi_n_3154 ,csa_tree_add_12_51_groupi_n_4388);
  or csa_tree_add_12_51_groupi_g17287(csa_tree_add_12_51_groupi_n_4476 ,csa_tree_add_12_51_groupi_n_3173 ,csa_tree_add_12_51_groupi_n_4387);
  or csa_tree_add_12_51_groupi_g17288(csa_tree_add_12_51_groupi_n_4475 ,csa_tree_add_12_51_groupi_n_3617 ,csa_tree_add_12_51_groupi_n_4377);
  xor csa_tree_add_12_51_groupi_g17289(csa_tree_add_12_51_groupi_n_4474 ,csa_tree_add_12_51_groupi_n_4324 ,in5[14]);
  xnor csa_tree_add_12_51_groupi_g17290(csa_tree_add_12_51_groupi_n_4473 ,csa_tree_add_12_51_groupi_n_4306 ,in5[11]);
  xnor csa_tree_add_12_51_groupi_g17291(csa_tree_add_12_51_groupi_n_4472 ,csa_tree_add_12_51_groupi_n_4142 ,csa_tree_add_12_51_groupi_n_4314);
  xor csa_tree_add_12_51_groupi_g17292(csa_tree_add_12_51_groupi_n_4471 ,csa_tree_add_12_51_groupi_n_4322 ,in5[5]);
  xnor csa_tree_add_12_51_groupi_g17293(csa_tree_add_12_51_groupi_n_4470 ,csa_tree_add_12_51_groupi_n_4313 ,in5[2]);
  xnor csa_tree_add_12_51_groupi_g17294(csa_tree_add_12_51_groupi_n_4469 ,csa_tree_add_12_51_groupi_n_4365 ,csa_tree_add_12_51_groupi_n_2163);
  xnor csa_tree_add_12_51_groupi_g17295(csa_tree_add_12_51_groupi_n_4468 ,csa_tree_add_12_51_groupi_n_4303 ,in5[8]);
  xnor csa_tree_add_12_51_groupi_g17296(csa_tree_add_12_51_groupi_n_4467 ,csa_tree_add_12_51_groupi_n_4361 ,csa_tree_add_12_51_groupi_n_4219);
  xnor csa_tree_add_12_51_groupi_g17297(csa_tree_add_12_51_groupi_n_4466 ,csa_tree_add_12_51_groupi_n_4224 ,csa_tree_add_12_51_groupi_n_4358);
  xnor csa_tree_add_12_51_groupi_g17298(csa_tree_add_12_51_groupi_n_4465 ,csa_tree_add_12_51_groupi_n_4357 ,csa_tree_add_12_51_groupi_n_4205);
  xnor csa_tree_add_12_51_groupi_g17299(csa_tree_add_12_51_groupi_n_4464 ,csa_tree_add_12_51_groupi_n_4136 ,csa_tree_add_12_51_groupi_n_4312);
  or csa_tree_add_12_51_groupi_g17300(csa_tree_add_12_51_groupi_n_4508 ,csa_tree_add_12_51_groupi_n_4354 ,csa_tree_add_12_51_groupi_n_4447);
  and csa_tree_add_12_51_groupi_g17301(csa_tree_add_12_51_groupi_n_4507 ,csa_tree_add_12_51_groupi_n_4186 ,csa_tree_add_12_51_groupi_n_4384);
  xnor csa_tree_add_12_51_groupi_g17302(csa_tree_add_12_51_groupi_n_4506 ,csa_tree_add_12_51_groupi_n_4315 ,csa_tree_add_12_51_groupi_n_4286);
  xnor csa_tree_add_12_51_groupi_g17303(csa_tree_add_12_51_groupi_n_4505 ,csa_tree_add_12_51_groupi_n_4325 ,csa_tree_add_12_51_groupi_n_4283);
  xnor csa_tree_add_12_51_groupi_g17304(csa_tree_add_12_51_groupi_n_4504 ,csa_tree_add_12_51_groupi_n_4319 ,csa_tree_add_12_51_groupi_n_4285);
  xnor csa_tree_add_12_51_groupi_g17305(csa_tree_add_12_51_groupi_n_4503 ,csa_tree_add_12_51_groupi_n_4317 ,csa_tree_add_12_51_groupi_n_4284);
  or csa_tree_add_12_51_groupi_g17306(csa_tree_add_12_51_groupi_n_4502 ,csa_tree_add_12_51_groupi_n_3799 ,csa_tree_add_12_51_groupi_n_4446);
  or csa_tree_add_12_51_groupi_g17307(csa_tree_add_12_51_groupi_n_4501 ,csa_tree_add_12_51_groupi_n_3800 ,csa_tree_add_12_51_groupi_n_4444);
  or csa_tree_add_12_51_groupi_g17308(csa_tree_add_12_51_groupi_n_4500 ,csa_tree_add_12_51_groupi_n_4296 ,csa_tree_add_12_51_groupi_n_4386);
  and csa_tree_add_12_51_groupi_g17309(csa_tree_add_12_51_groupi_n_4499 ,csa_tree_add_12_51_groupi_n_4254 ,csa_tree_add_12_51_groupi_n_4385);
  xnor csa_tree_add_12_51_groupi_g17310(csa_tree_add_12_51_groupi_n_4498 ,csa_tree_add_12_51_groupi_n_4366 ,csa_tree_add_12_51_groupi_n_11);
  or csa_tree_add_12_51_groupi_g17311(csa_tree_add_12_51_groupi_n_4496 ,csa_tree_add_12_51_groupi_n_4202 ,csa_tree_add_12_51_groupi_n_4383);
  xnor csa_tree_add_12_51_groupi_g17312(csa_tree_add_12_51_groupi_n_4495 ,csa_tree_add_12_51_groupi_n_4363 ,csa_tree_add_12_51_groupi_n_12);
  xnor csa_tree_add_12_51_groupi_g17313(csa_tree_add_12_51_groupi_n_4493 ,csa_tree_add_12_51_groupi_n_4364 ,csa_tree_add_12_51_groupi_n_10);
  xnor csa_tree_add_12_51_groupi_g17314(csa_tree_add_12_51_groupi_n_4491 ,csa_tree_add_12_51_groupi_n_4237 ,csa_tree_add_12_51_groupi_n_4287);
  xnor csa_tree_add_12_51_groupi_g17315(csa_tree_add_12_51_groupi_n_4490 ,csa_tree_add_12_51_groupi_n_4227 ,csa_tree_add_12_51_groupi_n_4291);
  or csa_tree_add_12_51_groupi_g17316(csa_tree_add_12_51_groupi_n_4488 ,csa_tree_add_12_51_groupi_n_4199 ,csa_tree_add_12_51_groupi_n_4382);
  xnor csa_tree_add_12_51_groupi_g17317(csa_tree_add_12_51_groupi_n_4487 ,csa_tree_add_12_51_groupi_n_4362 ,csa_tree_add_12_51_groupi_n_2558);
  or csa_tree_add_12_51_groupi_g17318(csa_tree_add_12_51_groupi_n_4456 ,in5[2] ,csa_tree_add_12_51_groupi_n_4313);
  and csa_tree_add_12_51_groupi_g17319(csa_tree_add_12_51_groupi_n_4455 ,csa_tree_add_12_51_groupi_n_3231 ,csa_tree_add_12_51_groupi_n_4307);
  and csa_tree_add_12_51_groupi_g17320(csa_tree_add_12_51_groupi_n_4454 ,in5[14] ,csa_tree_add_12_51_groupi_n_4302);
  nor csa_tree_add_12_51_groupi_g17321(csa_tree_add_12_51_groupi_n_4453 ,in5[14] ,csa_tree_add_12_51_groupi_n_4302);
  and csa_tree_add_12_51_groupi_g17322(csa_tree_add_12_51_groupi_n_4452 ,csa_tree_add_12_51_groupi_n_3512 ,csa_tree_add_12_51_groupi_n_4300);
  and csa_tree_add_12_51_groupi_g17323(csa_tree_add_12_51_groupi_n_4451 ,in5[8] ,csa_tree_add_12_51_groupi_n_4303);
  or csa_tree_add_12_51_groupi_g17324(csa_tree_add_12_51_groupi_n_4450 ,in5[8] ,csa_tree_add_12_51_groupi_n_4303);
  and csa_tree_add_12_51_groupi_g17325(csa_tree_add_12_51_groupi_n_4449 ,csa_tree_add_12_51_groupi_n_4357 ,csa_tree_add_12_51_groupi_n_4352);
  and csa_tree_add_12_51_groupi_g17326(csa_tree_add_12_51_groupi_n_4448 ,csa_tree_add_12_51_groupi_n_4360 ,csa_tree_add_12_51_groupi_n_4351);
  and csa_tree_add_12_51_groupi_g17327(csa_tree_add_12_51_groupi_n_4447 ,csa_tree_add_12_51_groupi_n_4365 ,csa_tree_add_12_51_groupi_n_4347);
  and csa_tree_add_12_51_groupi_g17328(csa_tree_add_12_51_groupi_n_4446 ,csa_tree_add_12_51_groupi_n_3798 ,csa_tree_add_12_51_groupi_n_4366);
  and csa_tree_add_12_51_groupi_g17329(csa_tree_add_12_51_groupi_n_4445 ,csa_tree_add_12_51_groupi_n_4278 ,csa_tree_add_12_51_groupi_n_4314);
  and csa_tree_add_12_51_groupi_g17330(csa_tree_add_12_51_groupi_n_4444 ,csa_tree_add_12_51_groupi_n_3801 ,csa_tree_add_12_51_groupi_n_4364);
  and csa_tree_add_12_51_groupi_g17331(csa_tree_add_12_51_groupi_n_4443 ,csa_tree_add_12_51_groupi_n_3802 ,csa_tree_add_12_51_groupi_n_4363);
  nor csa_tree_add_12_51_groupi_g17332(csa_tree_add_12_51_groupi_n_4442 ,csa_tree_add_12_51_groupi_n_4184 ,csa_tree_add_12_51_groupi_n_4330);
  and csa_tree_add_12_51_groupi_g17333(csa_tree_add_12_51_groupi_n_4441 ,csa_tree_add_12_51_groupi_n_4358 ,csa_tree_add_12_51_groupi_n_4294);
  or csa_tree_add_12_51_groupi_g17334(csa_tree_add_12_51_groupi_n_4440 ,csa_tree_add_12_51_groupi_n_4136 ,csa_tree_add_12_51_groupi_n_4312);
  and csa_tree_add_12_51_groupi_g17335(csa_tree_add_12_51_groupi_n_4439 ,in5[5] ,csa_tree_add_12_51_groupi_n_4304);
  and csa_tree_add_12_51_groupi_g17336(csa_tree_add_12_51_groupi_n_4438 ,csa_tree_add_12_51_groupi_n_4136 ,csa_tree_add_12_51_groupi_n_4312);
  or csa_tree_add_12_51_groupi_g17337(csa_tree_add_12_51_groupi_n_4437 ,csa_tree_add_12_51_groupi_n_2421 ,csa_tree_add_12_51_groupi_n_4362);
  or csa_tree_add_12_51_groupi_g17338(csa_tree_add_12_51_groupi_n_4436 ,in5[11] ,csa_tree_add_12_51_groupi_n_4306);
  and csa_tree_add_12_51_groupi_g17339(csa_tree_add_12_51_groupi_n_4435 ,in5[2] ,csa_tree_add_12_51_groupi_n_4313);
  nor csa_tree_add_12_51_groupi_g17340(csa_tree_add_12_51_groupi_n_4434 ,in5[5] ,csa_tree_add_12_51_groupi_n_4304);
  and csa_tree_add_12_51_groupi_g17341(csa_tree_add_12_51_groupi_n_4433 ,csa_tree_add_12_51_groupi_n_4359 ,csa_tree_add_12_51_groupi_n_4343);
  and csa_tree_add_12_51_groupi_g17342(csa_tree_add_12_51_groupi_n_4432 ,in5[11] ,csa_tree_add_12_51_groupi_n_4306);
  nor csa_tree_add_12_51_groupi_g17343(csa_tree_add_12_51_groupi_n_4431 ,csa_tree_add_12_51_groupi_n_4071 ,csa_tree_add_12_51_groupi_n_4332);
  nor csa_tree_add_12_51_groupi_g17344(csa_tree_add_12_51_groupi_n_4430 ,csa_tree_add_12_51_groupi_n_3909 ,csa_tree_add_12_51_groupi_n_4334);
  nor csa_tree_add_12_51_groupi_g17345(csa_tree_add_12_51_groupi_n_4429 ,csa_tree_add_12_51_groupi_n_3889 ,csa_tree_add_12_51_groupi_n_4335);
  nor csa_tree_add_12_51_groupi_g17346(csa_tree_add_12_51_groupi_n_4428 ,csa_tree_add_12_51_groupi_n_4053 ,csa_tree_add_12_51_groupi_n_4329);
  nor csa_tree_add_12_51_groupi_g17347(csa_tree_add_12_51_groupi_n_4427 ,csa_tree_add_12_51_groupi_n_4055 ,csa_tree_add_12_51_groupi_n_4328);
  nor csa_tree_add_12_51_groupi_g17348(csa_tree_add_12_51_groupi_n_4426 ,csa_tree_add_12_51_groupi_n_3897 ,csa_tree_add_12_51_groupi_n_4336);
  nor csa_tree_add_12_51_groupi_g17349(csa_tree_add_12_51_groupi_n_4425 ,csa_tree_add_12_51_groupi_n_3836 ,csa_tree_add_12_51_groupi_n_4341);
  nor csa_tree_add_12_51_groupi_g17350(csa_tree_add_12_51_groupi_n_4424 ,csa_tree_add_12_51_groupi_n_3471 ,csa_tree_add_12_51_groupi_n_4292);
  nor csa_tree_add_12_51_groupi_g17351(csa_tree_add_12_51_groupi_n_4423 ,csa_tree_add_12_51_groupi_n_3443 ,csa_tree_add_12_51_groupi_n_4297);
  nor csa_tree_add_12_51_groupi_g17352(csa_tree_add_12_51_groupi_n_4422 ,csa_tree_add_12_51_groupi_n_3450 ,csa_tree_add_12_51_groupi_n_4298);
  nor csa_tree_add_12_51_groupi_g17353(csa_tree_add_12_51_groupi_n_4421 ,csa_tree_add_12_51_groupi_n_3835 ,csa_tree_add_12_51_groupi_n_4344);
  nor csa_tree_add_12_51_groupi_g17354(csa_tree_add_12_51_groupi_n_4420 ,csa_tree_add_12_51_groupi_n_3874 ,csa_tree_add_12_51_groupi_n_4340);
  nor csa_tree_add_12_51_groupi_g17355(csa_tree_add_12_51_groupi_n_4419 ,csa_tree_add_12_51_groupi_n_4056 ,csa_tree_add_12_51_groupi_n_4327);
  nor csa_tree_add_12_51_groupi_g17356(csa_tree_add_12_51_groupi_n_4418 ,csa_tree_add_12_51_groupi_n_3877 ,csa_tree_add_12_51_groupi_n_4339);
  nor csa_tree_add_12_51_groupi_g17357(csa_tree_add_12_51_groupi_n_4417 ,csa_tree_add_12_51_groupi_n_4040 ,csa_tree_add_12_51_groupi_n_4326);
  or csa_tree_add_12_51_groupi_g17358(csa_tree_add_12_51_groupi_n_4463 ,csa_tree_add_12_51_groupi_n_3821 ,csa_tree_add_12_51_groupi_n_4333);
  and csa_tree_add_12_51_groupi_g17359(csa_tree_add_12_51_groupi_n_4462 ,csa_tree_add_12_51_groupi_n_4262 ,csa_tree_add_12_51_groupi_n_4350);
  or csa_tree_add_12_51_groupi_g17360(csa_tree_add_12_51_groupi_n_4461 ,csa_tree_add_12_51_groupi_n_3484 ,csa_tree_add_12_51_groupi_n_4346);
  or csa_tree_add_12_51_groupi_g17361(csa_tree_add_12_51_groupi_n_4460 ,csa_tree_add_12_51_groupi_n_3487 ,csa_tree_add_12_51_groupi_n_4348);
  or csa_tree_add_12_51_groupi_g17362(csa_tree_add_12_51_groupi_n_4459 ,csa_tree_add_12_51_groupi_n_3491 ,csa_tree_add_12_51_groupi_n_4355);
  or csa_tree_add_12_51_groupi_g17363(csa_tree_add_12_51_groupi_n_4458 ,csa_tree_add_12_51_groupi_n_3495 ,csa_tree_add_12_51_groupi_n_4349);
  or csa_tree_add_12_51_groupi_g17364(csa_tree_add_12_51_groupi_n_4457 ,csa_tree_add_12_51_groupi_n_3492 ,csa_tree_add_12_51_groupi_n_4342);
  not csa_tree_add_12_51_groupi_g17365(csa_tree_add_12_51_groupi_n_4401 ,csa_tree_add_12_51_groupi_n_4402);
  not csa_tree_add_12_51_groupi_g17366(csa_tree_add_12_51_groupi_n_4397 ,csa_tree_add_12_51_groupi_n_4396);
  or csa_tree_add_12_51_groupi_g17367(csa_tree_add_12_51_groupi_n_4393 ,csa_tree_add_12_51_groupi_n_3514 ,csa_tree_add_12_51_groupi_n_4310);
  or csa_tree_add_12_51_groupi_g17368(csa_tree_add_12_51_groupi_n_4392 ,csa_tree_add_12_51_groupi_n_3231 ,csa_tree_add_12_51_groupi_n_4307);
  and csa_tree_add_12_51_groupi_g17369(csa_tree_add_12_51_groupi_n_4391 ,csa_tree_add_12_51_groupi_n_3514 ,csa_tree_add_12_51_groupi_n_4310);
  or csa_tree_add_12_51_groupi_g17370(csa_tree_add_12_51_groupi_n_4390 ,csa_tree_add_12_51_groupi_n_3512 ,csa_tree_add_12_51_groupi_n_4300);
  nor csa_tree_add_12_51_groupi_g17371(csa_tree_add_12_51_groupi_n_4389 ,csa_tree_add_12_51_groupi_n_1583 ,csa_tree_add_12_51_groupi_n_1019);
  nor csa_tree_add_12_51_groupi_g17372(csa_tree_add_12_51_groupi_n_4388 ,csa_tree_add_12_51_groupi_n_1592 ,csa_tree_add_12_51_groupi_n_1022);
  nor csa_tree_add_12_51_groupi_g17373(csa_tree_add_12_51_groupi_n_4387 ,csa_tree_add_12_51_groupi_n_1604 ,csa_tree_add_12_51_groupi_n_157);
  and csa_tree_add_12_51_groupi_g17374(csa_tree_add_12_51_groupi_n_4386 ,csa_tree_add_12_51_groupi_n_4361 ,csa_tree_add_12_51_groupi_n_4295);
  or csa_tree_add_12_51_groupi_g17375(csa_tree_add_12_51_groupi_n_4385 ,csa_tree_add_12_51_groupi_n_4270 ,csa_tree_add_12_51_groupi_n_4316);
  or csa_tree_add_12_51_groupi_g17376(csa_tree_add_12_51_groupi_n_4384 ,csa_tree_add_12_51_groupi_n_4194 ,csa_tree_add_12_51_groupi_n_4320);
  and csa_tree_add_12_51_groupi_g17377(csa_tree_add_12_51_groupi_n_4383 ,csa_tree_add_12_51_groupi_n_4201 ,csa_tree_add_12_51_groupi_n_4325);
  and csa_tree_add_12_51_groupi_g17378(csa_tree_add_12_51_groupi_n_4382 ,csa_tree_add_12_51_groupi_n_4200 ,csa_tree_add_12_51_groupi_n_4317);
  nor csa_tree_add_12_51_groupi_g17379(csa_tree_add_12_51_groupi_n_4381 ,csa_tree_add_12_51_groupi_n_1628 ,csa_tree_add_12_51_groupi_n_1019);
  nor csa_tree_add_12_51_groupi_g17380(csa_tree_add_12_51_groupi_n_4380 ,csa_tree_add_12_51_groupi_n_1640 ,csa_tree_add_12_51_groupi_n_1020);
  nor csa_tree_add_12_51_groupi_g17381(csa_tree_add_12_51_groupi_n_4379 ,csa_tree_add_12_51_groupi_n_1616 ,csa_tree_add_12_51_groupi_n_1023);
  nor csa_tree_add_12_51_groupi_g17382(csa_tree_add_12_51_groupi_n_4378 ,csa_tree_add_12_51_groupi_n_1655 ,csa_tree_add_12_51_groupi_n_831);
  nor csa_tree_add_12_51_groupi_g17383(csa_tree_add_12_51_groupi_n_4377 ,csa_tree_add_12_51_groupi_n_1622 ,csa_tree_add_12_51_groupi_n_830);
  nor csa_tree_add_12_51_groupi_g17384(csa_tree_add_12_51_groupi_n_4376 ,csa_tree_add_12_51_groupi_n_1634 ,csa_tree_add_12_51_groupi_n_1020);
  nor csa_tree_add_12_51_groupi_g17385(csa_tree_add_12_51_groupi_n_4375 ,csa_tree_add_12_51_groupi_n_1610 ,csa_tree_add_12_51_groupi_n_830);
  nor csa_tree_add_12_51_groupi_g17386(csa_tree_add_12_51_groupi_n_4374 ,csa_tree_add_12_51_groupi_n_1586 ,csa_tree_add_12_51_groupi_n_1023);
  nor csa_tree_add_12_51_groupi_g17387(csa_tree_add_12_51_groupi_n_4373 ,csa_tree_add_12_51_groupi_n_1646 ,csa_tree_add_12_51_groupi_n_1022);
  nor csa_tree_add_12_51_groupi_g17388(csa_tree_add_12_51_groupi_n_4372 ,csa_tree_add_12_51_groupi_n_1664 ,csa_tree_add_12_51_groupi_n_1977);
  nor csa_tree_add_12_51_groupi_g17389(csa_tree_add_12_51_groupi_n_4371 ,csa_tree_add_12_51_groupi_n_1679 ,csa_tree_add_12_51_groupi_n_831);
  nor csa_tree_add_12_51_groupi_g17390(csa_tree_add_12_51_groupi_n_4370 ,csa_tree_add_12_51_groupi_n_1598 ,csa_tree_add_12_51_groupi_n_157);
  xnor csa_tree_add_12_51_groupi_g17391(csa_tree_add_12_51_groupi_n_4369 ,csa_tree_add_12_51_groupi_n_4222 ,csa_tree_add_12_51_groupi_n_4232);
  xnor csa_tree_add_12_51_groupi_g17392(csa_tree_add_12_51_groupi_n_4368 ,csa_tree_add_12_51_groupi_n_4231 ,csa_tree_add_12_51_groupi_n_4226);
  xnor csa_tree_add_12_51_groupi_g17393(csa_tree_add_12_51_groupi_n_4367 ,csa_tree_add_12_51_groupi_n_4182 ,csa_tree_add_12_51_groupi_n_4230);
  xnor csa_tree_add_12_51_groupi_g17394(csa_tree_add_12_51_groupi_n_4416 ,csa_tree_add_12_51_groupi_n_4240 ,csa_tree_add_12_51_groupi_n_1930);
  xnor csa_tree_add_12_51_groupi_g17395(csa_tree_add_12_51_groupi_n_4415 ,csa_tree_add_12_51_groupi_n_4247 ,in2[5]);
  xnor csa_tree_add_12_51_groupi_g17396(csa_tree_add_12_51_groupi_n_4414 ,csa_tree_add_12_51_groupi_n_4245 ,in3[2]);
  xnor csa_tree_add_12_51_groupi_g17397(csa_tree_add_12_51_groupi_n_4413 ,csa_tree_add_12_51_groupi_n_4251 ,in4[11]);
  xnor csa_tree_add_12_51_groupi_g17398(csa_tree_add_12_51_groupi_n_4412 ,csa_tree_add_12_51_groupi_n_4250 ,in2[11]);
  xnor csa_tree_add_12_51_groupi_g17399(csa_tree_add_12_51_groupi_n_4411 ,csa_tree_add_12_51_groupi_n_4235 ,csa_tree_add_12_51_groupi_n_3562);
  xnor csa_tree_add_12_51_groupi_g17400(csa_tree_add_12_51_groupi_n_4410 ,csa_tree_add_12_51_groupi_n_4242 ,in3[8]);
  xnor csa_tree_add_12_51_groupi_g17401(csa_tree_add_12_51_groupi_n_4409 ,csa_tree_add_12_51_groupi_n_4249 ,in3[11]);
  xnor csa_tree_add_12_51_groupi_g17402(csa_tree_add_12_51_groupi_n_4408 ,csa_tree_add_12_51_groupi_n_4243 ,in2[2]);
  xnor csa_tree_add_12_51_groupi_g17403(csa_tree_add_12_51_groupi_n_4407 ,csa_tree_add_12_51_groupi_n_4252 ,in3[5]);
  xnor csa_tree_add_12_51_groupi_g17404(csa_tree_add_12_51_groupi_n_4406 ,csa_tree_add_12_51_groupi_n_4248 ,in4[2]);
  xnor csa_tree_add_12_51_groupi_g17405(csa_tree_add_12_51_groupi_n_4405 ,csa_tree_add_12_51_groupi_n_4233 ,csa_tree_add_12_51_groupi_n_3560);
  xnor csa_tree_add_12_51_groupi_g17406(csa_tree_add_12_51_groupi_n_4404 ,csa_tree_add_12_51_groupi_n_4253 ,in2[8]);
  xnor csa_tree_add_12_51_groupi_g17407(csa_tree_add_12_51_groupi_n_4403 ,csa_tree_add_12_51_groupi_n_4239 ,in4[8]);
  xnor csa_tree_add_12_51_groupi_g17408(csa_tree_add_12_51_groupi_n_4402 ,csa_tree_add_12_51_groupi_n_4281 ,csa_tree_add_12_51_groupi_n_3981);
  xnor csa_tree_add_12_51_groupi_g17409(csa_tree_add_12_51_groupi_n_4400 ,csa_tree_add_12_51_groupi_n_4234 ,csa_tree_add_12_51_groupi_n_3564);
  xnor csa_tree_add_12_51_groupi_g17410(csa_tree_add_12_51_groupi_n_4399 ,csa_tree_add_12_51_groupi_n_4236 ,csa_tree_add_12_51_groupi_n_3559);
  xnor csa_tree_add_12_51_groupi_g17411(csa_tree_add_12_51_groupi_n_4398 ,csa_tree_add_12_51_groupi_n_4238 ,csa_tree_add_12_51_groupi_n_3561);
  xnor csa_tree_add_12_51_groupi_g17412(csa_tree_add_12_51_groupi_n_4396 ,csa_tree_add_12_51_groupi_n_4246 ,in2[14]);
  xnor csa_tree_add_12_51_groupi_g17413(csa_tree_add_12_51_groupi_n_4395 ,csa_tree_add_12_51_groupi_n_4244 ,in4[14]);
  xnor csa_tree_add_12_51_groupi_g17414(csa_tree_add_12_51_groupi_n_4394 ,csa_tree_add_12_51_groupi_n_4241 ,in4[5]);
  and csa_tree_add_12_51_groupi_g17415(csa_tree_add_12_51_groupi_n_4356 ,csa_tree_add_12_51_groupi_n_4204 ,csa_tree_add_12_51_groupi_n_4205);
  and csa_tree_add_12_51_groupi_g17416(csa_tree_add_12_51_groupi_n_4355 ,csa_tree_add_12_51_groupi_n_3485 ,csa_tree_add_12_51_groupi_n_4233);
  and csa_tree_add_12_51_groupi_g17417(csa_tree_add_12_51_groupi_n_4354 ,csa_tree_add_12_51_groupi_n_2153 ,csa_tree_add_12_51_groupi_n_4228);
  and csa_tree_add_12_51_groupi_g17418(csa_tree_add_12_51_groupi_n_4353 ,csa_tree_add_12_51_groupi_n_4231 ,csa_tree_add_12_51_groupi_n_4226);
  or csa_tree_add_12_51_groupi_g17419(csa_tree_add_12_51_groupi_n_4352 ,csa_tree_add_12_51_groupi_n_4204 ,csa_tree_add_12_51_groupi_n_4205);
  or csa_tree_add_12_51_groupi_g17420(csa_tree_add_12_51_groupi_n_4351 ,csa_tree_add_12_51_groupi_n_4231 ,csa_tree_add_12_51_groupi_n_4226);
  or csa_tree_add_12_51_groupi_g17421(csa_tree_add_12_51_groupi_n_4350 ,csa_tree_add_12_51_groupi_n_4263 ,csa_tree_add_12_51_groupi_n_4237);
  and csa_tree_add_12_51_groupi_g17422(csa_tree_add_12_51_groupi_n_4349 ,csa_tree_add_12_51_groupi_n_3489 ,csa_tree_add_12_51_groupi_n_4234);
  and csa_tree_add_12_51_groupi_g17423(csa_tree_add_12_51_groupi_n_4348 ,csa_tree_add_12_51_groupi_n_3490 ,csa_tree_add_12_51_groupi_n_4236);
  or csa_tree_add_12_51_groupi_g17424(csa_tree_add_12_51_groupi_n_4347 ,csa_tree_add_12_51_groupi_n_2153 ,csa_tree_add_12_51_groupi_n_4228);
  and csa_tree_add_12_51_groupi_g17425(csa_tree_add_12_51_groupi_n_4346 ,csa_tree_add_12_51_groupi_n_3486 ,csa_tree_add_12_51_groupi_n_4235);
  and csa_tree_add_12_51_groupi_g17426(csa_tree_add_12_51_groupi_n_4345 ,csa_tree_add_12_51_groupi_n_4222 ,csa_tree_add_12_51_groupi_n_4232);
  or csa_tree_add_12_51_groupi_g17427(csa_tree_add_12_51_groupi_n_4344 ,csa_tree_add_12_51_groupi_n_3694 ,csa_tree_add_12_51_groupi_n_4187);
  or csa_tree_add_12_51_groupi_g17428(csa_tree_add_12_51_groupi_n_4343 ,csa_tree_add_12_51_groupi_n_4222 ,csa_tree_add_12_51_groupi_n_4232);
  and csa_tree_add_12_51_groupi_g17429(csa_tree_add_12_51_groupi_n_4342 ,csa_tree_add_12_51_groupi_n_3493 ,csa_tree_add_12_51_groupi_n_4238);
  or csa_tree_add_12_51_groupi_g17430(csa_tree_add_12_51_groupi_n_4341 ,csa_tree_add_12_51_groupi_n_3626 ,csa_tree_add_12_51_groupi_n_4188);
  or csa_tree_add_12_51_groupi_g17431(csa_tree_add_12_51_groupi_n_4340 ,csa_tree_add_12_51_groupi_n_3717 ,csa_tree_add_12_51_groupi_n_4191);
  or csa_tree_add_12_51_groupi_g17432(csa_tree_add_12_51_groupi_n_4339 ,csa_tree_add_12_51_groupi_n_3699 ,csa_tree_add_12_51_groupi_n_4192);
  nor csa_tree_add_12_51_groupi_g17433(csa_tree_add_12_51_groupi_n_4338 ,csa_tree_add_12_51_groupi_n_4182 ,csa_tree_add_12_51_groupi_n_4230);
  or csa_tree_add_12_51_groupi_g17434(csa_tree_add_12_51_groupi_n_4337 ,csa_tree_add_12_51_groupi_n_4181 ,csa_tree_add_12_51_groupi_n_4229);
  or csa_tree_add_12_51_groupi_g17435(csa_tree_add_12_51_groupi_n_4336 ,csa_tree_add_12_51_groupi_n_3651 ,csa_tree_add_12_51_groupi_n_4195);
  or csa_tree_add_12_51_groupi_g17436(csa_tree_add_12_51_groupi_n_4335 ,csa_tree_add_12_51_groupi_n_3719 ,csa_tree_add_12_51_groupi_n_4196);
  or csa_tree_add_12_51_groupi_g17437(csa_tree_add_12_51_groupi_n_4334 ,csa_tree_add_12_51_groupi_n_3733 ,csa_tree_add_12_51_groupi_n_4197);
  and csa_tree_add_12_51_groupi_g17438(csa_tree_add_12_51_groupi_n_4333 ,csa_tree_add_12_51_groupi_n_3823 ,csa_tree_add_12_51_groupi_n_4281);
  or csa_tree_add_12_51_groupi_g17439(csa_tree_add_12_51_groupi_n_4332 ,csa_tree_add_12_51_groupi_n_3291 ,csa_tree_add_12_51_groupi_n_4193);
  and csa_tree_add_12_51_groupi_g17440(csa_tree_add_12_51_groupi_n_4331 ,csa_tree_add_12_51_groupi_n_3517 ,csa_tree_add_12_51_groupi_n_4227);
  nor csa_tree_add_12_51_groupi_g17441(csa_tree_add_12_51_groupi_n_4330 ,csa_tree_add_12_51_groupi_n_3517 ,csa_tree_add_12_51_groupi_n_4227);
  or csa_tree_add_12_51_groupi_g17442(csa_tree_add_12_51_groupi_n_4329 ,csa_tree_add_12_51_groupi_n_3396 ,csa_tree_add_12_51_groupi_n_4198);
  or csa_tree_add_12_51_groupi_g17443(csa_tree_add_12_51_groupi_n_4328 ,csa_tree_add_12_51_groupi_n_3380 ,csa_tree_add_12_51_groupi_n_4203);
  or csa_tree_add_12_51_groupi_g17444(csa_tree_add_12_51_groupi_n_4327 ,csa_tree_add_12_51_groupi_n_3317 ,csa_tree_add_12_51_groupi_n_4190);
  or csa_tree_add_12_51_groupi_g17445(csa_tree_add_12_51_groupi_n_4326 ,csa_tree_add_12_51_groupi_n_3273 ,csa_tree_add_12_51_groupi_n_4189);
  or csa_tree_add_12_51_groupi_g17446(csa_tree_add_12_51_groupi_n_4366 ,csa_tree_add_12_51_groupi_n_3826 ,csa_tree_add_12_51_groupi_n_4264);
  or csa_tree_add_12_51_groupi_g17447(csa_tree_add_12_51_groupi_n_4365 ,csa_tree_add_12_51_groupi_n_3818 ,csa_tree_add_12_51_groupi_n_4271);
  or csa_tree_add_12_51_groupi_g17448(csa_tree_add_12_51_groupi_n_4364 ,csa_tree_add_12_51_groupi_n_3822 ,csa_tree_add_12_51_groupi_n_4269);
  or csa_tree_add_12_51_groupi_g17449(csa_tree_add_12_51_groupi_n_4363 ,csa_tree_add_12_51_groupi_n_3828 ,csa_tree_add_12_51_groupi_n_4272);
  and csa_tree_add_12_51_groupi_g17450(csa_tree_add_12_51_groupi_n_4362 ,csa_tree_add_12_51_groupi_n_2435 ,csa_tree_add_12_51_groupi_n_4273);
  or csa_tree_add_12_51_groupi_g17451(csa_tree_add_12_51_groupi_n_4361 ,csa_tree_add_12_51_groupi_n_3963 ,csa_tree_add_12_51_groupi_n_4277);
  or csa_tree_add_12_51_groupi_g17452(csa_tree_add_12_51_groupi_n_4360 ,csa_tree_add_12_51_groupi_n_3960 ,csa_tree_add_12_51_groupi_n_4279);
  or csa_tree_add_12_51_groupi_g17453(csa_tree_add_12_51_groupi_n_4359 ,csa_tree_add_12_51_groupi_n_3965 ,csa_tree_add_12_51_groupi_n_4274);
  or csa_tree_add_12_51_groupi_g17454(csa_tree_add_12_51_groupi_n_4358 ,csa_tree_add_12_51_groupi_n_3969 ,csa_tree_add_12_51_groupi_n_4276);
  or csa_tree_add_12_51_groupi_g17455(csa_tree_add_12_51_groupi_n_4357 ,csa_tree_add_12_51_groupi_n_3964 ,csa_tree_add_12_51_groupi_n_4280);
  not csa_tree_add_12_51_groupi_g17456(csa_tree_add_12_51_groupi_n_4320 ,csa_tree_add_12_51_groupi_n_4319);
  not csa_tree_add_12_51_groupi_g17457(csa_tree_add_12_51_groupi_n_4316 ,csa_tree_add_12_51_groupi_n_4315);
  or csa_tree_add_12_51_groupi_g17458(csa_tree_add_12_51_groupi_n_4298 ,csa_tree_add_12_51_groupi_n_3024 ,csa_tree_add_12_51_groupi_n_4256);
  or csa_tree_add_12_51_groupi_g17459(csa_tree_add_12_51_groupi_n_4297 ,csa_tree_add_12_51_groupi_n_3012 ,csa_tree_add_12_51_groupi_n_4257);
  nor csa_tree_add_12_51_groupi_g17460(csa_tree_add_12_51_groupi_n_4296 ,csa_tree_add_12_51_groupi_n_4221 ,csa_tree_add_12_51_groupi_n_4219);
  or csa_tree_add_12_51_groupi_g17461(csa_tree_add_12_51_groupi_n_4295 ,csa_tree_add_12_51_groupi_n_4220 ,csa_tree_add_12_51_groupi_n_8);
  or csa_tree_add_12_51_groupi_g17462(csa_tree_add_12_51_groupi_n_4294 ,csa_tree_add_12_51_groupi_n_5 ,csa_tree_add_12_51_groupi_n_4223);
  nor csa_tree_add_12_51_groupi_g17463(csa_tree_add_12_51_groupi_n_4293 ,csa_tree_add_12_51_groupi_n_4225 ,csa_tree_add_12_51_groupi_n_4224);
  or csa_tree_add_12_51_groupi_g17464(csa_tree_add_12_51_groupi_n_4292 ,csa_tree_add_12_51_groupi_n_3067 ,csa_tree_add_12_51_groupi_n_4255);
  xor csa_tree_add_12_51_groupi_g17465(csa_tree_add_12_51_groupi_n_4291 ,csa_tree_add_12_51_groupi_n_3517 ,csa_tree_add_12_51_groupi_n_4184);
  xnor csa_tree_add_12_51_groupi_g17466(csa_tree_add_12_51_groupi_n_4290 ,csa_tree_add_12_51_groupi_n_3521 ,csa_tree_add_12_51_groupi_n_4173);
  xnor csa_tree_add_12_51_groupi_g17467(csa_tree_add_12_51_groupi_n_4289 ,csa_tree_add_12_51_groupi_n_3232 ,csa_tree_add_12_51_groupi_n_4180);
  xnor csa_tree_add_12_51_groupi_g17468(csa_tree_add_12_51_groupi_n_4288 ,csa_tree_add_12_51_groupi_n_3516 ,csa_tree_add_12_51_groupi_n_4175);
  xnor csa_tree_add_12_51_groupi_g17469(csa_tree_add_12_51_groupi_n_4287 ,csa_tree_add_12_51_groupi_n_3542 ,csa_tree_add_12_51_groupi_n_4179);
  xnor csa_tree_add_12_51_groupi_g17470(csa_tree_add_12_51_groupi_n_4286 ,csa_tree_add_12_51_groupi_n_4128 ,csa_tree_add_12_51_groupi_n_4141);
  xnor csa_tree_add_12_51_groupi_g17471(csa_tree_add_12_51_groupi_n_4285 ,csa_tree_add_12_51_groupi_n_4134 ,csa_tree_add_12_51_groupi_n_4140);
  xnor csa_tree_add_12_51_groupi_g17472(csa_tree_add_12_51_groupi_n_4284 ,csa_tree_add_12_51_groupi_n_4130 ,csa_tree_add_12_51_groupi_n_4131);
  xnor csa_tree_add_12_51_groupi_g17473(csa_tree_add_12_51_groupi_n_4283 ,csa_tree_add_12_51_groupi_n_4137 ,csa_tree_add_12_51_groupi_n_4132);
  xnor csa_tree_add_12_51_groupi_g17474(csa_tree_add_12_51_groupi_n_4282 ,csa_tree_add_12_51_groupi_n_2757 ,csa_tree_add_12_51_groupi_n_4177);
  xnor csa_tree_add_12_51_groupi_g17475(csa_tree_add_12_51_groupi_n_4325 ,csa_tree_add_12_51_groupi_n_4145 ,csa_tree_add_12_51_groupi_n_3984);
  xnor csa_tree_add_12_51_groupi_g17476(csa_tree_add_12_51_groupi_n_4324 ,csa_tree_add_12_51_groupi_n_4153 ,csa_tree_add_12_51_groupi_n_2367);
  xnor csa_tree_add_12_51_groupi_g17477(csa_tree_add_12_51_groupi_n_4323 ,csa_tree_add_12_51_groupi_n_4156 ,in2[2]);
  xnor csa_tree_add_12_51_groupi_g17478(csa_tree_add_12_51_groupi_n_4322 ,csa_tree_add_12_51_groupi_n_4154 ,csa_tree_add_12_51_groupi_n_2362);
  xnor csa_tree_add_12_51_groupi_g17479(csa_tree_add_12_51_groupi_n_4321 ,csa_tree_add_12_51_groupi_n_4152 ,in2[8]);
  xnor csa_tree_add_12_51_groupi_g17480(csa_tree_add_12_51_groupi_n_4319 ,csa_tree_add_12_51_groupi_n_4144 ,csa_tree_add_12_51_groupi_n_3987);
  xnor csa_tree_add_12_51_groupi_g17481(csa_tree_add_12_51_groupi_n_4318 ,csa_tree_add_12_51_groupi_n_4160 ,in3[11]);
  xnor csa_tree_add_12_51_groupi_g17482(csa_tree_add_12_51_groupi_n_4317 ,csa_tree_add_12_51_groupi_n_4147 ,csa_tree_add_12_51_groupi_n_3983);
  xnor csa_tree_add_12_51_groupi_g17483(csa_tree_add_12_51_groupi_n_4315 ,csa_tree_add_12_51_groupi_n_4148 ,csa_tree_add_12_51_groupi_n_3986);
  xnor csa_tree_add_12_51_groupi_g17484(csa_tree_add_12_51_groupi_n_4314 ,csa_tree_add_12_51_groupi_n_4149 ,csa_tree_add_12_51_groupi_n_3985);
  xnor csa_tree_add_12_51_groupi_g17485(csa_tree_add_12_51_groupi_n_4313 ,csa_tree_add_12_51_groupi_n_4158 ,in4[2]);
  xnor csa_tree_add_12_51_groupi_g17486(csa_tree_add_12_51_groupi_n_4312 ,csa_tree_add_12_51_groupi_n_4185 ,csa_tree_add_12_51_groupi_n_3979);
  xnor csa_tree_add_12_51_groupi_g17487(csa_tree_add_12_51_groupi_n_4311 ,csa_tree_add_12_51_groupi_n_4155 ,in3[8]);
  xnor csa_tree_add_12_51_groupi_g17488(csa_tree_add_12_51_groupi_n_4310 ,csa_tree_add_12_51_groupi_n_4150 ,csa_tree_add_12_51_groupi_n_3980);
  xnor csa_tree_add_12_51_groupi_g17489(csa_tree_add_12_51_groupi_n_4309 ,csa_tree_add_12_51_groupi_n_4157 ,in3[2]);
  xnor csa_tree_add_12_51_groupi_g17490(csa_tree_add_12_51_groupi_n_4308 ,csa_tree_add_12_51_groupi_n_4159 ,in2[11]);
  xnor csa_tree_add_12_51_groupi_g17491(csa_tree_add_12_51_groupi_n_4307 ,csa_tree_add_12_51_groupi_n_4146 ,csa_tree_add_12_51_groupi_n_3976);
  xnor csa_tree_add_12_51_groupi_g17492(csa_tree_add_12_51_groupi_n_4306 ,csa_tree_add_12_51_groupi_n_4161 ,in4[11]);
  xnor csa_tree_add_12_51_groupi_g17493(csa_tree_add_12_51_groupi_n_4305 ,csa_tree_add_12_51_groupi_n_4164 ,in2[5]);
  xnor csa_tree_add_12_51_groupi_g17494(csa_tree_add_12_51_groupi_n_4304 ,csa_tree_add_12_51_groupi_n_4163 ,in4[5]);
  xnor csa_tree_add_12_51_groupi_g17495(csa_tree_add_12_51_groupi_n_4303 ,csa_tree_add_12_51_groupi_n_4165 ,in4[8]);
  xnor csa_tree_add_12_51_groupi_g17496(csa_tree_add_12_51_groupi_n_4302 ,csa_tree_add_12_51_groupi_n_4162 ,in4[14]);
  xnor csa_tree_add_12_51_groupi_g17497(csa_tree_add_12_51_groupi_n_4301 ,csa_tree_add_12_51_groupi_n_4151 ,in3[14]);
  xnor csa_tree_add_12_51_groupi_g17498(csa_tree_add_12_51_groupi_n_4300 ,csa_tree_add_12_51_groupi_n_4143 ,csa_tree_add_12_51_groupi_n_3978);
  xnor csa_tree_add_12_51_groupi_g17499(csa_tree_add_12_51_groupi_n_4299 ,csa_tree_add_12_51_groupi_n_4183 ,csa_tree_add_12_51_groupi_n_2562);
  and csa_tree_add_12_51_groupi_g17500(csa_tree_add_12_51_groupi_n_4280 ,csa_tree_add_12_51_groupi_n_3961 ,csa_tree_add_12_51_groupi_n_4147);
  and csa_tree_add_12_51_groupi_g17501(csa_tree_add_12_51_groupi_n_4279 ,csa_tree_add_12_51_groupi_n_3959 ,csa_tree_add_12_51_groupi_n_4144);
  or csa_tree_add_12_51_groupi_g17502(csa_tree_add_12_51_groupi_n_4278 ,csa_tree_add_12_51_groupi_n_4138 ,csa_tree_add_12_51_groupi_n_4142);
  and csa_tree_add_12_51_groupi_g17503(csa_tree_add_12_51_groupi_n_4277 ,csa_tree_add_12_51_groupi_n_3958 ,csa_tree_add_12_51_groupi_n_4145);
  and csa_tree_add_12_51_groupi_g17504(csa_tree_add_12_51_groupi_n_4276 ,csa_tree_add_12_51_groupi_n_3867 ,csa_tree_add_12_51_groupi_n_4149);
  and csa_tree_add_12_51_groupi_g17505(csa_tree_add_12_51_groupi_n_4275 ,csa_tree_add_12_51_groupi_n_4138 ,csa_tree_add_12_51_groupi_n_4142);
  and csa_tree_add_12_51_groupi_g17506(csa_tree_add_12_51_groupi_n_4274 ,csa_tree_add_12_51_groupi_n_3968 ,csa_tree_add_12_51_groupi_n_4148);
  or csa_tree_add_12_51_groupi_g17507(csa_tree_add_12_51_groupi_n_4273 ,csa_tree_add_12_51_groupi_n_2424 ,csa_tree_add_12_51_groupi_n_4183);
  and csa_tree_add_12_51_groupi_g17508(csa_tree_add_12_51_groupi_n_4272 ,csa_tree_add_12_51_groupi_n_3829 ,csa_tree_add_12_51_groupi_n_4146);
  and csa_tree_add_12_51_groupi_g17509(csa_tree_add_12_51_groupi_n_4271 ,csa_tree_add_12_51_groupi_n_3819 ,csa_tree_add_12_51_groupi_n_4185);
  nor csa_tree_add_12_51_groupi_g17510(csa_tree_add_12_51_groupi_n_4270 ,csa_tree_add_12_51_groupi_n_4128 ,csa_tree_add_12_51_groupi_n_4141);
  and csa_tree_add_12_51_groupi_g17511(csa_tree_add_12_51_groupi_n_4269 ,csa_tree_add_12_51_groupi_n_3824 ,csa_tree_add_12_51_groupi_n_4143);
  or csa_tree_add_12_51_groupi_g17512(csa_tree_add_12_51_groupi_n_4268 ,csa_tree_add_12_51_groupi_n_3521 ,csa_tree_add_12_51_groupi_n_4173);
  and csa_tree_add_12_51_groupi_g17513(csa_tree_add_12_51_groupi_n_4267 ,csa_tree_add_12_51_groupi_n_3232 ,csa_tree_add_12_51_groupi_n_4180);
  or csa_tree_add_12_51_groupi_g17514(csa_tree_add_12_51_groupi_n_4266 ,csa_tree_add_12_51_groupi_n_3232 ,csa_tree_add_12_51_groupi_n_4180);
  and csa_tree_add_12_51_groupi_g17515(csa_tree_add_12_51_groupi_n_4265 ,csa_tree_add_12_51_groupi_n_3521 ,csa_tree_add_12_51_groupi_n_4173);
  and csa_tree_add_12_51_groupi_g17516(csa_tree_add_12_51_groupi_n_4264 ,csa_tree_add_12_51_groupi_n_3827 ,csa_tree_add_12_51_groupi_n_4150);
  nor csa_tree_add_12_51_groupi_g17517(csa_tree_add_12_51_groupi_n_4263 ,csa_tree_add_12_51_groupi_n_3542 ,csa_tree_add_12_51_groupi_n_4178);
  or csa_tree_add_12_51_groupi_g17518(csa_tree_add_12_51_groupi_n_4262 ,csa_tree_add_12_51_groupi_n_3541 ,csa_tree_add_12_51_groupi_n_4179);
  nor csa_tree_add_12_51_groupi_g17519(csa_tree_add_12_51_groupi_n_4261 ,csa_tree_add_12_51_groupi_n_3515 ,csa_tree_add_12_51_groupi_n_4175);
  or csa_tree_add_12_51_groupi_g17520(csa_tree_add_12_51_groupi_n_4260 ,csa_tree_add_12_51_groupi_n_3516 ,csa_tree_add_12_51_groupi_n_4174);
  nor csa_tree_add_12_51_groupi_g17521(csa_tree_add_12_51_groupi_n_4259 ,csa_tree_add_12_51_groupi_n_2757 ,csa_tree_add_12_51_groupi_n_4176);
  or csa_tree_add_12_51_groupi_g17522(csa_tree_add_12_51_groupi_n_4258 ,csa_tree_add_12_51_groupi_n_2756 ,csa_tree_add_12_51_groupi_n_4177);
  nor csa_tree_add_12_51_groupi_g17523(csa_tree_add_12_51_groupi_n_4257 ,csa_tree_add_12_51_groupi_n_1590 ,csa_tree_add_12_51_groupi_n_995);
  nor csa_tree_add_12_51_groupi_g17524(csa_tree_add_12_51_groupi_n_4256 ,csa_tree_add_12_51_groupi_n_1602 ,csa_tree_add_12_51_groupi_n_998);
  nor csa_tree_add_12_51_groupi_g17525(csa_tree_add_12_51_groupi_n_4255 ,csa_tree_add_12_51_groupi_n_1581 ,csa_tree_add_12_51_groupi_n_155);
  or csa_tree_add_12_51_groupi_g17526(csa_tree_add_12_51_groupi_n_4254 ,csa_tree_add_12_51_groupi_n_4127 ,csa_tree_add_12_51_groupi_n_7);
  nor csa_tree_add_12_51_groupi_g17527(csa_tree_add_12_51_groupi_n_4253 ,csa_tree_add_12_51_groupi_n_3887 ,csa_tree_add_12_51_groupi_n_4125);
  nor csa_tree_add_12_51_groupi_g17528(csa_tree_add_12_51_groupi_n_4252 ,csa_tree_add_12_51_groupi_n_4073 ,csa_tree_add_12_51_groupi_n_4172);
  nor csa_tree_add_12_51_groupi_g17529(csa_tree_add_12_51_groupi_n_4251 ,csa_tree_add_12_51_groupi_n_3833 ,csa_tree_add_12_51_groupi_n_4121);
  nor csa_tree_add_12_51_groupi_g17530(csa_tree_add_12_51_groupi_n_4250 ,csa_tree_add_12_51_groupi_n_3840 ,csa_tree_add_12_51_groupi_n_4120);
  nor csa_tree_add_12_51_groupi_g17531(csa_tree_add_12_51_groupi_n_4249 ,csa_tree_add_12_51_groupi_n_3860 ,csa_tree_add_12_51_groupi_n_4123);
  nor csa_tree_add_12_51_groupi_g17532(csa_tree_add_12_51_groupi_n_4248 ,csa_tree_add_12_51_groupi_n_3478 ,csa_tree_add_12_51_groupi_n_4119);
  nor csa_tree_add_12_51_groupi_g17533(csa_tree_add_12_51_groupi_n_4247 ,csa_tree_add_12_51_groupi_n_4082 ,csa_tree_add_12_51_groupi_n_4168);
  nor csa_tree_add_12_51_groupi_g17534(csa_tree_add_12_51_groupi_n_4246 ,csa_tree_add_12_51_groupi_n_3924 ,csa_tree_add_12_51_groupi_n_4171);
  nor csa_tree_add_12_51_groupi_g17535(csa_tree_add_12_51_groupi_n_4245 ,csa_tree_add_12_51_groupi_n_3474 ,csa_tree_add_12_51_groupi_n_4118);
  nor csa_tree_add_12_51_groupi_g17536(csa_tree_add_12_51_groupi_n_4244 ,csa_tree_add_12_51_groupi_n_3903 ,csa_tree_add_12_51_groupi_n_4170);
  nor csa_tree_add_12_51_groupi_g17537(csa_tree_add_12_51_groupi_n_4243 ,csa_tree_add_12_51_groupi_n_3477 ,csa_tree_add_12_51_groupi_n_4117);
  nor csa_tree_add_12_51_groupi_g17538(csa_tree_add_12_51_groupi_n_4242 ,csa_tree_add_12_51_groupi_n_3871 ,csa_tree_add_12_51_groupi_n_4124);
  nor csa_tree_add_12_51_groupi_g17539(csa_tree_add_12_51_groupi_n_4241 ,csa_tree_add_12_51_groupi_n_4081 ,csa_tree_add_12_51_groupi_n_4169);
  nor csa_tree_add_12_51_groupi_g17540(csa_tree_add_12_51_groupi_n_4240 ,csa_tree_add_12_51_groupi_n_3970 ,csa_tree_add_12_51_groupi_n_4122);
  nor csa_tree_add_12_51_groupi_g17541(csa_tree_add_12_51_groupi_n_4239 ,csa_tree_add_12_51_groupi_n_3923 ,csa_tree_add_12_51_groupi_n_4166);
  or csa_tree_add_12_51_groupi_g17542(csa_tree_add_12_51_groupi_n_4281 ,csa_tree_add_12_51_groupi_n_3825 ,csa_tree_add_12_51_groupi_n_4167);
  not csa_tree_add_12_51_groupi_g17543(csa_tree_add_12_51_groupi_n_4229 ,csa_tree_add_12_51_groupi_n_4230);
  not csa_tree_add_12_51_groupi_g17544(csa_tree_add_12_51_groupi_n_4225 ,csa_tree_add_12_51_groupi_n_5);
  not csa_tree_add_12_51_groupi_g17545(csa_tree_add_12_51_groupi_n_4224 ,csa_tree_add_12_51_groupi_n_4223);
  not csa_tree_add_12_51_groupi_g17546(csa_tree_add_12_51_groupi_n_4221 ,csa_tree_add_12_51_groupi_n_4220);
  not csa_tree_add_12_51_groupi_g17547(csa_tree_add_12_51_groupi_n_4219 ,csa_tree_add_12_51_groupi_n_8);
  not csa_tree_add_12_51_groupi_g17548(csa_tree_add_12_51_groupi_n_4217 ,csa_tree_add_12_51_groupi_n_4218);
  not csa_tree_add_12_51_groupi_g17549(csa_tree_add_12_51_groupi_n_4215 ,csa_tree_add_12_51_groupi_n_4216);
  not csa_tree_add_12_51_groupi_g17550(csa_tree_add_12_51_groupi_n_4213 ,csa_tree_add_12_51_groupi_n_4214);
  not csa_tree_add_12_51_groupi_g17551(csa_tree_add_12_51_groupi_n_4210 ,csa_tree_add_12_51_groupi_n_4211);
  not csa_tree_add_12_51_groupi_g17552(csa_tree_add_12_51_groupi_n_4208 ,csa_tree_add_12_51_groupi_n_4209);
  not csa_tree_add_12_51_groupi_g17553(csa_tree_add_12_51_groupi_n_4206 ,csa_tree_add_12_51_groupi_n_4207);
  nor csa_tree_add_12_51_groupi_g17554(csa_tree_add_12_51_groupi_n_4203 ,csa_tree_add_12_51_groupi_n_1608 ,csa_tree_add_12_51_groupi_n_995);
  and csa_tree_add_12_51_groupi_g17555(csa_tree_add_12_51_groupi_n_4202 ,csa_tree_add_12_51_groupi_n_4137 ,csa_tree_add_12_51_groupi_n_4132);
  or csa_tree_add_12_51_groupi_g17556(csa_tree_add_12_51_groupi_n_4201 ,csa_tree_add_12_51_groupi_n_4137 ,csa_tree_add_12_51_groupi_n_4132);
  or csa_tree_add_12_51_groupi_g17557(csa_tree_add_12_51_groupi_n_4200 ,csa_tree_add_12_51_groupi_n_4130 ,csa_tree_add_12_51_groupi_n_4131);
  and csa_tree_add_12_51_groupi_g17558(csa_tree_add_12_51_groupi_n_4199 ,csa_tree_add_12_51_groupi_n_4130 ,csa_tree_add_12_51_groupi_n_4131);
  nor csa_tree_add_12_51_groupi_g17559(csa_tree_add_12_51_groupi_n_4198 ,csa_tree_add_12_51_groupi_n_1596 ,csa_tree_add_12_51_groupi_n_996);
  nor csa_tree_add_12_51_groupi_g17560(csa_tree_add_12_51_groupi_n_4197 ,csa_tree_add_12_51_groupi_n_1620 ,csa_tree_add_12_51_groupi_n_999);
  nor csa_tree_add_12_51_groupi_g17561(csa_tree_add_12_51_groupi_n_4196 ,csa_tree_add_12_51_groupi_n_1689 ,csa_tree_add_12_51_groupi_n_936);
  nor csa_tree_add_12_51_groupi_g17562(csa_tree_add_12_51_groupi_n_4195 ,csa_tree_add_12_51_groupi_n_1614 ,csa_tree_add_12_51_groupi_n_935);
  nor csa_tree_add_12_51_groupi_g17563(csa_tree_add_12_51_groupi_n_4194 ,csa_tree_add_12_51_groupi_n_4134 ,csa_tree_add_12_51_groupi_n_4140);
  nor csa_tree_add_12_51_groupi_g17564(csa_tree_add_12_51_groupi_n_4193 ,csa_tree_add_12_51_groupi_n_1650 ,csa_tree_add_12_51_groupi_n_996);
  nor csa_tree_add_12_51_groupi_g17565(csa_tree_add_12_51_groupi_n_4192 ,csa_tree_add_12_51_groupi_n_1644 ,csa_tree_add_12_51_groupi_n_935);
  nor csa_tree_add_12_51_groupi_g17566(csa_tree_add_12_51_groupi_n_4191 ,csa_tree_add_12_51_groupi_n_1638 ,csa_tree_add_12_51_groupi_n_999);
  nor csa_tree_add_12_51_groupi_g17567(csa_tree_add_12_51_groupi_n_4190 ,csa_tree_add_12_51_groupi_n_1632 ,csa_tree_add_12_51_groupi_n_998);
  nor csa_tree_add_12_51_groupi_g17568(csa_tree_add_12_51_groupi_n_4189 ,csa_tree_add_12_51_groupi_n_1671 ,csa_tree_add_12_51_groupi_n_1968);
  nor csa_tree_add_12_51_groupi_g17569(csa_tree_add_12_51_groupi_n_4188 ,csa_tree_add_12_51_groupi_n_1659 ,csa_tree_add_12_51_groupi_n_936);
  nor csa_tree_add_12_51_groupi_g17570(csa_tree_add_12_51_groupi_n_4187 ,csa_tree_add_12_51_groupi_n_1626 ,csa_tree_add_12_51_groupi_n_155);
  or csa_tree_add_12_51_groupi_g17571(csa_tree_add_12_51_groupi_n_4186 ,csa_tree_add_12_51_groupi_n_4133 ,csa_tree_add_12_51_groupi_n_4139);
  xnor csa_tree_add_12_51_groupi_g17572(csa_tree_add_12_51_groupi_n_4238 ,csa_tree_add_12_51_groupi_n_4049 ,in3[14]);
  xnor csa_tree_add_12_51_groupi_g17573(csa_tree_add_12_51_groupi_n_4237 ,csa_tree_add_12_51_groupi_n_3557 ,csa_tree_add_12_51_groupi_n_3995);
  xnor csa_tree_add_12_51_groupi_g17574(csa_tree_add_12_51_groupi_n_4236 ,csa_tree_add_12_51_groupi_n_118 ,csa_tree_add_12_51_groupi_n_3999);
  xnor csa_tree_add_12_51_groupi_g17575(csa_tree_add_12_51_groupi_n_4235 ,csa_tree_add_12_51_groupi_n_4051 ,in2[11]);
  xnor csa_tree_add_12_51_groupi_g17576(csa_tree_add_12_51_groupi_n_4234 ,csa_tree_add_12_51_groupi_n_4000 ,in2[5]);
  xnor csa_tree_add_12_51_groupi_g17577(csa_tree_add_12_51_groupi_n_4233 ,csa_tree_add_12_51_groupi_n_4045 ,in4[8]);
  xnor csa_tree_add_12_51_groupi_g17578(csa_tree_add_12_51_groupi_n_4232 ,csa_tree_add_12_51_groupi_n_4050 ,in3[11]);
  xnor csa_tree_add_12_51_groupi_g17579(csa_tree_add_12_51_groupi_n_4231 ,csa_tree_add_12_51_groupi_n_4046 ,in2[8]);
  xnor csa_tree_add_12_51_groupi_g17580(csa_tree_add_12_51_groupi_n_4230 ,csa_tree_add_12_51_groupi_n_3554 ,csa_tree_add_12_51_groupi_n_3975);
  xnor csa_tree_add_12_51_groupi_g17581(csa_tree_add_12_51_groupi_n_4228 ,csa_tree_add_12_51_groupi_n_4116 ,csa_tree_add_12_51_groupi_n_3977);
  xnor csa_tree_add_12_51_groupi_g17582(csa_tree_add_12_51_groupi_n_4227 ,csa_tree_add_12_51_groupi_n_3558 ,csa_tree_add_12_51_groupi_n_3982);
  xnor csa_tree_add_12_51_groupi_g17583(csa_tree_add_12_51_groupi_n_4226 ,csa_tree_add_12_51_groupi_n_4048 ,in3[8]);
  xnor csa_tree_add_12_51_groupi_g17585(csa_tree_add_12_51_groupi_n_4223 ,csa_tree_add_12_51_groupi_n_1959 ,csa_tree_add_12_51_groupi_n_3974);
  xnor csa_tree_add_12_51_groupi_g17586(csa_tree_add_12_51_groupi_n_4222 ,csa_tree_add_12_51_groupi_n_4052 ,in4[11]);
  xnor csa_tree_add_12_51_groupi_g17587(csa_tree_add_12_51_groupi_n_4220 ,csa_tree_add_12_51_groupi_n_1936 ,csa_tree_add_12_51_groupi_n_3997);
  xnor csa_tree_add_12_51_groupi_g17589(csa_tree_add_12_51_groupi_n_4218 ,csa_tree_add_12_51_groupi_n_3551 ,csa_tree_add_12_51_groupi_n_3988);
  xnor csa_tree_add_12_51_groupi_g17590(csa_tree_add_12_51_groupi_n_4216 ,csa_tree_add_12_51_groupi_n_3255 ,csa_tree_add_12_51_groupi_n_3989);
  xnor csa_tree_add_12_51_groupi_g17591(csa_tree_add_12_51_groupi_n_4214 ,csa_tree_add_12_51_groupi_n_3552 ,csa_tree_add_12_51_groupi_n_3991);
  xnor csa_tree_add_12_51_groupi_g17592(csa_tree_add_12_51_groupi_n_4212 ,csa_tree_add_12_51_groupi_n_3254 ,csa_tree_add_12_51_groupi_n_3990);
  xnor csa_tree_add_12_51_groupi_g17593(csa_tree_add_12_51_groupi_n_4211 ,csa_tree_add_12_51_groupi_n_3253 ,csa_tree_add_12_51_groupi_n_3992);
  xnor csa_tree_add_12_51_groupi_g17594(csa_tree_add_12_51_groupi_n_4209 ,csa_tree_add_12_51_groupi_n_3553 ,csa_tree_add_12_51_groupi_n_3993);
  xnor csa_tree_add_12_51_groupi_g17595(csa_tree_add_12_51_groupi_n_4207 ,csa_tree_add_12_51_groupi_n_3556 ,csa_tree_add_12_51_groupi_n_3994);
  xnor csa_tree_add_12_51_groupi_g17596(csa_tree_add_12_51_groupi_n_4205 ,csa_tree_add_12_51_groupi_n_4044 ,in2[14]);
  xnor csa_tree_add_12_51_groupi_g17597(csa_tree_add_12_51_groupi_n_4204 ,csa_tree_add_12_51_groupi_n_4047 ,in4[14]);
  not csa_tree_add_12_51_groupi_g17598(csa_tree_add_12_51_groupi_n_4181 ,csa_tree_add_12_51_groupi_n_4182);
  not csa_tree_add_12_51_groupi_g17599(csa_tree_add_12_51_groupi_n_4179 ,csa_tree_add_12_51_groupi_n_4178);
  not csa_tree_add_12_51_groupi_g17600(csa_tree_add_12_51_groupi_n_4176 ,csa_tree_add_12_51_groupi_n_4177);
  not csa_tree_add_12_51_groupi_g17601(csa_tree_add_12_51_groupi_n_4175 ,csa_tree_add_12_51_groupi_n_4174);
  or csa_tree_add_12_51_groupi_g17602(csa_tree_add_12_51_groupi_n_4172 ,csa_tree_add_12_51_groupi_n_3358 ,csa_tree_add_12_51_groupi_n_4003);
  or csa_tree_add_12_51_groupi_g17603(csa_tree_add_12_51_groupi_n_4171 ,csa_tree_add_12_51_groupi_n_3751 ,csa_tree_add_12_51_groupi_n_4002);
  or csa_tree_add_12_51_groupi_g17604(csa_tree_add_12_51_groupi_n_4170 ,csa_tree_add_12_51_groupi_n_3760 ,csa_tree_add_12_51_groupi_n_4006);
  or csa_tree_add_12_51_groupi_g17605(csa_tree_add_12_51_groupi_n_4169 ,csa_tree_add_12_51_groupi_n_3270 ,csa_tree_add_12_51_groupi_n_4008);
  or csa_tree_add_12_51_groupi_g17606(csa_tree_add_12_51_groupi_n_4168 ,csa_tree_add_12_51_groupi_n_3275 ,csa_tree_add_12_51_groupi_n_4031);
  and csa_tree_add_12_51_groupi_g17607(csa_tree_add_12_51_groupi_n_4167 ,csa_tree_add_12_51_groupi_n_3820 ,csa_tree_add_12_51_groupi_n_4116);
  or csa_tree_add_12_51_groupi_g17608(csa_tree_add_12_51_groupi_n_4166 ,csa_tree_add_12_51_groupi_n_3755 ,csa_tree_add_12_51_groupi_n_4004);
  nor csa_tree_add_12_51_groupi_g17609(csa_tree_add_12_51_groupi_n_4165 ,csa_tree_add_12_51_groupi_n_3942 ,csa_tree_add_12_51_groupi_n_4021);
  nor csa_tree_add_12_51_groupi_g17610(csa_tree_add_12_51_groupi_n_4164 ,csa_tree_add_12_51_groupi_n_4088 ,csa_tree_add_12_51_groupi_n_4029);
  nor csa_tree_add_12_51_groupi_g17611(csa_tree_add_12_51_groupi_n_4163 ,csa_tree_add_12_51_groupi_n_4090 ,csa_tree_add_12_51_groupi_n_4030);
  nor csa_tree_add_12_51_groupi_g17612(csa_tree_add_12_51_groupi_n_4162 ,csa_tree_add_12_51_groupi_n_3940 ,csa_tree_add_12_51_groupi_n_4024);
  nor csa_tree_add_12_51_groupi_g17613(csa_tree_add_12_51_groupi_n_4161 ,csa_tree_add_12_51_groupi_n_3929 ,csa_tree_add_12_51_groupi_n_4018);
  nor csa_tree_add_12_51_groupi_g17614(csa_tree_add_12_51_groupi_n_4160 ,csa_tree_add_12_51_groupi_n_3933 ,csa_tree_add_12_51_groupi_n_4017);
  nor csa_tree_add_12_51_groupi_g17615(csa_tree_add_12_51_groupi_n_4159 ,csa_tree_add_12_51_groupi_n_4089 ,csa_tree_add_12_51_groupi_n_4028);
  nor csa_tree_add_12_51_groupi_g17616(csa_tree_add_12_51_groupi_n_4158 ,csa_tree_add_12_51_groupi_n_3483 ,csa_tree_add_12_51_groupi_n_4014);
  nor csa_tree_add_12_51_groupi_g17617(csa_tree_add_12_51_groupi_n_4157 ,csa_tree_add_12_51_groupi_n_3482 ,csa_tree_add_12_51_groupi_n_4015);
  nor csa_tree_add_12_51_groupi_g17618(csa_tree_add_12_51_groupi_n_4156 ,csa_tree_add_12_51_groupi_n_3481 ,csa_tree_add_12_51_groupi_n_4013);
  nor csa_tree_add_12_51_groupi_g17619(csa_tree_add_12_51_groupi_n_4155 ,csa_tree_add_12_51_groupi_n_3938 ,csa_tree_add_12_51_groupi_n_4019);
  nor csa_tree_add_12_51_groupi_g17620(csa_tree_add_12_51_groupi_n_4154 ,csa_tree_add_12_51_groupi_n_3944 ,csa_tree_add_12_51_groupi_n_4016);
  nor csa_tree_add_12_51_groupi_g17621(csa_tree_add_12_51_groupi_n_4153 ,csa_tree_add_12_51_groupi_n_3945 ,csa_tree_add_12_51_groupi_n_4023);
  nor csa_tree_add_12_51_groupi_g17622(csa_tree_add_12_51_groupi_n_4152 ,csa_tree_add_12_51_groupi_n_3946 ,csa_tree_add_12_51_groupi_n_4020);
  nor csa_tree_add_12_51_groupi_g17623(csa_tree_add_12_51_groupi_n_4151 ,csa_tree_add_12_51_groupi_n_3935 ,csa_tree_add_12_51_groupi_n_4022);
  or csa_tree_add_12_51_groupi_g17624(csa_tree_add_12_51_groupi_n_4185 ,csa_tree_add_12_51_groupi_n_3817 ,csa_tree_add_12_51_groupi_n_4093);
  and csa_tree_add_12_51_groupi_g17625(csa_tree_add_12_51_groupi_n_4184 ,csa_tree_add_12_51_groupi_n_3883 ,csa_tree_add_12_51_groupi_n_4099);
  and csa_tree_add_12_51_groupi_g17626(csa_tree_add_12_51_groupi_n_4183 ,csa_tree_add_12_51_groupi_n_2420 ,csa_tree_add_12_51_groupi_n_4112);
  or csa_tree_add_12_51_groupi_g17627(csa_tree_add_12_51_groupi_n_4182 ,csa_tree_add_12_51_groupi_n_3962 ,csa_tree_add_12_51_groupi_n_4113);
  or csa_tree_add_12_51_groupi_g17628(csa_tree_add_12_51_groupi_n_4180 ,csa_tree_add_12_51_groupi_n_3805 ,csa_tree_add_12_51_groupi_n_4087);
  or csa_tree_add_12_51_groupi_g17629(csa_tree_add_12_51_groupi_n_4178 ,csa_tree_add_12_51_groupi_n_3436 ,csa_tree_add_12_51_groupi_n_4102);
  or csa_tree_add_12_51_groupi_g17630(csa_tree_add_12_51_groupi_n_4177 ,csa_tree_add_12_51_groupi_n_3814 ,csa_tree_add_12_51_groupi_n_4092);
  or csa_tree_add_12_51_groupi_g17631(csa_tree_add_12_51_groupi_n_4174 ,csa_tree_add_12_51_groupi_n_3807 ,csa_tree_add_12_51_groupi_n_4115);
  or csa_tree_add_12_51_groupi_g17632(csa_tree_add_12_51_groupi_n_4173 ,csa_tree_add_12_51_groupi_n_3810 ,csa_tree_add_12_51_groupi_n_4091);
  not csa_tree_add_12_51_groupi_g17633(csa_tree_add_12_51_groupi_n_4141 ,csa_tree_add_12_51_groupi_n_7);
  not csa_tree_add_12_51_groupi_g17634(csa_tree_add_12_51_groupi_n_4140 ,csa_tree_add_12_51_groupi_n_4139);
  not csa_tree_add_12_51_groupi_g17635(csa_tree_add_12_51_groupi_n_4134 ,csa_tree_add_12_51_groupi_n_4133);
  not csa_tree_add_12_51_groupi_g17637(csa_tree_add_12_51_groupi_n_4128 ,csa_tree_add_12_51_groupi_n_4127);
  or csa_tree_add_12_51_groupi_g17638(csa_tree_add_12_51_groupi_n_4125 ,csa_tree_add_12_51_groupi_n_3744 ,csa_tree_add_12_51_groupi_n_4005);
  or csa_tree_add_12_51_groupi_g17639(csa_tree_add_12_51_groupi_n_4124 ,csa_tree_add_12_51_groupi_n_3743 ,csa_tree_add_12_51_groupi_n_4001);
  or csa_tree_add_12_51_groupi_g17640(csa_tree_add_12_51_groupi_n_4123 ,csa_tree_add_12_51_groupi_n_3753 ,csa_tree_add_12_51_groupi_n_4009);
  or csa_tree_add_12_51_groupi_g17641(csa_tree_add_12_51_groupi_n_4122 ,csa_tree_add_12_51_groupi_n_3758 ,csa_tree_add_12_51_groupi_n_4007);
  or csa_tree_add_12_51_groupi_g17642(csa_tree_add_12_51_groupi_n_4121 ,csa_tree_add_12_51_groupi_n_3741 ,csa_tree_add_12_51_groupi_n_4033);
  or csa_tree_add_12_51_groupi_g17643(csa_tree_add_12_51_groupi_n_4120 ,csa_tree_add_12_51_groupi_n_3745 ,csa_tree_add_12_51_groupi_n_4032);
  or csa_tree_add_12_51_groupi_g17644(csa_tree_add_12_51_groupi_n_4119 ,csa_tree_add_12_51_groupi_n_3119 ,csa_tree_add_12_51_groupi_n_4011);
  or csa_tree_add_12_51_groupi_g17645(csa_tree_add_12_51_groupi_n_4118 ,csa_tree_add_12_51_groupi_n_3159 ,csa_tree_add_12_51_groupi_n_4010);
  or csa_tree_add_12_51_groupi_g17646(csa_tree_add_12_51_groupi_n_4117 ,csa_tree_add_12_51_groupi_n_3059 ,csa_tree_add_12_51_groupi_n_4012);
  or csa_tree_add_12_51_groupi_g17647(csa_tree_add_12_51_groupi_n_4150 ,csa_tree_add_12_51_groupi_n_3791 ,csa_tree_add_12_51_groupi_n_4025);
  xnor csa_tree_add_12_51_groupi_g17648(csa_tree_add_12_51_groupi_n_4149 ,csa_tree_add_12_51_groupi_n_3768 ,in2[2]);
  xnor csa_tree_add_12_51_groupi_g17649(csa_tree_add_12_51_groupi_n_4148 ,csa_tree_add_12_51_groupi_n_3779 ,in4[11]);
  xnor csa_tree_add_12_51_groupi_g17650(csa_tree_add_12_51_groupi_n_4147 ,csa_tree_add_12_51_groupi_n_3777 ,in3[14]);
  or csa_tree_add_12_51_groupi_g17651(csa_tree_add_12_51_groupi_n_4146 ,csa_tree_add_12_51_groupi_n_3790 ,csa_tree_add_12_51_groupi_n_4026);
  xnor csa_tree_add_12_51_groupi_g17652(csa_tree_add_12_51_groupi_n_4145 ,csa_tree_add_12_51_groupi_n_3772 ,in2[5]);
  xnor csa_tree_add_12_51_groupi_g17653(csa_tree_add_12_51_groupi_n_4144 ,csa_tree_add_12_51_groupi_n_3769 ,in2[8]);
  or csa_tree_add_12_51_groupi_g17654(csa_tree_add_12_51_groupi_n_4143 ,csa_tree_add_12_51_groupi_n_3794 ,csa_tree_add_12_51_groupi_n_4027);
  xnor csa_tree_add_12_51_groupi_g17655(csa_tree_add_12_51_groupi_n_4142 ,csa_tree_add_12_51_groupi_n_3767 ,in3[2]);
  xnor csa_tree_add_12_51_groupi_g17657(csa_tree_add_12_51_groupi_n_4139 ,csa_tree_add_12_51_groupi_n_98 ,csa_tree_add_12_51_groupi_n_3778);
  xnor csa_tree_add_12_51_groupi_g17658(csa_tree_add_12_51_groupi_n_4138 ,csa_tree_add_12_51_groupi_n_3766 ,in4[2]);
  xnor csa_tree_add_12_51_groupi_g17659(csa_tree_add_12_51_groupi_n_4137 ,csa_tree_add_12_51_groupi_n_3780 ,in4[5]);
  xnor csa_tree_add_12_51_groupi_g17660(csa_tree_add_12_51_groupi_n_4136 ,csa_tree_add_12_51_groupi_n_3550 ,csa_tree_add_12_51_groupi_n_3566);
  xnor csa_tree_add_12_51_groupi_g17661(csa_tree_add_12_51_groupi_n_4135 ,csa_tree_add_12_51_groupi_n_3765 ,csa_tree_add_12_51_groupi_n_3563);
  xnor csa_tree_add_12_51_groupi_g17662(csa_tree_add_12_51_groupi_n_4133 ,csa_tree_add_12_51_groupi_n_1938 ,csa_tree_add_12_51_groupi_n_3773);
  xnor csa_tree_add_12_51_groupi_g17663(csa_tree_add_12_51_groupi_n_4132 ,csa_tree_add_12_51_groupi_n_3775 ,in3[5]);
  xnor csa_tree_add_12_51_groupi_g17664(csa_tree_add_12_51_groupi_n_4131 ,csa_tree_add_12_51_groupi_n_3771 ,in2[14]);
  xnor csa_tree_add_12_51_groupi_g17665(csa_tree_add_12_51_groupi_n_4130 ,csa_tree_add_12_51_groupi_n_3776 ,in4[14]);
  xnor csa_tree_add_12_51_groupi_g17666(csa_tree_add_12_51_groupi_n_4129 ,csa_tree_add_12_51_groupi_n_2755 ,csa_tree_add_12_51_groupi_n_3565);
  xnor csa_tree_add_12_51_groupi_g17667(csa_tree_add_12_51_groupi_n_4127 ,csa_tree_add_12_51_groupi_n_1920 ,csa_tree_add_12_51_groupi_n_3770);
  xnor csa_tree_add_12_51_groupi_g17668(csa_tree_add_12_51_groupi_n_4126 ,csa_tree_add_12_51_groupi_n_3971 ,csa_tree_add_12_51_groupi_n_2559);
  and csa_tree_add_12_51_groupi_g17669(csa_tree_add_12_51_groupi_n_4115 ,csa_tree_add_12_51_groupi_n_3551 ,csa_tree_add_12_51_groupi_n_3808);
  or csa_tree_add_12_51_groupi_g17670(csa_tree_add_12_51_groupi_n_4114 ,csa_tree_add_12_51_groupi_n_3003 ,csa_tree_add_12_51_groupi_n_3707);
  and csa_tree_add_12_51_groupi_g17671(csa_tree_add_12_51_groupi_n_4113 ,csa_tree_add_12_51_groupi_n_3557 ,csa_tree_add_12_51_groupi_n_3967);
  or csa_tree_add_12_51_groupi_g17672(csa_tree_add_12_51_groupi_n_4112 ,csa_tree_add_12_51_groupi_n_2425 ,csa_tree_add_12_51_groupi_n_3971);
  or csa_tree_add_12_51_groupi_g17673(csa_tree_add_12_51_groupi_n_4111 ,csa_tree_add_12_51_groupi_n_3028 ,csa_tree_add_12_51_groupi_n_3590);
  or csa_tree_add_12_51_groupi_g17674(csa_tree_add_12_51_groupi_n_4110 ,csa_tree_add_12_51_groupi_n_3111 ,csa_tree_add_12_51_groupi_n_3662);
  or csa_tree_add_12_51_groupi_g17675(csa_tree_add_12_51_groupi_n_4109 ,csa_tree_add_12_51_groupi_n_3075 ,csa_tree_add_12_51_groupi_n_3604);
  or csa_tree_add_12_51_groupi_g17676(csa_tree_add_12_51_groupi_n_4108 ,csa_tree_add_12_51_groupi_n_3031 ,csa_tree_add_12_51_groupi_n_3638);
  or csa_tree_add_12_51_groupi_g17677(csa_tree_add_12_51_groupi_n_4107 ,csa_tree_add_12_51_groupi_n_3071 ,csa_tree_add_12_51_groupi_n_3678);
  or csa_tree_add_12_51_groupi_g17678(csa_tree_add_12_51_groupi_n_4106 ,csa_tree_add_12_51_groupi_n_3086 ,csa_tree_add_12_51_groupi_n_3686);
  or csa_tree_add_12_51_groupi_g17679(csa_tree_add_12_51_groupi_n_4105 ,csa_tree_add_12_51_groupi_n_3054 ,csa_tree_add_12_51_groupi_n_3650);
  or csa_tree_add_12_51_groupi_g17680(csa_tree_add_12_51_groupi_n_4104 ,csa_tree_add_12_51_groupi_n_3107 ,csa_tree_add_12_51_groupi_n_3652);
  or csa_tree_add_12_51_groupi_g17681(csa_tree_add_12_51_groupi_n_4103 ,csa_tree_add_12_51_groupi_n_3044 ,csa_tree_add_12_51_groupi_n_3670);
  nor csa_tree_add_12_51_groupi_g17682(csa_tree_add_12_51_groupi_n_4102 ,csa_tree_add_12_51_groupi_n_3437 ,csa_tree_add_12_51_groupi_n_3765);
  or csa_tree_add_12_51_groupi_g17683(csa_tree_add_12_51_groupi_n_4101 ,csa_tree_add_12_51_groupi_n_3343 ,csa_tree_add_12_51_groupi_n_3629);
  or csa_tree_add_12_51_groupi_g17684(csa_tree_add_12_51_groupi_n_4100 ,csa_tree_add_12_51_groupi_n_3356 ,csa_tree_add_12_51_groupi_n_3605);
  or csa_tree_add_12_51_groupi_g17685(csa_tree_add_12_51_groupi_n_4099 ,csa_tree_add_12_51_groupi_n_3555 ,csa_tree_add_12_51_groupi_n_3884);
  or csa_tree_add_12_51_groupi_g17686(csa_tree_add_12_51_groupi_n_4098 ,csa_tree_add_12_51_groupi_n_3297 ,csa_tree_add_12_51_groupi_n_3689);
  or csa_tree_add_12_51_groupi_g17687(csa_tree_add_12_51_groupi_n_4097 ,csa_tree_add_12_51_groupi_n_3279 ,csa_tree_add_12_51_groupi_n_3632);
  or csa_tree_add_12_51_groupi_g17688(csa_tree_add_12_51_groupi_n_4096 ,csa_tree_add_12_51_groupi_n_3281 ,csa_tree_add_12_51_groupi_n_3620);
  or csa_tree_add_12_51_groupi_g17689(csa_tree_add_12_51_groupi_n_4095 ,csa_tree_add_12_51_groupi_n_3271 ,csa_tree_add_12_51_groupi_n_3732);
  or csa_tree_add_12_51_groupi_g17690(csa_tree_add_12_51_groupi_n_4094 ,csa_tree_add_12_51_groupi_n_3352 ,csa_tree_add_12_51_groupi_n_3606);
  and csa_tree_add_12_51_groupi_g17691(csa_tree_add_12_51_groupi_n_4093 ,csa_tree_add_12_51_groupi_n_3558 ,csa_tree_add_12_51_groupi_n_3816);
  and csa_tree_add_12_51_groupi_g17692(csa_tree_add_12_51_groupi_n_4092 ,csa_tree_add_12_51_groupi_n_3556 ,csa_tree_add_12_51_groupi_n_3815);
  and csa_tree_add_12_51_groupi_g17693(csa_tree_add_12_51_groupi_n_4091 ,csa_tree_add_12_51_groupi_n_3253 ,csa_tree_add_12_51_groupi_n_3809);
  or csa_tree_add_12_51_groupi_g17694(csa_tree_add_12_51_groupi_n_4090 ,csa_tree_add_12_51_groupi_n_3176 ,csa_tree_add_12_51_groupi_n_3782);
  or csa_tree_add_12_51_groupi_g17695(csa_tree_add_12_51_groupi_n_4089 ,csa_tree_add_12_51_groupi_n_3192 ,csa_tree_add_12_51_groupi_n_3781);
  or csa_tree_add_12_51_groupi_g17696(csa_tree_add_12_51_groupi_n_4088 ,csa_tree_add_12_51_groupi_n_3185 ,csa_tree_add_12_51_groupi_n_3762);
  and csa_tree_add_12_51_groupi_g17697(csa_tree_add_12_51_groupi_n_4087 ,csa_tree_add_12_51_groupi_n_3553 ,csa_tree_add_12_51_groupi_n_3806);
  or csa_tree_add_12_51_groupi_g17698(csa_tree_add_12_51_groupi_n_4086 ,csa_tree_add_12_51_groupi_n_3178 ,csa_tree_add_12_51_groupi_n_3722);
  or csa_tree_add_12_51_groupi_g17699(csa_tree_add_12_51_groupi_n_4085 ,csa_tree_add_12_51_groupi_n_3179 ,csa_tree_add_12_51_groupi_n_3734);
  or csa_tree_add_12_51_groupi_g17700(csa_tree_add_12_51_groupi_n_4084 ,csa_tree_add_12_51_groupi_n_3174 ,csa_tree_add_12_51_groupi_n_3598);
  or csa_tree_add_12_51_groupi_g17701(csa_tree_add_12_51_groupi_n_4083 ,csa_tree_add_12_51_groupi_n_3201 ,csa_tree_add_12_51_groupi_n_3700);
  or csa_tree_add_12_51_groupi_g17702(csa_tree_add_12_51_groupi_n_4082 ,csa_tree_add_12_51_groupi_n_3043 ,csa_tree_add_12_51_groupi_n_3742);
  or csa_tree_add_12_51_groupi_g17703(csa_tree_add_12_51_groupi_n_4081 ,csa_tree_add_12_51_groupi_n_2998 ,csa_tree_add_12_51_groupi_n_3756);
  or csa_tree_add_12_51_groupi_g17704(csa_tree_add_12_51_groupi_n_4080 ,csa_tree_add_12_51_groupi_n_3184 ,csa_tree_add_12_51_groupi_n_3594);
  or csa_tree_add_12_51_groupi_g17705(csa_tree_add_12_51_groupi_n_4079 ,csa_tree_add_12_51_groupi_n_3183 ,csa_tree_add_12_51_groupi_n_3639);
  or csa_tree_add_12_51_groupi_g17706(csa_tree_add_12_51_groupi_n_4078 ,csa_tree_add_12_51_groupi_n_3191 ,csa_tree_add_12_51_groupi_n_3637);
  or csa_tree_add_12_51_groupi_g17707(csa_tree_add_12_51_groupi_n_4077 ,csa_tree_add_12_51_groupi_n_3189 ,csa_tree_add_12_51_groupi_n_3593);
  or csa_tree_add_12_51_groupi_g17708(csa_tree_add_12_51_groupi_n_4076 ,csa_tree_add_12_51_groupi_n_3203 ,csa_tree_add_12_51_groupi_n_3631);
  or csa_tree_add_12_51_groupi_g17709(csa_tree_add_12_51_groupi_n_4075 ,csa_tree_add_12_51_groupi_n_3175 ,csa_tree_add_12_51_groupi_n_3655);
  or csa_tree_add_12_51_groupi_g17710(csa_tree_add_12_51_groupi_n_4074 ,csa_tree_add_12_51_groupi_n_3181 ,csa_tree_add_12_51_groupi_n_3710);
  or csa_tree_add_12_51_groupi_g17711(csa_tree_add_12_51_groupi_n_4073 ,csa_tree_add_12_51_groupi_n_3045 ,csa_tree_add_12_51_groupi_n_3740);
  or csa_tree_add_12_51_groupi_g17712(csa_tree_add_12_51_groupi_n_4072 ,csa_tree_add_12_51_groupi_n_3199 ,csa_tree_add_12_51_groupi_n_3654);
  or csa_tree_add_12_51_groupi_g17713(csa_tree_add_12_51_groupi_n_4071 ,csa_tree_add_12_51_groupi_n_3076 ,csa_tree_add_12_51_groupi_n_3619);
  or csa_tree_add_12_51_groupi_g17714(csa_tree_add_12_51_groupi_n_4070 ,csa_tree_add_12_51_groupi_n_3081 ,csa_tree_add_12_51_groupi_n_3705);
  or csa_tree_add_12_51_groupi_g17715(csa_tree_add_12_51_groupi_n_4069 ,csa_tree_add_12_51_groupi_n_3078 ,csa_tree_add_12_51_groupi_n_3634);
  or csa_tree_add_12_51_groupi_g17716(csa_tree_add_12_51_groupi_n_4068 ,csa_tree_add_12_51_groupi_n_2983 ,csa_tree_add_12_51_groupi_n_3642);
  or csa_tree_add_12_51_groupi_g17717(csa_tree_add_12_51_groupi_n_4067 ,csa_tree_add_12_51_groupi_n_3007 ,csa_tree_add_12_51_groupi_n_3611);
  or csa_tree_add_12_51_groupi_g17718(csa_tree_add_12_51_groupi_n_4066 ,csa_tree_add_12_51_groupi_n_3165 ,csa_tree_add_12_51_groupi_n_3588);
  or csa_tree_add_12_51_groupi_g17719(csa_tree_add_12_51_groupi_n_4065 ,csa_tree_add_12_51_groupi_n_3048 ,csa_tree_add_12_51_groupi_n_3625);
  or csa_tree_add_12_51_groupi_g17720(csa_tree_add_12_51_groupi_n_4064 ,csa_tree_add_12_51_groupi_n_2995 ,csa_tree_add_12_51_groupi_n_3712);
  or csa_tree_add_12_51_groupi_g17721(csa_tree_add_12_51_groupi_n_4063 ,csa_tree_add_12_51_groupi_n_3011 ,csa_tree_add_12_51_groupi_n_3669);
  or csa_tree_add_12_51_groupi_g17722(csa_tree_add_12_51_groupi_n_4062 ,csa_tree_add_12_51_groupi_n_3056 ,csa_tree_add_12_51_groupi_n_3667);
  or csa_tree_add_12_51_groupi_g17723(csa_tree_add_12_51_groupi_n_4061 ,csa_tree_add_12_51_groupi_n_2992 ,csa_tree_add_12_51_groupi_n_3683);
  or csa_tree_add_12_51_groupi_g17724(csa_tree_add_12_51_groupi_n_4060 ,csa_tree_add_12_51_groupi_n_3033 ,csa_tree_add_12_51_groupi_n_3682);
  or csa_tree_add_12_51_groupi_g17725(csa_tree_add_12_51_groupi_n_4059 ,csa_tree_add_12_51_groupi_n_2994 ,csa_tree_add_12_51_groupi_n_3616);
  or csa_tree_add_12_51_groupi_g17726(csa_tree_add_12_51_groupi_n_4058 ,csa_tree_add_12_51_groupi_n_3055 ,csa_tree_add_12_51_groupi_n_3718);
  or csa_tree_add_12_51_groupi_g17727(csa_tree_add_12_51_groupi_n_4057 ,csa_tree_add_12_51_groupi_n_3069 ,csa_tree_add_12_51_groupi_n_3706);
  or csa_tree_add_12_51_groupi_g17728(csa_tree_add_12_51_groupi_n_4056 ,csa_tree_add_12_51_groupi_n_3060 ,csa_tree_add_12_51_groupi_n_3724);
  or csa_tree_add_12_51_groupi_g17729(csa_tree_add_12_51_groupi_n_4055 ,csa_tree_add_12_51_groupi_n_3127 ,csa_tree_add_12_51_groupi_n_3610);
  or csa_tree_add_12_51_groupi_g17730(csa_tree_add_12_51_groupi_n_4054 ,csa_tree_add_12_51_groupi_n_3021 ,csa_tree_add_12_51_groupi_n_3687);
  or csa_tree_add_12_51_groupi_g17731(csa_tree_add_12_51_groupi_n_4053 ,csa_tree_add_12_51_groupi_n_3133 ,csa_tree_add_12_51_groupi_n_3729);
  nor csa_tree_add_12_51_groupi_g17732(csa_tree_add_12_51_groupi_n_4052 ,csa_tree_add_12_51_groupi_n_3226 ,csa_tree_add_12_51_groupi_n_3948);
  nor csa_tree_add_12_51_groupi_g17733(csa_tree_add_12_51_groupi_n_4051 ,csa_tree_add_12_51_groupi_n_3227 ,csa_tree_add_12_51_groupi_n_3949);
  nor csa_tree_add_12_51_groupi_g17734(csa_tree_add_12_51_groupi_n_4050 ,csa_tree_add_12_51_groupi_n_3221 ,csa_tree_add_12_51_groupi_n_3951);
  nor csa_tree_add_12_51_groupi_g17735(csa_tree_add_12_51_groupi_n_4049 ,csa_tree_add_12_51_groupi_n_3222 ,csa_tree_add_12_51_groupi_n_3950);
  nor csa_tree_add_12_51_groupi_g17736(csa_tree_add_12_51_groupi_n_4048 ,csa_tree_add_12_51_groupi_n_3225 ,csa_tree_add_12_51_groupi_n_3952);
  nor csa_tree_add_12_51_groupi_g17737(csa_tree_add_12_51_groupi_n_4047 ,csa_tree_add_12_51_groupi_n_3084 ,csa_tree_add_12_51_groupi_n_3956);
  nor csa_tree_add_12_51_groupi_g17738(csa_tree_add_12_51_groupi_n_4046 ,csa_tree_add_12_51_groupi_n_2963 ,csa_tree_add_12_51_groupi_n_3954);
  nor csa_tree_add_12_51_groupi_g17739(csa_tree_add_12_51_groupi_n_4045 ,csa_tree_add_12_51_groupi_n_2962 ,csa_tree_add_12_51_groupi_n_3953);
  nor csa_tree_add_12_51_groupi_g17740(csa_tree_add_12_51_groupi_n_4044 ,csa_tree_add_12_51_groupi_n_3220 ,csa_tree_add_12_51_groupi_n_3955);
  or csa_tree_add_12_51_groupi_g17741(csa_tree_add_12_51_groupi_n_4116 ,csa_tree_add_12_51_groupi_n_3494 ,csa_tree_add_12_51_groupi_n_3966);
  or csa_tree_add_12_51_groupi_g17742(csa_tree_add_12_51_groupi_n_4043 ,csa_tree_add_12_51_groupi_n_3160 ,csa_tree_add_12_51_groupi_n_3623);
  or csa_tree_add_12_51_groupi_g17743(csa_tree_add_12_51_groupi_n_4042 ,csa_tree_add_12_51_groupi_n_3157 ,csa_tree_add_12_51_groupi_n_3622);
  or csa_tree_add_12_51_groupi_g17744(csa_tree_add_12_51_groupi_n_4041 ,csa_tree_add_12_51_groupi_n_3019 ,csa_tree_add_12_51_groupi_n_3621);
  or csa_tree_add_12_51_groupi_g17745(csa_tree_add_12_51_groupi_n_4040 ,csa_tree_add_12_51_groupi_n_3062 ,csa_tree_add_12_51_groupi_n_3673);
  or csa_tree_add_12_51_groupi_g17746(csa_tree_add_12_51_groupi_n_4039 ,csa_tree_add_12_51_groupi_n_3036 ,csa_tree_add_12_51_groupi_n_3609);
  or csa_tree_add_12_51_groupi_g17747(csa_tree_add_12_51_groupi_n_4038 ,csa_tree_add_12_51_groupi_n_3017 ,csa_tree_add_12_51_groupi_n_3645);
  or csa_tree_add_12_51_groupi_g17748(csa_tree_add_12_51_groupi_n_4037 ,csa_tree_add_12_51_groupi_n_3008 ,csa_tree_add_12_51_groupi_n_3692);
  or csa_tree_add_12_51_groupi_g17749(csa_tree_add_12_51_groupi_n_4036 ,csa_tree_add_12_51_groupi_n_3135 ,csa_tree_add_12_51_groupi_n_3721);
  or csa_tree_add_12_51_groupi_g17750(csa_tree_add_12_51_groupi_n_4035 ,csa_tree_add_12_51_groupi_n_3092 ,csa_tree_add_12_51_groupi_n_3589);
  or csa_tree_add_12_51_groupi_g17751(csa_tree_add_12_51_groupi_n_4034 ,csa_tree_add_12_51_groupi_n_3085 ,csa_tree_add_12_51_groupi_n_3646);
  nor csa_tree_add_12_51_groupi_g17752(csa_tree_add_12_51_groupi_n_4033 ,csa_tree_add_12_51_groupi_n_64 ,csa_tree_add_12_51_groupi_n_818);
  nor csa_tree_add_12_51_groupi_g17753(csa_tree_add_12_51_groupi_n_4032 ,csa_tree_add_12_51_groupi_n_31 ,csa_tree_add_12_51_groupi_n_821);
  nor csa_tree_add_12_51_groupi_g17754(csa_tree_add_12_51_groupi_n_4031 ,csa_tree_add_12_51_groupi_n_25 ,csa_tree_add_12_51_groupi_n_173);
  or csa_tree_add_12_51_groupi_g17755(csa_tree_add_12_51_groupi_n_4030 ,csa_tree_add_12_51_groupi_n_3290 ,csa_tree_add_12_51_groupi_n_3567);
  or csa_tree_add_12_51_groupi_g17756(csa_tree_add_12_51_groupi_n_4029 ,csa_tree_add_12_51_groupi_n_3308 ,csa_tree_add_12_51_groupi_n_3571);
  or csa_tree_add_12_51_groupi_g17757(csa_tree_add_12_51_groupi_n_4028 ,csa_tree_add_12_51_groupi_n_3265 ,csa_tree_add_12_51_groupi_n_3568);
  and csa_tree_add_12_51_groupi_g17758(csa_tree_add_12_51_groupi_n_4027 ,csa_tree_add_12_51_groupi_n_3552 ,csa_tree_add_12_51_groupi_n_3793);
  and csa_tree_add_12_51_groupi_g17759(csa_tree_add_12_51_groupi_n_4026 ,csa_tree_add_12_51_groupi_n_3254 ,csa_tree_add_12_51_groupi_n_3792);
  and csa_tree_add_12_51_groupi_g17760(csa_tree_add_12_51_groupi_n_4025 ,csa_tree_add_12_51_groupi_n_3255 ,csa_tree_add_12_51_groupi_n_3789);
  or csa_tree_add_12_51_groupi_g17761(csa_tree_add_12_51_groupi_n_4024 ,csa_tree_add_12_51_groupi_n_3813 ,csa_tree_add_12_51_groupi_n_3578);
  or csa_tree_add_12_51_groupi_g17762(csa_tree_add_12_51_groupi_n_4023 ,csa_tree_add_12_51_groupi_n_3788 ,csa_tree_add_12_51_groupi_n_3576);
  or csa_tree_add_12_51_groupi_g17763(csa_tree_add_12_51_groupi_n_4022 ,csa_tree_add_12_51_groupi_n_3787 ,csa_tree_add_12_51_groupi_n_3569);
  or csa_tree_add_12_51_groupi_g17764(csa_tree_add_12_51_groupi_n_4021 ,csa_tree_add_12_51_groupi_n_3784 ,csa_tree_add_12_51_groupi_n_3573);
  or csa_tree_add_12_51_groupi_g17765(csa_tree_add_12_51_groupi_n_4020 ,csa_tree_add_12_51_groupi_n_3957 ,csa_tree_add_12_51_groupi_n_3575);
  or csa_tree_add_12_51_groupi_g17766(csa_tree_add_12_51_groupi_n_4019 ,csa_tree_add_12_51_groupi_n_3795 ,csa_tree_add_12_51_groupi_n_3570);
  or csa_tree_add_12_51_groupi_g17767(csa_tree_add_12_51_groupi_n_4018 ,csa_tree_add_12_51_groupi_n_3811 ,csa_tree_add_12_51_groupi_n_3577);
  or csa_tree_add_12_51_groupi_g17768(csa_tree_add_12_51_groupi_n_4017 ,csa_tree_add_12_51_groupi_n_3812 ,csa_tree_add_12_51_groupi_n_3572);
  or csa_tree_add_12_51_groupi_g17769(csa_tree_add_12_51_groupi_n_4016 ,csa_tree_add_12_51_groupi_n_3783 ,csa_tree_add_12_51_groupi_n_3574);
  or csa_tree_add_12_51_groupi_g17770(csa_tree_add_12_51_groupi_n_4015 ,csa_tree_add_12_51_groupi_n_3131 ,csa_tree_add_12_51_groupi_n_3581);
  or csa_tree_add_12_51_groupi_g17771(csa_tree_add_12_51_groupi_n_4014 ,csa_tree_add_12_51_groupi_n_3015 ,csa_tree_add_12_51_groupi_n_3579);
  or csa_tree_add_12_51_groupi_g17772(csa_tree_add_12_51_groupi_n_4013 ,csa_tree_add_12_51_groupi_n_2986 ,csa_tree_add_12_51_groupi_n_3580);
  nor csa_tree_add_12_51_groupi_g17773(csa_tree_add_12_51_groupi_n_4012 ,csa_tree_add_12_51_groupi_n_43 ,csa_tree_add_12_51_groupi_n_818);
  nor csa_tree_add_12_51_groupi_g17774(csa_tree_add_12_51_groupi_n_4011 ,csa_tree_add_12_51_groupi_n_37 ,csa_tree_add_12_51_groupi_n_819);
  nor csa_tree_add_12_51_groupi_g17775(csa_tree_add_12_51_groupi_n_4010 ,csa_tree_add_12_51_groupi_n_28 ,csa_tree_add_12_51_groupi_n_822);
  nor csa_tree_add_12_51_groupi_g17776(csa_tree_add_12_51_groupi_n_4009 ,csa_tree_add_12_51_groupi_n_58 ,csa_tree_add_12_51_groupi_n_849);
  nor csa_tree_add_12_51_groupi_g17777(csa_tree_add_12_51_groupi_n_4008 ,csa_tree_add_12_51_groupi_n_55 ,csa_tree_add_12_51_groupi_n_848);
  nor csa_tree_add_12_51_groupi_g17778(csa_tree_add_12_51_groupi_n_4007 ,csa_tree_add_12_51_groupi_n_22 ,csa_tree_add_12_51_groupi_n_819);
  nor csa_tree_add_12_51_groupi_g17779(csa_tree_add_12_51_groupi_n_4006 ,csa_tree_add_12_51_groupi_n_46 ,csa_tree_add_12_51_groupi_n_848);
  nor csa_tree_add_12_51_groupi_g17780(csa_tree_add_12_51_groupi_n_4005 ,csa_tree_add_12_51_groupi_n_49 ,csa_tree_add_12_51_groupi_n_822);
  nor csa_tree_add_12_51_groupi_g17781(csa_tree_add_12_51_groupi_n_4004 ,csa_tree_add_12_51_groupi_n_40 ,csa_tree_add_12_51_groupi_n_821);
  nor csa_tree_add_12_51_groupi_g17782(csa_tree_add_12_51_groupi_n_4003 ,csa_tree_add_12_51_groupi_n_61 ,csa_tree_add_12_51_groupi_n_1992);
  nor csa_tree_add_12_51_groupi_g17783(csa_tree_add_12_51_groupi_n_4002 ,csa_tree_add_12_51_groupi_n_52 ,csa_tree_add_12_51_groupi_n_849);
  nor csa_tree_add_12_51_groupi_g17784(csa_tree_add_12_51_groupi_n_4001 ,csa_tree_add_12_51_groupi_n_34 ,csa_tree_add_12_51_groupi_n_173);
  nor csa_tree_add_12_51_groupi_g17785(csa_tree_add_12_51_groupi_n_4000 ,csa_tree_add_12_51_groupi_n_3217 ,csa_tree_add_12_51_groupi_n_3804);
  or csa_tree_add_12_51_groupi_g17786(csa_tree_add_12_51_groupi_n_3999 ,csa_tree_add_12_51_groupi_n_3187 ,csa_tree_add_12_51_groupi_n_3660);
  or csa_tree_add_12_51_groupi_g17787(csa_tree_add_12_51_groupi_n_3998 ,csa_tree_add_12_51_groupi_n_3198 ,csa_tree_add_12_51_groupi_n_3786);
  or csa_tree_add_12_51_groupi_g17788(csa_tree_add_12_51_groupi_n_3997 ,csa_tree_add_12_51_groupi_n_3409 ,csa_tree_add_12_51_groupi_n_3796);
  or csa_tree_add_12_51_groupi_g17789(csa_tree_add_12_51_groupi_n_3996 ,csa_tree_add_12_51_groupi_n_3419 ,csa_tree_add_12_51_groupi_n_3797);
  xnor csa_tree_add_12_51_groupi_g17790(csa_tree_add_12_51_groupi_n_3995 ,csa_tree_add_12_51_groupi_n_3527 ,csa_tree_add_12_51_groupi_n_3544);
  xnor csa_tree_add_12_51_groupi_g17791(csa_tree_add_12_51_groupi_n_3994 ,csa_tree_add_12_51_groupi_n_3536 ,csa_tree_add_12_51_groupi_n_3238);
  xnor csa_tree_add_12_51_groupi_g17792(csa_tree_add_12_51_groupi_n_3993 ,csa_tree_add_12_51_groupi_n_3547 ,csa_tree_add_12_51_groupi_n_3236);
  xnor csa_tree_add_12_51_groupi_g17793(csa_tree_add_12_51_groupi_n_3992 ,csa_tree_add_12_51_groupi_n_3524 ,csa_tree_add_12_51_groupi_n_3240);
  xnor csa_tree_add_12_51_groupi_g17794(csa_tree_add_12_51_groupi_n_3991 ,csa_tree_add_12_51_groupi_n_2959 ,csa_tree_add_12_51_groupi_n_3520);
  xnor csa_tree_add_12_51_groupi_g17795(csa_tree_add_12_51_groupi_n_3990 ,csa_tree_add_12_51_groupi_n_2955 ,csa_tree_add_12_51_groupi_n_3518);
  xnor csa_tree_add_12_51_groupi_g17796(csa_tree_add_12_51_groupi_n_3989 ,csa_tree_add_12_51_groupi_n_2951 ,csa_tree_add_12_51_groupi_n_3539);
  xnor csa_tree_add_12_51_groupi_g17797(csa_tree_add_12_51_groupi_n_3988 ,csa_tree_add_12_51_groupi_n_3234 ,csa_tree_add_12_51_groupi_n_3510);
  xnor csa_tree_add_12_51_groupi_g17798(csa_tree_add_12_51_groupi_n_3987 ,csa_tree_add_12_51_groupi_n_3241 ,in2[8]);
  xnor csa_tree_add_12_51_groupi_g17799(csa_tree_add_12_51_groupi_n_3986 ,csa_tree_add_12_51_groupi_n_3243 ,in3[11]);
  xnor csa_tree_add_12_51_groupi_g17800(csa_tree_add_12_51_groupi_n_3985 ,csa_tree_add_12_51_groupi_n_3242 ,in2[2]);
  xnor csa_tree_add_12_51_groupi_g17801(csa_tree_add_12_51_groupi_n_3984 ,csa_tree_add_12_51_groupi_n_3244 ,in3[5]);
  xnor csa_tree_add_12_51_groupi_g17802(csa_tree_add_12_51_groupi_n_3983 ,csa_tree_add_12_51_groupi_n_3245 ,in4[14]);
  xnor csa_tree_add_12_51_groupi_g17806(csa_tree_add_12_51_groupi_n_3982 ,csa_tree_add_12_51_groupi_n_3252 ,csa_tree_add_12_51_groupi_n_3246);
  xnor csa_tree_add_12_51_groupi_g17807(csa_tree_add_12_51_groupi_n_3981 ,csa_tree_add_12_51_groupi_n_3549 ,csa_tree_add_12_51_groupi_n_3251);
  xnor csa_tree_add_12_51_groupi_g17808(csa_tree_add_12_51_groupi_n_3980 ,csa_tree_add_12_51_groupi_n_3540 ,csa_tree_add_12_51_groupi_n_3545);
  xnor csa_tree_add_12_51_groupi_g17809(csa_tree_add_12_51_groupi_n_3979 ,csa_tree_add_12_51_groupi_n_3525 ,csa_tree_add_12_51_groupi_n_3250);
  xnor csa_tree_add_12_51_groupi_g17810(csa_tree_add_12_51_groupi_n_3978 ,csa_tree_add_12_51_groupi_n_3537 ,csa_tree_add_12_51_groupi_n_3249);
  xnor csa_tree_add_12_51_groupi_g17811(csa_tree_add_12_51_groupi_n_3977 ,csa_tree_add_12_51_groupi_n_3522 ,csa_tree_add_12_51_groupi_n_3248);
  xnor csa_tree_add_12_51_groupi_g17812(csa_tree_add_12_51_groupi_n_3976 ,csa_tree_add_12_51_groupi_n_3528 ,csa_tree_add_12_51_groupi_n_3548);
  xnor csa_tree_add_12_51_groupi_g17813(csa_tree_add_12_51_groupi_n_3975 ,csa_tree_add_12_51_groupi_n_3534 ,csa_tree_add_12_51_groupi_n_3532);
  or csa_tree_add_12_51_groupi_g17814(csa_tree_add_12_51_groupi_n_3974 ,csa_tree_add_12_51_groupi_n_3186 ,csa_tree_add_12_51_groupi_n_3785);
  not csa_tree_add_12_51_groupi_g17815(csa_tree_add_12_51_groupi_n_3973 ,csa_tree_add_12_51_groupi_n_3972);
  or csa_tree_add_12_51_groupi_g17816(csa_tree_add_12_51_groupi_n_3970 ,csa_tree_add_12_51_groupi_n_3005 ,csa_tree_add_12_51_groupi_n_3305);
  and csa_tree_add_12_51_groupi_g17817(csa_tree_add_12_51_groupi_n_3969 ,in2[2] ,csa_tree_add_12_51_groupi_n_3242);
  or csa_tree_add_12_51_groupi_g17818(csa_tree_add_12_51_groupi_n_3968 ,in3[11] ,csa_tree_add_12_51_groupi_n_3243);
  or csa_tree_add_12_51_groupi_g17819(csa_tree_add_12_51_groupi_n_3967 ,csa_tree_add_12_51_groupi_n_3526 ,csa_tree_add_12_51_groupi_n_3544);
  and csa_tree_add_12_51_groupi_g17820(csa_tree_add_12_51_groupi_n_3966 ,csa_tree_add_12_51_groupi_n_3488 ,csa_tree_add_12_51_groupi_n_3550);
  and csa_tree_add_12_51_groupi_g17821(csa_tree_add_12_51_groupi_n_3965 ,in3[11] ,csa_tree_add_12_51_groupi_n_3243);
  and csa_tree_add_12_51_groupi_g17822(csa_tree_add_12_51_groupi_n_3964 ,in4[14] ,csa_tree_add_12_51_groupi_n_3245);
  and csa_tree_add_12_51_groupi_g17823(csa_tree_add_12_51_groupi_n_3963 ,in3[5] ,csa_tree_add_12_51_groupi_n_3244);
  nor csa_tree_add_12_51_groupi_g17824(csa_tree_add_12_51_groupi_n_3962 ,csa_tree_add_12_51_groupi_n_3527 ,csa_tree_add_12_51_groupi_n_3543);
  or csa_tree_add_12_51_groupi_g17825(csa_tree_add_12_51_groupi_n_3961 ,in4[14] ,csa_tree_add_12_51_groupi_n_3245);
  and csa_tree_add_12_51_groupi_g17826(csa_tree_add_12_51_groupi_n_3960 ,in2[8] ,csa_tree_add_12_51_groupi_n_3241);
  or csa_tree_add_12_51_groupi_g17827(csa_tree_add_12_51_groupi_n_3959 ,in2[8] ,csa_tree_add_12_51_groupi_n_3241);
  or csa_tree_add_12_51_groupi_g17828(csa_tree_add_12_51_groupi_n_3958 ,in3[5] ,csa_tree_add_12_51_groupi_n_3244);
  nor csa_tree_add_12_51_groupi_g17829(csa_tree_add_12_51_groupi_n_3957 ,csa_tree_add_12_51_groupi_n_1503 ,csa_tree_add_12_51_groupi_n_133);
  or csa_tree_add_12_51_groupi_g17830(csa_tree_add_12_51_groupi_n_3956 ,csa_tree_add_12_51_groupi_n_3213 ,csa_tree_add_12_51_groupi_n_3414);
  or csa_tree_add_12_51_groupi_g17831(csa_tree_add_12_51_groupi_n_3955 ,csa_tree_add_12_51_groupi_n_3209 ,csa_tree_add_12_51_groupi_n_3421);
  or csa_tree_add_12_51_groupi_g17832(csa_tree_add_12_51_groupi_n_3954 ,csa_tree_add_12_51_groupi_n_3214 ,csa_tree_add_12_51_groupi_n_3423);
  or csa_tree_add_12_51_groupi_g17833(csa_tree_add_12_51_groupi_n_3953 ,csa_tree_add_12_51_groupi_n_3210 ,csa_tree_add_12_51_groupi_n_3422);
  or csa_tree_add_12_51_groupi_g17834(csa_tree_add_12_51_groupi_n_3952 ,csa_tree_add_12_51_groupi_n_3215 ,csa_tree_add_12_51_groupi_n_3406);
  or csa_tree_add_12_51_groupi_g17835(csa_tree_add_12_51_groupi_n_3951 ,csa_tree_add_12_51_groupi_n_3218 ,csa_tree_add_12_51_groupi_n_3407);
  or csa_tree_add_12_51_groupi_g17836(csa_tree_add_12_51_groupi_n_3950 ,csa_tree_add_12_51_groupi_n_3211 ,csa_tree_add_12_51_groupi_n_3404);
  or csa_tree_add_12_51_groupi_g17837(csa_tree_add_12_51_groupi_n_3949 ,csa_tree_add_12_51_groupi_n_3207 ,csa_tree_add_12_51_groupi_n_3401);
  or csa_tree_add_12_51_groupi_g17838(csa_tree_add_12_51_groupi_n_3948 ,csa_tree_add_12_51_groupi_n_3216 ,csa_tree_add_12_51_groupi_n_3400);
  or csa_tree_add_12_51_groupi_g17839(csa_tree_add_12_51_groupi_n_3947 ,csa_tree_add_12_51_groupi_n_3147 ,csa_tree_add_12_51_groupi_n_3417);
  or csa_tree_add_12_51_groupi_g17840(csa_tree_add_12_51_groupi_n_3946 ,csa_tree_add_12_51_groupi_n_3188 ,csa_tree_add_12_51_groupi_n_3348);
  or csa_tree_add_12_51_groupi_g17841(csa_tree_add_12_51_groupi_n_3945 ,csa_tree_add_12_51_groupi_n_3193 ,csa_tree_add_12_51_groupi_n_3365);
  or csa_tree_add_12_51_groupi_g17842(csa_tree_add_12_51_groupi_n_3944 ,csa_tree_add_12_51_groupi_n_3194 ,csa_tree_add_12_51_groupi_n_3338);
  or csa_tree_add_12_51_groupi_g17843(csa_tree_add_12_51_groupi_n_3943 ,csa_tree_add_12_51_groupi_n_2993 ,csa_tree_add_12_51_groupi_n_3416);
  or csa_tree_add_12_51_groupi_g17844(csa_tree_add_12_51_groupi_n_3942 ,csa_tree_add_12_51_groupi_n_3182 ,csa_tree_add_12_51_groupi_n_3342);
  or csa_tree_add_12_51_groupi_g17845(csa_tree_add_12_51_groupi_n_3941 ,csa_tree_add_12_51_groupi_n_3156 ,csa_tree_add_12_51_groupi_n_3420);
  or csa_tree_add_12_51_groupi_g17846(csa_tree_add_12_51_groupi_n_3940 ,csa_tree_add_12_51_groupi_n_3197 ,csa_tree_add_12_51_groupi_n_3398);
  or csa_tree_add_12_51_groupi_g17847(csa_tree_add_12_51_groupi_n_3939 ,csa_tree_add_12_51_groupi_n_3100 ,csa_tree_add_12_51_groupi_n_3418);
  or csa_tree_add_12_51_groupi_g17848(csa_tree_add_12_51_groupi_n_3938 ,csa_tree_add_12_51_groupi_n_3202 ,csa_tree_add_12_51_groupi_n_3325);
  or csa_tree_add_12_51_groupi_g17849(csa_tree_add_12_51_groupi_n_3937 ,csa_tree_add_12_51_groupi_n_3170 ,csa_tree_add_12_51_groupi_n_3411);
  or csa_tree_add_12_51_groupi_g17850(csa_tree_add_12_51_groupi_n_3936 ,csa_tree_add_12_51_groupi_n_3161 ,csa_tree_add_12_51_groupi_n_3410);
  or csa_tree_add_12_51_groupi_g17851(csa_tree_add_12_51_groupi_n_3935 ,csa_tree_add_12_51_groupi_n_3195 ,csa_tree_add_12_51_groupi_n_3324);
  or csa_tree_add_12_51_groupi_g17852(csa_tree_add_12_51_groupi_n_3934 ,csa_tree_add_12_51_groupi_n_3057 ,csa_tree_add_12_51_groupi_n_3405);
  or csa_tree_add_12_51_groupi_g17853(csa_tree_add_12_51_groupi_n_3933 ,csa_tree_add_12_51_groupi_n_3177 ,csa_tree_add_12_51_groupi_n_3286);
  or csa_tree_add_12_51_groupi_g17854(csa_tree_add_12_51_groupi_n_3932 ,csa_tree_add_12_51_groupi_n_2984 ,csa_tree_add_12_51_groupi_n_3413);
  or csa_tree_add_12_51_groupi_g17855(csa_tree_add_12_51_groupi_n_3931 ,csa_tree_add_12_51_groupi_n_3130 ,csa_tree_add_12_51_groupi_n_3403);
  or csa_tree_add_12_51_groupi_g17856(csa_tree_add_12_51_groupi_n_3930 ,csa_tree_add_12_51_groupi_n_3116 ,csa_tree_add_12_51_groupi_n_3402);
  or csa_tree_add_12_51_groupi_g17857(csa_tree_add_12_51_groupi_n_3929 ,csa_tree_add_12_51_groupi_n_3200 ,csa_tree_add_12_51_groupi_n_3429);
  or csa_tree_add_12_51_groupi_g17858(csa_tree_add_12_51_groupi_n_3928 ,csa_tree_add_12_51_groupi_n_3026 ,csa_tree_add_12_51_groupi_n_3346);
  or csa_tree_add_12_51_groupi_g17859(csa_tree_add_12_51_groupi_n_3927 ,csa_tree_add_12_51_groupi_n_2997 ,csa_tree_add_12_51_groupi_n_3340);
  or csa_tree_add_12_51_groupi_g17860(csa_tree_add_12_51_groupi_n_3926 ,csa_tree_add_12_51_groupi_n_2982 ,csa_tree_add_12_51_groupi_n_3369);
  or csa_tree_add_12_51_groupi_g17861(csa_tree_add_12_51_groupi_n_3925 ,csa_tree_add_12_51_groupi_n_3120 ,csa_tree_add_12_51_groupi_n_3389);
  or csa_tree_add_12_51_groupi_g17862(csa_tree_add_12_51_groupi_n_3924 ,csa_tree_add_12_51_groupi_n_2996 ,csa_tree_add_12_51_groupi_n_3378);
  or csa_tree_add_12_51_groupi_g17863(csa_tree_add_12_51_groupi_n_3923 ,csa_tree_add_12_51_groupi_n_3047 ,csa_tree_add_12_51_groupi_n_3354);
  or csa_tree_add_12_51_groupi_g17864(csa_tree_add_12_51_groupi_n_3922 ,csa_tree_add_12_51_groupi_n_3001 ,csa_tree_add_12_51_groupi_n_3375);
  or csa_tree_add_12_51_groupi_g17865(csa_tree_add_12_51_groupi_n_3921 ,csa_tree_add_12_51_groupi_n_3145 ,csa_tree_add_12_51_groupi_n_3344);
  or csa_tree_add_12_51_groupi_g17866(csa_tree_add_12_51_groupi_n_3920 ,csa_tree_add_12_51_groupi_n_3150 ,csa_tree_add_12_51_groupi_n_3397);
  or csa_tree_add_12_51_groupi_g17867(csa_tree_add_12_51_groupi_n_3919 ,csa_tree_add_12_51_groupi_n_3002 ,csa_tree_add_12_51_groupi_n_3374);
  or csa_tree_add_12_51_groupi_g17868(csa_tree_add_12_51_groupi_n_3918 ,csa_tree_add_12_51_groupi_n_3061 ,csa_tree_add_12_51_groupi_n_3390);
  or csa_tree_add_12_51_groupi_g17869(csa_tree_add_12_51_groupi_n_3917 ,csa_tree_add_12_51_groupi_n_3168 ,csa_tree_add_12_51_groupi_n_3360);
  or csa_tree_add_12_51_groupi_g17870(csa_tree_add_12_51_groupi_n_3916 ,csa_tree_add_12_51_groupi_n_3117 ,csa_tree_add_12_51_groupi_n_3382);
  or csa_tree_add_12_51_groupi_g17871(csa_tree_add_12_51_groupi_n_3915 ,csa_tree_add_12_51_groupi_n_3088 ,csa_tree_add_12_51_groupi_n_3377);
  or csa_tree_add_12_51_groupi_g17872(csa_tree_add_12_51_groupi_n_3914 ,csa_tree_add_12_51_groupi_n_3106 ,csa_tree_add_12_51_groupi_n_3345);
  or csa_tree_add_12_51_groupi_g17873(csa_tree_add_12_51_groupi_n_3913 ,csa_tree_add_12_51_groupi_n_3000 ,csa_tree_add_12_51_groupi_n_3341);
  or csa_tree_add_12_51_groupi_g17874(csa_tree_add_12_51_groupi_n_3912 ,csa_tree_add_12_51_groupi_n_3040 ,csa_tree_add_12_51_groupi_n_3393);
  or csa_tree_add_12_51_groupi_g17875(csa_tree_add_12_51_groupi_n_3911 ,csa_tree_add_12_51_groupi_n_3068 ,csa_tree_add_12_51_groupi_n_3366);
  or csa_tree_add_12_51_groupi_g17876(csa_tree_add_12_51_groupi_n_3910 ,csa_tree_add_12_51_groupi_n_3166 ,csa_tree_add_12_51_groupi_n_3353);
  or csa_tree_add_12_51_groupi_g17877(csa_tree_add_12_51_groupi_n_3909 ,csa_tree_add_12_51_groupi_n_3096 ,csa_tree_add_12_51_groupi_n_3394);
  or csa_tree_add_12_51_groupi_g17878(csa_tree_add_12_51_groupi_n_3908 ,csa_tree_add_12_51_groupi_n_3053 ,csa_tree_add_12_51_groupi_n_3370);
  or csa_tree_add_12_51_groupi_g17879(csa_tree_add_12_51_groupi_n_3907 ,csa_tree_add_12_51_groupi_n_3141 ,csa_tree_add_12_51_groupi_n_3337);
  or csa_tree_add_12_51_groupi_g17880(csa_tree_add_12_51_groupi_n_3906 ,csa_tree_add_12_51_groupi_n_3101 ,csa_tree_add_12_51_groupi_n_3351);
  or csa_tree_add_12_51_groupi_g17881(csa_tree_add_12_51_groupi_n_3905 ,csa_tree_add_12_51_groupi_n_3169 ,csa_tree_add_12_51_groupi_n_3379);
  or csa_tree_add_12_51_groupi_g17882(csa_tree_add_12_51_groupi_n_3904 ,csa_tree_add_12_51_groupi_n_3077 ,csa_tree_add_12_51_groupi_n_3381);
  or csa_tree_add_12_51_groupi_g17883(csa_tree_add_12_51_groupi_n_3903 ,csa_tree_add_12_51_groupi_n_3013 ,csa_tree_add_12_51_groupi_n_3391);
  or csa_tree_add_12_51_groupi_g17884(csa_tree_add_12_51_groupi_n_3902 ,csa_tree_add_12_51_groupi_n_3167 ,csa_tree_add_12_51_groupi_n_3371);
  or csa_tree_add_12_51_groupi_g17885(csa_tree_add_12_51_groupi_n_3901 ,csa_tree_add_12_51_groupi_n_2980 ,csa_tree_add_12_51_groupi_n_3336);
  or csa_tree_add_12_51_groupi_g17886(csa_tree_add_12_51_groupi_n_3900 ,csa_tree_add_12_51_groupi_n_3138 ,csa_tree_add_12_51_groupi_n_3349);
  or csa_tree_add_12_51_groupi_g17887(csa_tree_add_12_51_groupi_n_3899 ,csa_tree_add_12_51_groupi_n_3042 ,csa_tree_add_12_51_groupi_n_3359);
  or csa_tree_add_12_51_groupi_g17888(csa_tree_add_12_51_groupi_n_3898 ,csa_tree_add_12_51_groupi_n_2987 ,csa_tree_add_12_51_groupi_n_3387);
  or csa_tree_add_12_51_groupi_g17889(csa_tree_add_12_51_groupi_n_3897 ,csa_tree_add_12_51_groupi_n_3103 ,csa_tree_add_12_51_groupi_n_3385);
  or csa_tree_add_12_51_groupi_g17890(csa_tree_add_12_51_groupi_n_3896 ,csa_tree_add_12_51_groupi_n_3022 ,csa_tree_add_12_51_groupi_n_3347);
  or csa_tree_add_12_51_groupi_g17891(csa_tree_add_12_51_groupi_n_3895 ,csa_tree_add_12_51_groupi_n_3014 ,csa_tree_add_12_51_groupi_n_3364);
  or csa_tree_add_12_51_groupi_g17892(csa_tree_add_12_51_groupi_n_3894 ,csa_tree_add_12_51_groupi_n_3050 ,csa_tree_add_12_51_groupi_n_3386);
  or csa_tree_add_12_51_groupi_g17893(csa_tree_add_12_51_groupi_n_3893 ,csa_tree_add_12_51_groupi_n_3029 ,csa_tree_add_12_51_groupi_n_3376);
  or csa_tree_add_12_51_groupi_g17894(csa_tree_add_12_51_groupi_n_3892 ,csa_tree_add_12_51_groupi_n_3027 ,csa_tree_add_12_51_groupi_n_3367);
  or csa_tree_add_12_51_groupi_g17895(csa_tree_add_12_51_groupi_n_3891 ,csa_tree_add_12_51_groupi_n_3136 ,csa_tree_add_12_51_groupi_n_3355);
  or csa_tree_add_12_51_groupi_g17896(csa_tree_add_12_51_groupi_n_3890 ,csa_tree_add_12_51_groupi_n_3090 ,csa_tree_add_12_51_groupi_n_3395);
  or csa_tree_add_12_51_groupi_g17897(csa_tree_add_12_51_groupi_n_3889 ,csa_tree_add_12_51_groupi_n_3066 ,csa_tree_add_12_51_groupi_n_3373);
  or csa_tree_add_12_51_groupi_g17898(csa_tree_add_12_51_groupi_n_3888 ,csa_tree_add_12_51_groupi_n_3039 ,csa_tree_add_12_51_groupi_n_3399);
  or csa_tree_add_12_51_groupi_g17899(csa_tree_add_12_51_groupi_n_3887 ,csa_tree_add_12_51_groupi_n_3139 ,csa_tree_add_12_51_groupi_n_3392);
  or csa_tree_add_12_51_groupi_g17900(csa_tree_add_12_51_groupi_n_3886 ,csa_tree_add_12_51_groupi_n_3079 ,csa_tree_add_12_51_groupi_n_3357);
  or csa_tree_add_12_51_groupi_g17901(csa_tree_add_12_51_groupi_n_3885 ,csa_tree_add_12_51_groupi_n_2981 ,csa_tree_add_12_51_groupi_n_3388);
  nor csa_tree_add_12_51_groupi_g17902(csa_tree_add_12_51_groupi_n_3884 ,csa_tree_add_12_51_groupi_n_3534 ,csa_tree_add_12_51_groupi_n_3532);
  or csa_tree_add_12_51_groupi_g17903(csa_tree_add_12_51_groupi_n_3883 ,csa_tree_add_12_51_groupi_n_3533 ,csa_tree_add_12_51_groupi_n_3531);
  or csa_tree_add_12_51_groupi_g17904(csa_tree_add_12_51_groupi_n_3882 ,csa_tree_add_12_51_groupi_n_3162 ,csa_tree_add_12_51_groupi_n_3328);
  or csa_tree_add_12_51_groupi_g17905(csa_tree_add_12_51_groupi_n_3881 ,csa_tree_add_12_51_groupi_n_2988 ,csa_tree_add_12_51_groupi_n_3326);
  or csa_tree_add_12_51_groupi_g17906(csa_tree_add_12_51_groupi_n_3880 ,csa_tree_add_12_51_groupi_n_3158 ,csa_tree_add_12_51_groupi_n_3331);
  or csa_tree_add_12_51_groupi_g17907(csa_tree_add_12_51_groupi_n_3879 ,csa_tree_add_12_51_groupi_n_3128 ,csa_tree_add_12_51_groupi_n_3276);
  or csa_tree_add_12_51_groupi_g17908(csa_tree_add_12_51_groupi_n_3878 ,csa_tree_add_12_51_groupi_n_3034 ,csa_tree_add_12_51_groupi_n_3318);
  or csa_tree_add_12_51_groupi_g17909(csa_tree_add_12_51_groupi_n_3877 ,csa_tree_add_12_51_groupi_n_3098 ,csa_tree_add_12_51_groupi_n_3309);
  or csa_tree_add_12_51_groupi_g17910(csa_tree_add_12_51_groupi_n_3876 ,csa_tree_add_12_51_groupi_n_2999 ,csa_tree_add_12_51_groupi_n_3310);
  or csa_tree_add_12_51_groupi_g17911(csa_tree_add_12_51_groupi_n_3875 ,csa_tree_add_12_51_groupi_n_3104 ,csa_tree_add_12_51_groupi_n_3314);
  or csa_tree_add_12_51_groupi_g17912(csa_tree_add_12_51_groupi_n_3874 ,csa_tree_add_12_51_groupi_n_3146 ,csa_tree_add_12_51_groupi_n_3283);
  or csa_tree_add_12_51_groupi_g17913(csa_tree_add_12_51_groupi_n_3873 ,csa_tree_add_12_51_groupi_n_3115 ,csa_tree_add_12_51_groupi_n_3299);
  or csa_tree_add_12_51_groupi_g17914(csa_tree_add_12_51_groupi_n_3872 ,csa_tree_add_12_51_groupi_n_3072 ,csa_tree_add_12_51_groupi_n_3330);
  or csa_tree_add_12_51_groupi_g17915(csa_tree_add_12_51_groupi_n_3871 ,csa_tree_add_12_51_groupi_n_3114 ,csa_tree_add_12_51_groupi_n_3295);
  or csa_tree_add_12_51_groupi_g17916(csa_tree_add_12_51_groupi_n_3870 ,csa_tree_add_12_51_groupi_n_3032 ,csa_tree_add_12_51_groupi_n_3316);
  or csa_tree_add_12_51_groupi_g17917(csa_tree_add_12_51_groupi_n_3869 ,csa_tree_add_12_51_groupi_n_3163 ,csa_tree_add_12_51_groupi_n_3282);
  or csa_tree_add_12_51_groupi_g17918(csa_tree_add_12_51_groupi_n_3868 ,csa_tree_add_12_51_groupi_n_3065 ,csa_tree_add_12_51_groupi_n_3301);
  or csa_tree_add_12_51_groupi_g17919(csa_tree_add_12_51_groupi_n_3867 ,in2[2] ,csa_tree_add_12_51_groupi_n_3242);
  or csa_tree_add_12_51_groupi_g17920(csa_tree_add_12_51_groupi_n_3866 ,csa_tree_add_12_51_groupi_n_3087 ,csa_tree_add_12_51_groupi_n_3334);
  or csa_tree_add_12_51_groupi_g17921(csa_tree_add_12_51_groupi_n_3865 ,csa_tree_add_12_51_groupi_n_3152 ,csa_tree_add_12_51_groupi_n_3289);
  or csa_tree_add_12_51_groupi_g17922(csa_tree_add_12_51_groupi_n_3864 ,csa_tree_add_12_51_groupi_n_3020 ,csa_tree_add_12_51_groupi_n_3327);
  or csa_tree_add_12_51_groupi_g17923(csa_tree_add_12_51_groupi_n_3863 ,csa_tree_add_12_51_groupi_n_3144 ,csa_tree_add_12_51_groupi_n_3320);
  or csa_tree_add_12_51_groupi_g17924(csa_tree_add_12_51_groupi_n_3862 ,csa_tree_add_12_51_groupi_n_3083 ,csa_tree_add_12_51_groupi_n_3278);
  or csa_tree_add_12_51_groupi_g17925(csa_tree_add_12_51_groupi_n_3861 ,csa_tree_add_12_51_groupi_n_3109 ,csa_tree_add_12_51_groupi_n_3332);
  or csa_tree_add_12_51_groupi_g17926(csa_tree_add_12_51_groupi_n_3860 ,csa_tree_add_12_51_groupi_n_3143 ,csa_tree_add_12_51_groupi_n_3284);
  or csa_tree_add_12_51_groupi_g17927(csa_tree_add_12_51_groupi_n_3859 ,csa_tree_add_12_51_groupi_n_3148 ,csa_tree_add_12_51_groupi_n_3277);
  or csa_tree_add_12_51_groupi_g17928(csa_tree_add_12_51_groupi_n_3858 ,csa_tree_add_12_51_groupi_n_3142 ,csa_tree_add_12_51_groupi_n_3293);
  or csa_tree_add_12_51_groupi_g17929(csa_tree_add_12_51_groupi_n_3857 ,csa_tree_add_12_51_groupi_n_3125 ,csa_tree_add_12_51_groupi_n_3313);
  or csa_tree_add_12_51_groupi_g17930(csa_tree_add_12_51_groupi_n_3856 ,csa_tree_add_12_51_groupi_n_3089 ,csa_tree_add_12_51_groupi_n_3321);
  or csa_tree_add_12_51_groupi_g17931(csa_tree_add_12_51_groupi_n_3855 ,csa_tree_add_12_51_groupi_n_3030 ,csa_tree_add_12_51_groupi_n_3303);
  or csa_tree_add_12_51_groupi_g17932(csa_tree_add_12_51_groupi_n_3854 ,csa_tree_add_12_51_groupi_n_3049 ,csa_tree_add_12_51_groupi_n_3274);
  or csa_tree_add_12_51_groupi_g17933(csa_tree_add_12_51_groupi_n_3853 ,csa_tree_add_12_51_groupi_n_3105 ,csa_tree_add_12_51_groupi_n_3272);
  or csa_tree_add_12_51_groupi_g17934(csa_tree_add_12_51_groupi_n_3852 ,csa_tree_add_12_51_groupi_n_3108 ,csa_tree_add_12_51_groupi_n_3315);
  or csa_tree_add_12_51_groupi_g17935(csa_tree_add_12_51_groupi_n_3851 ,csa_tree_add_12_51_groupi_n_3228 ,csa_tree_add_12_51_groupi_n_3319);
  or csa_tree_add_12_51_groupi_g17936(csa_tree_add_12_51_groupi_n_3850 ,csa_tree_add_12_51_groupi_n_3153 ,csa_tree_add_12_51_groupi_n_3322);
  or csa_tree_add_12_51_groupi_g17937(csa_tree_add_12_51_groupi_n_3849 ,csa_tree_add_12_51_groupi_n_3151 ,csa_tree_add_12_51_groupi_n_3292);
  or csa_tree_add_12_51_groupi_g17938(csa_tree_add_12_51_groupi_n_3848 ,csa_tree_add_12_51_groupi_n_3171 ,csa_tree_add_12_51_groupi_n_3300);
  or csa_tree_add_12_51_groupi_g17939(csa_tree_add_12_51_groupi_n_3847 ,csa_tree_add_12_51_groupi_n_3149 ,csa_tree_add_12_51_groupi_n_3329);
  or csa_tree_add_12_51_groupi_g17940(csa_tree_add_12_51_groupi_n_3846 ,csa_tree_add_12_51_groupi_n_3051 ,csa_tree_add_12_51_groupi_n_3430);
  or csa_tree_add_12_51_groupi_g17941(csa_tree_add_12_51_groupi_n_3845 ,csa_tree_add_12_51_groupi_n_3006 ,csa_tree_add_12_51_groupi_n_3261);
  or csa_tree_add_12_51_groupi_g17942(csa_tree_add_12_51_groupi_n_3844 ,csa_tree_add_12_51_groupi_n_3038 ,csa_tree_add_12_51_groupi_n_3425);
  or csa_tree_add_12_51_groupi_g17943(csa_tree_add_12_51_groupi_n_3843 ,csa_tree_add_12_51_groupi_n_3010 ,csa_tree_add_12_51_groupi_n_3264);
  or csa_tree_add_12_51_groupi_g17944(csa_tree_add_12_51_groupi_n_3842 ,csa_tree_add_12_51_groupi_n_3121 ,csa_tree_add_12_51_groupi_n_3426);
  or csa_tree_add_12_51_groupi_g17945(csa_tree_add_12_51_groupi_n_3841 ,csa_tree_add_12_51_groupi_n_3129 ,csa_tree_add_12_51_groupi_n_3268);
  or csa_tree_add_12_51_groupi_g17946(csa_tree_add_12_51_groupi_n_3840 ,csa_tree_add_12_51_groupi_n_3123 ,csa_tree_add_12_51_groupi_n_3427);
  or csa_tree_add_12_51_groupi_g17947(csa_tree_add_12_51_groupi_n_3839 ,csa_tree_add_12_51_groupi_n_3118 ,csa_tree_add_12_51_groupi_n_3434);
  or csa_tree_add_12_51_groupi_g17948(csa_tree_add_12_51_groupi_n_3838 ,csa_tree_add_12_51_groupi_n_2990 ,csa_tree_add_12_51_groupi_n_3433);
  or csa_tree_add_12_51_groupi_g17949(csa_tree_add_12_51_groupi_n_3837 ,csa_tree_add_12_51_groupi_n_2991 ,csa_tree_add_12_51_groupi_n_3257);
  or csa_tree_add_12_51_groupi_g17950(csa_tree_add_12_51_groupi_n_3836 ,csa_tree_add_12_51_groupi_n_3064 ,csa_tree_add_12_51_groupi_n_3424);
  or csa_tree_add_12_51_groupi_g17951(csa_tree_add_12_51_groupi_n_3835 ,csa_tree_add_12_51_groupi_n_3009 ,csa_tree_add_12_51_groupi_n_3262);
  or csa_tree_add_12_51_groupi_g17952(csa_tree_add_12_51_groupi_n_3834 ,csa_tree_add_12_51_groupi_n_3063 ,csa_tree_add_12_51_groupi_n_3260);
  or csa_tree_add_12_51_groupi_g17953(csa_tree_add_12_51_groupi_n_3833 ,csa_tree_add_12_51_groupi_n_3137 ,csa_tree_add_12_51_groupi_n_3428);
  or csa_tree_add_12_51_groupi_g17954(csa_tree_add_12_51_groupi_n_3832 ,csa_tree_add_12_51_groupi_n_3025 ,csa_tree_add_12_51_groupi_n_3269);
  or csa_tree_add_12_51_groupi_g17955(csa_tree_add_12_51_groupi_n_3831 ,csa_tree_add_12_51_groupi_n_3126 ,csa_tree_add_12_51_groupi_n_3432);
  or csa_tree_add_12_51_groupi_g17956(csa_tree_add_12_51_groupi_n_3830 ,csa_tree_add_12_51_groupi_n_2989 ,csa_tree_add_12_51_groupi_n_3431);
  or csa_tree_add_12_51_groupi_g17957(csa_tree_add_12_51_groupi_n_3829 ,csa_tree_add_12_51_groupi_n_3528 ,csa_tree_add_12_51_groupi_n_3548);
  and csa_tree_add_12_51_groupi_g17958(csa_tree_add_12_51_groupi_n_3828 ,csa_tree_add_12_51_groupi_n_3528 ,csa_tree_add_12_51_groupi_n_3548);
  or csa_tree_add_12_51_groupi_g17959(csa_tree_add_12_51_groupi_n_3827 ,csa_tree_add_12_51_groupi_n_3540 ,csa_tree_add_12_51_groupi_n_3545);
  and csa_tree_add_12_51_groupi_g17960(csa_tree_add_12_51_groupi_n_3826 ,csa_tree_add_12_51_groupi_n_3540 ,csa_tree_add_12_51_groupi_n_3545);
  and csa_tree_add_12_51_groupi_g17961(csa_tree_add_12_51_groupi_n_3825 ,csa_tree_add_12_51_groupi_n_3522 ,csa_tree_add_12_51_groupi_n_3248);
  or csa_tree_add_12_51_groupi_g17962(csa_tree_add_12_51_groupi_n_3824 ,csa_tree_add_12_51_groupi_n_3537 ,csa_tree_add_12_51_groupi_n_3249);
  or csa_tree_add_12_51_groupi_g17963(csa_tree_add_12_51_groupi_n_3823 ,csa_tree_add_12_51_groupi_n_3549 ,csa_tree_add_12_51_groupi_n_3251);
  and csa_tree_add_12_51_groupi_g17964(csa_tree_add_12_51_groupi_n_3822 ,csa_tree_add_12_51_groupi_n_3537 ,csa_tree_add_12_51_groupi_n_3249);
  and csa_tree_add_12_51_groupi_g17965(csa_tree_add_12_51_groupi_n_3821 ,csa_tree_add_12_51_groupi_n_3549 ,csa_tree_add_12_51_groupi_n_3251);
  or csa_tree_add_12_51_groupi_g17966(csa_tree_add_12_51_groupi_n_3820 ,csa_tree_add_12_51_groupi_n_3522 ,csa_tree_add_12_51_groupi_n_3248);
  or csa_tree_add_12_51_groupi_g17967(csa_tree_add_12_51_groupi_n_3819 ,csa_tree_add_12_51_groupi_n_3525 ,csa_tree_add_12_51_groupi_n_3250);
  and csa_tree_add_12_51_groupi_g17968(csa_tree_add_12_51_groupi_n_3818 ,csa_tree_add_12_51_groupi_n_3525 ,csa_tree_add_12_51_groupi_n_3250);
  and csa_tree_add_12_51_groupi_g17969(csa_tree_add_12_51_groupi_n_3817 ,csa_tree_add_12_51_groupi_n_3252 ,csa_tree_add_12_51_groupi_n_3246);
  or csa_tree_add_12_51_groupi_g17970(csa_tree_add_12_51_groupi_n_3816 ,csa_tree_add_12_51_groupi_n_3252 ,csa_tree_add_12_51_groupi_n_3246);
  or csa_tree_add_12_51_groupi_g17971(csa_tree_add_12_51_groupi_n_3815 ,csa_tree_add_12_51_groupi_n_3536 ,csa_tree_add_12_51_groupi_n_3237);
  nor csa_tree_add_12_51_groupi_g17972(csa_tree_add_12_51_groupi_n_3814 ,csa_tree_add_12_51_groupi_n_3535 ,csa_tree_add_12_51_groupi_n_3238);
  nor csa_tree_add_12_51_groupi_g17973(csa_tree_add_12_51_groupi_n_3813 ,csa_tree_add_12_51_groupi_n_1089 ,csa_tree_add_12_51_groupi_n_143);
  nor csa_tree_add_12_51_groupi_g17974(csa_tree_add_12_51_groupi_n_3812 ,csa_tree_add_12_51_groupi_n_1170 ,csa_tree_add_12_51_groupi_n_142);
  nor csa_tree_add_12_51_groupi_g17975(csa_tree_add_12_51_groupi_n_3811 ,csa_tree_add_12_51_groupi_n_456 ,csa_tree_add_12_51_groupi_n_903);
  nor csa_tree_add_12_51_groupi_g17976(csa_tree_add_12_51_groupi_n_3810 ,csa_tree_add_12_51_groupi_n_3523 ,csa_tree_add_12_51_groupi_n_3240);
  or csa_tree_add_12_51_groupi_g17977(csa_tree_add_12_51_groupi_n_3809 ,csa_tree_add_12_51_groupi_n_3524 ,csa_tree_add_12_51_groupi_n_3239);
  or csa_tree_add_12_51_groupi_g17978(csa_tree_add_12_51_groupi_n_3808 ,csa_tree_add_12_51_groupi_n_2163 ,csa_tree_add_12_51_groupi_n_3233);
  nor csa_tree_add_12_51_groupi_g17979(csa_tree_add_12_51_groupi_n_3807 ,csa_tree_add_12_51_groupi_n_3509 ,csa_tree_add_12_51_groupi_n_3234);
  or csa_tree_add_12_51_groupi_g17980(csa_tree_add_12_51_groupi_n_3806 ,csa_tree_add_12_51_groupi_n_3547 ,csa_tree_add_12_51_groupi_n_3235);
  nor csa_tree_add_12_51_groupi_g17981(csa_tree_add_12_51_groupi_n_3805 ,csa_tree_add_12_51_groupi_n_3546 ,csa_tree_add_12_51_groupi_n_3236);
  or csa_tree_add_12_51_groupi_g17982(csa_tree_add_12_51_groupi_n_3804 ,csa_tree_add_12_51_groupi_n_3408 ,csa_tree_add_12_51_groupi_n_3223);
  and csa_tree_add_12_51_groupi_g17983(csa_tree_add_12_51_groupi_n_3803 ,csa_tree_add_12_51_groupi_n_3530 ,csa_tree_add_12_51_groupi_n_1914);
  or csa_tree_add_12_51_groupi_g17984(csa_tree_add_12_51_groupi_n_3802 ,csa_tree_add_12_51_groupi_n_3530 ,csa_tree_add_12_51_groupi_n_1914);
  or csa_tree_add_12_51_groupi_g17985(csa_tree_add_12_51_groupi_n_3801 ,csa_tree_add_12_51_groupi_n_1910 ,csa_tree_add_12_51_groupi_n_3529);
  and csa_tree_add_12_51_groupi_g17986(csa_tree_add_12_51_groupi_n_3800 ,csa_tree_add_12_51_groupi_n_1910 ,csa_tree_add_12_51_groupi_n_3529);
  and csa_tree_add_12_51_groupi_g17987(csa_tree_add_12_51_groupi_n_3799 ,csa_tree_add_12_51_groupi_n_1912 ,csa_tree_add_12_51_groupi_n_3247);
  or csa_tree_add_12_51_groupi_g17988(csa_tree_add_12_51_groupi_n_3798 ,csa_tree_add_12_51_groupi_n_1912 ,csa_tree_add_12_51_groupi_n_3247);
  or csa_tree_add_12_51_groupi_g17989(csa_tree_add_12_51_groupi_n_3797 ,csa_tree_add_12_51_groupi_n_3208 ,csa_tree_add_12_51_groupi_n_3219);
  or csa_tree_add_12_51_groupi_g17990(csa_tree_add_12_51_groupi_n_3796 ,csa_tree_add_12_51_groupi_n_3212 ,csa_tree_add_12_51_groupi_n_3224);
  nor csa_tree_add_12_51_groupi_g17991(csa_tree_add_12_51_groupi_n_3795 ,csa_tree_add_12_51_groupi_n_451 ,csa_tree_add_12_51_groupi_n_1236);
  nor csa_tree_add_12_51_groupi_g17992(csa_tree_add_12_51_groupi_n_3794 ,csa_tree_add_12_51_groupi_n_2959 ,csa_tree_add_12_51_groupi_n_3519);
  or csa_tree_add_12_51_groupi_g17993(csa_tree_add_12_51_groupi_n_3793 ,csa_tree_add_12_51_groupi_n_2958 ,csa_tree_add_12_51_groupi_n_3520);
  or csa_tree_add_12_51_groupi_g17994(csa_tree_add_12_51_groupi_n_3792 ,csa_tree_add_12_51_groupi_n_2955 ,csa_tree_add_12_51_groupi_n_3518);
  nor csa_tree_add_12_51_groupi_g17995(csa_tree_add_12_51_groupi_n_3791 ,csa_tree_add_12_51_groupi_n_2951 ,csa_tree_add_12_51_groupi_n_3538);
  and csa_tree_add_12_51_groupi_g17996(csa_tree_add_12_51_groupi_n_3790 ,csa_tree_add_12_51_groupi_n_2955 ,csa_tree_add_12_51_groupi_n_3518);
  or csa_tree_add_12_51_groupi_g17997(csa_tree_add_12_51_groupi_n_3789 ,csa_tree_add_12_51_groupi_n_2950 ,csa_tree_add_12_51_groupi_n_3539);
  nor csa_tree_add_12_51_groupi_g17998(csa_tree_add_12_51_groupi_n_3788 ,csa_tree_add_12_51_groupi_n_1527 ,csa_tree_add_12_51_groupi_n_699);
  nor csa_tree_add_12_51_groupi_g17999(csa_tree_add_12_51_groupi_n_3787 ,csa_tree_add_12_51_groupi_n_1227 ,csa_tree_add_12_51_groupi_n_146);
  or csa_tree_add_12_51_groupi_g18000(csa_tree_add_12_51_groupi_n_3786 ,csa_tree_add_12_51_groupi_n_2673 ,csa_tree_add_12_51_groupi_n_2966);
  or csa_tree_add_12_51_groupi_g18001(csa_tree_add_12_51_groupi_n_3785 ,csa_tree_add_12_51_groupi_n_2678 ,csa_tree_add_12_51_groupi_n_2964);
  nor csa_tree_add_12_51_groupi_g18002(csa_tree_add_12_51_groupi_n_3784 ,csa_tree_add_12_51_groupi_n_1476 ,csa_tree_add_12_51_groupi_n_127);
  nor csa_tree_add_12_51_groupi_g18003(csa_tree_add_12_51_groupi_n_3783 ,csa_tree_add_12_51_groupi_n_1152 ,csa_tree_add_12_51_groupi_n_130);
  nor csa_tree_add_12_51_groupi_g18004(csa_tree_add_12_51_groupi_n_3782 ,csa_tree_add_12_51_groupi_n_1320 ,csa_tree_add_12_51_groupi_n_137);
  nor csa_tree_add_12_51_groupi_g18005(csa_tree_add_12_51_groupi_n_3781 ,csa_tree_add_12_51_groupi_n_1359 ,csa_tree_add_12_51_groupi_n_295);
  or csa_tree_add_12_51_groupi_g18006(csa_tree_add_12_51_groupi_n_3780 ,csa_tree_add_12_51_groupi_n_131 ,csa_tree_add_12_51_groupi_n_2969);
  or csa_tree_add_12_51_groupi_g18007(csa_tree_add_12_51_groupi_n_3779 ,csa_tree_add_12_51_groupi_n_149 ,csa_tree_add_12_51_groupi_n_2968);
  or csa_tree_add_12_51_groupi_g18008(csa_tree_add_12_51_groupi_n_3778 ,csa_tree_add_12_51_groupi_n_146 ,csa_tree_add_12_51_groupi_n_2971);
  or csa_tree_add_12_51_groupi_g18009(csa_tree_add_12_51_groupi_n_3777 ,csa_tree_add_12_51_groupi_n_700 ,csa_tree_add_12_51_groupi_n_2973);
  or csa_tree_add_12_51_groupi_g18010(csa_tree_add_12_51_groupi_n_3776 ,csa_tree_add_12_51_groupi_n_1047 ,csa_tree_add_12_51_groupi_n_2978);
  or csa_tree_add_12_51_groupi_g18011(csa_tree_add_12_51_groupi_n_3775 ,csa_tree_add_12_51_groupi_n_229 ,csa_tree_add_12_51_groupi_n_2974);
  or csa_tree_add_12_51_groupi_g18012(csa_tree_add_12_51_groupi_n_3774 ,csa_tree_add_12_51_groupi_n_134 ,csa_tree_add_12_51_groupi_n_2970);
  or csa_tree_add_12_51_groupi_g18013(csa_tree_add_12_51_groupi_n_3773 ,csa_tree_add_12_51_groupi_n_457 ,csa_tree_add_12_51_groupi_n_2977);
  or csa_tree_add_12_51_groupi_g18014(csa_tree_add_12_51_groupi_n_3772 ,csa_tree_add_12_51_groupi_n_451 ,csa_tree_add_12_51_groupi_n_2972);
  or csa_tree_add_12_51_groupi_g18015(csa_tree_add_12_51_groupi_n_3771 ,csa_tree_add_12_51_groupi_n_1050 ,csa_tree_add_12_51_groupi_n_2975);
  or csa_tree_add_12_51_groupi_g18016(csa_tree_add_12_51_groupi_n_3770 ,csa_tree_add_12_51_groupi_n_409 ,csa_tree_add_12_51_groupi_n_2967);
  or csa_tree_add_12_51_groupi_g18017(csa_tree_add_12_51_groupi_n_3769 ,csa_tree_add_12_51_groupi_n_128 ,csa_tree_add_12_51_groupi_n_2976);
  and csa_tree_add_12_51_groupi_g18018(csa_tree_add_12_51_groupi_n_3972 ,csa_tree_add_12_51_groupi_n_2828 ,csa_tree_add_12_51_groupi_n_3435);
  or csa_tree_add_12_51_groupi_g18019(csa_tree_add_12_51_groupi_n_3768 ,csa_tree_add_12_51_groupi_n_140 ,csa_tree_add_12_51_groupi_n_3205);
  or csa_tree_add_12_51_groupi_g18020(csa_tree_add_12_51_groupi_n_3767 ,csa_tree_add_12_51_groupi_n_137 ,csa_tree_add_12_51_groupi_n_3204);
  or csa_tree_add_12_51_groupi_g18021(csa_tree_add_12_51_groupi_n_3766 ,csa_tree_add_12_51_groupi_n_143 ,csa_tree_add_12_51_groupi_n_3206);
  and csa_tree_add_12_51_groupi_g18022(csa_tree_add_12_51_groupi_n_3971 ,csa_tree_add_12_51_groupi_n_2426 ,csa_tree_add_12_51_groupi_n_3480);
  nor csa_tree_add_12_51_groupi_g18023(csa_tree_add_12_51_groupi_n_3763 ,csa_tree_add_12_51_groupi_n_549 ,csa_tree_add_12_51_groupi_n_1182);
  nor csa_tree_add_12_51_groupi_g18024(csa_tree_add_12_51_groupi_n_3762 ,csa_tree_add_12_51_groupi_n_1173 ,csa_tree_add_12_51_groupi_n_295);
  nor csa_tree_add_12_51_groupi_g18025(csa_tree_add_12_51_groupi_n_3761 ,csa_tree_add_12_51_groupi_n_697 ,csa_tree_add_12_51_groupi_n_957);
  nor csa_tree_add_12_51_groupi_g18026(csa_tree_add_12_51_groupi_n_3760 ,csa_tree_add_12_51_groupi_n_531 ,csa_tree_add_12_51_groupi_n_870);
  nor csa_tree_add_12_51_groupi_g18027(csa_tree_add_12_51_groupi_n_3759 ,csa_tree_add_12_51_groupi_n_1691 ,csa_tree_add_12_51_groupi_n_1181);
  nor csa_tree_add_12_51_groupi_g18028(csa_tree_add_12_51_groupi_n_3758 ,csa_tree_add_12_51_groupi_n_1802 ,csa_tree_add_12_51_groupi_n_873);
  nor csa_tree_add_12_51_groupi_g18029(csa_tree_add_12_51_groupi_n_3757 ,csa_tree_add_12_51_groupi_n_1692 ,csa_tree_add_12_51_groupi_n_1226);
  nor csa_tree_add_12_51_groupi_g18030(csa_tree_add_12_51_groupi_n_3756 ,csa_tree_add_12_51_groupi_n_1572 ,csa_tree_add_12_51_groupi_n_887);
  nor csa_tree_add_12_51_groupi_g18031(csa_tree_add_12_51_groupi_n_3755 ,csa_tree_add_12_51_groupi_n_1803 ,csa_tree_add_12_51_groupi_n_1154);
  nor csa_tree_add_12_51_groupi_g18032(csa_tree_add_12_51_groupi_n_3754 ,csa_tree_add_12_51_groupi_n_1092 ,csa_tree_add_12_51_groupi_n_462);
  nor csa_tree_add_12_51_groupi_g18033(csa_tree_add_12_51_groupi_n_3753 ,csa_tree_add_12_51_groupi_n_1806 ,csa_tree_add_12_51_groupi_n_1166);
  nor csa_tree_add_12_51_groupi_g18034(csa_tree_add_12_51_groupi_n_3752 ,csa_tree_add_12_51_groupi_n_1146 ,csa_tree_add_12_51_groupi_n_310);
  nor csa_tree_add_12_51_groupi_g18035(csa_tree_add_12_51_groupi_n_3751 ,csa_tree_add_12_51_groupi_n_1524 ,csa_tree_add_12_51_groupi_n_232);
  nor csa_tree_add_12_51_groupi_g18036(csa_tree_add_12_51_groupi_n_3750 ,csa_tree_add_12_51_groupi_n_1077 ,csa_tree_add_12_51_groupi_n_220);
  nor csa_tree_add_12_51_groupi_g18037(csa_tree_add_12_51_groupi_n_3749 ,csa_tree_add_12_51_groupi_n_1140 ,csa_tree_add_12_51_groupi_n_289);
  nor csa_tree_add_12_51_groupi_g18038(csa_tree_add_12_51_groupi_n_3748 ,csa_tree_add_12_51_groupi_n_1386 ,csa_tree_add_12_51_groupi_n_372);
  nor csa_tree_add_12_51_groupi_g18039(csa_tree_add_12_51_groupi_n_3747 ,csa_tree_add_12_51_groupi_n_696 ,csa_tree_add_12_51_groupi_n_927);
  nor csa_tree_add_12_51_groupi_g18040(csa_tree_add_12_51_groupi_n_3746 ,csa_tree_add_12_51_groupi_n_505 ,csa_tree_add_12_51_groupi_n_876);
  nor csa_tree_add_12_51_groupi_g18041(csa_tree_add_12_51_groupi_n_3745 ,csa_tree_add_12_51_groupi_n_1223 ,csa_tree_add_12_51_groupi_n_208);
  nor csa_tree_add_12_51_groupi_g18042(csa_tree_add_12_51_groupi_n_3744 ,csa_tree_add_12_51_groupi_n_1311 ,csa_tree_add_12_51_groupi_n_421);
  nor csa_tree_add_12_51_groupi_g18043(csa_tree_add_12_51_groupi_n_3743 ,csa_tree_add_12_51_groupi_n_1467 ,csa_tree_add_12_51_groupi_n_1373);
  nor csa_tree_add_12_51_groupi_g18044(csa_tree_add_12_51_groupi_n_3742 ,csa_tree_add_12_51_groupi_n_1470 ,csa_tree_add_12_51_groupi_n_1175);
  nor csa_tree_add_12_51_groupi_g18045(csa_tree_add_12_51_groupi_n_3741 ,csa_tree_add_12_51_groupi_n_532 ,csa_tree_add_12_51_groupi_n_902);
  nor csa_tree_add_12_51_groupi_g18046(csa_tree_add_12_51_groupi_n_3740 ,csa_tree_add_12_51_groupi_n_658 ,csa_tree_add_12_51_groupi_n_1151);
  nor csa_tree_add_12_51_groupi_g18047(csa_tree_add_12_51_groupi_n_3739 ,csa_tree_add_12_51_groupi_n_694 ,csa_tree_add_12_51_groupi_n_1260);
  nor csa_tree_add_12_51_groupi_g18048(csa_tree_add_12_51_groupi_n_3738 ,csa_tree_add_12_51_groupi_n_1509 ,csa_tree_add_12_51_groupi_n_307);
  nor csa_tree_add_12_51_groupi_g18049(csa_tree_add_12_51_groupi_n_3737 ,csa_tree_add_12_51_groupi_n_528 ,csa_tree_add_12_51_groupi_n_873);
  nor csa_tree_add_12_51_groupi_g18050(csa_tree_add_12_51_groupi_n_3736 ,csa_tree_add_12_51_groupi_n_514 ,csa_tree_add_12_51_groupi_n_963);
  nor csa_tree_add_12_51_groupi_g18051(csa_tree_add_12_51_groupi_n_3735 ,csa_tree_add_12_51_groupi_n_537 ,csa_tree_add_12_51_groupi_n_1248);
  nor csa_tree_add_12_51_groupi_g18052(csa_tree_add_12_51_groupi_n_3734 ,csa_tree_add_12_51_groupi_n_1809 ,csa_tree_add_12_51_groupi_n_1550);
  nor csa_tree_add_12_51_groupi_g18053(csa_tree_add_12_51_groupi_n_3733 ,csa_tree_add_12_51_groupi_n_573 ,csa_tree_add_12_51_groupi_n_879);
  nor csa_tree_add_12_51_groupi_g18054(csa_tree_add_12_51_groupi_n_3732 ,csa_tree_add_12_51_groupi_n_1697 ,csa_tree_add_12_51_groupi_n_872);
  nor csa_tree_add_12_51_groupi_g18055(csa_tree_add_12_51_groupi_n_3731 ,csa_tree_add_12_51_groupi_n_648 ,csa_tree_add_12_51_groupi_n_962);
  nor csa_tree_add_12_51_groupi_g18056(csa_tree_add_12_51_groupi_n_3730 ,csa_tree_add_12_51_groupi_n_595 ,csa_tree_add_12_51_groupi_n_870);
  nor csa_tree_add_12_51_groupi_g18057(csa_tree_add_12_51_groupi_n_3729 ,csa_tree_add_12_51_groupi_n_1736 ,csa_tree_add_12_51_groupi_n_1080);
  nor csa_tree_add_12_51_groupi_g18058(csa_tree_add_12_51_groupi_n_3728 ,csa_tree_add_12_51_groupi_n_556 ,csa_tree_add_12_51_groupi_n_926);
  nor csa_tree_add_12_51_groupi_g18059(csa_tree_add_12_51_groupi_n_3727 ,csa_tree_add_12_51_groupi_n_652 ,csa_tree_add_12_51_groupi_n_1143);
  nor csa_tree_add_12_51_groupi_g18060(csa_tree_add_12_51_groupi_n_3726 ,csa_tree_add_12_51_groupi_n_1566 ,csa_tree_add_12_51_groupi_n_878);
  nor csa_tree_add_12_51_groupi_g18061(csa_tree_add_12_51_groupi_n_3725 ,csa_tree_add_12_51_groupi_n_585 ,csa_tree_add_12_51_groupi_n_1088);
  nor csa_tree_add_12_51_groupi_g18062(csa_tree_add_12_51_groupi_n_3724 ,csa_tree_add_12_51_groupi_n_1734 ,csa_tree_add_12_51_groupi_n_1104);
  nor csa_tree_add_12_51_groupi_g18063(csa_tree_add_12_51_groupi_n_3723 ,csa_tree_add_12_51_groupi_n_636 ,csa_tree_add_12_51_groupi_n_1137);
  nor csa_tree_add_12_51_groupi_g18064(csa_tree_add_12_51_groupi_n_3722 ,csa_tree_add_12_51_groupi_n_678 ,csa_tree_add_12_51_groupi_n_1386);
  nor csa_tree_add_12_51_groupi_g18065(csa_tree_add_12_51_groupi_n_3721 ,csa_tree_add_12_51_groupi_n_610 ,csa_tree_add_12_51_groupi_n_1325);
  nor csa_tree_add_12_51_groupi_g18066(csa_tree_add_12_51_groupi_n_3720 ,csa_tree_add_12_51_groupi_n_1758 ,csa_tree_add_12_51_groupi_n_956);
  nor csa_tree_add_12_51_groupi_g18067(csa_tree_add_12_51_groupi_n_3719 ,csa_tree_add_12_51_groupi_n_1737 ,csa_tree_add_12_51_groupi_n_1157);
  nor csa_tree_add_12_51_groupi_g18068(csa_tree_add_12_51_groupi_n_3718 ,csa_tree_add_12_51_groupi_n_579 ,csa_tree_add_12_51_groupi_n_1103);
  nor csa_tree_add_12_51_groupi_g18069(csa_tree_add_12_51_groupi_n_3717 ,csa_tree_add_12_51_groupi_n_1740 ,csa_tree_add_12_51_groupi_n_1169);
  nor csa_tree_add_12_51_groupi_g18070(csa_tree_add_12_51_groupi_n_3716 ,csa_tree_add_12_51_groupi_n_615 ,csa_tree_add_12_51_groupi_n_1158);
  nor csa_tree_add_12_51_groupi_g18071(csa_tree_add_12_51_groupi_n_3715 ,csa_tree_add_12_51_groupi_n_589 ,csa_tree_add_12_51_groupi_n_1170);
  nor csa_tree_add_12_51_groupi_g18072(csa_tree_add_12_51_groupi_n_3714 ,csa_tree_add_12_51_groupi_n_1761 ,csa_tree_add_12_51_groupi_n_1142);
  nor csa_tree_add_12_51_groupi_g18073(csa_tree_add_12_51_groupi_n_3713 ,csa_tree_add_12_51_groupi_n_1794 ,csa_tree_add_12_51_groupi_n_1089);
  nor csa_tree_add_12_51_groupi_g18074(csa_tree_add_12_51_groupi_n_3712 ,csa_tree_add_12_51_groupi_n_1707 ,csa_tree_add_12_51_groupi_n_902);
  nor csa_tree_add_12_51_groupi_g18075(csa_tree_add_12_51_groupi_n_3711 ,csa_tree_add_12_51_groupi_n_640 ,csa_tree_add_12_51_groupi_n_1365);
  nor csa_tree_add_12_51_groupi_g18076(csa_tree_add_12_51_groupi_n_3710 ,csa_tree_add_12_51_groupi_n_1812 ,csa_tree_add_12_51_groupi_n_1260);
  nor csa_tree_add_12_51_groupi_g18077(csa_tree_add_12_51_groupi_n_3709 ,csa_tree_add_12_51_groupi_n_1749 ,csa_tree_add_12_51_groupi_n_1364);
  nor csa_tree_add_12_51_groupi_g18078(csa_tree_add_12_51_groupi_n_3708 ,csa_tree_add_12_51_groupi_n_1772 ,csa_tree_add_12_51_groupi_n_876);
  nor csa_tree_add_12_51_groupi_g18079(csa_tree_add_12_51_groupi_n_3707 ,csa_tree_add_12_51_groupi_n_1710 ,csa_tree_add_12_51_groupi_n_1359);
  nor csa_tree_add_12_51_groupi_g18080(csa_tree_add_12_51_groupi_n_3706 ,csa_tree_add_12_51_groupi_n_1770 ,csa_tree_add_12_51_groupi_n_1167);
  nor csa_tree_add_12_51_groupi_g18081(csa_tree_add_12_51_groupi_n_3705 ,csa_tree_add_12_51_groupi_n_1782 ,csa_tree_add_12_51_groupi_n_1319);
  nor csa_tree_add_12_51_groupi_g18082(csa_tree_add_12_51_groupi_n_3704 ,csa_tree_add_12_51_groupi_n_1704 ,csa_tree_add_12_51_groupi_n_1088);
  nor csa_tree_add_12_51_groupi_g18083(csa_tree_add_12_51_groupi_n_3703 ,csa_tree_add_12_51_groupi_n_1785 ,csa_tree_add_12_51_groupi_n_903);
  nor csa_tree_add_12_51_groupi_g18084(csa_tree_add_12_51_groupi_n_3702 ,csa_tree_add_12_51_groupi_n_514 ,csa_tree_add_12_51_groupi_n_1526);
  nor csa_tree_add_12_51_groupi_g18085(csa_tree_add_12_51_groupi_n_3701 ,csa_tree_add_12_51_groupi_n_1767 ,csa_tree_add_12_51_groupi_n_875);
  nor csa_tree_add_12_51_groupi_g18086(csa_tree_add_12_51_groupi_n_3700 ,csa_tree_add_12_51_groupi_n_1779 ,csa_tree_add_12_51_groupi_n_1079);
  nor csa_tree_add_12_51_groupi_g18087(csa_tree_add_12_51_groupi_n_3699 ,csa_tree_add_12_51_groupi_n_1374 ,csa_tree_add_12_51_groupi_n_468);
  nor csa_tree_add_12_51_groupi_g18088(csa_tree_add_12_51_groupi_n_3698 ,csa_tree_add_12_51_groupi_n_1797 ,csa_tree_add_12_51_groupi_n_1169);
  nor csa_tree_add_12_51_groupi_g18089(csa_tree_add_12_51_groupi_n_3697 ,csa_tree_add_12_51_groupi_n_1176 ,csa_tree_add_12_51_groupi_n_186);
  nor csa_tree_add_12_51_groupi_g18090(csa_tree_add_12_51_groupi_n_3696 ,csa_tree_add_12_51_groupi_n_1773 ,csa_tree_add_12_51_groupi_n_1136);
  nor csa_tree_add_12_51_groupi_g18091(csa_tree_add_12_51_groupi_n_3695 ,csa_tree_add_12_51_groupi_n_567 ,csa_tree_add_12_51_groupi_n_1475);
  nor csa_tree_add_12_51_groupi_g18092(csa_tree_add_12_51_groupi_n_3694 ,csa_tree_add_12_51_groupi_n_1358 ,csa_tree_add_12_51_groupi_n_274);
  nor csa_tree_add_12_51_groupi_g18093(csa_tree_add_12_51_groupi_n_3693 ,csa_tree_add_12_51_groupi_n_1800 ,csa_tree_add_12_51_groupi_n_1116);
  nor csa_tree_add_12_51_groupi_g18094(csa_tree_add_12_51_groupi_n_3692 ,csa_tree_add_12_51_groupi_n_558 ,csa_tree_add_12_51_groupi_n_1152);
  nor csa_tree_add_12_51_groupi_g18095(csa_tree_add_12_51_groupi_n_3691 ,csa_tree_add_12_51_groupi_n_1527 ,csa_tree_add_12_51_groupi_n_214);
  nor csa_tree_add_12_51_groupi_g18096(csa_tree_add_12_51_groupi_n_3690 ,csa_tree_add_12_51_groupi_n_1727 ,csa_tree_add_12_51_groupi_n_875);
  nor csa_tree_add_12_51_groupi_g18097(csa_tree_add_12_51_groupi_n_3689 ,csa_tree_add_12_51_groupi_n_1745 ,csa_tree_add_12_51_groupi_n_1166);
  nor csa_tree_add_12_51_groupi_g18098(csa_tree_add_12_51_groupi_n_3688 ,csa_tree_add_12_51_groupi_n_1752 ,csa_tree_add_12_51_groupi_n_1310);
  nor csa_tree_add_12_51_groupi_g18099(csa_tree_add_12_51_groupi_n_3687 ,csa_tree_add_12_51_groupi_n_1725 ,csa_tree_add_12_51_groupi_n_1508);
  nor csa_tree_add_12_51_groupi_g18100(csa_tree_add_12_51_groupi_n_3686 ,csa_tree_add_12_51_groupi_n_1695 ,csa_tree_add_12_51_groupi_n_1502);
  nor csa_tree_add_12_51_groupi_g18101(csa_tree_add_12_51_groupi_n_3685 ,csa_tree_add_12_51_groupi_n_1116 ,csa_tree_add_12_51_groupi_n_243);
  nor csa_tree_add_12_51_groupi_g18102(csa_tree_add_12_51_groupi_n_3684 ,csa_tree_add_12_51_groupi_n_1764 ,csa_tree_add_12_51_groupi_n_1115);
  nor csa_tree_add_12_51_groupi_g18103(csa_tree_add_12_51_groupi_n_3683 ,csa_tree_add_12_51_groupi_n_1755 ,csa_tree_add_12_51_groupi_n_1358);
  nor csa_tree_add_12_51_groupi_g18104(csa_tree_add_12_51_groupi_n_3682 ,csa_tree_add_12_51_groupi_n_1776 ,csa_tree_add_12_51_groupi_n_1181);
  nor csa_tree_add_12_51_groupi_g18105(csa_tree_add_12_51_groupi_n_3681 ,csa_tree_add_12_51_groupi_n_1728 ,csa_tree_add_12_51_groupi_n_1523);
  nor csa_tree_add_12_51_groupi_g18106(csa_tree_add_12_51_groupi_n_3680 ,csa_tree_add_12_51_groupi_n_1743 ,csa_tree_add_12_51_groupi_n_1223);
  nor csa_tree_add_12_51_groupi_g18107(csa_tree_add_12_51_groupi_n_3679 ,csa_tree_add_12_51_groupi_n_1247 ,csa_tree_add_12_51_groupi_n_291);
  nor csa_tree_add_12_51_groupi_g18108(csa_tree_add_12_51_groupi_n_3678 ,csa_tree_add_12_51_groupi_n_1746 ,csa_tree_add_12_51_groupi_n_1178);
  nor csa_tree_add_12_51_groupi_g18109(csa_tree_add_12_51_groupi_n_3677 ,csa_tree_add_12_51_groupi_n_1698 ,csa_tree_add_12_51_groupi_n_1149);
  nor csa_tree_add_12_51_groupi_g18110(csa_tree_add_12_51_groupi_n_3676 ,csa_tree_add_12_51_groupi_n_1722 ,csa_tree_add_12_51_groupi_n_1115);
  nor csa_tree_add_12_51_groupi_g18111(csa_tree_add_12_51_groupi_n_3675 ,csa_tree_add_12_51_groupi_n_1788 ,csa_tree_add_12_51_groupi_n_1224);
  nor csa_tree_add_12_51_groupi_g18112(csa_tree_add_12_51_groupi_n_3674 ,csa_tree_add_12_51_groupi_n_1509 ,csa_tree_add_12_51_groupi_n_357);
  nor csa_tree_add_12_51_groupi_g18113(csa_tree_add_12_51_groupi_n_3673 ,csa_tree_add_12_51_groupi_n_1179 ,csa_tree_add_12_51_groupi_n_225);
  nor csa_tree_add_12_51_groupi_g18114(csa_tree_add_12_51_groupi_n_3672 ,csa_tree_add_12_51_groupi_n_1236 ,csa_tree_add_12_51_groupi_n_433);
  nor csa_tree_add_12_51_groupi_g18115(csa_tree_add_12_51_groupi_n_3671 ,csa_tree_add_12_51_groupi_n_1476 ,csa_tree_add_12_51_groupi_n_418);
  nor csa_tree_add_12_51_groupi_g18116(csa_tree_add_12_51_groupi_n_3670 ,csa_tree_add_12_51_groupi_n_1731 ,csa_tree_add_12_51_groupi_n_1385);
  nor csa_tree_add_12_51_groupi_g18117(csa_tree_add_12_51_groupi_n_3669 ,csa_tree_add_12_51_groupi_n_1320 ,csa_tree_add_12_51_groupi_n_366);
  nor csa_tree_add_12_51_groupi_g18118(csa_tree_add_12_51_groupi_n_3668 ,csa_tree_add_12_51_groupi_n_1475 ,csa_tree_add_12_51_groupi_n_237);
  nor csa_tree_add_12_51_groupi_g18119(csa_tree_add_12_51_groupi_n_3667 ,csa_tree_add_12_51_groupi_n_1715 ,csa_tree_add_12_51_groupi_n_1179);
  nor csa_tree_add_12_51_groupi_g18120(csa_tree_add_12_51_groupi_n_3666 ,csa_tree_add_12_51_groupi_n_1701 ,csa_tree_add_12_51_groupi_n_1079);
  nor csa_tree_add_12_51_groupi_g18121(csa_tree_add_12_51_groupi_n_3665 ,csa_tree_add_12_51_groupi_n_1713 ,csa_tree_add_12_51_groupi_n_1259);
  nor csa_tree_add_12_51_groupi_g18122(csa_tree_add_12_51_groupi_n_3664 ,csa_tree_add_12_51_groupi_n_1503 ,csa_tree_add_12_51_groupi_n_334);
  nor csa_tree_add_12_51_groupi_g18123(csa_tree_add_12_51_groupi_n_3663 ,csa_tree_add_12_51_groupi_n_1364 ,csa_tree_add_12_51_groupi_n_340);
  nor csa_tree_add_12_51_groupi_g18124(csa_tree_add_12_51_groupi_n_3662 ,csa_tree_add_12_51_groupi_n_1157 ,csa_tree_add_12_51_groupi_n_198);
  nor csa_tree_add_12_51_groupi_g18125(csa_tree_add_12_51_groupi_n_3661 ,csa_tree_add_12_51_groupi_n_1182 ,csa_tree_add_12_51_groupi_n_301);
  or csa_tree_add_12_51_groupi_g18126(csa_tree_add_12_51_groupi_n_3660 ,csa_tree_add_12_51_groupi_n_2677 ,csa_tree_add_12_51_groupi_n_2965);
  nor csa_tree_add_12_51_groupi_g18127(csa_tree_add_12_51_groupi_n_3659 ,csa_tree_add_12_51_groupi_n_1406 ,csa_tree_add_12_51_groupi_n_1151);
  nor csa_tree_add_12_51_groupi_g18128(csa_tree_add_12_51_groupi_n_3658 ,csa_tree_add_12_51_groupi_n_1259 ,csa_tree_add_12_51_groupi_n_184);
  nor csa_tree_add_12_51_groupi_g18129(csa_tree_add_12_51_groupi_n_3657 ,csa_tree_add_12_51_groupi_n_1716 ,csa_tree_add_12_51_groupi_n_1145);
  nor csa_tree_add_12_51_groupi_g18130(csa_tree_add_12_51_groupi_n_3656 ,csa_tree_add_12_51_groupi_n_1719 ,csa_tree_add_12_51_groupi_n_869);
  nor csa_tree_add_12_51_groupi_g18131(csa_tree_add_12_51_groupi_n_3655 ,csa_tree_add_12_51_groupi_n_1791 ,csa_tree_add_12_51_groupi_n_1235);
  nor csa_tree_add_12_51_groupi_g18132(csa_tree_add_12_51_groupi_n_3654 ,csa_tree_add_12_51_groupi_n_1365 ,csa_tree_add_12_51_groupi_n_390);
  nor csa_tree_add_12_51_groupi_g18133(csa_tree_add_12_51_groupi_n_3653 ,csa_tree_add_12_51_groupi_n_1526 ,csa_tree_add_12_51_groupi_n_369);
  nor csa_tree_add_12_51_groupi_g18134(csa_tree_add_12_51_groupi_n_3652 ,csa_tree_add_12_51_groupi_n_1385 ,csa_tree_add_12_51_groupi_n_430);
  nor csa_tree_add_12_51_groupi_g18135(csa_tree_add_12_51_groupi_n_3651 ,csa_tree_add_12_51_groupi_n_1419 ,csa_tree_add_12_51_groupi_n_1310);
  nor csa_tree_add_12_51_groupi_g18136(csa_tree_add_12_51_groupi_n_3650 ,csa_tree_add_12_51_groupi_n_1080 ,csa_tree_add_12_51_groupi_n_397);
  nor csa_tree_add_12_51_groupi_g18137(csa_tree_add_12_51_groupi_n_3649 ,csa_tree_add_12_51_groupi_n_583 ,csa_tree_add_12_51_groupi_n_1149);
  nor csa_tree_add_12_51_groupi_g18138(csa_tree_add_12_51_groupi_n_3648 ,csa_tree_add_12_51_groupi_n_1502 ,csa_tree_add_12_51_groupi_n_204);
  nor csa_tree_add_12_51_groupi_g18139(csa_tree_add_12_51_groupi_n_3647 ,csa_tree_add_12_51_groupi_n_1440 ,csa_tree_add_12_51_groupi_n_1235);
  nor csa_tree_add_12_51_groupi_g18140(csa_tree_add_12_51_groupi_n_3646 ,csa_tree_add_12_51_groupi_n_1551 ,csa_tree_add_12_51_groupi_n_393);
  nor csa_tree_add_12_51_groupi_g18141(csa_tree_add_12_51_groupi_n_3645 ,csa_tree_add_12_51_groupi_n_1508 ,csa_tree_add_12_51_groupi_n_426);
  nor csa_tree_add_12_51_groupi_g18142(csa_tree_add_12_51_groupi_n_3644 ,csa_tree_add_12_51_groupi_n_1523 ,csa_tree_add_12_51_groupi_n_252);
  nor csa_tree_add_12_51_groupi_g18143(csa_tree_add_12_51_groupi_n_3643 ,csa_tree_add_12_51_groupi_n_523 ,csa_tree_add_12_51_groupi_n_1226);
  nor csa_tree_add_12_51_groupi_g18144(csa_tree_add_12_51_groupi_n_3642 ,csa_tree_add_12_51_groupi_n_1155 ,csa_tree_add_12_51_groupi_n_190);
  nor csa_tree_add_12_51_groupi_g18145(csa_tree_add_12_51_groupi_n_3641 ,csa_tree_add_12_51_groupi_n_1373 ,csa_tree_add_12_51_groupi_n_363);
  nor csa_tree_add_12_51_groupi_g18146(csa_tree_add_12_51_groupi_n_3640 ,csa_tree_add_12_51_groupi_n_1326 ,csa_tree_add_12_51_groupi_n_283);
  nor csa_tree_add_12_51_groupi_g18147(csa_tree_add_12_51_groupi_n_3639 ,csa_tree_add_12_51_groupi_n_1104 ,csa_tree_add_12_51_groupi_n_264);
  nor csa_tree_add_12_51_groupi_g18148(csa_tree_add_12_51_groupi_n_3638 ,csa_tree_add_12_51_groupi_n_493 ,csa_tree_add_12_51_groupi_n_1374);
  nor csa_tree_add_12_51_groupi_g18149(csa_tree_add_12_51_groupi_n_3637 ,csa_tree_add_12_51_groupi_n_1148 ,csa_tree_add_12_51_groupi_n_192);
  nor csa_tree_add_12_51_groupi_g18150(csa_tree_add_12_51_groupi_n_3636 ,csa_tree_add_12_51_groupi_n_1167 ,csa_tree_add_12_51_groupi_n_379);
  nor csa_tree_add_12_51_groupi_g18151(csa_tree_add_12_51_groupi_n_3635 ,csa_tree_add_12_51_groupi_n_1325 ,csa_tree_add_12_51_groupi_n_276);
  nor csa_tree_add_12_51_groupi_g18152(csa_tree_add_12_51_groupi_n_3634 ,csa_tree_add_12_51_groupi_n_547 ,csa_tree_add_12_51_groupi_n_1224);
  nor csa_tree_add_12_51_groupi_g18153(csa_tree_add_12_51_groupi_n_3633 ,csa_tree_add_12_51_groupi_n_1455 ,csa_tree_add_12_51_groupi_n_1175);
  nor csa_tree_add_12_51_groupi_g18154(csa_tree_add_12_51_groupi_n_3632 ,csa_tree_add_12_51_groupi_n_1410 ,csa_tree_add_12_51_groupi_n_1085);
  nor csa_tree_add_12_51_groupi_g18155(csa_tree_add_12_51_groupi_n_3631 ,csa_tree_add_12_51_groupi_n_1473 ,csa_tree_add_12_51_groupi_n_1139);
  nor csa_tree_add_12_51_groupi_g18156(csa_tree_add_12_51_groupi_n_3630 ,csa_tree_add_12_51_groupi_n_1458 ,csa_tree_add_12_51_groupi_n_963);
  nor csa_tree_add_12_51_groupi_g18157(csa_tree_add_12_51_groupi_n_3629 ,csa_tree_add_12_51_groupi_n_1311 ,csa_tree_add_12_51_groupi_n_403);
  nor csa_tree_add_12_51_groupi_g18158(csa_tree_add_12_51_groupi_n_3628 ,csa_tree_add_12_51_groupi_n_1404 ,csa_tree_add_12_51_groupi_n_1139);
  nor csa_tree_add_12_51_groupi_g18159(csa_tree_add_12_51_groupi_n_3627 ,csa_tree_add_12_51_groupi_n_616 ,csa_tree_add_12_51_groupi_n_1326);
  nor csa_tree_add_12_51_groupi_g18160(csa_tree_add_12_51_groupi_n_3626 ,csa_tree_add_12_51_groupi_n_1422 ,csa_tree_add_12_51_groupi_n_1248);
  nor csa_tree_add_12_51_groupi_g18161(csa_tree_add_12_51_groupi_n_3625 ,csa_tree_add_12_51_groupi_n_619 ,csa_tree_add_12_51_groupi_n_1148);
  nor csa_tree_add_12_51_groupi_g18162(csa_tree_add_12_51_groupi_n_3624 ,csa_tree_add_12_51_groupi_n_1431 ,csa_tree_add_12_51_groupi_n_879);
  nor csa_tree_add_12_51_groupi_g18163(csa_tree_add_12_51_groupi_n_3623 ,csa_tree_add_12_51_groupi_n_1524 ,csa_tree_add_12_51_groupi_n_349);
  nor csa_tree_add_12_51_groupi_g18164(csa_tree_add_12_51_groupi_n_3622 ,csa_tree_add_12_51_groupi_n_1434 ,csa_tree_add_12_51_groupi_n_1178);
  nor csa_tree_add_12_51_groupi_g18165(csa_tree_add_12_51_groupi_n_3621 ,csa_tree_add_12_51_groupi_n_586 ,csa_tree_add_12_51_groupi_n_1076);
  nor csa_tree_add_12_51_groupi_g18166(csa_tree_add_12_51_groupi_n_3620 ,csa_tree_add_12_51_groupi_n_682 ,csa_tree_add_12_51_groupi_n_1227);
  nor csa_tree_add_12_51_groupi_g18167(csa_tree_add_12_51_groupi_n_3619 ,csa_tree_add_12_51_groupi_n_574 ,csa_tree_add_12_51_groupi_n_1085);
  nor csa_tree_add_12_51_groupi_g18168(csa_tree_add_12_51_groupi_n_3618 ,csa_tree_add_12_51_groupi_n_1461 ,csa_tree_add_12_51_groupi_n_1172);
  nor csa_tree_add_12_51_groupi_g18169(csa_tree_add_12_51_groupi_n_3617 ,csa_tree_add_12_51_groupi_n_1427 ,csa_tree_add_12_51_groupi_n_1158);
  nor csa_tree_add_12_51_groupi_g18170(csa_tree_add_12_51_groupi_n_3616 ,csa_tree_add_12_51_groupi_n_580 ,csa_tree_add_12_51_groupi_n_1076);
  nor csa_tree_add_12_51_groupi_g18171(csa_tree_add_12_51_groupi_n_3615 ,csa_tree_add_12_51_groupi_n_1398 ,csa_tree_add_12_51_groupi_n_1091);
  nor csa_tree_add_12_51_groupi_g18172(csa_tree_add_12_51_groupi_n_3614 ,csa_tree_add_12_51_groupi_n_1137 ,csa_tree_add_12_51_groupi_n_466);
  nor csa_tree_add_12_51_groupi_g18173(csa_tree_add_12_51_groupi_n_3613 ,csa_tree_add_12_51_groupi_n_538 ,csa_tree_add_12_51_groupi_n_1145);
  nor csa_tree_add_12_51_groupi_g18174(csa_tree_add_12_51_groupi_n_3612 ,csa_tree_add_12_51_groupi_n_1086 ,csa_tree_add_12_51_groupi_n_346);
  nor csa_tree_add_12_51_groupi_g18175(csa_tree_add_12_51_groupi_n_3611 ,csa_tree_add_12_51_groupi_n_1551 ,csa_tree_add_12_51_groupi_n_375);
  nor csa_tree_add_12_51_groupi_g18176(csa_tree_add_12_51_groupi_n_3610 ,csa_tree_add_12_51_groupi_n_577 ,csa_tree_add_12_51_groupi_n_1077);
  nor csa_tree_add_12_51_groupi_g18177(csa_tree_add_12_51_groupi_n_3609 ,csa_tree_add_12_51_groupi_n_1751 ,csa_tree_add_12_51_groupi_n_1319);
  nor csa_tree_add_12_51_groupi_g18178(csa_tree_add_12_51_groupi_n_3608 ,csa_tree_add_12_51_groupi_n_484 ,csa_tree_add_12_51_groupi_n_926);
  nor csa_tree_add_12_51_groupi_g18179(csa_tree_add_12_51_groupi_n_3607 ,csa_tree_add_12_51_groupi_n_1550 ,csa_tree_add_12_51_groupi_n_478);
  nor csa_tree_add_12_51_groupi_g18180(csa_tree_add_12_51_groupi_n_3606 ,csa_tree_add_12_51_groupi_n_1143 ,csa_tree_add_12_51_groupi_n_445);
  nor csa_tree_add_12_51_groupi_g18181(csa_tree_add_12_51_groupi_n_3605 ,csa_tree_add_12_51_groupi_n_529 ,csa_tree_add_12_51_groupi_n_1140);
  nor csa_tree_add_12_51_groupi_g18182(csa_tree_add_12_51_groupi_n_3604 ,csa_tree_add_12_51_groupi_n_1269 ,csa_tree_add_12_51_groupi_n_1091);
  nor csa_tree_add_12_51_groupi_g18183(csa_tree_add_12_51_groupi_n_3603 ,csa_tree_add_12_51_groupi_n_1413 ,csa_tree_add_12_51_groupi_n_962);
  nor csa_tree_add_12_51_groupi_g18184(csa_tree_add_12_51_groupi_n_3602 ,csa_tree_add_12_51_groupi_n_550 ,csa_tree_add_12_51_groupi_n_1155);
  nor csa_tree_add_12_51_groupi_g18185(csa_tree_add_12_51_groupi_n_3601 ,csa_tree_add_12_51_groupi_n_1416 ,csa_tree_add_12_51_groupi_n_927);
  nor csa_tree_add_12_51_groupi_g18186(csa_tree_add_12_51_groupi_n_3600 ,csa_tree_add_12_51_groupi_n_568 ,csa_tree_add_12_51_groupi_n_1176);
  nor csa_tree_add_12_51_groupi_g18187(csa_tree_add_12_51_groupi_n_3599 ,csa_tree_add_12_51_groupi_n_649 ,csa_tree_add_12_51_groupi_n_887);
  nor csa_tree_add_12_51_groupi_g18188(csa_tree_add_12_51_groupi_n_3598 ,csa_tree_add_12_51_groupi_n_667 ,csa_tree_add_12_51_groupi_n_1146);
  nor csa_tree_add_12_51_groupi_g18189(csa_tree_add_12_51_groupi_n_3597 ,csa_tree_add_12_51_groupi_n_571 ,csa_tree_add_12_51_groupi_n_888);
  nor csa_tree_add_12_51_groupi_g18190(csa_tree_add_12_51_groupi_n_3596 ,csa_tree_add_12_51_groupi_n_661 ,csa_tree_add_12_51_groupi_n_1173);
  nor csa_tree_add_12_51_groupi_g18191(csa_tree_add_12_51_groupi_n_3595 ,csa_tree_add_12_51_groupi_n_637 ,csa_tree_add_12_51_groupi_n_1092);
  nor csa_tree_add_12_51_groupi_g18192(csa_tree_add_12_51_groupi_n_3594 ,csa_tree_add_12_51_groupi_n_679 ,csa_tree_add_12_51_groupi_n_1172);
  nor csa_tree_add_12_51_groupi_g18193(csa_tree_add_12_51_groupi_n_3593 ,csa_tree_add_12_51_groupi_n_634 ,csa_tree_add_12_51_groupi_n_878);
  nor csa_tree_add_12_51_groupi_g18194(csa_tree_add_12_51_groupi_n_3592 ,csa_tree_add_12_51_groupi_n_625 ,csa_tree_add_12_51_groupi_n_1086);
  nor csa_tree_add_12_51_groupi_g18195(csa_tree_add_12_51_groupi_n_3591 ,csa_tree_add_12_51_groupi_n_1569 ,csa_tree_add_12_51_groupi_n_1142);
  nor csa_tree_add_12_51_groupi_g18196(csa_tree_add_12_51_groupi_n_3590 ,csa_tree_add_12_51_groupi_n_607 ,csa_tree_add_12_51_groupi_n_869);
  nor csa_tree_add_12_51_groupi_g18197(csa_tree_add_12_51_groupi_n_3589 ,csa_tree_add_12_51_groupi_n_610 ,csa_tree_add_12_51_groupi_n_1154);
  nor csa_tree_add_12_51_groupi_g18198(csa_tree_add_12_51_groupi_n_3588 ,csa_tree_add_12_51_groupi_n_1709 ,csa_tree_add_12_51_groupi_n_956);
  nor csa_tree_add_12_51_groupi_g18199(csa_tree_add_12_51_groupi_n_3587 ,csa_tree_add_12_51_groupi_n_559 ,csa_tree_add_12_51_groupi_n_1247);
  nor csa_tree_add_12_51_groupi_g18200(csa_tree_add_12_51_groupi_n_3586 ,csa_tree_add_12_51_groupi_n_595 ,csa_tree_add_12_51_groupi_n_888);
  nor csa_tree_add_12_51_groupi_g18201(csa_tree_add_12_51_groupi_n_3585 ,csa_tree_add_12_51_groupi_n_652 ,csa_tree_add_12_51_groupi_n_872);
  nor csa_tree_add_12_51_groupi_g18202(csa_tree_add_12_51_groupi_n_3584 ,csa_tree_add_12_51_groupi_n_673 ,csa_tree_add_12_51_groupi_n_1136);
  nor csa_tree_add_12_51_groupi_g18203(csa_tree_add_12_51_groupi_n_3583 ,csa_tree_add_12_51_groupi_n_541 ,csa_tree_add_12_51_groupi_n_1103);
  nor csa_tree_add_12_51_groupi_g18204(csa_tree_add_12_51_groupi_n_3582 ,csa_tree_add_12_51_groupi_n_1784 ,csa_tree_add_12_51_groupi_n_957);
  nor csa_tree_add_12_51_groupi_g18205(csa_tree_add_12_51_groupi_n_3581 ,csa_tree_add_12_51_groupi_n_1605 ,csa_tree_add_12_51_groupi_n_1037);
  nor csa_tree_add_12_51_groupi_g18206(csa_tree_add_12_51_groupi_n_3580 ,csa_tree_add_12_51_groupi_n_1593 ,csa_tree_add_12_51_groupi_n_1040);
  nor csa_tree_add_12_51_groupi_g18207(csa_tree_add_12_51_groupi_n_3579 ,csa_tree_add_12_51_groupi_n_1584 ,csa_tree_add_12_51_groupi_n_169);
  nor csa_tree_add_12_51_groupi_g18208(csa_tree_add_12_51_groupi_n_3578 ,csa_tree_add_12_51_groupi_n_1617 ,csa_tree_add_12_51_groupi_n_1037);
  nor csa_tree_add_12_51_groupi_g18209(csa_tree_add_12_51_groupi_n_3577 ,csa_tree_add_12_51_groupi_n_1599 ,csa_tree_add_12_51_groupi_n_1038);
  nor csa_tree_add_12_51_groupi_g18210(csa_tree_add_12_51_groupi_n_3576 ,csa_tree_add_12_51_groupi_n_1656 ,csa_tree_add_12_51_groupi_n_1041);
  nor csa_tree_add_12_51_groupi_g18211(csa_tree_add_12_51_groupi_n_3575 ,csa_tree_add_12_51_groupi_n_1641 ,csa_tree_add_12_51_groupi_n_894);
  nor csa_tree_add_12_51_groupi_g18212(csa_tree_add_12_51_groupi_n_3574 ,csa_tree_add_12_51_groupi_n_1629 ,csa_tree_add_12_51_groupi_n_893);
  nor csa_tree_add_12_51_groupi_g18213(csa_tree_add_12_51_groupi_n_3573 ,csa_tree_add_12_51_groupi_n_1623 ,csa_tree_add_12_51_groupi_n_1038);
  nor csa_tree_add_12_51_groupi_g18214(csa_tree_add_12_51_groupi_n_3572 ,csa_tree_add_12_51_groupi_n_1611 ,csa_tree_add_12_51_groupi_n_893);
  nor csa_tree_add_12_51_groupi_g18215(csa_tree_add_12_51_groupi_n_3571 ,csa_tree_add_12_51_groupi_n_1647 ,csa_tree_add_12_51_groupi_n_1041);
  nor csa_tree_add_12_51_groupi_g18216(csa_tree_add_12_51_groupi_n_3570 ,csa_tree_add_12_51_groupi_n_1635 ,csa_tree_add_12_51_groupi_n_1040);
  nor csa_tree_add_12_51_groupi_g18217(csa_tree_add_12_51_groupi_n_3569 ,csa_tree_add_12_51_groupi_n_1665 ,csa_tree_add_12_51_groupi_n_2007);
  nor csa_tree_add_12_51_groupi_g18218(csa_tree_add_12_51_groupi_n_3568 ,csa_tree_add_12_51_groupi_n_1680 ,csa_tree_add_12_51_groupi_n_894);
  nor csa_tree_add_12_51_groupi_g18219(csa_tree_add_12_51_groupi_n_3567 ,csa_tree_add_12_51_groupi_n_1587 ,csa_tree_add_12_51_groupi_n_169);
  xnor csa_tree_add_12_51_groupi_g18220(csa_tree_add_12_51_groupi_n_3566 ,csa_tree_add_12_51_groupi_n_2468 ,csa_tree_add_12_51_groupi_n_2949);
  xnor csa_tree_add_12_51_groupi_g18221(csa_tree_add_12_51_groupi_n_3565 ,csa_tree_add_12_51_groupi_n_2961 ,csa_tree_add_12_51_groupi_n_2758);
  xnor csa_tree_add_12_51_groupi_g18222(csa_tree_add_12_51_groupi_n_3564 ,csa_tree_add_12_51_groupi_n_2956 ,in5[4]);
  xnor csa_tree_add_12_51_groupi_g18223(csa_tree_add_12_51_groupi_n_3563 ,csa_tree_add_12_51_groupi_n_2869 ,csa_tree_add_12_51_groupi_n_2868);
  xnor csa_tree_add_12_51_groupi_g18224(csa_tree_add_12_51_groupi_n_3562 ,csa_tree_add_12_51_groupi_n_2954 ,in5[10]);
  xnor csa_tree_add_12_51_groupi_g18225(csa_tree_add_12_51_groupi_n_3561 ,csa_tree_add_12_51_groupi_n_2953 ,in5[13]);
  xnor csa_tree_add_12_51_groupi_g18226(csa_tree_add_12_51_groupi_n_3560 ,csa_tree_add_12_51_groupi_n_2957 ,in5[7]);
  xnor csa_tree_add_12_51_groupi_g18227(csa_tree_add_12_51_groupi_n_3559 ,csa_tree_add_12_51_groupi_n_2952 ,in5[1]);
  xnor csa_tree_add_12_51_groupi_g18228(csa_tree_add_12_51_groupi_n_3765 ,csa_tree_add_12_51_groupi_n_2870 ,in5[15]);
  xnor csa_tree_add_12_51_groupi_g18229(csa_tree_add_12_51_groupi_n_3764 ,csa_tree_add_12_51_groupi_n_2960 ,csa_tree_add_12_51_groupi_n_2561);
  not csa_tree_add_12_51_groupi_g18230(csa_tree_add_12_51_groupi_n_3555 ,csa_tree_add_12_51_groupi_n_3554);
  not csa_tree_add_12_51_groupi_g18231(csa_tree_add_12_51_groupi_n_3546 ,csa_tree_add_12_51_groupi_n_3547);
  not csa_tree_add_12_51_groupi_g18232(csa_tree_add_12_51_groupi_n_3543 ,csa_tree_add_12_51_groupi_n_3544);
  not csa_tree_add_12_51_groupi_g18233(csa_tree_add_12_51_groupi_n_3541 ,csa_tree_add_12_51_groupi_n_3542);
  not csa_tree_add_12_51_groupi_g18234(csa_tree_add_12_51_groupi_n_3538 ,csa_tree_add_12_51_groupi_n_3539);
  not csa_tree_add_12_51_groupi_g18235(csa_tree_add_12_51_groupi_n_3535 ,csa_tree_add_12_51_groupi_n_3536);
  not csa_tree_add_12_51_groupi_g18236(csa_tree_add_12_51_groupi_n_3533 ,csa_tree_add_12_51_groupi_n_3534);
  not csa_tree_add_12_51_groupi_g18237(csa_tree_add_12_51_groupi_n_3531 ,csa_tree_add_12_51_groupi_n_3532);
  not csa_tree_add_12_51_groupi_g18238(csa_tree_add_12_51_groupi_n_3526 ,csa_tree_add_12_51_groupi_n_3527);
  not csa_tree_add_12_51_groupi_g18239(csa_tree_add_12_51_groupi_n_3523 ,csa_tree_add_12_51_groupi_n_3524);
  not csa_tree_add_12_51_groupi_g18240(csa_tree_add_12_51_groupi_n_3519 ,csa_tree_add_12_51_groupi_n_3520);
  not csa_tree_add_12_51_groupi_g18241(csa_tree_add_12_51_groupi_n_3515 ,csa_tree_add_12_51_groupi_n_3516);
  not csa_tree_add_12_51_groupi_g18242(csa_tree_add_12_51_groupi_n_3514 ,csa_tree_add_12_51_groupi_n_3513);
  not csa_tree_add_12_51_groupi_g18243(csa_tree_add_12_51_groupi_n_3512 ,csa_tree_add_12_51_groupi_n_3511);
  not csa_tree_add_12_51_groupi_g18244(csa_tree_add_12_51_groupi_n_3509 ,csa_tree_add_12_51_groupi_n_3510);
  nor csa_tree_add_12_51_groupi_g18245(csa_tree_add_12_51_groupi_n_3496 ,csa_tree_add_12_51_groupi_n_1799 ,csa_tree_add_12_51_groupi_n_1488);
  and csa_tree_add_12_51_groupi_g18246(csa_tree_add_12_51_groupi_n_3495 ,in5[4] ,csa_tree_add_12_51_groupi_n_2956);
  and csa_tree_add_12_51_groupi_g18247(csa_tree_add_12_51_groupi_n_3494 ,csa_tree_add_12_51_groupi_n_2468 ,csa_tree_add_12_51_groupi_n_2161);
  or csa_tree_add_12_51_groupi_g18248(csa_tree_add_12_51_groupi_n_3493 ,in5[13] ,csa_tree_add_12_51_groupi_n_2953);
  and csa_tree_add_12_51_groupi_g18249(csa_tree_add_12_51_groupi_n_3492 ,in5[13] ,csa_tree_add_12_51_groupi_n_2953);
  and csa_tree_add_12_51_groupi_g18250(csa_tree_add_12_51_groupi_n_3491 ,in5[7] ,csa_tree_add_12_51_groupi_n_2957);
  or csa_tree_add_12_51_groupi_g18251(csa_tree_add_12_51_groupi_n_3490 ,in5[1] ,csa_tree_add_12_51_groupi_n_2952);
  or csa_tree_add_12_51_groupi_g18252(csa_tree_add_12_51_groupi_n_3489 ,in5[4] ,csa_tree_add_12_51_groupi_n_2956);
  or csa_tree_add_12_51_groupi_g18253(csa_tree_add_12_51_groupi_n_3488 ,csa_tree_add_12_51_groupi_n_2468 ,csa_tree_add_12_51_groupi_n_2949);
  and csa_tree_add_12_51_groupi_g18254(csa_tree_add_12_51_groupi_n_3487 ,in5[1] ,csa_tree_add_12_51_groupi_n_2952);
  or csa_tree_add_12_51_groupi_g18255(csa_tree_add_12_51_groupi_n_3486 ,in5[10] ,csa_tree_add_12_51_groupi_n_2954);
  or csa_tree_add_12_51_groupi_g18256(csa_tree_add_12_51_groupi_n_3485 ,in5[7] ,csa_tree_add_12_51_groupi_n_2957);
  and csa_tree_add_12_51_groupi_g18257(csa_tree_add_12_51_groupi_n_3484 ,in5[10] ,csa_tree_add_12_51_groupi_n_2954);
  or csa_tree_add_12_51_groupi_g18258(csa_tree_add_12_51_groupi_n_3483 ,csa_tree_add_12_51_groupi_n_2670 ,csa_tree_add_12_51_groupi_n_2897);
  or csa_tree_add_12_51_groupi_g18259(csa_tree_add_12_51_groupi_n_3482 ,csa_tree_add_12_51_groupi_n_2666 ,csa_tree_add_12_51_groupi_n_2889);
  or csa_tree_add_12_51_groupi_g18260(csa_tree_add_12_51_groupi_n_3481 ,csa_tree_add_12_51_groupi_n_2669 ,csa_tree_add_12_51_groupi_n_2902);
  or csa_tree_add_12_51_groupi_g18261(csa_tree_add_12_51_groupi_n_3480 ,csa_tree_add_12_51_groupi_n_2442 ,csa_tree_add_12_51_groupi_n_2960);
  or csa_tree_add_12_51_groupi_g18262(csa_tree_add_12_51_groupi_n_3479 ,csa_tree_add_12_51_groupi_n_2664 ,csa_tree_add_12_51_groupi_n_2864);
  or csa_tree_add_12_51_groupi_g18263(csa_tree_add_12_51_groupi_n_3478 ,csa_tree_add_12_51_groupi_n_2602 ,csa_tree_add_12_51_groupi_n_2885);
  or csa_tree_add_12_51_groupi_g18264(csa_tree_add_12_51_groupi_n_3477 ,csa_tree_add_12_51_groupi_n_2691 ,csa_tree_add_12_51_groupi_n_2882);
  or csa_tree_add_12_51_groupi_g18265(csa_tree_add_12_51_groupi_n_3476 ,csa_tree_add_12_51_groupi_n_2668 ,csa_tree_add_12_51_groupi_n_2830);
  or csa_tree_add_12_51_groupi_g18266(csa_tree_add_12_51_groupi_n_3475 ,csa_tree_add_12_51_groupi_n_2672 ,csa_tree_add_12_51_groupi_n_2883);
  or csa_tree_add_12_51_groupi_g18267(csa_tree_add_12_51_groupi_n_3474 ,csa_tree_add_12_51_groupi_n_2599 ,csa_tree_add_12_51_groupi_n_2905);
  or csa_tree_add_12_51_groupi_g18268(csa_tree_add_12_51_groupi_n_3473 ,csa_tree_add_12_51_groupi_n_2618 ,csa_tree_add_12_51_groupi_n_2831);
  or csa_tree_add_12_51_groupi_g18269(csa_tree_add_12_51_groupi_n_3472 ,csa_tree_add_12_51_groupi_n_2580 ,csa_tree_add_12_51_groupi_n_2861);
  or csa_tree_add_12_51_groupi_g18270(csa_tree_add_12_51_groupi_n_3471 ,csa_tree_add_12_51_groupi_n_2593 ,csa_tree_add_12_51_groupi_n_2859);
  or csa_tree_add_12_51_groupi_g18271(csa_tree_add_12_51_groupi_n_3470 ,csa_tree_add_12_51_groupi_n_2577 ,csa_tree_add_12_51_groupi_n_2856);
  or csa_tree_add_12_51_groupi_g18272(csa_tree_add_12_51_groupi_n_3469 ,csa_tree_add_12_51_groupi_n_2710 ,csa_tree_add_12_51_groupi_n_2834);
  or csa_tree_add_12_51_groupi_g18273(csa_tree_add_12_51_groupi_n_3468 ,csa_tree_add_12_51_groupi_n_2687 ,csa_tree_add_12_51_groupi_n_2839);
  or csa_tree_add_12_51_groupi_g18274(csa_tree_add_12_51_groupi_n_3467 ,csa_tree_add_12_51_groupi_n_2589 ,csa_tree_add_12_51_groupi_n_2835);
  or csa_tree_add_12_51_groupi_g18275(csa_tree_add_12_51_groupi_n_3466 ,csa_tree_add_12_51_groupi_n_2605 ,csa_tree_add_12_51_groupi_n_2866);
  or csa_tree_add_12_51_groupi_g18276(csa_tree_add_12_51_groupi_n_3465 ,csa_tree_add_12_51_groupi_n_2607 ,csa_tree_add_12_51_groupi_n_2840);
  or csa_tree_add_12_51_groupi_g18277(csa_tree_add_12_51_groupi_n_3464 ,csa_tree_add_12_51_groupi_n_2606 ,csa_tree_add_12_51_groupi_n_2852);
  or csa_tree_add_12_51_groupi_g18278(csa_tree_add_12_51_groupi_n_3463 ,csa_tree_add_12_51_groupi_n_2611 ,csa_tree_add_12_51_groupi_n_2833);
  or csa_tree_add_12_51_groupi_g18279(csa_tree_add_12_51_groupi_n_3462 ,csa_tree_add_12_51_groupi_n_2601 ,csa_tree_add_12_51_groupi_n_2836);
  or csa_tree_add_12_51_groupi_g18280(csa_tree_add_12_51_groupi_n_3461 ,csa_tree_add_12_51_groupi_n_2636 ,csa_tree_add_12_51_groupi_n_2860);
  or csa_tree_add_12_51_groupi_g18281(csa_tree_add_12_51_groupi_n_3460 ,csa_tree_add_12_51_groupi_n_2600 ,csa_tree_add_12_51_groupi_n_2858);
  or csa_tree_add_12_51_groupi_g18282(csa_tree_add_12_51_groupi_n_3459 ,csa_tree_add_12_51_groupi_n_2634 ,csa_tree_add_12_51_groupi_n_2847);
  or csa_tree_add_12_51_groupi_g18283(csa_tree_add_12_51_groupi_n_3458 ,csa_tree_add_12_51_groupi_n_2734 ,csa_tree_add_12_51_groupi_n_2841);
  or csa_tree_add_12_51_groupi_g18284(csa_tree_add_12_51_groupi_n_3457 ,csa_tree_add_12_51_groupi_n_2635 ,csa_tree_add_12_51_groupi_n_2865);
  or csa_tree_add_12_51_groupi_g18285(csa_tree_add_12_51_groupi_n_3456 ,csa_tree_add_12_51_groupi_n_2613 ,csa_tree_add_12_51_groupi_n_2845);
  or csa_tree_add_12_51_groupi_g18286(csa_tree_add_12_51_groupi_n_3455 ,csa_tree_add_12_51_groupi_n_2709 ,csa_tree_add_12_51_groupi_n_2849);
  or csa_tree_add_12_51_groupi_g18287(csa_tree_add_12_51_groupi_n_3454 ,csa_tree_add_12_51_groupi_n_2586 ,csa_tree_add_12_51_groupi_n_2844);
  or csa_tree_add_12_51_groupi_g18288(csa_tree_add_12_51_groupi_n_3453 ,csa_tree_add_12_51_groupi_n_2596 ,csa_tree_add_12_51_groupi_n_2863);
  or csa_tree_add_12_51_groupi_g18289(csa_tree_add_12_51_groupi_n_3452 ,csa_tree_add_12_51_groupi_n_2612 ,csa_tree_add_12_51_groupi_n_2857);
  or csa_tree_add_12_51_groupi_g18290(csa_tree_add_12_51_groupi_n_3451 ,csa_tree_add_12_51_groupi_n_2592 ,csa_tree_add_12_51_groupi_n_2862);
  or csa_tree_add_12_51_groupi_g18291(csa_tree_add_12_51_groupi_n_3450 ,csa_tree_add_12_51_groupi_n_2625 ,csa_tree_add_12_51_groupi_n_2850);
  or csa_tree_add_12_51_groupi_g18292(csa_tree_add_12_51_groupi_n_3449 ,csa_tree_add_12_51_groupi_n_2621 ,csa_tree_add_12_51_groupi_n_2837);
  or csa_tree_add_12_51_groupi_g18293(csa_tree_add_12_51_groupi_n_3448 ,csa_tree_add_12_51_groupi_n_2579 ,csa_tree_add_12_51_groupi_n_2838);
  or csa_tree_add_12_51_groupi_g18294(csa_tree_add_12_51_groupi_n_3447 ,csa_tree_add_12_51_groupi_n_2617 ,csa_tree_add_12_51_groupi_n_2842);
  or csa_tree_add_12_51_groupi_g18295(csa_tree_add_12_51_groupi_n_3446 ,csa_tree_add_12_51_groupi_n_2743 ,csa_tree_add_12_51_groupi_n_2853);
  or csa_tree_add_12_51_groupi_g18296(csa_tree_add_12_51_groupi_n_3445 ,csa_tree_add_12_51_groupi_n_2624 ,csa_tree_add_12_51_groupi_n_2823);
  or csa_tree_add_12_51_groupi_g18297(csa_tree_add_12_51_groupi_n_3444 ,csa_tree_add_12_51_groupi_n_2594 ,csa_tree_add_12_51_groupi_n_2855);
  or csa_tree_add_12_51_groupi_g18298(csa_tree_add_12_51_groupi_n_3443 ,csa_tree_add_12_51_groupi_n_2694 ,csa_tree_add_12_51_groupi_n_2851);
  or csa_tree_add_12_51_groupi_g18299(csa_tree_add_12_51_groupi_n_3442 ,csa_tree_add_12_51_groupi_n_2603 ,csa_tree_add_12_51_groupi_n_2854);
  or csa_tree_add_12_51_groupi_g18300(csa_tree_add_12_51_groupi_n_3441 ,csa_tree_add_12_51_groupi_n_2604 ,csa_tree_add_12_51_groupi_n_2848);
  or csa_tree_add_12_51_groupi_g18301(csa_tree_add_12_51_groupi_n_3440 ,csa_tree_add_12_51_groupi_n_2690 ,csa_tree_add_12_51_groupi_n_2846);
  or csa_tree_add_12_51_groupi_g18302(csa_tree_add_12_51_groupi_n_3439 ,csa_tree_add_12_51_groupi_n_2622 ,csa_tree_add_12_51_groupi_n_2832);
  or csa_tree_add_12_51_groupi_g18303(csa_tree_add_12_51_groupi_n_3438 ,csa_tree_add_12_51_groupi_n_2629 ,csa_tree_add_12_51_groupi_n_2843);
  and csa_tree_add_12_51_groupi_g18304(csa_tree_add_12_51_groupi_n_3437 ,csa_tree_add_12_51_groupi_n_2869 ,csa_tree_add_12_51_groupi_n_2868);
  nor csa_tree_add_12_51_groupi_g18305(csa_tree_add_12_51_groupi_n_3436 ,csa_tree_add_12_51_groupi_n_2869 ,csa_tree_add_12_51_groupi_n_2868);
  or csa_tree_add_12_51_groupi_g18306(csa_tree_add_12_51_groupi_n_3435 ,csa_tree_add_12_51_groupi_n_2961 ,csa_tree_add_12_51_groupi_n_2829);
  nor csa_tree_add_12_51_groupi_g18307(csa_tree_add_12_51_groupi_n_3434 ,csa_tree_add_12_51_groupi_n_1730 ,csa_tree_add_12_51_groupi_n_1341);
  nor csa_tree_add_12_51_groupi_g18308(csa_tree_add_12_51_groupi_n_3433 ,csa_tree_add_12_51_groupi_n_1574 ,csa_tree_add_12_51_groupi_n_262);
  nor csa_tree_add_12_51_groupi_g18309(csa_tree_add_12_51_groupi_n_3432 ,csa_tree_add_12_51_groupi_n_1754 ,csa_tree_add_12_51_groupi_n_1119);
  nor csa_tree_add_12_51_groupi_g18310(csa_tree_add_12_51_groupi_n_3431 ,csa_tree_add_12_51_groupi_n_1685 ,csa_tree_add_12_51_groupi_n_199);
  nor csa_tree_add_12_51_groupi_g18311(csa_tree_add_12_51_groupi_n_3430 ,csa_tree_add_12_51_groupi_n_1775 ,csa_tree_add_12_51_groupi_n_1497);
  nor csa_tree_add_12_51_groupi_g18312(csa_tree_add_12_51_groupi_n_3429 ,csa_tree_add_12_51_groupi_n_1739 ,csa_tree_add_12_51_groupi_n_1302);
  nor csa_tree_add_12_51_groupi_g18313(csa_tree_add_12_51_groupi_n_3428 ,csa_tree_add_12_51_groupi_n_1721 ,csa_tree_add_12_51_groupi_n_1520);
  nor csa_tree_add_12_51_groupi_g18314(csa_tree_add_12_51_groupi_n_3427 ,csa_tree_add_12_51_groupi_n_1118 ,csa_tree_add_12_51_groupi_n_268);
  nor csa_tree_add_12_51_groupi_g18315(csa_tree_add_12_51_groupi_n_3426 ,csa_tree_add_12_51_groupi_n_646 ,csa_tree_add_12_51_groupi_n_1301);
  nor csa_tree_add_12_51_groupi_g18316(csa_tree_add_12_51_groupi_n_3425 ,csa_tree_add_12_51_groupi_n_1305 ,csa_tree_add_12_51_groupi_n_292);
  nor csa_tree_add_12_51_groupi_g18317(csa_tree_add_12_51_groupi_n_3424 ,csa_tree_add_12_51_groupi_n_1718 ,csa_tree_add_12_51_groupi_n_1340);
  nor csa_tree_add_12_51_groupi_g18318(csa_tree_add_12_51_groupi_n_3423 ,csa_tree_add_12_51_groupi_n_1805 ,csa_tree_add_12_51_groupi_n_1542);
  nor csa_tree_add_12_51_groupi_g18319(csa_tree_add_12_51_groupi_n_3422 ,csa_tree_add_12_51_groupi_n_1134 ,csa_tree_add_12_51_groupi_n_436);
  nor csa_tree_add_12_51_groupi_g18320(csa_tree_add_12_51_groupi_n_3421 ,csa_tree_add_12_51_groupi_n_1674 ,csa_tree_add_12_51_groupi_n_259);
  nor csa_tree_add_12_51_groupi_g18321(csa_tree_add_12_51_groupi_n_3420 ,csa_tree_add_12_51_groupi_n_1095 ,csa_tree_add_12_51_groupi_n_309);
  nor csa_tree_add_12_51_groupi_g18322(csa_tree_add_12_51_groupi_n_3419 ,csa_tree_add_12_51_groupi_n_1536 ,csa_tree_add_12_51_groupi_n_421);
  nor csa_tree_add_12_51_groupi_g18323(csa_tree_add_12_51_groupi_n_3418 ,csa_tree_add_12_51_groupi_n_1194 ,csa_tree_add_12_51_groupi_n_220);
  nor csa_tree_add_12_51_groupi_g18324(csa_tree_add_12_51_groupi_n_3417 ,csa_tree_add_12_51_groupi_n_1131 ,csa_tree_add_12_51_groupi_n_337);
  nor csa_tree_add_12_51_groupi_g18325(csa_tree_add_12_51_groupi_n_3416 ,csa_tree_add_12_51_groupi_n_864 ,csa_tree_add_12_51_groupi_n_217);
  nor csa_tree_add_12_51_groupi_g18326(csa_tree_add_12_51_groupi_n_3415 ,csa_tree_add_12_51_groupi_n_1668 ,csa_tree_add_12_51_groupi_n_1265);
  nor csa_tree_add_12_51_groupi_g18327(csa_tree_add_12_51_groupi_n_3414 ,csa_tree_add_12_51_groupi_n_481 ,csa_tree_add_12_51_groupi_n_1338);
  nor csa_tree_add_12_51_groupi_g18328(csa_tree_add_12_51_groupi_n_3413 ,csa_tree_add_12_51_groupi_n_504 ,csa_tree_add_12_51_groupi_n_915);
  nor csa_tree_add_12_51_groupi_g18329(csa_tree_add_12_51_groupi_n_3412 ,csa_tree_add_12_51_groupi_n_694 ,csa_tree_add_12_51_groupi_n_1197);
  nor csa_tree_add_12_51_groupi_g18330(csa_tree_add_12_51_groupi_n_3411 ,csa_tree_add_12_51_groupi_n_1554 ,csa_tree_add_12_51_groupi_n_307);
  nor csa_tree_add_12_51_groupi_g18331(csa_tree_add_12_51_groupi_n_3410 ,csa_tree_add_12_51_groupi_n_1395 ,csa_tree_add_12_51_groupi_n_322);
  nor csa_tree_add_12_51_groupi_g18332(csa_tree_add_12_51_groupi_n_3409 ,csa_tree_add_12_51_groupi_n_526 ,csa_tree_add_12_51_groupi_n_1212);
  nor csa_tree_add_12_51_groupi_g18333(csa_tree_add_12_51_groupi_n_3408 ,csa_tree_add_12_51_groupi_n_1572 ,csa_tree_add_12_51_groupi_n_858);
  nor csa_tree_add_12_51_groupi_g18334(csa_tree_add_12_51_groupi_n_3407 ,csa_tree_add_12_51_groupi_n_1803 ,csa_tree_add_12_51_groupi_n_1206);
  nor csa_tree_add_12_51_groupi_g18335(csa_tree_add_12_51_groupi_n_3406 ,csa_tree_add_12_51_groupi_n_664 ,csa_tree_add_12_51_groupi_n_1124);
  nor csa_tree_add_12_51_groupi_g18336(csa_tree_add_12_51_groupi_n_3405 ,csa_tree_add_12_51_groupi_n_1293 ,csa_tree_add_12_51_groupi_n_304);
  nor csa_tree_add_12_51_groupi_g18337(csa_tree_add_12_51_groupi_n_3404 ,csa_tree_add_12_51_groupi_n_1392 ,csa_tree_add_12_51_groupi_n_232);
  nor csa_tree_add_12_51_groupi_g18338(csa_tree_add_12_51_groupi_n_3403 ,csa_tree_add_12_51_groupi_n_1341 ,csa_tree_add_12_51_groupi_n_337);
  nor csa_tree_add_12_51_groupi_g18339(csa_tree_add_12_51_groupi_n_3402 ,csa_tree_add_12_51_groupi_n_1575 ,csa_tree_add_12_51_groupi_n_217);
  nor csa_tree_add_12_51_groupi_g18340(csa_tree_add_12_51_groupi_n_3401 ,csa_tree_add_12_51_groupi_n_1686 ,csa_tree_add_12_51_groupi_n_208);
  nor csa_tree_add_12_51_groupi_g18341(csa_tree_add_12_51_groupi_n_3400 ,csa_tree_add_12_51_groupi_n_1521 ,csa_tree_add_12_51_groupi_n_256);
  nor csa_tree_add_12_51_groupi_g18342(csa_tree_add_12_51_groupi_n_3399 ,csa_tree_add_12_51_groupi_n_1539 ,csa_tree_add_12_51_groupi_n_313);
  nor csa_tree_add_12_51_groupi_g18343(csa_tree_add_12_51_groupi_n_3398 ,csa_tree_add_12_51_groupi_n_1560 ,csa_tree_add_12_51_groupi_n_424);
  nor csa_tree_add_12_51_groupi_g18344(csa_tree_add_12_51_groupi_n_3397 ,csa_tree_add_12_51_groupi_n_604 ,csa_tree_add_12_51_groupi_n_1064);
  nor csa_tree_add_12_51_groupi_g18345(csa_tree_add_12_51_groupi_n_3396 ,csa_tree_add_12_51_groupi_n_939 ,csa_tree_add_12_51_groupi_n_427);
  nor csa_tree_add_12_51_groupi_g18346(csa_tree_add_12_51_groupi_n_3395 ,csa_tree_add_12_51_groupi_n_1563 ,csa_tree_add_12_51_groupi_n_406);
  nor csa_tree_add_12_51_groupi_g18347(csa_tree_add_12_51_groupi_n_3394 ,csa_tree_add_12_51_groupi_n_918 ,csa_tree_add_12_51_groupi_n_379);
  nor csa_tree_add_12_51_groupi_g18348(csa_tree_add_12_51_groupi_n_3393 ,csa_tree_add_12_51_groupi_n_1541 ,csa_tree_add_12_51_groupi_n_355);
  nor csa_tree_add_12_51_groupi_g18349(csa_tree_add_12_51_groupi_n_3392 ,csa_tree_add_12_51_groupi_n_1190 ,csa_tree_add_12_51_groupi_n_286);
  nor csa_tree_add_12_51_groupi_g18350(csa_tree_add_12_51_groupi_n_3391 ,csa_tree_add_12_51_groupi_n_1337 ,csa_tree_add_12_51_groupi_n_349);
  nor csa_tree_add_12_51_groupi_g18351(csa_tree_add_12_51_groupi_n_3390 ,csa_tree_add_12_51_groupi_n_1667 ,csa_tree_add_12_51_groupi_n_250);
  nor csa_tree_add_12_51_groupi_g18352(csa_tree_add_12_51_groupi_n_3389 ,csa_tree_add_12_51_groupi_n_598 ,csa_tree_add_12_51_groupi_n_1065);
  nor csa_tree_add_12_51_groupi_g18353(csa_tree_add_12_51_groupi_n_3388 ,csa_tree_add_12_51_groupi_n_670 ,csa_tree_add_12_51_groupi_n_1191);
  nor csa_tree_add_12_51_groupi_g18354(csa_tree_add_12_51_groupi_n_3387 ,csa_tree_add_12_51_groupi_n_1545 ,csa_tree_add_12_51_groupi_n_376);
  nor csa_tree_add_12_51_groupi_g18355(csa_tree_add_12_51_groupi_n_3386 ,csa_tree_add_12_51_groupi_n_1544 ,csa_tree_add_12_51_groupi_n_187);
  nor csa_tree_add_12_51_groupi_g18356(csa_tree_add_12_51_groupi_n_3385 ,csa_tree_add_12_51_groupi_n_1542 ,csa_tree_add_12_51_groupi_n_277);
  nor csa_tree_add_12_51_groupi_g18357(csa_tree_add_12_51_groupi_n_3384 ,csa_tree_add_12_51_groupi_n_1538 ,csa_tree_add_12_51_groupi_n_202);
  nor csa_tree_add_12_51_groupi_g18358(csa_tree_add_12_51_groupi_n_3383 ,csa_tree_add_12_51_groupi_n_1536 ,csa_tree_add_12_51_groupi_n_343);
  nor csa_tree_add_12_51_groupi_g18359(csa_tree_add_12_51_groupi_n_3382 ,csa_tree_add_12_51_groupi_n_1560 ,csa_tree_add_12_51_groupi_n_241);
  nor csa_tree_add_12_51_groupi_g18360(csa_tree_add_12_51_groupi_n_3381 ,csa_tree_add_12_51_groupi_n_921 ,csa_tree_add_12_51_groupi_n_193);
  nor csa_tree_add_12_51_groupi_g18361(csa_tree_add_12_51_groupi_n_3380 ,csa_tree_add_12_51_groupi_n_1410 ,csa_tree_add_12_51_groupi_n_1539);
  nor csa_tree_add_12_51_groupi_g18362(csa_tree_add_12_51_groupi_n_3379 ,csa_tree_add_12_51_groupi_n_544 ,csa_tree_add_12_51_groupi_n_1559);
  nor csa_tree_add_12_51_groupi_g18363(csa_tree_add_12_51_groupi_n_3378 ,csa_tree_add_12_51_groupi_n_681 ,csa_tree_add_12_51_groupi_n_1131);
  nor csa_tree_add_12_51_groupi_g18364(csa_tree_add_12_51_groupi_n_3377 ,csa_tree_add_12_51_groupi_n_1668 ,csa_tree_add_12_51_groupi_n_196);
  nor csa_tree_add_12_51_groupi_g18365(csa_tree_add_12_51_groupi_n_3376 ,csa_tree_add_12_51_groupi_n_643 ,csa_tree_add_12_51_groupi_n_1535);
  nor csa_tree_add_12_51_groupi_g18366(csa_tree_add_12_51_groupi_n_3375 ,csa_tree_add_12_51_groupi_n_1559 ,csa_tree_add_12_51_groupi_n_205);
  nor csa_tree_add_12_51_groupi_g18367(csa_tree_add_12_51_groupi_n_3374 ,csa_tree_add_12_51_groupi_n_1535 ,csa_tree_add_12_51_groupi_n_301);
  nor csa_tree_add_12_51_groupi_g18368(csa_tree_add_12_51_groupi_n_3373 ,csa_tree_add_12_51_groupi_n_1268 ,csa_tree_add_12_51_groupi_n_1134);
  nor csa_tree_add_12_51_groupi_g18369(csa_tree_add_12_51_groupi_n_3372 ,csa_tree_add_12_51_groupi_n_552 ,csa_tree_add_12_51_groupi_n_1545);
  nor csa_tree_add_12_51_groupi_g18370(csa_tree_add_12_51_groupi_n_3371 ,csa_tree_add_12_51_groupi_n_1541 ,csa_tree_add_12_51_groupi_n_235);
  nor csa_tree_add_12_51_groupi_g18371(csa_tree_add_12_51_groupi_n_3370 ,csa_tree_add_12_51_groupi_n_1673 ,csa_tree_add_12_51_groupi_n_346);
  nor csa_tree_add_12_51_groupi_g18372(csa_tree_add_12_51_groupi_n_3369 ,csa_tree_add_12_51_groupi_n_1563 ,csa_tree_add_12_51_groupi_n_298);
  nor csa_tree_add_12_51_groupi_g18373(csa_tree_add_12_51_groupi_n_3368 ,csa_tree_add_12_51_groupi_n_1065 ,csa_tree_add_12_51_groupi_n_430);
  nor csa_tree_add_12_51_groupi_g18374(csa_tree_add_12_51_groupi_n_3367 ,csa_tree_add_12_51_groupi_n_1487 ,csa_tree_add_12_51_groupi_n_412);
  nor csa_tree_add_12_51_groupi_g18375(csa_tree_add_12_51_groupi_n_3366 ,csa_tree_add_12_51_groupi_n_1412 ,csa_tree_add_12_51_groupi_n_1094);
  nor csa_tree_add_12_51_groupi_g18376(csa_tree_add_12_51_groupi_n_3365 ,csa_tree_add_12_51_groupi_n_1674 ,csa_tree_add_12_51_groupi_n_400);
  nor csa_tree_add_12_51_groupi_g18377(csa_tree_add_12_51_groupi_n_3364 ,csa_tree_add_12_51_groupi_n_1562 ,csa_tree_add_12_51_groupi_n_415);
  nor csa_tree_add_12_51_groupi_g18378(csa_tree_add_12_51_groupi_n_3363 ,csa_tree_add_12_51_groupi_n_1488 ,csa_tree_add_12_51_groupi_n_328);
  nor csa_tree_add_12_51_groupi_g18379(csa_tree_add_12_51_groupi_n_3362 ,csa_tree_add_12_51_groupi_n_1538 ,csa_tree_add_12_51_groupi_n_340);
  nor csa_tree_add_12_51_groupi_g18380(csa_tree_add_12_51_groupi_n_3361 ,csa_tree_add_12_51_groupi_n_1431 ,csa_tree_add_12_51_groupi_n_1095);
  nor csa_tree_add_12_51_groupi_g18381(csa_tree_add_12_51_groupi_n_3360 ,csa_tree_add_12_51_groupi_n_1487 ,csa_tree_add_12_51_groupi_n_325);
  nor csa_tree_add_12_51_groupi_g18382(csa_tree_add_12_51_groupi_n_3359 ,csa_tree_add_12_51_groupi_n_627 ,csa_tree_add_12_51_groupi_n_939);
  nor csa_tree_add_12_51_groupi_g18383(csa_tree_add_12_51_groupi_n_3358 ,csa_tree_add_12_51_groupi_n_1428 ,csa_tree_add_12_51_groupi_n_1064);
  nor csa_tree_add_12_51_groupi_g18384(csa_tree_add_12_51_groupi_n_3357 ,csa_tree_add_12_51_groupi_n_1667 ,csa_tree_add_12_51_groupi_n_244);
  nor csa_tree_add_12_51_groupi_g18385(csa_tree_add_12_51_groupi_n_3356 ,csa_tree_add_12_51_groupi_n_1443 ,csa_tree_add_12_51_groupi_n_1193);
  nor csa_tree_add_12_51_groupi_g18386(csa_tree_add_12_51_groupi_n_3355 ,csa_tree_add_12_51_groupi_n_1473 ,csa_tree_add_12_51_groupi_n_1562);
  nor csa_tree_add_12_51_groupi_g18387(csa_tree_add_12_51_groupi_n_3354 ,csa_tree_add_12_51_groupi_n_1743 ,csa_tree_add_12_51_groupi_n_1133);
  nor csa_tree_add_12_51_groupi_g18388(csa_tree_add_12_51_groupi_n_3353 ,csa_tree_add_12_51_groupi_n_1433 ,csa_tree_add_12_51_groupi_n_917);
  nor csa_tree_add_12_51_groupi_g18389(csa_tree_add_12_51_groupi_n_3352 ,csa_tree_add_12_51_groupi_n_1685 ,csa_tree_add_12_51_groupi_n_384);
  nor csa_tree_add_12_51_groupi_g18390(csa_tree_add_12_51_groupi_n_3351 ,csa_tree_add_12_51_groupi_n_1673 ,csa_tree_add_12_51_groupi_n_382);
  nor csa_tree_add_12_51_groupi_g18391(csa_tree_add_12_51_groupi_n_3350 ,csa_tree_add_12_51_groupi_n_1338 ,csa_tree_add_12_51_groupi_n_253);
  nor csa_tree_add_12_51_groupi_g18392(csa_tree_add_12_51_groupi_n_3349 ,csa_tree_add_12_51_groupi_n_1544 ,csa_tree_add_12_51_groupi_n_210);
  nor csa_tree_add_12_51_groupi_g18393(csa_tree_add_12_51_groupi_n_3348 ,csa_tree_add_12_51_groupi_n_1191 ,csa_tree_add_12_51_groupi_n_226);
  nor csa_tree_add_12_51_groupi_g18394(csa_tree_add_12_51_groupi_n_3347 ,csa_tree_add_12_51_groupi_n_1436 ,csa_tree_add_12_51_groupi_n_1094);
  nor csa_tree_add_12_51_groupi_g18395(csa_tree_add_12_51_groupi_n_3346 ,csa_tree_add_12_51_groupi_n_1407 ,csa_tree_add_12_51_groupi_n_938);
  nor csa_tree_add_12_51_groupi_g18396(csa_tree_add_12_51_groupi_n_3345 ,csa_tree_add_12_51_groupi_n_1454 ,csa_tree_add_12_51_groupi_n_1337);
  nor csa_tree_add_12_51_groupi_g18397(csa_tree_add_12_51_groupi_n_3344 ,csa_tree_add_12_51_groupi_n_1439 ,csa_tree_add_12_51_groupi_n_1130);
  nor csa_tree_add_12_51_groupi_g18398(csa_tree_add_12_51_groupi_n_3343 ,csa_tree_add_12_51_groupi_n_1749 ,csa_tree_add_12_51_groupi_n_1194);
  nor csa_tree_add_12_51_groupi_g18399(csa_tree_add_12_51_groupi_n_3342 ,csa_tree_add_12_51_groupi_n_1418 ,csa_tree_add_12_51_groupi_n_920);
  nor csa_tree_add_12_51_groupi_g18400(csa_tree_add_12_51_groupi_n_3341 ,csa_tree_add_12_51_groupi_n_523 ,csa_tree_add_12_51_groupi_n_921);
  nor csa_tree_add_12_51_groupi_g18401(csa_tree_add_12_51_groupi_n_3340 ,csa_tree_add_12_51_groupi_n_483 ,csa_tree_add_12_51_groupi_n_863);
  nor csa_tree_add_12_51_groupi_g18402(csa_tree_add_12_51_groupi_n_3339 ,csa_tree_add_12_51_groupi_n_1725 ,csa_tree_add_12_51_groupi_n_1130);
  nor csa_tree_add_12_51_groupi_g18403(csa_tree_add_12_51_groupi_n_3338 ,csa_tree_add_12_51_groupi_n_1421 ,csa_tree_add_12_51_groupi_n_864);
  nor csa_tree_add_12_51_groupi_g18404(csa_tree_add_12_51_groupi_n_3337 ,csa_tree_add_12_51_groupi_n_1809 ,csa_tree_add_12_51_groupi_n_1193);
  nor csa_tree_add_12_51_groupi_g18405(csa_tree_add_12_51_groupi_n_3336 ,csa_tree_add_12_51_groupi_n_1400 ,csa_tree_add_12_51_groupi_n_1133);
  nor csa_tree_add_12_51_groupi_g18406(csa_tree_add_12_51_groupi_n_3335 ,csa_tree_add_12_51_groupi_n_547 ,csa_tree_add_12_51_groupi_n_918);
  nor csa_tree_add_12_51_groupi_g18407(csa_tree_add_12_51_groupi_n_3334 ,csa_tree_add_12_51_groupi_n_589 ,csa_tree_add_12_51_groupi_n_1256);
  nor csa_tree_add_12_51_groupi_g18408(csa_tree_add_12_51_groupi_n_3333 ,csa_tree_add_12_51_groupi_n_1770 ,csa_tree_add_12_51_groupi_n_857);
  nor csa_tree_add_12_51_groupi_g18409(csa_tree_add_12_51_groupi_n_3332 ,csa_tree_add_12_51_groupi_n_517 ,csa_tree_add_12_51_groupi_n_914);
  nor csa_tree_add_12_51_groupi_g18410(csa_tree_add_12_51_groupi_n_3331 ,csa_tree_add_12_51_groupi_n_1445 ,csa_tree_add_12_51_groupi_n_1199);
  nor csa_tree_add_12_51_groupi_g18411(csa_tree_add_12_51_groupi_n_3330 ,csa_tree_add_12_51_groupi_n_1728 ,csa_tree_add_12_51_groupi_n_1553);
  nor csa_tree_add_12_51_groupi_g18412(csa_tree_add_12_51_groupi_n_3329 ,csa_tree_add_12_51_groupi_n_1794 ,csa_tree_add_12_51_groupi_n_1289);
  nor csa_tree_add_12_51_groupi_g18413(csa_tree_add_12_51_groupi_n_3328 ,csa_tree_add_12_51_groupi_n_601 ,csa_tree_add_12_51_groupi_n_912);
  nor csa_tree_add_12_51_groupi_g18414(csa_tree_add_12_51_groupi_n_3327 ,csa_tree_add_12_51_groupi_n_1695 ,csa_tree_add_12_51_groupi_n_1290);
  nor csa_tree_add_12_51_groupi_g18415(csa_tree_add_12_51_groupi_n_3326 ,csa_tree_add_12_51_groupi_n_1566 ,csa_tree_add_12_51_groupi_n_855);
  nor csa_tree_add_12_51_groupi_g18416(csa_tree_add_12_51_groupi_n_3325 ,csa_tree_add_12_51_groupi_n_1734 ,csa_tree_add_12_51_groupi_n_1125);
  nor csa_tree_add_12_51_groupi_g18417(csa_tree_add_12_51_groupi_n_3324 ,csa_tree_add_12_51_groupi_n_1737 ,csa_tree_add_12_51_groupi_n_1391);
  nor csa_tree_add_12_51_groupi_g18418(csa_tree_add_12_51_groupi_n_3323 ,csa_tree_add_12_51_groupi_n_1812 ,csa_tree_add_12_51_groupi_n_1211);
  nor csa_tree_add_12_51_groupi_g18419(csa_tree_add_12_51_groupi_n_3322 ,csa_tree_add_12_51_groupi_n_1568 ,csa_tree_add_12_51_groupi_n_1206);
  nor csa_tree_add_12_51_groupi_g18420(csa_tree_add_12_51_groupi_n_3321 ,csa_tree_add_12_51_groupi_n_520 ,csa_tree_add_12_51_groupi_n_858);
  nor csa_tree_add_12_51_groupi_g18421(csa_tree_add_12_51_groupi_n_3320 ,csa_tree_add_12_51_groupi_n_1758 ,csa_tree_add_12_51_groupi_n_1254);
  nor csa_tree_add_12_51_groupi_g18422(csa_tree_add_12_51_groupi_n_3319 ,csa_tree_add_12_51_groupi_n_592 ,csa_tree_add_12_51_groupi_n_854);
  nor csa_tree_add_12_51_groupi_g18423(csa_tree_add_12_51_groupi_n_3318 ,csa_tree_add_12_51_groupi_n_1782 ,csa_tree_add_12_51_groupi_n_1127);
  nor csa_tree_add_12_51_groupi_g18424(csa_tree_add_12_51_groupi_n_3317 ,csa_tree_add_12_51_groupi_n_1713 ,csa_tree_add_12_51_groupi_n_1209);
  nor csa_tree_add_12_51_groupi_g18425(csa_tree_add_12_51_groupi_n_3316 ,csa_tree_add_12_51_groupi_n_1779 ,csa_tree_add_12_51_groupi_n_1203);
  nor csa_tree_add_12_51_groupi_g18426(csa_tree_add_12_51_groupi_n_3315 ,csa_tree_add_12_51_groupi_n_1197 ,csa_tree_add_12_51_groupi_n_330);
  nor csa_tree_add_12_51_groupi_g18427(csa_tree_add_12_51_groupi_n_3314 ,csa_tree_add_12_51_groupi_n_1773 ,csa_tree_add_12_51_groupi_n_1128);
  nor csa_tree_add_12_51_groupi_g18428(csa_tree_add_12_51_groupi_n_3313 ,csa_tree_add_12_51_groupi_n_1547 ,csa_tree_add_12_51_groupi_n_184);
  nor csa_tree_add_12_51_groupi_g18429(csa_tree_add_12_51_groupi_n_3312 ,csa_tree_add_12_51_groupi_n_1791 ,csa_tree_add_12_51_groupi_n_855);
  nor csa_tree_add_12_51_groupi_g18430(csa_tree_add_12_51_groupi_n_3311 ,csa_tree_add_12_51_groupi_n_1200 ,csa_tree_add_12_51_groupi_n_465);
  nor csa_tree_add_12_51_groupi_g18431(csa_tree_add_12_51_groupi_n_3310 ,csa_tree_add_12_51_groupi_n_1767 ,csa_tree_add_12_51_groupi_n_1256);
  nor csa_tree_add_12_51_groupi_g18432(csa_tree_add_12_51_groupi_n_3309 ,csa_tree_add_12_51_groupi_n_1716 ,csa_tree_add_12_51_groupi_n_914);
  nor csa_tree_add_12_51_groupi_g18433(csa_tree_add_12_51_groupi_n_3308 ,csa_tree_add_12_51_groupi_n_613 ,csa_tree_add_12_51_groupi_n_857);
  nor csa_tree_add_12_51_groupi_g18434(csa_tree_add_12_51_groupi_n_3307 ,csa_tree_add_12_51_groupi_n_1403 ,csa_tree_add_12_51_groupi_n_1548);
  nor csa_tree_add_12_51_groupi_g18435(csa_tree_add_12_51_groupi_n_3306 ,csa_tree_add_12_51_groupi_n_1128 ,csa_tree_add_12_51_groupi_n_364);
  nor csa_tree_add_12_51_groupi_g18436(csa_tree_add_12_51_groupi_n_3305 ,csa_tree_add_12_51_groupi_n_1746 ,csa_tree_add_12_51_groupi_n_1257);
  nor csa_tree_add_12_51_groupi_g18437(csa_tree_add_12_51_groupi_n_3304 ,csa_tree_add_12_51_groupi_n_631 ,csa_tree_add_12_51_groupi_n_1200);
  nor csa_tree_add_12_51_groupi_g18438(csa_tree_add_12_51_groupi_n_3303 ,csa_tree_add_12_51_groupi_n_1394 ,csa_tree_add_12_51_groupi_n_249);
  nor csa_tree_add_12_51_groupi_g18439(csa_tree_add_12_51_groupi_n_3302 ,csa_tree_add_12_51_groupi_n_1797 ,csa_tree_add_12_51_groupi_n_915);
  nor csa_tree_add_12_51_groupi_g18440(csa_tree_add_12_51_groupi_n_3301 ,csa_tree_add_12_51_groupi_n_640 ,csa_tree_add_12_51_groupi_n_1394);
  nor csa_tree_add_12_51_groupi_g18441(csa_tree_add_12_51_groupi_n_3300 ,csa_tree_add_12_51_groupi_n_655 ,csa_tree_add_12_51_groupi_n_1199);
  nor csa_tree_add_12_51_groupi_g18442(csa_tree_add_12_51_groupi_n_3299 ,csa_tree_add_12_51_groupi_n_1707 ,csa_tree_add_12_51_groupi_n_911);
  nor csa_tree_add_12_51_groupi_g18443(csa_tree_add_12_51_groupi_n_3298 ,csa_tree_add_12_51_groupi_n_1554 ,csa_tree_add_12_51_groupi_n_199);
  nor csa_tree_add_12_51_groupi_g18444(csa_tree_add_12_51_groupi_n_3297 ,csa_tree_add_12_51_groupi_n_1547 ,csa_tree_add_12_51_groupi_n_354);
  nor csa_tree_add_12_51_groupi_g18445(csa_tree_add_12_51_groupi_n_3296 ,csa_tree_add_12_51_groupi_n_1761 ,csa_tree_add_12_51_groupi_n_1196);
  nor csa_tree_add_12_51_groupi_g18446(csa_tree_add_12_51_groupi_n_3295 ,csa_tree_add_12_51_groupi_n_565 ,csa_tree_add_12_51_groupi_n_1127);
  nor csa_tree_add_12_51_groupi_g18447(csa_tree_add_12_51_groupi_n_3294 ,csa_tree_add_12_51_groupi_n_556 ,csa_tree_add_12_51_groupi_n_1212);
  nor csa_tree_add_12_51_groupi_g18448(csa_tree_add_12_51_groupi_n_3293 ,csa_tree_add_12_51_groupi_n_1698 ,csa_tree_add_12_51_groupi_n_1395);
  nor csa_tree_add_12_51_groupi_g18449(csa_tree_add_12_51_groupi_n_3292 ,csa_tree_add_12_51_groupi_n_1701 ,csa_tree_add_12_51_groupi_n_1196);
  nor csa_tree_add_12_51_groupi_g18450(csa_tree_add_12_51_groupi_n_3291 ,csa_tree_add_12_51_groupi_n_562 ,csa_tree_add_12_51_groupi_n_1392);
  nor csa_tree_add_12_51_groupi_g18451(csa_tree_add_12_51_groupi_n_3290 ,csa_tree_add_12_51_groupi_n_1208 ,csa_tree_add_12_51_groupi_n_424);
  nor csa_tree_add_12_51_groupi_g18452(csa_tree_add_12_51_groupi_n_3289 ,csa_tree_add_12_51_groupi_n_1764 ,csa_tree_add_12_51_groupi_n_1124);
  nor csa_tree_add_12_51_groupi_g18453(csa_tree_add_12_51_groupi_n_3288 ,csa_tree_add_12_51_groupi_n_1553 ,csa_tree_add_12_51_groupi_n_441);
  nor csa_tree_add_12_51_groupi_g18454(csa_tree_add_12_51_groupi_n_3287 ,csa_tree_add_12_51_groupi_n_1293 ,csa_tree_add_12_51_groupi_n_376);
  nor csa_tree_add_12_51_groupi_g18455(csa_tree_add_12_51_groupi_n_3286 ,csa_tree_add_12_51_groupi_n_1202 ,csa_tree_add_12_51_groupi_n_399);
  nor csa_tree_add_12_51_groupi_g18456(csa_tree_add_12_51_groupi_n_3285 ,csa_tree_add_12_51_groupi_n_1704 ,csa_tree_add_12_51_groupi_n_854);
  nor csa_tree_add_12_51_groupi_g18457(csa_tree_add_12_51_groupi_n_3284 ,csa_tree_add_12_51_groupi_n_1548 ,csa_tree_add_12_51_groupi_n_267);
  nor csa_tree_add_12_51_groupi_g18458(csa_tree_add_12_51_groupi_n_3283 ,csa_tree_add_12_51_groupi_n_1205 ,csa_tree_add_12_51_groupi_n_270);
  nor csa_tree_add_12_51_groupi_g18459(csa_tree_add_12_51_groupi_n_3282 ,csa_tree_add_12_51_groupi_n_912 ,csa_tree_add_12_51_groupi_n_201);
  nor csa_tree_add_12_51_groupi_g18460(csa_tree_add_12_51_groupi_n_3281 ,csa_tree_add_12_51_groupi_n_1257 ,csa_tree_add_12_51_groupi_n_429);
  nor csa_tree_add_12_51_groupi_g18461(csa_tree_add_12_51_groupi_n_3280 ,csa_tree_add_12_51_groupi_n_1203 ,csa_tree_add_12_51_groupi_n_300);
  nor csa_tree_add_12_51_groupi_g18462(csa_tree_add_12_51_groupi_n_3279 ,csa_tree_add_12_51_groupi_n_1253 ,csa_tree_add_12_51_groupi_n_342);
  nor csa_tree_add_12_51_groupi_g18463(csa_tree_add_12_51_groupi_n_3278 ,csa_tree_add_12_51_groupi_n_1391 ,csa_tree_add_12_51_groupi_n_411);
  nor csa_tree_add_12_51_groupi_g18464(csa_tree_add_12_51_groupi_n_3277 ,csa_tree_add_12_51_groupi_n_1788 ,csa_tree_add_12_51_groupi_n_1205);
  nor csa_tree_add_12_51_groupi_g18465(csa_tree_add_12_51_groupi_n_3276 ,csa_tree_add_12_51_groupi_n_1289 ,csa_tree_add_12_51_groupi_n_402);
  nor csa_tree_add_12_51_groupi_g18466(csa_tree_add_12_51_groupi_n_3275 ,csa_tree_add_12_51_groupi_n_1292 ,csa_tree_add_12_51_groupi_n_285);
  nor csa_tree_add_12_51_groupi_g18467(csa_tree_add_12_51_groupi_n_3274 ,csa_tree_add_12_51_groupi_n_1125 ,csa_tree_add_12_51_groupi_n_471);
  nor csa_tree_add_12_51_groupi_g18468(csa_tree_add_12_51_groupi_n_3273 ,csa_tree_add_12_51_groupi_n_1290 ,csa_tree_add_12_51_groupi_n_351);
  nor csa_tree_add_12_51_groupi_g18469(csa_tree_add_12_51_groupi_n_3272 ,csa_tree_add_12_51_groupi_n_1211 ,csa_tree_add_12_51_groupi_n_234);
  nor csa_tree_add_12_51_groupi_g18470(csa_tree_add_12_51_groupi_n_3271 ,csa_tree_add_12_51_groupi_n_1254 ,csa_tree_add_12_51_groupi_n_406);
  nor csa_tree_add_12_51_groupi_g18471(csa_tree_add_12_51_groupi_n_3270 ,csa_tree_add_12_51_groupi_n_1209 ,csa_tree_add_12_51_groupi_n_318);
  nor csa_tree_add_12_51_groupi_g18472(csa_tree_add_12_51_groupi_n_3269 ,csa_tree_add_12_51_groupi_n_1574 ,csa_tree_add_12_51_groupi_n_327);
  nor csa_tree_add_12_51_groupi_g18473(csa_tree_add_12_51_groupi_n_3268 ,csa_tree_add_12_51_groupi_n_1686 ,csa_tree_add_12_51_groupi_n_345);
  nor csa_tree_add_12_51_groupi_g18474(csa_tree_add_12_51_groupi_n_3267 ,csa_tree_add_12_51_groupi_n_1119 ,csa_tree_add_12_51_groupi_n_414);
  nor csa_tree_add_12_51_groupi_g18475(csa_tree_add_12_51_groupi_n_3266 ,csa_tree_add_12_51_groupi_n_1520 ,csa_tree_add_12_51_groupi_n_360);
  nor csa_tree_add_12_51_groupi_g18476(csa_tree_add_12_51_groupi_n_3265 ,csa_tree_add_12_51_groupi_n_1575 ,csa_tree_add_12_51_groupi_n_279);
  nor csa_tree_add_12_51_groupi_g18477(csa_tree_add_12_51_groupi_n_3264 ,csa_tree_add_12_51_groupi_n_1340 ,csa_tree_add_12_51_groupi_n_438);
  nor csa_tree_add_12_51_groupi_g18478(csa_tree_add_12_51_groupi_n_3263 ,csa_tree_add_12_51_groupi_n_1497 ,csa_tree_add_12_51_groupi_n_297);
  nor csa_tree_add_12_51_groupi_g18479(csa_tree_add_12_51_groupi_n_3262 ,csa_tree_add_12_51_groupi_n_1496 ,csa_tree_add_12_51_groupi_n_453);
  nor csa_tree_add_12_51_groupi_g18480(csa_tree_add_12_51_groupi_n_3261 ,csa_tree_add_12_51_groupi_n_1302 ,csa_tree_add_12_51_groupi_n_324);
  nor csa_tree_add_12_51_groupi_g18481(csa_tree_add_12_51_groupi_n_3260 ,csa_tree_add_12_51_groupi_n_1521 ,csa_tree_add_12_51_groupi_n_381);
  nor csa_tree_add_12_51_groupi_g18482(csa_tree_add_12_51_groupi_n_3259 ,csa_tree_add_12_51_groupi_n_1496 ,csa_tree_add_12_51_groupi_n_459);
  nor csa_tree_add_12_51_groupi_g18483(csa_tree_add_12_51_groupi_n_3258 ,csa_tree_add_12_51_groupi_n_1305 ,csa_tree_add_12_51_groupi_n_211);
  nor csa_tree_add_12_51_groupi_g18484(csa_tree_add_12_51_groupi_n_3257 ,csa_tree_add_12_51_groupi_n_1304 ,csa_tree_add_12_51_groupi_n_316);
  nor csa_tree_add_12_51_groupi_g18485(csa_tree_add_12_51_groupi_n_3256 ,csa_tree_add_12_51_groupi_n_1301 ,csa_tree_add_12_51_groupi_n_385);
  or csa_tree_add_12_51_groupi_g18486(csa_tree_add_12_51_groupi_n_3558 ,csa_tree_add_12_51_groupi_n_2706 ,csa_tree_add_12_51_groupi_n_2795);
  or csa_tree_add_12_51_groupi_g18487(csa_tree_add_12_51_groupi_n_3557 ,csa_tree_add_12_51_groupi_n_2674 ,csa_tree_add_12_51_groupi_n_2822);
  or csa_tree_add_12_51_groupi_g18488(csa_tree_add_12_51_groupi_n_3556 ,csa_tree_add_12_51_groupi_n_2610 ,csa_tree_add_12_51_groupi_n_2826);
  or csa_tree_add_12_51_groupi_g18489(csa_tree_add_12_51_groupi_n_3554 ,csa_tree_add_12_51_groupi_n_2667 ,csa_tree_add_12_51_groupi_n_2803);
  or csa_tree_add_12_51_groupi_g18490(csa_tree_add_12_51_groupi_n_3553 ,csa_tree_add_12_51_groupi_n_2688 ,csa_tree_add_12_51_groupi_n_2819);
  or csa_tree_add_12_51_groupi_g18491(csa_tree_add_12_51_groupi_n_3552 ,csa_tree_add_12_51_groupi_n_2598 ,csa_tree_add_12_51_groupi_n_2812);
  or csa_tree_add_12_51_groupi_g18492(csa_tree_add_12_51_groupi_n_3551 ,csa_tree_add_12_51_groupi_n_2633 ,csa_tree_add_12_51_groupi_n_2790);
  or csa_tree_add_12_51_groupi_g18493(csa_tree_add_12_51_groupi_n_3550 ,csa_tree_add_12_51_groupi_n_2574 ,csa_tree_add_12_51_groupi_n_2800);
  or csa_tree_add_12_51_groupi_g18494(csa_tree_add_12_51_groupi_n_3549 ,csa_tree_add_12_51_groupi_n_2632 ,csa_tree_add_12_51_groupi_n_2808);
  or csa_tree_add_12_51_groupi_g18495(csa_tree_add_12_51_groupi_n_3548 ,csa_tree_add_12_51_groupi_n_2623 ,csa_tree_add_12_51_groupi_n_2815);
  or csa_tree_add_12_51_groupi_g18496(csa_tree_add_12_51_groupi_n_3547 ,csa_tree_add_12_51_groupi_n_2713 ,csa_tree_add_12_51_groupi_n_2814);
  or csa_tree_add_12_51_groupi_g18497(csa_tree_add_12_51_groupi_n_3545 ,csa_tree_add_12_51_groupi_n_2628 ,csa_tree_add_12_51_groupi_n_2783);
  or csa_tree_add_12_51_groupi_g18498(csa_tree_add_12_51_groupi_n_3544 ,csa_tree_add_12_51_groupi_n_2676 ,csa_tree_add_12_51_groupi_n_2824);
  or csa_tree_add_12_51_groupi_g18499(csa_tree_add_12_51_groupi_n_3542 ,csa_tree_add_12_51_groupi_n_2675 ,csa_tree_add_12_51_groupi_n_2867);
  or csa_tree_add_12_51_groupi_g18500(csa_tree_add_12_51_groupi_n_3540 ,csa_tree_add_12_51_groupi_n_2582 ,csa_tree_add_12_51_groupi_n_2792);
  or csa_tree_add_12_51_groupi_g18501(csa_tree_add_12_51_groupi_n_3539 ,csa_tree_add_12_51_groupi_n_2620 ,csa_tree_add_12_51_groupi_n_2816);
  or csa_tree_add_12_51_groupi_g18502(csa_tree_add_12_51_groupi_n_3537 ,csa_tree_add_12_51_groupi_n_2619 ,csa_tree_add_12_51_groupi_n_2788);
  or csa_tree_add_12_51_groupi_g18503(csa_tree_add_12_51_groupi_n_3536 ,csa_tree_add_12_51_groupi_n_2576 ,csa_tree_add_12_51_groupi_n_2821);
  or csa_tree_add_12_51_groupi_g18504(csa_tree_add_12_51_groupi_n_3534 ,csa_tree_add_12_51_groupi_n_2671 ,csa_tree_add_12_51_groupi_n_2813);
  or csa_tree_add_12_51_groupi_g18505(csa_tree_add_12_51_groupi_n_3532 ,csa_tree_add_12_51_groupi_n_2665 ,csa_tree_add_12_51_groupi_n_2787);
  or csa_tree_add_12_51_groupi_g18506(csa_tree_add_12_51_groupi_n_3530 ,csa_tree_add_12_51_groupi_n_2627 ,csa_tree_add_12_51_groupi_n_2825);
  or csa_tree_add_12_51_groupi_g18507(csa_tree_add_12_51_groupi_n_3529 ,csa_tree_add_12_51_groupi_n_2715 ,csa_tree_add_12_51_groupi_n_2798);
  or csa_tree_add_12_51_groupi_g18508(csa_tree_add_12_51_groupi_n_3528 ,csa_tree_add_12_51_groupi_n_2584 ,csa_tree_add_12_51_groupi_n_2786);
  or csa_tree_add_12_51_groupi_g18509(csa_tree_add_12_51_groupi_n_3527 ,csa_tree_add_12_51_groupi_n_2417 ,csa_tree_add_12_51_groupi_n_2871);
  or csa_tree_add_12_51_groupi_g18510(csa_tree_add_12_51_groupi_n_3525 ,csa_tree_add_12_51_groupi_n_2608 ,csa_tree_add_12_51_groupi_n_2818);
  or csa_tree_add_12_51_groupi_g18511(csa_tree_add_12_51_groupi_n_3524 ,csa_tree_add_12_51_groupi_n_2597 ,csa_tree_add_12_51_groupi_n_2789);
  or csa_tree_add_12_51_groupi_g18512(csa_tree_add_12_51_groupi_n_3522 ,csa_tree_add_12_51_groupi_n_2631 ,csa_tree_add_12_51_groupi_n_2817);
  or csa_tree_add_12_51_groupi_g18513(csa_tree_add_12_51_groupi_n_3521 ,csa_tree_add_12_51_groupi_n_2578 ,csa_tree_add_12_51_groupi_n_2810);
  or csa_tree_add_12_51_groupi_g18514(csa_tree_add_12_51_groupi_n_3520 ,csa_tree_add_12_51_groupi_n_2609 ,csa_tree_add_12_51_groupi_n_2805);
  or csa_tree_add_12_51_groupi_g18515(csa_tree_add_12_51_groupi_n_3518 ,csa_tree_add_12_51_groupi_n_2590 ,csa_tree_add_12_51_groupi_n_2802);
  or csa_tree_add_12_51_groupi_g18516(csa_tree_add_12_51_groupi_n_3517 ,csa_tree_add_12_51_groupi_n_2581 ,csa_tree_add_12_51_groupi_n_2797);
  or csa_tree_add_12_51_groupi_g18517(csa_tree_add_12_51_groupi_n_3516 ,csa_tree_add_12_51_groupi_n_2735 ,csa_tree_add_12_51_groupi_n_2820);
  or csa_tree_add_12_51_groupi_g18518(csa_tree_add_12_51_groupi_n_3513 ,csa_tree_add_12_51_groupi_n_2615 ,csa_tree_add_12_51_groupi_n_2827);
  or csa_tree_add_12_51_groupi_g18519(csa_tree_add_12_51_groupi_n_3511 ,csa_tree_add_12_51_groupi_n_2595 ,csa_tree_add_12_51_groupi_n_2809);
  or csa_tree_add_12_51_groupi_g18520(csa_tree_add_12_51_groupi_n_3510 ,csa_tree_add_12_51_groupi_n_2626 ,csa_tree_add_12_51_groupi_n_2794);
  and csa_tree_add_12_51_groupi_g18521(csa_tree_add_12_51_groupi_n_3508 ,csa_tree_add_12_51_groupi_n_2872 ,csa_tree_add_12_51_groupi_n_2888);
  and csa_tree_add_12_51_groupi_g18522(csa_tree_add_12_51_groupi_n_3507 ,csa_tree_add_12_51_groupi_n_2874 ,csa_tree_add_12_51_groupi_n_2879);
  and csa_tree_add_12_51_groupi_g18523(csa_tree_add_12_51_groupi_n_3506 ,csa_tree_add_12_51_groupi_n_2881 ,csa_tree_add_12_51_groupi_n_2895);
  and csa_tree_add_12_51_groupi_g18524(csa_tree_add_12_51_groupi_n_3505 ,csa_tree_add_12_51_groupi_n_2900 ,csa_tree_add_12_51_groupi_n_2886);
  and csa_tree_add_12_51_groupi_g18525(csa_tree_add_12_51_groupi_n_3504 ,csa_tree_add_12_51_groupi_n_2890 ,csa_tree_add_12_51_groupi_n_2884);
  and csa_tree_add_12_51_groupi_g18526(csa_tree_add_12_51_groupi_n_3503 ,csa_tree_add_12_51_groupi_n_2887 ,csa_tree_add_12_51_groupi_n_2891);
  and csa_tree_add_12_51_groupi_g18527(csa_tree_add_12_51_groupi_n_3502 ,csa_tree_add_12_51_groupi_n_2876 ,csa_tree_add_12_51_groupi_n_2898);
  and csa_tree_add_12_51_groupi_g18528(csa_tree_add_12_51_groupi_n_3501 ,csa_tree_add_12_51_groupi_n_2880 ,csa_tree_add_12_51_groupi_n_2906);
  and csa_tree_add_12_51_groupi_g18529(csa_tree_add_12_51_groupi_n_3500 ,csa_tree_add_12_51_groupi_n_2903 ,csa_tree_add_12_51_groupi_n_2892);
  and csa_tree_add_12_51_groupi_g18530(csa_tree_add_12_51_groupi_n_3499 ,csa_tree_add_12_51_groupi_n_2896 ,csa_tree_add_12_51_groupi_n_2904);
  and csa_tree_add_12_51_groupi_g18531(csa_tree_add_12_51_groupi_n_3498 ,csa_tree_add_12_51_groupi_n_2873 ,csa_tree_add_12_51_groupi_n_2893);
  and csa_tree_add_12_51_groupi_g18532(csa_tree_add_12_51_groupi_n_3497 ,csa_tree_add_12_51_groupi_n_2899 ,csa_tree_add_12_51_groupi_n_2894);
  not csa_tree_add_12_51_groupi_g18533(csa_tree_add_12_51_groupi_n_3240 ,csa_tree_add_12_51_groupi_n_3239);
  not csa_tree_add_12_51_groupi_g18534(csa_tree_add_12_51_groupi_n_3238 ,csa_tree_add_12_51_groupi_n_3237);
  not csa_tree_add_12_51_groupi_g18535(csa_tree_add_12_51_groupi_n_3236 ,csa_tree_add_12_51_groupi_n_3235);
  not csa_tree_add_12_51_groupi_g18536(csa_tree_add_12_51_groupi_n_3233 ,csa_tree_add_12_51_groupi_n_3234);
  not csa_tree_add_12_51_groupi_g18537(csa_tree_add_12_51_groupi_n_3231 ,csa_tree_add_12_51_groupi_n_3230);
  nor csa_tree_add_12_51_groupi_g18538(csa_tree_add_12_51_groupi_n_3228 ,csa_tree_add_12_51_groupi_n_553 ,csa_tree_add_12_51_groupi_n_897);
  nor csa_tree_add_12_51_groupi_g18539(csa_tree_add_12_51_groupi_n_3227 ,csa_tree_add_12_51_groupi_n_66 ,csa_tree_add_12_51_groupi_n_836);
  nor csa_tree_add_12_51_groupi_g18540(csa_tree_add_12_51_groupi_n_3226 ,csa_tree_add_12_51_groupi_n_92 ,csa_tree_add_12_51_groupi_n_833);
  nor csa_tree_add_12_51_groupi_g18541(csa_tree_add_12_51_groupi_n_3225 ,csa_tree_add_12_51_groupi_n_78 ,csa_tree_add_12_51_groupi_n_167);
  nor csa_tree_add_12_51_groupi_g18542(csa_tree_add_12_51_groupi_n_3224 ,csa_tree_add_12_51_groupi_n_82 ,csa_tree_add_12_51_groupi_n_836);
  nor csa_tree_add_12_51_groupi_g18543(csa_tree_add_12_51_groupi_n_3223 ,csa_tree_add_12_51_groupi_n_86 ,csa_tree_add_12_51_groupi_n_837);
  nor csa_tree_add_12_51_groupi_g18544(csa_tree_add_12_51_groupi_n_3222 ,csa_tree_add_12_51_groupi_n_72 ,csa_tree_add_12_51_groupi_n_834);
  nor csa_tree_add_12_51_groupi_g18545(csa_tree_add_12_51_groupi_n_3221 ,csa_tree_add_12_51_groupi_n_76 ,csa_tree_add_12_51_groupi_n_852);
  nor csa_tree_add_12_51_groupi_g18546(csa_tree_add_12_51_groupi_n_3220 ,csa_tree_add_12_51_groupi_n_90 ,csa_tree_add_12_51_groupi_n_1995);
  nor csa_tree_add_12_51_groupi_g18547(csa_tree_add_12_51_groupi_n_3219 ,csa_tree_add_12_51_groupi_n_70 ,csa_tree_add_12_51_groupi_n_833);
  nor csa_tree_add_12_51_groupi_g18548(csa_tree_add_12_51_groupi_n_3218 ,csa_tree_add_12_51_groupi_n_1383 ,csa_tree_add_12_51_groupi_n_136);
  nor csa_tree_add_12_51_groupi_g18549(csa_tree_add_12_51_groupi_n_3217 ,csa_tree_add_12_51_groupi_n_1377 ,csa_tree_add_12_51_groupi_n_139);
  nor csa_tree_add_12_51_groupi_g18550(csa_tree_add_12_51_groupi_n_3216 ,csa_tree_add_12_51_groupi_n_1275 ,csa_tree_add_12_51_groupi_n_128);
  nor csa_tree_add_12_51_groupi_g18551(csa_tree_add_12_51_groupi_n_3215 ,csa_tree_add_12_51_groupi_n_1512 ,csa_tree_add_12_51_groupi_n_145);
  nor csa_tree_add_12_51_groupi_g18552(csa_tree_add_12_51_groupi_n_3214 ,csa_tree_add_12_51_groupi_n_1515 ,csa_tree_add_12_51_groupi_n_228);
  nor csa_tree_add_12_51_groupi_g18553(csa_tree_add_12_51_groupi_n_3213 ,csa_tree_add_12_51_groupi_n_450 ,csa_tree_add_12_51_groupi_n_954);
  nor csa_tree_add_12_51_groupi_g18554(csa_tree_add_12_51_groupi_n_3212 ,csa_tree_add_12_51_groupi_n_457 ,csa_tree_add_12_51_groupi_n_1164);
  nor csa_tree_add_12_51_groupi_g18555(csa_tree_add_12_51_groupi_n_3211 ,csa_tree_add_12_51_groupi_n_1188 ,csa_tree_add_12_51_groupi_n_294);
  nor csa_tree_add_12_51_groupi_g18556(csa_tree_add_12_51_groupi_n_3210 ,csa_tree_add_12_51_groupi_n_1233 ,csa_tree_add_12_51_groupi_n_134);
  nor csa_tree_add_12_51_groupi_g18557(csa_tree_add_12_51_groupi_n_3209 ,csa_tree_add_12_51_groupi_n_1506 ,csa_tree_add_12_51_groupi_n_131);
  nor csa_tree_add_12_51_groupi_g18558(csa_tree_add_12_51_groupi_n_3208 ,csa_tree_add_12_51_groupi_n_1368 ,csa_tree_add_12_51_groupi_n_149);
  nor csa_tree_add_12_51_groupi_g18559(csa_tree_add_12_51_groupi_n_3207 ,csa_tree_add_12_51_groupi_n_1662 ,csa_tree_add_12_51_groupi_n_409);
  and csa_tree_add_12_51_groupi_g18560(csa_tree_add_12_51_groupi_n_3206 ,csa_tree_add_12_51_groupi_n_37 ,csa_tree_add_12_51_groupi_n_705);
  and csa_tree_add_12_51_groupi_g18561(csa_tree_add_12_51_groupi_n_3205 ,csa_tree_add_12_51_groupi_n_43 ,csa_tree_add_12_51_groupi_n_702);
  and csa_tree_add_12_51_groupi_g18562(csa_tree_add_12_51_groupi_n_3204 ,csa_tree_add_12_51_groupi_n_28 ,csa_tree_add_12_51_groupi_n_905);
  nor csa_tree_add_12_51_groupi_g18563(csa_tree_add_12_51_groupi_n_3203 ,csa_tree_add_12_51_groupi_n_697 ,csa_tree_add_12_51_groupi_n_1068);
  nor csa_tree_add_12_51_groupi_g18564(csa_tree_add_12_51_groupi_n_3202 ,csa_tree_add_12_51_groupi_n_1466 ,csa_tree_add_12_51_groupi_n_933);
  nor csa_tree_add_12_51_groupi_g18565(csa_tree_add_12_51_groupi_n_3201 ,csa_tree_add_12_51_groupi_n_1263 ,csa_tree_add_12_51_groupi_n_975);
  nor csa_tree_add_12_51_groupi_g18566(csa_tree_add_12_51_groupi_n_3200 ,csa_tree_add_12_51_groupi_n_1469 ,csa_tree_add_12_51_groupi_n_882);
  nor csa_tree_add_12_51_groupi_g18567(csa_tree_add_12_51_groupi_n_3199 ,csa_tree_add_12_51_groupi_n_1692 ,csa_tree_add_12_51_groupi_n_890);
  nor csa_tree_add_12_51_groupi_g18568(csa_tree_add_12_51_groupi_n_3198 ,csa_tree_add_12_51_groupi_n_1805 ,csa_tree_add_12_51_groupi_n_705);
  nor csa_tree_add_12_51_groupi_g18569(csa_tree_add_12_51_groupi_n_3197 ,csa_tree_add_12_51_groupi_n_657 ,csa_tree_add_12_51_groupi_n_1100);
  nor csa_tree_add_12_51_groupi_g18570(csa_tree_add_12_51_groupi_n_3196 ,csa_tree_add_12_51_groupi_n_1122 ,csa_tree_add_12_51_groupi_n_306);
  nor csa_tree_add_12_51_groupi_g18571(csa_tree_add_12_51_groupi_n_3195 ,csa_tree_add_12_51_groupi_n_1806 ,csa_tree_add_12_51_groupi_n_1187);
  nor csa_tree_add_12_51_groupi_g18572(csa_tree_add_12_51_groupi_n_3194 ,csa_tree_add_12_51_groupi_n_1281 ,csa_tree_add_12_51_groupi_n_435);
  nor csa_tree_add_12_51_groupi_g18573(csa_tree_add_12_51_groupi_n_3193 ,csa_tree_add_12_51_groupi_n_1479 ,csa_tree_add_12_51_groupi_n_207);
  nor csa_tree_add_12_51_groupi_g18574(csa_tree_add_12_51_groupi_n_3192 ,csa_tree_add_12_51_groupi_n_1533 ,csa_tree_add_12_51_groupi_n_420);
  nor csa_tree_add_12_51_groupi_g18575(csa_tree_add_12_51_groupi_n_3191 ,csa_tree_add_12_51_groupi_n_1230 ,csa_tree_add_12_51_groupi_n_310);
  nor csa_tree_add_12_51_groupi_g18576(csa_tree_add_12_51_groupi_n_3190 ,csa_tree_add_12_51_groupi_n_1299 ,csa_tree_add_12_51_groupi_n_219);
  nor csa_tree_add_12_51_groupi_g18577(csa_tree_add_12_51_groupi_n_3189 ,csa_tree_add_12_51_groupi_n_1314 ,csa_tree_add_12_51_groupi_n_336);
  nor csa_tree_add_12_51_groupi_g18578(csa_tree_add_12_51_groupi_n_3188 ,csa_tree_add_12_51_groupi_n_481 ,csa_tree_add_12_51_groupi_n_1515);
  nor csa_tree_add_12_51_groupi_g18579(csa_tree_add_12_51_groupi_n_3187 ,csa_tree_add_12_51_groupi_n_526 ,csa_tree_add_12_51_groupi_n_1055);
  nor csa_tree_add_12_51_groupi_g18580(csa_tree_add_12_51_groupi_n_3186 ,csa_tree_add_12_51_groupi_n_1571 ,csa_tree_add_12_51_groupi_n_1346);
  nor csa_tree_add_12_51_groupi_g18581(csa_tree_add_12_51_groupi_n_3185 ,csa_tree_add_12_51_groupi_n_1802 ,csa_tree_add_12_51_groupi_n_896);
  nor csa_tree_add_12_51_groupi_g18582(csa_tree_add_12_51_groupi_n_3184 ,csa_tree_add_12_51_groupi_n_1239 ,csa_tree_add_12_51_groupi_n_373);
  nor csa_tree_add_12_51_groupi_g18583(csa_tree_add_12_51_groupi_n_3183 ,csa_tree_add_12_51_groupi_n_1266 ,csa_tree_add_12_51_groupi_n_924);
  nor csa_tree_add_12_51_groupi_g18584(csa_tree_add_12_51_groupi_n_3182 ,csa_tree_add_12_51_groupi_n_664 ,csa_tree_add_12_51_groupi_n_1481);
  nor csa_tree_add_12_51_groupi_g18585(csa_tree_add_12_51_groupi_n_3181 ,csa_tree_add_12_51_groupi_n_505 ,csa_tree_add_12_51_groupi_n_1233);
  nor csa_tree_add_12_51_groupi_g18586(csa_tree_add_12_51_groupi_n_3180 ,csa_tree_add_12_51_groupi_n_1691 ,csa_tree_add_12_51_groupi_n_1107);
  nor csa_tree_add_12_51_groupi_g18587(csa_tree_add_12_51_groupi_n_3179 ,csa_tree_add_12_51_groupi_n_1242 ,csa_tree_add_12_51_groupi_n_463);
  nor csa_tree_add_12_51_groupi_g18588(csa_tree_add_12_51_groupi_n_3178 ,csa_tree_add_12_51_groupi_n_1272 ,csa_tree_add_12_51_groupi_n_321);
  nor csa_tree_add_12_51_groupi_g18589(csa_tree_add_12_51_groupi_n_3177 ,csa_tree_add_12_51_groupi_n_1244 ,csa_tree_add_12_51_groupi_n_231);
  nor csa_tree_add_12_51_groupi_g18590(csa_tree_add_12_51_groupi_n_3176 ,csa_tree_add_12_51_groupi_n_1163 ,csa_tree_add_12_51_groupi_n_258);
  nor csa_tree_add_12_51_groupi_g18591(csa_tree_add_12_51_groupi_n_3175 ,csa_tree_add_12_51_groupi_n_1323 ,csa_tree_add_12_51_groupi_n_303);
  nor csa_tree_add_12_51_groupi_g18592(csa_tree_add_12_51_groupi_n_3174 ,csa_tree_add_12_51_groupi_n_1557 ,csa_tree_add_12_51_groupi_n_288);
  nor csa_tree_add_12_51_groupi_g18593(csa_tree_add_12_51_groupi_n_3173 ,csa_tree_add_12_51_groupi_n_1448 ,csa_tree_add_12_51_groupi_n_906);
  nor csa_tree_add_12_51_groupi_g18594(csa_tree_add_12_51_groupi_n_3172 ,csa_tree_add_12_51_groupi_n_1413 ,csa_tree_add_12_51_groupi_n_702);
  nor csa_tree_add_12_51_groupi_g18595(csa_tree_add_12_51_groupi_n_3171 ,csa_tree_add_12_51_groupi_n_570 ,csa_tree_add_12_51_groupi_n_923);
  nor csa_tree_add_12_51_groupi_g18596(csa_tree_add_12_51_groupi_n_3170 ,csa_tree_add_12_51_groupi_n_498 ,csa_tree_add_12_51_groupi_n_1241);
  nor csa_tree_add_12_51_groupi_g18597(csa_tree_add_12_51_groupi_n_3169 ,csa_tree_add_12_51_groupi_n_1437 ,csa_tree_add_12_51_groupi_n_972);
  nor csa_tree_add_12_51_groupi_g18598(csa_tree_add_12_51_groupi_n_3168 ,csa_tree_add_12_51_groupi_n_1401 ,csa_tree_add_12_51_groupi_n_1058);
  nor csa_tree_add_12_51_groupi_g18599(csa_tree_add_12_51_groupi_n_3167 ,csa_tree_add_12_51_groupi_n_508 ,csa_tree_add_12_51_groupi_n_1068);
  nor csa_tree_add_12_51_groupi_g18600(csa_tree_add_12_51_groupi_n_3166 ,csa_tree_add_12_51_groupi_n_1463 ,csa_tree_add_12_51_groupi_n_1052);
  nor csa_tree_add_12_51_groupi_g18601(csa_tree_add_12_51_groupi_n_3165 ,csa_tree_add_12_51_groupi_n_622 ,csa_tree_add_12_51_groupi_n_1241);
  nor csa_tree_add_12_51_groupi_g18602(csa_tree_add_12_51_groupi_n_3164 ,csa_tree_add_12_51_groupi_n_502 ,csa_tree_add_12_51_groupi_n_703);
  nor csa_tree_add_12_51_groupi_g18603(csa_tree_add_12_51_groupi_n_3163 ,csa_tree_add_12_51_groupi_n_520 ,csa_tree_add_12_51_groupi_n_1332);
  nor csa_tree_add_12_51_groupi_g18604(csa_tree_add_12_51_groupi_n_3162 ,csa_tree_add_12_51_groupi_n_1452 ,csa_tree_add_12_51_groupi_n_932);
  nor csa_tree_add_12_51_groupi_g18605(csa_tree_add_12_51_groupi_n_3161 ,csa_tree_add_12_51_groupi_n_666 ,csa_tree_add_12_51_groupi_n_1109);
  nor csa_tree_add_12_51_groupi_g18606(csa_tree_add_12_51_groupi_n_3160 ,csa_tree_add_12_51_groupi_n_495 ,csa_tree_add_12_51_groupi_n_1052);
  nor csa_tree_add_12_51_groupi_g18607(csa_tree_add_12_51_groupi_n_3159 ,csa_tree_add_12_51_groupi_n_1424 ,csa_tree_add_12_51_groupi_n_1121);
  nor csa_tree_add_12_51_groupi_g18608(csa_tree_add_12_51_groupi_n_3158 ,csa_tree_add_12_51_groupi_n_1398 ,csa_tree_add_12_51_groupi_n_924);
  nor csa_tree_add_12_51_groupi_g18609(csa_tree_add_12_51_groupi_n_3157 ,csa_tree_add_12_51_groupi_n_643 ,csa_tree_add_12_51_groupi_n_1239);
  nor csa_tree_add_12_51_groupi_g18610(csa_tree_add_12_51_groupi_n_3156 ,csa_tree_add_12_51_groupi_n_1790 ,csa_tree_add_12_51_groupi_n_1058);
  nor csa_tree_add_12_51_groupi_g18611(csa_tree_add_12_51_groupi_n_3155 ,csa_tree_add_12_51_groupi_n_1446 ,csa_tree_add_12_51_groupi_n_706);
  nor csa_tree_add_12_51_groupi_g18612(csa_tree_add_12_51_groupi_n_3154 ,csa_tree_add_12_51_groupi_n_631 ,csa_tree_add_12_51_groupi_n_1106);
  nor csa_tree_add_12_51_groupi_g18613(csa_tree_add_12_51_groupi_n_3153 ,csa_tree_add_12_51_groupi_n_544 ,csa_tree_add_12_51_groupi_n_1244);
  nor csa_tree_add_12_51_groupi_g18614(csa_tree_add_12_51_groupi_n_3152 ,csa_tree_add_12_51_groupi_n_540 ,csa_tree_add_12_51_groupi_n_1323);
  nor csa_tree_add_12_51_groupi_g18615(csa_tree_add_12_51_groupi_n_3151 ,csa_tree_add_12_51_groupi_n_1760 ,csa_tree_add_12_51_groupi_n_1160);
  nor csa_tree_add_12_51_groupi_g18616(csa_tree_add_12_51_groupi_n_3150 ,csa_tree_add_12_51_groupi_n_1700 ,csa_tree_add_12_51_groupi_n_1280);
  nor csa_tree_add_12_51_groupi_g18617(csa_tree_add_12_51_groupi_n_3149 ,csa_tree_add_12_51_groupi_n_1763 ,csa_tree_add_12_51_groupi_n_896);
  nor csa_tree_add_12_51_groupi_g18618(csa_tree_add_12_51_groupi_n_3148 ,csa_tree_add_12_51_groupi_n_1434 ,csa_tree_add_12_51_groupi_n_1383);
  nor csa_tree_add_12_51_groupi_g18619(csa_tree_add_12_51_groupi_n_3147 ,csa_tree_add_12_51_groupi_n_633 ,csa_tree_add_12_51_groupi_n_1313);
  nor csa_tree_add_12_51_groupi_g18620(csa_tree_add_12_51_groupi_n_3146 ,csa_tree_add_12_51_groupi_n_687 ,csa_tree_add_12_51_groupi_n_1382);
  nor csa_tree_add_12_51_groupi_g18621(csa_tree_add_12_51_groupi_n_3145 ,csa_tree_add_12_51_groupi_n_534 ,csa_tree_add_12_51_groupi_n_1313);
  nor csa_tree_add_12_51_groupi_g18622(csa_tree_add_12_51_groupi_n_3144 ,csa_tree_add_12_51_groupi_n_487 ,csa_tree_add_12_51_groupi_n_891);
  nor csa_tree_add_12_51_groupi_g18623(csa_tree_add_12_51_groupi_n_3143 ,csa_tree_add_12_51_groupi_n_676 ,csa_tree_add_12_51_groupi_n_1245);
  nor csa_tree_add_12_51_groupi_g18624(csa_tree_add_12_51_groupi_n_3142 ,csa_tree_add_12_51_groupi_n_594 ,csa_tree_add_12_51_groupi_n_1187);
  nor csa_tree_add_12_51_groupi_g18625(csa_tree_add_12_51_groupi_n_3141 ,csa_tree_add_12_51_groupi_n_1785 ,csa_tree_add_12_51_groupi_n_1484);
  nor csa_tree_add_12_51_groupi_g18626(csa_tree_add_12_51_groupi_n_3140 ,csa_tree_add_12_51_groupi_n_645 ,csa_tree_add_12_51_groupi_n_1062);
  nor csa_tree_add_12_51_groupi_g18627(csa_tree_add_12_51_groupi_n_3139 ,csa_tree_add_12_51_groupi_n_685 ,csa_tree_add_12_51_groupi_n_1328);
  nor csa_tree_add_12_51_groupi_g18628(csa_tree_add_12_51_groupi_n_3138 ,csa_tree_add_12_51_groupi_n_597 ,csa_tree_add_12_51_groupi_n_1328);
  nor csa_tree_add_12_51_groupi_g18629(csa_tree_add_12_51_groupi_n_3137 ,csa_tree_add_12_51_groupi_n_1739 ,csa_tree_add_12_51_groupi_n_1098);
  nor csa_tree_add_12_51_groupi_g18630(csa_tree_add_12_51_groupi_n_3136 ,csa_tree_add_12_51_groupi_n_1787 ,csa_tree_add_12_51_groupi_n_1505);
  nor csa_tree_add_12_51_groupi_g18631(csa_tree_add_12_51_groupi_n_3135 ,csa_tree_add_12_51_groupi_n_655 ,csa_tree_add_12_51_groupi_n_1322);
  nor csa_tree_add_12_51_groupi_g18632(csa_tree_add_12_51_groupi_n_3134 ,csa_tree_add_12_51_groupi_n_1703 ,csa_tree_add_12_51_groupi_n_1493);
  nor csa_tree_add_12_51_groupi_g18633(csa_tree_add_12_51_groupi_n_3133 ,csa_tree_add_12_51_groupi_n_565 ,csa_tree_add_12_51_groupi_n_971);
  nor csa_tree_add_12_51_groupi_g18634(csa_tree_add_12_51_groupi_n_3132 ,csa_tree_add_12_51_groupi_n_490 ,csa_tree_add_12_51_groupi_n_1245);
  nor csa_tree_add_12_51_groupi_g18635(csa_tree_add_12_51_groupi_n_3131 ,csa_tree_add_12_51_groupi_n_576 ,csa_tree_add_12_51_groupi_n_951);
  nor csa_tree_add_12_51_groupi_g18636(csa_tree_add_12_51_groupi_n_3130 ,csa_tree_add_12_51_groupi_n_1097 ,csa_tree_add_12_51_groupi_n_250);
  nor csa_tree_add_12_51_groupi_g18637(csa_tree_add_12_51_groupi_n_3129 ,csa_tree_add_12_51_groupi_n_1530 ,csa_tree_add_12_51_groupi_n_247);
  nor csa_tree_add_12_51_groupi_g18638(csa_tree_add_12_51_groupi_n_3128 ,csa_tree_add_12_51_groupi_n_1113 ,csa_tree_add_12_51_groupi_n_394);
  nor csa_tree_add_12_51_groupi_g18639(csa_tree_add_12_51_groupi_n_3127 ,csa_tree_add_12_51_groupi_n_606 ,csa_tree_add_12_51_groupi_n_1277);
  nor csa_tree_add_12_51_groupi_g18640(csa_tree_add_12_51_groupi_n_3126 ,csa_tree_add_12_51_groupi_n_1796 ,csa_tree_add_12_51_groupi_n_1529);
  nor csa_tree_add_12_51_groupi_g18641(csa_tree_add_12_51_groupi_n_3125 ,csa_tree_add_12_51_groupi_n_1800 ,csa_tree_add_12_51_groupi_n_1242);
  nor csa_tree_add_12_51_groupi_g18642(csa_tree_add_12_51_groupi_n_3124 ,csa_tree_add_12_51_groupi_n_1299 ,csa_tree_add_12_51_groupi_n_235);
  nor csa_tree_add_12_51_groupi_g18643(csa_tree_add_12_51_groupi_n_3123 ,csa_tree_add_12_51_groupi_n_613 ,csa_tree_add_12_51_groupi_n_1556);
  nor csa_tree_add_12_51_groupi_g18644(csa_tree_add_12_51_groupi_n_3122 ,csa_tree_add_12_51_groupi_n_628 ,csa_tree_add_12_51_groupi_n_950);
  nor csa_tree_add_12_51_groupi_g18645(csa_tree_add_12_51_groupi_n_3121 ,csa_tree_add_12_51_groupi_n_1271 ,csa_tree_add_12_51_groupi_n_238);
  nor csa_tree_add_12_51_groupi_g18646(csa_tree_add_12_51_groupi_n_3120 ,csa_tree_add_12_51_groupi_n_1710 ,csa_tree_add_12_51_groupi_n_1229);
  nor csa_tree_add_12_51_groupi_g18647(csa_tree_add_12_51_groupi_n_3119 ,csa_tree_add_12_51_groupi_n_1722 ,csa_tree_add_12_51_groupi_n_1298);
  nor csa_tree_add_12_51_groupi_g18648(csa_tree_add_12_51_groupi_n_3118 ,csa_tree_add_12_51_groupi_n_618 ,csa_tree_add_12_51_groupi_n_1272);
  nor csa_tree_add_12_51_groupi_g18649(csa_tree_add_12_51_groupi_n_3117 ,csa_tree_add_12_51_groupi_n_1100 ,csa_tree_add_12_51_groupi_n_447);
  nor csa_tree_add_12_51_groupi_g18650(csa_tree_add_12_51_groupi_n_3116 ,csa_tree_add_12_51_groupi_n_1661 ,csa_tree_add_12_51_groupi_n_202);
  nor csa_tree_add_12_51_groupi_g18651(csa_tree_add_12_51_groupi_n_3115 ,csa_tree_add_12_51_groupi_n_601 ,csa_tree_add_12_51_groupi_n_1511);
  nor csa_tree_add_12_51_groupi_g18652(csa_tree_add_12_51_groupi_n_3114 ,csa_tree_add_12_51_groupi_n_1512 ,csa_tree_add_12_51_groupi_n_423);
  nor csa_tree_add_12_51_groupi_g18653(csa_tree_add_12_51_groupi_n_3113 ,csa_tree_add_12_51_groupi_n_1493 ,csa_tree_add_12_51_groupi_n_189);
  nor csa_tree_add_12_51_groupi_g18654(csa_tree_add_12_51_groupi_n_3112 ,csa_tree_add_12_51_groupi_n_609 ,csa_tree_add_12_51_groupi_n_1347);
  nor csa_tree_add_12_51_groupi_g18655(csa_tree_add_12_51_groupi_n_3111 ,csa_tree_add_12_51_groupi_n_592 ,csa_tree_add_12_51_groupi_n_1371);
  nor csa_tree_add_12_51_groupi_g18656(csa_tree_add_12_51_groupi_n_3110 ,csa_tree_add_12_51_groupi_n_1295 ,csa_tree_add_12_51_groupi_n_405);
  nor csa_tree_add_12_51_groupi_g18657(csa_tree_add_12_51_groupi_n_3109 ,csa_tree_add_12_51_groupi_n_1322 ,csa_tree_add_12_51_groupi_n_442);
  nor csa_tree_add_12_51_groupi_g18658(csa_tree_add_12_51_groupi_n_3108 ,csa_tree_add_12_51_groupi_n_1161 ,csa_tree_add_12_51_groupi_n_315);
  nor csa_tree_add_12_51_groupi_g18659(csa_tree_add_12_51_groupi_n_3107 ,csa_tree_add_12_51_groupi_n_624 ,csa_tree_add_12_51_groupi_n_1274);
  nor csa_tree_add_12_51_groupi_g18660(csa_tree_add_12_51_groupi_n_3106 ,csa_tree_add_12_51_groupi_n_1752 ,csa_tree_add_12_51_groupi_n_953);
  nor csa_tree_add_12_51_groupi_g18661(csa_tree_add_12_51_groupi_n_3105 ,csa_tree_add_12_51_groupi_n_1755 ,csa_tree_add_12_51_groupi_n_1161);
  nor csa_tree_add_12_51_groupi_g18662(csa_tree_add_12_51_groupi_n_3104 ,csa_tree_add_12_51_groupi_n_562 ,csa_tree_add_12_51_groupi_n_932);
  nor csa_tree_add_12_51_groupi_g18663(csa_tree_add_12_51_groupi_n_3103 ,csa_tree_add_12_51_groupi_n_1329 ,csa_tree_add_12_51_groupi_n_333);
  nor csa_tree_add_12_51_groupi_g18664(csa_tree_add_12_51_groupi_n_3102 ,csa_tree_add_12_51_groupi_n_1106 ,csa_tree_add_12_51_groupi_n_331);
  nor csa_tree_add_12_51_groupi_g18665(csa_tree_add_12_51_groupi_n_3101 ,csa_tree_add_12_51_groupi_n_1506 ,csa_tree_add_12_51_groupi_n_183);
  nor csa_tree_add_12_51_groupi_g18666(csa_tree_add_12_51_groupi_n_3100 ,csa_tree_add_12_51_groupi_n_1514 ,csa_tree_add_12_51_groupi_n_460);
  nor csa_tree_add_12_51_groupi_g18667(csa_tree_add_12_51_groupi_n_3099 ,csa_tree_add_12_51_groupi_n_1460 ,csa_tree_add_12_51_groupi_n_1107);
  nor csa_tree_add_12_51_groupi_g18668(csa_tree_add_12_51_groupi_n_3098 ,csa_tree_add_12_51_groupi_n_1511 ,csa_tree_add_12_51_groupi_n_286);
  nor csa_tree_add_12_51_groupi_g18669(csa_tree_add_12_51_groupi_n_3097 ,csa_tree_add_12_51_groupi_n_603 ,csa_tree_add_12_51_groupi_n_1184);
  nor csa_tree_add_12_51_groupi_g18670(csa_tree_add_12_51_groupi_n_3096 ,csa_tree_add_12_51_groupi_n_1314 ,csa_tree_add_12_51_groupi_n_348);
  nor csa_tree_add_12_51_groupi_g18671(csa_tree_add_12_51_groupi_n_3095 ,csa_tree_add_12_51_groupi_n_1346 ,csa_tree_add_12_51_groupi_n_240);
  nor csa_tree_add_12_51_groupi_g18672(csa_tree_add_12_51_groupi_n_3094 ,csa_tree_add_12_51_groupi_n_1347 ,csa_tree_add_12_51_groupi_n_472);
  nor csa_tree_add_12_51_groupi_g18673(csa_tree_add_12_51_groupi_n_3093 ,csa_tree_add_12_51_groupi_n_1731 ,csa_tree_add_12_51_groupi_n_1295);
  nor csa_tree_add_12_51_groupi_g18674(csa_tree_add_12_51_groupi_n_3092 ,csa_tree_add_12_51_groupi_n_1464 ,csa_tree_add_12_51_groupi_n_1370);
  nor csa_tree_add_12_51_groupi_g18675(csa_tree_add_12_51_groupi_n_3091 ,csa_tree_add_12_51_groupi_n_1776 ,csa_tree_add_12_51_groupi_n_1188);
  nor csa_tree_add_12_51_groupi_g18676(csa_tree_add_12_51_groupi_n_3090 ,csa_tree_add_12_51_groupi_n_1478 ,csa_tree_add_12_51_groupi_n_195);
  nor csa_tree_add_12_51_groupi_g18677(csa_tree_add_12_51_groupi_n_3089 ,csa_tree_add_12_51_groupi_n_507 ,csa_tree_add_12_51_groupi_n_897);
  nor csa_tree_add_12_51_groupi_g18678(csa_tree_add_12_51_groupi_n_3088 ,csa_tree_add_12_51_groupi_n_1401 ,csa_tree_add_12_51_groupi_n_1101);
  nor csa_tree_add_12_51_groupi_g18679(csa_tree_add_12_51_groupi_n_3087 ,csa_tree_add_12_51_groupi_n_1793 ,csa_tree_add_12_51_groupi_n_1185);
  nor csa_tree_add_12_51_groupi_g18680(csa_tree_add_12_51_groupi_n_3086 ,csa_tree_add_12_51_groupi_n_1514 ,csa_tree_add_12_51_groupi_n_475);
  nor csa_tree_add_12_51_groupi_g18681(csa_tree_add_12_51_groupi_n_3085 ,csa_tree_add_12_51_groupi_n_1382 ,csa_tree_add_12_51_groupi_n_477);
  nor csa_tree_add_12_51_groupi_g18682(csa_tree_add_12_51_groupi_n_3084 ,csa_tree_add_12_51_groupi_n_88 ,csa_tree_add_12_51_groupi_n_852);
  nor csa_tree_add_12_51_groupi_g18683(csa_tree_add_12_51_groupi_n_3083 ,csa_tree_add_12_51_groupi_n_1185 ,csa_tree_add_12_51_groupi_n_261);
  nor csa_tree_add_12_51_groupi_g18684(csa_tree_add_12_51_groupi_n_3082 ,csa_tree_add_12_51_groupi_n_1056 ,csa_tree_add_12_51_groupi_n_417);
  nor csa_tree_add_12_51_groupi_g18685(csa_tree_add_12_51_groupi_n_3081 ,csa_tree_add_12_51_groupi_n_1472 ,csa_tree_add_12_51_groupi_n_1163);
  nor csa_tree_add_12_51_groupi_g18686(csa_tree_add_12_51_groupi_n_3080 ,csa_tree_add_12_51_groupi_n_1808 ,csa_tree_add_12_51_groupi_n_1122);
  nor csa_tree_add_12_51_groupi_g18687(csa_tree_add_12_51_groupi_n_3079 ,csa_tree_add_12_51_groupi_n_669 ,csa_tree_add_12_51_groupi_n_1101);
  nor csa_tree_add_12_51_groupi_g18688(csa_tree_add_12_51_groupi_n_3078 ,csa_tree_add_12_51_groupi_n_1661 ,csa_tree_add_12_51_groupi_n_222);
  nor csa_tree_add_12_51_groupi_g18689(csa_tree_add_12_51_groupi_n_3077 ,csa_tree_add_12_51_groupi_n_1371 ,csa_tree_add_12_51_groupi_n_382);
  nor csa_tree_add_12_51_groupi_g18690(csa_tree_add_12_51_groupi_n_3076 ,csa_tree_add_12_51_groupi_n_1425 ,csa_tree_add_12_51_groupi_n_891);
  nor csa_tree_add_12_51_groupi_g18691(csa_tree_add_12_51_groupi_n_3075 ,csa_tree_add_12_51_groupi_n_1505 ,csa_tree_add_12_51_groupi_n_367);
  nor csa_tree_add_12_51_groupi_g18692(csa_tree_add_12_51_groupi_n_3074 ,csa_tree_add_12_51_groupi_n_502 ,csa_tree_add_12_51_groupi_n_951);
  nor csa_tree_add_12_51_groupi_g18693(csa_tree_add_12_51_groupi_n_3073 ,csa_tree_add_12_51_groupi_n_1662 ,csa_tree_add_12_51_groupi_n_213);
  nor csa_tree_add_12_51_groupi_g18694(csa_tree_add_12_51_groupi_n_3072 ,csa_tree_add_12_51_groupi_n_1380 ,csa_tree_add_12_51_groupi_n_388);
  nor csa_tree_add_12_51_groupi_g18695(csa_tree_add_12_51_groupi_n_3071 ,csa_tree_add_12_51_groupi_n_672 ,csa_tree_add_12_51_groupi_n_1113);
  nor csa_tree_add_12_51_groupi_g18696(csa_tree_add_12_51_groupi_n_3070 ,csa_tree_add_12_51_groupi_n_651 ,csa_tree_add_12_51_groupi_n_1067);
  nor csa_tree_add_12_51_groupi_g18697(csa_tree_add_12_51_groupi_n_3069 ,csa_tree_add_12_51_groupi_n_1379 ,csa_tree_add_12_51_groupi_n_444);
  nor csa_tree_add_12_51_groupi_g18698(csa_tree_add_12_51_groupi_n_3068 ,csa_tree_add_12_51_groupi_n_1370 ,csa_tree_add_12_51_groupi_n_439);
  nor csa_tree_add_12_51_groupi_g18699(csa_tree_add_12_51_groupi_n_3067 ,csa_tree_add_12_51_groupi_n_1719 ,csa_tree_add_12_51_groupi_n_1296);
  nor csa_tree_add_12_51_groupi_g18700(csa_tree_add_12_51_groupi_n_3066 ,csa_tree_add_12_51_groupi_n_688 ,csa_tree_add_12_51_groupi_n_1232);
  nor csa_tree_add_12_51_groupi_g18701(csa_tree_add_12_51_groupi_n_3065 ,csa_tree_add_12_51_groupi_n_510 ,csa_tree_add_12_51_groupi_n_1184);
  nor csa_tree_add_12_51_groupi_g18702(csa_tree_add_12_51_groupi_n_3064 ,csa_tree_add_12_51_groupi_n_1742 ,csa_tree_add_12_51_groupi_n_1271);
  nor csa_tree_add_12_51_groupi_g18703(csa_tree_add_12_51_groupi_n_3063 ,csa_tree_add_12_51_groupi_n_1748 ,csa_tree_add_12_51_groupi_n_1275);
  nor csa_tree_add_12_51_groupi_g18704(csa_tree_add_12_51_groupi_n_3062 ,csa_tree_add_12_51_groupi_n_1745 ,csa_tree_add_12_51_groupi_n_1112);
  nor csa_tree_add_12_51_groupi_g18705(csa_tree_add_12_51_groupi_n_3061 ,csa_tree_add_12_51_groupi_n_1458 ,csa_tree_add_12_51_groupi_n_954);
  nor csa_tree_add_12_51_groupi_g18706(csa_tree_add_12_51_groupi_n_3060 ,csa_tree_add_12_51_groupi_n_564 ,csa_tree_add_12_51_groupi_n_1164);
  nor csa_tree_add_12_51_groupi_g18707(csa_tree_add_12_51_groupi_n_3059 ,csa_tree_add_12_51_groupi_n_1494 ,csa_tree_add_12_51_groupi_n_268);
  nor csa_tree_add_12_51_groupi_g18708(csa_tree_add_12_51_groupi_n_3058 ,csa_tree_add_12_51_groupi_n_522 ,csa_tree_add_12_51_groupi_n_706);
  nor csa_tree_add_12_51_groupi_g18709(csa_tree_add_12_51_groupi_n_3057 ,csa_tree_add_12_51_groupi_n_1811 ,csa_tree_add_12_51_groupi_n_1238);
  nor csa_tree_add_12_51_groupi_g18710(csa_tree_add_12_51_groupi_n_3056 ,csa_tree_add_12_51_groupi_n_1452 ,csa_tree_add_12_51_groupi_n_1112);
  nor csa_tree_add_12_51_groupi_g18711(csa_tree_add_12_51_groupi_n_3055 ,csa_tree_add_12_51_groupi_n_1316 ,csa_tree_add_12_51_groupi_n_427);
  nor csa_tree_add_12_51_groupi_g18712(csa_tree_add_12_51_groupi_n_3054 ,csa_tree_add_12_51_groupi_n_1778 ,csa_tree_add_12_51_groupi_n_972);
  nor csa_tree_add_12_51_groupi_g18713(csa_tree_add_12_51_groupi_n_3053 ,csa_tree_add_12_51_groupi_n_516 ,csa_tree_add_12_51_groupi_n_1478);
  nor csa_tree_add_12_51_groupi_g18714(csa_tree_add_12_51_groupi_n_3052 ,csa_tree_add_12_51_groupi_n_1437 ,csa_tree_add_12_51_groupi_n_1298);
  nor csa_tree_add_12_51_groupi_g18715(csa_tree_add_12_51_groupi_n_3051 ,csa_tree_add_12_51_groupi_n_1557 ,csa_tree_add_12_51_groupi_n_378);
  nor csa_tree_add_12_51_groupi_g18716(csa_tree_add_12_51_groupi_n_3050 ,csa_tree_add_12_51_groupi_n_1329 ,csa_tree_add_12_51_groupi_n_415);
  nor csa_tree_add_12_51_groupi_g18717(csa_tree_add_12_51_groupi_n_3049 ,csa_tree_add_12_51_groupi_n_1331 ,csa_tree_add_12_51_groupi_n_339);
  nor csa_tree_add_12_51_groupi_g18718(csa_tree_add_12_51_groupi_n_3048 ,csa_tree_add_12_51_groupi_n_690 ,csa_tree_add_12_51_groupi_n_1230);
  nor csa_tree_add_12_51_groupi_g18719(csa_tree_add_12_51_groupi_n_3047 ,csa_tree_add_12_51_groupi_n_1482 ,csa_tree_add_12_51_groupi_n_273);
  nor csa_tree_add_12_51_groupi_g18720(csa_tree_add_12_51_groupi_n_3046 ,csa_tree_add_12_51_groupi_n_1442 ,csa_tree_add_12_51_groupi_n_703);
  nor csa_tree_add_12_51_groupi_g18721(csa_tree_add_12_51_groupi_n_3045 ,csa_tree_add_12_51_groupi_n_1367 ,csa_tree_add_12_51_groupi_n_280);
  nor csa_tree_add_12_51_groupi_g18722(csa_tree_add_12_51_groupi_n_3044 ,csa_tree_add_12_51_groupi_n_1407 ,csa_tree_add_12_51_groupi_n_882);
  nor csa_tree_add_12_51_groupi_g18723(csa_tree_add_12_51_groupi_n_3043 ,csa_tree_add_12_51_groupi_n_1419 ,csa_tree_add_12_51_groupi_n_1238);
  nor csa_tree_add_12_51_groupi_g18724(csa_tree_add_12_51_groupi_n_3042 ,csa_tree_add_12_51_groupi_n_1769 ,csa_tree_add_12_51_groupi_n_953);
  nor csa_tree_add_12_51_groupi_g18725(csa_tree_add_12_51_groupi_n_3041 ,csa_tree_add_12_51_groupi_n_1790 ,csa_tree_add_12_51_groupi_n_1056);
  nor csa_tree_add_12_51_groupi_g18726(csa_tree_add_12_51_groupi_n_3040 ,csa_tree_add_12_51_groupi_n_1484 ,csa_tree_add_12_51_groupi_n_454);
  nor csa_tree_add_12_51_groupi_g18727(csa_tree_add_12_51_groupi_n_3039 ,csa_tree_add_12_51_groupi_n_654 ,csa_tree_add_12_51_groupi_n_1367);
  nor csa_tree_add_12_51_groupi_g18728(csa_tree_add_12_51_groupi_n_3038 ,csa_tree_add_12_51_groupi_n_1274 ,csa_tree_add_12_51_groupi_n_448);
  nor csa_tree_add_12_51_groupi_g18729(csa_tree_add_12_51_groupi_n_3037 ,csa_tree_add_12_51_groupi_n_1694 ,csa_tree_add_12_51_groupi_n_1061);
  nor csa_tree_add_12_51_groupi_g18730(csa_tree_add_12_51_groupi_n_3036 ,csa_tree_add_12_51_groupi_n_1781 ,csa_tree_add_12_51_groupi_n_1160);
  nor csa_tree_add_12_51_groupi_g18731(csa_tree_add_12_51_groupi_n_3035 ,csa_tree_add_12_51_groupi_n_905 ,csa_tree_add_12_51_groupi_n_370);
  nor csa_tree_add_12_51_groupi_g18732(csa_tree_add_12_51_groupi_n_3034 ,csa_tree_add_12_51_groupi_n_588 ,csa_tree_add_12_51_groupi_n_1331);
  nor csa_tree_add_12_51_groupi_g18733(csa_tree_add_12_51_groupi_n_3033 ,csa_tree_add_12_51_groupi_n_1416 ,csa_tree_add_12_51_groupi_n_1377);
  nor csa_tree_add_12_51_groupi_g18734(csa_tree_add_12_51_groupi_n_3032 ,csa_tree_add_12_51_groupi_n_639 ,csa_tree_add_12_51_groupi_n_1380);
  nor csa_tree_add_12_51_groupi_g18735(csa_tree_add_12_51_groupi_n_3031 ,csa_tree_add_12_51_groupi_n_661 ,csa_tree_add_12_51_groupi_n_933);
  nor csa_tree_add_12_51_groupi_g18736(csa_tree_add_12_51_groupi_n_3030 ,csa_tree_add_12_51_groupi_n_642 ,csa_tree_add_12_51_groupi_n_890);
  nor csa_tree_add_12_51_groupi_g18737(csa_tree_add_12_51_groupi_n_3029 ,csa_tree_add_12_51_groupi_n_591 ,csa_tree_add_12_51_groupi_n_1368);
  nor csa_tree_add_12_51_groupi_g18738(csa_tree_add_12_51_groupi_n_3028 ,csa_tree_add_12_51_groupi_n_1409 ,csa_tree_add_12_51_groupi_n_974);
  nor csa_tree_add_12_51_groupi_g18739(csa_tree_add_12_51_groupi_n_3027 ,csa_tree_add_12_51_groupi_n_1724 ,csa_tree_add_12_51_groupi_n_1232);
  nor csa_tree_add_12_51_groupi_g18740(csa_tree_add_12_51_groupi_n_3026 ,csa_tree_add_12_51_groupi_n_1727 ,csa_tree_add_12_51_groupi_n_974);
  nor csa_tree_add_12_51_groupi_g18741(csa_tree_add_12_51_groupi_n_3025 ,csa_tree_add_12_51_groupi_n_1529 ,csa_tree_add_12_51_groupi_n_292);
  nor csa_tree_add_12_51_groupi_g18742(csa_tree_add_12_51_groupi_n_3024 ,csa_tree_add_12_51_groupi_n_489 ,csa_tree_add_12_51_groupi_n_906);
  nor csa_tree_add_12_51_groupi_g18743(csa_tree_add_12_51_groupi_n_3023 ,csa_tree_add_12_51_groupi_n_1712 ,csa_tree_add_12_51_groupi_n_1110);
  nor csa_tree_add_12_51_groupi_g18744(csa_tree_add_12_51_groupi_n_3022 ,csa_tree_add_12_51_groupi_n_487 ,csa_tree_add_12_51_groupi_n_1059);
  nor csa_tree_add_12_51_groupi_g18745(csa_tree_add_12_51_groupi_n_3021 ,csa_tree_add_12_51_groupi_n_1706 ,csa_tree_add_12_51_groupi_n_1316);
  nor csa_tree_add_12_51_groupi_g18746(csa_tree_add_12_51_groupi_n_3020 ,csa_tree_add_12_51_groupi_n_1440 ,csa_tree_add_12_51_groupi_n_1376);
  nor csa_tree_add_12_51_groupi_g18747(csa_tree_add_12_51_groupi_n_3019 ,csa_tree_add_12_51_groupi_n_1278 ,csa_tree_add_12_51_groupi_n_432);
  nor csa_tree_add_12_51_groupi_g18748(csa_tree_add_12_51_groupi_n_3018 ,csa_tree_add_12_51_groupi_n_1697 ,csa_tree_add_12_51_groupi_n_1121);
  nor csa_tree_add_12_51_groupi_g18749(csa_tree_add_12_51_groupi_n_3017 ,csa_tree_add_12_51_groupi_n_1772 ,csa_tree_add_12_51_groupi_n_1317);
  nor csa_tree_add_12_51_groupi_g18750(csa_tree_add_12_51_groupi_n_3016 ,csa_tree_add_12_51_groupi_n_1061 ,csa_tree_add_12_51_groupi_n_313);
  nor csa_tree_add_12_51_groupi_g18751(csa_tree_add_12_51_groupi_n_3015 ,csa_tree_add_12_51_groupi_n_1422 ,csa_tree_add_12_51_groupi_n_1062);
  nor csa_tree_add_12_51_groupi_g18752(csa_tree_add_12_51_groupi_n_3014 ,csa_tree_add_12_51_groupi_n_600 ,csa_tree_add_12_51_groupi_n_1053);
  nor csa_tree_add_12_51_groupi_g18753(csa_tree_add_12_51_groupi_n_3013 ,csa_tree_add_12_51_groupi_n_1733 ,csa_tree_add_12_51_groupi_n_975);
  nor csa_tree_add_12_51_groupi_g18754(csa_tree_add_12_51_groupi_n_3012 ,csa_tree_add_12_51_groupi_n_1715 ,csa_tree_add_12_51_groupi_n_1055);
  nor csa_tree_add_12_51_groupi_g18755(csa_tree_add_12_51_groupi_n_3011 ,csa_tree_add_12_51_groupi_n_1317 ,csa_tree_add_12_51_groupi_n_262);
  nor csa_tree_add_12_51_groupi_g18756(csa_tree_add_12_51_groupi_n_3010 ,csa_tree_add_12_51_groupi_n_561 ,csa_tree_add_12_51_groupi_n_1097);
  nor csa_tree_add_12_51_groupi_g18757(csa_tree_add_12_51_groupi_n_3009 ,csa_tree_add_12_51_groupi_n_1556 ,csa_tree_add_12_51_groupi_n_282);
  nor csa_tree_add_12_51_groupi_g18758(csa_tree_add_12_51_groupi_n_3008 ,csa_tree_add_12_51_groupi_n_630 ,csa_tree_add_12_51_groupi_n_1229);
  nor csa_tree_add_12_51_groupi_g18759(csa_tree_add_12_51_groupi_n_3007 ,csa_tree_add_12_51_groupi_n_555 ,csa_tree_add_12_51_groupi_n_1379);
  nor csa_tree_add_12_51_groupi_g18760(csa_tree_add_12_51_groupi_n_3006 ,csa_tree_add_12_51_groupi_n_543 ,csa_tree_add_12_51_groupi_n_881);
  nor csa_tree_add_12_51_groupi_g18761(csa_tree_add_12_51_groupi_n_3005 ,csa_tree_add_12_51_groupi_n_1736 ,csa_tree_add_12_51_groupi_n_1110);
  nor csa_tree_add_12_51_groupi_g18762(csa_tree_add_12_51_groupi_n_3004 ,csa_tree_add_12_51_groupi_n_1703 ,csa_tree_add_12_51_groupi_n_950);
  nor csa_tree_add_12_51_groupi_g18763(csa_tree_add_12_51_groupi_n_3003 ,csa_tree_add_12_51_groupi_n_1565 ,csa_tree_add_12_51_groupi_n_1532);
  nor csa_tree_add_12_51_groupi_g18764(csa_tree_add_12_51_groupi_n_3002 ,csa_tree_add_12_51_groupi_n_1757 ,csa_tree_add_12_51_groupi_n_1278);
  nor csa_tree_add_12_51_groupi_g18765(csa_tree_add_12_51_groupi_n_3001 ,csa_tree_add_12_51_groupi_n_513 ,csa_tree_add_12_51_groupi_n_971);
  nor csa_tree_add_12_51_groupi_g18766(csa_tree_add_12_51_groupi_n_3000 ,csa_tree_add_12_51_groupi_n_1482 ,csa_tree_add_12_51_groupi_n_271);
  nor csa_tree_add_12_51_groupi_g18767(csa_tree_add_12_51_groupi_n_2999 ,csa_tree_add_12_51_groupi_n_1109 ,csa_tree_add_12_51_groupi_n_246);
  nor csa_tree_add_12_51_groupi_g18768(csa_tree_add_12_51_groupi_n_2998 ,csa_tree_add_12_51_groupi_n_1740 ,csa_tree_add_12_51_groupi_n_923);
  nor csa_tree_add_12_51_groupi_g18769(csa_tree_add_12_51_groupi_n_2997 ,csa_tree_add_12_51_groupi_n_1766 ,csa_tree_add_12_51_groupi_n_1281);
  nor csa_tree_add_12_51_groupi_g18770(csa_tree_add_12_51_groupi_n_2996 ,csa_tree_add_12_51_groupi_n_1053 ,csa_tree_add_12_51_groupi_n_469);
  nor csa_tree_add_12_51_groupi_g18771(csa_tree_add_12_51_groupi_n_2995 ,csa_tree_add_12_51_groupi_n_1760 ,csa_tree_add_12_51_groupi_n_1098);
  nor csa_tree_add_12_51_groupi_g18772(csa_tree_add_12_51_groupi_n_2994 ,csa_tree_add_12_51_groupi_n_1277 ,csa_tree_add_12_51_groupi_n_352);
  nor csa_tree_add_12_51_groupi_g18773(csa_tree_add_12_51_groupi_n_2993 ,csa_tree_add_12_51_groupi_n_1280 ,csa_tree_add_12_51_groupi_n_391);
  nor csa_tree_add_12_51_groupi_g18774(csa_tree_add_12_51_groupi_n_2992 ,csa_tree_add_12_51_groupi_n_1532 ,csa_tree_add_12_51_groupi_n_238);
  nor csa_tree_add_12_51_groupi_g18775(csa_tree_add_12_51_groupi_n_2991 ,csa_tree_add_12_51_groupi_n_1763 ,csa_tree_add_12_51_groupi_n_881);
  nor csa_tree_add_12_51_groupi_g18776(csa_tree_add_12_51_groupi_n_2990 ,csa_tree_add_12_51_groupi_n_1533 ,csa_tree_add_12_51_groupi_n_367);
  nor csa_tree_add_12_51_groupi_g18777(csa_tree_add_12_51_groupi_n_2989 ,csa_tree_add_12_51_groupi_n_1530 ,csa_tree_add_12_51_groupi_n_196);
  nor csa_tree_add_12_51_groupi_g18778(csa_tree_add_12_51_groupi_n_2988 ,csa_tree_add_12_51_groupi_n_1376 ,csa_tree_add_12_51_groupi_n_412);
  nor csa_tree_add_12_51_groupi_g18779(csa_tree_add_12_51_groupi_n_2987 ,csa_tree_add_12_51_groupi_n_1485 ,csa_tree_add_12_51_groupi_n_388);
  nor csa_tree_add_12_51_groupi_g18780(csa_tree_add_12_51_groupi_n_2986 ,csa_tree_add_12_51_groupi_n_1494 ,csa_tree_add_12_51_groupi_n_400);
  nor csa_tree_add_12_51_groupi_g18781(csa_tree_add_12_51_groupi_n_2985 ,csa_tree_add_12_51_groupi_n_1067 ,csa_tree_add_12_51_groupi_n_394);
  nor csa_tree_add_12_51_groupi_g18782(csa_tree_add_12_51_groupi_n_2984 ,csa_tree_add_12_51_groupi_n_1332 ,csa_tree_add_12_51_groupi_n_265);
  nor csa_tree_add_12_51_groupi_g18783(csa_tree_add_12_51_groupi_n_2983 ,csa_tree_add_12_51_groupi_n_1481 ,csa_tree_add_12_51_groupi_n_474);
  nor csa_tree_add_12_51_groupi_g18784(csa_tree_add_12_51_groupi_n_2982 ,csa_tree_add_12_51_groupi_n_1479 ,csa_tree_add_12_51_groupi_n_187);
  nor csa_tree_add_12_51_groupi_g18785(csa_tree_add_12_51_groupi_n_2981 ,csa_tree_add_12_51_groupi_n_1485 ,csa_tree_add_12_51_groupi_n_223);
  nor csa_tree_add_12_51_groupi_g18786(csa_tree_add_12_51_groupi_n_2980 ,csa_tree_add_12_51_groupi_n_1059 ,csa_tree_add_12_51_groupi_n_244);
  nor csa_tree_add_12_51_groupi_g18787(csa_tree_add_12_51_groupi_n_2979 ,csa_tree_add_12_51_groupi_n_1296 ,csa_tree_add_12_51_groupi_n_358);
  and csa_tree_add_12_51_groupi_g18788(csa_tree_add_12_51_groupi_n_2978 ,csa_tree_add_12_51_groupi_n_46 ,csa_tree_add_12_51_groupi_n_938);
  and csa_tree_add_12_51_groupi_g18789(csa_tree_add_12_51_groupi_n_2977 ,csa_tree_add_12_51_groupi_n_40 ,csa_tree_add_12_51_groupi_n_920);
  and csa_tree_add_12_51_groupi_g18790(csa_tree_add_12_51_groupi_n_2976 ,csa_tree_add_12_51_groupi_n_49 ,csa_tree_add_12_51_groupi_n_1190);
  and csa_tree_add_12_51_groupi_g18791(csa_tree_add_12_51_groupi_n_2975 ,csa_tree_add_12_51_groupi_n_52 ,csa_tree_add_12_51_groupi_n_917);
  and csa_tree_add_12_51_groupi_g18792(csa_tree_add_12_51_groupi_n_2974 ,csa_tree_add_12_51_groupi_n_61 ,csa_tree_add_12_51_groupi_n_863);
  and csa_tree_add_12_51_groupi_g18793(csa_tree_add_12_51_groupi_n_2973 ,csa_tree_add_12_51_groupi_n_22 ,csa_tree_add_12_51_groupi_n_1253);
  and csa_tree_add_12_51_groupi_g18794(csa_tree_add_12_51_groupi_n_2972 ,csa_tree_add_12_51_groupi_n_25 ,csa_tree_add_12_51_groupi_n_1292);
  and csa_tree_add_12_51_groupi_g18795(csa_tree_add_12_51_groupi_n_2971 ,csa_tree_add_12_51_groupi_n_34 ,csa_tree_add_12_51_groupi_n_911);
  and csa_tree_add_12_51_groupi_g18796(csa_tree_add_12_51_groupi_n_2970 ,csa_tree_add_12_51_groupi_n_58 ,csa_tree_add_12_51_groupi_n_1202);
  and csa_tree_add_12_51_groupi_g18797(csa_tree_add_12_51_groupi_n_2969 ,csa_tree_add_12_51_groupi_n_55 ,csa_tree_add_12_51_groupi_n_1208);
  and csa_tree_add_12_51_groupi_g18798(csa_tree_add_12_51_groupi_n_2968 ,csa_tree_add_12_51_groupi_n_64 ,csa_tree_add_12_51_groupi_n_1304);
  and csa_tree_add_12_51_groupi_g18799(csa_tree_add_12_51_groupi_n_2967 ,csa_tree_add_12_51_groupi_n_31 ,csa_tree_add_12_51_groupi_n_1118);
  nor csa_tree_add_12_51_groupi_g18800(csa_tree_add_12_51_groupi_n_2966 ,csa_tree_add_12_51_groupi_n_68 ,csa_tree_add_12_51_groupi_n_837);
  nor csa_tree_add_12_51_groupi_g18801(csa_tree_add_12_51_groupi_n_2965 ,csa_tree_add_12_51_groupi_n_74 ,csa_tree_add_12_51_groupi_n_834);
  nor csa_tree_add_12_51_groupi_g18802(csa_tree_add_12_51_groupi_n_2964 ,csa_tree_add_12_51_groupi_n_80 ,csa_tree_add_12_51_groupi_n_851);
  nor csa_tree_add_12_51_groupi_g18803(csa_tree_add_12_51_groupi_n_2963 ,csa_tree_add_12_51_groupi_n_84 ,csa_tree_add_12_51_groupi_n_167);
  nor csa_tree_add_12_51_groupi_g18804(csa_tree_add_12_51_groupi_n_2962 ,csa_tree_add_12_51_groupi_n_94 ,csa_tree_add_12_51_groupi_n_851);
  or csa_tree_add_12_51_groupi_g18805(csa_tree_add_12_51_groupi_n_3255 ,csa_tree_add_12_51_groupi_n_2588 ,csa_tree_add_12_51_groupi_n_2784);
  or csa_tree_add_12_51_groupi_g18806(csa_tree_add_12_51_groupi_n_3254 ,csa_tree_add_12_51_groupi_n_2587 ,csa_tree_add_12_51_groupi_n_2799);
  or csa_tree_add_12_51_groupi_g18807(csa_tree_add_12_51_groupi_n_3253 ,csa_tree_add_12_51_groupi_n_2585 ,csa_tree_add_12_51_groupi_n_2793);
  or csa_tree_add_12_51_groupi_g18808(csa_tree_add_12_51_groupi_n_3252 ,csa_tree_add_12_51_groupi_n_2614 ,csa_tree_add_12_51_groupi_n_2796);
  or csa_tree_add_12_51_groupi_g18809(csa_tree_add_12_51_groupi_n_3251 ,csa_tree_add_12_51_groupi_n_2702 ,csa_tree_add_12_51_groupi_n_2807);
  or csa_tree_add_12_51_groupi_g18810(csa_tree_add_12_51_groupi_n_3250 ,csa_tree_add_12_51_groupi_n_2717 ,csa_tree_add_12_51_groupi_n_2806);
  or csa_tree_add_12_51_groupi_g18811(csa_tree_add_12_51_groupi_n_3249 ,csa_tree_add_12_51_groupi_n_2575 ,csa_tree_add_12_51_groupi_n_2801);
  or csa_tree_add_12_51_groupi_g18812(csa_tree_add_12_51_groupi_n_3248 ,csa_tree_add_12_51_groupi_n_2616 ,csa_tree_add_12_51_groupi_n_2811);
  or csa_tree_add_12_51_groupi_g18813(csa_tree_add_12_51_groupi_n_3247 ,csa_tree_add_12_51_groupi_n_2583 ,csa_tree_add_12_51_groupi_n_2785);
  or csa_tree_add_12_51_groupi_g18814(csa_tree_add_12_51_groupi_n_3246 ,csa_tree_add_12_51_groupi_n_2901 ,csa_tree_add_12_51_groupi_n_2351);
  xnor csa_tree_add_12_51_groupi_g18815(csa_tree_add_12_51_groupi_n_3245 ,csa_tree_add_12_51_groupi_n_2572 ,in2[14]);
  xnor csa_tree_add_12_51_groupi_g18816(csa_tree_add_12_51_groupi_n_3244 ,csa_tree_add_12_51_groupi_n_2553 ,in2[5]);
  xnor csa_tree_add_12_51_groupi_g18817(csa_tree_add_12_51_groupi_n_3243 ,csa_tree_add_12_51_groupi_n_2554 ,in4[11]);
  xnor csa_tree_add_12_51_groupi_g18818(csa_tree_add_12_51_groupi_n_3242 ,csa_tree_add_12_51_groupi_n_2552 ,in4[2]);
  xnor csa_tree_add_12_51_groupi_g18819(csa_tree_add_12_51_groupi_n_3241 ,csa_tree_add_12_51_groupi_n_2573 ,in3[8]);
  xnor csa_tree_add_12_51_groupi_g18820(csa_tree_add_12_51_groupi_n_3239 ,csa_tree_add_12_51_groupi_n_2361 ,csa_tree_add_12_51_groupi_n_2551);
  xnor csa_tree_add_12_51_groupi_g18821(csa_tree_add_12_51_groupi_n_3237 ,csa_tree_add_12_51_groupi_n_1916 ,csa_tree_add_12_51_groupi_n_2571);
  xnor csa_tree_add_12_51_groupi_g18822(csa_tree_add_12_51_groupi_n_3235 ,csa_tree_add_12_51_groupi_n_1944 ,csa_tree_add_12_51_groupi_n_2556);
  xnor csa_tree_add_12_51_groupi_g18823(csa_tree_add_12_51_groupi_n_3234 ,csa_tree_add_12_51_groupi_n_2555 ,in2[5]);
  or csa_tree_add_12_51_groupi_g18824(csa_tree_add_12_51_groupi_n_3232 ,csa_tree_add_12_51_groupi_n_2630 ,csa_tree_add_12_51_groupi_n_2791);
  or csa_tree_add_12_51_groupi_g18825(csa_tree_add_12_51_groupi_n_3230 ,csa_tree_add_12_51_groupi_n_2591 ,csa_tree_add_12_51_groupi_n_2804);
  xnor csa_tree_add_12_51_groupi_g18826(csa_tree_add_12_51_groupi_n_3229 ,csa_tree_add_12_51_groupi_n_2467 ,csa_tree_add_12_51_groupi_n_2565);
  not csa_tree_add_12_51_groupi_g18827(csa_tree_add_12_51_groupi_n_2958 ,csa_tree_add_12_51_groupi_n_2959);
  not csa_tree_add_12_51_groupi_g18828(csa_tree_add_12_51_groupi_n_2950 ,csa_tree_add_12_51_groupi_n_2951);
  or csa_tree_add_12_51_groupi_g18830(csa_tree_add_12_51_groupi_n_2906 ,in2[11] ,csa_tree_add_12_51_groupi_n_2725);
  nor csa_tree_add_12_51_groupi_g18831(csa_tree_add_12_51_groupi_n_2905 ,csa_tree_add_12_51_groupi_n_1335 ,csa_tree_add_12_51_groupi_n_255);
  or csa_tree_add_12_51_groupi_g18832(csa_tree_add_12_51_groupi_n_2904 ,in3[2] ,csa_tree_add_12_51_groupi_n_2744);
  or csa_tree_add_12_51_groupi_g18833(csa_tree_add_12_51_groupi_n_2903 ,csa_tree_add_12_51_groupi_n_1932 ,csa_tree_add_12_51_groupi_n_2737);
  nor csa_tree_add_12_51_groupi_g18834(csa_tree_add_12_51_groupi_n_2902 ,csa_tree_add_12_51_groupi_n_229 ,csa_tree_add_12_51_groupi_n_987);
  nor csa_tree_add_12_51_groupi_g18835(csa_tree_add_12_51_groupi_n_2901 ,in3[2] ,csa_tree_add_12_51_groupi_n_2649);
  or csa_tree_add_12_51_groupi_g18836(csa_tree_add_12_51_groupi_n_2900 ,csa_tree_add_12_51_groupi_n_117 ,csa_tree_add_12_51_groupi_n_2728);
  or csa_tree_add_12_51_groupi_g18837(csa_tree_add_12_51_groupi_n_2899 ,csa_tree_add_12_51_groupi_n_2402 ,csa_tree_add_12_51_groupi_n_2749);
  or csa_tree_add_12_51_groupi_g18838(csa_tree_add_12_51_groupi_n_2898 ,in4[11] ,csa_tree_add_12_51_groupi_n_2746);
  nor csa_tree_add_12_51_groupi_g18839(csa_tree_add_12_51_groupi_n_2897 ,csa_tree_add_12_51_groupi_n_1047 ,csa_tree_add_12_51_groupi_n_1251);
  or csa_tree_add_12_51_groupi_g18840(csa_tree_add_12_51_groupi_n_2896 ,csa_tree_add_12_51_groupi_n_122 ,csa_tree_add_12_51_groupi_n_2698);
  or csa_tree_add_12_51_groupi_g18841(csa_tree_add_12_51_groupi_n_2895 ,in4[2] ,csa_tree_add_12_51_groupi_n_2738);
  or csa_tree_add_12_51_groupi_g18842(csa_tree_add_12_51_groupi_n_2894 ,in2[5] ,csa_tree_add_12_51_groupi_n_2741);
  or csa_tree_add_12_51_groupi_g18843(csa_tree_add_12_51_groupi_n_2893 ,in2[8] ,csa_tree_add_12_51_groupi_n_2742);
  or csa_tree_add_12_51_groupi_g18844(csa_tree_add_12_51_groupi_n_2892 ,in4[5] ,csa_tree_add_12_51_groupi_n_2731);
  or csa_tree_add_12_51_groupi_g18845(csa_tree_add_12_51_groupi_n_2891 ,in3[11] ,csa_tree_add_12_51_groupi_n_2729);
  or csa_tree_add_12_51_groupi_g18846(csa_tree_add_12_51_groupi_n_2890 ,csa_tree_add_12_51_groupi_n_125 ,csa_tree_add_12_51_groupi_n_2730);
  nor csa_tree_add_12_51_groupi_g18847(csa_tree_add_12_51_groupi_n_2889 ,csa_tree_add_12_51_groupi_n_1049 ,csa_tree_add_12_51_groupi_n_1083);
  or csa_tree_add_12_51_groupi_g18848(csa_tree_add_12_51_groupi_n_2888 ,in3[5] ,csa_tree_add_12_51_groupi_n_2736);
  or csa_tree_add_12_51_groupi_g18849(csa_tree_add_12_51_groupi_n_2887 ,csa_tree_add_12_51_groupi_n_1892 ,csa_tree_add_12_51_groupi_n_2750);
  or csa_tree_add_12_51_groupi_g18850(csa_tree_add_12_51_groupi_n_2886 ,in2[2] ,csa_tree_add_12_51_groupi_n_2748);
  nor csa_tree_add_12_51_groupi_g18851(csa_tree_add_12_51_groupi_n_2885 ,csa_tree_add_12_51_groupi_n_1467 ,csa_tree_add_12_51_groupi_n_1074);
  or csa_tree_add_12_51_groupi_g18852(csa_tree_add_12_51_groupi_n_2884 ,in4[8] ,csa_tree_add_12_51_groupi_n_2727);
  nor csa_tree_add_12_51_groupi_g18853(csa_tree_add_12_51_groupi_n_2883 ,csa_tree_add_12_51_groupi_n_1334 ,csa_tree_add_12_51_groupi_n_193);
  nor csa_tree_add_12_51_groupi_g18854(csa_tree_add_12_51_groupi_n_2882 ,csa_tree_add_12_51_groupi_n_1470 ,csa_tree_add_12_51_groupi_n_941);
  or csa_tree_add_12_51_groupi_g18855(csa_tree_add_12_51_groupi_n_2881 ,csa_tree_add_12_51_groupi_n_1951 ,csa_tree_add_12_51_groupi_n_2740);
  or csa_tree_add_12_51_groupi_g18856(csa_tree_add_12_51_groupi_n_2880 ,csa_tree_add_12_51_groupi_n_1947 ,csa_tree_add_12_51_groupi_n_2726);
  or csa_tree_add_12_51_groupi_g18857(csa_tree_add_12_51_groupi_n_2879 ,in3[8] ,csa_tree_add_12_51_groupi_n_2733);
  nor csa_tree_add_12_51_groupi_g18858(csa_tree_add_12_51_groupi_n_2878 ,csa_tree_add_12_51_groupi_n_1491 ,csa_tree_add_12_51_groupi_n_373);
  nor csa_tree_add_12_51_groupi_g18859(csa_tree_add_12_51_groupi_n_2877 ,csa_tree_add_12_51_groupi_n_1266 ,csa_tree_add_12_51_groupi_n_1251);
  or csa_tree_add_12_51_groupi_g18860(csa_tree_add_12_51_groupi_n_2876 ,csa_tree_add_12_51_groupi_n_2365 ,csa_tree_add_12_51_groupi_n_2739);
  nor csa_tree_add_12_51_groupi_g18861(csa_tree_add_12_51_groupi_n_2875 ,csa_tree_add_12_51_groupi_n_1262 ,csa_tree_add_12_51_groupi_n_984);
  or csa_tree_add_12_51_groupi_g18862(csa_tree_add_12_51_groupi_n_2874 ,csa_tree_add_12_51_groupi_n_98 ,csa_tree_add_12_51_groupi_n_2747);
  or csa_tree_add_12_51_groupi_g18863(csa_tree_add_12_51_groupi_n_2873 ,csa_tree_add_12_51_groupi_n_1949 ,csa_tree_add_12_51_groupi_n_2745);
  or csa_tree_add_12_51_groupi_g18864(csa_tree_add_12_51_groupi_n_2872 ,csa_tree_add_12_51_groupi_n_1894 ,csa_tree_add_12_51_groupi_n_2732);
  and csa_tree_add_12_51_groupi_g18865(csa_tree_add_12_51_groupi_n_2961 ,csa_tree_add_12_51_groupi_n_2451 ,csa_tree_add_12_51_groupi_n_2682);
  and csa_tree_add_12_51_groupi_g18866(csa_tree_add_12_51_groupi_n_2960 ,csa_tree_add_12_51_groupi_n_2439 ,csa_tree_add_12_51_groupi_n_2685);
  and csa_tree_add_12_51_groupi_g18867(csa_tree_add_12_51_groupi_n_2959 ,csa_tree_add_12_51_groupi_n_2443 ,csa_tree_add_12_51_groupi_n_2679);
  or csa_tree_add_12_51_groupi_g18868(csa_tree_add_12_51_groupi_n_2957 ,csa_tree_add_12_51_groupi_n_2446 ,csa_tree_add_12_51_groupi_n_2720);
  or csa_tree_add_12_51_groupi_g18869(csa_tree_add_12_51_groupi_n_2956 ,csa_tree_add_12_51_groupi_n_2474 ,csa_tree_add_12_51_groupi_n_2722);
  or csa_tree_add_12_51_groupi_g18870(csa_tree_add_12_51_groupi_n_2955 ,csa_tree_add_12_51_groupi_n_2473 ,csa_tree_add_12_51_groupi_n_2681);
  or csa_tree_add_12_51_groupi_g18871(csa_tree_add_12_51_groupi_n_2954 ,csa_tree_add_12_51_groupi_n_2471 ,csa_tree_add_12_51_groupi_n_2723);
  or csa_tree_add_12_51_groupi_g18872(csa_tree_add_12_51_groupi_n_2953 ,csa_tree_add_12_51_groupi_n_2453 ,csa_tree_add_12_51_groupi_n_2724);
  or csa_tree_add_12_51_groupi_g18873(csa_tree_add_12_51_groupi_n_2952 ,csa_tree_add_12_51_groupi_n_2449 ,csa_tree_add_12_51_groupi_n_2721);
  and csa_tree_add_12_51_groupi_g18874(csa_tree_add_12_51_groupi_n_2951 ,csa_tree_add_12_51_groupi_n_2472 ,csa_tree_add_12_51_groupi_n_2680);
  or csa_tree_add_12_51_groupi_g18875(csa_tree_add_12_51_groupi_n_2949 ,csa_tree_add_12_51_groupi_n_1960 ,csa_tree_add_12_51_groupi_n_2648);
  and csa_tree_add_12_51_groupi_g18876(csa_tree_add_12_51_groupi_n_2948 ,csa_tree_add_12_51_groupi_n_2693 ,csa_tree_add_12_51_groupi_n_2703);
  or csa_tree_add_12_51_groupi_g18877(csa_tree_add_12_51_groupi_n_2947 ,csa_tree_add_12_51_groupi_n_2380 ,csa_tree_add_12_51_groupi_n_2658);
  and csa_tree_add_12_51_groupi_g18878(csa_tree_add_12_51_groupi_n_2946 ,csa_tree_add_12_51_groupi_n_2708 ,csa_tree_add_12_51_groupi_n_2718);
  and csa_tree_add_12_51_groupi_g18879(csa_tree_add_12_51_groupi_n_2945 ,csa_tree_add_12_51_groupi_n_2716 ,csa_tree_add_12_51_groupi_n_2686);
  and csa_tree_add_12_51_groupi_g18880(csa_tree_add_12_51_groupi_n_2944 ,csa_tree_add_12_51_groupi_n_2704 ,csa_tree_add_12_51_groupi_n_2751);
  and csa_tree_add_12_51_groupi_g18881(csa_tree_add_12_51_groupi_n_2943 ,csa_tree_add_12_51_groupi_n_2707 ,csa_tree_add_12_51_groupi_n_2714);
  or csa_tree_add_12_51_groupi_g18882(csa_tree_add_12_51_groupi_n_2942 ,csa_tree_add_12_51_groupi_n_2383 ,csa_tree_add_12_51_groupi_n_2662);
  or csa_tree_add_12_51_groupi_g18883(csa_tree_add_12_51_groupi_n_2941 ,csa_tree_add_12_51_groupi_n_2382 ,csa_tree_add_12_51_groupi_n_2660);
  or csa_tree_add_12_51_groupi_g18884(csa_tree_add_12_51_groupi_n_2940 ,csa_tree_add_12_51_groupi_n_2645 ,csa_tree_add_12_51_groupi_n_2767);
  or csa_tree_add_12_51_groupi_g18885(csa_tree_add_12_51_groupi_n_2939 ,csa_tree_add_12_51_groupi_n_2646 ,csa_tree_add_12_51_groupi_n_2775);
  and csa_tree_add_12_51_groupi_g18886(csa_tree_add_12_51_groupi_n_2938 ,csa_tree_add_12_51_groupi_n_2711 ,csa_tree_add_12_51_groupi_n_2683);
  or csa_tree_add_12_51_groupi_g18887(csa_tree_add_12_51_groupi_n_2937 ,csa_tree_add_12_51_groupi_n_2656 ,csa_tree_add_12_51_groupi_n_2779);
  and csa_tree_add_12_51_groupi_g18888(csa_tree_add_12_51_groupi_n_2936 ,csa_tree_add_12_51_groupi_n_2696 ,csa_tree_add_12_51_groupi_n_2719);
  or csa_tree_add_12_51_groupi_g18889(csa_tree_add_12_51_groupi_n_2935 ,csa_tree_add_12_51_groupi_n_2647 ,csa_tree_add_12_51_groupi_n_2761);
  and csa_tree_add_12_51_groupi_g18890(csa_tree_add_12_51_groupi_n_2934 ,csa_tree_add_12_51_groupi_n_2701 ,csa_tree_add_12_51_groupi_n_2700);
  and csa_tree_add_12_51_groupi_g18891(csa_tree_add_12_51_groupi_n_2933 ,csa_tree_add_12_51_groupi_n_2689 ,csa_tree_add_12_51_groupi_n_2684);
  or csa_tree_add_12_51_groupi_g18892(csa_tree_add_12_51_groupi_n_2932 ,csa_tree_add_12_51_groupi_n_2644 ,csa_tree_add_12_51_groupi_n_2771);
  and csa_tree_add_12_51_groupi_g18893(csa_tree_add_12_51_groupi_n_2931 ,csa_tree_add_12_51_groupi_n_2697 ,csa_tree_add_12_51_groupi_n_2692);
  or csa_tree_add_12_51_groupi_g18894(csa_tree_add_12_51_groupi_n_2930 ,csa_tree_add_12_51_groupi_n_2654 ,csa_tree_add_12_51_groupi_n_2765);
  and csa_tree_add_12_51_groupi_g18895(csa_tree_add_12_51_groupi_n_2929 ,csa_tree_add_12_51_groupi_n_2699 ,csa_tree_add_12_51_groupi_n_2705);
  or csa_tree_add_12_51_groupi_g18896(csa_tree_add_12_51_groupi_n_2928 ,csa_tree_add_12_51_groupi_n_2652 ,csa_tree_add_12_51_groupi_n_2769);
  and csa_tree_add_12_51_groupi_g18897(csa_tree_add_12_51_groupi_n_2927 ,csa_tree_add_12_51_groupi_n_2712 ,csa_tree_add_12_51_groupi_n_2695);
  or csa_tree_add_12_51_groupi_g18898(csa_tree_add_12_51_groupi_n_2926 ,csa_tree_add_12_51_groupi_n_2657 ,csa_tree_add_12_51_groupi_n_2777);
  or csa_tree_add_12_51_groupi_g18899(csa_tree_add_12_51_groupi_n_2925 ,csa_tree_add_12_51_groupi_n_2653 ,csa_tree_add_12_51_groupi_n_2759);
  or csa_tree_add_12_51_groupi_g18900(csa_tree_add_12_51_groupi_n_2924 ,csa_tree_add_12_51_groupi_n_2650 ,csa_tree_add_12_51_groupi_n_2781);
  or csa_tree_add_12_51_groupi_g18901(csa_tree_add_12_51_groupi_n_2923 ,csa_tree_add_12_51_groupi_n_2655 ,csa_tree_add_12_51_groupi_n_2763);
  or csa_tree_add_12_51_groupi_g18902(csa_tree_add_12_51_groupi_n_2922 ,csa_tree_add_12_51_groupi_n_2651 ,csa_tree_add_12_51_groupi_n_2773);
  or csa_tree_add_12_51_groupi_g18903(csa_tree_add_12_51_groupi_n_2921 ,csa_tree_add_12_51_groupi_n_2772 ,csa_tree_add_12_51_groupi_n_2644);
  or csa_tree_add_12_51_groupi_g18904(csa_tree_add_12_51_groupi_n_2920 ,csa_tree_add_12_51_groupi_n_2782 ,csa_tree_add_12_51_groupi_n_2650);
  or csa_tree_add_12_51_groupi_g18905(csa_tree_add_12_51_groupi_n_2919 ,csa_tree_add_12_51_groupi_n_2764 ,csa_tree_add_12_51_groupi_n_2655);
  or csa_tree_add_12_51_groupi_g18906(csa_tree_add_12_51_groupi_n_2918 ,csa_tree_add_12_51_groupi_n_2760 ,csa_tree_add_12_51_groupi_n_2653);
  or csa_tree_add_12_51_groupi_g18907(csa_tree_add_12_51_groupi_n_2917 ,csa_tree_add_12_51_groupi_n_2774 ,csa_tree_add_12_51_groupi_n_2651);
  or csa_tree_add_12_51_groupi_g18908(csa_tree_add_12_51_groupi_n_2916 ,csa_tree_add_12_51_groupi_n_2766 ,csa_tree_add_12_51_groupi_n_2654);
  or csa_tree_add_12_51_groupi_g18909(csa_tree_add_12_51_groupi_n_2915 ,csa_tree_add_12_51_groupi_n_2770 ,csa_tree_add_12_51_groupi_n_2652);
  or csa_tree_add_12_51_groupi_g18910(csa_tree_add_12_51_groupi_n_2914 ,csa_tree_add_12_51_groupi_n_2778 ,csa_tree_add_12_51_groupi_n_2657);
  or csa_tree_add_12_51_groupi_g18911(csa_tree_add_12_51_groupi_n_2913 ,csa_tree_add_12_51_groupi_n_2768 ,csa_tree_add_12_51_groupi_n_2645);
  or csa_tree_add_12_51_groupi_g18912(csa_tree_add_12_51_groupi_n_2912 ,csa_tree_add_12_51_groupi_n_2780 ,csa_tree_add_12_51_groupi_n_2656);
  or csa_tree_add_12_51_groupi_g18913(csa_tree_add_12_51_groupi_n_2911 ,csa_tree_add_12_51_groupi_n_2776 ,csa_tree_add_12_51_groupi_n_2646);
  or csa_tree_add_12_51_groupi_g18914(csa_tree_add_12_51_groupi_n_2910 ,csa_tree_add_12_51_groupi_n_2762 ,csa_tree_add_12_51_groupi_n_2647);
  or csa_tree_add_12_51_groupi_g18915(csa_tree_add_12_51_groupi_n_2909 ,csa_tree_add_12_51_groupi_n_2380 ,csa_tree_add_12_51_groupi_n_2659);
  or csa_tree_add_12_51_groupi_g18916(csa_tree_add_12_51_groupi_n_2908 ,csa_tree_add_12_51_groupi_n_2382 ,csa_tree_add_12_51_groupi_n_2661);
  or csa_tree_add_12_51_groupi_g18917(csa_tree_add_12_51_groupi_n_2907 ,csa_tree_add_12_51_groupi_n_2383 ,csa_tree_add_12_51_groupi_n_2663);
  not csa_tree_add_12_51_groupi_g18918(csa_tree_add_12_51_groupi_n_2871 ,csa_tree_add_12_51_groupi_n_2870);
  nor csa_tree_add_12_51_groupi_g18919(csa_tree_add_12_51_groupi_n_2867 ,csa_tree_add_12_51_groupi_n_532 ,csa_tree_add_12_51_groupi_n_2193);
  nor csa_tree_add_12_51_groupi_g18920(csa_tree_add_12_51_groupi_n_2866 ,csa_tree_add_12_51_groupi_n_1343 ,csa_tree_add_12_51_groupi_n_241);
  nor csa_tree_add_12_51_groupi_g18921(csa_tree_add_12_51_groupi_n_2865 ,csa_tree_add_12_51_groupi_n_1490 ,csa_tree_add_12_51_groupi_n_361);
  nor csa_tree_add_12_51_groupi_g18922(csa_tree_add_12_51_groupi_n_2864 ,csa_tree_add_12_51_groupi_n_499 ,csa_tree_add_12_51_groupi_n_884);
  nor csa_tree_add_12_51_groupi_g18923(csa_tree_add_12_51_groupi_n_2863 ,csa_tree_add_12_51_groupi_n_1074 ,csa_tree_add_12_51_groupi_n_397);
  nor csa_tree_add_12_51_groupi_g18924(csa_tree_add_12_51_groupi_n_2862 ,csa_tree_add_12_51_groupi_n_1518 ,csa_tree_add_12_51_groupi_n_277);
  nor csa_tree_add_12_51_groupi_g18925(csa_tree_add_12_51_groupi_n_2861 ,csa_tree_add_12_51_groupi_n_1389 ,csa_tree_add_12_51_groupi_n_325);
  nor csa_tree_add_12_51_groupi_g18926(csa_tree_add_12_51_groupi_n_2860 ,csa_tree_add_12_51_groupi_n_1344 ,csa_tree_add_12_51_groupi_n_319);
  nor csa_tree_add_12_51_groupi_g18927(csa_tree_add_12_51_groupi_n_2859 ,csa_tree_add_12_51_groupi_n_1250 ,csa_tree_add_12_51_groupi_n_280);
  nor csa_tree_add_12_51_groupi_g18928(csa_tree_add_12_51_groupi_n_2858 ,csa_tree_add_12_51_groupi_n_1443 ,csa_tree_add_12_51_groupi_n_1517);
  nor csa_tree_add_12_51_groupi_g18929(csa_tree_add_12_51_groupi_n_2857 ,csa_tree_add_12_51_groupi_n_508 ,csa_tree_add_12_51_groupi_n_1335);
  nor csa_tree_add_12_51_groupi_g18930(csa_tree_add_12_51_groupi_n_2856 ,csa_tree_add_12_51_groupi_n_682 ,csa_tree_add_12_51_groupi_n_1334);
  nor csa_tree_add_12_51_groupi_g18931(csa_tree_add_12_51_groupi_n_2855 ,csa_tree_add_12_51_groupi_n_1517 ,csa_tree_add_12_51_groupi_n_211);
  nor csa_tree_add_12_51_groupi_g18932(csa_tree_add_12_51_groupi_n_2854 ,csa_tree_add_12_51_groupi_n_535 ,csa_tree_add_12_51_groupi_n_983);
  nor csa_tree_add_12_51_groupi_g18933(csa_tree_add_12_51_groupi_n_2853 ,csa_tree_add_12_51_groupi_n_1082 ,csa_tree_add_12_51_groupi_n_385);
  nor csa_tree_add_12_51_groupi_g18934(csa_tree_add_12_51_groupi_n_2852 ,csa_tree_add_12_51_groupi_n_1518 ,csa_tree_add_12_51_groupi_n_253);
  nor csa_tree_add_12_51_groupi_g18935(csa_tree_add_12_51_groupi_n_2851 ,csa_tree_add_12_51_groupi_n_675 ,csa_tree_add_12_51_groupi_n_987);
  nor csa_tree_add_12_51_groupi_g18936(csa_tree_add_12_51_groupi_n_2850 ,csa_tree_add_12_51_groupi_n_685 ,csa_tree_add_12_51_groupi_n_1082);
  nor csa_tree_add_12_51_groupi_g18937(csa_tree_add_12_51_groupi_n_2849 ,csa_tree_add_12_51_groupi_n_1388 ,csa_tree_add_12_51_groupi_n_343);
  nor csa_tree_add_12_51_groupi_g18938(csa_tree_add_12_51_groupi_n_2848 ,csa_tree_add_12_51_groupi_n_496 ,csa_tree_add_12_51_groupi_n_1389);
  nor csa_tree_add_12_51_groupi_g18939(csa_tree_add_12_51_groupi_n_2847 ,csa_tree_add_12_51_groupi_n_492 ,csa_tree_add_12_51_groupi_n_984);
  nor csa_tree_add_12_51_groupi_g18940(csa_tree_add_12_51_groupi_n_2846 ,csa_tree_add_12_51_groupi_n_490 ,csa_tree_add_12_51_groupi_n_986);
  nor csa_tree_add_12_51_groupi_g18941(csa_tree_add_12_51_groupi_n_2845 ,csa_tree_add_12_51_groupi_n_1404 ,csa_tree_add_12_51_groupi_n_1388);
  nor csa_tree_add_12_51_groupi_g18942(csa_tree_add_12_51_groupi_n_2844 ,csa_tree_add_12_51_groupi_n_1449 ,csa_tree_add_12_51_groupi_n_884);
  nor csa_tree_add_12_51_groupi_g18943(csa_tree_add_12_51_groupi_n_2843 ,csa_tree_add_12_51_groupi_n_546 ,csa_tree_add_12_51_groupi_n_986);
  nor csa_tree_add_12_51_groupi_g18944(csa_tree_add_12_51_groupi_n_2842 ,csa_tree_add_12_51_groupi_n_691 ,csa_tree_add_12_51_groupi_n_942);
  nor csa_tree_add_12_51_groupi_g18945(csa_tree_add_12_51_groupi_n_2841 ,csa_tree_add_12_51_groupi_n_688 ,csa_tree_add_12_51_groupi_n_1250);
  nor csa_tree_add_12_51_groupi_g18946(csa_tree_add_12_51_groupi_n_2840 ,csa_tree_add_12_51_groupi_n_511 ,csa_tree_add_12_51_groupi_n_1073);
  nor csa_tree_add_12_51_groupi_g18947(csa_tree_add_12_51_groupi_n_2839 ,csa_tree_add_12_51_groupi_n_1455 ,csa_tree_add_12_51_groupi_n_983);
  nor csa_tree_add_12_51_groupi_g18948(csa_tree_add_12_51_groupi_n_2838 ,csa_tree_add_12_51_groupi_n_517 ,csa_tree_add_12_51_groupi_n_885);
  nor csa_tree_add_12_51_groupi_g18949(csa_tree_add_12_51_groupi_n_2837 ,csa_tree_add_12_51_groupi_n_628 ,csa_tree_add_12_51_groupi_n_1083);
  nor csa_tree_add_12_51_groupi_g18950(csa_tree_add_12_51_groupi_n_2836 ,csa_tree_add_12_51_groupi_n_1491 ,csa_tree_add_12_51_groupi_n_205);
  nor csa_tree_add_12_51_groupi_g18951(csa_tree_add_12_51_groupi_n_2835 ,csa_tree_add_12_51_groupi_n_519 ,csa_tree_add_12_51_groupi_n_1490);
  nor csa_tree_add_12_51_groupi_g18952(csa_tree_add_12_51_groupi_n_2834 ,csa_tree_add_12_51_groupi_n_583 ,csa_tree_add_12_51_groupi_n_942);
  nor csa_tree_add_12_51_groupi_g18953(csa_tree_add_12_51_groupi_n_2833 ,csa_tree_add_12_51_groupi_n_553 ,csa_tree_add_12_51_groupi_n_885);
  nor csa_tree_add_12_51_groupi_g18954(csa_tree_add_12_51_groupi_n_2832 ,csa_tree_add_12_51_groupi_n_1464 ,csa_tree_add_12_51_groupi_n_1344);
  nor csa_tree_add_12_51_groupi_g18955(csa_tree_add_12_51_groupi_n_2831 ,csa_tree_add_12_51_groupi_n_1446 ,csa_tree_add_12_51_groupi_n_1343);
  nor csa_tree_add_12_51_groupi_g18956(csa_tree_add_12_51_groupi_n_2830 ,csa_tree_add_12_51_groupi_n_667 ,csa_tree_add_12_51_groupi_n_941);
  and csa_tree_add_12_51_groupi_g18957(csa_tree_add_12_51_groupi_n_2829 ,csa_tree_add_12_51_groupi_n_2758 ,csa_tree_add_12_51_groupi_n_2755);
  or csa_tree_add_12_51_groupi_g18958(csa_tree_add_12_51_groupi_n_2828 ,csa_tree_add_12_51_groupi_n_2758 ,csa_tree_add_12_51_groupi_n_2755);
  nor csa_tree_add_12_51_groupi_g18959(csa_tree_add_12_51_groupi_n_2827 ,csa_tree_add_12_51_groupi_n_622 ,csa_tree_add_12_51_groupi_n_867);
  nor csa_tree_add_12_51_groupi_g18960(csa_tree_add_12_51_groupi_n_2826 ,csa_tree_add_12_51_groupi_n_693 ,csa_tree_add_12_51_groupi_n_981);
  nor csa_tree_add_12_51_groupi_g18961(csa_tree_add_12_51_groupi_n_2825 ,csa_tree_add_12_51_groupi_n_463 ,csa_tree_add_12_51_groupi_n_2189);
  nor csa_tree_add_12_51_groupi_g18962(csa_tree_add_12_51_groupi_n_2824 ,csa_tree_add_12_51_groupi_n_658 ,csa_tree_add_12_51_groupi_n_966);
  nor csa_tree_add_12_51_groupi_g18963(csa_tree_add_12_51_groupi_n_2823 ,csa_tree_add_12_51_groupi_n_529 ,csa_tree_add_12_51_groupi_n_1073);
  nor csa_tree_add_12_51_groupi_g18964(csa_tree_add_12_51_groupi_n_2822 ,csa_tree_add_12_51_groupi_n_663 ,csa_tree_add_12_51_groupi_n_969);
  nor csa_tree_add_12_51_groupi_g18965(csa_tree_add_12_51_groupi_n_2821 ,csa_tree_add_12_51_groupi_n_1071 ,csa_tree_add_12_51_groupi_n_322);
  nor csa_tree_add_12_51_groupi_g18966(csa_tree_add_12_51_groupi_n_2820 ,csa_tree_add_12_51_groupi_n_550 ,csa_tree_add_12_51_groupi_n_980);
  nor csa_tree_add_12_51_groupi_g18967(csa_tree_add_12_51_groupi_n_2819 ,csa_tree_add_12_51_groupi_n_538 ,csa_tree_add_12_51_groupi_n_709);
  nor csa_tree_add_12_51_groupi_g18968(csa_tree_add_12_51_groupi_n_2818 ,csa_tree_add_12_51_groupi_n_559 ,csa_tree_add_12_51_groupi_n_708);
  nor csa_tree_add_12_51_groupi_g18969(csa_tree_add_12_51_groupi_n_2817 ,csa_tree_add_12_51_groupi_n_616 ,csa_tree_add_12_51_groupi_n_981);
  nor csa_tree_add_12_51_groupi_g18970(csa_tree_add_12_51_groupi_n_2816 ,csa_tree_add_12_51_groupi_n_1709 ,csa_tree_add_12_51_groupi_n_712);
  nor csa_tree_add_12_51_groupi_g18971(csa_tree_add_12_51_groupi_n_2815 ,csa_tree_add_12_51_groupi_n_679 ,csa_tree_add_12_51_groupi_n_711);
  nor csa_tree_add_12_51_groupi_g18972(csa_tree_add_12_51_groupi_n_2814 ,csa_tree_add_12_51_groupi_n_541 ,csa_tree_add_12_51_groupi_n_1070);
  nor csa_tree_add_12_51_groupi_g18973(csa_tree_add_12_51_groupi_n_2813 ,csa_tree_add_12_51_groupi_n_574 ,csa_tree_add_12_51_groupi_n_980);
  nor csa_tree_add_12_51_groupi_g18974(csa_tree_add_12_51_groupi_n_2812 ,csa_tree_add_12_51_groupi_n_1568 ,csa_tree_add_12_51_groupi_n_1071);
  nor csa_tree_add_12_51_groupi_g18975(csa_tree_add_12_51_groupi_n_2811 ,csa_tree_add_12_51_groupi_n_619 ,csa_tree_add_12_51_groupi_n_2186);
  nor csa_tree_add_12_51_groupi_g18976(csa_tree_add_12_51_groupi_n_2810 ,csa_tree_add_12_51_groupi_n_637 ,csa_tree_add_12_51_groupi_n_977);
  nor csa_tree_add_12_51_groupi_g18977(csa_tree_add_12_51_groupi_n_2809 ,csa_tree_add_12_51_groupi_n_649 ,csa_tree_add_12_51_groupi_n_978);
  nor csa_tree_add_12_51_groupi_g18978(csa_tree_add_12_51_groupi_n_2808 ,csa_tree_add_12_51_groupi_n_568 ,csa_tree_add_12_51_groupi_n_867);
  nor csa_tree_add_12_51_groupi_g18979(csa_tree_add_12_51_groupi_n_2807 ,csa_tree_add_12_51_groupi_n_625 ,csa_tree_add_12_51_groupi_n_2190);
  nor csa_tree_add_12_51_groupi_g18980(csa_tree_add_12_51_groupi_n_2806 ,csa_tree_add_12_51_groupi_n_673 ,csa_tree_add_12_51_groupi_n_2186);
  nor csa_tree_add_12_51_groupi_g18981(csa_tree_add_12_51_groupi_n_2805 ,csa_tree_add_12_51_groupi_n_1766 ,csa_tree_add_12_51_groupi_n_978);
  nor csa_tree_add_12_51_groupi_g18982(csa_tree_add_12_51_groupi_n_2804 ,csa_tree_add_12_51_groupi_n_634 ,csa_tree_add_12_51_groupi_n_2187);
  nor csa_tree_add_12_51_groupi_g18983(csa_tree_add_12_51_groupi_n_2803 ,csa_tree_add_12_51_groupi_n_577 ,csa_tree_add_12_51_groupi_n_1070);
  nor csa_tree_add_12_51_groupi_g18984(csa_tree_add_12_51_groupi_n_2802 ,csa_tree_add_12_51_groupi_n_1784 ,csa_tree_add_12_51_groupi_n_866);
  nor csa_tree_add_12_51_groupi_g18985(csa_tree_add_12_51_groupi_n_2801 ,csa_tree_add_12_51_groupi_n_1796 ,csa_tree_add_12_51_groupi_n_2187);
  nor csa_tree_add_12_51_groupi_g18986(csa_tree_add_12_51_groupi_n_2800 ,csa_tree_add_12_51_groupi_n_1718 ,csa_tree_add_12_51_groupi_n_712);
  nor csa_tree_add_12_51_groupi_g18987(csa_tree_add_12_51_groupi_n_2799 ,csa_tree_add_12_51_groupi_n_1787 ,csa_tree_add_12_51_groupi_n_2192);
  nor csa_tree_add_12_51_groupi_g18988(csa_tree_add_12_51_groupi_n_2798 ,csa_tree_add_12_51_groupi_n_586 ,csa_tree_add_12_51_groupi_n_866);
  nor csa_tree_add_12_51_groupi_g18989(csa_tree_add_12_51_groupi_n_2797 ,csa_tree_add_12_51_groupi_n_580 ,csa_tree_add_12_51_groupi_n_709);
  nor csa_tree_add_12_51_groupi_g18990(csa_tree_add_12_51_groupi_n_2796 ,csa_tree_add_12_51_groupi_n_607 ,csa_tree_add_12_51_groupi_n_2157);
  nor csa_tree_add_12_51_groupi_g18991(csa_tree_add_12_51_groupi_n_2795 ,csa_tree_add_12_51_groupi_n_1721 ,csa_tree_add_12_51_groupi_n_968);
  nor csa_tree_add_12_51_groupi_g18992(csa_tree_add_12_51_groupi_n_2794 ,csa_tree_add_12_51_groupi_n_1775 ,csa_tree_add_12_51_groupi_n_968);
  nor csa_tree_add_12_51_groupi_g18993(csa_tree_add_12_51_groupi_n_2793 ,csa_tree_add_12_51_groupi_n_1751 ,csa_tree_add_12_51_groupi_n_2642);
  nor csa_tree_add_12_51_groupi_g18994(csa_tree_add_12_51_groupi_n_2792 ,csa_tree_add_12_51_groupi_n_1757 ,csa_tree_add_12_51_groupi_n_977);
  nor csa_tree_add_12_51_groupi_g18995(csa_tree_add_12_51_groupi_n_2791 ,csa_tree_add_12_51_groupi_n_604 ,csa_tree_add_12_51_groupi_n_2189);
  nor csa_tree_add_12_51_groupi_g18996(csa_tree_add_12_51_groupi_n_2790 ,csa_tree_add_12_51_groupi_n_1730 ,csa_tree_add_12_51_groupi_n_965);
  nor csa_tree_add_12_51_groupi_g18997(csa_tree_add_12_51_groupi_n_2789 ,csa_tree_add_12_51_groupi_n_1754 ,csa_tree_add_12_51_groupi_n_965);
  nor csa_tree_add_12_51_groupi_g18998(csa_tree_add_12_51_groupi_n_2788 ,csa_tree_add_12_51_groupi_n_1799 ,csa_tree_add_12_51_groupi_n_969);
  nor csa_tree_add_12_51_groupi_g18999(csa_tree_add_12_51_groupi_n_2787 ,csa_tree_add_12_51_groupi_n_612 ,csa_tree_add_12_51_groupi_n_2190);
  nor csa_tree_add_12_51_groupi_g19000(csa_tree_add_12_51_groupi_n_2786 ,csa_tree_add_12_51_groupi_n_646 ,csa_tree_add_12_51_groupi_n_966);
  nor csa_tree_add_12_51_groupi_g19001(csa_tree_add_12_51_groupi_n_2785 ,csa_tree_add_12_51_groupi_n_1700 ,csa_tree_add_12_51_groupi_n_2157);
  nor csa_tree_add_12_51_groupi_g19002(csa_tree_add_12_51_groupi_n_2784 ,csa_tree_add_12_51_groupi_n_670 ,csa_tree_add_12_51_groupi_n_2193);
  nor csa_tree_add_12_51_groupi_g19003(csa_tree_add_12_51_groupi_n_2783 ,csa_tree_add_12_51_groupi_n_598 ,csa_tree_add_12_51_groupi_n_2192);
  and csa_tree_add_12_51_groupi_g19004(csa_tree_add_12_51_groupi_n_2870 ,in1[0] ,csa_tree_add_12_51_groupi_n_1908);
  or csa_tree_add_12_51_groupi_g19005(csa_tree_add_12_51_groupi_n_2869 ,csa_tree_add_12_51_groupi_n_1049 ,csa_tree_add_12_51_groupi_n_708);
  or csa_tree_add_12_51_groupi_g19006(csa_tree_add_12_51_groupi_n_2868 ,csa_tree_add_12_51_groupi_n_699 ,csa_tree_add_12_51_groupi_n_711);
  not csa_tree_add_12_51_groupi_g19007(csa_tree_add_12_51_groupi_n_2782 ,csa_tree_add_12_51_groupi_n_2781);
  not csa_tree_add_12_51_groupi_g19008(csa_tree_add_12_51_groupi_n_2780 ,csa_tree_add_12_51_groupi_n_2779);
  not csa_tree_add_12_51_groupi_g19009(csa_tree_add_12_51_groupi_n_2778 ,csa_tree_add_12_51_groupi_n_2777);
  not csa_tree_add_12_51_groupi_g19010(csa_tree_add_12_51_groupi_n_2776 ,csa_tree_add_12_51_groupi_n_2775);
  not csa_tree_add_12_51_groupi_g19011(csa_tree_add_12_51_groupi_n_2774 ,csa_tree_add_12_51_groupi_n_2773);
  not csa_tree_add_12_51_groupi_g19012(csa_tree_add_12_51_groupi_n_2772 ,csa_tree_add_12_51_groupi_n_2771);
  not csa_tree_add_12_51_groupi_g19013(csa_tree_add_12_51_groupi_n_2770 ,csa_tree_add_12_51_groupi_n_2769);
  not csa_tree_add_12_51_groupi_g19014(csa_tree_add_12_51_groupi_n_2768 ,csa_tree_add_12_51_groupi_n_2767);
  not csa_tree_add_12_51_groupi_g19015(csa_tree_add_12_51_groupi_n_2766 ,csa_tree_add_12_51_groupi_n_2765);
  not csa_tree_add_12_51_groupi_g19016(csa_tree_add_12_51_groupi_n_2764 ,csa_tree_add_12_51_groupi_n_2763);
  not csa_tree_add_12_51_groupi_g19017(csa_tree_add_12_51_groupi_n_2762 ,csa_tree_add_12_51_groupi_n_2761);
  not csa_tree_add_12_51_groupi_g19018(csa_tree_add_12_51_groupi_n_2760 ,csa_tree_add_12_51_groupi_n_2759);
  not csa_tree_add_12_51_groupi_g19019(csa_tree_add_12_51_groupi_n_2757 ,csa_tree_add_12_51_groupi_n_2756);
  or csa_tree_add_12_51_groupi_g19020(csa_tree_add_12_51_groupi_n_2751 ,in3[11] ,csa_tree_add_12_51_groupi_n_2502);
  or csa_tree_add_12_51_groupi_g19021(csa_tree_add_12_51_groupi_n_2750 ,csa_tree_add_12_51_groupi_n_2368 ,csa_tree_add_12_51_groupi_n_2547);
  or csa_tree_add_12_51_groupi_g19022(csa_tree_add_12_51_groupi_n_2749 ,csa_tree_add_12_51_groupi_n_2372 ,csa_tree_add_12_51_groupi_n_2509);
  or csa_tree_add_12_51_groupi_g19023(csa_tree_add_12_51_groupi_n_2748 ,in2[3] ,csa_tree_add_12_51_groupi_n_2534);
  or csa_tree_add_12_51_groupi_g19024(csa_tree_add_12_51_groupi_n_2747 ,csa_tree_add_12_51_groupi_n_2377 ,csa_tree_add_12_51_groupi_n_2521);
  or csa_tree_add_12_51_groupi_g19025(csa_tree_add_12_51_groupi_n_2746 ,in4[12] ,csa_tree_add_12_51_groupi_n_2540);
  or csa_tree_add_12_51_groupi_g19026(csa_tree_add_12_51_groupi_n_2745 ,csa_tree_add_12_51_groupi_n_2370 ,csa_tree_add_12_51_groupi_n_2537);
  or csa_tree_add_12_51_groupi_g19027(csa_tree_add_12_51_groupi_n_2744 ,in3[3] ,csa_tree_add_12_51_groupi_n_2512);
  nor csa_tree_add_12_51_groupi_g19028(csa_tree_add_12_51_groupi_n_2743 ,csa_tree_add_12_51_groupi_n_1652 ,csa_tree_add_12_51_groupi_n_247);
  or csa_tree_add_12_51_groupi_g19029(csa_tree_add_12_51_groupi_n_2742 ,in2[9] ,csa_tree_add_12_51_groupi_n_2524);
  or csa_tree_add_12_51_groupi_g19030(csa_tree_add_12_51_groupi_n_2741 ,in2[6] ,csa_tree_add_12_51_groupi_n_2476);
  or csa_tree_add_12_51_groupi_g19031(csa_tree_add_12_51_groupi_n_2740 ,csa_tree_add_12_51_groupi_n_2406 ,csa_tree_add_12_51_groupi_n_2531);
  or csa_tree_add_12_51_groupi_g19032(csa_tree_add_12_51_groupi_n_2739 ,csa_tree_add_12_51_groupi_n_2405 ,csa_tree_add_12_51_groupi_n_2543);
  or csa_tree_add_12_51_groupi_g19033(csa_tree_add_12_51_groupi_n_2738 ,in4[3] ,csa_tree_add_12_51_groupi_n_2528);
  or csa_tree_add_12_51_groupi_g19034(csa_tree_add_12_51_groupi_n_2737 ,csa_tree_add_12_51_groupi_n_2374 ,csa_tree_add_12_51_groupi_n_2469);
  or csa_tree_add_12_51_groupi_g19035(csa_tree_add_12_51_groupi_n_2736 ,in3[6] ,csa_tree_add_12_51_groupi_n_2514);
  nor csa_tree_add_12_51_groupi_g19036(csa_tree_add_12_51_groupi_n_2735 ,csa_tree_add_12_51_groupi_n_466 ,csa_tree_add_12_51_groupi_n_2169);
  nor csa_tree_add_12_51_groupi_g19037(csa_tree_add_12_51_groupi_n_2734 ,csa_tree_add_12_51_groupi_n_1221 ,csa_tree_add_12_51_groupi_n_271);
  or csa_tree_add_12_51_groupi_g19038(csa_tree_add_12_51_groupi_n_2733 ,in3[9] ,csa_tree_add_12_51_groupi_n_2520);
  or csa_tree_add_12_51_groupi_g19039(csa_tree_add_12_51_groupi_n_2732 ,csa_tree_add_12_51_groupi_n_2371 ,csa_tree_add_12_51_groupi_n_2515);
  or csa_tree_add_12_51_groupi_g19040(csa_tree_add_12_51_groupi_n_2731 ,in4[6] ,csa_tree_add_12_51_groupi_n_2508);
  or csa_tree_add_12_51_groupi_g19041(csa_tree_add_12_51_groupi_n_2730 ,csa_tree_add_12_51_groupi_n_2375 ,csa_tree_add_12_51_groupi_n_2525);
  or csa_tree_add_12_51_groupi_g19042(csa_tree_add_12_51_groupi_n_2729 ,in3[12] ,csa_tree_add_12_51_groupi_n_2550);
  or csa_tree_add_12_51_groupi_g19043(csa_tree_add_12_51_groupi_n_2728 ,csa_tree_add_12_51_groupi_n_2376 ,csa_tree_add_12_51_groupi_n_2529);
  or csa_tree_add_12_51_groupi_g19044(csa_tree_add_12_51_groupi_n_2727 ,in4[9] ,csa_tree_add_12_51_groupi_n_2536);
  or csa_tree_add_12_51_groupi_g19045(csa_tree_add_12_51_groupi_n_2726 ,csa_tree_add_12_51_groupi_n_2369 ,csa_tree_add_12_51_groupi_n_2545);
  or csa_tree_add_12_51_groupi_g19046(csa_tree_add_12_51_groupi_n_2725 ,in2[12] ,csa_tree_add_12_51_groupi_n_2542);
  and csa_tree_add_12_51_groupi_g19047(csa_tree_add_12_51_groupi_n_2724 ,in5[12] ,csa_tree_add_12_51_groupi_n_2452);
  nor csa_tree_add_12_51_groupi_g19048(csa_tree_add_12_51_groupi_n_2723 ,csa_tree_add_12_51_groupi_n_2416 ,csa_tree_add_12_51_groupi_n_2473);
  and csa_tree_add_12_51_groupi_g19049(csa_tree_add_12_51_groupi_n_2722 ,in5[3] ,csa_tree_add_12_51_groupi_n_2472);
  and csa_tree_add_12_51_groupi_g19050(csa_tree_add_12_51_groupi_n_2721 ,in5[0] ,csa_tree_add_12_51_groupi_n_2448);
  and csa_tree_add_12_51_groupi_g19051(csa_tree_add_12_51_groupi_n_2720 ,in5[6] ,csa_tree_add_12_51_groupi_n_2445);
  or csa_tree_add_12_51_groupi_g19052(csa_tree_add_12_51_groupi_n_2719 ,in2[8] ,csa_tree_add_12_51_groupi_n_2501);
  or csa_tree_add_12_51_groupi_g19053(csa_tree_add_12_51_groupi_n_2718 ,in3[8] ,csa_tree_add_12_51_groupi_n_2499);
  nor csa_tree_add_12_51_groupi_g19054(csa_tree_add_12_51_groupi_n_2717 ,csa_tree_add_12_51_groupi_n_1286 ,csa_tree_add_12_51_groupi_n_334);
  or csa_tree_add_12_51_groupi_g19055(csa_tree_add_12_51_groupi_n_2716 ,csa_tree_add_12_51_groupi_n_1941 ,csa_tree_add_12_51_groupi_n_2487);
  nor csa_tree_add_12_51_groupi_g19056(csa_tree_add_12_51_groupi_n_2715 ,csa_tree_add_12_51_groupi_n_448 ,csa_tree_add_12_51_groupi_n_2196);
  or csa_tree_add_12_51_groupi_g19057(csa_tree_add_12_51_groupi_n_2714 ,in3[5] ,csa_tree_add_12_51_groupi_n_2489);
  nor csa_tree_add_12_51_groupi_g19058(csa_tree_add_12_51_groupi_n_2713 ,csa_tree_add_12_51_groupi_n_442 ,csa_tree_add_12_51_groupi_n_2198);
  or csa_tree_add_12_51_groupi_g19059(csa_tree_add_12_51_groupi_n_2712 ,csa_tree_add_12_51_groupi_n_1921 ,csa_tree_add_12_51_groupi_n_2492);
  or csa_tree_add_12_51_groupi_g19060(csa_tree_add_12_51_groupi_n_2711 ,csa_tree_add_12_51_groupi_n_1935 ,csa_tree_add_12_51_groupi_n_2503);
  nor csa_tree_add_12_51_groupi_g19061(csa_tree_add_12_51_groupi_n_2710 ,csa_tree_add_12_51_groupi_n_1682 ,csa_tree_add_12_51_groupi_n_298);
  nor csa_tree_add_12_51_groupi_g19062(csa_tree_add_12_51_groupi_n_2709 ,csa_tree_add_12_51_groupi_n_1353 ,csa_tree_add_12_51_groupi_n_214);
  or csa_tree_add_12_51_groupi_g19063(csa_tree_add_12_51_groupi_n_2708 ,csa_tree_add_12_51_groupi_n_1945 ,csa_tree_add_12_51_groupi_n_2494);
  or csa_tree_add_12_51_groupi_g19064(csa_tree_add_12_51_groupi_n_2707 ,csa_tree_add_12_51_groupi_n_1903 ,csa_tree_add_12_51_groupi_n_2491);
  nor csa_tree_add_12_51_groupi_g19065(csa_tree_add_12_51_groupi_n_2706 ,csa_tree_add_12_51_groupi_n_469 ,csa_tree_add_12_51_groupi_n_2201);
  or csa_tree_add_12_51_groupi_g19066(csa_tree_add_12_51_groupi_n_2705 ,in4[8] ,csa_tree_add_12_51_groupi_n_2486);
  or csa_tree_add_12_51_groupi_g19067(csa_tree_add_12_51_groupi_n_2704 ,csa_tree_add_12_51_groupi_n_1896 ,csa_tree_add_12_51_groupi_n_2496);
  or csa_tree_add_12_51_groupi_g19068(csa_tree_add_12_51_groupi_n_2703 ,in2[5] ,csa_tree_add_12_51_groupi_n_2483);
  nor csa_tree_add_12_51_groupi_g19069(csa_tree_add_12_51_groupi_n_2702 ,csa_tree_add_12_51_groupi_n_1286 ,csa_tree_add_12_51_groupi_n_355);
  or csa_tree_add_12_51_groupi_g19070(csa_tree_add_12_51_groupi_n_2701 ,csa_tree_add_12_51_groupi_n_122 ,csa_tree_add_12_51_groupi_n_2484);
  or csa_tree_add_12_51_groupi_g19071(csa_tree_add_12_51_groupi_n_2700 ,in3[2] ,csa_tree_add_12_51_groupi_n_2490);
  or csa_tree_add_12_51_groupi_g19072(csa_tree_add_12_51_groupi_n_2699 ,csa_tree_add_12_51_groupi_n_125 ,csa_tree_add_12_51_groupi_n_2495);
  or csa_tree_add_12_51_groupi_g19073(csa_tree_add_12_51_groupi_n_2698 ,csa_tree_add_12_51_groupi_n_2373 ,csa_tree_add_12_51_groupi_n_2517);
  or csa_tree_add_12_51_groupi_g19074(csa_tree_add_12_51_groupi_n_2697 ,csa_tree_add_12_51_groupi_n_1926 ,csa_tree_add_12_51_groupi_n_2498);
  or csa_tree_add_12_51_groupi_g19075(csa_tree_add_12_51_groupi_n_2696 ,csa_tree_add_12_51_groupi_n_114 ,csa_tree_add_12_51_groupi_n_2500);
  or csa_tree_add_12_51_groupi_g19076(csa_tree_add_12_51_groupi_n_2695 ,in2[11] ,csa_tree_add_12_51_groupi_n_2485);
  nor csa_tree_add_12_51_groupi_g19077(csa_tree_add_12_51_groupi_n_2694 ,csa_tree_add_12_51_groupi_n_1499 ,csa_tree_add_12_51_groupi_n_283);
  or csa_tree_add_12_51_groupi_g19078(csa_tree_add_12_51_groupi_n_2693 ,csa_tree_add_12_51_groupi_n_2402 ,csa_tree_add_12_51_groupi_n_2481);
  or csa_tree_add_12_51_groupi_g19079(csa_tree_add_12_51_groupi_n_2692 ,in4[2] ,csa_tree_add_12_51_groupi_n_2493);
  nor csa_tree_add_12_51_groupi_g19080(csa_tree_add_12_51_groupi_n_2691 ,csa_tree_add_12_51_groupi_n_1682 ,csa_tree_add_12_51_groupi_n_274);
  nor csa_tree_add_12_51_groupi_g19081(csa_tree_add_12_51_groupi_n_2690 ,csa_tree_add_12_51_groupi_n_1499 ,csa_tree_add_12_51_groupi_n_387);
  or csa_tree_add_12_51_groupi_g19082(csa_tree_add_12_51_groupi_n_2689 ,csa_tree_add_12_51_groupi_n_2365 ,csa_tree_add_12_51_groupi_n_2488);
  nor csa_tree_add_12_51_groupi_g19083(csa_tree_add_12_51_groupi_n_2688 ,csa_tree_add_12_51_groupi_n_472 ,csa_tree_add_12_51_groupi_n_2168);
  nor csa_tree_add_12_51_groupi_g19084(csa_tree_add_12_51_groupi_n_2687 ,csa_tree_add_12_51_groupi_n_1307 ,csa_tree_add_12_51_groupi_n_391);
  or csa_tree_add_12_51_groupi_g19085(csa_tree_add_12_51_groupi_n_2686 ,in2[2] ,csa_tree_add_12_51_groupi_n_2480);
  or csa_tree_add_12_51_groupi_g19086(csa_tree_add_12_51_groupi_n_2685 ,csa_tree_add_12_51_groupi_n_2467 ,csa_tree_add_12_51_groupi_n_2438);
  or csa_tree_add_12_51_groupi_g19087(csa_tree_add_12_51_groupi_n_2684 ,in4[11] ,csa_tree_add_12_51_groupi_n_2497);
  or csa_tree_add_12_51_groupi_g19088(csa_tree_add_12_51_groupi_n_2683 ,in4[5] ,csa_tree_add_12_51_groupi_n_2482);
  or csa_tree_add_12_51_groupi_g19089(csa_tree_add_12_51_groupi_n_2682 ,in3[14] ,csa_tree_add_12_51_groupi_n_2450);
  nor csa_tree_add_12_51_groupi_g19090(csa_tree_add_12_51_groupi_n_2681 ,in3[11] ,csa_tree_add_12_51_groupi_n_2471);
  or csa_tree_add_12_51_groupi_g19091(csa_tree_add_12_51_groupi_n_2680 ,in3[5] ,csa_tree_add_12_51_groupi_n_2474);
  or csa_tree_add_12_51_groupi_g19092(csa_tree_add_12_51_groupi_n_2679 ,in3[8] ,csa_tree_add_12_51_groupi_n_2444);
  nor csa_tree_add_12_51_groupi_g19093(csa_tree_add_12_51_groupi_n_2678 ,csa_tree_add_12_51_groupi_n_1350 ,csa_tree_add_12_51_groupi_n_140);
  nor csa_tree_add_12_51_groupi_g19094(csa_tree_add_12_51_groupi_n_2677 ,csa_tree_add_12_51_groupi_n_1683 ,csa_tree_add_12_51_groupi_n_148);
  nor csa_tree_add_12_51_groupi_g19095(csa_tree_add_12_51_groupi_n_2676 ,csa_tree_add_12_51_groupi_n_408 ,csa_tree_add_12_51_groupi_n_2172);
  nor csa_tree_add_12_51_groupi_g19096(csa_tree_add_12_51_groupi_n_2675 ,csa_tree_add_12_51_groupi_n_1578 ,csa_tree_add_12_51_groupi_n_700);
  nor csa_tree_add_12_51_groupi_g19097(csa_tree_add_12_51_groupi_n_2674 ,csa_tree_add_12_51_groupi_n_1046 ,csa_tree_add_12_51_groupi_n_2199);
  nor csa_tree_add_12_51_groupi_g19098(csa_tree_add_12_51_groupi_n_2673 ,csa_tree_add_12_51_groupi_n_1050 ,csa_tree_add_12_51_groupi_n_1356);
  nor csa_tree_add_12_51_groupi_g19099(csa_tree_add_12_51_groupi_n_2672 ,csa_tree_add_12_51_groupi_n_1653 ,csa_tree_add_12_51_groupi_n_304);
  nor csa_tree_add_12_51_groupi_g19100(csa_tree_add_12_51_groupi_n_2671 ,csa_tree_add_12_51_groupi_n_436 ,csa_tree_add_12_51_groupi_n_2168);
  nor csa_tree_add_12_51_groupi_g19101(csa_tree_add_12_51_groupi_n_2670 ,csa_tree_add_12_51_groupi_n_1353 ,csa_tree_add_12_51_groupi_n_259);
  nor csa_tree_add_12_51_groupi_g19102(csa_tree_add_12_51_groupi_n_2669 ,csa_tree_add_12_51_groupi_n_1683 ,csa_tree_add_12_51_groupi_n_256);
  nor csa_tree_add_12_51_groupi_g19103(csa_tree_add_12_51_groupi_n_2668 ,csa_tree_add_12_51_groupi_n_1677 ,csa_tree_add_12_51_groupi_n_289);
  nor csa_tree_add_12_51_groupi_g19104(csa_tree_add_12_51_groupi_n_2667 ,csa_tree_add_12_51_groupi_n_480 ,csa_tree_add_12_51_groupi_n_2201);
  nor csa_tree_add_12_51_groupi_g19105(csa_tree_add_12_51_groupi_n_2666 ,csa_tree_add_12_51_groupi_n_525 ,csa_tree_add_12_51_groupi_n_1350);
  nor csa_tree_add_12_51_groupi_g19106(csa_tree_add_12_51_groupi_n_2665 ,csa_tree_add_12_51_groupi_n_1815 ,csa_tree_add_12_51_groupi_n_1571);
  nor csa_tree_add_12_51_groupi_g19107(csa_tree_add_12_51_groupi_n_2664 ,csa_tree_add_12_51_groupi_n_1218 ,csa_tree_add_12_51_groupi_n_216);
  or csa_tree_add_12_51_groupi_g19108(csa_tree_add_12_51_groupi_n_2781 ,csa_tree_add_12_51_groupi_n_2530 ,csa_tree_add_12_51_groupi_n_2533);
  or csa_tree_add_12_51_groupi_g19109(csa_tree_add_12_51_groupi_n_2779 ,csa_tree_add_12_51_groupi_n_2510 ,csa_tree_add_12_51_groupi_n_2475);
  or csa_tree_add_12_51_groupi_g19110(csa_tree_add_12_51_groupi_n_2777 ,csa_tree_add_12_51_groupi_n_2538 ,csa_tree_add_12_51_groupi_n_2523);
  or csa_tree_add_12_51_groupi_g19111(csa_tree_add_12_51_groupi_n_2775 ,csa_tree_add_12_51_groupi_n_2518 ,csa_tree_add_12_51_groupi_n_2511);
  or csa_tree_add_12_51_groupi_g19112(csa_tree_add_12_51_groupi_n_2773 ,csa_tree_add_12_51_groupi_n_2516 ,csa_tree_add_12_51_groupi_n_2513);
  or csa_tree_add_12_51_groupi_g19113(csa_tree_add_12_51_groupi_n_2771 ,csa_tree_add_12_51_groupi_n_2470 ,csa_tree_add_12_51_groupi_n_2507);
  or csa_tree_add_12_51_groupi_g19114(csa_tree_add_12_51_groupi_n_2769 ,csa_tree_add_12_51_groupi_n_2532 ,csa_tree_add_12_51_groupi_n_2527);
  or csa_tree_add_12_51_groupi_g19115(csa_tree_add_12_51_groupi_n_2767 ,csa_tree_add_12_51_groupi_n_2546 ,csa_tree_add_12_51_groupi_n_2541);
  or csa_tree_add_12_51_groupi_g19116(csa_tree_add_12_51_groupi_n_2765 ,csa_tree_add_12_51_groupi_n_2522 ,csa_tree_add_12_51_groupi_n_2519);
  or csa_tree_add_12_51_groupi_g19117(csa_tree_add_12_51_groupi_n_2763 ,csa_tree_add_12_51_groupi_n_2526 ,csa_tree_add_12_51_groupi_n_2535);
  or csa_tree_add_12_51_groupi_g19118(csa_tree_add_12_51_groupi_n_2761 ,csa_tree_add_12_51_groupi_n_2544 ,csa_tree_add_12_51_groupi_n_2539);
  or csa_tree_add_12_51_groupi_g19119(csa_tree_add_12_51_groupi_n_2759 ,csa_tree_add_12_51_groupi_n_2548 ,csa_tree_add_12_51_groupi_n_2549);
  or csa_tree_add_12_51_groupi_g19120(csa_tree_add_12_51_groupi_n_2758 ,csa_tree_add_12_51_groupi_n_1262 ,csa_tree_add_12_51_groupi_n_2165);
  and csa_tree_add_12_51_groupi_g19121(csa_tree_add_12_51_groupi_n_2756 ,in1[15] ,csa_tree_add_12_51_groupi_n_1905);
  or csa_tree_add_12_51_groupi_g19122(csa_tree_add_12_51_groupi_n_2755 ,csa_tree_add_12_51_groupi_n_1265 ,csa_tree_add_12_51_groupi_n_19);
  or csa_tree_add_12_51_groupi_g19123(csa_tree_add_12_51_groupi_n_2754 ,in3[0] ,csa_tree_add_12_51_groupi_n_2479);
  or csa_tree_add_12_51_groupi_g19124(csa_tree_add_12_51_groupi_n_2753 ,in2[0] ,csa_tree_add_12_51_groupi_n_2478);
  or csa_tree_add_12_51_groupi_g19125(csa_tree_add_12_51_groupi_n_2752 ,in4[0] ,csa_tree_add_12_51_groupi_n_2477);
  not csa_tree_add_12_51_groupi_g19126(csa_tree_add_12_51_groupi_n_2663 ,csa_tree_add_12_51_groupi_n_2662);
  not csa_tree_add_12_51_groupi_g19127(csa_tree_add_12_51_groupi_n_2661 ,csa_tree_add_12_51_groupi_n_2660);
  not csa_tree_add_12_51_groupi_g19128(csa_tree_add_12_51_groupi_n_2659 ,csa_tree_add_12_51_groupi_n_2658);
  not csa_tree_add_12_51_groupi_g19129(csa_tree_add_12_51_groupi_n_2649 ,csa_tree_add_12_51_groupi_n_2648);
  not csa_tree_add_12_51_groupi_g19130(csa_tree_add_12_51_groupi_n_2642 ,csa_tree_add_12_51_groupi_n_2641);
  not csa_tree_add_12_51_groupi_g19131(csa_tree_add_12_51_groupi_n_2640 ,csa_tree_add_12_51_groupi_n_1908);
  not csa_tree_add_12_51_groupi_g19133(csa_tree_add_12_51_groupi_n_2639 ,csa_tree_add_12_51_groupi_n_2641);
  nor csa_tree_add_12_51_groupi_g19134(csa_tree_add_12_51_groupi_n_2636 ,csa_tree_add_12_51_groupi_n_1677 ,csa_tree_add_12_51_groupi_n_352);
  nor csa_tree_add_12_51_groupi_g19135(csa_tree_add_12_51_groupi_n_2635 ,csa_tree_add_12_51_groupi_n_1214 ,csa_tree_add_12_51_groupi_n_418);
  nor csa_tree_add_12_51_groupi_g19136(csa_tree_add_12_51_groupi_n_2634 ,csa_tree_add_12_51_groupi_n_1676 ,csa_tree_add_12_51_groupi_n_403);
  nor csa_tree_add_12_51_groupi_g19137(csa_tree_add_12_51_groupi_n_2633 ,csa_tree_add_12_51_groupi_n_439 ,csa_tree_add_12_51_groupi_n_2166);
  nor csa_tree_add_12_51_groupi_g19138(csa_tree_add_12_51_groupi_n_2632 ,csa_tree_add_12_51_groupi_n_1449 ,csa_tree_add_12_51_groupi_n_2202);
  nor csa_tree_add_12_51_groupi_g19139(csa_tree_add_12_51_groupi_n_2631 ,csa_tree_add_12_51_groupi_n_454 ,csa_tree_add_12_51_groupi_n_2165);
  nor csa_tree_add_12_51_groupi_g19140(csa_tree_add_12_51_groupi_n_2630 ,csa_tree_add_12_51_groupi_n_1578 ,csa_tree_add_12_51_groupi_n_190);
  nor csa_tree_add_12_51_groupi_g19141(csa_tree_add_12_51_groupi_n_2629 ,csa_tree_add_12_51_groupi_n_1500 ,csa_tree_add_12_51_groupi_n_223);
  nor csa_tree_add_12_51_groupi_g19142(csa_tree_add_12_51_groupi_n_2628 ,csa_tree_add_12_51_groupi_n_1815 ,csa_tree_add_12_51_groupi_n_358);
  nor csa_tree_add_12_51_groupi_g19143(csa_tree_add_12_51_groupi_n_2627 ,csa_tree_add_12_51_groupi_n_1283 ,csa_tree_add_12_51_groupi_n_265);
  nor csa_tree_add_12_51_groupi_g19144(csa_tree_add_12_51_groupi_n_2626 ,csa_tree_add_12_51_groupi_n_496 ,csa_tree_add_12_51_groupi_n_2202);
  nor csa_tree_add_12_51_groupi_g19145(csa_tree_add_12_51_groupi_n_2625 ,csa_tree_add_12_51_groupi_n_1653 ,csa_tree_add_12_51_groupi_n_319);
  nor csa_tree_add_12_51_groupi_g19146(csa_tree_add_12_51_groupi_n_2624 ,csa_tree_add_12_51_groupi_n_493 ,csa_tree_add_12_51_groupi_n_1220);
  nor csa_tree_add_12_51_groupi_g19147(csa_tree_add_12_51_groupi_n_2623 ,csa_tree_add_12_51_groupi_n_433 ,csa_tree_add_12_51_groupi_n_2199);
  nor csa_tree_add_12_51_groupi_g19148(csa_tree_add_12_51_groupi_n_2622 ,csa_tree_add_12_51_groupi_n_1676 ,csa_tree_add_12_51_groupi_n_331);
  nor csa_tree_add_12_51_groupi_g19149(csa_tree_add_12_51_groupi_n_2621 ,csa_tree_add_12_51_groupi_n_1361 ,csa_tree_add_12_51_groupi_n_361);
  nor csa_tree_add_12_51_groupi_g19150(csa_tree_add_12_51_groupi_n_2620 ,csa_tree_add_12_51_groupi_n_445 ,csa_tree_add_12_51_groupi_n_2160);
  nor csa_tree_add_12_51_groupi_g19151(csa_tree_add_12_51_groupi_n_2619 ,csa_tree_add_12_51_groupi_n_475 ,csa_tree_add_12_51_groupi_n_2159);
  nor csa_tree_add_12_51_groupi_g19152(csa_tree_add_12_51_groupi_n_2618 ,csa_tree_add_12_51_groupi_n_1308 ,csa_tree_add_12_51_groupi_n_370);
  nor csa_tree_add_12_51_groupi_g19153(csa_tree_add_12_51_groupi_n_2617 ,csa_tree_add_12_51_groupi_n_535 ,csa_tree_add_12_51_groupi_n_1308);
  nor csa_tree_add_12_51_groupi_g19154(csa_tree_add_12_51_groupi_n_2616 ,csa_tree_add_12_51_groupi_n_1577 ,csa_tree_add_12_51_groupi_n_1269);
  nor csa_tree_add_12_51_groupi_g19155(csa_tree_add_12_51_groupi_n_2615 ,csa_tree_add_12_51_groupi_n_486 ,csa_tree_add_12_51_groupi_n_2198);
  nor csa_tree_add_12_51_groupi_g19156(csa_tree_add_12_51_groupi_n_2614 ,csa_tree_add_12_51_groupi_n_1284 ,csa_tree_add_12_51_groupi_n_226);
  nor csa_tree_add_12_51_groupi_g19157(csa_tree_add_12_51_groupi_n_2613 ,csa_tree_add_12_51_groupi_n_582 ,csa_tree_add_12_51_groupi_n_1221);
  nor csa_tree_add_12_51_groupi_g19158(csa_tree_add_12_51_groupi_n_2612 ,csa_tree_add_12_51_groupi_n_1652 ,csa_tree_add_12_51_groupi_n_328);
  nor csa_tree_add_12_51_groupi_g19159(csa_tree_add_12_51_groupi_n_2611 ,csa_tree_add_12_51_groupi_n_1355 ,csa_tree_add_12_51_groupi_n_312);
  nor csa_tree_add_12_51_groupi_g19160(csa_tree_add_12_51_groupi_n_2610 ,csa_tree_add_12_51_groupi_n_460 ,csa_tree_add_12_51_groupi_n_2171);
  nor csa_tree_add_12_51_groupi_g19161(csa_tree_add_12_51_groupi_n_2609 ,csa_tree_add_12_51_groupi_n_1397 ,csa_tree_add_12_51_groupi_n_2174);
  nor csa_tree_add_12_51_groupi_g19162(csa_tree_add_12_51_groupi_n_2608 ,csa_tree_add_12_51_groupi_n_1425 ,csa_tree_add_12_51_groupi_n_2172);
  nor csa_tree_add_12_51_groupi_g19163(csa_tree_add_12_51_groupi_n_2607 ,csa_tree_add_12_51_groupi_n_1356 ,csa_tree_add_12_51_groupi_n_396);
  nor csa_tree_add_12_51_groupi_g19164(csa_tree_add_12_51_groupi_n_2606 ,csa_tree_add_12_51_groupi_n_691 ,csa_tree_add_12_51_groupi_n_1361);
  nor csa_tree_add_12_51_groupi_g19165(csa_tree_add_12_51_groupi_n_2605 ,csa_tree_add_12_51_groupi_n_501 ,csa_tree_add_12_51_groupi_n_1500);
  nor csa_tree_add_12_51_groupi_g19166(csa_tree_add_12_51_groupi_n_2604 ,csa_tree_add_12_51_groupi_n_1451 ,csa_tree_add_12_51_groupi_n_1355);
  nor csa_tree_add_12_51_groupi_g19167(csa_tree_add_12_51_groupi_n_2603 ,csa_tree_add_12_51_groupi_n_621 ,csa_tree_add_12_51_groupi_n_1307);
  nor csa_tree_add_12_51_groupi_g19168(csa_tree_add_12_51_groupi_n_2602 ,csa_tree_add_12_51_groupi_n_676 ,csa_tree_add_12_51_groupi_n_1217);
  nor csa_tree_add_12_51_groupi_g19169(csa_tree_add_12_51_groupi_n_2601 ,csa_tree_add_12_51_groupi_n_1362 ,csa_tree_add_12_51_groupi_n_364);
  nor csa_tree_add_12_51_groupi_g19170(csa_tree_add_12_51_groupi_n_2600 ,csa_tree_add_12_51_groupi_n_1349 ,csa_tree_add_12_51_groupi_n_316);
  nor csa_tree_add_12_51_groupi_g19171(csa_tree_add_12_51_groupi_n_2599 ,csa_tree_add_12_51_groupi_n_684 ,csa_tree_add_12_51_groupi_n_1362);
  nor csa_tree_add_12_51_groupi_g19172(csa_tree_add_12_51_groupi_n_2598 ,csa_tree_add_12_51_groupi_n_1694 ,csa_tree_add_12_51_groupi_n_2196);
  nor csa_tree_add_12_51_groupi_g19173(csa_tree_add_12_51_groupi_n_2597 ,csa_tree_add_12_51_groupi_n_1461 ,csa_tree_add_12_51_groupi_n_2171);
  nor csa_tree_add_12_51_groupi_g19174(csa_tree_add_12_51_groupi_n_2596 ,csa_tree_add_12_51_groupi_n_499 ,csa_tree_add_12_51_groupi_n_1220);
  nor csa_tree_add_12_51_groupi_g19175(csa_tree_add_12_51_groupi_n_2595 ,csa_tree_add_12_51_groupi_n_478 ,csa_tree_add_12_51_groupi_n_2169);
  nor csa_tree_add_12_51_groupi_g19176(csa_tree_add_12_51_groupi_n_2594 ,csa_tree_add_12_51_groupi_n_571 ,csa_tree_add_12_51_groupi_n_1215);
  nor csa_tree_add_12_51_groupi_g19177(csa_tree_add_12_51_groupi_n_2593 ,csa_tree_add_12_51_groupi_n_1428 ,csa_tree_add_12_51_groupi_n_1218);
  nor csa_tree_add_12_51_groupi_g19178(csa_tree_add_12_51_groupi_n_2592 ,csa_tree_add_12_51_groupi_n_1769 ,csa_tree_add_12_51_groupi_n_1215);
  nor csa_tree_add_12_51_groupi_g19179(csa_tree_add_12_51_groupi_n_2591 ,csa_tree_add_12_51_groupi_n_1457 ,csa_tree_add_12_51_groupi_n_1287);
  nor csa_tree_add_12_51_groupi_g19180(csa_tree_add_12_51_groupi_n_2590 ,csa_tree_add_12_51_groupi_n_1430 ,csa_tree_add_12_51_groupi_n_2160);
  nor csa_tree_add_12_51_groupi_g19181(csa_tree_add_12_51_groupi_n_2589 ,csa_tree_add_12_51_groupi_n_1808 ,csa_tree_add_12_51_groupi_n_1349);
  nor csa_tree_add_12_51_groupi_g19182(csa_tree_add_12_51_groupi_n_2588 ,csa_tree_add_12_51_groupi_n_1415 ,csa_tree_add_12_51_groupi_n_1284);
  nor csa_tree_add_12_51_groupi_g19183(csa_tree_add_12_51_groupi_n_2587 ,csa_tree_add_12_51_groupi_n_511 ,csa_tree_add_12_51_groupi_n_1283);
  nor csa_tree_add_12_51_groupi_g19184(csa_tree_add_12_51_groupi_n_2586 ,csa_tree_add_12_51_groupi_n_1724 ,csa_tree_add_12_51_groupi_n_1352);
  nor csa_tree_add_12_51_groupi_g19185(csa_tree_add_12_51_groupi_n_2585 ,csa_tree_add_12_51_groupi_n_484 ,csa_tree_add_12_51_groupi_n_1287);
  nor csa_tree_add_12_51_groupi_g19186(csa_tree_add_12_51_groupi_n_2584 ,csa_tree_add_12_51_groupi_n_1781 ,csa_tree_add_12_51_groupi_n_2175);
  nor csa_tree_add_12_51_groupi_g19187(csa_tree_add_12_51_groupi_n_2583 ,csa_tree_add_12_51_groupi_n_1814 ,csa_tree_add_12_51_groupi_n_1565);
  nor csa_tree_add_12_51_groupi_g19188(csa_tree_add_12_51_groupi_n_2582 ,csa_tree_add_12_51_groupi_n_1706 ,csa_tree_add_12_51_groupi_n_2166);
  nor csa_tree_add_12_51_groupi_g19189(csa_tree_add_12_51_groupi_n_2581 ,csa_tree_add_12_51_groupi_n_1733 ,csa_tree_add_12_51_groupi_n_2175);
  nor csa_tree_add_12_51_groupi_g19190(csa_tree_add_12_51_groupi_n_2580 ,csa_tree_add_12_51_groupi_n_1793 ,csa_tree_add_12_51_groupi_n_1217);
  nor csa_tree_add_12_51_groupi_g19191(csa_tree_add_12_51_groupi_n_2579 ,csa_tree_add_12_51_groupi_n_660 ,csa_tree_add_12_51_groupi_n_1352);
  nor csa_tree_add_12_51_groupi_g19192(csa_tree_add_12_51_groupi_n_2578 ,csa_tree_add_12_51_groupi_n_1748 ,csa_tree_add_12_51_groupi_n_2174);
  nor csa_tree_add_12_51_groupi_g19193(csa_tree_add_12_51_groupi_n_2577 ,csa_tree_add_12_51_groupi_n_1712 ,csa_tree_add_12_51_groupi_n_1214);
  nor csa_tree_add_12_51_groupi_g19194(csa_tree_add_12_51_groupi_n_2576 ,csa_tree_add_12_51_groupi_n_1811 ,csa_tree_add_12_51_groupi_n_2195);
  nor csa_tree_add_12_51_groupi_g19195(csa_tree_add_12_51_groupi_n_2575 ,csa_tree_add_12_51_groupi_n_1577 ,csa_tree_add_12_51_groupi_n_1569);
  nor csa_tree_add_12_51_groupi_g19196(csa_tree_add_12_51_groupi_n_2574 ,csa_tree_add_12_51_groupi_n_1742 ,csa_tree_add_12_51_groupi_n_2195);
  xnor csa_tree_add_12_51_groupi_g19197(csa_tree_add_12_51_groupi_n_2573 ,in4[8] ,in5[6]);
  xnor csa_tree_add_12_51_groupi_g19198(csa_tree_add_12_51_groupi_n_2572 ,in3[14] ,in5[12]);
  xnor csa_tree_add_12_51_groupi_g19199(csa_tree_add_12_51_groupi_n_2571 ,in4[14] ,in3[14]);
  xnor csa_tree_add_12_51_groupi_g19200(csa_tree_add_12_51_groupi_n_2662 ,csa_tree_add_12_51_groupi_n_120 ,in4[1]);
  xnor csa_tree_add_12_51_groupi_g19201(csa_tree_add_12_51_groupi_n_2660 ,csa_tree_add_12_51_groupi_n_110 ,in2[1]);
  xnor csa_tree_add_12_51_groupi_g19202(csa_tree_add_12_51_groupi_n_2658 ,csa_tree_add_12_51_groupi_n_106 ,in3[1]);
  xnor csa_tree_add_12_51_groupi_g19203(csa_tree_add_12_51_groupi_n_2570 ,in1[13] ,in1[12]);
  xnor csa_tree_add_12_51_groupi_g19204(csa_tree_add_12_51_groupi_n_2569 ,in1[8] ,in1[7]);
  xnor csa_tree_add_12_51_groupi_g19205(csa_tree_add_12_51_groupi_n_2568 ,in1[15] ,in1[14]);
  xnor csa_tree_add_12_51_groupi_g19206(csa_tree_add_12_51_groupi_n_2567 ,in1[12] ,in1[11]);
  xnor csa_tree_add_12_51_groupi_g19207(csa_tree_add_12_51_groupi_n_2566 ,in1[10] ,in1[9]);
  xnor csa_tree_add_12_51_groupi_g19208(csa_tree_add_12_51_groupi_n_2565 ,in1[2] ,in1[1]);
  xnor csa_tree_add_12_51_groupi_g19209(csa_tree_add_12_51_groupi_n_2564 ,in1[14] ,in1[13]);
  xnor csa_tree_add_12_51_groupi_g19210(csa_tree_add_12_51_groupi_n_2563 ,in1[9] ,in1[8]);
  xnor csa_tree_add_12_51_groupi_g19211(csa_tree_add_12_51_groupi_n_2562 ,in1[5] ,in1[4]);
  xnor csa_tree_add_12_51_groupi_g19212(csa_tree_add_12_51_groupi_n_2561 ,in1[3] ,in1[2]);
  xnor csa_tree_add_12_51_groupi_g19213(csa_tree_add_12_51_groupi_n_2560 ,in1[7] ,in1[6]);
  xnor csa_tree_add_12_51_groupi_g19214(csa_tree_add_12_51_groupi_n_2559 ,in1[4] ,in1[3]);
  xnor csa_tree_add_12_51_groupi_g19215(csa_tree_add_12_51_groupi_n_2558 ,in1[6] ,in1[5]);
  xnor csa_tree_add_12_51_groupi_g19216(csa_tree_add_12_51_groupi_n_2557 ,in1[11] ,in1[10]);
  xnor csa_tree_add_12_51_groupi_g19217(csa_tree_add_12_51_groupi_n_2657 ,in2[9] ,in2[8]);
  xnor csa_tree_add_12_51_groupi_g19218(csa_tree_add_12_51_groupi_n_2656 ,in2[6] ,in2[5]);
  xnor csa_tree_add_12_51_groupi_g19219(csa_tree_add_12_51_groupi_n_2655 ,in4[9] ,in4[8]);
  xnor csa_tree_add_12_51_groupi_g19220(csa_tree_add_12_51_groupi_n_2556 ,in4[8] ,in2[8]);
  xnor csa_tree_add_12_51_groupi_g19221(csa_tree_add_12_51_groupi_n_2654 ,in3[9] ,in3[8]);
  xnor csa_tree_add_12_51_groupi_g19222(csa_tree_add_12_51_groupi_n_2653 ,in3[12] ,in3[11]);
  xnor csa_tree_add_12_51_groupi_g19223(csa_tree_add_12_51_groupi_n_2555 ,in4[5] ,in3[5]);
  xnor csa_tree_add_12_51_groupi_g19224(csa_tree_add_12_51_groupi_n_2652 ,in4[3] ,in4[2]);
  xnor csa_tree_add_12_51_groupi_g19225(csa_tree_add_12_51_groupi_n_2651 ,in3[6] ,in3[5]);
  xnor csa_tree_add_12_51_groupi_g19226(csa_tree_add_12_51_groupi_n_2650 ,in2[3] ,in2[2]);
  xnor csa_tree_add_12_51_groupi_g19227(csa_tree_add_12_51_groupi_n_2648 ,csa_tree_add_12_51_groupi_n_1926 ,in2[2]);
  xnor csa_tree_add_12_51_groupi_g19228(csa_tree_add_12_51_groupi_n_2554 ,in2[11] ,in5[9]);
  xnor csa_tree_add_12_51_groupi_g19229(csa_tree_add_12_51_groupi_n_2647 ,in4[12] ,in4[11]);
  xnor csa_tree_add_12_51_groupi_g19230(csa_tree_add_12_51_groupi_n_2646 ,in3[3] ,in3[2]);
  xnor csa_tree_add_12_51_groupi_g19231(csa_tree_add_12_51_groupi_n_2553 ,in4[5] ,in5[3]);
  xnor csa_tree_add_12_51_groupi_g19232(csa_tree_add_12_51_groupi_n_2645 ,in2[12] ,in2[11]);
  xnor csa_tree_add_12_51_groupi_g19233(csa_tree_add_12_51_groupi_n_2552 ,in3[2] ,in5[0]);
  xnor csa_tree_add_12_51_groupi_g19234(csa_tree_add_12_51_groupi_n_2551 ,in4[11] ,in2[11]);
  xnor csa_tree_add_12_51_groupi_g19235(csa_tree_add_12_51_groupi_n_2644 ,in4[6] ,in4[5]);
  xnor csa_tree_add_12_51_groupi_g19236(csa_tree_add_12_51_groupi_n_2643 ,in1[1] ,in1[0]);
  and csa_tree_add_12_51_groupi_g19237(csa_tree_add_12_51_groupi_n_2641 ,csa_tree_add_12_51_groupi_n_19 ,csa_tree_add_12_51_groupi_n_2457);
  or csa_tree_add_12_51_groupi_g19238(csa_tree_add_12_51_groupi_n_2638 ,csa_tree_add_12_51_groupi_n_1907 ,csa_tree_add_12_51_groupi_n_2455);
  or csa_tree_add_12_51_groupi_g19239(csa_tree_add_12_51_groupi_n_2637 ,csa_tree_add_12_51_groupi_n_1906 ,csa_tree_add_12_51_groupi_n_2454);
  not csa_tree_add_12_51_groupi_g19240(csa_tree_add_12_51_groupi_n_2550 ,csa_tree_add_12_51_groupi_n_2549);
  not csa_tree_add_12_51_groupi_g19241(csa_tree_add_12_51_groupi_n_2548 ,csa_tree_add_12_51_groupi_n_2547);
  not csa_tree_add_12_51_groupi_g19242(csa_tree_add_12_51_groupi_n_2546 ,csa_tree_add_12_51_groupi_n_2545);
  not csa_tree_add_12_51_groupi_g19243(csa_tree_add_12_51_groupi_n_2544 ,csa_tree_add_12_51_groupi_n_2543);
  not csa_tree_add_12_51_groupi_g19244(csa_tree_add_12_51_groupi_n_2542 ,csa_tree_add_12_51_groupi_n_2541);
  not csa_tree_add_12_51_groupi_g19245(csa_tree_add_12_51_groupi_n_2540 ,csa_tree_add_12_51_groupi_n_2539);
  not csa_tree_add_12_51_groupi_g19246(csa_tree_add_12_51_groupi_n_2538 ,csa_tree_add_12_51_groupi_n_2537);
  not csa_tree_add_12_51_groupi_g19247(csa_tree_add_12_51_groupi_n_2536 ,csa_tree_add_12_51_groupi_n_2535);
  not csa_tree_add_12_51_groupi_g19248(csa_tree_add_12_51_groupi_n_2534 ,csa_tree_add_12_51_groupi_n_2533);
  not csa_tree_add_12_51_groupi_g19249(csa_tree_add_12_51_groupi_n_2532 ,csa_tree_add_12_51_groupi_n_2531);
  not csa_tree_add_12_51_groupi_g19250(csa_tree_add_12_51_groupi_n_2530 ,csa_tree_add_12_51_groupi_n_2529);
  not csa_tree_add_12_51_groupi_g19251(csa_tree_add_12_51_groupi_n_2528 ,csa_tree_add_12_51_groupi_n_2527);
  not csa_tree_add_12_51_groupi_g19252(csa_tree_add_12_51_groupi_n_2526 ,csa_tree_add_12_51_groupi_n_2525);
  not csa_tree_add_12_51_groupi_g19253(csa_tree_add_12_51_groupi_n_2524 ,csa_tree_add_12_51_groupi_n_2523);
  not csa_tree_add_12_51_groupi_g19254(csa_tree_add_12_51_groupi_n_2522 ,csa_tree_add_12_51_groupi_n_2521);
  not csa_tree_add_12_51_groupi_g19255(csa_tree_add_12_51_groupi_n_2520 ,csa_tree_add_12_51_groupi_n_2519);
  not csa_tree_add_12_51_groupi_g19256(csa_tree_add_12_51_groupi_n_2518 ,csa_tree_add_12_51_groupi_n_2517);
  not csa_tree_add_12_51_groupi_g19257(csa_tree_add_12_51_groupi_n_2516 ,csa_tree_add_12_51_groupi_n_2515);
  not csa_tree_add_12_51_groupi_g19258(csa_tree_add_12_51_groupi_n_2514 ,csa_tree_add_12_51_groupi_n_2513);
  not csa_tree_add_12_51_groupi_g19259(csa_tree_add_12_51_groupi_n_2512 ,csa_tree_add_12_51_groupi_n_2511);
  not csa_tree_add_12_51_groupi_g19260(csa_tree_add_12_51_groupi_n_2510 ,csa_tree_add_12_51_groupi_n_2509);
  not csa_tree_add_12_51_groupi_g19261(csa_tree_add_12_51_groupi_n_2508 ,csa_tree_add_12_51_groupi_n_2507);
  or csa_tree_add_12_51_groupi_g19262(csa_tree_add_12_51_groupi_n_2503 ,csa_tree_add_12_51_groupi_n_2374 ,in4[7]);
  or csa_tree_add_12_51_groupi_g19263(csa_tree_add_12_51_groupi_n_2502 ,csa_tree_add_12_51_groupi_n_2413 ,in3[12]);
  or csa_tree_add_12_51_groupi_g19264(csa_tree_add_12_51_groupi_n_2501 ,csa_tree_add_12_51_groupi_n_2408 ,in2[9]);
  or csa_tree_add_12_51_groupi_g19265(csa_tree_add_12_51_groupi_n_2500 ,csa_tree_add_12_51_groupi_n_2370 ,in2[10]);
  or csa_tree_add_12_51_groupi_g19266(csa_tree_add_12_51_groupi_n_2499 ,csa_tree_add_12_51_groupi_n_2414 ,in3[9]);
  or csa_tree_add_12_51_groupi_g19267(csa_tree_add_12_51_groupi_n_2498 ,csa_tree_add_12_51_groupi_n_2406 ,in4[4]);
  or csa_tree_add_12_51_groupi_g19268(csa_tree_add_12_51_groupi_n_2497 ,csa_tree_add_12_51_groupi_n_2409 ,in4[12]);
  or csa_tree_add_12_51_groupi_g19269(csa_tree_add_12_51_groupi_n_2496 ,csa_tree_add_12_51_groupi_n_2368 ,in3[13]);
  or csa_tree_add_12_51_groupi_g19270(csa_tree_add_12_51_groupi_n_2495 ,csa_tree_add_12_51_groupi_n_2375 ,in4[10]);
  or csa_tree_add_12_51_groupi_g19271(csa_tree_add_12_51_groupi_n_2494 ,csa_tree_add_12_51_groupi_n_2377 ,in3[10]);
  or csa_tree_add_12_51_groupi_g19272(csa_tree_add_12_51_groupi_n_2493 ,csa_tree_add_12_51_groupi_n_2378 ,in4[3]);
  or csa_tree_add_12_51_groupi_g19273(csa_tree_add_12_51_groupi_n_2492 ,csa_tree_add_12_51_groupi_n_2369 ,in2[13]);
  or csa_tree_add_12_51_groupi_g19274(csa_tree_add_12_51_groupi_n_2491 ,csa_tree_add_12_51_groupi_n_2371 ,in3[7]);
  or csa_tree_add_12_51_groupi_g19275(csa_tree_add_12_51_groupi_n_2490 ,csa_tree_add_12_51_groupi_n_2410 ,in3[3]);
  or csa_tree_add_12_51_groupi_g19276(csa_tree_add_12_51_groupi_n_2489 ,csa_tree_add_12_51_groupi_n_2379 ,in3[6]);
  or csa_tree_add_12_51_groupi_g19277(csa_tree_add_12_51_groupi_n_2488 ,csa_tree_add_12_51_groupi_n_2405 ,in4[13]);
  or csa_tree_add_12_51_groupi_g19278(csa_tree_add_12_51_groupi_n_2487 ,csa_tree_add_12_51_groupi_n_2376 ,in2[4]);
  or csa_tree_add_12_51_groupi_g19279(csa_tree_add_12_51_groupi_n_2486 ,csa_tree_add_12_51_groupi_n_2381 ,in4[9]);
  or csa_tree_add_12_51_groupi_g19280(csa_tree_add_12_51_groupi_n_2485 ,csa_tree_add_12_51_groupi_n_2407 ,in2[12]);
  or csa_tree_add_12_51_groupi_g19281(csa_tree_add_12_51_groupi_n_2484 ,csa_tree_add_12_51_groupi_n_2373 ,in3[4]);
  or csa_tree_add_12_51_groupi_g19282(csa_tree_add_12_51_groupi_n_2483 ,csa_tree_add_12_51_groupi_n_2411 ,in2[6]);
  or csa_tree_add_12_51_groupi_g19283(csa_tree_add_12_51_groupi_n_2482 ,csa_tree_add_12_51_groupi_n_2412 ,in4[6]);
  or csa_tree_add_12_51_groupi_g19284(csa_tree_add_12_51_groupi_n_2481 ,csa_tree_add_12_51_groupi_n_2372 ,in2[7]);
  or csa_tree_add_12_51_groupi_g19285(csa_tree_add_12_51_groupi_n_2480 ,csa_tree_add_12_51_groupi_n_2384 ,in2[3]);
  and csa_tree_add_12_51_groupi_g19286(csa_tree_add_12_51_groupi_n_2549 ,in3[14] ,csa_tree_add_12_51_groupi_n_2413);
  or csa_tree_add_12_51_groupi_g19287(csa_tree_add_12_51_groupi_n_2547 ,csa_tree_add_12_51_groupi_n_2413 ,in3[14]);
  or csa_tree_add_12_51_groupi_g19288(csa_tree_add_12_51_groupi_n_2545 ,csa_tree_add_12_51_groupi_n_2407 ,in2[14]);
  or csa_tree_add_12_51_groupi_g19289(csa_tree_add_12_51_groupi_n_2543 ,csa_tree_add_12_51_groupi_n_2409 ,in4[14]);
  and csa_tree_add_12_51_groupi_g19290(csa_tree_add_12_51_groupi_n_2541 ,in2[14] ,csa_tree_add_12_51_groupi_n_2407);
  and csa_tree_add_12_51_groupi_g19291(csa_tree_add_12_51_groupi_n_2539 ,in4[14] ,csa_tree_add_12_51_groupi_n_2409);
  or csa_tree_add_12_51_groupi_g19292(csa_tree_add_12_51_groupi_n_2537 ,csa_tree_add_12_51_groupi_n_2408 ,in2[11]);
  and csa_tree_add_12_51_groupi_g19293(csa_tree_add_12_51_groupi_n_2535 ,in4[11] ,csa_tree_add_12_51_groupi_n_2381);
  and csa_tree_add_12_51_groupi_g19294(csa_tree_add_12_51_groupi_n_2533 ,in2[5] ,csa_tree_add_12_51_groupi_n_2384);
  or csa_tree_add_12_51_groupi_g19295(csa_tree_add_12_51_groupi_n_2531 ,csa_tree_add_12_51_groupi_n_2378 ,in4[5]);
  or csa_tree_add_12_51_groupi_g19296(csa_tree_add_12_51_groupi_n_2529 ,csa_tree_add_12_51_groupi_n_2384 ,in2[5]);
  and csa_tree_add_12_51_groupi_g19297(csa_tree_add_12_51_groupi_n_2527 ,in4[5] ,csa_tree_add_12_51_groupi_n_2378);
  or csa_tree_add_12_51_groupi_g19298(csa_tree_add_12_51_groupi_n_2525 ,csa_tree_add_12_51_groupi_n_2381 ,in4[11]);
  and csa_tree_add_12_51_groupi_g19299(csa_tree_add_12_51_groupi_n_2523 ,in2[11] ,csa_tree_add_12_51_groupi_n_2408);
  or csa_tree_add_12_51_groupi_g19300(csa_tree_add_12_51_groupi_n_2479 ,csa_tree_add_12_51_groupi_n_100 ,in3[1]);
  or csa_tree_add_12_51_groupi_g19301(csa_tree_add_12_51_groupi_n_2521 ,csa_tree_add_12_51_groupi_n_2414 ,in3[11]);
  and csa_tree_add_12_51_groupi_g19302(csa_tree_add_12_51_groupi_n_2519 ,in3[11] ,csa_tree_add_12_51_groupi_n_2414);
  or csa_tree_add_12_51_groupi_g19303(csa_tree_add_12_51_groupi_n_2517 ,csa_tree_add_12_51_groupi_n_2410 ,in3[5]);
  or csa_tree_add_12_51_groupi_g19304(csa_tree_add_12_51_groupi_n_2478 ,csa_tree_add_12_51_groupi_n_1942 ,in2[1]);
  or csa_tree_add_12_51_groupi_g19305(csa_tree_add_12_51_groupi_n_2477 ,csa_tree_add_12_51_groupi_n_1951 ,in4[1]);
  or csa_tree_add_12_51_groupi_g19306(csa_tree_add_12_51_groupi_n_2515 ,csa_tree_add_12_51_groupi_n_2379 ,in3[8]);
  and csa_tree_add_12_51_groupi_g19307(csa_tree_add_12_51_groupi_n_2513 ,in3[8] ,csa_tree_add_12_51_groupi_n_2379);
  and csa_tree_add_12_51_groupi_g19308(csa_tree_add_12_51_groupi_n_2511 ,in3[5] ,csa_tree_add_12_51_groupi_n_2410);
  or csa_tree_add_12_51_groupi_g19309(csa_tree_add_12_51_groupi_n_2509 ,csa_tree_add_12_51_groupi_n_2411 ,in2[8]);
  and csa_tree_add_12_51_groupi_g19310(csa_tree_add_12_51_groupi_n_2507 ,in4[8] ,csa_tree_add_12_51_groupi_n_2412);
  or csa_tree_add_12_51_groupi_g19311(csa_tree_add_12_51_groupi_n_2506 ,csa_tree_add_12_51_groupi_n_2415 ,in4[0]);
  or csa_tree_add_12_51_groupi_g19312(csa_tree_add_12_51_groupi_n_2505 ,csa_tree_add_12_51_groupi_n_2385 ,in3[0]);
  or csa_tree_add_12_51_groupi_g19313(csa_tree_add_12_51_groupi_n_2504 ,csa_tree_add_12_51_groupi_n_2386 ,in2[0]);
  not csa_tree_add_12_51_groupi_g19314(csa_tree_add_12_51_groupi_n_2476 ,csa_tree_add_12_51_groupi_n_2475);
  not csa_tree_add_12_51_groupi_g19315(csa_tree_add_12_51_groupi_n_2470 ,csa_tree_add_12_51_groupi_n_2469);
  not csa_tree_add_12_51_groupi_g19317(csa_tree_add_12_51_groupi_n_2465 ,csa_tree_add_12_51_groupi_n_1906);
  not csa_tree_add_12_51_groupi_g19319(csa_tree_add_12_51_groupi_n_2464 ,csa_tree_add_12_51_groupi_n_1905);
  not csa_tree_add_12_51_groupi_g19320(csa_tree_add_12_51_groupi_n_2462 ,csa_tree_add_12_51_groupi_n_1907);
  not csa_tree_add_12_51_groupi_g19322(csa_tree_add_12_51_groupi_n_2461 ,csa_tree_add_12_51_groupi_n_2460);
  or csa_tree_add_12_51_groupi_g19324(csa_tree_add_12_51_groupi_n_2459 ,csa_tree_add_12_51_groupi_n_1406 ,csa_tree_add_12_51_groupi_n_1412);
  nor csa_tree_add_12_51_groupi_g19325(csa_tree_add_12_51_groupi_n_2458 ,in1[11] ,in1[10]);
  or csa_tree_add_12_51_groupi_g19326(csa_tree_add_12_51_groupi_n_2457 ,in3[15] ,in3[14]);
  or csa_tree_add_12_51_groupi_g19327(csa_tree_add_12_51_groupi_n_2456 ,csa_tree_add_12_51_groupi_n_1460 ,csa_tree_add_12_51_groupi_n_1442);
  nor csa_tree_add_12_51_groupi_g19328(csa_tree_add_12_51_groupi_n_2455 ,in4[15] ,in4[14]);
  nor csa_tree_add_12_51_groupi_g19329(csa_tree_add_12_51_groupi_n_2454 ,in2[15] ,in2[14]);
  nor csa_tree_add_12_51_groupi_g19330(csa_tree_add_12_51_groupi_n_2453 ,csa_tree_add_12_51_groupi_n_1955 ,csa_tree_add_12_51_groupi_n_1899);
  or csa_tree_add_12_51_groupi_g19331(csa_tree_add_12_51_groupi_n_2452 ,in2[14] ,in3[14]);
  or csa_tree_add_12_51_groupi_g19332(csa_tree_add_12_51_groupi_n_2451 ,in4[14] ,in2[14]);
  nor csa_tree_add_12_51_groupi_g19333(csa_tree_add_12_51_groupi_n_2450 ,csa_tree_add_12_51_groupi_n_1918 ,csa_tree_add_12_51_groupi_n_1916);
  nor csa_tree_add_12_51_groupi_g19334(csa_tree_add_12_51_groupi_n_2449 ,csa_tree_add_12_51_groupi_n_123 ,csa_tree_add_12_51_groupi_n_1927);
  or csa_tree_add_12_51_groupi_g19335(csa_tree_add_12_51_groupi_n_2448 ,in4[2] ,in3[2]);
  nor csa_tree_add_12_51_groupi_g19336(csa_tree_add_12_51_groupi_n_2447 ,in1[7] ,in1[6]);
  nor csa_tree_add_12_51_groupi_g19337(csa_tree_add_12_51_groupi_n_2446 ,csa_tree_add_12_51_groupi_n_1957 ,csa_tree_add_12_51_groupi_n_1953);
  or csa_tree_add_12_51_groupi_g19338(csa_tree_add_12_51_groupi_n_2445 ,in4[8] ,in3[8]);
  nor csa_tree_add_12_51_groupi_g19339(csa_tree_add_12_51_groupi_n_2444 ,csa_tree_add_12_51_groupi_n_1938 ,csa_tree_add_12_51_groupi_n_1924);
  or csa_tree_add_12_51_groupi_g19340(csa_tree_add_12_51_groupi_n_2443 ,in4[8] ,in2[8]);
  nor csa_tree_add_12_51_groupi_g19341(csa_tree_add_12_51_groupi_n_2442 ,in1[3] ,in1[2]);
  nor csa_tree_add_12_51_groupi_g19342(csa_tree_add_12_51_groupi_n_2441 ,csa_tree_add_12_51_groupi_n_1778 ,csa_tree_add_12_51_groupi_n_1263);
  nor csa_tree_add_12_51_groupi_g19343(csa_tree_add_12_51_groupi_n_2440 ,in1[15] ,in1[14]);
  or csa_tree_add_12_51_groupi_g19344(csa_tree_add_12_51_groupi_n_2439 ,csa_tree_add_12_51_groupi_n_1418 ,csa_tree_add_12_51_groupi_n_1466);
  nor csa_tree_add_12_51_groupi_g19345(csa_tree_add_12_51_groupi_n_2438 ,in1[2] ,in1[1]);
  nor csa_tree_add_12_51_groupi_g19346(csa_tree_add_12_51_groupi_n_2437 ,in1[13] ,in1[12]);
  or csa_tree_add_12_51_groupi_g19347(csa_tree_add_12_51_groupi_n_2436 ,csa_tree_add_12_51_groupi_n_1472 ,csa_tree_add_12_51_groupi_n_1454);
  or csa_tree_add_12_51_groupi_g19348(csa_tree_add_12_51_groupi_n_2435 ,csa_tree_add_12_51_groupi_n_1448 ,csa_tree_add_12_51_groupi_n_1409);
  or csa_tree_add_12_51_groupi_g19349(csa_tree_add_12_51_groupi_n_2434 ,csa_tree_add_12_51_groupi_n_1457 ,csa_tree_add_12_51_groupi_n_1430);
  nor csa_tree_add_12_51_groupi_g19350(csa_tree_add_12_51_groupi_n_2433 ,in1[10] ,in1[9]);
  nor csa_tree_add_12_51_groupi_g19351(csa_tree_add_12_51_groupi_n_2432 ,in1[12] ,in1[11]);
  nor csa_tree_add_12_51_groupi_g19352(csa_tree_add_12_51_groupi_n_2431 ,in1[14] ,in1[13]);
  or csa_tree_add_12_51_groupi_g19353(csa_tree_add_12_51_groupi_n_2430 ,csa_tree_add_12_51_groupi_n_1415 ,csa_tree_add_12_51_groupi_n_1451);
  nor csa_tree_add_12_51_groupi_g19354(csa_tree_add_12_51_groupi_n_2429 ,in1[8] ,in1[7]);
  or csa_tree_add_12_51_groupi_g19355(csa_tree_add_12_51_groupi_n_2428 ,csa_tree_add_12_51_groupi_n_1436 ,csa_tree_add_12_51_groupi_n_1403);
  or csa_tree_add_12_51_groupi_g19356(csa_tree_add_12_51_groupi_n_2427 ,csa_tree_add_12_51_groupi_n_1445 ,csa_tree_add_12_51_groupi_n_1400);
  or csa_tree_add_12_51_groupi_g19357(csa_tree_add_12_51_groupi_n_2426 ,csa_tree_add_12_51_groupi_n_1424 ,csa_tree_add_12_51_groupi_n_1421);
  nor csa_tree_add_12_51_groupi_g19358(csa_tree_add_12_51_groupi_n_2425 ,in1[4] ,in1[3]);
  nor csa_tree_add_12_51_groupi_g19359(csa_tree_add_12_51_groupi_n_2424 ,in1[5] ,in1[4]);
  or csa_tree_add_12_51_groupi_g19360(csa_tree_add_12_51_groupi_n_2423 ,csa_tree_add_12_51_groupi_n_1433 ,csa_tree_add_12_51_groupi_n_1463);
  or csa_tree_add_12_51_groupi_g19361(csa_tree_add_12_51_groupi_n_2422 ,csa_tree_add_12_51_groupi_n_1397 ,csa_tree_add_12_51_groupi_n_1439);
  nor csa_tree_add_12_51_groupi_g19362(csa_tree_add_12_51_groupi_n_2421 ,in1[6] ,in1[5]);
  or csa_tree_add_12_51_groupi_g19363(csa_tree_add_12_51_groupi_n_2420 ,csa_tree_add_12_51_groupi_n_1268 ,csa_tree_add_12_51_groupi_n_1427);
  nor csa_tree_add_12_51_groupi_g19364(csa_tree_add_12_51_groupi_n_2419 ,in1[9] ,in1[8]);
  and csa_tree_add_12_51_groupi_g19365(csa_tree_add_12_51_groupi_n_2475 ,in2[8] ,csa_tree_add_12_51_groupi_n_2411);
  and csa_tree_add_12_51_groupi_g19366(csa_tree_add_12_51_groupi_n_2474 ,in4[5] ,in2[5]);
  and csa_tree_add_12_51_groupi_g19367(csa_tree_add_12_51_groupi_n_2473 ,csa_tree_add_12_51_groupi_n_2365 ,csa_tree_add_12_51_groupi_n_112);
  or csa_tree_add_12_51_groupi_g19368(csa_tree_add_12_51_groupi_n_2472 ,in4[5] ,in2[5]);
  and csa_tree_add_12_51_groupi_g19369(csa_tree_add_12_51_groupi_n_2471 ,in4[11] ,in2[11]);
  or csa_tree_add_12_51_groupi_g19370(csa_tree_add_12_51_groupi_n_2469 ,csa_tree_add_12_51_groupi_n_2412 ,in4[8]);
  and csa_tree_add_12_51_groupi_g19371(csa_tree_add_12_51_groupi_n_2468 ,csa_tree_add_12_51_groupi_n_120 ,csa_tree_add_12_51_groupi_n_104);
  or csa_tree_add_12_51_groupi_g19372(csa_tree_add_12_51_groupi_n_2467 ,csa_tree_add_12_51_groupi_n_1469 ,csa_tree_add_12_51_groupi_n_1046);
  and csa_tree_add_12_51_groupi_g19373(csa_tree_add_12_51_groupi_n_2466 ,in2[15] ,in2[14]);
  or csa_tree_add_12_51_groupi_g19374(csa_tree_add_12_51_groupi_n_2463 ,csa_tree_add_12_51_groupi_n_2418 ,csa_tree_add_12_51_groupi_n_108);
  and csa_tree_add_12_51_groupi_g19375(csa_tree_add_12_51_groupi_n_2460 ,in4[15] ,in4[14]);
  not csa_tree_add_12_51_groupi_g19376(csa_tree_add_12_51_groupi_n_2418 ,in3[15]);
  not csa_tree_add_12_51_groupi_g19377(csa_tree_add_12_51_groupi_n_2417 ,in5[15]);
  not csa_tree_add_12_51_groupi_g19378(csa_tree_add_12_51_groupi_n_2416 ,in5[9]);
  not csa_tree_add_12_51_groupi_g19379(csa_tree_add_12_51_groupi_n_2415 ,in4[1]);
  not csa_tree_add_12_51_groupi_g19380(csa_tree_add_12_51_groupi_n_2414 ,in3[10]);
  not csa_tree_add_12_51_groupi_g19381(csa_tree_add_12_51_groupi_n_2413 ,in3[13]);
  not csa_tree_add_12_51_groupi_g19382(csa_tree_add_12_51_groupi_n_2412 ,in4[7]);
  not csa_tree_add_12_51_groupi_g19383(csa_tree_add_12_51_groupi_n_2411 ,in2[7]);
  not csa_tree_add_12_51_groupi_g19384(csa_tree_add_12_51_groupi_n_2410 ,in3[4]);
  not csa_tree_add_12_51_groupi_g19385(csa_tree_add_12_51_groupi_n_2409 ,in4[13]);
  not csa_tree_add_12_51_groupi_g19386(csa_tree_add_12_51_groupi_n_2408 ,in2[10]);
  not csa_tree_add_12_51_groupi_g19387(csa_tree_add_12_51_groupi_n_2407 ,in2[13]);
  not csa_tree_add_12_51_groupi_g19388(csa_tree_add_12_51_groupi_n_2406 ,in4[3]);
  not csa_tree_add_12_51_groupi_g19389(csa_tree_add_12_51_groupi_n_2405 ,in4[12]);
  not csa_tree_add_12_51_groupi_g19390(csa_tree_add_12_51_groupi_n_2404 ,in3[14]);
  not csa_tree_add_12_51_groupi_g19391(csa_tree_add_12_51_groupi_n_2403 ,in2[11]);
  not csa_tree_add_12_51_groupi_g19392(csa_tree_add_12_51_groupi_n_2402 ,in2[5]);
  not csa_tree_add_12_51_groupi_g19393(csa_tree_add_12_51_groupi_n_2401 ,in4[5]);
  not csa_tree_add_12_51_groupi_g19394(csa_tree_add_12_51_groupi_n_2400 ,in3[8]);
  not csa_tree_add_12_51_groupi_g19395(csa_tree_add_12_51_groupi_n_2399 ,in2[2]);
  not csa_tree_add_12_51_groupi_g19396(csa_tree_add_12_51_groupi_n_2398 ,in4[8]);
  not csa_tree_add_12_51_groupi_g19397(csa_tree_add_12_51_groupi_n_2397 ,in2[8]);
  not csa_tree_add_12_51_groupi_g19398(csa_tree_add_12_51_groupi_n_2396 ,in1[15]);
  not csa_tree_add_12_51_groupi_g19399(csa_tree_add_12_51_groupi_n_2395 ,in1[1]);
  not csa_tree_add_12_51_groupi_g19400(csa_tree_add_12_51_groupi_n_2394 ,in1[11]);
  not csa_tree_add_12_51_groupi_g19401(csa_tree_add_12_51_groupi_n_2393 ,in1[13]);
  not csa_tree_add_12_51_groupi_g19402(csa_tree_add_12_51_groupi_n_2392 ,in1[14]);
  not csa_tree_add_12_51_groupi_g19403(csa_tree_add_12_51_groupi_n_2391 ,in1[5]);
  not csa_tree_add_12_51_groupi_g19404(csa_tree_add_12_51_groupi_n_2390 ,in1[10]);
  not csa_tree_add_12_51_groupi_g19405(csa_tree_add_12_51_groupi_n_2389 ,in1[8]);
  not csa_tree_add_12_51_groupi_g19406(csa_tree_add_12_51_groupi_n_2388 ,in1[12]);
  not csa_tree_add_12_51_groupi_g19407(csa_tree_add_12_51_groupi_n_2387 ,in1[3]);
  not csa_tree_add_12_51_groupi_g19408(csa_tree_add_12_51_groupi_n_2386 ,in2[1]);
  not csa_tree_add_12_51_groupi_g19409(csa_tree_add_12_51_groupi_n_2385 ,in3[1]);
  not csa_tree_add_12_51_groupi_g19410(csa_tree_add_12_51_groupi_n_2384 ,in2[4]);
  not csa_tree_add_12_51_groupi_g19411(csa_tree_add_12_51_groupi_n_2383 ,in4[0]);
  not csa_tree_add_12_51_groupi_g19412(csa_tree_add_12_51_groupi_n_2382 ,in2[0]);
  not csa_tree_add_12_51_groupi_g19413(csa_tree_add_12_51_groupi_n_2381 ,in4[10]);
  not csa_tree_add_12_51_groupi_g19414(csa_tree_add_12_51_groupi_n_2380 ,in3[0]);
  not csa_tree_add_12_51_groupi_g19415(csa_tree_add_12_51_groupi_n_2379 ,in3[7]);
  not csa_tree_add_12_51_groupi_g19416(csa_tree_add_12_51_groupi_n_2378 ,in4[4]);
  not csa_tree_add_12_51_groupi_g19417(csa_tree_add_12_51_groupi_n_2377 ,in3[9]);
  not csa_tree_add_12_51_groupi_g19418(csa_tree_add_12_51_groupi_n_2376 ,in2[3]);
  not csa_tree_add_12_51_groupi_g19419(csa_tree_add_12_51_groupi_n_2375 ,in4[9]);
  not csa_tree_add_12_51_groupi_g19420(csa_tree_add_12_51_groupi_n_2374 ,in4[6]);
  not csa_tree_add_12_51_groupi_g19421(csa_tree_add_12_51_groupi_n_2373 ,in3[3]);
  not csa_tree_add_12_51_groupi_g19422(csa_tree_add_12_51_groupi_n_2372 ,in2[6]);
  not csa_tree_add_12_51_groupi_g19423(csa_tree_add_12_51_groupi_n_2371 ,in3[6]);
  not csa_tree_add_12_51_groupi_g19424(csa_tree_add_12_51_groupi_n_2370 ,in2[9]);
  not csa_tree_add_12_51_groupi_g19425(csa_tree_add_12_51_groupi_n_2369 ,in2[12]);
  not csa_tree_add_12_51_groupi_g19426(csa_tree_add_12_51_groupi_n_2368 ,in3[12]);
  not csa_tree_add_12_51_groupi_g19427(csa_tree_add_12_51_groupi_n_2367 ,in2[14]);
  not csa_tree_add_12_51_groupi_g19428(csa_tree_add_12_51_groupi_n_2366 ,in4[14]);
  not csa_tree_add_12_51_groupi_g19429(csa_tree_add_12_51_groupi_n_2365 ,in4[11]);
  not csa_tree_add_12_51_groupi_g19430(csa_tree_add_12_51_groupi_n_2364 ,in3[2]);
  not csa_tree_add_12_51_groupi_g19431(csa_tree_add_12_51_groupi_n_2363 ,in4[2]);
  not csa_tree_add_12_51_groupi_g19432(csa_tree_add_12_51_groupi_n_2362 ,in3[5]);
  not csa_tree_add_12_51_groupi_g19433(csa_tree_add_12_51_groupi_n_2361 ,in3[11]);
  not csa_tree_add_12_51_groupi_g19434(csa_tree_add_12_51_groupi_n_2360 ,in1[0]);
  not csa_tree_add_12_51_groupi_g19435(csa_tree_add_12_51_groupi_n_2359 ,in1[2]);
  not csa_tree_add_12_51_groupi_g19436(csa_tree_add_12_51_groupi_n_2358 ,in1[6]);
  not csa_tree_add_12_51_groupi_g19437(csa_tree_add_12_51_groupi_n_2357 ,in1[4]);
  not csa_tree_add_12_51_groupi_g19438(csa_tree_add_12_51_groupi_n_2356 ,in1[7]);
  not csa_tree_add_12_51_groupi_g19439(csa_tree_add_12_51_groupi_n_2355 ,in1[9]);
  not csa_tree_add_12_51_groupi_drc_bufs(csa_tree_add_12_51_groupi_n_2346 ,csa_tree_add_12_51_groupi_n_723);
  not csa_tree_add_12_51_groupi_drc_bufs19440(csa_tree_add_12_51_groupi_n_2345 ,csa_tree_add_12_51_groupi_n_725);
  not csa_tree_add_12_51_groupi_drc_bufs19441(csa_tree_add_12_51_groupi_n_2344 ,csa_tree_add_12_51_groupi_n_724);
  not csa_tree_add_12_51_groupi_drc_bufs19442(csa_tree_add_12_51_groupi_n_2343 ,csa_tree_add_12_51_groupi_n_726);
  not csa_tree_add_12_51_groupi_drc_bufs19443(csa_tree_add_12_51_groupi_n_2342 ,csa_tree_add_12_51_groupi_n_723);
  not csa_tree_add_12_51_groupi_drc_bufs19444(csa_tree_add_12_51_groupi_n_2341 ,csa_tree_add_12_51_groupi_n_725);
  not csa_tree_add_12_51_groupi_drc_bufs19445(csa_tree_add_12_51_groupi_n_2340 ,csa_tree_add_12_51_groupi_n_724);
  not csa_tree_add_12_51_groupi_drc_bufs19446(csa_tree_add_12_51_groupi_n_2339 ,csa_tree_add_12_51_groupi_n_726);
  not csa_tree_add_12_51_groupi_drc_bufs19447(csa_tree_add_12_51_groupi_n_2338 ,csa_tree_add_12_51_groupi_n_2392);
  not csa_tree_add_12_51_groupi_drc_bufs19453(csa_tree_add_12_51_groupi_n_2337 ,csa_tree_add_12_51_groupi_n_781);
  not csa_tree_add_12_51_groupi_drc_bufs19454(csa_tree_add_12_51_groupi_n_2336 ,csa_tree_add_12_51_groupi_n_783);
  not csa_tree_add_12_51_groupi_drc_bufs19455(csa_tree_add_12_51_groupi_n_2335 ,csa_tree_add_12_51_groupi_n_782);
  not csa_tree_add_12_51_groupi_drc_bufs19456(csa_tree_add_12_51_groupi_n_2334 ,csa_tree_add_12_51_groupi_n_784);
  not csa_tree_add_12_51_groupi_drc_bufs19457(csa_tree_add_12_51_groupi_n_2333 ,csa_tree_add_12_51_groupi_n_781);
  not csa_tree_add_12_51_groupi_drc_bufs19458(csa_tree_add_12_51_groupi_n_2332 ,csa_tree_add_12_51_groupi_n_783);
  not csa_tree_add_12_51_groupi_drc_bufs19459(csa_tree_add_12_51_groupi_n_2331 ,csa_tree_add_12_51_groupi_n_782);
  not csa_tree_add_12_51_groupi_drc_bufs19460(csa_tree_add_12_51_groupi_n_2330 ,csa_tree_add_12_51_groupi_n_784);
  not csa_tree_add_12_51_groupi_drc_bufs19461(csa_tree_add_12_51_groupi_n_2329 ,csa_tree_add_12_51_groupi_n_2395);
  not csa_tree_add_12_51_groupi_drc_bufs19467(csa_tree_add_12_51_groupi_n_2328 ,csa_tree_add_12_51_groupi_n_776);
  not csa_tree_add_12_51_groupi_drc_bufs19468(csa_tree_add_12_51_groupi_n_2327 ,csa_tree_add_12_51_groupi_n_778);
  not csa_tree_add_12_51_groupi_drc_bufs19469(csa_tree_add_12_51_groupi_n_2326 ,csa_tree_add_12_51_groupi_n_777);
  not csa_tree_add_12_51_groupi_drc_bufs19470(csa_tree_add_12_51_groupi_n_2325 ,csa_tree_add_12_51_groupi_n_779);
  not csa_tree_add_12_51_groupi_drc_bufs19471(csa_tree_add_12_51_groupi_n_2324 ,csa_tree_add_12_51_groupi_n_776);
  not csa_tree_add_12_51_groupi_drc_bufs19472(csa_tree_add_12_51_groupi_n_2323 ,csa_tree_add_12_51_groupi_n_778);
  not csa_tree_add_12_51_groupi_drc_bufs19473(csa_tree_add_12_51_groupi_n_2322 ,csa_tree_add_12_51_groupi_n_777);
  not csa_tree_add_12_51_groupi_drc_bufs19474(csa_tree_add_12_51_groupi_n_2321 ,csa_tree_add_12_51_groupi_n_779);
  not csa_tree_add_12_51_groupi_drc_bufs19475(csa_tree_add_12_51_groupi_n_2320 ,csa_tree_add_12_51_groupi_n_2394);
  not csa_tree_add_12_51_groupi_drc_bufs19481(csa_tree_add_12_51_groupi_n_2319 ,csa_tree_add_12_51_groupi_n_771);
  not csa_tree_add_12_51_groupi_drc_bufs19482(csa_tree_add_12_51_groupi_n_2318 ,csa_tree_add_12_51_groupi_n_773);
  not csa_tree_add_12_51_groupi_drc_bufs19483(csa_tree_add_12_51_groupi_n_2317 ,csa_tree_add_12_51_groupi_n_772);
  not csa_tree_add_12_51_groupi_drc_bufs19484(csa_tree_add_12_51_groupi_n_2316 ,csa_tree_add_12_51_groupi_n_774);
  not csa_tree_add_12_51_groupi_drc_bufs19485(csa_tree_add_12_51_groupi_n_2315 ,csa_tree_add_12_51_groupi_n_771);
  not csa_tree_add_12_51_groupi_drc_bufs19486(csa_tree_add_12_51_groupi_n_2314 ,csa_tree_add_12_51_groupi_n_773);
  not csa_tree_add_12_51_groupi_drc_bufs19487(csa_tree_add_12_51_groupi_n_2313 ,csa_tree_add_12_51_groupi_n_772);
  not csa_tree_add_12_51_groupi_drc_bufs19488(csa_tree_add_12_51_groupi_n_2312 ,csa_tree_add_12_51_groupi_n_774);
  not csa_tree_add_12_51_groupi_drc_bufs19489(csa_tree_add_12_51_groupi_n_2311 ,csa_tree_add_12_51_groupi_n_2393);
  not csa_tree_add_12_51_groupi_drc_bufs19495(csa_tree_add_12_51_groupi_n_2310 ,csa_tree_add_12_51_groupi_n_766);
  not csa_tree_add_12_51_groupi_drc_bufs19496(csa_tree_add_12_51_groupi_n_2309 ,csa_tree_add_12_51_groupi_n_768);
  not csa_tree_add_12_51_groupi_drc_bufs19497(csa_tree_add_12_51_groupi_n_2308 ,csa_tree_add_12_51_groupi_n_767);
  not csa_tree_add_12_51_groupi_drc_bufs19498(csa_tree_add_12_51_groupi_n_2307 ,csa_tree_add_12_51_groupi_n_769);
  not csa_tree_add_12_51_groupi_drc_bufs19499(csa_tree_add_12_51_groupi_n_2306 ,csa_tree_add_12_51_groupi_n_766);
  not csa_tree_add_12_51_groupi_drc_bufs19500(csa_tree_add_12_51_groupi_n_2305 ,csa_tree_add_12_51_groupi_n_768);
  not csa_tree_add_12_51_groupi_drc_bufs19501(csa_tree_add_12_51_groupi_n_2304 ,csa_tree_add_12_51_groupi_n_767);
  not csa_tree_add_12_51_groupi_drc_bufs19502(csa_tree_add_12_51_groupi_n_2303 ,csa_tree_add_12_51_groupi_n_769);
  not csa_tree_add_12_51_groupi_drc_bufs19503(csa_tree_add_12_51_groupi_n_2302 ,csa_tree_add_12_51_groupi_n_2391);
  not csa_tree_add_12_51_groupi_drc_bufs19509(csa_tree_add_12_51_groupi_n_2301 ,csa_tree_add_12_51_groupi_n_761);
  not csa_tree_add_12_51_groupi_drc_bufs19510(csa_tree_add_12_51_groupi_n_2300 ,csa_tree_add_12_51_groupi_n_763);
  not csa_tree_add_12_51_groupi_drc_bufs19511(csa_tree_add_12_51_groupi_n_2299 ,csa_tree_add_12_51_groupi_n_762);
  not csa_tree_add_12_51_groupi_drc_bufs19512(csa_tree_add_12_51_groupi_n_2298 ,csa_tree_add_12_51_groupi_n_764);
  not csa_tree_add_12_51_groupi_drc_bufs19513(csa_tree_add_12_51_groupi_n_2297 ,csa_tree_add_12_51_groupi_n_761);
  not csa_tree_add_12_51_groupi_drc_bufs19514(csa_tree_add_12_51_groupi_n_2296 ,csa_tree_add_12_51_groupi_n_763);
  not csa_tree_add_12_51_groupi_drc_bufs19515(csa_tree_add_12_51_groupi_n_2295 ,csa_tree_add_12_51_groupi_n_762);
  not csa_tree_add_12_51_groupi_drc_bufs19516(csa_tree_add_12_51_groupi_n_2294 ,csa_tree_add_12_51_groupi_n_764);
  not csa_tree_add_12_51_groupi_drc_bufs19517(csa_tree_add_12_51_groupi_n_2293 ,csa_tree_add_12_51_groupi_n_2390);
  not csa_tree_add_12_51_groupi_drc_bufs19523(csa_tree_add_12_51_groupi_n_2292 ,csa_tree_add_12_51_groupi_n_758);
  not csa_tree_add_12_51_groupi_drc_bufs19524(csa_tree_add_12_51_groupi_n_2291 ,csa_tree_add_12_51_groupi_n_714);
  not csa_tree_add_12_51_groupi_drc_bufs19525(csa_tree_add_12_51_groupi_n_2290 ,csa_tree_add_12_51_groupi_n_759);
  not csa_tree_add_12_51_groupi_drc_bufs19526(csa_tree_add_12_51_groupi_n_2289 ,csa_tree_add_12_51_groupi_n_715);
  not csa_tree_add_12_51_groupi_drc_bufs19527(csa_tree_add_12_51_groupi_n_2288 ,csa_tree_add_12_51_groupi_n_758);
  not csa_tree_add_12_51_groupi_drc_bufs19528(csa_tree_add_12_51_groupi_n_2287 ,csa_tree_add_12_51_groupi_n_714);
  not csa_tree_add_12_51_groupi_drc_bufs19529(csa_tree_add_12_51_groupi_n_2286 ,csa_tree_add_12_51_groupi_n_759);
  not csa_tree_add_12_51_groupi_drc_bufs19530(csa_tree_add_12_51_groupi_n_2285 ,csa_tree_add_12_51_groupi_n_715);
  not csa_tree_add_12_51_groupi_drc_bufs19531(csa_tree_add_12_51_groupi_n_2284 ,csa_tree_add_12_51_groupi_n_2389);
  not csa_tree_add_12_51_groupi_drc_bufs19537(csa_tree_add_12_51_groupi_n_2283 ,csa_tree_add_12_51_groupi_n_720);
  not csa_tree_add_12_51_groupi_drc_bufs19538(csa_tree_add_12_51_groupi_n_2282 ,csa_tree_add_12_51_groupi_n_787);
  not csa_tree_add_12_51_groupi_drc_bufs19539(csa_tree_add_12_51_groupi_n_2281 ,csa_tree_add_12_51_groupi_n_721);
  not csa_tree_add_12_51_groupi_drc_bufs19540(csa_tree_add_12_51_groupi_n_2280 ,csa_tree_add_12_51_groupi_n_788);
  not csa_tree_add_12_51_groupi_drc_bufs19541(csa_tree_add_12_51_groupi_n_2279 ,csa_tree_add_12_51_groupi_n_720);
  not csa_tree_add_12_51_groupi_drc_bufs19542(csa_tree_add_12_51_groupi_n_2278 ,csa_tree_add_12_51_groupi_n_787);
  not csa_tree_add_12_51_groupi_drc_bufs19543(csa_tree_add_12_51_groupi_n_2277 ,csa_tree_add_12_51_groupi_n_721);
  not csa_tree_add_12_51_groupi_drc_bufs19544(csa_tree_add_12_51_groupi_n_2276 ,csa_tree_add_12_51_groupi_n_788);
  not csa_tree_add_12_51_groupi_drc_bufs19545(csa_tree_add_12_51_groupi_n_2275 ,csa_tree_add_12_51_groupi_n_2388);
  not csa_tree_add_12_51_groupi_drc_bufs19551(csa_tree_add_12_51_groupi_n_2274 ,csa_tree_add_12_51_groupi_n_754);
  not csa_tree_add_12_51_groupi_drc_bufs19552(csa_tree_add_12_51_groupi_n_2273 ,csa_tree_add_12_51_groupi_n_756);
  not csa_tree_add_12_51_groupi_drc_bufs19553(csa_tree_add_12_51_groupi_n_2272 ,csa_tree_add_12_51_groupi_n_755);
  not csa_tree_add_12_51_groupi_drc_bufs19554(csa_tree_add_12_51_groupi_n_2271 ,csa_tree_add_12_51_groupi_n_757);
  not csa_tree_add_12_51_groupi_drc_bufs19555(csa_tree_add_12_51_groupi_n_2270 ,csa_tree_add_12_51_groupi_n_754);
  not csa_tree_add_12_51_groupi_drc_bufs19556(csa_tree_add_12_51_groupi_n_2269 ,csa_tree_add_12_51_groupi_n_756);
  not csa_tree_add_12_51_groupi_drc_bufs19557(csa_tree_add_12_51_groupi_n_2268 ,csa_tree_add_12_51_groupi_n_755);
  not csa_tree_add_12_51_groupi_drc_bufs19558(csa_tree_add_12_51_groupi_n_2267 ,csa_tree_add_12_51_groupi_n_757);
  not csa_tree_add_12_51_groupi_drc_bufs19559(csa_tree_add_12_51_groupi_n_2266 ,csa_tree_add_12_51_groupi_n_2387);
  not csa_tree_add_12_51_groupi_drc_bufs19565(csa_tree_add_12_51_groupi_n_2265 ,csa_tree_add_12_51_groupi_n_751);
  not csa_tree_add_12_51_groupi_drc_bufs19566(csa_tree_add_12_51_groupi_n_2264 ,csa_tree_add_12_51_groupi_n_717);
  not csa_tree_add_12_51_groupi_drc_bufs19567(csa_tree_add_12_51_groupi_n_2263 ,csa_tree_add_12_51_groupi_n_752);
  not csa_tree_add_12_51_groupi_drc_bufs19568(csa_tree_add_12_51_groupi_n_2262 ,csa_tree_add_12_51_groupi_n_718);
  not csa_tree_add_12_51_groupi_drc_bufs19569(csa_tree_add_12_51_groupi_n_2261 ,csa_tree_add_12_51_groupi_n_751);
  not csa_tree_add_12_51_groupi_drc_bufs19570(csa_tree_add_12_51_groupi_n_2260 ,csa_tree_add_12_51_groupi_n_717);
  not csa_tree_add_12_51_groupi_drc_bufs19571(csa_tree_add_12_51_groupi_n_2259 ,csa_tree_add_12_51_groupi_n_752);
  not csa_tree_add_12_51_groupi_drc_bufs19572(csa_tree_add_12_51_groupi_n_2258 ,csa_tree_add_12_51_groupi_n_718);
  not csa_tree_add_12_51_groupi_drc_bufs19573(csa_tree_add_12_51_groupi_n_2257 ,csa_tree_add_12_51_groupi_n_2359);
  not csa_tree_add_12_51_groupi_drc_bufs19579(csa_tree_add_12_51_groupi_n_2256 ,csa_tree_add_12_51_groupi_n_747);
  not csa_tree_add_12_51_groupi_drc_bufs19580(csa_tree_add_12_51_groupi_n_2255 ,csa_tree_add_12_51_groupi_n_749);
  not csa_tree_add_12_51_groupi_drc_bufs19581(csa_tree_add_12_51_groupi_n_2254 ,csa_tree_add_12_51_groupi_n_748);
  not csa_tree_add_12_51_groupi_drc_bufs19582(csa_tree_add_12_51_groupi_n_2253 ,csa_tree_add_12_51_groupi_n_750);
  not csa_tree_add_12_51_groupi_drc_bufs19583(csa_tree_add_12_51_groupi_n_2252 ,csa_tree_add_12_51_groupi_n_747);
  not csa_tree_add_12_51_groupi_drc_bufs19584(csa_tree_add_12_51_groupi_n_2251 ,csa_tree_add_12_51_groupi_n_749);
  not csa_tree_add_12_51_groupi_drc_bufs19585(csa_tree_add_12_51_groupi_n_2250 ,csa_tree_add_12_51_groupi_n_748);
  not csa_tree_add_12_51_groupi_drc_bufs19586(csa_tree_add_12_51_groupi_n_2249 ,csa_tree_add_12_51_groupi_n_750);
  not csa_tree_add_12_51_groupi_drc_bufs19587(csa_tree_add_12_51_groupi_n_2248 ,csa_tree_add_12_51_groupi_n_2358);
  not csa_tree_add_12_51_groupi_drc_bufs19593(csa_tree_add_12_51_groupi_n_2247 ,csa_tree_add_12_51_groupi_n_744);
  not csa_tree_add_12_51_groupi_drc_bufs19594(csa_tree_add_12_51_groupi_n_2246 ,csa_tree_add_12_51_groupi_n_791);
  not csa_tree_add_12_51_groupi_drc_bufs19595(csa_tree_add_12_51_groupi_n_2245 ,csa_tree_add_12_51_groupi_n_745);
  not csa_tree_add_12_51_groupi_drc_bufs19596(csa_tree_add_12_51_groupi_n_2244 ,csa_tree_add_12_51_groupi_n_792);
  not csa_tree_add_12_51_groupi_drc_bufs19597(csa_tree_add_12_51_groupi_n_2243 ,csa_tree_add_12_51_groupi_n_744);
  not csa_tree_add_12_51_groupi_drc_bufs19598(csa_tree_add_12_51_groupi_n_2242 ,csa_tree_add_12_51_groupi_n_791);
  not csa_tree_add_12_51_groupi_drc_bufs19599(csa_tree_add_12_51_groupi_n_2241 ,csa_tree_add_12_51_groupi_n_745);
  not csa_tree_add_12_51_groupi_drc_bufs19600(csa_tree_add_12_51_groupi_n_2240 ,csa_tree_add_12_51_groupi_n_792);
  not csa_tree_add_12_51_groupi_drc_bufs19601(csa_tree_add_12_51_groupi_n_2239 ,csa_tree_add_12_51_groupi_n_2357);
  not csa_tree_add_12_51_groupi_drc_bufs19607(csa_tree_add_12_51_groupi_n_2238 ,csa_tree_add_12_51_groupi_n_739);
  not csa_tree_add_12_51_groupi_drc_bufs19608(csa_tree_add_12_51_groupi_n_2237 ,csa_tree_add_12_51_groupi_n_741);
  not csa_tree_add_12_51_groupi_drc_bufs19609(csa_tree_add_12_51_groupi_n_2236 ,csa_tree_add_12_51_groupi_n_740);
  not csa_tree_add_12_51_groupi_drc_bufs19610(csa_tree_add_12_51_groupi_n_2235 ,csa_tree_add_12_51_groupi_n_742);
  not csa_tree_add_12_51_groupi_drc_bufs19611(csa_tree_add_12_51_groupi_n_2234 ,csa_tree_add_12_51_groupi_n_739);
  not csa_tree_add_12_51_groupi_drc_bufs19612(csa_tree_add_12_51_groupi_n_2233 ,csa_tree_add_12_51_groupi_n_741);
  not csa_tree_add_12_51_groupi_drc_bufs19613(csa_tree_add_12_51_groupi_n_2232 ,csa_tree_add_12_51_groupi_n_740);
  not csa_tree_add_12_51_groupi_drc_bufs19614(csa_tree_add_12_51_groupi_n_2231 ,csa_tree_add_12_51_groupi_n_742);
  not csa_tree_add_12_51_groupi_drc_bufs19615(csa_tree_add_12_51_groupi_n_2230 ,csa_tree_add_12_51_groupi_n_2356);
  not csa_tree_add_12_51_groupi_drc_bufs19621(csa_tree_add_12_51_groupi_n_2229 ,csa_tree_add_12_51_groupi_n_736);
  not csa_tree_add_12_51_groupi_drc_bufs19622(csa_tree_add_12_51_groupi_n_2228 ,csa_tree_add_12_51_groupi_n_789);
  not csa_tree_add_12_51_groupi_drc_bufs19623(csa_tree_add_12_51_groupi_n_2227 ,csa_tree_add_12_51_groupi_n_737);
  not csa_tree_add_12_51_groupi_drc_bufs19624(csa_tree_add_12_51_groupi_n_2226 ,csa_tree_add_12_51_groupi_n_790);
  not csa_tree_add_12_51_groupi_drc_bufs19625(csa_tree_add_12_51_groupi_n_2225 ,csa_tree_add_12_51_groupi_n_736);
  not csa_tree_add_12_51_groupi_drc_bufs19626(csa_tree_add_12_51_groupi_n_2224 ,csa_tree_add_12_51_groupi_n_789);
  not csa_tree_add_12_51_groupi_drc_bufs19627(csa_tree_add_12_51_groupi_n_2223 ,csa_tree_add_12_51_groupi_n_737);
  not csa_tree_add_12_51_groupi_drc_bufs19628(csa_tree_add_12_51_groupi_n_2222 ,csa_tree_add_12_51_groupi_n_790);
  not csa_tree_add_12_51_groupi_drc_bufs19629(csa_tree_add_12_51_groupi_n_2221 ,csa_tree_add_12_51_groupi_n_2355);
  not csa_tree_add_12_51_groupi_drc_bufs19635(csa_tree_add_12_51_groupi_n_2220 ,csa_tree_add_12_51_groupi_n_731);
  not csa_tree_add_12_51_groupi_drc_bufs19636(csa_tree_add_12_51_groupi_n_2219 ,csa_tree_add_12_51_groupi_n_733);
  not csa_tree_add_12_51_groupi_drc_bufs19637(csa_tree_add_12_51_groupi_n_2218 ,csa_tree_add_12_51_groupi_n_732);
  not csa_tree_add_12_51_groupi_drc_bufs19638(csa_tree_add_12_51_groupi_n_2217 ,csa_tree_add_12_51_groupi_n_734);
  not csa_tree_add_12_51_groupi_drc_bufs19639(csa_tree_add_12_51_groupi_n_2216 ,csa_tree_add_12_51_groupi_n_731);
  not csa_tree_add_12_51_groupi_drc_bufs19640(csa_tree_add_12_51_groupi_n_2215 ,csa_tree_add_12_51_groupi_n_733);
  not csa_tree_add_12_51_groupi_drc_bufs19641(csa_tree_add_12_51_groupi_n_2214 ,csa_tree_add_12_51_groupi_n_732);
  not csa_tree_add_12_51_groupi_drc_bufs19642(csa_tree_add_12_51_groupi_n_2213 ,csa_tree_add_12_51_groupi_n_734);
  not csa_tree_add_12_51_groupi_drc_bufs19643(csa_tree_add_12_51_groupi_n_2212 ,csa_tree_add_12_51_groupi_n_2396);
  not csa_tree_add_12_51_groupi_drc_bufs19649(csa_tree_add_12_51_groupi_n_2211 ,csa_tree_add_12_51_groupi_n_728);
  not csa_tree_add_12_51_groupi_drc_bufs19650(csa_tree_add_12_51_groupi_n_2210 ,csa_tree_add_12_51_groupi_n_785);
  not csa_tree_add_12_51_groupi_drc_bufs19651(csa_tree_add_12_51_groupi_n_2209 ,csa_tree_add_12_51_groupi_n_729);
  not csa_tree_add_12_51_groupi_drc_bufs19652(csa_tree_add_12_51_groupi_n_2208 ,csa_tree_add_12_51_groupi_n_786);
  not csa_tree_add_12_51_groupi_drc_bufs19653(csa_tree_add_12_51_groupi_n_2207 ,csa_tree_add_12_51_groupi_n_728);
  not csa_tree_add_12_51_groupi_drc_bufs19654(csa_tree_add_12_51_groupi_n_2206 ,csa_tree_add_12_51_groupi_n_785);
  not csa_tree_add_12_51_groupi_drc_bufs19655(csa_tree_add_12_51_groupi_n_2205 ,csa_tree_add_12_51_groupi_n_729);
  not csa_tree_add_12_51_groupi_drc_bufs19656(csa_tree_add_12_51_groupi_n_2204 ,csa_tree_add_12_51_groupi_n_786);
  not csa_tree_add_12_51_groupi_drc_bufs19657(csa_tree_add_12_51_groupi_n_2203 ,csa_tree_add_12_51_groupi_n_2360);
  not csa_tree_add_12_51_groupi_drc_bufs21080(csa_tree_add_12_51_groupi_n_2202 ,csa_tree_add_12_51_groupi_n_2200);
  not csa_tree_add_12_51_groupi_drc_bufs21081(csa_tree_add_12_51_groupi_n_2201 ,csa_tree_add_12_51_groupi_n_2200);
  not csa_tree_add_12_51_groupi_drc_bufs21082(csa_tree_add_12_51_groupi_n_2200 ,csa_tree_add_12_51_groupi_n_2348);
  not csa_tree_add_12_51_groupi_drc_bufs21084(csa_tree_add_12_51_groupi_n_2199 ,csa_tree_add_12_51_groupi_n_2197);
  not csa_tree_add_12_51_groupi_drc_bufs21085(csa_tree_add_12_51_groupi_n_2198 ,csa_tree_add_12_51_groupi_n_2197);
  not csa_tree_add_12_51_groupi_drc_bufs21086(csa_tree_add_12_51_groupi_n_2197 ,csa_tree_add_12_51_groupi_n_2465);
  not csa_tree_add_12_51_groupi_drc_bufs21088(csa_tree_add_12_51_groupi_n_2196 ,csa_tree_add_12_51_groupi_n_2194);
  not csa_tree_add_12_51_groupi_drc_bufs21089(csa_tree_add_12_51_groupi_n_2195 ,csa_tree_add_12_51_groupi_n_2194);
  not csa_tree_add_12_51_groupi_drc_bufs21090(csa_tree_add_12_51_groupi_n_2194 ,csa_tree_add_12_51_groupi_n_2464);
  not csa_tree_add_12_51_groupi_drc_bufs21092(csa_tree_add_12_51_groupi_n_2193 ,csa_tree_add_12_51_groupi_n_2191);
  not csa_tree_add_12_51_groupi_drc_bufs21093(csa_tree_add_12_51_groupi_n_2192 ,csa_tree_add_12_51_groupi_n_2191);
  not csa_tree_add_12_51_groupi_drc_bufs21094(csa_tree_add_12_51_groupi_n_2191 ,csa_tree_add_12_51_groupi_n_2639);
  not csa_tree_add_12_51_groupi_drc_bufs21096(csa_tree_add_12_51_groupi_n_2190 ,csa_tree_add_12_51_groupi_n_2188);
  not csa_tree_add_12_51_groupi_drc_bufs21097(csa_tree_add_12_51_groupi_n_2189 ,csa_tree_add_12_51_groupi_n_2188);
  not csa_tree_add_12_51_groupi_drc_bufs21098(csa_tree_add_12_51_groupi_n_2188 ,csa_tree_add_12_51_groupi_n_2640);
  not csa_tree_add_12_51_groupi_drc_bufs21100(csa_tree_add_12_51_groupi_n_2187 ,csa_tree_add_12_51_groupi_n_2185);
  not csa_tree_add_12_51_groupi_drc_bufs21101(csa_tree_add_12_51_groupi_n_2186 ,csa_tree_add_12_51_groupi_n_2185);
  not csa_tree_add_12_51_groupi_drc_bufs21102(csa_tree_add_12_51_groupi_n_2185 ,csa_tree_add_12_51_groupi_n_2350);
  not csa_tree_add_12_51_groupi_drc_bufs21104(csa_tree_add_12_51_groupi_n_2184 ,csa_tree_add_12_51_groupi_n_2182);
  not csa_tree_add_12_51_groupi_drc_bufs21105(csa_tree_add_12_51_groupi_n_2183 ,csa_tree_add_12_51_groupi_n_2182);
  not csa_tree_add_12_51_groupi_drc_bufs21106(csa_tree_add_12_51_groupi_n_2182 ,csa_tree_add_12_51_groupi_n_2353);
  not csa_tree_add_12_51_groupi_drc_bufs21108(csa_tree_add_12_51_groupi_n_2181 ,csa_tree_add_12_51_groupi_n_2179);
  not csa_tree_add_12_51_groupi_drc_bufs21109(csa_tree_add_12_51_groupi_n_2180 ,csa_tree_add_12_51_groupi_n_2179);
  not csa_tree_add_12_51_groupi_drc_bufs21110(csa_tree_add_12_51_groupi_n_2179 ,csa_tree_add_12_51_groupi_n_6161);
  not csa_tree_add_12_51_groupi_drc_bufs21112(csa_tree_add_12_51_groupi_n_2178 ,csa_tree_add_12_51_groupi_n_2176);
  not csa_tree_add_12_51_groupi_drc_bufs21113(csa_tree_add_12_51_groupi_n_2177 ,csa_tree_add_12_51_groupi_n_2176);
  not csa_tree_add_12_51_groupi_drc_bufs21114(csa_tree_add_12_51_groupi_n_2176 ,csa_tree_add_12_51_groupi_n_6162);
  not csa_tree_add_12_51_groupi_drc_bufs21116(csa_tree_add_12_51_groupi_n_2175 ,csa_tree_add_12_51_groupi_n_2173);
  not csa_tree_add_12_51_groupi_drc_bufs21117(csa_tree_add_12_51_groupi_n_2174 ,csa_tree_add_12_51_groupi_n_2173);
  not csa_tree_add_12_51_groupi_drc_bufs21118(csa_tree_add_12_51_groupi_n_2173 ,csa_tree_add_12_51_groupi_n_2461);
  not csa_tree_add_12_51_groupi_drc_bufs21120(csa_tree_add_12_51_groupi_n_2172 ,csa_tree_add_12_51_groupi_n_2170);
  not csa_tree_add_12_51_groupi_drc_bufs21121(csa_tree_add_12_51_groupi_n_2171 ,csa_tree_add_12_51_groupi_n_2170);
  not csa_tree_add_12_51_groupi_drc_bufs21122(csa_tree_add_12_51_groupi_n_2170 ,csa_tree_add_12_51_groupi_n_2347);
  not csa_tree_add_12_51_groupi_drc_bufs21124(csa_tree_add_12_51_groupi_n_2169 ,csa_tree_add_12_51_groupi_n_2167);
  not csa_tree_add_12_51_groupi_drc_bufs21125(csa_tree_add_12_51_groupi_n_2168 ,csa_tree_add_12_51_groupi_n_2167);
  not csa_tree_add_12_51_groupi_drc_bufs21126(csa_tree_add_12_51_groupi_n_2167 ,csa_tree_add_12_51_groupi_n_2462);
  not csa_tree_add_12_51_groupi_drc_bufs21128(csa_tree_add_12_51_groupi_n_2166 ,csa_tree_add_12_51_groupi_n_2164);
  not csa_tree_add_12_51_groupi_drc_bufs21129(csa_tree_add_12_51_groupi_n_2165 ,csa_tree_add_12_51_groupi_n_2164);
  not csa_tree_add_12_51_groupi_drc_bufs21130(csa_tree_add_12_51_groupi_n_2164 ,csa_tree_add_12_51_groupi_n_2461);
  not csa_tree_add_12_51_groupi_drc_bufs21133(csa_tree_add_12_51_groupi_n_2163 ,csa_tree_add_12_51_groupi_n_2162);
  not csa_tree_add_12_51_groupi_drc_bufs21134(csa_tree_add_12_51_groupi_n_2162 ,csa_tree_add_12_51_groupi_n_3510);
  not csa_tree_add_12_51_groupi_drc_bufs21137(csa_tree_add_12_51_groupi_n_2161 ,csa_tree_add_12_51_groupi_n_2351);
  not csa_tree_add_12_51_groupi_drc_bufs21138(csa_tree_add_12_51_groupi_n_2351 ,csa_tree_add_12_51_groupi_n_2949);
  not csa_tree_add_12_51_groupi_drc_bufs21140(csa_tree_add_12_51_groupi_n_2160 ,csa_tree_add_12_51_groupi_n_2158);
  not csa_tree_add_12_51_groupi_drc_bufs21141(csa_tree_add_12_51_groupi_n_2159 ,csa_tree_add_12_51_groupi_n_2158);
  not csa_tree_add_12_51_groupi_drc_bufs21142(csa_tree_add_12_51_groupi_n_2158 ,csa_tree_add_12_51_groupi_n_2349);
  not csa_tree_add_12_51_groupi_drc_bufs21159(csa_tree_add_12_51_groupi_n_2157 ,csa_tree_add_12_51_groupi_n_2156);
  not csa_tree_add_12_51_groupi_drc_bufs21161(csa_tree_add_12_51_groupi_n_2156 ,csa_tree_add_12_51_groupi_n_2642);
  not csa_tree_add_12_51_groupi_drc_bufs21163(csa_tree_add_12_51_groupi_n_2155 ,csa_tree_add_12_51_groupi_n_2154);
  not csa_tree_add_12_51_groupi_drc_bufs21165(csa_tree_add_12_51_groupi_n_2154 ,csa_tree_add_12_51_groupi_n_6164);
  not csa_tree_add_12_51_groupi_drc_bufs21393(csa_tree_add_12_51_groupi_n_2153 ,csa_tree_add_12_51_groupi_n_2152);
  not csa_tree_add_12_51_groupi_drc_bufs21394(csa_tree_add_12_51_groupi_n_2152 ,csa_tree_add_12_51_groupi_n_3509);
  not csa_tree_add_12_51_groupi_drc_bufs21415(csa_tree_add_12_51_groupi_n_2151 ,csa_tree_add_12_51_groupi_n_2354);
  not csa_tree_add_12_51_groupi_drc_bufs21416(csa_tree_add_12_51_groupi_n_2354 ,csa_tree_add_12_51_groupi_n_6937);
  not csa_tree_add_12_51_groupi_drc_bufs21419(csa_tree_add_12_51_groupi_n_2150 ,csa_tree_add_12_51_groupi_n_2352);
  not csa_tree_add_12_51_groupi_drc_bufs21420(csa_tree_add_12_51_groupi_n_2352 ,csa_tree_add_12_51_groupi_n_4129);
  not csa_tree_add_12_51_groupi_drc_bufs21497(csa_tree_add_12_51_groupi_n_2149 ,csa_tree_add_12_51_groupi_n_2147);
  not csa_tree_add_12_51_groupi_drc_bufs21498(csa_tree_add_12_51_groupi_n_2148 ,csa_tree_add_12_51_groupi_n_2147);
  not csa_tree_add_12_51_groupi_drc_bufs21499(csa_tree_add_12_51_groupi_n_2147 ,csa_tree_add_12_51_groupi_n_2921);
  not csa_tree_add_12_51_groupi_drc_bufs21502(csa_tree_add_12_51_groupi_n_2146 ,csa_tree_add_12_51_groupi_n_2144);
  not csa_tree_add_12_51_groupi_drc_bufs21503(csa_tree_add_12_51_groupi_n_2145 ,csa_tree_add_12_51_groupi_n_2144);
  not csa_tree_add_12_51_groupi_drc_bufs21504(csa_tree_add_12_51_groupi_n_2144 ,csa_tree_add_12_51_groupi_n_2920);
  not csa_tree_add_12_51_groupi_drc_bufs21507(csa_tree_add_12_51_groupi_n_2143 ,csa_tree_add_12_51_groupi_n_2141);
  not csa_tree_add_12_51_groupi_drc_bufs21508(csa_tree_add_12_51_groupi_n_2142 ,csa_tree_add_12_51_groupi_n_2141);
  not csa_tree_add_12_51_groupi_drc_bufs21509(csa_tree_add_12_51_groupi_n_2141 ,csa_tree_add_12_51_groupi_n_2919);
  not csa_tree_add_12_51_groupi_drc_bufs21512(csa_tree_add_12_51_groupi_n_2140 ,csa_tree_add_12_51_groupi_n_2138);
  not csa_tree_add_12_51_groupi_drc_bufs21513(csa_tree_add_12_51_groupi_n_2139 ,csa_tree_add_12_51_groupi_n_2138);
  not csa_tree_add_12_51_groupi_drc_bufs21514(csa_tree_add_12_51_groupi_n_2138 ,csa_tree_add_12_51_groupi_n_2918);
  not csa_tree_add_12_51_groupi_drc_bufs21517(csa_tree_add_12_51_groupi_n_2137 ,csa_tree_add_12_51_groupi_n_2135);
  not csa_tree_add_12_51_groupi_drc_bufs21518(csa_tree_add_12_51_groupi_n_2136 ,csa_tree_add_12_51_groupi_n_2135);
  not csa_tree_add_12_51_groupi_drc_bufs21519(csa_tree_add_12_51_groupi_n_2135 ,csa_tree_add_12_51_groupi_n_2917);
  not csa_tree_add_12_51_groupi_drc_bufs21522(csa_tree_add_12_51_groupi_n_2134 ,csa_tree_add_12_51_groupi_n_2132);
  not csa_tree_add_12_51_groupi_drc_bufs21523(csa_tree_add_12_51_groupi_n_2133 ,csa_tree_add_12_51_groupi_n_2132);
  not csa_tree_add_12_51_groupi_drc_bufs21524(csa_tree_add_12_51_groupi_n_2132 ,csa_tree_add_12_51_groupi_n_2916);
  not csa_tree_add_12_51_groupi_drc_bufs21527(csa_tree_add_12_51_groupi_n_2131 ,csa_tree_add_12_51_groupi_n_2129);
  not csa_tree_add_12_51_groupi_drc_bufs21528(csa_tree_add_12_51_groupi_n_2130 ,csa_tree_add_12_51_groupi_n_2129);
  not csa_tree_add_12_51_groupi_drc_bufs21529(csa_tree_add_12_51_groupi_n_2129 ,csa_tree_add_12_51_groupi_n_2915);
  not csa_tree_add_12_51_groupi_drc_bufs21532(csa_tree_add_12_51_groupi_n_2128 ,csa_tree_add_12_51_groupi_n_2126);
  not csa_tree_add_12_51_groupi_drc_bufs21533(csa_tree_add_12_51_groupi_n_2127 ,csa_tree_add_12_51_groupi_n_2126);
  not csa_tree_add_12_51_groupi_drc_bufs21534(csa_tree_add_12_51_groupi_n_2126 ,csa_tree_add_12_51_groupi_n_2914);
  not csa_tree_add_12_51_groupi_drc_bufs21537(csa_tree_add_12_51_groupi_n_2125 ,csa_tree_add_12_51_groupi_n_2123);
  not csa_tree_add_12_51_groupi_drc_bufs21538(csa_tree_add_12_51_groupi_n_2124 ,csa_tree_add_12_51_groupi_n_2123);
  not csa_tree_add_12_51_groupi_drc_bufs21539(csa_tree_add_12_51_groupi_n_2123 ,csa_tree_add_12_51_groupi_n_2913);
  not csa_tree_add_12_51_groupi_drc_bufs21542(csa_tree_add_12_51_groupi_n_2122 ,csa_tree_add_12_51_groupi_n_2120);
  not csa_tree_add_12_51_groupi_drc_bufs21543(csa_tree_add_12_51_groupi_n_2121 ,csa_tree_add_12_51_groupi_n_2120);
  not csa_tree_add_12_51_groupi_drc_bufs21544(csa_tree_add_12_51_groupi_n_2120 ,csa_tree_add_12_51_groupi_n_2912);
  not csa_tree_add_12_51_groupi_drc_bufs21547(csa_tree_add_12_51_groupi_n_2119 ,csa_tree_add_12_51_groupi_n_2117);
  not csa_tree_add_12_51_groupi_drc_bufs21548(csa_tree_add_12_51_groupi_n_2118 ,csa_tree_add_12_51_groupi_n_2117);
  not csa_tree_add_12_51_groupi_drc_bufs21549(csa_tree_add_12_51_groupi_n_2117 ,csa_tree_add_12_51_groupi_n_2911);
  not csa_tree_add_12_51_groupi_drc_bufs21552(csa_tree_add_12_51_groupi_n_2116 ,csa_tree_add_12_51_groupi_n_2114);
  not csa_tree_add_12_51_groupi_drc_bufs21553(csa_tree_add_12_51_groupi_n_2115 ,csa_tree_add_12_51_groupi_n_2114);
  not csa_tree_add_12_51_groupi_drc_bufs21554(csa_tree_add_12_51_groupi_n_2114 ,csa_tree_add_12_51_groupi_n_2909);
  not csa_tree_add_12_51_groupi_drc_bufs21557(csa_tree_add_12_51_groupi_n_2113 ,csa_tree_add_12_51_groupi_n_2111);
  not csa_tree_add_12_51_groupi_drc_bufs21558(csa_tree_add_12_51_groupi_n_2112 ,csa_tree_add_12_51_groupi_n_2111);
  not csa_tree_add_12_51_groupi_drc_bufs21559(csa_tree_add_12_51_groupi_n_2111 ,csa_tree_add_12_51_groupi_n_2910);
  not csa_tree_add_12_51_groupi_drc_bufs21562(csa_tree_add_12_51_groupi_n_2110 ,csa_tree_add_12_51_groupi_n_2108);
  not csa_tree_add_12_51_groupi_drc_bufs21563(csa_tree_add_12_51_groupi_n_2109 ,csa_tree_add_12_51_groupi_n_2108);
  not csa_tree_add_12_51_groupi_drc_bufs21564(csa_tree_add_12_51_groupi_n_2108 ,csa_tree_add_12_51_groupi_n_2908);
  not csa_tree_add_12_51_groupi_drc_bufs21567(csa_tree_add_12_51_groupi_n_2107 ,csa_tree_add_12_51_groupi_n_2105);
  not csa_tree_add_12_51_groupi_drc_bufs21568(csa_tree_add_12_51_groupi_n_2106 ,csa_tree_add_12_51_groupi_n_2105);
  not csa_tree_add_12_51_groupi_drc_bufs21569(csa_tree_add_12_51_groupi_n_2105 ,csa_tree_add_12_51_groupi_n_2907);
  not csa_tree_add_12_51_groupi_drc_bufs21622(csa_tree_add_12_51_groupi_n_2104 ,csa_tree_add_12_51_groupi_n_2103);
  not csa_tree_add_12_51_groupi_drc_bufs21624(csa_tree_add_12_51_groupi_n_2103 ,csa_tree_add_12_51_groupi_n_2936);
  not csa_tree_add_12_51_groupi_drc_bufs21667(csa_tree_add_12_51_groupi_n_2102 ,csa_tree_add_12_51_groupi_n_2101);
  not csa_tree_add_12_51_groupi_drc_bufs21669(csa_tree_add_12_51_groupi_n_2101 ,csa_tree_add_12_51_groupi_n_2504);
  not csa_tree_add_12_51_groupi_drc_bufs21672(csa_tree_add_12_51_groupi_n_2100 ,csa_tree_add_12_51_groupi_n_2099);
  not csa_tree_add_12_51_groupi_drc_bufs21674(csa_tree_add_12_51_groupi_n_2099 ,csa_tree_add_12_51_groupi_n_2923);
  not csa_tree_add_12_51_groupi_drc_bufs21677(csa_tree_add_12_51_groupi_n_2098 ,csa_tree_add_12_51_groupi_n_2097);
  not csa_tree_add_12_51_groupi_drc_bufs21679(csa_tree_add_12_51_groupi_n_2097 ,csa_tree_add_12_51_groupi_n_2926);
  not csa_tree_add_12_51_groupi_drc_bufs21697(csa_tree_add_12_51_groupi_n_2096 ,csa_tree_add_12_51_groupi_n_2095);
  not csa_tree_add_12_51_groupi_drc_bufs21699(csa_tree_add_12_51_groupi_n_2095 ,csa_tree_add_12_51_groupi_n_2463);
  not csa_tree_add_12_51_groupi_drc_bufs21702(csa_tree_add_12_51_groupi_n_2094 ,csa_tree_add_12_51_groupi_n_2093);
  not csa_tree_add_12_51_groupi_drc_bufs21704(csa_tree_add_12_51_groupi_n_2093 ,csa_tree_add_12_51_groupi_n_2754);
  not csa_tree_add_12_51_groupi_drc_bufs21712(csa_tree_add_12_51_groupi_n_2092 ,csa_tree_add_12_51_groupi_n_2091);
  not csa_tree_add_12_51_groupi_drc_bufs21714(csa_tree_add_12_51_groupi_n_2091 ,csa_tree_add_12_51_groupi_n_2948);
  not csa_tree_add_12_51_groupi_drc_bufs21732(csa_tree_add_12_51_groupi_n_2090 ,csa_tree_add_12_51_groupi_n_2089);
  not csa_tree_add_12_51_groupi_drc_bufs21734(csa_tree_add_12_51_groupi_n_2089 ,csa_tree_add_12_51_groupi_n_2927);
  not csa_tree_add_12_51_groupi_drc_bufs21747(csa_tree_add_12_51_groupi_n_2088 ,csa_tree_add_12_51_groupi_n_2087);
  not csa_tree_add_12_51_groupi_drc_bufs21749(csa_tree_add_12_51_groupi_n_2087 ,csa_tree_add_12_51_groupi_n_2925);
  not csa_tree_add_12_51_groupi_drc_bufs21767(csa_tree_add_12_51_groupi_n_2086 ,csa_tree_add_12_51_groupi_n_2085);
  not csa_tree_add_12_51_groupi_drc_bufs21769(csa_tree_add_12_51_groupi_n_2085 ,csa_tree_add_12_51_groupi_n_2946);
  not csa_tree_add_12_51_groupi_drc_bufs21782(csa_tree_add_12_51_groupi_n_2084 ,csa_tree_add_12_51_groupi_n_2083);
  not csa_tree_add_12_51_groupi_drc_bufs21784(csa_tree_add_12_51_groupi_n_2083 ,csa_tree_add_12_51_groupi_n_2938);
  not csa_tree_add_12_51_groupi_drc_bufs21792(csa_tree_add_12_51_groupi_n_2082 ,csa_tree_add_12_51_groupi_n_2081);
  not csa_tree_add_12_51_groupi_drc_bufs21794(csa_tree_add_12_51_groupi_n_2081 ,csa_tree_add_12_51_groupi_n_2934);
  not csa_tree_add_12_51_groupi_drc_bufs21812(csa_tree_add_12_51_groupi_n_2080 ,csa_tree_add_12_51_groupi_n_2079);
  not csa_tree_add_12_51_groupi_drc_bufs21814(csa_tree_add_12_51_groupi_n_2079 ,csa_tree_add_12_51_groupi_n_2506);
  not csa_tree_add_12_51_groupi_drc_bufs21817(csa_tree_add_12_51_groupi_n_2078 ,csa_tree_add_12_51_groupi_n_2077);
  not csa_tree_add_12_51_groupi_drc_bufs21819(csa_tree_add_12_51_groupi_n_2077 ,csa_tree_add_12_51_groupi_n_2505);
  not csa_tree_add_12_51_groupi_drc_bufs21827(csa_tree_add_12_51_groupi_n_2076 ,csa_tree_add_12_51_groupi_n_2075);
  not csa_tree_add_12_51_groupi_drc_bufs21829(csa_tree_add_12_51_groupi_n_2075 ,csa_tree_add_12_51_groupi_n_2930);
  not csa_tree_add_12_51_groupi_drc_bufs21832(csa_tree_add_12_51_groupi_n_2074 ,csa_tree_add_12_51_groupi_n_2073);
  not csa_tree_add_12_51_groupi_drc_bufs21834(csa_tree_add_12_51_groupi_n_2073 ,csa_tree_add_12_51_groupi_n_2928);
  not csa_tree_add_12_51_groupi_drc_bufs21847(csa_tree_add_12_51_groupi_n_2072 ,csa_tree_add_12_51_groupi_n_2071);
  not csa_tree_add_12_51_groupi_drc_bufs21849(csa_tree_add_12_51_groupi_n_2071 ,csa_tree_add_12_51_groupi_n_2937);
  not csa_tree_add_12_51_groupi_drc_bufs21852(csa_tree_add_12_51_groupi_n_2070 ,csa_tree_add_12_51_groupi_n_2069);
  not csa_tree_add_12_51_groupi_drc_bufs21854(csa_tree_add_12_51_groupi_n_2069 ,csa_tree_add_12_51_groupi_n_2935);
  not csa_tree_add_12_51_groupi_drc_bufs21862(csa_tree_add_12_51_groupi_n_2068 ,csa_tree_add_12_51_groupi_n_2067);
  not csa_tree_add_12_51_groupi_drc_bufs21864(csa_tree_add_12_51_groupi_n_2067 ,csa_tree_add_12_51_groupi_n_2943);
  not csa_tree_add_12_51_groupi_drc_bufs21872(csa_tree_add_12_51_groupi_n_2066 ,csa_tree_add_12_51_groupi_n_2065);
  not csa_tree_add_12_51_groupi_drc_bufs21874(csa_tree_add_12_51_groupi_n_2065 ,csa_tree_add_12_51_groupi_n_3505);
  not csa_tree_add_12_51_groupi_drc_bufs21877(csa_tree_add_12_51_groupi_n_2064 ,csa_tree_add_12_51_groupi_n_2063);
  not csa_tree_add_12_51_groupi_drc_bufs21879(csa_tree_add_12_51_groupi_n_2063 ,csa_tree_add_12_51_groupi_n_3508);
  not csa_tree_add_12_51_groupi_drc_bufs21882(csa_tree_add_12_51_groupi_n_2062 ,csa_tree_add_12_51_groupi_n_2061);
  not csa_tree_add_12_51_groupi_drc_bufs21884(csa_tree_add_12_51_groupi_n_2061 ,csa_tree_add_12_51_groupi_n_3507);
  not csa_tree_add_12_51_groupi_drc_bufs21892(csa_tree_add_12_51_groupi_n_2060 ,csa_tree_add_12_51_groupi_n_2059);
  not csa_tree_add_12_51_groupi_drc_bufs21894(csa_tree_add_12_51_groupi_n_2059 ,csa_tree_add_12_51_groupi_n_2931);
  not csa_tree_add_12_51_groupi_drc_bufs21897(csa_tree_add_12_51_groupi_n_2058 ,csa_tree_add_12_51_groupi_n_2057);
  not csa_tree_add_12_51_groupi_drc_bufs21899(csa_tree_add_12_51_groupi_n_2057 ,csa_tree_add_12_51_groupi_n_3500);
  not csa_tree_add_12_51_groupi_drc_bufs21907(csa_tree_add_12_51_groupi_n_2056 ,csa_tree_add_12_51_groupi_n_2055);
  not csa_tree_add_12_51_groupi_drc_bufs21909(csa_tree_add_12_51_groupi_n_2055 ,csa_tree_add_12_51_groupi_n_3498);
  not csa_tree_add_12_51_groupi_drc_bufs21912(csa_tree_add_12_51_groupi_n_2054 ,csa_tree_add_12_51_groupi_n_2053);
  not csa_tree_add_12_51_groupi_drc_bufs21914(csa_tree_add_12_51_groupi_n_2053 ,csa_tree_add_12_51_groupi_n_3497);
  not csa_tree_add_12_51_groupi_drc_bufs21917(csa_tree_add_12_51_groupi_n_2052 ,csa_tree_add_12_51_groupi_n_2051);
  not csa_tree_add_12_51_groupi_drc_bufs21919(csa_tree_add_12_51_groupi_n_2051 ,csa_tree_add_12_51_groupi_n_2932);
  not csa_tree_add_12_51_groupi_drc_bufs21922(csa_tree_add_12_51_groupi_n_2050 ,csa_tree_add_12_51_groupi_n_2049);
  not csa_tree_add_12_51_groupi_drc_bufs21924(csa_tree_add_12_51_groupi_n_2049 ,csa_tree_add_12_51_groupi_n_2940);
  not csa_tree_add_12_51_groupi_drc_bufs21932(csa_tree_add_12_51_groupi_n_2048 ,csa_tree_add_12_51_groupi_n_2047);
  not csa_tree_add_12_51_groupi_drc_bufs21934(csa_tree_add_12_51_groupi_n_2047 ,csa_tree_add_12_51_groupi_n_2922);
  not csa_tree_add_12_51_groupi_drc_bufs21937(csa_tree_add_12_51_groupi_n_2046 ,csa_tree_add_12_51_groupi_n_2045);
  not csa_tree_add_12_51_groupi_drc_bufs21939(csa_tree_add_12_51_groupi_n_2045 ,csa_tree_add_12_51_groupi_n_2947);
  not csa_tree_add_12_51_groupi_drc_bufs21942(csa_tree_add_12_51_groupi_n_2044 ,csa_tree_add_12_51_groupi_n_2043);
  not csa_tree_add_12_51_groupi_drc_bufs21944(csa_tree_add_12_51_groupi_n_2043 ,csa_tree_add_12_51_groupi_n_3504);
  not csa_tree_add_12_51_groupi_drc_bufs21947(csa_tree_add_12_51_groupi_n_2042 ,csa_tree_add_12_51_groupi_n_2041);
  not csa_tree_add_12_51_groupi_drc_bufs21949(csa_tree_add_12_51_groupi_n_2041 ,csa_tree_add_12_51_groupi_n_2945);
  not csa_tree_add_12_51_groupi_drc_bufs21952(csa_tree_add_12_51_groupi_n_2040 ,csa_tree_add_12_51_groupi_n_2039);
  not csa_tree_add_12_51_groupi_drc_bufs21954(csa_tree_add_12_51_groupi_n_2039 ,csa_tree_add_12_51_groupi_n_2944);
  not csa_tree_add_12_51_groupi_drc_bufs21957(csa_tree_add_12_51_groupi_n_2038 ,csa_tree_add_12_51_groupi_n_2037);
  not csa_tree_add_12_51_groupi_drc_bufs21959(csa_tree_add_12_51_groupi_n_2037 ,csa_tree_add_12_51_groupi_n_3506);
  not csa_tree_add_12_51_groupi_drc_bufs21967(csa_tree_add_12_51_groupi_n_2036 ,csa_tree_add_12_51_groupi_n_2035);
  not csa_tree_add_12_51_groupi_drc_bufs21969(csa_tree_add_12_51_groupi_n_2035 ,csa_tree_add_12_51_groupi_n_2929);
  not csa_tree_add_12_51_groupi_drc_bufs21972(csa_tree_add_12_51_groupi_n_2034 ,csa_tree_add_12_51_groupi_n_2033);
  not csa_tree_add_12_51_groupi_drc_bufs21974(csa_tree_add_12_51_groupi_n_2033 ,csa_tree_add_12_51_groupi_n_3501);
  not csa_tree_add_12_51_groupi_drc_bufs21982(csa_tree_add_12_51_groupi_n_2032 ,csa_tree_add_12_51_groupi_n_2031);
  not csa_tree_add_12_51_groupi_drc_bufs21984(csa_tree_add_12_51_groupi_n_2031 ,csa_tree_add_12_51_groupi_n_3503);
  not csa_tree_add_12_51_groupi_drc_bufs21987(csa_tree_add_12_51_groupi_n_2030 ,csa_tree_add_12_51_groupi_n_2029);
  not csa_tree_add_12_51_groupi_drc_bufs21989(csa_tree_add_12_51_groupi_n_2029 ,csa_tree_add_12_51_groupi_n_3502);
  not csa_tree_add_12_51_groupi_drc_bufs21992(csa_tree_add_12_51_groupi_n_2028 ,csa_tree_add_12_51_groupi_n_2027);
  not csa_tree_add_12_51_groupi_drc_bufs21994(csa_tree_add_12_51_groupi_n_2027 ,csa_tree_add_12_51_groupi_n_3499);
  not csa_tree_add_12_51_groupi_drc_bufs21997(csa_tree_add_12_51_groupi_n_2026 ,csa_tree_add_12_51_groupi_n_2025);
  not csa_tree_add_12_51_groupi_drc_bufs21999(csa_tree_add_12_51_groupi_n_2025 ,csa_tree_add_12_51_groupi_n_2752);
  not csa_tree_add_12_51_groupi_drc_bufs22007(csa_tree_add_12_51_groupi_n_2024 ,csa_tree_add_12_51_groupi_n_2023);
  not csa_tree_add_12_51_groupi_drc_bufs22009(csa_tree_add_12_51_groupi_n_2023 ,csa_tree_add_12_51_groupi_n_2939);
  not csa_tree_add_12_51_groupi_drc_bufs22012(csa_tree_add_12_51_groupi_n_2022 ,csa_tree_add_12_51_groupi_n_2021);
  not csa_tree_add_12_51_groupi_drc_bufs22014(csa_tree_add_12_51_groupi_n_2021 ,csa_tree_add_12_51_groupi_n_2924);
  not csa_tree_add_12_51_groupi_drc_bufs22017(csa_tree_add_12_51_groupi_n_2020 ,csa_tree_add_12_51_groupi_n_2019);
  not csa_tree_add_12_51_groupi_drc_bufs22019(csa_tree_add_12_51_groupi_n_2019 ,csa_tree_add_12_51_groupi_n_2942);
  not csa_tree_add_12_51_groupi_drc_bufs22022(csa_tree_add_12_51_groupi_n_2018 ,csa_tree_add_12_51_groupi_n_2017);
  not csa_tree_add_12_51_groupi_drc_bufs22024(csa_tree_add_12_51_groupi_n_2017 ,csa_tree_add_12_51_groupi_n_2941);
  not csa_tree_add_12_51_groupi_drc_bufs22107(csa_tree_add_12_51_groupi_n_2016 ,csa_tree_add_12_51_groupi_n_2015);
  not csa_tree_add_12_51_groupi_drc_bufs22109(csa_tree_add_12_51_groupi_n_2015 ,csa_tree_add_12_51_groupi_n_2753);
  not csa_tree_add_12_51_groupi_drc_bufs22117(csa_tree_add_12_51_groupi_n_2014 ,csa_tree_add_12_51_groupi_n_2013);
  not csa_tree_add_12_51_groupi_drc_bufs22119(csa_tree_add_12_51_groupi_n_2013 ,csa_tree_add_12_51_groupi_n_2933);
  not csa_tree_add_12_51_groupi_drc_bufs22122(csa_tree_add_12_51_groupi_n_2012 ,csa_tree_add_12_51_groupi_n_2011);
  not csa_tree_add_12_51_groupi_drc_bufs22124(csa_tree_add_12_51_groupi_n_2011 ,csa_tree_add_12_51_groupi_n_2637);
  not csa_tree_add_12_51_groupi_drc_bufs22127(csa_tree_add_12_51_groupi_n_2010 ,csa_tree_add_12_51_groupi_n_2009);
  not csa_tree_add_12_51_groupi_drc_bufs22129(csa_tree_add_12_51_groupi_n_2009 ,csa_tree_add_12_51_groupi_n_2638);
  not csa_tree_add_12_51_groupi_drc_bufs22516(csa_tree_add_12_51_groupi_n_2008 ,csa_tree_add_12_51_groupi_n_2006);
  not csa_tree_add_12_51_groupi_drc_bufs22517(csa_tree_add_12_51_groupi_n_2007 ,csa_tree_add_12_51_groupi_n_2006);
  not csa_tree_add_12_51_groupi_drc_bufs22518(csa_tree_add_12_51_groupi_n_2006 ,csa_tree_add_12_51_groupi_n_3229);
  not csa_tree_add_12_51_groupi_drc_bufs22520(csa_tree_add_12_51_groupi_n_2005 ,csa_tree_add_12_51_groupi_n_2003);
  not csa_tree_add_12_51_groupi_drc_bufs22521(csa_tree_add_12_51_groupi_n_2004 ,csa_tree_add_12_51_groupi_n_2003);
  not csa_tree_add_12_51_groupi_drc_bufs22522(csa_tree_add_12_51_groupi_n_2003 ,csa_tree_add_12_51_groupi_n_5175);
  not csa_tree_add_12_51_groupi_drc_bufs22524(csa_tree_add_12_51_groupi_n_2002 ,csa_tree_add_12_51_groupi_n_2000);
  not csa_tree_add_12_51_groupi_drc_bufs22525(csa_tree_add_12_51_groupi_n_2001 ,csa_tree_add_12_51_groupi_n_2000);
  not csa_tree_add_12_51_groupi_drc_bufs22526(csa_tree_add_12_51_groupi_n_2000 ,csa_tree_add_12_51_groupi_n_6024);
  not csa_tree_add_12_51_groupi_drc_bufs22528(csa_tree_add_12_51_groupi_n_1999 ,csa_tree_add_12_51_groupi_n_1997);
  not csa_tree_add_12_51_groupi_drc_bufs22529(csa_tree_add_12_51_groupi_n_1998 ,csa_tree_add_12_51_groupi_n_1997);
  not csa_tree_add_12_51_groupi_drc_bufs22530(csa_tree_add_12_51_groupi_n_1997 ,csa_tree_add_12_51_groupi_n_5842);
  not csa_tree_add_12_51_groupi_drc_bufs22532(csa_tree_add_12_51_groupi_n_1996 ,csa_tree_add_12_51_groupi_n_1994);
  not csa_tree_add_12_51_groupi_drc_bufs22533(csa_tree_add_12_51_groupi_n_1995 ,csa_tree_add_12_51_groupi_n_1994);
  not csa_tree_add_12_51_groupi_drc_bufs22534(csa_tree_add_12_51_groupi_n_1994 ,csa_tree_add_12_51_groupi_n_2643);
  not csa_tree_add_12_51_groupi_drc_bufs22536(csa_tree_add_12_51_groupi_n_1993 ,csa_tree_add_12_51_groupi_n_1991);
  not csa_tree_add_12_51_groupi_drc_bufs22537(csa_tree_add_12_51_groupi_n_1992 ,csa_tree_add_12_51_groupi_n_1991);
  not csa_tree_add_12_51_groupi_drc_bufs22538(csa_tree_add_12_51_groupi_n_1991 ,csa_tree_add_12_51_groupi_n_3764);
  not csa_tree_add_12_51_groupi_drc_bufs22540(csa_tree_add_12_51_groupi_n_1990 ,csa_tree_add_12_51_groupi_n_1988);
  not csa_tree_add_12_51_groupi_drc_bufs22541(csa_tree_add_12_51_groupi_n_1989 ,csa_tree_add_12_51_groupi_n_1988);
  not csa_tree_add_12_51_groupi_drc_bufs22542(csa_tree_add_12_51_groupi_n_1988 ,csa_tree_add_12_51_groupi_n_5020);
  not csa_tree_add_12_51_groupi_drc_bufs22544(csa_tree_add_12_51_groupi_n_1987 ,csa_tree_add_12_51_groupi_n_1985);
  not csa_tree_add_12_51_groupi_drc_bufs22545(csa_tree_add_12_51_groupi_n_1986 ,csa_tree_add_12_51_groupi_n_1985);
  not csa_tree_add_12_51_groupi_drc_bufs22546(csa_tree_add_12_51_groupi_n_1985 ,csa_tree_add_12_51_groupi_n_5676);
  not csa_tree_add_12_51_groupi_drc_bufs22548(csa_tree_add_12_51_groupi_n_1984 ,csa_tree_add_12_51_groupi_n_1982);
  not csa_tree_add_12_51_groupi_drc_bufs22549(csa_tree_add_12_51_groupi_n_1983 ,csa_tree_add_12_51_groupi_n_1982);
  not csa_tree_add_12_51_groupi_drc_bufs22550(csa_tree_add_12_51_groupi_n_1982 ,csa_tree_add_12_51_groupi_n_4839);
  not csa_tree_add_12_51_groupi_drc_bufs22552(csa_tree_add_12_51_groupi_n_1981 ,csa_tree_add_12_51_groupi_n_1979);
  not csa_tree_add_12_51_groupi_drc_bufs22553(csa_tree_add_12_51_groupi_n_1980 ,csa_tree_add_12_51_groupi_n_1979);
  not csa_tree_add_12_51_groupi_drc_bufs22554(csa_tree_add_12_51_groupi_n_1979 ,csa_tree_add_12_51_groupi_n_4665);
  not csa_tree_add_12_51_groupi_drc_bufs22556(csa_tree_add_12_51_groupi_n_1978 ,csa_tree_add_12_51_groupi_n_1976);
  not csa_tree_add_12_51_groupi_drc_bufs22557(csa_tree_add_12_51_groupi_n_1977 ,csa_tree_add_12_51_groupi_n_1976);
  not csa_tree_add_12_51_groupi_drc_bufs22558(csa_tree_add_12_51_groupi_n_1976 ,csa_tree_add_12_51_groupi_n_4299);
  not csa_tree_add_12_51_groupi_drc_bufs22560(csa_tree_add_12_51_groupi_n_1975 ,csa_tree_add_12_51_groupi_n_1973);
  not csa_tree_add_12_51_groupi_drc_bufs22561(csa_tree_add_12_51_groupi_n_1974 ,csa_tree_add_12_51_groupi_n_1973);
  not csa_tree_add_12_51_groupi_drc_bufs22562(csa_tree_add_12_51_groupi_n_1973 ,csa_tree_add_12_51_groupi_n_5499);
  not csa_tree_add_12_51_groupi_drc_bufs22564(csa_tree_add_12_51_groupi_n_1972 ,csa_tree_add_12_51_groupi_n_1970);
  not csa_tree_add_12_51_groupi_drc_bufs22565(csa_tree_add_12_51_groupi_n_1971 ,csa_tree_add_12_51_groupi_n_1970);
  not csa_tree_add_12_51_groupi_drc_bufs22566(csa_tree_add_12_51_groupi_n_1970 ,csa_tree_add_12_51_groupi_n_5346);
  not csa_tree_add_12_51_groupi_drc_bufs22568(csa_tree_add_12_51_groupi_n_1969 ,csa_tree_add_12_51_groupi_n_1967);
  not csa_tree_add_12_51_groupi_drc_bufs22569(csa_tree_add_12_51_groupi_n_1968 ,csa_tree_add_12_51_groupi_n_1967);
  not csa_tree_add_12_51_groupi_drc_bufs22570(csa_tree_add_12_51_groupi_n_1967 ,csa_tree_add_12_51_groupi_n_4126);
  not csa_tree_add_12_51_groupi_drc_bufs22572(csa_tree_add_12_51_groupi_n_1966 ,csa_tree_add_12_51_groupi_n_1964);
  not csa_tree_add_12_51_groupi_drc_bufs22573(csa_tree_add_12_51_groupi_n_1965 ,csa_tree_add_12_51_groupi_n_1964);
  not csa_tree_add_12_51_groupi_drc_bufs22574(csa_tree_add_12_51_groupi_n_1964 ,csa_tree_add_12_51_groupi_n_4487);
  not csa_tree_add_12_51_groupi_drc_bufs22576(csa_tree_add_12_51_groupi_n_1963 ,csa_tree_add_12_51_groupi_n_1961);
  not csa_tree_add_12_51_groupi_drc_bufs22577(csa_tree_add_12_51_groupi_n_1962 ,csa_tree_add_12_51_groupi_n_1961);
  not csa_tree_add_12_51_groupi_drc_bufs22578(csa_tree_add_12_51_groupi_n_1961 ,csa_tree_add_12_51_groupi_n_6206);
  not csa_tree_add_12_51_groupi_drc_bufs22792(csa_tree_add_12_51_groupi_n_1960 ,csa_tree_add_12_51_groupi_n_1958);
  not csa_tree_add_12_51_groupi_drc_bufs22793(csa_tree_add_12_51_groupi_n_1959 ,csa_tree_add_12_51_groupi_n_1958);
  not csa_tree_add_12_51_groupi_drc_bufs22794(csa_tree_add_12_51_groupi_n_1958 ,csa_tree_add_12_51_groupi_n_2364);
  not csa_tree_add_12_51_groupi_drc_bufs22801(csa_tree_add_12_51_groupi_n_1957 ,csa_tree_add_12_51_groupi_n_1956);
  not csa_tree_add_12_51_groupi_drc_bufs22802(csa_tree_add_12_51_groupi_n_1956 ,csa_tree_add_12_51_groupi_n_2398);
  not csa_tree_add_12_51_groupi_drc_bufs22804(csa_tree_add_12_51_groupi_n_1955 ,csa_tree_add_12_51_groupi_n_1954);
  not csa_tree_add_12_51_groupi_drc_bufs22806(csa_tree_add_12_51_groupi_n_1954 ,csa_tree_add_12_51_groupi_n_2404);
  not csa_tree_add_12_51_groupi_drc_bufs22808(csa_tree_add_12_51_groupi_n_1953 ,csa_tree_add_12_51_groupi_n_1952);
  not csa_tree_add_12_51_groupi_drc_bufs22810(csa_tree_add_12_51_groupi_n_1952 ,csa_tree_add_12_51_groupi_n_2400);
  not csa_tree_add_12_51_groupi_drc_bufs22813(csa_tree_add_12_51_groupi_n_1951 ,csa_tree_add_12_51_groupi_n_1950);
  not csa_tree_add_12_51_groupi_drc_bufs22814(csa_tree_add_12_51_groupi_n_1950 ,csa_tree_add_12_51_groupi_n_2363);
  not csa_tree_add_12_51_groupi_drc_bufs22817(csa_tree_add_12_51_groupi_n_1949 ,csa_tree_add_12_51_groupi_n_1948);
  not csa_tree_add_12_51_groupi_drc_bufs22818(csa_tree_add_12_51_groupi_n_1948 ,csa_tree_add_12_51_groupi_n_2397);
  not csa_tree_add_12_51_groupi_drc_bufs22821(csa_tree_add_12_51_groupi_n_1947 ,csa_tree_add_12_51_groupi_n_1946);
  not csa_tree_add_12_51_groupi_drc_bufs22822(csa_tree_add_12_51_groupi_n_1946 ,csa_tree_add_12_51_groupi_n_2403);
  not csa_tree_add_12_51_groupi_drc_bufs22824(csa_tree_add_12_51_groupi_n_1945 ,csa_tree_add_12_51_groupi_n_1943);
  not csa_tree_add_12_51_groupi_drc_bufs22825(csa_tree_add_12_51_groupi_n_1944 ,csa_tree_add_12_51_groupi_n_1943);
  not csa_tree_add_12_51_groupi_drc_bufs22826(csa_tree_add_12_51_groupi_n_1943 ,csa_tree_add_12_51_groupi_n_2400);
  not csa_tree_add_12_51_groupi_drc_bufs22828(csa_tree_add_12_51_groupi_n_1942 ,csa_tree_add_12_51_groupi_n_1940);
  not csa_tree_add_12_51_groupi_drc_bufs22829(csa_tree_add_12_51_groupi_n_1941 ,csa_tree_add_12_51_groupi_n_1940);
  not csa_tree_add_12_51_groupi_drc_bufs22830(csa_tree_add_12_51_groupi_n_1940 ,csa_tree_add_12_51_groupi_n_2399);
  not csa_tree_add_12_51_groupi_drc_bufs22832(csa_tree_add_12_51_groupi_n_1939 ,csa_tree_add_12_51_groupi_n_1937);
  not csa_tree_add_12_51_groupi_drc_bufs22833(csa_tree_add_12_51_groupi_n_1938 ,csa_tree_add_12_51_groupi_n_1937);
  not csa_tree_add_12_51_groupi_drc_bufs22834(csa_tree_add_12_51_groupi_n_1937 ,csa_tree_add_12_51_groupi_n_2398);
  not csa_tree_add_12_51_groupi_drc_bufs22836(csa_tree_add_12_51_groupi_n_1936 ,csa_tree_add_12_51_groupi_n_1934);
  not csa_tree_add_12_51_groupi_drc_bufs22837(csa_tree_add_12_51_groupi_n_1935 ,csa_tree_add_12_51_groupi_n_1934);
  not csa_tree_add_12_51_groupi_drc_bufs22838(csa_tree_add_12_51_groupi_n_1934 ,csa_tree_add_12_51_groupi_n_2401);
  not csa_tree_add_12_51_groupi_drc_bufs22840(csa_tree_add_12_51_groupi_n_1933 ,csa_tree_add_12_51_groupi_n_1931);
  not csa_tree_add_12_51_groupi_drc_bufs22841(csa_tree_add_12_51_groupi_n_1932 ,csa_tree_add_12_51_groupi_n_1931);
  not csa_tree_add_12_51_groupi_drc_bufs22842(csa_tree_add_12_51_groupi_n_1931 ,csa_tree_add_12_51_groupi_n_2401);
  not csa_tree_add_12_51_groupi_drc_bufs22844(csa_tree_add_12_51_groupi_n_1930 ,csa_tree_add_12_51_groupi_n_1928);
  not csa_tree_add_12_51_groupi_drc_bufs22845(csa_tree_add_12_51_groupi_n_1929 ,csa_tree_add_12_51_groupi_n_1928);
  not csa_tree_add_12_51_groupi_drc_bufs22846(csa_tree_add_12_51_groupi_n_1928 ,csa_tree_add_12_51_groupi_n_2404);
  not csa_tree_add_12_51_groupi_drc_bufs22848(csa_tree_add_12_51_groupi_n_1927 ,csa_tree_add_12_51_groupi_n_1925);
  not csa_tree_add_12_51_groupi_drc_bufs22849(csa_tree_add_12_51_groupi_n_1926 ,csa_tree_add_12_51_groupi_n_1925);
  not csa_tree_add_12_51_groupi_drc_bufs22850(csa_tree_add_12_51_groupi_n_1925 ,csa_tree_add_12_51_groupi_n_2363);
  not csa_tree_add_12_51_groupi_drc_bufs22852(csa_tree_add_12_51_groupi_n_1924 ,csa_tree_add_12_51_groupi_n_1922);
  not csa_tree_add_12_51_groupi_drc_bufs22853(csa_tree_add_12_51_groupi_n_1923 ,csa_tree_add_12_51_groupi_n_1922);
  not csa_tree_add_12_51_groupi_drc_bufs22854(csa_tree_add_12_51_groupi_n_1922 ,csa_tree_add_12_51_groupi_n_2397);
  not csa_tree_add_12_51_groupi_drc_bufs22856(csa_tree_add_12_51_groupi_n_1921 ,csa_tree_add_12_51_groupi_n_1919);
  not csa_tree_add_12_51_groupi_drc_bufs22857(csa_tree_add_12_51_groupi_n_1920 ,csa_tree_add_12_51_groupi_n_1919);
  not csa_tree_add_12_51_groupi_drc_bufs22858(csa_tree_add_12_51_groupi_n_1919 ,csa_tree_add_12_51_groupi_n_2403);
  not csa_tree_add_12_51_groupi_drc_bufs22860(csa_tree_add_12_51_groupi_n_1918 ,csa_tree_add_12_51_groupi_n_1917);
  not csa_tree_add_12_51_groupi_drc_bufs22862(csa_tree_add_12_51_groupi_n_1917 ,csa_tree_add_12_51_groupi_n_2366);
  not csa_tree_add_12_51_groupi_drc_bufs22864(csa_tree_add_12_51_groupi_n_1916 ,csa_tree_add_12_51_groupi_n_1915);
  not csa_tree_add_12_51_groupi_drc_bufs22866(csa_tree_add_12_51_groupi_n_1915 ,csa_tree_add_12_51_groupi_n_2367);
  not csa_tree_add_12_51_groupi_drc_bufs22872(csa_tree_add_12_51_groupi_n_1914 ,csa_tree_add_12_51_groupi_n_1913);
  not csa_tree_add_12_51_groupi_drc_bufs22873(csa_tree_add_12_51_groupi_n_1913 ,csa_tree_add_12_51_groupi_n_3230);
  not csa_tree_add_12_51_groupi_drc_bufs22876(csa_tree_add_12_51_groupi_n_1912 ,csa_tree_add_12_51_groupi_n_1911);
  not csa_tree_add_12_51_groupi_drc_bufs22877(csa_tree_add_12_51_groupi_n_1911 ,csa_tree_add_12_51_groupi_n_3513);
  not csa_tree_add_12_51_groupi_drc_bufs22880(csa_tree_add_12_51_groupi_n_1910 ,csa_tree_add_12_51_groupi_n_1909);
  not csa_tree_add_12_51_groupi_drc_bufs22881(csa_tree_add_12_51_groupi_n_1909 ,csa_tree_add_12_51_groupi_n_3511);
  not csa_tree_add_12_51_groupi_drc_bufs22883(csa_tree_add_12_51_groupi_n_1908 ,csa_tree_add_12_51_groupi_n_2350);
  not csa_tree_add_12_51_groupi_drc_bufs22885(csa_tree_add_12_51_groupi_n_2350 ,csa_tree_add_12_51_groupi_n_2641);
  not csa_tree_add_12_51_groupi_drc_bufs22887(csa_tree_add_12_51_groupi_n_1907 ,csa_tree_add_12_51_groupi_n_2347);
  not csa_tree_add_12_51_groupi_drc_bufs22889(csa_tree_add_12_51_groupi_n_2347 ,csa_tree_add_12_51_groupi_n_2460);
  not csa_tree_add_12_51_groupi_drc_bufs22891(csa_tree_add_12_51_groupi_n_1906 ,csa_tree_add_12_51_groupi_n_2348);
  not csa_tree_add_12_51_groupi_drc_bufs22893(csa_tree_add_12_51_groupi_n_2348 ,csa_tree_add_12_51_groupi_n_2466);
  not csa_tree_add_12_51_groupi_drc_bufs22895(csa_tree_add_12_51_groupi_n_1905 ,csa_tree_add_12_51_groupi_n_2349);
  not csa_tree_add_12_51_groupi_drc_bufs22897(csa_tree_add_12_51_groupi_n_2349 ,csa_tree_add_12_51_groupi_n_2466);
  not csa_tree_add_12_51_groupi_drc_bufs22899(csa_tree_add_12_51_groupi_n_1904 ,csa_tree_add_12_51_groupi_n_2353);
  not csa_tree_add_12_51_groupi_drc_bufs22901(csa_tree_add_12_51_groupi_n_2353 ,csa_tree_add_12_51_groupi_n_6163);
  not csa_tree_add_12_51_groupi_drc_bufs22904(csa_tree_add_12_51_groupi_n_1903 ,csa_tree_add_12_51_groupi_n_1902);
  not csa_tree_add_12_51_groupi_drc_bufs22905(csa_tree_add_12_51_groupi_n_1902 ,csa_tree_add_12_51_groupi_n_2362);
  not csa_tree_add_12_51_groupi_drc_bufs22908(csa_tree_add_12_51_groupi_n_1901 ,csa_tree_add_12_51_groupi_n_1900);
  not csa_tree_add_12_51_groupi_drc_bufs22909(csa_tree_add_12_51_groupi_n_1900 ,csa_tree_add_12_51_groupi_n_2366);
  not csa_tree_add_12_51_groupi_drc_bufs22917(csa_tree_add_12_51_groupi_n_1899 ,csa_tree_add_12_51_groupi_n_1897);
  not csa_tree_add_12_51_groupi_drc_bufs22918(csa_tree_add_12_51_groupi_n_1898 ,csa_tree_add_12_51_groupi_n_1897);
  not csa_tree_add_12_51_groupi_drc_bufs22919(csa_tree_add_12_51_groupi_n_1897 ,csa_tree_add_12_51_groupi_n_2367);
  not csa_tree_add_12_51_groupi_drc_bufs22928(csa_tree_add_12_51_groupi_n_1896 ,csa_tree_add_12_51_groupi_n_1895);
  not csa_tree_add_12_51_groupi_drc_bufs22930(csa_tree_add_12_51_groupi_n_1895 ,csa_tree_add_12_51_groupi_n_2361);
  not csa_tree_add_12_51_groupi_drc_bufs22932(csa_tree_add_12_51_groupi_n_1894 ,csa_tree_add_12_51_groupi_n_1893);
  not csa_tree_add_12_51_groupi_drc_bufs22934(csa_tree_add_12_51_groupi_n_1893 ,csa_tree_add_12_51_groupi_n_2362);
  not csa_tree_add_12_51_groupi_drc_bufs22936(csa_tree_add_12_51_groupi_n_1892 ,csa_tree_add_12_51_groupi_n_1891);
  not csa_tree_add_12_51_groupi_drc_bufs22938(csa_tree_add_12_51_groupi_n_1891 ,csa_tree_add_12_51_groupi_n_2361);
  not csa_tree_add_12_51_groupi_drc_bufs22940(csa_tree_add_12_51_groupi_n_1890 ,csa_tree_add_12_51_groupi_n_1888);
  not csa_tree_add_12_51_groupi_drc_bufs22941(csa_tree_add_12_51_groupi_n_1889 ,csa_tree_add_12_51_groupi_n_1888);
  not csa_tree_add_12_51_groupi_drc_bufs22942(csa_tree_add_12_51_groupi_n_1888 ,csa_tree_add_12_51_groupi_n_2921);
  not csa_tree_add_12_51_groupi_drc_bufs22944(csa_tree_add_12_51_groupi_n_1887 ,csa_tree_add_12_51_groupi_n_1885);
  not csa_tree_add_12_51_groupi_drc_bufs22945(csa_tree_add_12_51_groupi_n_1886 ,csa_tree_add_12_51_groupi_n_1885);
  not csa_tree_add_12_51_groupi_drc_bufs22946(csa_tree_add_12_51_groupi_n_1885 ,csa_tree_add_12_51_groupi_n_2919);
  not csa_tree_add_12_51_groupi_drc_bufs22948(csa_tree_add_12_51_groupi_n_1884 ,csa_tree_add_12_51_groupi_n_1882);
  not csa_tree_add_12_51_groupi_drc_bufs22949(csa_tree_add_12_51_groupi_n_1883 ,csa_tree_add_12_51_groupi_n_1882);
  not csa_tree_add_12_51_groupi_drc_bufs22950(csa_tree_add_12_51_groupi_n_1882 ,csa_tree_add_12_51_groupi_n_2917);
  not csa_tree_add_12_51_groupi_drc_bufs22952(csa_tree_add_12_51_groupi_n_1881 ,csa_tree_add_12_51_groupi_n_1879);
  not csa_tree_add_12_51_groupi_drc_bufs22953(csa_tree_add_12_51_groupi_n_1880 ,csa_tree_add_12_51_groupi_n_1879);
  not csa_tree_add_12_51_groupi_drc_bufs22954(csa_tree_add_12_51_groupi_n_1879 ,csa_tree_add_12_51_groupi_n_2913);
  not csa_tree_add_12_51_groupi_drc_bufs22956(csa_tree_add_12_51_groupi_n_1878 ,csa_tree_add_12_51_groupi_n_1876);
  not csa_tree_add_12_51_groupi_drc_bufs22957(csa_tree_add_12_51_groupi_n_1877 ,csa_tree_add_12_51_groupi_n_1876);
  not csa_tree_add_12_51_groupi_drc_bufs22958(csa_tree_add_12_51_groupi_n_1876 ,csa_tree_add_12_51_groupi_n_2912);
  not csa_tree_add_12_51_groupi_drc_bufs22960(csa_tree_add_12_51_groupi_n_1875 ,csa_tree_add_12_51_groupi_n_1873);
  not csa_tree_add_12_51_groupi_drc_bufs22961(csa_tree_add_12_51_groupi_n_1874 ,csa_tree_add_12_51_groupi_n_1873);
  not csa_tree_add_12_51_groupi_drc_bufs22962(csa_tree_add_12_51_groupi_n_1873 ,csa_tree_add_12_51_groupi_n_2916);
  not csa_tree_add_12_51_groupi_drc_bufs22964(csa_tree_add_12_51_groupi_n_1872 ,csa_tree_add_12_51_groupi_n_1870);
  not csa_tree_add_12_51_groupi_drc_bufs22965(csa_tree_add_12_51_groupi_n_1871 ,csa_tree_add_12_51_groupi_n_1870);
  not csa_tree_add_12_51_groupi_drc_bufs22966(csa_tree_add_12_51_groupi_n_1870 ,csa_tree_add_12_51_groupi_n_2911);
  not csa_tree_add_12_51_groupi_drc_bufs22968(csa_tree_add_12_51_groupi_n_1869 ,csa_tree_add_12_51_groupi_n_1867);
  not csa_tree_add_12_51_groupi_drc_bufs22969(csa_tree_add_12_51_groupi_n_1868 ,csa_tree_add_12_51_groupi_n_1867);
  not csa_tree_add_12_51_groupi_drc_bufs22970(csa_tree_add_12_51_groupi_n_1867 ,csa_tree_add_12_51_groupi_n_2910);
  not csa_tree_add_12_51_groupi_drc_bufs22972(csa_tree_add_12_51_groupi_n_1866 ,csa_tree_add_12_51_groupi_n_1864);
  not csa_tree_add_12_51_groupi_drc_bufs22973(csa_tree_add_12_51_groupi_n_1865 ,csa_tree_add_12_51_groupi_n_1864);
  not csa_tree_add_12_51_groupi_drc_bufs22974(csa_tree_add_12_51_groupi_n_1864 ,csa_tree_add_12_51_groupi_n_2920);
  not csa_tree_add_12_51_groupi_drc_bufs22976(csa_tree_add_12_51_groupi_n_1863 ,csa_tree_add_12_51_groupi_n_1861);
  not csa_tree_add_12_51_groupi_drc_bufs22977(csa_tree_add_12_51_groupi_n_1862 ,csa_tree_add_12_51_groupi_n_1861);
  not csa_tree_add_12_51_groupi_drc_bufs22978(csa_tree_add_12_51_groupi_n_1861 ,csa_tree_add_12_51_groupi_n_2915);
  not csa_tree_add_12_51_groupi_drc_bufs22980(csa_tree_add_12_51_groupi_n_1860 ,csa_tree_add_12_51_groupi_n_1858);
  not csa_tree_add_12_51_groupi_drc_bufs22981(csa_tree_add_12_51_groupi_n_1859 ,csa_tree_add_12_51_groupi_n_1858);
  not csa_tree_add_12_51_groupi_drc_bufs22982(csa_tree_add_12_51_groupi_n_1858 ,csa_tree_add_12_51_groupi_n_2909);
  not csa_tree_add_12_51_groupi_drc_bufs22984(csa_tree_add_12_51_groupi_n_1857 ,csa_tree_add_12_51_groupi_n_1855);
  not csa_tree_add_12_51_groupi_drc_bufs22985(csa_tree_add_12_51_groupi_n_1856 ,csa_tree_add_12_51_groupi_n_1855);
  not csa_tree_add_12_51_groupi_drc_bufs22986(csa_tree_add_12_51_groupi_n_1855 ,csa_tree_add_12_51_groupi_n_2908);
  not csa_tree_add_12_51_groupi_drc_bufs22988(csa_tree_add_12_51_groupi_n_1854 ,csa_tree_add_12_51_groupi_n_1852);
  not csa_tree_add_12_51_groupi_drc_bufs22989(csa_tree_add_12_51_groupi_n_1853 ,csa_tree_add_12_51_groupi_n_1852);
  not csa_tree_add_12_51_groupi_drc_bufs22990(csa_tree_add_12_51_groupi_n_1852 ,csa_tree_add_12_51_groupi_n_2918);
  not csa_tree_add_12_51_groupi_drc_bufs22992(csa_tree_add_12_51_groupi_n_1851 ,csa_tree_add_12_51_groupi_n_1849);
  not csa_tree_add_12_51_groupi_drc_bufs22993(csa_tree_add_12_51_groupi_n_1850 ,csa_tree_add_12_51_groupi_n_1849);
  not csa_tree_add_12_51_groupi_drc_bufs22994(csa_tree_add_12_51_groupi_n_1849 ,csa_tree_add_12_51_groupi_n_2907);
  not csa_tree_add_12_51_groupi_drc_bufs22996(csa_tree_add_12_51_groupi_n_1848 ,csa_tree_add_12_51_groupi_n_1846);
  not csa_tree_add_12_51_groupi_drc_bufs22997(csa_tree_add_12_51_groupi_n_1847 ,csa_tree_add_12_51_groupi_n_1846);
  not csa_tree_add_12_51_groupi_drc_bufs22998(csa_tree_add_12_51_groupi_n_1846 ,csa_tree_add_12_51_groupi_n_2914);
  not csa_tree_add_12_51_groupi_drc_bufs23001(csa_tree_add_12_51_groupi_n_1845 ,csa_tree_add_12_51_groupi_n_1844);
  not csa_tree_add_12_51_groupi_drc_bufs23002(csa_tree_add_12_51_groupi_n_1844 ,csa_tree_add_12_51_groupi_n_2146);
  not csa_tree_add_12_51_groupi_drc_bufs23005(csa_tree_add_12_51_groupi_n_1843 ,csa_tree_add_12_51_groupi_n_1842);
  not csa_tree_add_12_51_groupi_drc_bufs23006(csa_tree_add_12_51_groupi_n_1842 ,csa_tree_add_12_51_groupi_n_2143);
  not csa_tree_add_12_51_groupi_drc_bufs23009(csa_tree_add_12_51_groupi_n_1841 ,csa_tree_add_12_51_groupi_n_1840);
  not csa_tree_add_12_51_groupi_drc_bufs23010(csa_tree_add_12_51_groupi_n_1840 ,csa_tree_add_12_51_groupi_n_2140);
  not csa_tree_add_12_51_groupi_drc_bufs23013(csa_tree_add_12_51_groupi_n_1839 ,csa_tree_add_12_51_groupi_n_1838);
  not csa_tree_add_12_51_groupi_drc_bufs23014(csa_tree_add_12_51_groupi_n_1838 ,csa_tree_add_12_51_groupi_n_2137);
  not csa_tree_add_12_51_groupi_drc_bufs23017(csa_tree_add_12_51_groupi_n_1837 ,csa_tree_add_12_51_groupi_n_1836);
  not csa_tree_add_12_51_groupi_drc_bufs23018(csa_tree_add_12_51_groupi_n_1836 ,csa_tree_add_12_51_groupi_n_2134);
  not csa_tree_add_12_51_groupi_drc_bufs23021(csa_tree_add_12_51_groupi_n_1835 ,csa_tree_add_12_51_groupi_n_1834);
  not csa_tree_add_12_51_groupi_drc_bufs23022(csa_tree_add_12_51_groupi_n_1834 ,csa_tree_add_12_51_groupi_n_2131);
  not csa_tree_add_12_51_groupi_drc_bufs23025(csa_tree_add_12_51_groupi_n_1833 ,csa_tree_add_12_51_groupi_n_1832);
  not csa_tree_add_12_51_groupi_drc_bufs23026(csa_tree_add_12_51_groupi_n_1832 ,csa_tree_add_12_51_groupi_n_2128);
  not csa_tree_add_12_51_groupi_drc_bufs23029(csa_tree_add_12_51_groupi_n_1831 ,csa_tree_add_12_51_groupi_n_1830);
  not csa_tree_add_12_51_groupi_drc_bufs23030(csa_tree_add_12_51_groupi_n_1830 ,csa_tree_add_12_51_groupi_n_2125);
  not csa_tree_add_12_51_groupi_drc_bufs23033(csa_tree_add_12_51_groupi_n_1829 ,csa_tree_add_12_51_groupi_n_1828);
  not csa_tree_add_12_51_groupi_drc_bufs23034(csa_tree_add_12_51_groupi_n_1828 ,csa_tree_add_12_51_groupi_n_2122);
  not csa_tree_add_12_51_groupi_drc_bufs23037(csa_tree_add_12_51_groupi_n_1827 ,csa_tree_add_12_51_groupi_n_1826);
  not csa_tree_add_12_51_groupi_drc_bufs23038(csa_tree_add_12_51_groupi_n_1826 ,csa_tree_add_12_51_groupi_n_2119);
  not csa_tree_add_12_51_groupi_drc_bufs23041(csa_tree_add_12_51_groupi_n_1825 ,csa_tree_add_12_51_groupi_n_1824);
  not csa_tree_add_12_51_groupi_drc_bufs23042(csa_tree_add_12_51_groupi_n_1824 ,csa_tree_add_12_51_groupi_n_2116);
  not csa_tree_add_12_51_groupi_drc_bufs23045(csa_tree_add_12_51_groupi_n_1823 ,csa_tree_add_12_51_groupi_n_1822);
  not csa_tree_add_12_51_groupi_drc_bufs23046(csa_tree_add_12_51_groupi_n_1822 ,csa_tree_add_12_51_groupi_n_2113);
  not csa_tree_add_12_51_groupi_drc_bufs23049(csa_tree_add_12_51_groupi_n_1821 ,csa_tree_add_12_51_groupi_n_1820);
  not csa_tree_add_12_51_groupi_drc_bufs23050(csa_tree_add_12_51_groupi_n_1820 ,csa_tree_add_12_51_groupi_n_2110);
  not csa_tree_add_12_51_groupi_drc_bufs23053(csa_tree_add_12_51_groupi_n_1819 ,csa_tree_add_12_51_groupi_n_1818);
  not csa_tree_add_12_51_groupi_drc_bufs23054(csa_tree_add_12_51_groupi_n_1818 ,csa_tree_add_12_51_groupi_n_2107);
  not csa_tree_add_12_51_groupi_drc_bufs23057(csa_tree_add_12_51_groupi_n_1817 ,csa_tree_add_12_51_groupi_n_1816);
  not csa_tree_add_12_51_groupi_drc_bufs23058(csa_tree_add_12_51_groupi_n_1816 ,csa_tree_add_12_51_groupi_n_2149);
  not csa_tree_add_12_51_groupi_drc_bufs23060(csa_tree_add_12_51_groupi_n_1815 ,csa_tree_add_12_51_groupi_n_1813);
  not csa_tree_add_12_51_groupi_drc_bufs23061(csa_tree_add_12_51_groupi_n_1814 ,csa_tree_add_12_51_groupi_n_1813);
  not csa_tree_add_12_51_groupi_drc_bufs23062(csa_tree_add_12_51_groupi_n_1813 ,csa_tree_add_12_51_groupi_n_2463);
  not csa_tree_add_12_51_groupi_drc_bufs23064(csa_tree_add_12_51_groupi_n_1812 ,csa_tree_add_12_51_groupi_n_1810);
  not csa_tree_add_12_51_groupi_drc_bufs23065(csa_tree_add_12_51_groupi_n_1811 ,csa_tree_add_12_51_groupi_n_1810);
  not csa_tree_add_12_51_groupi_drc_bufs23066(csa_tree_add_12_51_groupi_n_1810 ,csa_tree_add_12_51_groupi_n_2344);
  not csa_tree_add_12_51_groupi_drc_bufs23068(csa_tree_add_12_51_groupi_n_1809 ,csa_tree_add_12_51_groupi_n_1807);
  not csa_tree_add_12_51_groupi_drc_bufs23069(csa_tree_add_12_51_groupi_n_1808 ,csa_tree_add_12_51_groupi_n_1807);
  not csa_tree_add_12_51_groupi_drc_bufs23070(csa_tree_add_12_51_groupi_n_1807 ,csa_tree_add_12_51_groupi_n_2343);
  not csa_tree_add_12_51_groupi_drc_bufs23072(csa_tree_add_12_51_groupi_n_1806 ,csa_tree_add_12_51_groupi_n_1804);
  not csa_tree_add_12_51_groupi_drc_bufs23073(csa_tree_add_12_51_groupi_n_1805 ,csa_tree_add_12_51_groupi_n_1804);
  not csa_tree_add_12_51_groupi_drc_bufs23074(csa_tree_add_12_51_groupi_n_1804 ,csa_tree_add_12_51_groupi_n_2337);
  not csa_tree_add_12_51_groupi_drc_bufs23076(csa_tree_add_12_51_groupi_n_1803 ,csa_tree_add_12_51_groupi_n_1801);
  not csa_tree_add_12_51_groupi_drc_bufs23077(csa_tree_add_12_51_groupi_n_1802 ,csa_tree_add_12_51_groupi_n_1801);
  not csa_tree_add_12_51_groupi_drc_bufs23078(csa_tree_add_12_51_groupi_n_1801 ,csa_tree_add_12_51_groupi_n_2336);
  not csa_tree_add_12_51_groupi_drc_bufs23080(csa_tree_add_12_51_groupi_n_1800 ,csa_tree_add_12_51_groupi_n_1798);
  not csa_tree_add_12_51_groupi_drc_bufs23081(csa_tree_add_12_51_groupi_n_1799 ,csa_tree_add_12_51_groupi_n_1798);
  not csa_tree_add_12_51_groupi_drc_bufs23082(csa_tree_add_12_51_groupi_n_1798 ,csa_tree_add_12_51_groupi_n_2328);
  not csa_tree_add_12_51_groupi_drc_bufs23084(csa_tree_add_12_51_groupi_n_1797 ,csa_tree_add_12_51_groupi_n_1795);
  not csa_tree_add_12_51_groupi_drc_bufs23085(csa_tree_add_12_51_groupi_n_1796 ,csa_tree_add_12_51_groupi_n_1795);
  not csa_tree_add_12_51_groupi_drc_bufs23086(csa_tree_add_12_51_groupi_n_1795 ,csa_tree_add_12_51_groupi_n_2327);
  not csa_tree_add_12_51_groupi_drc_bufs23088(csa_tree_add_12_51_groupi_n_1794 ,csa_tree_add_12_51_groupi_n_1792);
  not csa_tree_add_12_51_groupi_drc_bufs23089(csa_tree_add_12_51_groupi_n_1793 ,csa_tree_add_12_51_groupi_n_1792);
  not csa_tree_add_12_51_groupi_drc_bufs23090(csa_tree_add_12_51_groupi_n_1792 ,csa_tree_add_12_51_groupi_n_2326);
  not csa_tree_add_12_51_groupi_drc_bufs23092(csa_tree_add_12_51_groupi_n_1791 ,csa_tree_add_12_51_groupi_n_1789);
  not csa_tree_add_12_51_groupi_drc_bufs23093(csa_tree_add_12_51_groupi_n_1790 ,csa_tree_add_12_51_groupi_n_1789);
  not csa_tree_add_12_51_groupi_drc_bufs23094(csa_tree_add_12_51_groupi_n_1789 ,csa_tree_add_12_51_groupi_n_2346);
  not csa_tree_add_12_51_groupi_drc_bufs23096(csa_tree_add_12_51_groupi_n_1788 ,csa_tree_add_12_51_groupi_n_1786);
  not csa_tree_add_12_51_groupi_drc_bufs23097(csa_tree_add_12_51_groupi_n_1787 ,csa_tree_add_12_51_groupi_n_1786);
  not csa_tree_add_12_51_groupi_drc_bufs23098(csa_tree_add_12_51_groupi_n_1786 ,csa_tree_add_12_51_groupi_n_2319);
  not csa_tree_add_12_51_groupi_drc_bufs23100(csa_tree_add_12_51_groupi_n_1785 ,csa_tree_add_12_51_groupi_n_1783);
  not csa_tree_add_12_51_groupi_drc_bufs23101(csa_tree_add_12_51_groupi_n_1784 ,csa_tree_add_12_51_groupi_n_1783);
  not csa_tree_add_12_51_groupi_drc_bufs23102(csa_tree_add_12_51_groupi_n_1783 ,csa_tree_add_12_51_groupi_n_2318);
  not csa_tree_add_12_51_groupi_drc_bufs23104(csa_tree_add_12_51_groupi_n_1782 ,csa_tree_add_12_51_groupi_n_1780);
  not csa_tree_add_12_51_groupi_drc_bufs23105(csa_tree_add_12_51_groupi_n_1781 ,csa_tree_add_12_51_groupi_n_1780);
  not csa_tree_add_12_51_groupi_drc_bufs23106(csa_tree_add_12_51_groupi_n_1780 ,csa_tree_add_12_51_groupi_n_2317);
  not csa_tree_add_12_51_groupi_drc_bufs23108(csa_tree_add_12_51_groupi_n_1779 ,csa_tree_add_12_51_groupi_n_1777);
  not csa_tree_add_12_51_groupi_drc_bufs23109(csa_tree_add_12_51_groupi_n_1778 ,csa_tree_add_12_51_groupi_n_1777);
  not csa_tree_add_12_51_groupi_drc_bufs23110(csa_tree_add_12_51_groupi_n_1777 ,csa_tree_add_12_51_groupi_n_2345);
  not csa_tree_add_12_51_groupi_drc_bufs23112(csa_tree_add_12_51_groupi_n_1776 ,csa_tree_add_12_51_groupi_n_1774);
  not csa_tree_add_12_51_groupi_drc_bufs23113(csa_tree_add_12_51_groupi_n_1775 ,csa_tree_add_12_51_groupi_n_1774);
  not csa_tree_add_12_51_groupi_drc_bufs23114(csa_tree_add_12_51_groupi_n_1774 ,csa_tree_add_12_51_groupi_n_2310);
  not csa_tree_add_12_51_groupi_drc_bufs23116(csa_tree_add_12_51_groupi_n_1773 ,csa_tree_add_12_51_groupi_n_1771);
  not csa_tree_add_12_51_groupi_drc_bufs23117(csa_tree_add_12_51_groupi_n_1772 ,csa_tree_add_12_51_groupi_n_1771);
  not csa_tree_add_12_51_groupi_drc_bufs23118(csa_tree_add_12_51_groupi_n_1771 ,csa_tree_add_12_51_groupi_n_2309);
  not csa_tree_add_12_51_groupi_drc_bufs23120(csa_tree_add_12_51_groupi_n_1770 ,csa_tree_add_12_51_groupi_n_1768);
  not csa_tree_add_12_51_groupi_drc_bufs23121(csa_tree_add_12_51_groupi_n_1769 ,csa_tree_add_12_51_groupi_n_1768);
  not csa_tree_add_12_51_groupi_drc_bufs23122(csa_tree_add_12_51_groupi_n_1768 ,csa_tree_add_12_51_groupi_n_2308);
  not csa_tree_add_12_51_groupi_drc_bufs23124(csa_tree_add_12_51_groupi_n_1767 ,csa_tree_add_12_51_groupi_n_1765);
  not csa_tree_add_12_51_groupi_drc_bufs23125(csa_tree_add_12_51_groupi_n_1766 ,csa_tree_add_12_51_groupi_n_1765);
  not csa_tree_add_12_51_groupi_drc_bufs23126(csa_tree_add_12_51_groupi_n_1765 ,csa_tree_add_12_51_groupi_n_2300);
  not csa_tree_add_12_51_groupi_drc_bufs23128(csa_tree_add_12_51_groupi_n_1764 ,csa_tree_add_12_51_groupi_n_1762);
  not csa_tree_add_12_51_groupi_drc_bufs23129(csa_tree_add_12_51_groupi_n_1763 ,csa_tree_add_12_51_groupi_n_1762);
  not csa_tree_add_12_51_groupi_drc_bufs23130(csa_tree_add_12_51_groupi_n_1762 ,csa_tree_add_12_51_groupi_n_2301);
  not csa_tree_add_12_51_groupi_drc_bufs23132(csa_tree_add_12_51_groupi_n_1761 ,csa_tree_add_12_51_groupi_n_1759);
  not csa_tree_add_12_51_groupi_drc_bufs23133(csa_tree_add_12_51_groupi_n_1760 ,csa_tree_add_12_51_groupi_n_1759);
  not csa_tree_add_12_51_groupi_drc_bufs23134(csa_tree_add_12_51_groupi_n_1759 ,csa_tree_add_12_51_groupi_n_2292);
  not csa_tree_add_12_51_groupi_drc_bufs23136(csa_tree_add_12_51_groupi_n_1758 ,csa_tree_add_12_51_groupi_n_1756);
  not csa_tree_add_12_51_groupi_drc_bufs23137(csa_tree_add_12_51_groupi_n_1757 ,csa_tree_add_12_51_groupi_n_1756);
  not csa_tree_add_12_51_groupi_drc_bufs23138(csa_tree_add_12_51_groupi_n_1756 ,csa_tree_add_12_51_groupi_n_2291);
  not csa_tree_add_12_51_groupi_drc_bufs23140(csa_tree_add_12_51_groupi_n_1755 ,csa_tree_add_12_51_groupi_n_1753);
  not csa_tree_add_12_51_groupi_drc_bufs23141(csa_tree_add_12_51_groupi_n_1754 ,csa_tree_add_12_51_groupi_n_1753);
  not csa_tree_add_12_51_groupi_drc_bufs23142(csa_tree_add_12_51_groupi_n_1753 ,csa_tree_add_12_51_groupi_n_2283);
  not csa_tree_add_12_51_groupi_drc_bufs23144(csa_tree_add_12_51_groupi_n_1752 ,csa_tree_add_12_51_groupi_n_1750);
  not csa_tree_add_12_51_groupi_drc_bufs23145(csa_tree_add_12_51_groupi_n_1751 ,csa_tree_add_12_51_groupi_n_1750);
  not csa_tree_add_12_51_groupi_drc_bufs23146(csa_tree_add_12_51_groupi_n_1750 ,csa_tree_add_12_51_groupi_n_2282);
  not csa_tree_add_12_51_groupi_drc_bufs23148(csa_tree_add_12_51_groupi_n_1749 ,csa_tree_add_12_51_groupi_n_1747);
  not csa_tree_add_12_51_groupi_drc_bufs23149(csa_tree_add_12_51_groupi_n_1748 ,csa_tree_add_12_51_groupi_n_1747);
  not csa_tree_add_12_51_groupi_drc_bufs23150(csa_tree_add_12_51_groupi_n_1747 ,csa_tree_add_12_51_groupi_n_2281);
  not csa_tree_add_12_51_groupi_drc_bufs23152(csa_tree_add_12_51_groupi_n_1746 ,csa_tree_add_12_51_groupi_n_1744);
  not csa_tree_add_12_51_groupi_drc_bufs23153(csa_tree_add_12_51_groupi_n_1745 ,csa_tree_add_12_51_groupi_n_1744);
  not csa_tree_add_12_51_groupi_drc_bufs23154(csa_tree_add_12_51_groupi_n_1744 ,csa_tree_add_12_51_groupi_n_2273);
  not csa_tree_add_12_51_groupi_drc_bufs23156(csa_tree_add_12_51_groupi_n_1743 ,csa_tree_add_12_51_groupi_n_1741);
  not csa_tree_add_12_51_groupi_drc_bufs23157(csa_tree_add_12_51_groupi_n_1742 ,csa_tree_add_12_51_groupi_n_1741);
  not csa_tree_add_12_51_groupi_drc_bufs23158(csa_tree_add_12_51_groupi_n_1741 ,csa_tree_add_12_51_groupi_n_2272);
  not csa_tree_add_12_51_groupi_drc_bufs23160(csa_tree_add_12_51_groupi_n_1740 ,csa_tree_add_12_51_groupi_n_1738);
  not csa_tree_add_12_51_groupi_drc_bufs23161(csa_tree_add_12_51_groupi_n_1739 ,csa_tree_add_12_51_groupi_n_1738);
  not csa_tree_add_12_51_groupi_drc_bufs23162(csa_tree_add_12_51_groupi_n_1738 ,csa_tree_add_12_51_groupi_n_2265);
  not csa_tree_add_12_51_groupi_drc_bufs23164(csa_tree_add_12_51_groupi_n_1737 ,csa_tree_add_12_51_groupi_n_1735);
  not csa_tree_add_12_51_groupi_drc_bufs23165(csa_tree_add_12_51_groupi_n_1736 ,csa_tree_add_12_51_groupi_n_1735);
  not csa_tree_add_12_51_groupi_drc_bufs23166(csa_tree_add_12_51_groupi_n_1735 ,csa_tree_add_12_51_groupi_n_2264);
  not csa_tree_add_12_51_groupi_drc_bufs23168(csa_tree_add_12_51_groupi_n_1734 ,csa_tree_add_12_51_groupi_n_1732);
  not csa_tree_add_12_51_groupi_drc_bufs23169(csa_tree_add_12_51_groupi_n_1733 ,csa_tree_add_12_51_groupi_n_1732);
  not csa_tree_add_12_51_groupi_drc_bufs23170(csa_tree_add_12_51_groupi_n_1732 ,csa_tree_add_12_51_groupi_n_2263);
  not csa_tree_add_12_51_groupi_drc_bufs23172(csa_tree_add_12_51_groupi_n_1731 ,csa_tree_add_12_51_groupi_n_1729);
  not csa_tree_add_12_51_groupi_drc_bufs23173(csa_tree_add_12_51_groupi_n_1730 ,csa_tree_add_12_51_groupi_n_1729);
  not csa_tree_add_12_51_groupi_drc_bufs23174(csa_tree_add_12_51_groupi_n_1729 ,csa_tree_add_12_51_groupi_n_2256);
  not csa_tree_add_12_51_groupi_drc_bufs23176(csa_tree_add_12_51_groupi_n_1728 ,csa_tree_add_12_51_groupi_n_1726);
  not csa_tree_add_12_51_groupi_drc_bufs23177(csa_tree_add_12_51_groupi_n_1727 ,csa_tree_add_12_51_groupi_n_1726);
  not csa_tree_add_12_51_groupi_drc_bufs23178(csa_tree_add_12_51_groupi_n_1726 ,csa_tree_add_12_51_groupi_n_2255);
  not csa_tree_add_12_51_groupi_drc_bufs23180(csa_tree_add_12_51_groupi_n_1725 ,csa_tree_add_12_51_groupi_n_1723);
  not csa_tree_add_12_51_groupi_drc_bufs23181(csa_tree_add_12_51_groupi_n_1724 ,csa_tree_add_12_51_groupi_n_1723);
  not csa_tree_add_12_51_groupi_drc_bufs23182(csa_tree_add_12_51_groupi_n_1723 ,csa_tree_add_12_51_groupi_n_2254);
  not csa_tree_add_12_51_groupi_drc_bufs23184(csa_tree_add_12_51_groupi_n_1722 ,csa_tree_add_12_51_groupi_n_1720);
  not csa_tree_add_12_51_groupi_drc_bufs23185(csa_tree_add_12_51_groupi_n_1721 ,csa_tree_add_12_51_groupi_n_1720);
  not csa_tree_add_12_51_groupi_drc_bufs23186(csa_tree_add_12_51_groupi_n_1720 ,csa_tree_add_12_51_groupi_n_2274);
  not csa_tree_add_12_51_groupi_drc_bufs23188(csa_tree_add_12_51_groupi_n_1719 ,csa_tree_add_12_51_groupi_n_1717);
  not csa_tree_add_12_51_groupi_drc_bufs23189(csa_tree_add_12_51_groupi_n_1718 ,csa_tree_add_12_51_groupi_n_1717);
  not csa_tree_add_12_51_groupi_drc_bufs23190(csa_tree_add_12_51_groupi_n_1717 ,csa_tree_add_12_51_groupi_n_2247);
  not csa_tree_add_12_51_groupi_drc_bufs23192(csa_tree_add_12_51_groupi_n_1716 ,csa_tree_add_12_51_groupi_n_1714);
  not csa_tree_add_12_51_groupi_drc_bufs23193(csa_tree_add_12_51_groupi_n_1715 ,csa_tree_add_12_51_groupi_n_1714);
  not csa_tree_add_12_51_groupi_drc_bufs23194(csa_tree_add_12_51_groupi_n_1714 ,csa_tree_add_12_51_groupi_n_2246);
  not csa_tree_add_12_51_groupi_drc_bufs23196(csa_tree_add_12_51_groupi_n_1713 ,csa_tree_add_12_51_groupi_n_1711);
  not csa_tree_add_12_51_groupi_drc_bufs23197(csa_tree_add_12_51_groupi_n_1712 ,csa_tree_add_12_51_groupi_n_1711);
  not csa_tree_add_12_51_groupi_drc_bufs23198(csa_tree_add_12_51_groupi_n_1711 ,csa_tree_add_12_51_groupi_n_2245);
  not csa_tree_add_12_51_groupi_drc_bufs23200(csa_tree_add_12_51_groupi_n_1710 ,csa_tree_add_12_51_groupi_n_1708);
  not csa_tree_add_12_51_groupi_drc_bufs23201(csa_tree_add_12_51_groupi_n_1709 ,csa_tree_add_12_51_groupi_n_1708);
  not csa_tree_add_12_51_groupi_drc_bufs23202(csa_tree_add_12_51_groupi_n_1708 ,csa_tree_add_12_51_groupi_n_2237);
  not csa_tree_add_12_51_groupi_drc_bufs23204(csa_tree_add_12_51_groupi_n_1707 ,csa_tree_add_12_51_groupi_n_1705);
  not csa_tree_add_12_51_groupi_drc_bufs23205(csa_tree_add_12_51_groupi_n_1706 ,csa_tree_add_12_51_groupi_n_1705);
  not csa_tree_add_12_51_groupi_drc_bufs23206(csa_tree_add_12_51_groupi_n_1705 ,csa_tree_add_12_51_groupi_n_2236);
  not csa_tree_add_12_51_groupi_drc_bufs23208(csa_tree_add_12_51_groupi_n_1704 ,csa_tree_add_12_51_groupi_n_1702);
  not csa_tree_add_12_51_groupi_drc_bufs23209(csa_tree_add_12_51_groupi_n_1703 ,csa_tree_add_12_51_groupi_n_1702);
  not csa_tree_add_12_51_groupi_drc_bufs23210(csa_tree_add_12_51_groupi_n_1702 ,csa_tree_add_12_51_groupi_n_2238);
  not csa_tree_add_12_51_groupi_drc_bufs23212(csa_tree_add_12_51_groupi_n_1701 ,csa_tree_add_12_51_groupi_n_1699);
  not csa_tree_add_12_51_groupi_drc_bufs23213(csa_tree_add_12_51_groupi_n_1700 ,csa_tree_add_12_51_groupi_n_1699);
  not csa_tree_add_12_51_groupi_drc_bufs23214(csa_tree_add_12_51_groupi_n_1699 ,csa_tree_add_12_51_groupi_n_2229);
  not csa_tree_add_12_51_groupi_drc_bufs23216(csa_tree_add_12_51_groupi_n_1698 ,csa_tree_add_12_51_groupi_n_1696);
  not csa_tree_add_12_51_groupi_drc_bufs23217(csa_tree_add_12_51_groupi_n_1697 ,csa_tree_add_12_51_groupi_n_1696);
  not csa_tree_add_12_51_groupi_drc_bufs23218(csa_tree_add_12_51_groupi_n_1696 ,csa_tree_add_12_51_groupi_n_2228);
  not csa_tree_add_12_51_groupi_drc_bufs23220(csa_tree_add_12_51_groupi_n_1695 ,csa_tree_add_12_51_groupi_n_1693);
  not csa_tree_add_12_51_groupi_drc_bufs23221(csa_tree_add_12_51_groupi_n_1694 ,csa_tree_add_12_51_groupi_n_1693);
  not csa_tree_add_12_51_groupi_drc_bufs23222(csa_tree_add_12_51_groupi_n_1693 ,csa_tree_add_12_51_groupi_n_2227);
  not csa_tree_add_12_51_groupi_drc_bufs23224(csa_tree_add_12_51_groupi_n_1692 ,csa_tree_add_12_51_groupi_n_1690);
  not csa_tree_add_12_51_groupi_drc_bufs23225(csa_tree_add_12_51_groupi_n_1691 ,csa_tree_add_12_51_groupi_n_1690);
  not csa_tree_add_12_51_groupi_drc_bufs23226(csa_tree_add_12_51_groupi_n_1690 ,csa_tree_add_12_51_groupi_n_2220);
  not csa_tree_add_12_51_groupi_drc_bufs23228(csa_tree_add_12_51_groupi_n_1689 ,csa_tree_add_12_51_groupi_n_1687);
  not csa_tree_add_12_51_groupi_drc_bufs23229(csa_tree_add_12_51_groupi_n_1688 ,csa_tree_add_12_51_groupi_n_1687);
  not csa_tree_add_12_51_groupi_drc_bufs23230(csa_tree_add_12_51_groupi_n_1687 ,csa_tree_add_12_51_groupi_n_2148);
  not csa_tree_add_12_51_groupi_drc_bufs23232(csa_tree_add_12_51_groupi_n_1686 ,csa_tree_add_12_51_groupi_n_1684);
  not csa_tree_add_12_51_groupi_drc_bufs23233(csa_tree_add_12_51_groupi_n_1685 ,csa_tree_add_12_51_groupi_n_1684);
  not csa_tree_add_12_51_groupi_drc_bufs23234(csa_tree_add_12_51_groupi_n_1684 ,csa_tree_add_12_51_groupi_n_2926);
  not csa_tree_add_12_51_groupi_drc_bufs23236(csa_tree_add_12_51_groupi_n_1683 ,csa_tree_add_12_51_groupi_n_1681);
  not csa_tree_add_12_51_groupi_drc_bufs23237(csa_tree_add_12_51_groupi_n_1682 ,csa_tree_add_12_51_groupi_n_1681);
  not csa_tree_add_12_51_groupi_drc_bufs23238(csa_tree_add_12_51_groupi_n_1681 ,csa_tree_add_12_51_groupi_n_2504);
  not csa_tree_add_12_51_groupi_drc_bufs23240(csa_tree_add_12_51_groupi_n_1680 ,csa_tree_add_12_51_groupi_n_1678);
  not csa_tree_add_12_51_groupi_drc_bufs23241(csa_tree_add_12_51_groupi_n_1679 ,csa_tree_add_12_51_groupi_n_1678);
  not csa_tree_add_12_51_groupi_drc_bufs23242(csa_tree_add_12_51_groupi_n_1678 ,csa_tree_add_12_51_groupi_n_2914);
  not csa_tree_add_12_51_groupi_drc_bufs23244(csa_tree_add_12_51_groupi_n_1677 ,csa_tree_add_12_51_groupi_n_1675);
  not csa_tree_add_12_51_groupi_drc_bufs23245(csa_tree_add_12_51_groupi_n_1676 ,csa_tree_add_12_51_groupi_n_1675);
  not csa_tree_add_12_51_groupi_drc_bufs23246(csa_tree_add_12_51_groupi_n_1675 ,csa_tree_add_12_51_groupi_n_2504);
  not csa_tree_add_12_51_groupi_drc_bufs23248(csa_tree_add_12_51_groupi_n_1674 ,csa_tree_add_12_51_groupi_n_1672);
  not csa_tree_add_12_51_groupi_drc_bufs23249(csa_tree_add_12_51_groupi_n_1673 ,csa_tree_add_12_51_groupi_n_1672);
  not csa_tree_add_12_51_groupi_drc_bufs23250(csa_tree_add_12_51_groupi_n_1672 ,csa_tree_add_12_51_groupi_n_2940);
  not csa_tree_add_12_51_groupi_drc_bufs23252(csa_tree_add_12_51_groupi_n_1671 ,csa_tree_add_12_51_groupi_n_1669);
  not csa_tree_add_12_51_groupi_drc_bufs23253(csa_tree_add_12_51_groupi_n_1670 ,csa_tree_add_12_51_groupi_n_1669);
  not csa_tree_add_12_51_groupi_drc_bufs23254(csa_tree_add_12_51_groupi_n_1669 ,csa_tree_add_12_51_groupi_n_2145);
  not csa_tree_add_12_51_groupi_drc_bufs23256(csa_tree_add_12_51_groupi_n_1668 ,csa_tree_add_12_51_groupi_n_1666);
  not csa_tree_add_12_51_groupi_drc_bufs23257(csa_tree_add_12_51_groupi_n_1667 ,csa_tree_add_12_51_groupi_n_1666);
  not csa_tree_add_12_51_groupi_drc_bufs23258(csa_tree_add_12_51_groupi_n_1666 ,csa_tree_add_12_51_groupi_n_2935);
  not csa_tree_add_12_51_groupi_drc_bufs23260(csa_tree_add_12_51_groupi_n_1665 ,csa_tree_add_12_51_groupi_n_1663);
  not csa_tree_add_12_51_groupi_drc_bufs23261(csa_tree_add_12_51_groupi_n_1664 ,csa_tree_add_12_51_groupi_n_1663);
  not csa_tree_add_12_51_groupi_drc_bufs23262(csa_tree_add_12_51_groupi_n_1663 ,csa_tree_add_12_51_groupi_n_2918);
  not csa_tree_add_12_51_groupi_drc_bufs23264(csa_tree_add_12_51_groupi_n_1662 ,csa_tree_add_12_51_groupi_n_1660);
  not csa_tree_add_12_51_groupi_drc_bufs23265(csa_tree_add_12_51_groupi_n_1661 ,csa_tree_add_12_51_groupi_n_1660);
  not csa_tree_add_12_51_groupi_drc_bufs23266(csa_tree_add_12_51_groupi_n_1660 ,csa_tree_add_12_51_groupi_n_2936);
  not csa_tree_add_12_51_groupi_drc_bufs23268(csa_tree_add_12_51_groupi_n_1659 ,csa_tree_add_12_51_groupi_n_1657);
  not csa_tree_add_12_51_groupi_drc_bufs23269(csa_tree_add_12_51_groupi_n_1658 ,csa_tree_add_12_51_groupi_n_1657);
  not csa_tree_add_12_51_groupi_drc_bufs23270(csa_tree_add_12_51_groupi_n_1657 ,csa_tree_add_12_51_groupi_n_2142);
  not csa_tree_add_12_51_groupi_drc_bufs23272(csa_tree_add_12_51_groupi_n_1656 ,csa_tree_add_12_51_groupi_n_1654);
  not csa_tree_add_12_51_groupi_drc_bufs23273(csa_tree_add_12_51_groupi_n_1655 ,csa_tree_add_12_51_groupi_n_1654);
  not csa_tree_add_12_51_groupi_drc_bufs23274(csa_tree_add_12_51_groupi_n_1654 ,csa_tree_add_12_51_groupi_n_2913);
  not csa_tree_add_12_51_groupi_drc_bufs23276(csa_tree_add_12_51_groupi_n_1653 ,csa_tree_add_12_51_groupi_n_1651);
  not csa_tree_add_12_51_groupi_drc_bufs23277(csa_tree_add_12_51_groupi_n_1652 ,csa_tree_add_12_51_groupi_n_1651);
  not csa_tree_add_12_51_groupi_drc_bufs23278(csa_tree_add_12_51_groupi_n_1651 ,csa_tree_add_12_51_groupi_n_2505);
  not csa_tree_add_12_51_groupi_drc_bufs23280(csa_tree_add_12_51_groupi_n_1650 ,csa_tree_add_12_51_groupi_n_1648);
  not csa_tree_add_12_51_groupi_drc_bufs23281(csa_tree_add_12_51_groupi_n_1649 ,csa_tree_add_12_51_groupi_n_1648);
  not csa_tree_add_12_51_groupi_drc_bufs23282(csa_tree_add_12_51_groupi_n_1648 ,csa_tree_add_12_51_groupi_n_2139);
  not csa_tree_add_12_51_groupi_drc_bufs23284(csa_tree_add_12_51_groupi_n_1647 ,csa_tree_add_12_51_groupi_n_1645);
  not csa_tree_add_12_51_groupi_drc_bufs23285(csa_tree_add_12_51_groupi_n_1646 ,csa_tree_add_12_51_groupi_n_1645);
  not csa_tree_add_12_51_groupi_drc_bufs23286(csa_tree_add_12_51_groupi_n_1645 ,csa_tree_add_12_51_groupi_n_2920);
  not csa_tree_add_12_51_groupi_drc_bufs23288(csa_tree_add_12_51_groupi_n_1644 ,csa_tree_add_12_51_groupi_n_1642);
  not csa_tree_add_12_51_groupi_drc_bufs23289(csa_tree_add_12_51_groupi_n_1643 ,csa_tree_add_12_51_groupi_n_1642);
  not csa_tree_add_12_51_groupi_drc_bufs23290(csa_tree_add_12_51_groupi_n_1642 ,csa_tree_add_12_51_groupi_n_2136);
  not csa_tree_add_12_51_groupi_drc_bufs23292(csa_tree_add_12_51_groupi_n_1641 ,csa_tree_add_12_51_groupi_n_1639);
  not csa_tree_add_12_51_groupi_drc_bufs23293(csa_tree_add_12_51_groupi_n_1640 ,csa_tree_add_12_51_groupi_n_1639);
  not csa_tree_add_12_51_groupi_drc_bufs23294(csa_tree_add_12_51_groupi_n_1639 ,csa_tree_add_12_51_groupi_n_2912);
  not csa_tree_add_12_51_groupi_drc_bufs23296(csa_tree_add_12_51_groupi_n_1638 ,csa_tree_add_12_51_groupi_n_1636);
  not csa_tree_add_12_51_groupi_drc_bufs23297(csa_tree_add_12_51_groupi_n_1637 ,csa_tree_add_12_51_groupi_n_1636);
  not csa_tree_add_12_51_groupi_drc_bufs23298(csa_tree_add_12_51_groupi_n_1636 ,csa_tree_add_12_51_groupi_n_2133);
  not csa_tree_add_12_51_groupi_drc_bufs23300(csa_tree_add_12_51_groupi_n_1635 ,csa_tree_add_12_51_groupi_n_1633);
  not csa_tree_add_12_51_groupi_drc_bufs23301(csa_tree_add_12_51_groupi_n_1634 ,csa_tree_add_12_51_groupi_n_1633);
  not csa_tree_add_12_51_groupi_drc_bufs23302(csa_tree_add_12_51_groupi_n_1633 ,csa_tree_add_12_51_groupi_n_2917);
  not csa_tree_add_12_51_groupi_drc_bufs23304(csa_tree_add_12_51_groupi_n_1632 ,csa_tree_add_12_51_groupi_n_1630);
  not csa_tree_add_12_51_groupi_drc_bufs23305(csa_tree_add_12_51_groupi_n_1631 ,csa_tree_add_12_51_groupi_n_1630);
  not csa_tree_add_12_51_groupi_drc_bufs23306(csa_tree_add_12_51_groupi_n_1630 ,csa_tree_add_12_51_groupi_n_2130);
  not csa_tree_add_12_51_groupi_drc_bufs23308(csa_tree_add_12_51_groupi_n_1629 ,csa_tree_add_12_51_groupi_n_1627);
  not csa_tree_add_12_51_groupi_drc_bufs23309(csa_tree_add_12_51_groupi_n_1628 ,csa_tree_add_12_51_groupi_n_1627);
  not csa_tree_add_12_51_groupi_drc_bufs23310(csa_tree_add_12_51_groupi_n_1627 ,csa_tree_add_12_51_groupi_n_2911);
  not csa_tree_add_12_51_groupi_drc_bufs23312(csa_tree_add_12_51_groupi_n_1626 ,csa_tree_add_12_51_groupi_n_1624);
  not csa_tree_add_12_51_groupi_drc_bufs23313(csa_tree_add_12_51_groupi_n_1625 ,csa_tree_add_12_51_groupi_n_1624);
  not csa_tree_add_12_51_groupi_drc_bufs23314(csa_tree_add_12_51_groupi_n_1624 ,csa_tree_add_12_51_groupi_n_2127);
  not csa_tree_add_12_51_groupi_drc_bufs23316(csa_tree_add_12_51_groupi_n_1623 ,csa_tree_add_12_51_groupi_n_1621);
  not csa_tree_add_12_51_groupi_drc_bufs23317(csa_tree_add_12_51_groupi_n_1622 ,csa_tree_add_12_51_groupi_n_1621);
  not csa_tree_add_12_51_groupi_drc_bufs23318(csa_tree_add_12_51_groupi_n_1621 ,csa_tree_add_12_51_groupi_n_2921);
  not csa_tree_add_12_51_groupi_drc_bufs23320(csa_tree_add_12_51_groupi_n_1620 ,csa_tree_add_12_51_groupi_n_1618);
  not csa_tree_add_12_51_groupi_drc_bufs23321(csa_tree_add_12_51_groupi_n_1619 ,csa_tree_add_12_51_groupi_n_1618);
  not csa_tree_add_12_51_groupi_drc_bufs23322(csa_tree_add_12_51_groupi_n_1618 ,csa_tree_add_12_51_groupi_n_2124);
  not csa_tree_add_12_51_groupi_drc_bufs23324(csa_tree_add_12_51_groupi_n_1617 ,csa_tree_add_12_51_groupi_n_1615);
  not csa_tree_add_12_51_groupi_drc_bufs23325(csa_tree_add_12_51_groupi_n_1616 ,csa_tree_add_12_51_groupi_n_1615);
  not csa_tree_add_12_51_groupi_drc_bufs23326(csa_tree_add_12_51_groupi_n_1615 ,csa_tree_add_12_51_groupi_n_2910);
  not csa_tree_add_12_51_groupi_drc_bufs23328(csa_tree_add_12_51_groupi_n_1614 ,csa_tree_add_12_51_groupi_n_1612);
  not csa_tree_add_12_51_groupi_drc_bufs23329(csa_tree_add_12_51_groupi_n_1613 ,csa_tree_add_12_51_groupi_n_1612);
  not csa_tree_add_12_51_groupi_drc_bufs23330(csa_tree_add_12_51_groupi_n_1612 ,csa_tree_add_12_51_groupi_n_2121);
  not csa_tree_add_12_51_groupi_drc_bufs23332(csa_tree_add_12_51_groupi_n_1611 ,csa_tree_add_12_51_groupi_n_1609);
  not csa_tree_add_12_51_groupi_drc_bufs23333(csa_tree_add_12_51_groupi_n_1610 ,csa_tree_add_12_51_groupi_n_1609);
  not csa_tree_add_12_51_groupi_drc_bufs23334(csa_tree_add_12_51_groupi_n_1609 ,csa_tree_add_12_51_groupi_n_2916);
  not csa_tree_add_12_51_groupi_drc_bufs23336(csa_tree_add_12_51_groupi_n_1608 ,csa_tree_add_12_51_groupi_n_1606);
  not csa_tree_add_12_51_groupi_drc_bufs23337(csa_tree_add_12_51_groupi_n_1607 ,csa_tree_add_12_51_groupi_n_1606);
  not csa_tree_add_12_51_groupi_drc_bufs23338(csa_tree_add_12_51_groupi_n_1606 ,csa_tree_add_12_51_groupi_n_2118);
  not csa_tree_add_12_51_groupi_drc_bufs23340(csa_tree_add_12_51_groupi_n_1605 ,csa_tree_add_12_51_groupi_n_1603);
  not csa_tree_add_12_51_groupi_drc_bufs23341(csa_tree_add_12_51_groupi_n_1604 ,csa_tree_add_12_51_groupi_n_1603);
  not csa_tree_add_12_51_groupi_drc_bufs23342(csa_tree_add_12_51_groupi_n_1603 ,csa_tree_add_12_51_groupi_n_2909);
  not csa_tree_add_12_51_groupi_drc_bufs23344(csa_tree_add_12_51_groupi_n_1602 ,csa_tree_add_12_51_groupi_n_1600);
  not csa_tree_add_12_51_groupi_drc_bufs23345(csa_tree_add_12_51_groupi_n_1601 ,csa_tree_add_12_51_groupi_n_1600);
  not csa_tree_add_12_51_groupi_drc_bufs23346(csa_tree_add_12_51_groupi_n_1600 ,csa_tree_add_12_51_groupi_n_2115);
  not csa_tree_add_12_51_groupi_drc_bufs23348(csa_tree_add_12_51_groupi_n_1599 ,csa_tree_add_12_51_groupi_n_1597);
  not csa_tree_add_12_51_groupi_drc_bufs23349(csa_tree_add_12_51_groupi_n_1598 ,csa_tree_add_12_51_groupi_n_1597);
  not csa_tree_add_12_51_groupi_drc_bufs23350(csa_tree_add_12_51_groupi_n_1597 ,csa_tree_add_12_51_groupi_n_2919);
  not csa_tree_add_12_51_groupi_drc_bufs23352(csa_tree_add_12_51_groupi_n_1596 ,csa_tree_add_12_51_groupi_n_1594);
  not csa_tree_add_12_51_groupi_drc_bufs23353(csa_tree_add_12_51_groupi_n_1595 ,csa_tree_add_12_51_groupi_n_1594);
  not csa_tree_add_12_51_groupi_drc_bufs23354(csa_tree_add_12_51_groupi_n_1594 ,csa_tree_add_12_51_groupi_n_2112);
  not csa_tree_add_12_51_groupi_drc_bufs23356(csa_tree_add_12_51_groupi_n_1593 ,csa_tree_add_12_51_groupi_n_1591);
  not csa_tree_add_12_51_groupi_drc_bufs23357(csa_tree_add_12_51_groupi_n_1592 ,csa_tree_add_12_51_groupi_n_1591);
  not csa_tree_add_12_51_groupi_drc_bufs23358(csa_tree_add_12_51_groupi_n_1591 ,csa_tree_add_12_51_groupi_n_2908);
  not csa_tree_add_12_51_groupi_drc_bufs23360(csa_tree_add_12_51_groupi_n_1590 ,csa_tree_add_12_51_groupi_n_1588);
  not csa_tree_add_12_51_groupi_drc_bufs23361(csa_tree_add_12_51_groupi_n_1589 ,csa_tree_add_12_51_groupi_n_1588);
  not csa_tree_add_12_51_groupi_drc_bufs23362(csa_tree_add_12_51_groupi_n_1588 ,csa_tree_add_12_51_groupi_n_2109);
  not csa_tree_add_12_51_groupi_drc_bufs23364(csa_tree_add_12_51_groupi_n_1587 ,csa_tree_add_12_51_groupi_n_1585);
  not csa_tree_add_12_51_groupi_drc_bufs23365(csa_tree_add_12_51_groupi_n_1586 ,csa_tree_add_12_51_groupi_n_1585);
  not csa_tree_add_12_51_groupi_drc_bufs23366(csa_tree_add_12_51_groupi_n_1585 ,csa_tree_add_12_51_groupi_n_2915);
  not csa_tree_add_12_51_groupi_drc_bufs23368(csa_tree_add_12_51_groupi_n_1584 ,csa_tree_add_12_51_groupi_n_1582);
  not csa_tree_add_12_51_groupi_drc_bufs23369(csa_tree_add_12_51_groupi_n_1583 ,csa_tree_add_12_51_groupi_n_1582);
  not csa_tree_add_12_51_groupi_drc_bufs23370(csa_tree_add_12_51_groupi_n_1582 ,csa_tree_add_12_51_groupi_n_2907);
  not csa_tree_add_12_51_groupi_drc_bufs23372(csa_tree_add_12_51_groupi_n_1581 ,csa_tree_add_12_51_groupi_n_1579);
  not csa_tree_add_12_51_groupi_drc_bufs23373(csa_tree_add_12_51_groupi_n_1580 ,csa_tree_add_12_51_groupi_n_1579);
  not csa_tree_add_12_51_groupi_drc_bufs23374(csa_tree_add_12_51_groupi_n_1579 ,csa_tree_add_12_51_groupi_n_2106);
  not csa_tree_add_12_51_groupi_drc_bufs23376(csa_tree_add_12_51_groupi_n_1578 ,csa_tree_add_12_51_groupi_n_1576);
  not csa_tree_add_12_51_groupi_drc_bufs23377(csa_tree_add_12_51_groupi_n_1577 ,csa_tree_add_12_51_groupi_n_1576);
  not csa_tree_add_12_51_groupi_drc_bufs23378(csa_tree_add_12_51_groupi_n_1576 ,csa_tree_add_12_51_groupi_n_2463);
  not csa_tree_add_12_51_groupi_drc_bufs23380(csa_tree_add_12_51_groupi_n_1575 ,csa_tree_add_12_51_groupi_n_1573);
  not csa_tree_add_12_51_groupi_drc_bufs23381(csa_tree_add_12_51_groupi_n_1574 ,csa_tree_add_12_51_groupi_n_1573);
  not csa_tree_add_12_51_groupi_drc_bufs23382(csa_tree_add_12_51_groupi_n_1573 ,csa_tree_add_12_51_groupi_n_2926);
  not csa_tree_add_12_51_groupi_drc_bufs23384(csa_tree_add_12_51_groupi_n_1572 ,csa_tree_add_12_51_groupi_n_1570);
  not csa_tree_add_12_51_groupi_drc_bufs23385(csa_tree_add_12_51_groupi_n_1571 ,csa_tree_add_12_51_groupi_n_1570);
  not csa_tree_add_12_51_groupi_drc_bufs23386(csa_tree_add_12_51_groupi_n_1570 ,csa_tree_add_12_51_groupi_n_2335);
  not csa_tree_add_12_51_groupi_drc_bufs23388(csa_tree_add_12_51_groupi_n_1569 ,csa_tree_add_12_51_groupi_n_1567);
  not csa_tree_add_12_51_groupi_drc_bufs23389(csa_tree_add_12_51_groupi_n_1568 ,csa_tree_add_12_51_groupi_n_1567);
  not csa_tree_add_12_51_groupi_drc_bufs23390(csa_tree_add_12_51_groupi_n_1567 ,csa_tree_add_12_51_groupi_n_2299);
  not csa_tree_add_12_51_groupi_drc_bufs23392(csa_tree_add_12_51_groupi_n_1566 ,csa_tree_add_12_51_groupi_n_1564);
  not csa_tree_add_12_51_groupi_drc_bufs23393(csa_tree_add_12_51_groupi_n_1565 ,csa_tree_add_12_51_groupi_n_1564);
  not csa_tree_add_12_51_groupi_drc_bufs23394(csa_tree_add_12_51_groupi_n_1564 ,csa_tree_add_12_51_groupi_n_2290);
  not csa_tree_add_12_51_groupi_drc_bufs23396(csa_tree_add_12_51_groupi_n_1563 ,csa_tree_add_12_51_groupi_n_1561);
  not csa_tree_add_12_51_groupi_drc_bufs23397(csa_tree_add_12_51_groupi_n_1562 ,csa_tree_add_12_51_groupi_n_1561);
  not csa_tree_add_12_51_groupi_drc_bufs23398(csa_tree_add_12_51_groupi_n_1561 ,csa_tree_add_12_51_groupi_n_2940);
  not csa_tree_add_12_51_groupi_drc_bufs23400(csa_tree_add_12_51_groupi_n_1560 ,csa_tree_add_12_51_groupi_n_1558);
  not csa_tree_add_12_51_groupi_drc_bufs23401(csa_tree_add_12_51_groupi_n_1559 ,csa_tree_add_12_51_groupi_n_1558);
  not csa_tree_add_12_51_groupi_drc_bufs23402(csa_tree_add_12_51_groupi_n_1558 ,csa_tree_add_12_51_groupi_n_2935);
  not csa_tree_add_12_51_groupi_drc_bufs23404(csa_tree_add_12_51_groupi_n_1557 ,csa_tree_add_12_51_groupi_n_1555);
  not csa_tree_add_12_51_groupi_drc_bufs23405(csa_tree_add_12_51_groupi_n_1556 ,csa_tree_add_12_51_groupi_n_1555);
  not csa_tree_add_12_51_groupi_drc_bufs23406(csa_tree_add_12_51_groupi_n_1555 ,csa_tree_add_12_51_groupi_n_2936);
  not csa_tree_add_12_51_groupi_drc_bufs23408(csa_tree_add_12_51_groupi_n_1554 ,csa_tree_add_12_51_groupi_n_1552);
  not csa_tree_add_12_51_groupi_drc_bufs23409(csa_tree_add_12_51_groupi_n_1553 ,csa_tree_add_12_51_groupi_n_1552);
  not csa_tree_add_12_51_groupi_drc_bufs23410(csa_tree_add_12_51_groupi_n_1552 ,csa_tree_add_12_51_groupi_n_2930);
  not csa_tree_add_12_51_groupi_drc_bufs23412(csa_tree_add_12_51_groupi_n_1551 ,csa_tree_add_12_51_groupi_n_1549);
  not csa_tree_add_12_51_groupi_drc_bufs23413(csa_tree_add_12_51_groupi_n_1550 ,csa_tree_add_12_51_groupi_n_1549);
  not csa_tree_add_12_51_groupi_drc_bufs23414(csa_tree_add_12_51_groupi_n_1549 ,csa_tree_add_12_51_groupi_n_3507);
  not csa_tree_add_12_51_groupi_drc_bufs23416(csa_tree_add_12_51_groupi_n_1548 ,csa_tree_add_12_51_groupi_n_1546);
  not csa_tree_add_12_51_groupi_drc_bufs23417(csa_tree_add_12_51_groupi_n_1547 ,csa_tree_add_12_51_groupi_n_1546);
  not csa_tree_add_12_51_groupi_drc_bufs23418(csa_tree_add_12_51_groupi_n_1546 ,csa_tree_add_12_51_groupi_n_2930);
  not csa_tree_add_12_51_groupi_drc_bufs23420(csa_tree_add_12_51_groupi_n_1545 ,csa_tree_add_12_51_groupi_n_1543);
  not csa_tree_add_12_51_groupi_drc_bufs23421(csa_tree_add_12_51_groupi_n_1544 ,csa_tree_add_12_51_groupi_n_1543);
  not csa_tree_add_12_51_groupi_drc_bufs23422(csa_tree_add_12_51_groupi_n_1543 ,csa_tree_add_12_51_groupi_n_2937);
  not csa_tree_add_12_51_groupi_drc_bufs23424(csa_tree_add_12_51_groupi_n_1542 ,csa_tree_add_12_51_groupi_n_1540);
  not csa_tree_add_12_51_groupi_drc_bufs23425(csa_tree_add_12_51_groupi_n_1541 ,csa_tree_add_12_51_groupi_n_1540);
  not csa_tree_add_12_51_groupi_drc_bufs23426(csa_tree_add_12_51_groupi_n_1540 ,csa_tree_add_12_51_groupi_n_2937);
  not csa_tree_add_12_51_groupi_drc_bufs23428(csa_tree_add_12_51_groupi_n_1539 ,csa_tree_add_12_51_groupi_n_1537);
  not csa_tree_add_12_51_groupi_drc_bufs23429(csa_tree_add_12_51_groupi_n_1538 ,csa_tree_add_12_51_groupi_n_1537);
  not csa_tree_add_12_51_groupi_drc_bufs23430(csa_tree_add_12_51_groupi_n_1537 ,csa_tree_add_12_51_groupi_n_2939);
  not csa_tree_add_12_51_groupi_drc_bufs23432(csa_tree_add_12_51_groupi_n_1536 ,csa_tree_add_12_51_groupi_n_1534);
  not csa_tree_add_12_51_groupi_drc_bufs23433(csa_tree_add_12_51_groupi_n_1535 ,csa_tree_add_12_51_groupi_n_1534);
  not csa_tree_add_12_51_groupi_drc_bufs23434(csa_tree_add_12_51_groupi_n_1534 ,csa_tree_add_12_51_groupi_n_2939);
  not csa_tree_add_12_51_groupi_drc_bufs23436(csa_tree_add_12_51_groupi_n_1533 ,csa_tree_add_12_51_groupi_n_1531);
  not csa_tree_add_12_51_groupi_drc_bufs23437(csa_tree_add_12_51_groupi_n_1532 ,csa_tree_add_12_51_groupi_n_1531);
  not csa_tree_add_12_51_groupi_drc_bufs23438(csa_tree_add_12_51_groupi_n_1531 ,csa_tree_add_12_51_groupi_n_2104);
  not csa_tree_add_12_51_groupi_drc_bufs23440(csa_tree_add_12_51_groupi_n_1530 ,csa_tree_add_12_51_groupi_n_1528);
  not csa_tree_add_12_51_groupi_drc_bufs23441(csa_tree_add_12_51_groupi_n_1529 ,csa_tree_add_12_51_groupi_n_1528);
  not csa_tree_add_12_51_groupi_drc_bufs23442(csa_tree_add_12_51_groupi_n_1528 ,csa_tree_add_12_51_groupi_n_2104);
  not csa_tree_add_12_51_groupi_drc_bufs23444(csa_tree_add_12_51_groupi_n_1527 ,csa_tree_add_12_51_groupi_n_1525);
  not csa_tree_add_12_51_groupi_drc_bufs23445(csa_tree_add_12_51_groupi_n_1526 ,csa_tree_add_12_51_groupi_n_1525);
  not csa_tree_add_12_51_groupi_drc_bufs23446(csa_tree_add_12_51_groupi_n_1525 ,csa_tree_add_12_51_groupi_n_3501);
  not csa_tree_add_12_51_groupi_drc_bufs23448(csa_tree_add_12_51_groupi_n_1524 ,csa_tree_add_12_51_groupi_n_1522);
  not csa_tree_add_12_51_groupi_drc_bufs23449(csa_tree_add_12_51_groupi_n_1523 ,csa_tree_add_12_51_groupi_n_1522);
  not csa_tree_add_12_51_groupi_drc_bufs23450(csa_tree_add_12_51_groupi_n_1522 ,csa_tree_add_12_51_groupi_n_3501);
  not csa_tree_add_12_51_groupi_drc_bufs23452(csa_tree_add_12_51_groupi_n_1521 ,csa_tree_add_12_51_groupi_n_1519);
  not csa_tree_add_12_51_groupi_drc_bufs23453(csa_tree_add_12_51_groupi_n_1520 ,csa_tree_add_12_51_groupi_n_1519);
  not csa_tree_add_12_51_groupi_drc_bufs23454(csa_tree_add_12_51_groupi_n_1519 ,csa_tree_add_12_51_groupi_n_2923);
  not csa_tree_add_12_51_groupi_drc_bufs23456(csa_tree_add_12_51_groupi_n_1518 ,csa_tree_add_12_51_groupi_n_1516);
  not csa_tree_add_12_51_groupi_drc_bufs23457(csa_tree_add_12_51_groupi_n_1517 ,csa_tree_add_12_51_groupi_n_1516);
  not csa_tree_add_12_51_groupi_drc_bufs23458(csa_tree_add_12_51_groupi_n_1516 ,csa_tree_add_12_51_groupi_n_2754);
  not csa_tree_add_12_51_groupi_drc_bufs23460(csa_tree_add_12_51_groupi_n_1515 ,csa_tree_add_12_51_groupi_n_1513);
  not csa_tree_add_12_51_groupi_drc_bufs23461(csa_tree_add_12_51_groupi_n_1514 ,csa_tree_add_12_51_groupi_n_1513);
  not csa_tree_add_12_51_groupi_drc_bufs23462(csa_tree_add_12_51_groupi_n_1513 ,csa_tree_add_12_51_groupi_n_2948);
  not csa_tree_add_12_51_groupi_drc_bufs23464(csa_tree_add_12_51_groupi_n_1512 ,csa_tree_add_12_51_groupi_n_1510);
  not csa_tree_add_12_51_groupi_drc_bufs23465(csa_tree_add_12_51_groupi_n_1511 ,csa_tree_add_12_51_groupi_n_1510);
  not csa_tree_add_12_51_groupi_drc_bufs23466(csa_tree_add_12_51_groupi_n_1510 ,csa_tree_add_12_51_groupi_n_2943);
  not csa_tree_add_12_51_groupi_drc_bufs23468(csa_tree_add_12_51_groupi_n_1509 ,csa_tree_add_12_51_groupi_n_1507);
  not csa_tree_add_12_51_groupi_drc_bufs23469(csa_tree_add_12_51_groupi_n_1508 ,csa_tree_add_12_51_groupi_n_1507);
  not csa_tree_add_12_51_groupi_drc_bufs23470(csa_tree_add_12_51_groupi_n_1507 ,csa_tree_add_12_51_groupi_n_3506);
  not csa_tree_add_12_51_groupi_drc_bufs23472(csa_tree_add_12_51_groupi_n_1506 ,csa_tree_add_12_51_groupi_n_1504);
  not csa_tree_add_12_51_groupi_drc_bufs23473(csa_tree_add_12_51_groupi_n_1505 ,csa_tree_add_12_51_groupi_n_1504);
  not csa_tree_add_12_51_groupi_drc_bufs23474(csa_tree_add_12_51_groupi_n_1504 ,csa_tree_add_12_51_groupi_n_2927);
  not csa_tree_add_12_51_groupi_drc_bufs23476(csa_tree_add_12_51_groupi_n_1503 ,csa_tree_add_12_51_groupi_n_1501);
  not csa_tree_add_12_51_groupi_drc_bufs23477(csa_tree_add_12_51_groupi_n_1502 ,csa_tree_add_12_51_groupi_n_1501);
  not csa_tree_add_12_51_groupi_drc_bufs23478(csa_tree_add_12_51_groupi_n_1501 ,csa_tree_add_12_51_groupi_n_3497);
  not csa_tree_add_12_51_groupi_drc_bufs23480(csa_tree_add_12_51_groupi_n_1500 ,csa_tree_add_12_51_groupi_n_1498);
  not csa_tree_add_12_51_groupi_drc_bufs23481(csa_tree_add_12_51_groupi_n_1499 ,csa_tree_add_12_51_groupi_n_1498);
  not csa_tree_add_12_51_groupi_drc_bufs23482(csa_tree_add_12_51_groupi_n_1498 ,csa_tree_add_12_51_groupi_n_2102);
  not csa_tree_add_12_51_groupi_drc_bufs23484(csa_tree_add_12_51_groupi_n_1497 ,csa_tree_add_12_51_groupi_n_1495);
  not csa_tree_add_12_51_groupi_drc_bufs23485(csa_tree_add_12_51_groupi_n_1496 ,csa_tree_add_12_51_groupi_n_1495);
  not csa_tree_add_12_51_groupi_drc_bufs23486(csa_tree_add_12_51_groupi_n_1495 ,csa_tree_add_12_51_groupi_n_2098);
  not csa_tree_add_12_51_groupi_drc_bufs23488(csa_tree_add_12_51_groupi_n_1494 ,csa_tree_add_12_51_groupi_n_1492);
  not csa_tree_add_12_51_groupi_drc_bufs23489(csa_tree_add_12_51_groupi_n_1493 ,csa_tree_add_12_51_groupi_n_1492);
  not csa_tree_add_12_51_groupi_drc_bufs23490(csa_tree_add_12_51_groupi_n_1492 ,csa_tree_add_12_51_groupi_n_2941);
  not csa_tree_add_12_51_groupi_drc_bufs23492(csa_tree_add_12_51_groupi_n_1491 ,csa_tree_add_12_51_groupi_n_1489);
  not csa_tree_add_12_51_groupi_drc_bufs23493(csa_tree_add_12_51_groupi_n_1490 ,csa_tree_add_12_51_groupi_n_1489);
  not csa_tree_add_12_51_groupi_drc_bufs23494(csa_tree_add_12_51_groupi_n_1489 ,csa_tree_add_12_51_groupi_n_2094);
  not csa_tree_add_12_51_groupi_drc_bufs23496(csa_tree_add_12_51_groupi_n_1488 ,csa_tree_add_12_51_groupi_n_1486);
  not csa_tree_add_12_51_groupi_drc_bufs23497(csa_tree_add_12_51_groupi_n_1487 ,csa_tree_add_12_51_groupi_n_1486);
  not csa_tree_add_12_51_groupi_drc_bufs23498(csa_tree_add_12_51_groupi_n_1486 ,csa_tree_add_12_51_groupi_n_2932);
  not csa_tree_add_12_51_groupi_drc_bufs23500(csa_tree_add_12_51_groupi_n_1485 ,csa_tree_add_12_51_groupi_n_1483);
  not csa_tree_add_12_51_groupi_drc_bufs23501(csa_tree_add_12_51_groupi_n_1484 ,csa_tree_add_12_51_groupi_n_1483);
  not csa_tree_add_12_51_groupi_drc_bufs23502(csa_tree_add_12_51_groupi_n_1483 ,csa_tree_add_12_51_groupi_n_2092);
  not csa_tree_add_12_51_groupi_drc_bufs23504(csa_tree_add_12_51_groupi_n_1482 ,csa_tree_add_12_51_groupi_n_1480);
  not csa_tree_add_12_51_groupi_drc_bufs23505(csa_tree_add_12_51_groupi_n_1481 ,csa_tree_add_12_51_groupi_n_1480);
  not csa_tree_add_12_51_groupi_drc_bufs23506(csa_tree_add_12_51_groupi_n_1480 ,csa_tree_add_12_51_groupi_n_2938);
  not csa_tree_add_12_51_groupi_drc_bufs23508(csa_tree_add_12_51_groupi_n_1479 ,csa_tree_add_12_51_groupi_n_1477);
  not csa_tree_add_12_51_groupi_drc_bufs23509(csa_tree_add_12_51_groupi_n_1478 ,csa_tree_add_12_51_groupi_n_1477);
  not csa_tree_add_12_51_groupi_drc_bufs23510(csa_tree_add_12_51_groupi_n_1477 ,csa_tree_add_12_51_groupi_n_2090);
  not csa_tree_add_12_51_groupi_drc_bufs23512(csa_tree_add_12_51_groupi_n_1476 ,csa_tree_add_12_51_groupi_n_1474);
  not csa_tree_add_12_51_groupi_drc_bufs23513(csa_tree_add_12_51_groupi_n_1475 ,csa_tree_add_12_51_groupi_n_1474);
  not csa_tree_add_12_51_groupi_drc_bufs23514(csa_tree_add_12_51_groupi_n_1474 ,csa_tree_add_12_51_groupi_n_3500);
  not csa_tree_add_12_51_groupi_drc_bufs23516(csa_tree_add_12_51_groupi_n_1473 ,csa_tree_add_12_51_groupi_n_1471);
  not csa_tree_add_12_51_groupi_drc_bufs23517(csa_tree_add_12_51_groupi_n_1472 ,csa_tree_add_12_51_groupi_n_1471);
  not csa_tree_add_12_51_groupi_drc_bufs23518(csa_tree_add_12_51_groupi_n_1471 ,csa_tree_add_12_51_groupi_n_2342);
  not csa_tree_add_12_51_groupi_drc_bufs23520(csa_tree_add_12_51_groupi_n_1470 ,csa_tree_add_12_51_groupi_n_1468);
  not csa_tree_add_12_51_groupi_drc_bufs23521(csa_tree_add_12_51_groupi_n_1469 ,csa_tree_add_12_51_groupi_n_1468);
  not csa_tree_add_12_51_groupi_drc_bufs23522(csa_tree_add_12_51_groupi_n_1468 ,csa_tree_add_12_51_groupi_n_2334);
  not csa_tree_add_12_51_groupi_drc_bufs23524(csa_tree_add_12_51_groupi_n_1467 ,csa_tree_add_12_51_groupi_n_1465);
  not csa_tree_add_12_51_groupi_drc_bufs23525(csa_tree_add_12_51_groupi_n_1466 ,csa_tree_add_12_51_groupi_n_1465);
  not csa_tree_add_12_51_groupi_drc_bufs23526(csa_tree_add_12_51_groupi_n_1465 ,csa_tree_add_12_51_groupi_n_2333);
  not csa_tree_add_12_51_groupi_drc_bufs23528(csa_tree_add_12_51_groupi_n_1464 ,csa_tree_add_12_51_groupi_n_1462);
  not csa_tree_add_12_51_groupi_drc_bufs23529(csa_tree_add_12_51_groupi_n_1463 ,csa_tree_add_12_51_groupi_n_1462);
  not csa_tree_add_12_51_groupi_drc_bufs23530(csa_tree_add_12_51_groupi_n_1462 ,csa_tree_add_12_51_groupi_n_2325);
  not csa_tree_add_12_51_groupi_drc_bufs23532(csa_tree_add_12_51_groupi_n_1461 ,csa_tree_add_12_51_groupi_n_1459);
  not csa_tree_add_12_51_groupi_drc_bufs23533(csa_tree_add_12_51_groupi_n_1460 ,csa_tree_add_12_51_groupi_n_1459);
  not csa_tree_add_12_51_groupi_drc_bufs23534(csa_tree_add_12_51_groupi_n_1459 ,csa_tree_add_12_51_groupi_n_2324);
  not csa_tree_add_12_51_groupi_drc_bufs23536(csa_tree_add_12_51_groupi_n_1458 ,csa_tree_add_12_51_groupi_n_1456);
  not csa_tree_add_12_51_groupi_drc_bufs23537(csa_tree_add_12_51_groupi_n_1457 ,csa_tree_add_12_51_groupi_n_1456);
  not csa_tree_add_12_51_groupi_drc_bufs23538(csa_tree_add_12_51_groupi_n_1456 ,csa_tree_add_12_51_groupi_n_2316);
  not csa_tree_add_12_51_groupi_drc_bufs23540(csa_tree_add_12_51_groupi_n_1455 ,csa_tree_add_12_51_groupi_n_1453);
  not csa_tree_add_12_51_groupi_drc_bufs23541(csa_tree_add_12_51_groupi_n_1454 ,csa_tree_add_12_51_groupi_n_1453);
  not csa_tree_add_12_51_groupi_drc_bufs23542(csa_tree_add_12_51_groupi_n_1453 ,csa_tree_add_12_51_groupi_n_2315);
  not csa_tree_add_12_51_groupi_drc_bufs23544(csa_tree_add_12_51_groupi_n_1452 ,csa_tree_add_12_51_groupi_n_1450);
  not csa_tree_add_12_51_groupi_drc_bufs23545(csa_tree_add_12_51_groupi_n_1451 ,csa_tree_add_12_51_groupi_n_1450);
  not csa_tree_add_12_51_groupi_drc_bufs23546(csa_tree_add_12_51_groupi_n_1450 ,csa_tree_add_12_51_groupi_n_2307);
  not csa_tree_add_12_51_groupi_drc_bufs23548(csa_tree_add_12_51_groupi_n_1449 ,csa_tree_add_12_51_groupi_n_1447);
  not csa_tree_add_12_51_groupi_drc_bufs23549(csa_tree_add_12_51_groupi_n_1448 ,csa_tree_add_12_51_groupi_n_1447);
  not csa_tree_add_12_51_groupi_drc_bufs23550(csa_tree_add_12_51_groupi_n_1447 ,csa_tree_add_12_51_groupi_n_2306);
  not csa_tree_add_12_51_groupi_drc_bufs23552(csa_tree_add_12_51_groupi_n_1446 ,csa_tree_add_12_51_groupi_n_1444);
  not csa_tree_add_12_51_groupi_drc_bufs23553(csa_tree_add_12_51_groupi_n_1445 ,csa_tree_add_12_51_groupi_n_1444);
  not csa_tree_add_12_51_groupi_drc_bufs23554(csa_tree_add_12_51_groupi_n_1444 ,csa_tree_add_12_51_groupi_n_2298);
  not csa_tree_add_12_51_groupi_drc_bufs23556(csa_tree_add_12_51_groupi_n_1443 ,csa_tree_add_12_51_groupi_n_1441);
  not csa_tree_add_12_51_groupi_drc_bufs23557(csa_tree_add_12_51_groupi_n_1442 ,csa_tree_add_12_51_groupi_n_1441);
  not csa_tree_add_12_51_groupi_drc_bufs23558(csa_tree_add_12_51_groupi_n_1441 ,csa_tree_add_12_51_groupi_n_2297);
  not csa_tree_add_12_51_groupi_drc_bufs23560(csa_tree_add_12_51_groupi_n_1440 ,csa_tree_add_12_51_groupi_n_1438);
  not csa_tree_add_12_51_groupi_drc_bufs23561(csa_tree_add_12_51_groupi_n_1439 ,csa_tree_add_12_51_groupi_n_1438);
  not csa_tree_add_12_51_groupi_drc_bufs23562(csa_tree_add_12_51_groupi_n_1438 ,csa_tree_add_12_51_groupi_n_2289);
  not csa_tree_add_12_51_groupi_drc_bufs23564(csa_tree_add_12_51_groupi_n_1437 ,csa_tree_add_12_51_groupi_n_1435);
  not csa_tree_add_12_51_groupi_drc_bufs23565(csa_tree_add_12_51_groupi_n_1436 ,csa_tree_add_12_51_groupi_n_1435);
  not csa_tree_add_12_51_groupi_drc_bufs23566(csa_tree_add_12_51_groupi_n_1435 ,csa_tree_add_12_51_groupi_n_2288);
  not csa_tree_add_12_51_groupi_drc_bufs23568(csa_tree_add_12_51_groupi_n_1434 ,csa_tree_add_12_51_groupi_n_1432);
  not csa_tree_add_12_51_groupi_drc_bufs23569(csa_tree_add_12_51_groupi_n_1433 ,csa_tree_add_12_51_groupi_n_1432);
  not csa_tree_add_12_51_groupi_drc_bufs23570(csa_tree_add_12_51_groupi_n_1432 ,csa_tree_add_12_51_groupi_n_2280);
  not csa_tree_add_12_51_groupi_drc_bufs23572(csa_tree_add_12_51_groupi_n_1431 ,csa_tree_add_12_51_groupi_n_1429);
  not csa_tree_add_12_51_groupi_drc_bufs23573(csa_tree_add_12_51_groupi_n_1430 ,csa_tree_add_12_51_groupi_n_1429);
  not csa_tree_add_12_51_groupi_drc_bufs23574(csa_tree_add_12_51_groupi_n_1429 ,csa_tree_add_12_51_groupi_n_2279);
  not csa_tree_add_12_51_groupi_drc_bufs23576(csa_tree_add_12_51_groupi_n_1428 ,csa_tree_add_12_51_groupi_n_1426);
  not csa_tree_add_12_51_groupi_drc_bufs23577(csa_tree_add_12_51_groupi_n_1427 ,csa_tree_add_12_51_groupi_n_1426);
  not csa_tree_add_12_51_groupi_drc_bufs23578(csa_tree_add_12_51_groupi_n_1426 ,csa_tree_add_12_51_groupi_n_2271);
  not csa_tree_add_12_51_groupi_drc_bufs23580(csa_tree_add_12_51_groupi_n_1425 ,csa_tree_add_12_51_groupi_n_1423);
  not csa_tree_add_12_51_groupi_drc_bufs23581(csa_tree_add_12_51_groupi_n_1424 ,csa_tree_add_12_51_groupi_n_1423);
  not csa_tree_add_12_51_groupi_drc_bufs23582(csa_tree_add_12_51_groupi_n_1423 ,csa_tree_add_12_51_groupi_n_2270);
  not csa_tree_add_12_51_groupi_drc_bufs23584(csa_tree_add_12_51_groupi_n_1422 ,csa_tree_add_12_51_groupi_n_1420);
  not csa_tree_add_12_51_groupi_drc_bufs23585(csa_tree_add_12_51_groupi_n_1421 ,csa_tree_add_12_51_groupi_n_1420);
  not csa_tree_add_12_51_groupi_drc_bufs23586(csa_tree_add_12_51_groupi_n_1420 ,csa_tree_add_12_51_groupi_n_2262);
  not csa_tree_add_12_51_groupi_drc_bufs23588(csa_tree_add_12_51_groupi_n_1419 ,csa_tree_add_12_51_groupi_n_1417);
  not csa_tree_add_12_51_groupi_drc_bufs23589(csa_tree_add_12_51_groupi_n_1418 ,csa_tree_add_12_51_groupi_n_1417);
  not csa_tree_add_12_51_groupi_drc_bufs23590(csa_tree_add_12_51_groupi_n_1417 ,csa_tree_add_12_51_groupi_n_2261);
  not csa_tree_add_12_51_groupi_drc_bufs23592(csa_tree_add_12_51_groupi_n_1416 ,csa_tree_add_12_51_groupi_n_1414);
  not csa_tree_add_12_51_groupi_drc_bufs23593(csa_tree_add_12_51_groupi_n_1415 ,csa_tree_add_12_51_groupi_n_1414);
  not csa_tree_add_12_51_groupi_drc_bufs23594(csa_tree_add_12_51_groupi_n_1414 ,csa_tree_add_12_51_groupi_n_2253);
  not csa_tree_add_12_51_groupi_drc_bufs23596(csa_tree_add_12_51_groupi_n_1413 ,csa_tree_add_12_51_groupi_n_1411);
  not csa_tree_add_12_51_groupi_drc_bufs23597(csa_tree_add_12_51_groupi_n_1412 ,csa_tree_add_12_51_groupi_n_1411);
  not csa_tree_add_12_51_groupi_drc_bufs23598(csa_tree_add_12_51_groupi_n_1411 ,csa_tree_add_12_51_groupi_n_2252);
  not csa_tree_add_12_51_groupi_drc_bufs23600(csa_tree_add_12_51_groupi_n_1410 ,csa_tree_add_12_51_groupi_n_1408);
  not csa_tree_add_12_51_groupi_drc_bufs23601(csa_tree_add_12_51_groupi_n_1409 ,csa_tree_add_12_51_groupi_n_1408);
  not csa_tree_add_12_51_groupi_drc_bufs23602(csa_tree_add_12_51_groupi_n_1408 ,csa_tree_add_12_51_groupi_n_2243);
  not csa_tree_add_12_51_groupi_drc_bufs23604(csa_tree_add_12_51_groupi_n_1407 ,csa_tree_add_12_51_groupi_n_1405);
  not csa_tree_add_12_51_groupi_drc_bufs23605(csa_tree_add_12_51_groupi_n_1406 ,csa_tree_add_12_51_groupi_n_1405);
  not csa_tree_add_12_51_groupi_drc_bufs23606(csa_tree_add_12_51_groupi_n_1405 ,csa_tree_add_12_51_groupi_n_2234);
  not csa_tree_add_12_51_groupi_drc_bufs23608(csa_tree_add_12_51_groupi_n_1404 ,csa_tree_add_12_51_groupi_n_1402);
  not csa_tree_add_12_51_groupi_drc_bufs23609(csa_tree_add_12_51_groupi_n_1403 ,csa_tree_add_12_51_groupi_n_1402);
  not csa_tree_add_12_51_groupi_drc_bufs23610(csa_tree_add_12_51_groupi_n_1402 ,csa_tree_add_12_51_groupi_n_2235);
  not csa_tree_add_12_51_groupi_drc_bufs23612(csa_tree_add_12_51_groupi_n_1401 ,csa_tree_add_12_51_groupi_n_1399);
  not csa_tree_add_12_51_groupi_drc_bufs23613(csa_tree_add_12_51_groupi_n_1400 ,csa_tree_add_12_51_groupi_n_1399);
  not csa_tree_add_12_51_groupi_drc_bufs23614(csa_tree_add_12_51_groupi_n_1399 ,csa_tree_add_12_51_groupi_n_2225);
  not csa_tree_add_12_51_groupi_drc_bufs23616(csa_tree_add_12_51_groupi_n_1398 ,csa_tree_add_12_51_groupi_n_1396);
  not csa_tree_add_12_51_groupi_drc_bufs23617(csa_tree_add_12_51_groupi_n_1397 ,csa_tree_add_12_51_groupi_n_1396);
  not csa_tree_add_12_51_groupi_drc_bufs23618(csa_tree_add_12_51_groupi_n_1396 ,csa_tree_add_12_51_groupi_n_2226);
  not csa_tree_add_12_51_groupi_drc_bufs23620(csa_tree_add_12_51_groupi_n_1395 ,csa_tree_add_12_51_groupi_n_1393);
  not csa_tree_add_12_51_groupi_drc_bufs23621(csa_tree_add_12_51_groupi_n_1394 ,csa_tree_add_12_51_groupi_n_1393);
  not csa_tree_add_12_51_groupi_drc_bufs23622(csa_tree_add_12_51_groupi_n_1393 ,csa_tree_add_12_51_groupi_n_2925);
  not csa_tree_add_12_51_groupi_drc_bufs23624(csa_tree_add_12_51_groupi_n_1392 ,csa_tree_add_12_51_groupi_n_1390);
  not csa_tree_add_12_51_groupi_drc_bufs23625(csa_tree_add_12_51_groupi_n_1391 ,csa_tree_add_12_51_groupi_n_1390);
  not csa_tree_add_12_51_groupi_drc_bufs23626(csa_tree_add_12_51_groupi_n_1390 ,csa_tree_add_12_51_groupi_n_2088);
  not csa_tree_add_12_51_groupi_drc_bufs23628(csa_tree_add_12_51_groupi_n_1389 ,csa_tree_add_12_51_groupi_n_1387);
  not csa_tree_add_12_51_groupi_drc_bufs23629(csa_tree_add_12_51_groupi_n_1388 ,csa_tree_add_12_51_groupi_n_1387);
  not csa_tree_add_12_51_groupi_drc_bufs23630(csa_tree_add_12_51_groupi_n_1387 ,csa_tree_add_12_51_groupi_n_2752);
  not csa_tree_add_12_51_groupi_drc_bufs23632(csa_tree_add_12_51_groupi_n_1386 ,csa_tree_add_12_51_groupi_n_1384);
  not csa_tree_add_12_51_groupi_drc_bufs23633(csa_tree_add_12_51_groupi_n_1385 ,csa_tree_add_12_51_groupi_n_1384);
  not csa_tree_add_12_51_groupi_drc_bufs23634(csa_tree_add_12_51_groupi_n_1384 ,csa_tree_add_12_51_groupi_n_3504);
  not csa_tree_add_12_51_groupi_drc_bufs23636(csa_tree_add_12_51_groupi_n_1383 ,csa_tree_add_12_51_groupi_n_1381);
  not csa_tree_add_12_51_groupi_drc_bufs23637(csa_tree_add_12_51_groupi_n_1382 ,csa_tree_add_12_51_groupi_n_1381);
  not csa_tree_add_12_51_groupi_drc_bufs23638(csa_tree_add_12_51_groupi_n_1381 ,csa_tree_add_12_51_groupi_n_2946);
  not csa_tree_add_12_51_groupi_drc_bufs23640(csa_tree_add_12_51_groupi_n_1380 ,csa_tree_add_12_51_groupi_n_1378);
  not csa_tree_add_12_51_groupi_drc_bufs23641(csa_tree_add_12_51_groupi_n_1379 ,csa_tree_add_12_51_groupi_n_1378);
  not csa_tree_add_12_51_groupi_drc_bufs23642(csa_tree_add_12_51_groupi_n_1378 ,csa_tree_add_12_51_groupi_n_2086);
  not csa_tree_add_12_51_groupi_drc_bufs23644(csa_tree_add_12_51_groupi_n_1377 ,csa_tree_add_12_51_groupi_n_1375);
  not csa_tree_add_12_51_groupi_drc_bufs23645(csa_tree_add_12_51_groupi_n_1376 ,csa_tree_add_12_51_groupi_n_1375);
  not csa_tree_add_12_51_groupi_drc_bufs23646(csa_tree_add_12_51_groupi_n_1375 ,csa_tree_add_12_51_groupi_n_2945);
  not csa_tree_add_12_51_groupi_drc_bufs23648(csa_tree_add_12_51_groupi_n_1374 ,csa_tree_add_12_51_groupi_n_1372);
  not csa_tree_add_12_51_groupi_drc_bufs23649(csa_tree_add_12_51_groupi_n_1373 ,csa_tree_add_12_51_groupi_n_1372);
  not csa_tree_add_12_51_groupi_drc_bufs23650(csa_tree_add_12_51_groupi_n_1372 ,csa_tree_add_12_51_groupi_n_3508);
  not csa_tree_add_12_51_groupi_drc_bufs23652(csa_tree_add_12_51_groupi_n_1371 ,csa_tree_add_12_51_groupi_n_1369);
  not csa_tree_add_12_51_groupi_drc_bufs23653(csa_tree_add_12_51_groupi_n_1370 ,csa_tree_add_12_51_groupi_n_1369);
  not csa_tree_add_12_51_groupi_drc_bufs23654(csa_tree_add_12_51_groupi_n_1369 ,csa_tree_add_12_51_groupi_n_2084);
  not csa_tree_add_12_51_groupi_drc_bufs23656(csa_tree_add_12_51_groupi_n_1368 ,csa_tree_add_12_51_groupi_n_1366);
  not csa_tree_add_12_51_groupi_drc_bufs23657(csa_tree_add_12_51_groupi_n_1367 ,csa_tree_add_12_51_groupi_n_1366);
  not csa_tree_add_12_51_groupi_drc_bufs23658(csa_tree_add_12_51_groupi_n_1366 ,csa_tree_add_12_51_groupi_n_2082);
  not csa_tree_add_12_51_groupi_drc_bufs23660(csa_tree_add_12_51_groupi_n_1365 ,csa_tree_add_12_51_groupi_n_1363);
  not csa_tree_add_12_51_groupi_drc_bufs23661(csa_tree_add_12_51_groupi_n_1364 ,csa_tree_add_12_51_groupi_n_1363);
  not csa_tree_add_12_51_groupi_drc_bufs23662(csa_tree_add_12_51_groupi_n_1363 ,csa_tree_add_12_51_groupi_n_3503);
  not csa_tree_add_12_51_groupi_drc_bufs23664(csa_tree_add_12_51_groupi_n_1362 ,csa_tree_add_12_51_groupi_n_1360);
  not csa_tree_add_12_51_groupi_drc_bufs23665(csa_tree_add_12_51_groupi_n_1361 ,csa_tree_add_12_51_groupi_n_1360);
  not csa_tree_add_12_51_groupi_drc_bufs23666(csa_tree_add_12_51_groupi_n_1360 ,csa_tree_add_12_51_groupi_n_2505);
  not csa_tree_add_12_51_groupi_drc_bufs23668(csa_tree_add_12_51_groupi_n_1359 ,csa_tree_add_12_51_groupi_n_1357);
  not csa_tree_add_12_51_groupi_drc_bufs23669(csa_tree_add_12_51_groupi_n_1358 ,csa_tree_add_12_51_groupi_n_1357);
  not csa_tree_add_12_51_groupi_drc_bufs23670(csa_tree_add_12_51_groupi_n_1357 ,csa_tree_add_12_51_groupi_n_3498);
  not csa_tree_add_12_51_groupi_drc_bufs23672(csa_tree_add_12_51_groupi_n_1356 ,csa_tree_add_12_51_groupi_n_1354);
  not csa_tree_add_12_51_groupi_drc_bufs23673(csa_tree_add_12_51_groupi_n_1355 ,csa_tree_add_12_51_groupi_n_1354);
  not csa_tree_add_12_51_groupi_drc_bufs23674(csa_tree_add_12_51_groupi_n_1354 ,csa_tree_add_12_51_groupi_n_2506);
  not csa_tree_add_12_51_groupi_drc_bufs23676(csa_tree_add_12_51_groupi_n_1353 ,csa_tree_add_12_51_groupi_n_1351);
  not csa_tree_add_12_51_groupi_drc_bufs23677(csa_tree_add_12_51_groupi_n_1352 ,csa_tree_add_12_51_groupi_n_1351);
  not csa_tree_add_12_51_groupi_drc_bufs23678(csa_tree_add_12_51_groupi_n_1351 ,csa_tree_add_12_51_groupi_n_2080);
  not csa_tree_add_12_51_groupi_drc_bufs23680(csa_tree_add_12_51_groupi_n_1350 ,csa_tree_add_12_51_groupi_n_1348);
  not csa_tree_add_12_51_groupi_drc_bufs23681(csa_tree_add_12_51_groupi_n_1349 ,csa_tree_add_12_51_groupi_n_1348);
  not csa_tree_add_12_51_groupi_drc_bufs23682(csa_tree_add_12_51_groupi_n_1348 ,csa_tree_add_12_51_groupi_n_2078);
  not csa_tree_add_12_51_groupi_drc_bufs23684(csa_tree_add_12_51_groupi_n_1347 ,csa_tree_add_12_51_groupi_n_1345);
  not csa_tree_add_12_51_groupi_drc_bufs23685(csa_tree_add_12_51_groupi_n_1346 ,csa_tree_add_12_51_groupi_n_1345);
  not csa_tree_add_12_51_groupi_drc_bufs23686(csa_tree_add_12_51_groupi_n_1345 ,csa_tree_add_12_51_groupi_n_2947);
  not csa_tree_add_12_51_groupi_drc_bufs23688(csa_tree_add_12_51_groupi_n_1344 ,csa_tree_add_12_51_groupi_n_1342);
  not csa_tree_add_12_51_groupi_drc_bufs23689(csa_tree_add_12_51_groupi_n_1343 ,csa_tree_add_12_51_groupi_n_1342);
  not csa_tree_add_12_51_groupi_drc_bufs23690(csa_tree_add_12_51_groupi_n_1342 ,csa_tree_add_12_51_groupi_n_2753);
  not csa_tree_add_12_51_groupi_drc_bufs23692(csa_tree_add_12_51_groupi_n_1341 ,csa_tree_add_12_51_groupi_n_1339);
  not csa_tree_add_12_51_groupi_drc_bufs23693(csa_tree_add_12_51_groupi_n_1340 ,csa_tree_add_12_51_groupi_n_1339);
  not csa_tree_add_12_51_groupi_drc_bufs23694(csa_tree_add_12_51_groupi_n_1339 ,csa_tree_add_12_51_groupi_n_2923);
  not csa_tree_add_12_51_groupi_drc_bufs23696(csa_tree_add_12_51_groupi_n_1338 ,csa_tree_add_12_51_groupi_n_1336);
  not csa_tree_add_12_51_groupi_drc_bufs23697(csa_tree_add_12_51_groupi_n_1337 ,csa_tree_add_12_51_groupi_n_1336);
  not csa_tree_add_12_51_groupi_drc_bufs23698(csa_tree_add_12_51_groupi_n_1336 ,csa_tree_add_12_51_groupi_n_2070);
  not csa_tree_add_12_51_groupi_drc_bufs23700(csa_tree_add_12_51_groupi_n_1335 ,csa_tree_add_12_51_groupi_n_1333);
  not csa_tree_add_12_51_groupi_drc_bufs23701(csa_tree_add_12_51_groupi_n_1334 ,csa_tree_add_12_51_groupi_n_1333);
  not csa_tree_add_12_51_groupi_drc_bufs23702(csa_tree_add_12_51_groupi_n_1333 ,csa_tree_add_12_51_groupi_n_2754);
  not csa_tree_add_12_51_groupi_drc_bufs23704(csa_tree_add_12_51_groupi_n_1332 ,csa_tree_add_12_51_groupi_n_1330);
  not csa_tree_add_12_51_groupi_drc_bufs23705(csa_tree_add_12_51_groupi_n_1331 ,csa_tree_add_12_51_groupi_n_1330);
  not csa_tree_add_12_51_groupi_drc_bufs23706(csa_tree_add_12_51_groupi_n_1330 ,csa_tree_add_12_51_groupi_n_2068);
  not csa_tree_add_12_51_groupi_drc_bufs23708(csa_tree_add_12_51_groupi_n_1329 ,csa_tree_add_12_51_groupi_n_1327);
  not csa_tree_add_12_51_groupi_drc_bufs23709(csa_tree_add_12_51_groupi_n_1328 ,csa_tree_add_12_51_groupi_n_1327);
  not csa_tree_add_12_51_groupi_drc_bufs23710(csa_tree_add_12_51_groupi_n_1327 ,csa_tree_add_12_51_groupi_n_2948);
  not csa_tree_add_12_51_groupi_drc_bufs23712(csa_tree_add_12_51_groupi_n_1326 ,csa_tree_add_12_51_groupi_n_1324);
  not csa_tree_add_12_51_groupi_drc_bufs23713(csa_tree_add_12_51_groupi_n_1325 ,csa_tree_add_12_51_groupi_n_1324);
  not csa_tree_add_12_51_groupi_drc_bufs23714(csa_tree_add_12_51_groupi_n_1324 ,csa_tree_add_12_51_groupi_n_2064);
  not csa_tree_add_12_51_groupi_drc_bufs23716(csa_tree_add_12_51_groupi_n_1323 ,csa_tree_add_12_51_groupi_n_1321);
  not csa_tree_add_12_51_groupi_drc_bufs23717(csa_tree_add_12_51_groupi_n_1322 ,csa_tree_add_12_51_groupi_n_1321);
  not csa_tree_add_12_51_groupi_drc_bufs23718(csa_tree_add_12_51_groupi_n_1321 ,csa_tree_add_12_51_groupi_n_2943);
  not csa_tree_add_12_51_groupi_drc_bufs23720(csa_tree_add_12_51_groupi_n_1320 ,csa_tree_add_12_51_groupi_n_1318);
  not csa_tree_add_12_51_groupi_drc_bufs23721(csa_tree_add_12_51_groupi_n_1319 ,csa_tree_add_12_51_groupi_n_1318);
  not csa_tree_add_12_51_groupi_drc_bufs23722(csa_tree_add_12_51_groupi_n_1318 ,csa_tree_add_12_51_groupi_n_3506);
  not csa_tree_add_12_51_groupi_drc_bufs23724(csa_tree_add_12_51_groupi_n_1317 ,csa_tree_add_12_51_groupi_n_1315);
  not csa_tree_add_12_51_groupi_drc_bufs23725(csa_tree_add_12_51_groupi_n_1316 ,csa_tree_add_12_51_groupi_n_1315);
  not csa_tree_add_12_51_groupi_drc_bufs23726(csa_tree_add_12_51_groupi_n_1315 ,csa_tree_add_12_51_groupi_n_2931);
  not csa_tree_add_12_51_groupi_drc_bufs23728(csa_tree_add_12_51_groupi_n_1314 ,csa_tree_add_12_51_groupi_n_1312);
  not csa_tree_add_12_51_groupi_drc_bufs23729(csa_tree_add_12_51_groupi_n_1313 ,csa_tree_add_12_51_groupi_n_1312);
  not csa_tree_add_12_51_groupi_drc_bufs23730(csa_tree_add_12_51_groupi_n_1312 ,csa_tree_add_12_51_groupi_n_2927);
  not csa_tree_add_12_51_groupi_drc_bufs23732(csa_tree_add_12_51_groupi_n_1311 ,csa_tree_add_12_51_groupi_n_1309);
  not csa_tree_add_12_51_groupi_drc_bufs23733(csa_tree_add_12_51_groupi_n_1310 ,csa_tree_add_12_51_groupi_n_1309);
  not csa_tree_add_12_51_groupi_drc_bufs23734(csa_tree_add_12_51_groupi_n_1309 ,csa_tree_add_12_51_groupi_n_3497);
  not csa_tree_add_12_51_groupi_drc_bufs23736(csa_tree_add_12_51_groupi_n_1308 ,csa_tree_add_12_51_groupi_n_1306);
  not csa_tree_add_12_51_groupi_drc_bufs23737(csa_tree_add_12_51_groupi_n_1307 ,csa_tree_add_12_51_groupi_n_1306);
  not csa_tree_add_12_51_groupi_drc_bufs23738(csa_tree_add_12_51_groupi_n_1306 ,csa_tree_add_12_51_groupi_n_2102);
  not csa_tree_add_12_51_groupi_drc_bufs23740(csa_tree_add_12_51_groupi_n_1305 ,csa_tree_add_12_51_groupi_n_1303);
  not csa_tree_add_12_51_groupi_drc_bufs23741(csa_tree_add_12_51_groupi_n_1304 ,csa_tree_add_12_51_groupi_n_1303);
  not csa_tree_add_12_51_groupi_drc_bufs23742(csa_tree_add_12_51_groupi_n_1303 ,csa_tree_add_12_51_groupi_n_2100);
  not csa_tree_add_12_51_groupi_drc_bufs23744(csa_tree_add_12_51_groupi_n_1302 ,csa_tree_add_12_51_groupi_n_1300);
  not csa_tree_add_12_51_groupi_drc_bufs23745(csa_tree_add_12_51_groupi_n_1301 ,csa_tree_add_12_51_groupi_n_1300);
  not csa_tree_add_12_51_groupi_drc_bufs23746(csa_tree_add_12_51_groupi_n_1300 ,csa_tree_add_12_51_groupi_n_2100);
  not csa_tree_add_12_51_groupi_drc_bufs23748(csa_tree_add_12_51_groupi_n_1299 ,csa_tree_add_12_51_groupi_n_1297);
  not csa_tree_add_12_51_groupi_drc_bufs23749(csa_tree_add_12_51_groupi_n_1298 ,csa_tree_add_12_51_groupi_n_1297);
  not csa_tree_add_12_51_groupi_drc_bufs23750(csa_tree_add_12_51_groupi_n_1297 ,csa_tree_add_12_51_groupi_n_2942);
  not csa_tree_add_12_51_groupi_drc_bufs23752(csa_tree_add_12_51_groupi_n_1296 ,csa_tree_add_12_51_groupi_n_1294);
  not csa_tree_add_12_51_groupi_drc_bufs23753(csa_tree_add_12_51_groupi_n_1295 ,csa_tree_add_12_51_groupi_n_1294);
  not csa_tree_add_12_51_groupi_drc_bufs23754(csa_tree_add_12_51_groupi_n_1294 ,csa_tree_add_12_51_groupi_n_2942);
  not csa_tree_add_12_51_groupi_drc_bufs23756(csa_tree_add_12_51_groupi_n_1293 ,csa_tree_add_12_51_groupi_n_1291);
  not csa_tree_add_12_51_groupi_drc_bufs23757(csa_tree_add_12_51_groupi_n_1292 ,csa_tree_add_12_51_groupi_n_1291);
  not csa_tree_add_12_51_groupi_drc_bufs23758(csa_tree_add_12_51_groupi_n_1291 ,csa_tree_add_12_51_groupi_n_2924);
  not csa_tree_add_12_51_groupi_drc_bufs23760(csa_tree_add_12_51_groupi_n_1290 ,csa_tree_add_12_51_groupi_n_1288);
  not csa_tree_add_12_51_groupi_drc_bufs23761(csa_tree_add_12_51_groupi_n_1289 ,csa_tree_add_12_51_groupi_n_1288);
  not csa_tree_add_12_51_groupi_drc_bufs23762(csa_tree_add_12_51_groupi_n_1288 ,csa_tree_add_12_51_groupi_n_2924);
  not csa_tree_add_12_51_groupi_drc_bufs23764(csa_tree_add_12_51_groupi_n_1287 ,csa_tree_add_12_51_groupi_n_1285);
  not csa_tree_add_12_51_groupi_drc_bufs23765(csa_tree_add_12_51_groupi_n_1286 ,csa_tree_add_12_51_groupi_n_1285);
  not csa_tree_add_12_51_groupi_drc_bufs23766(csa_tree_add_12_51_groupi_n_1285 ,csa_tree_add_12_51_groupi_n_2096);
  not csa_tree_add_12_51_groupi_drc_bufs23768(csa_tree_add_12_51_groupi_n_1284 ,csa_tree_add_12_51_groupi_n_1282);
  not csa_tree_add_12_51_groupi_drc_bufs23769(csa_tree_add_12_51_groupi_n_1283 ,csa_tree_add_12_51_groupi_n_1282);
  not csa_tree_add_12_51_groupi_drc_bufs23770(csa_tree_add_12_51_groupi_n_1282 ,csa_tree_add_12_51_groupi_n_2096);
  not csa_tree_add_12_51_groupi_drc_bufs23772(csa_tree_add_12_51_groupi_n_1281 ,csa_tree_add_12_51_groupi_n_1279);
  not csa_tree_add_12_51_groupi_drc_bufs23773(csa_tree_add_12_51_groupi_n_1280 ,csa_tree_add_12_51_groupi_n_1279);
  not csa_tree_add_12_51_groupi_drc_bufs23774(csa_tree_add_12_51_groupi_n_1279 ,csa_tree_add_12_51_groupi_n_2934);
  not csa_tree_add_12_51_groupi_drc_bufs23776(csa_tree_add_12_51_groupi_n_1278 ,csa_tree_add_12_51_groupi_n_1276);
  not csa_tree_add_12_51_groupi_drc_bufs23777(csa_tree_add_12_51_groupi_n_1277 ,csa_tree_add_12_51_groupi_n_1276);
  not csa_tree_add_12_51_groupi_drc_bufs23778(csa_tree_add_12_51_groupi_n_1276 ,csa_tree_add_12_51_groupi_n_2934);
  not csa_tree_add_12_51_groupi_drc_bufs23780(csa_tree_add_12_51_groupi_n_1275 ,csa_tree_add_12_51_groupi_n_1273);
  not csa_tree_add_12_51_groupi_drc_bufs23781(csa_tree_add_12_51_groupi_n_1274 ,csa_tree_add_12_51_groupi_n_1273);
  not csa_tree_add_12_51_groupi_drc_bufs23782(csa_tree_add_12_51_groupi_n_1273 ,csa_tree_add_12_51_groupi_n_2929);
  not csa_tree_add_12_51_groupi_drc_bufs23784(csa_tree_add_12_51_groupi_n_1272 ,csa_tree_add_12_51_groupi_n_1270);
  not csa_tree_add_12_51_groupi_drc_bufs23785(csa_tree_add_12_51_groupi_n_1271 ,csa_tree_add_12_51_groupi_n_1270);
  not csa_tree_add_12_51_groupi_drc_bufs23786(csa_tree_add_12_51_groupi_n_1270 ,csa_tree_add_12_51_groupi_n_2929);
  not csa_tree_add_12_51_groupi_drc_bufs23788(csa_tree_add_12_51_groupi_n_1269 ,csa_tree_add_12_51_groupi_n_1267);
  not csa_tree_add_12_51_groupi_drc_bufs23789(csa_tree_add_12_51_groupi_n_1268 ,csa_tree_add_12_51_groupi_n_1267);
  not csa_tree_add_12_51_groupi_drc_bufs23790(csa_tree_add_12_51_groupi_n_1267 ,csa_tree_add_12_51_groupi_n_2244);
  not csa_tree_add_12_51_groupi_drc_bufs23792(csa_tree_add_12_51_groupi_n_1266 ,csa_tree_add_12_51_groupi_n_1264);
  not csa_tree_add_12_51_groupi_drc_bufs23793(csa_tree_add_12_51_groupi_n_1265 ,csa_tree_add_12_51_groupi_n_1264);
  not csa_tree_add_12_51_groupi_drc_bufs23794(csa_tree_add_12_51_groupi_n_1264 ,csa_tree_add_12_51_groupi_n_2218);
  not csa_tree_add_12_51_groupi_drc_bufs23796(csa_tree_add_12_51_groupi_n_1263 ,csa_tree_add_12_51_groupi_n_1261);
  not csa_tree_add_12_51_groupi_drc_bufs23797(csa_tree_add_12_51_groupi_n_1262 ,csa_tree_add_12_51_groupi_n_1261);
  not csa_tree_add_12_51_groupi_drc_bufs23798(csa_tree_add_12_51_groupi_n_1261 ,csa_tree_add_12_51_groupi_n_2219);
  not csa_tree_add_12_51_groupi_drc_bufs23800(csa_tree_add_12_51_groupi_n_1260 ,csa_tree_add_12_51_groupi_n_1258);
  not csa_tree_add_12_51_groupi_drc_bufs23801(csa_tree_add_12_51_groupi_n_1259 ,csa_tree_add_12_51_groupi_n_1258);
  not csa_tree_add_12_51_groupi_drc_bufs23802(csa_tree_add_12_51_groupi_n_1258 ,csa_tree_add_12_51_groupi_n_3500);
  not csa_tree_add_12_51_groupi_drc_bufs23804(csa_tree_add_12_51_groupi_n_1257 ,csa_tree_add_12_51_groupi_n_1255);
  not csa_tree_add_12_51_groupi_drc_bufs23805(csa_tree_add_12_51_groupi_n_1256 ,csa_tree_add_12_51_groupi_n_1255);
  not csa_tree_add_12_51_groupi_drc_bufs23806(csa_tree_add_12_51_groupi_n_1255 ,csa_tree_add_12_51_groupi_n_2925);
  not csa_tree_add_12_51_groupi_drc_bufs23808(csa_tree_add_12_51_groupi_n_1254 ,csa_tree_add_12_51_groupi_n_1252);
  not csa_tree_add_12_51_groupi_drc_bufs23809(csa_tree_add_12_51_groupi_n_1253 ,csa_tree_add_12_51_groupi_n_1252);
  not csa_tree_add_12_51_groupi_drc_bufs23810(csa_tree_add_12_51_groupi_n_1252 ,csa_tree_add_12_51_groupi_n_2088);
  not csa_tree_add_12_51_groupi_drc_bufs23812(csa_tree_add_12_51_groupi_n_1251 ,csa_tree_add_12_51_groupi_n_1249);
  not csa_tree_add_12_51_groupi_drc_bufs23813(csa_tree_add_12_51_groupi_n_1250 ,csa_tree_add_12_51_groupi_n_1249);
  not csa_tree_add_12_51_groupi_drc_bufs23814(csa_tree_add_12_51_groupi_n_1249 ,csa_tree_add_12_51_groupi_n_2752);
  not csa_tree_add_12_51_groupi_drc_bufs23816(csa_tree_add_12_51_groupi_n_1248 ,csa_tree_add_12_51_groupi_n_1246);
  not csa_tree_add_12_51_groupi_drc_bufs23817(csa_tree_add_12_51_groupi_n_1247 ,csa_tree_add_12_51_groupi_n_1246);
  not csa_tree_add_12_51_groupi_drc_bufs23818(csa_tree_add_12_51_groupi_n_1246 ,csa_tree_add_12_51_groupi_n_3504);
  not csa_tree_add_12_51_groupi_drc_bufs23820(csa_tree_add_12_51_groupi_n_1245 ,csa_tree_add_12_51_groupi_n_1243);
  not csa_tree_add_12_51_groupi_drc_bufs23821(csa_tree_add_12_51_groupi_n_1244 ,csa_tree_add_12_51_groupi_n_1243);
  not csa_tree_add_12_51_groupi_drc_bufs23822(csa_tree_add_12_51_groupi_n_1243 ,csa_tree_add_12_51_groupi_n_2946);
  not csa_tree_add_12_51_groupi_drc_bufs23824(csa_tree_add_12_51_groupi_n_1242 ,csa_tree_add_12_51_groupi_n_1240);
  not csa_tree_add_12_51_groupi_drc_bufs23825(csa_tree_add_12_51_groupi_n_1241 ,csa_tree_add_12_51_groupi_n_1240);
  not csa_tree_add_12_51_groupi_drc_bufs23826(csa_tree_add_12_51_groupi_n_1240 ,csa_tree_add_12_51_groupi_n_2086);
  not csa_tree_add_12_51_groupi_drc_bufs23828(csa_tree_add_12_51_groupi_n_1239 ,csa_tree_add_12_51_groupi_n_1237);
  not csa_tree_add_12_51_groupi_drc_bufs23829(csa_tree_add_12_51_groupi_n_1238 ,csa_tree_add_12_51_groupi_n_1237);
  not csa_tree_add_12_51_groupi_drc_bufs23830(csa_tree_add_12_51_groupi_n_1237 ,csa_tree_add_12_51_groupi_n_2945);
  not csa_tree_add_12_51_groupi_drc_bufs23832(csa_tree_add_12_51_groupi_n_1236 ,csa_tree_add_12_51_groupi_n_1234);
  not csa_tree_add_12_51_groupi_drc_bufs23833(csa_tree_add_12_51_groupi_n_1235 ,csa_tree_add_12_51_groupi_n_1234);
  not csa_tree_add_12_51_groupi_drc_bufs23834(csa_tree_add_12_51_groupi_n_1234 ,csa_tree_add_12_51_groupi_n_3508);
  not csa_tree_add_12_51_groupi_drc_bufs23836(csa_tree_add_12_51_groupi_n_1233 ,csa_tree_add_12_51_groupi_n_1231);
  not csa_tree_add_12_51_groupi_drc_bufs23837(csa_tree_add_12_51_groupi_n_1232 ,csa_tree_add_12_51_groupi_n_1231);
  not csa_tree_add_12_51_groupi_drc_bufs23838(csa_tree_add_12_51_groupi_n_1231 ,csa_tree_add_12_51_groupi_n_2084);
  not csa_tree_add_12_51_groupi_drc_bufs23840(csa_tree_add_12_51_groupi_n_1230 ,csa_tree_add_12_51_groupi_n_1228);
  not csa_tree_add_12_51_groupi_drc_bufs23841(csa_tree_add_12_51_groupi_n_1229 ,csa_tree_add_12_51_groupi_n_1228);
  not csa_tree_add_12_51_groupi_drc_bufs23842(csa_tree_add_12_51_groupi_n_1228 ,csa_tree_add_12_51_groupi_n_2082);
  not csa_tree_add_12_51_groupi_drc_bufs23844(csa_tree_add_12_51_groupi_n_1227 ,csa_tree_add_12_51_groupi_n_1225);
  not csa_tree_add_12_51_groupi_drc_bufs23845(csa_tree_add_12_51_groupi_n_1226 ,csa_tree_add_12_51_groupi_n_1225);
  not csa_tree_add_12_51_groupi_drc_bufs23846(csa_tree_add_12_51_groupi_n_1225 ,csa_tree_add_12_51_groupi_n_3503);
  not csa_tree_add_12_51_groupi_drc_bufs23848(csa_tree_add_12_51_groupi_n_1224 ,csa_tree_add_12_51_groupi_n_1222);
  not csa_tree_add_12_51_groupi_drc_bufs23849(csa_tree_add_12_51_groupi_n_1223 ,csa_tree_add_12_51_groupi_n_1222);
  not csa_tree_add_12_51_groupi_drc_bufs23850(csa_tree_add_12_51_groupi_n_1222 ,csa_tree_add_12_51_groupi_n_3498);
  not csa_tree_add_12_51_groupi_drc_bufs23852(csa_tree_add_12_51_groupi_n_1221 ,csa_tree_add_12_51_groupi_n_1219);
  not csa_tree_add_12_51_groupi_drc_bufs23853(csa_tree_add_12_51_groupi_n_1220 ,csa_tree_add_12_51_groupi_n_1219);
  not csa_tree_add_12_51_groupi_drc_bufs23854(csa_tree_add_12_51_groupi_n_1219 ,csa_tree_add_12_51_groupi_n_2506);
  not csa_tree_add_12_51_groupi_drc_bufs23856(csa_tree_add_12_51_groupi_n_1218 ,csa_tree_add_12_51_groupi_n_1216);
  not csa_tree_add_12_51_groupi_drc_bufs23857(csa_tree_add_12_51_groupi_n_1217 ,csa_tree_add_12_51_groupi_n_1216);
  not csa_tree_add_12_51_groupi_drc_bufs23858(csa_tree_add_12_51_groupi_n_1216 ,csa_tree_add_12_51_groupi_n_2080);
  not csa_tree_add_12_51_groupi_drc_bufs23860(csa_tree_add_12_51_groupi_n_1215 ,csa_tree_add_12_51_groupi_n_1213);
  not csa_tree_add_12_51_groupi_drc_bufs23861(csa_tree_add_12_51_groupi_n_1214 ,csa_tree_add_12_51_groupi_n_1213);
  not csa_tree_add_12_51_groupi_drc_bufs23862(csa_tree_add_12_51_groupi_n_1213 ,csa_tree_add_12_51_groupi_n_2078);
  not csa_tree_add_12_51_groupi_drc_bufs23864(csa_tree_add_12_51_groupi_n_1212 ,csa_tree_add_12_51_groupi_n_1210);
  not csa_tree_add_12_51_groupi_drc_bufs23865(csa_tree_add_12_51_groupi_n_1211 ,csa_tree_add_12_51_groupi_n_1210);
  not csa_tree_add_12_51_groupi_drc_bufs23866(csa_tree_add_12_51_groupi_n_1210 ,csa_tree_add_12_51_groupi_n_2928);
  not csa_tree_add_12_51_groupi_drc_bufs23868(csa_tree_add_12_51_groupi_n_1209 ,csa_tree_add_12_51_groupi_n_1207);
  not csa_tree_add_12_51_groupi_drc_bufs23869(csa_tree_add_12_51_groupi_n_1208 ,csa_tree_add_12_51_groupi_n_1207);
  not csa_tree_add_12_51_groupi_drc_bufs23870(csa_tree_add_12_51_groupi_n_1207 ,csa_tree_add_12_51_groupi_n_2928);
  not csa_tree_add_12_51_groupi_drc_bufs23872(csa_tree_add_12_51_groupi_n_1206 ,csa_tree_add_12_51_groupi_n_1204);
  not csa_tree_add_12_51_groupi_drc_bufs23873(csa_tree_add_12_51_groupi_n_1205 ,csa_tree_add_12_51_groupi_n_1204);
  not csa_tree_add_12_51_groupi_drc_bufs23874(csa_tree_add_12_51_groupi_n_1204 ,csa_tree_add_12_51_groupi_n_2076);
  not csa_tree_add_12_51_groupi_drc_bufs23876(csa_tree_add_12_51_groupi_n_1203 ,csa_tree_add_12_51_groupi_n_1201);
  not csa_tree_add_12_51_groupi_drc_bufs23877(csa_tree_add_12_51_groupi_n_1202 ,csa_tree_add_12_51_groupi_n_1201);
  not csa_tree_add_12_51_groupi_drc_bufs23878(csa_tree_add_12_51_groupi_n_1201 ,csa_tree_add_12_51_groupi_n_2076);
  not csa_tree_add_12_51_groupi_drc_bufs23880(csa_tree_add_12_51_groupi_n_1200 ,csa_tree_add_12_51_groupi_n_1198);
  not csa_tree_add_12_51_groupi_drc_bufs23881(csa_tree_add_12_51_groupi_n_1199 ,csa_tree_add_12_51_groupi_n_1198);
  not csa_tree_add_12_51_groupi_drc_bufs23882(csa_tree_add_12_51_groupi_n_1198 ,csa_tree_add_12_51_groupi_n_2074);
  not csa_tree_add_12_51_groupi_drc_bufs23884(csa_tree_add_12_51_groupi_n_1197 ,csa_tree_add_12_51_groupi_n_1195);
  not csa_tree_add_12_51_groupi_drc_bufs23885(csa_tree_add_12_51_groupi_n_1196 ,csa_tree_add_12_51_groupi_n_1195);
  not csa_tree_add_12_51_groupi_drc_bufs23886(csa_tree_add_12_51_groupi_n_1195 ,csa_tree_add_12_51_groupi_n_2074);
  not csa_tree_add_12_51_groupi_drc_bufs23888(csa_tree_add_12_51_groupi_n_1194 ,csa_tree_add_12_51_groupi_n_1192);
  not csa_tree_add_12_51_groupi_drc_bufs23889(csa_tree_add_12_51_groupi_n_1193 ,csa_tree_add_12_51_groupi_n_1192);
  not csa_tree_add_12_51_groupi_drc_bufs23890(csa_tree_add_12_51_groupi_n_1192 ,csa_tree_add_12_51_groupi_n_2072);
  not csa_tree_add_12_51_groupi_drc_bufs23892(csa_tree_add_12_51_groupi_n_1191 ,csa_tree_add_12_51_groupi_n_1189);
  not csa_tree_add_12_51_groupi_drc_bufs23893(csa_tree_add_12_51_groupi_n_1190 ,csa_tree_add_12_51_groupi_n_1189);
  not csa_tree_add_12_51_groupi_drc_bufs23894(csa_tree_add_12_51_groupi_n_1189 ,csa_tree_add_12_51_groupi_n_2072);
  not csa_tree_add_12_51_groupi_drc_bufs23896(csa_tree_add_12_51_groupi_n_1188 ,csa_tree_add_12_51_groupi_n_1186);
  not csa_tree_add_12_51_groupi_drc_bufs23897(csa_tree_add_12_51_groupi_n_1187 ,csa_tree_add_12_51_groupi_n_1186);
  not csa_tree_add_12_51_groupi_drc_bufs23898(csa_tree_add_12_51_groupi_n_1186 ,csa_tree_add_12_51_groupi_n_2944);
  not csa_tree_add_12_51_groupi_drc_bufs23900(csa_tree_add_12_51_groupi_n_1185 ,csa_tree_add_12_51_groupi_n_1183);
  not csa_tree_add_12_51_groupi_drc_bufs23901(csa_tree_add_12_51_groupi_n_1184 ,csa_tree_add_12_51_groupi_n_1183);
  not csa_tree_add_12_51_groupi_drc_bufs23902(csa_tree_add_12_51_groupi_n_1183 ,csa_tree_add_12_51_groupi_n_2944);
  not csa_tree_add_12_51_groupi_drc_bufs23904(csa_tree_add_12_51_groupi_n_1182 ,csa_tree_add_12_51_groupi_n_1180);
  not csa_tree_add_12_51_groupi_drc_bufs23905(csa_tree_add_12_51_groupi_n_1181 ,csa_tree_add_12_51_groupi_n_1180);
  not csa_tree_add_12_51_groupi_drc_bufs23906(csa_tree_add_12_51_groupi_n_1180 ,csa_tree_add_12_51_groupi_n_3505);
  not csa_tree_add_12_51_groupi_drc_bufs23908(csa_tree_add_12_51_groupi_n_1179 ,csa_tree_add_12_51_groupi_n_1177);
  not csa_tree_add_12_51_groupi_drc_bufs23909(csa_tree_add_12_51_groupi_n_1178 ,csa_tree_add_12_51_groupi_n_1177);
  not csa_tree_add_12_51_groupi_drc_bufs23910(csa_tree_add_12_51_groupi_n_1177 ,csa_tree_add_12_51_groupi_n_3505);
  not csa_tree_add_12_51_groupi_drc_bufs23912(csa_tree_add_12_51_groupi_n_1176 ,csa_tree_add_12_51_groupi_n_1174);
  not csa_tree_add_12_51_groupi_drc_bufs23913(csa_tree_add_12_51_groupi_n_1175 ,csa_tree_add_12_51_groupi_n_1174);
  not csa_tree_add_12_51_groupi_drc_bufs23914(csa_tree_add_12_51_groupi_n_1174 ,csa_tree_add_12_51_groupi_n_2066);
  not csa_tree_add_12_51_groupi_drc_bufs23916(csa_tree_add_12_51_groupi_n_1173 ,csa_tree_add_12_51_groupi_n_1171);
  not csa_tree_add_12_51_groupi_drc_bufs23917(csa_tree_add_12_51_groupi_n_1172 ,csa_tree_add_12_51_groupi_n_1171);
  not csa_tree_add_12_51_groupi_drc_bufs23918(csa_tree_add_12_51_groupi_n_1171 ,csa_tree_add_12_51_groupi_n_2066);
  not csa_tree_add_12_51_groupi_drc_bufs23920(csa_tree_add_12_51_groupi_n_1170 ,csa_tree_add_12_51_groupi_n_1168);
  not csa_tree_add_12_51_groupi_drc_bufs23921(csa_tree_add_12_51_groupi_n_1169 ,csa_tree_add_12_51_groupi_n_1168);
  not csa_tree_add_12_51_groupi_drc_bufs23922(csa_tree_add_12_51_groupi_n_1168 ,csa_tree_add_12_51_groupi_n_2062);
  not csa_tree_add_12_51_groupi_drc_bufs23924(csa_tree_add_12_51_groupi_n_1167 ,csa_tree_add_12_51_groupi_n_1165);
  not csa_tree_add_12_51_groupi_drc_bufs23925(csa_tree_add_12_51_groupi_n_1166 ,csa_tree_add_12_51_groupi_n_1165);
  not csa_tree_add_12_51_groupi_drc_bufs23926(csa_tree_add_12_51_groupi_n_1165 ,csa_tree_add_12_51_groupi_n_2062);
  not csa_tree_add_12_51_groupi_drc_bufs23928(csa_tree_add_12_51_groupi_n_1164 ,csa_tree_add_12_51_groupi_n_1162);
  not csa_tree_add_12_51_groupi_drc_bufs23929(csa_tree_add_12_51_groupi_n_1163 ,csa_tree_add_12_51_groupi_n_1162);
  not csa_tree_add_12_51_groupi_drc_bufs23930(csa_tree_add_12_51_groupi_n_1162 ,csa_tree_add_12_51_groupi_n_2060);
  not csa_tree_add_12_51_groupi_drc_bufs23932(csa_tree_add_12_51_groupi_n_1161 ,csa_tree_add_12_51_groupi_n_1159);
  not csa_tree_add_12_51_groupi_drc_bufs23933(csa_tree_add_12_51_groupi_n_1160 ,csa_tree_add_12_51_groupi_n_1159);
  not csa_tree_add_12_51_groupi_drc_bufs23934(csa_tree_add_12_51_groupi_n_1159 ,csa_tree_add_12_51_groupi_n_2060);
  not csa_tree_add_12_51_groupi_drc_bufs23936(csa_tree_add_12_51_groupi_n_1158 ,csa_tree_add_12_51_groupi_n_1156);
  not csa_tree_add_12_51_groupi_drc_bufs23937(csa_tree_add_12_51_groupi_n_1157 ,csa_tree_add_12_51_groupi_n_1156);
  not csa_tree_add_12_51_groupi_drc_bufs23938(csa_tree_add_12_51_groupi_n_1156 ,csa_tree_add_12_51_groupi_n_2058);
  not csa_tree_add_12_51_groupi_drc_bufs23940(csa_tree_add_12_51_groupi_n_1155 ,csa_tree_add_12_51_groupi_n_1153);
  not csa_tree_add_12_51_groupi_drc_bufs23941(csa_tree_add_12_51_groupi_n_1154 ,csa_tree_add_12_51_groupi_n_1153);
  not csa_tree_add_12_51_groupi_drc_bufs23942(csa_tree_add_12_51_groupi_n_1153 ,csa_tree_add_12_51_groupi_n_2058);
  not csa_tree_add_12_51_groupi_drc_bufs23944(csa_tree_add_12_51_groupi_n_1152 ,csa_tree_add_12_51_groupi_n_1150);
  not csa_tree_add_12_51_groupi_drc_bufs23945(csa_tree_add_12_51_groupi_n_1151 ,csa_tree_add_12_51_groupi_n_1150);
  not csa_tree_add_12_51_groupi_drc_bufs23946(csa_tree_add_12_51_groupi_n_1150 ,csa_tree_add_12_51_groupi_n_3499);
  not csa_tree_add_12_51_groupi_drc_bufs23948(csa_tree_add_12_51_groupi_n_1149 ,csa_tree_add_12_51_groupi_n_1147);
  not csa_tree_add_12_51_groupi_drc_bufs23949(csa_tree_add_12_51_groupi_n_1148 ,csa_tree_add_12_51_groupi_n_1147);
  not csa_tree_add_12_51_groupi_drc_bufs23950(csa_tree_add_12_51_groupi_n_1147 ,csa_tree_add_12_51_groupi_n_3499);
  not csa_tree_add_12_51_groupi_drc_bufs23952(csa_tree_add_12_51_groupi_n_1146 ,csa_tree_add_12_51_groupi_n_1144);
  not csa_tree_add_12_51_groupi_drc_bufs23953(csa_tree_add_12_51_groupi_n_1145 ,csa_tree_add_12_51_groupi_n_1144);
  not csa_tree_add_12_51_groupi_drc_bufs23954(csa_tree_add_12_51_groupi_n_1144 ,csa_tree_add_12_51_groupi_n_2056);
  not csa_tree_add_12_51_groupi_drc_bufs23956(csa_tree_add_12_51_groupi_n_1143 ,csa_tree_add_12_51_groupi_n_1141);
  not csa_tree_add_12_51_groupi_drc_bufs23957(csa_tree_add_12_51_groupi_n_1142 ,csa_tree_add_12_51_groupi_n_1141);
  not csa_tree_add_12_51_groupi_drc_bufs23958(csa_tree_add_12_51_groupi_n_1141 ,csa_tree_add_12_51_groupi_n_2056);
  not csa_tree_add_12_51_groupi_drc_bufs23960(csa_tree_add_12_51_groupi_n_1140 ,csa_tree_add_12_51_groupi_n_1138);
  not csa_tree_add_12_51_groupi_drc_bufs23961(csa_tree_add_12_51_groupi_n_1139 ,csa_tree_add_12_51_groupi_n_1138);
  not csa_tree_add_12_51_groupi_drc_bufs23962(csa_tree_add_12_51_groupi_n_1138 ,csa_tree_add_12_51_groupi_n_2054);
  not csa_tree_add_12_51_groupi_drc_bufs23964(csa_tree_add_12_51_groupi_n_1137 ,csa_tree_add_12_51_groupi_n_1135);
  not csa_tree_add_12_51_groupi_drc_bufs23965(csa_tree_add_12_51_groupi_n_1136 ,csa_tree_add_12_51_groupi_n_1135);
  not csa_tree_add_12_51_groupi_drc_bufs23966(csa_tree_add_12_51_groupi_n_1135 ,csa_tree_add_12_51_groupi_n_2054);
  not csa_tree_add_12_51_groupi_drc_bufs23968(csa_tree_add_12_51_groupi_n_1134 ,csa_tree_add_12_51_groupi_n_1132);
  not csa_tree_add_12_51_groupi_drc_bufs23969(csa_tree_add_12_51_groupi_n_1133 ,csa_tree_add_12_51_groupi_n_1132);
  not csa_tree_add_12_51_groupi_drc_bufs23970(csa_tree_add_12_51_groupi_n_1132 ,csa_tree_add_12_51_groupi_n_2052);
  not csa_tree_add_12_51_groupi_drc_bufs23972(csa_tree_add_12_51_groupi_n_1131 ,csa_tree_add_12_51_groupi_n_1129);
  not csa_tree_add_12_51_groupi_drc_bufs23973(csa_tree_add_12_51_groupi_n_1130 ,csa_tree_add_12_51_groupi_n_1129);
  not csa_tree_add_12_51_groupi_drc_bufs23974(csa_tree_add_12_51_groupi_n_1129 ,csa_tree_add_12_51_groupi_n_2050);
  not csa_tree_add_12_51_groupi_drc_bufs23976(csa_tree_add_12_51_groupi_n_1128 ,csa_tree_add_12_51_groupi_n_1126);
  not csa_tree_add_12_51_groupi_drc_bufs23977(csa_tree_add_12_51_groupi_n_1127 ,csa_tree_add_12_51_groupi_n_1126);
  not csa_tree_add_12_51_groupi_drc_bufs23978(csa_tree_add_12_51_groupi_n_1126 ,csa_tree_add_12_51_groupi_n_2922);
  not csa_tree_add_12_51_groupi_drc_bufs23980(csa_tree_add_12_51_groupi_n_1125 ,csa_tree_add_12_51_groupi_n_1123);
  not csa_tree_add_12_51_groupi_drc_bufs23981(csa_tree_add_12_51_groupi_n_1124 ,csa_tree_add_12_51_groupi_n_1123);
  not csa_tree_add_12_51_groupi_drc_bufs23982(csa_tree_add_12_51_groupi_n_1123 ,csa_tree_add_12_51_groupi_n_2048);
  not csa_tree_add_12_51_groupi_drc_bufs23984(csa_tree_add_12_51_groupi_n_1122 ,csa_tree_add_12_51_groupi_n_1120);
  not csa_tree_add_12_51_groupi_drc_bufs23985(csa_tree_add_12_51_groupi_n_1121 ,csa_tree_add_12_51_groupi_n_1120);
  not csa_tree_add_12_51_groupi_drc_bufs23986(csa_tree_add_12_51_groupi_n_1120 ,csa_tree_add_12_51_groupi_n_2046);
  not csa_tree_add_12_51_groupi_drc_bufs23988(csa_tree_add_12_51_groupi_n_1119 ,csa_tree_add_12_51_groupi_n_1117);
  not csa_tree_add_12_51_groupi_drc_bufs23989(csa_tree_add_12_51_groupi_n_1118 ,csa_tree_add_12_51_groupi_n_1117);
  not csa_tree_add_12_51_groupi_drc_bufs23990(csa_tree_add_12_51_groupi_n_1117 ,csa_tree_add_12_51_groupi_n_2098);
  not csa_tree_add_12_51_groupi_drc_bufs23992(csa_tree_add_12_51_groupi_n_1116 ,csa_tree_add_12_51_groupi_n_1114);
  not csa_tree_add_12_51_groupi_drc_bufs23993(csa_tree_add_12_51_groupi_n_1115 ,csa_tree_add_12_51_groupi_n_1114);
  not csa_tree_add_12_51_groupi_drc_bufs23994(csa_tree_add_12_51_groupi_n_1114 ,csa_tree_add_12_51_groupi_n_2044);
  not csa_tree_add_12_51_groupi_drc_bufs23996(csa_tree_add_12_51_groupi_n_1113 ,csa_tree_add_12_51_groupi_n_1111);
  not csa_tree_add_12_51_groupi_drc_bufs23997(csa_tree_add_12_51_groupi_n_1112 ,csa_tree_add_12_51_groupi_n_1111);
  not csa_tree_add_12_51_groupi_drc_bufs23998(csa_tree_add_12_51_groupi_n_1111 ,csa_tree_add_12_51_groupi_n_2042);
  not csa_tree_add_12_51_groupi_drc_bufs24000(csa_tree_add_12_51_groupi_n_1110 ,csa_tree_add_12_51_groupi_n_1108);
  not csa_tree_add_12_51_groupi_drc_bufs24001(csa_tree_add_12_51_groupi_n_1109 ,csa_tree_add_12_51_groupi_n_1108);
  not csa_tree_add_12_51_groupi_drc_bufs24002(csa_tree_add_12_51_groupi_n_1108 ,csa_tree_add_12_51_groupi_n_2040);
  not csa_tree_add_12_51_groupi_drc_bufs24004(csa_tree_add_12_51_groupi_n_1107 ,csa_tree_add_12_51_groupi_n_1105);
  not csa_tree_add_12_51_groupi_drc_bufs24005(csa_tree_add_12_51_groupi_n_1106 ,csa_tree_add_12_51_groupi_n_1105);
  not csa_tree_add_12_51_groupi_drc_bufs24006(csa_tree_add_12_51_groupi_n_1105 ,csa_tree_add_12_51_groupi_n_2941);
  not csa_tree_add_12_51_groupi_drc_bufs24008(csa_tree_add_12_51_groupi_n_1104 ,csa_tree_add_12_51_groupi_n_1102);
  not csa_tree_add_12_51_groupi_drc_bufs24009(csa_tree_add_12_51_groupi_n_1103 ,csa_tree_add_12_51_groupi_n_1102);
  not csa_tree_add_12_51_groupi_drc_bufs24010(csa_tree_add_12_51_groupi_n_1102 ,csa_tree_add_12_51_groupi_n_2038);
  not csa_tree_add_12_51_groupi_drc_bufs24012(csa_tree_add_12_51_groupi_n_1101 ,csa_tree_add_12_51_groupi_n_1099);
  not csa_tree_add_12_51_groupi_drc_bufs24013(csa_tree_add_12_51_groupi_n_1100 ,csa_tree_add_12_51_groupi_n_1099);
  not csa_tree_add_12_51_groupi_drc_bufs24014(csa_tree_add_12_51_groupi_n_1099 ,csa_tree_add_12_51_groupi_n_2933);
  not csa_tree_add_12_51_groupi_drc_bufs24016(csa_tree_add_12_51_groupi_n_1098 ,csa_tree_add_12_51_groupi_n_1096);
  not csa_tree_add_12_51_groupi_drc_bufs24017(csa_tree_add_12_51_groupi_n_1097 ,csa_tree_add_12_51_groupi_n_1096);
  not csa_tree_add_12_51_groupi_drc_bufs24018(csa_tree_add_12_51_groupi_n_1096 ,csa_tree_add_12_51_groupi_n_2036);
  not csa_tree_add_12_51_groupi_drc_bufs24020(csa_tree_add_12_51_groupi_n_1095 ,csa_tree_add_12_51_groupi_n_1093);
  not csa_tree_add_12_51_groupi_drc_bufs24021(csa_tree_add_12_51_groupi_n_1094 ,csa_tree_add_12_51_groupi_n_1093);
  not csa_tree_add_12_51_groupi_drc_bufs24022(csa_tree_add_12_51_groupi_n_1093 ,csa_tree_add_12_51_groupi_n_2932);
  not csa_tree_add_12_51_groupi_drc_bufs24024(csa_tree_add_12_51_groupi_n_1092 ,csa_tree_add_12_51_groupi_n_1090);
  not csa_tree_add_12_51_groupi_drc_bufs24025(csa_tree_add_12_51_groupi_n_1091 ,csa_tree_add_12_51_groupi_n_1090);
  not csa_tree_add_12_51_groupi_drc_bufs24026(csa_tree_add_12_51_groupi_n_1090 ,csa_tree_add_12_51_groupi_n_2034);
  not csa_tree_add_12_51_groupi_drc_bufs24028(csa_tree_add_12_51_groupi_n_1089 ,csa_tree_add_12_51_groupi_n_1087);
  not csa_tree_add_12_51_groupi_drc_bufs24029(csa_tree_add_12_51_groupi_n_1088 ,csa_tree_add_12_51_groupi_n_1087);
  not csa_tree_add_12_51_groupi_drc_bufs24030(csa_tree_add_12_51_groupi_n_1087 ,csa_tree_add_12_51_groupi_n_3502);
  not csa_tree_add_12_51_groupi_drc_bufs24032(csa_tree_add_12_51_groupi_n_1086 ,csa_tree_add_12_51_groupi_n_1084);
  not csa_tree_add_12_51_groupi_drc_bufs24033(csa_tree_add_12_51_groupi_n_1085 ,csa_tree_add_12_51_groupi_n_1084);
  not csa_tree_add_12_51_groupi_drc_bufs24034(csa_tree_add_12_51_groupi_n_1084 ,csa_tree_add_12_51_groupi_n_2032);
  not csa_tree_add_12_51_groupi_drc_bufs24036(csa_tree_add_12_51_groupi_n_1083 ,csa_tree_add_12_51_groupi_n_1081);
  not csa_tree_add_12_51_groupi_drc_bufs24037(csa_tree_add_12_51_groupi_n_1082 ,csa_tree_add_12_51_groupi_n_1081);
  not csa_tree_add_12_51_groupi_drc_bufs24038(csa_tree_add_12_51_groupi_n_1081 ,csa_tree_add_12_51_groupi_n_2094);
  not csa_tree_add_12_51_groupi_drc_bufs24040(csa_tree_add_12_51_groupi_n_1080 ,csa_tree_add_12_51_groupi_n_1078);
  not csa_tree_add_12_51_groupi_drc_bufs24041(csa_tree_add_12_51_groupi_n_1079 ,csa_tree_add_12_51_groupi_n_1078);
  not csa_tree_add_12_51_groupi_drc_bufs24042(csa_tree_add_12_51_groupi_n_1078 ,csa_tree_add_12_51_groupi_n_2030);
  not csa_tree_add_12_51_groupi_drc_bufs24044(csa_tree_add_12_51_groupi_n_1077 ,csa_tree_add_12_51_groupi_n_1075);
  not csa_tree_add_12_51_groupi_drc_bufs24045(csa_tree_add_12_51_groupi_n_1076 ,csa_tree_add_12_51_groupi_n_1075);
  not csa_tree_add_12_51_groupi_drc_bufs24046(csa_tree_add_12_51_groupi_n_1075 ,csa_tree_add_12_51_groupi_n_2028);
  not csa_tree_add_12_51_groupi_drc_bufs24048(csa_tree_add_12_51_groupi_n_1074 ,csa_tree_add_12_51_groupi_n_1072);
  not csa_tree_add_12_51_groupi_drc_bufs24049(csa_tree_add_12_51_groupi_n_1073 ,csa_tree_add_12_51_groupi_n_1072);
  not csa_tree_add_12_51_groupi_drc_bufs24050(csa_tree_add_12_51_groupi_n_1072 ,csa_tree_add_12_51_groupi_n_2026);
  not csa_tree_add_12_51_groupi_drc_bufs24052(csa_tree_add_12_51_groupi_n_1071 ,csa_tree_add_12_51_groupi_n_1069);
  not csa_tree_add_12_51_groupi_drc_bufs24053(csa_tree_add_12_51_groupi_n_1070 ,csa_tree_add_12_51_groupi_n_1069);
  not csa_tree_add_12_51_groupi_drc_bufs24054(csa_tree_add_12_51_groupi_n_1069 ,csa_tree_add_12_51_groupi_n_2637);
  not csa_tree_add_12_51_groupi_drc_bufs24056(csa_tree_add_12_51_groupi_n_1068 ,csa_tree_add_12_51_groupi_n_1066);
  not csa_tree_add_12_51_groupi_drc_bufs24057(csa_tree_add_12_51_groupi_n_1067 ,csa_tree_add_12_51_groupi_n_1066);
  not csa_tree_add_12_51_groupi_drc_bufs24058(csa_tree_add_12_51_groupi_n_1066 ,csa_tree_add_12_51_groupi_n_2092);
  not csa_tree_add_12_51_groupi_drc_bufs24060(csa_tree_add_12_51_groupi_n_1065 ,csa_tree_add_12_51_groupi_n_1063);
  not csa_tree_add_12_51_groupi_drc_bufs24061(csa_tree_add_12_51_groupi_n_1064 ,csa_tree_add_12_51_groupi_n_1063);
  not csa_tree_add_12_51_groupi_drc_bufs24062(csa_tree_add_12_51_groupi_n_1063 ,csa_tree_add_12_51_groupi_n_2024);
  not csa_tree_add_12_51_groupi_drc_bufs24064(csa_tree_add_12_51_groupi_n_1062 ,csa_tree_add_12_51_groupi_n_1060);
  not csa_tree_add_12_51_groupi_drc_bufs24065(csa_tree_add_12_51_groupi_n_1061 ,csa_tree_add_12_51_groupi_n_1060);
  not csa_tree_add_12_51_groupi_drc_bufs24066(csa_tree_add_12_51_groupi_n_1060 ,csa_tree_add_12_51_groupi_n_2020);
  not csa_tree_add_12_51_groupi_drc_bufs24068(csa_tree_add_12_51_groupi_n_1059 ,csa_tree_add_12_51_groupi_n_1057);
  not csa_tree_add_12_51_groupi_drc_bufs24069(csa_tree_add_12_51_groupi_n_1058 ,csa_tree_add_12_51_groupi_n_1057);
  not csa_tree_add_12_51_groupi_drc_bufs24070(csa_tree_add_12_51_groupi_n_1057 ,csa_tree_add_12_51_groupi_n_2938);
  not csa_tree_add_12_51_groupi_drc_bufs24072(csa_tree_add_12_51_groupi_n_1056 ,csa_tree_add_12_51_groupi_n_1054);
  not csa_tree_add_12_51_groupi_drc_bufs24073(csa_tree_add_12_51_groupi_n_1055 ,csa_tree_add_12_51_groupi_n_1054);
  not csa_tree_add_12_51_groupi_drc_bufs24074(csa_tree_add_12_51_groupi_n_1054 ,csa_tree_add_12_51_groupi_n_2018);
  not csa_tree_add_12_51_groupi_drc_bufs24076(csa_tree_add_12_51_groupi_n_1053 ,csa_tree_add_12_51_groupi_n_1051);
  not csa_tree_add_12_51_groupi_drc_bufs24077(csa_tree_add_12_51_groupi_n_1052 ,csa_tree_add_12_51_groupi_n_1051);
  not csa_tree_add_12_51_groupi_drc_bufs24078(csa_tree_add_12_51_groupi_n_1051 ,csa_tree_add_12_51_groupi_n_2090);
  not csa_tree_add_12_51_groupi_drc_bufs24080(csa_tree_add_12_51_groupi_n_1050 ,csa_tree_add_12_51_groupi_n_1048);
  not csa_tree_add_12_51_groupi_drc_bufs24081(csa_tree_add_12_51_groupi_n_1049 ,csa_tree_add_12_51_groupi_n_1048);
  not csa_tree_add_12_51_groupi_drc_bufs24082(csa_tree_add_12_51_groupi_n_1048 ,csa_tree_add_12_51_groupi_n_2210);
  not csa_tree_add_12_51_groupi_drc_bufs24084(csa_tree_add_12_51_groupi_n_1047 ,csa_tree_add_12_51_groupi_n_1045);
  not csa_tree_add_12_51_groupi_drc_bufs24085(csa_tree_add_12_51_groupi_n_1046 ,csa_tree_add_12_51_groupi_n_1045);
  not csa_tree_add_12_51_groupi_drc_bufs24086(csa_tree_add_12_51_groupi_n_1045 ,csa_tree_add_12_51_groupi_n_2209);
  not csa_tree_add_12_51_groupi_drc_bufs24088(csa_tree_add_12_51_groupi_n_1044 ,csa_tree_add_12_51_groupi_n_1042);
  not csa_tree_add_12_51_groupi_drc_bufs24089(csa_tree_add_12_51_groupi_n_1043 ,csa_tree_add_12_51_groupi_n_1042);
  not csa_tree_add_12_51_groupi_drc_bufs24090(csa_tree_add_12_51_groupi_n_1042 ,csa_tree_add_12_51_groupi_n_4839);
  not csa_tree_add_12_51_groupi_drc_bufs24092(csa_tree_add_12_51_groupi_n_1041 ,csa_tree_add_12_51_groupi_n_1039);
  not csa_tree_add_12_51_groupi_drc_bufs24093(csa_tree_add_12_51_groupi_n_1040 ,csa_tree_add_12_51_groupi_n_1039);
  not csa_tree_add_12_51_groupi_drc_bufs24094(csa_tree_add_12_51_groupi_n_1039 ,csa_tree_add_12_51_groupi_n_3229);
  not csa_tree_add_12_51_groupi_drc_bufs24096(csa_tree_add_12_51_groupi_n_1038 ,csa_tree_add_12_51_groupi_n_1036);
  not csa_tree_add_12_51_groupi_drc_bufs24097(csa_tree_add_12_51_groupi_n_1037 ,csa_tree_add_12_51_groupi_n_1036);
  not csa_tree_add_12_51_groupi_drc_bufs24098(csa_tree_add_12_51_groupi_n_1036 ,csa_tree_add_12_51_groupi_n_3229);
  not csa_tree_add_12_51_groupi_drc_bufs24100(csa_tree_add_12_51_groupi_n_1035 ,csa_tree_add_12_51_groupi_n_1033);
  not csa_tree_add_12_51_groupi_drc_bufs24101(csa_tree_add_12_51_groupi_n_1034 ,csa_tree_add_12_51_groupi_n_1033);
  not csa_tree_add_12_51_groupi_drc_bufs24102(csa_tree_add_12_51_groupi_n_1033 ,csa_tree_add_12_51_groupi_n_4665);
  not csa_tree_add_12_51_groupi_drc_bufs24104(csa_tree_add_12_51_groupi_n_1032 ,csa_tree_add_12_51_groupi_n_1030);
  not csa_tree_add_12_51_groupi_drc_bufs24105(csa_tree_add_12_51_groupi_n_1031 ,csa_tree_add_12_51_groupi_n_1030);
  not csa_tree_add_12_51_groupi_drc_bufs24106(csa_tree_add_12_51_groupi_n_1030 ,csa_tree_add_12_51_groupi_n_4665);
  not csa_tree_add_12_51_groupi_drc_bufs24108(csa_tree_add_12_51_groupi_n_1029 ,csa_tree_add_12_51_groupi_n_1027);
  not csa_tree_add_12_51_groupi_drc_bufs24109(csa_tree_add_12_51_groupi_n_1028 ,csa_tree_add_12_51_groupi_n_1027);
  not csa_tree_add_12_51_groupi_drc_bufs24110(csa_tree_add_12_51_groupi_n_1027 ,csa_tree_add_12_51_groupi_n_4487);
  not csa_tree_add_12_51_groupi_drc_bufs24112(csa_tree_add_12_51_groupi_n_1026 ,csa_tree_add_12_51_groupi_n_1024);
  not csa_tree_add_12_51_groupi_drc_bufs24113(csa_tree_add_12_51_groupi_n_1025 ,csa_tree_add_12_51_groupi_n_1024);
  not csa_tree_add_12_51_groupi_drc_bufs24114(csa_tree_add_12_51_groupi_n_1024 ,csa_tree_add_12_51_groupi_n_4487);
  not csa_tree_add_12_51_groupi_drc_bufs24116(csa_tree_add_12_51_groupi_n_1023 ,csa_tree_add_12_51_groupi_n_1021);
  not csa_tree_add_12_51_groupi_drc_bufs24117(csa_tree_add_12_51_groupi_n_1022 ,csa_tree_add_12_51_groupi_n_1021);
  not csa_tree_add_12_51_groupi_drc_bufs24118(csa_tree_add_12_51_groupi_n_1021 ,csa_tree_add_12_51_groupi_n_4299);
  not csa_tree_add_12_51_groupi_drc_bufs24120(csa_tree_add_12_51_groupi_n_1020 ,csa_tree_add_12_51_groupi_n_1018);
  not csa_tree_add_12_51_groupi_drc_bufs24121(csa_tree_add_12_51_groupi_n_1019 ,csa_tree_add_12_51_groupi_n_1018);
  not csa_tree_add_12_51_groupi_drc_bufs24122(csa_tree_add_12_51_groupi_n_1018 ,csa_tree_add_12_51_groupi_n_4299);
  not csa_tree_add_12_51_groupi_drc_bufs24124(csa_tree_add_12_51_groupi_n_1017 ,csa_tree_add_12_51_groupi_n_1015);
  not csa_tree_add_12_51_groupi_drc_bufs24125(csa_tree_add_12_51_groupi_n_1016 ,csa_tree_add_12_51_groupi_n_1015);
  not csa_tree_add_12_51_groupi_drc_bufs24126(csa_tree_add_12_51_groupi_n_1015 ,csa_tree_add_12_51_groupi_n_6024);
  not csa_tree_add_12_51_groupi_drc_bufs24128(csa_tree_add_12_51_groupi_n_1014 ,csa_tree_add_12_51_groupi_n_1012);
  not csa_tree_add_12_51_groupi_drc_bufs24129(csa_tree_add_12_51_groupi_n_1013 ,csa_tree_add_12_51_groupi_n_1012);
  not csa_tree_add_12_51_groupi_drc_bufs24130(csa_tree_add_12_51_groupi_n_1012 ,csa_tree_add_12_51_groupi_n_6024);
  not csa_tree_add_12_51_groupi_drc_bufs24132(csa_tree_add_12_51_groupi_n_1011 ,csa_tree_add_12_51_groupi_n_1009);
  not csa_tree_add_12_51_groupi_drc_bufs24133(csa_tree_add_12_51_groupi_n_1010 ,csa_tree_add_12_51_groupi_n_1009);
  not csa_tree_add_12_51_groupi_drc_bufs24134(csa_tree_add_12_51_groupi_n_1009 ,csa_tree_add_12_51_groupi_n_5499);
  not csa_tree_add_12_51_groupi_drc_bufs24136(csa_tree_add_12_51_groupi_n_1008 ,csa_tree_add_12_51_groupi_n_1006);
  not csa_tree_add_12_51_groupi_drc_bufs24137(csa_tree_add_12_51_groupi_n_1007 ,csa_tree_add_12_51_groupi_n_1006);
  not csa_tree_add_12_51_groupi_drc_bufs24138(csa_tree_add_12_51_groupi_n_1006 ,csa_tree_add_12_51_groupi_n_5499);
  not csa_tree_add_12_51_groupi_drc_bufs24140(csa_tree_add_12_51_groupi_n_1005 ,csa_tree_add_12_51_groupi_n_1003);
  not csa_tree_add_12_51_groupi_drc_bufs24141(csa_tree_add_12_51_groupi_n_1004 ,csa_tree_add_12_51_groupi_n_1003);
  not csa_tree_add_12_51_groupi_drc_bufs24142(csa_tree_add_12_51_groupi_n_1003 ,csa_tree_add_12_51_groupi_n_5346);
  not csa_tree_add_12_51_groupi_drc_bufs24144(csa_tree_add_12_51_groupi_n_1002 ,csa_tree_add_12_51_groupi_n_1000);
  not csa_tree_add_12_51_groupi_drc_bufs24145(csa_tree_add_12_51_groupi_n_1001 ,csa_tree_add_12_51_groupi_n_1000);
  not csa_tree_add_12_51_groupi_drc_bufs24146(csa_tree_add_12_51_groupi_n_1000 ,csa_tree_add_12_51_groupi_n_5346);
  not csa_tree_add_12_51_groupi_drc_bufs24148(csa_tree_add_12_51_groupi_n_999 ,csa_tree_add_12_51_groupi_n_997);
  not csa_tree_add_12_51_groupi_drc_bufs24149(csa_tree_add_12_51_groupi_n_998 ,csa_tree_add_12_51_groupi_n_997);
  not csa_tree_add_12_51_groupi_drc_bufs24150(csa_tree_add_12_51_groupi_n_997 ,csa_tree_add_12_51_groupi_n_4126);
  not csa_tree_add_12_51_groupi_drc_bufs24152(csa_tree_add_12_51_groupi_n_996 ,csa_tree_add_12_51_groupi_n_994);
  not csa_tree_add_12_51_groupi_drc_bufs24153(csa_tree_add_12_51_groupi_n_995 ,csa_tree_add_12_51_groupi_n_994);
  not csa_tree_add_12_51_groupi_drc_bufs24154(csa_tree_add_12_51_groupi_n_994 ,csa_tree_add_12_51_groupi_n_4126);
  not csa_tree_add_12_51_groupi_drc_bufs24156(csa_tree_add_12_51_groupi_n_993 ,csa_tree_add_12_51_groupi_n_991);
  not csa_tree_add_12_51_groupi_drc_bufs24157(csa_tree_add_12_51_groupi_n_992 ,csa_tree_add_12_51_groupi_n_991);
  not csa_tree_add_12_51_groupi_drc_bufs24158(csa_tree_add_12_51_groupi_n_991 ,csa_tree_add_12_51_groupi_n_6206);
  not csa_tree_add_12_51_groupi_drc_bufs24160(csa_tree_add_12_51_groupi_n_990 ,csa_tree_add_12_51_groupi_n_988);
  not csa_tree_add_12_51_groupi_drc_bufs24161(csa_tree_add_12_51_groupi_n_989 ,csa_tree_add_12_51_groupi_n_988);
  not csa_tree_add_12_51_groupi_drc_bufs24162(csa_tree_add_12_51_groupi_n_988 ,csa_tree_add_12_51_groupi_n_6206);
  not csa_tree_add_12_51_groupi_drc_bufs24164(csa_tree_add_12_51_groupi_n_987 ,csa_tree_add_12_51_groupi_n_985);
  not csa_tree_add_12_51_groupi_drc_bufs24165(csa_tree_add_12_51_groupi_n_986 ,csa_tree_add_12_51_groupi_n_985);
  not csa_tree_add_12_51_groupi_drc_bufs24166(csa_tree_add_12_51_groupi_n_985 ,csa_tree_add_12_51_groupi_n_2016);
  not csa_tree_add_12_51_groupi_drc_bufs24168(csa_tree_add_12_51_groupi_n_984 ,csa_tree_add_12_51_groupi_n_982);
  not csa_tree_add_12_51_groupi_drc_bufs24169(csa_tree_add_12_51_groupi_n_983 ,csa_tree_add_12_51_groupi_n_982);
  not csa_tree_add_12_51_groupi_drc_bufs24170(csa_tree_add_12_51_groupi_n_982 ,csa_tree_add_12_51_groupi_n_2016);
  not csa_tree_add_12_51_groupi_drc_bufs24172(csa_tree_add_12_51_groupi_n_981 ,csa_tree_add_12_51_groupi_n_979);
  not csa_tree_add_12_51_groupi_drc_bufs24173(csa_tree_add_12_51_groupi_n_980 ,csa_tree_add_12_51_groupi_n_979);
  not csa_tree_add_12_51_groupi_drc_bufs24174(csa_tree_add_12_51_groupi_n_979 ,csa_tree_add_12_51_groupi_n_2638);
  not csa_tree_add_12_51_groupi_drc_bufs24176(csa_tree_add_12_51_groupi_n_978 ,csa_tree_add_12_51_groupi_n_976);
  not csa_tree_add_12_51_groupi_drc_bufs24177(csa_tree_add_12_51_groupi_n_977 ,csa_tree_add_12_51_groupi_n_976);
  not csa_tree_add_12_51_groupi_drc_bufs24178(csa_tree_add_12_51_groupi_n_976 ,csa_tree_add_12_51_groupi_n_2638);
  not csa_tree_add_12_51_groupi_drc_bufs24180(csa_tree_add_12_51_groupi_n_975 ,csa_tree_add_12_51_groupi_n_973);
  not csa_tree_add_12_51_groupi_drc_bufs24181(csa_tree_add_12_51_groupi_n_974 ,csa_tree_add_12_51_groupi_n_973);
  not csa_tree_add_12_51_groupi_drc_bufs24182(csa_tree_add_12_51_groupi_n_973 ,csa_tree_add_12_51_groupi_n_2014);
  not csa_tree_add_12_51_groupi_drc_bufs24184(csa_tree_add_12_51_groupi_n_972 ,csa_tree_add_12_51_groupi_n_970);
  not csa_tree_add_12_51_groupi_drc_bufs24185(csa_tree_add_12_51_groupi_n_971 ,csa_tree_add_12_51_groupi_n_970);
  not csa_tree_add_12_51_groupi_drc_bufs24186(csa_tree_add_12_51_groupi_n_970 ,csa_tree_add_12_51_groupi_n_2014);
  not csa_tree_add_12_51_groupi_drc_bufs24188(csa_tree_add_12_51_groupi_n_969 ,csa_tree_add_12_51_groupi_n_967);
  not csa_tree_add_12_51_groupi_drc_bufs24189(csa_tree_add_12_51_groupi_n_968 ,csa_tree_add_12_51_groupi_n_967);
  not csa_tree_add_12_51_groupi_drc_bufs24190(csa_tree_add_12_51_groupi_n_967 ,csa_tree_add_12_51_groupi_n_2012);
  not csa_tree_add_12_51_groupi_drc_bufs24192(csa_tree_add_12_51_groupi_n_966 ,csa_tree_add_12_51_groupi_n_964);
  not csa_tree_add_12_51_groupi_drc_bufs24193(csa_tree_add_12_51_groupi_n_965 ,csa_tree_add_12_51_groupi_n_964);
  not csa_tree_add_12_51_groupi_drc_bufs24194(csa_tree_add_12_51_groupi_n_964 ,csa_tree_add_12_51_groupi_n_2010);
  not csa_tree_add_12_51_groupi_drc_bufs24196(csa_tree_add_12_51_groupi_n_963 ,csa_tree_add_12_51_groupi_n_961);
  not csa_tree_add_12_51_groupi_drc_bufs24197(csa_tree_add_12_51_groupi_n_962 ,csa_tree_add_12_51_groupi_n_961);
  not csa_tree_add_12_51_groupi_drc_bufs24198(csa_tree_add_12_51_groupi_n_961 ,csa_tree_add_12_51_groupi_n_2028);
  not csa_tree_add_12_51_groupi_drc_bufs24200(csa_tree_add_12_51_groupi_n_960 ,csa_tree_add_12_51_groupi_n_958);
  not csa_tree_add_12_51_groupi_drc_bufs24201(csa_tree_add_12_51_groupi_n_959 ,csa_tree_add_12_51_groupi_n_958);
  not csa_tree_add_12_51_groupi_drc_bufs24202(csa_tree_add_12_51_groupi_n_958 ,csa_tree_add_12_51_groupi_n_1963);
  not csa_tree_add_12_51_groupi_drc_bufs24204(csa_tree_add_12_51_groupi_n_957 ,csa_tree_add_12_51_groupi_n_955);
  not csa_tree_add_12_51_groupi_drc_bufs24205(csa_tree_add_12_51_groupi_n_956 ,csa_tree_add_12_51_groupi_n_955);
  not csa_tree_add_12_51_groupi_drc_bufs24206(csa_tree_add_12_51_groupi_n_955 ,csa_tree_add_12_51_groupi_n_3507);
  not csa_tree_add_12_51_groupi_drc_bufs24208(csa_tree_add_12_51_groupi_n_954 ,csa_tree_add_12_51_groupi_n_952);
  not csa_tree_add_12_51_groupi_drc_bufs24209(csa_tree_add_12_51_groupi_n_953 ,csa_tree_add_12_51_groupi_n_952);
  not csa_tree_add_12_51_groupi_drc_bufs24210(csa_tree_add_12_51_groupi_n_952 ,csa_tree_add_12_51_groupi_n_2933);
  not csa_tree_add_12_51_groupi_drc_bufs24212(csa_tree_add_12_51_groupi_n_951 ,csa_tree_add_12_51_groupi_n_949);
  not csa_tree_add_12_51_groupi_drc_bufs24213(csa_tree_add_12_51_groupi_n_950 ,csa_tree_add_12_51_groupi_n_949);
  not csa_tree_add_12_51_groupi_drc_bufs24214(csa_tree_add_12_51_groupi_n_949 ,csa_tree_add_12_51_groupi_n_2947);
  not csa_tree_add_12_51_groupi_drc_bufs24216(csa_tree_add_12_51_groupi_n_948 ,csa_tree_add_12_51_groupi_n_946);
  not csa_tree_add_12_51_groupi_drc_bufs24217(csa_tree_add_12_51_groupi_n_947 ,csa_tree_add_12_51_groupi_n_946);
  not csa_tree_add_12_51_groupi_drc_bufs24218(csa_tree_add_12_51_groupi_n_946 ,csa_tree_add_12_51_groupi_n_1972);
  not csa_tree_add_12_51_groupi_drc_bufs24220(csa_tree_add_12_51_groupi_n_945 ,csa_tree_add_12_51_groupi_n_943);
  not csa_tree_add_12_51_groupi_drc_bufs24221(csa_tree_add_12_51_groupi_n_944 ,csa_tree_add_12_51_groupi_n_943);
  not csa_tree_add_12_51_groupi_drc_bufs24222(csa_tree_add_12_51_groupi_n_943 ,csa_tree_add_12_51_groupi_n_1981);
  not csa_tree_add_12_51_groupi_drc_bufs24224(csa_tree_add_12_51_groupi_n_942 ,csa_tree_add_12_51_groupi_n_940);
  not csa_tree_add_12_51_groupi_drc_bufs24225(csa_tree_add_12_51_groupi_n_941 ,csa_tree_add_12_51_groupi_n_940);
  not csa_tree_add_12_51_groupi_drc_bufs24226(csa_tree_add_12_51_groupi_n_940 ,csa_tree_add_12_51_groupi_n_2753);
  not csa_tree_add_12_51_groupi_drc_bufs24228(csa_tree_add_12_51_groupi_n_939 ,csa_tree_add_12_51_groupi_n_937);
  not csa_tree_add_12_51_groupi_drc_bufs24229(csa_tree_add_12_51_groupi_n_938 ,csa_tree_add_12_51_groupi_n_937);
  not csa_tree_add_12_51_groupi_drc_bufs24230(csa_tree_add_12_51_groupi_n_937 ,csa_tree_add_12_51_groupi_n_2070);
  not csa_tree_add_12_51_groupi_drc_bufs24232(csa_tree_add_12_51_groupi_n_936 ,csa_tree_add_12_51_groupi_n_934);
  not csa_tree_add_12_51_groupi_drc_bufs24233(csa_tree_add_12_51_groupi_n_935 ,csa_tree_add_12_51_groupi_n_934);
  not csa_tree_add_12_51_groupi_drc_bufs24234(csa_tree_add_12_51_groupi_n_934 ,csa_tree_add_12_51_groupi_n_1969);
  not csa_tree_add_12_51_groupi_drc_bufs24236(csa_tree_add_12_51_groupi_n_933 ,csa_tree_add_12_51_groupi_n_931);
  not csa_tree_add_12_51_groupi_drc_bufs24237(csa_tree_add_12_51_groupi_n_932 ,csa_tree_add_12_51_groupi_n_931);
  not csa_tree_add_12_51_groupi_drc_bufs24238(csa_tree_add_12_51_groupi_n_931 ,csa_tree_add_12_51_groupi_n_2068);
  not csa_tree_add_12_51_groupi_drc_bufs24240(csa_tree_add_12_51_groupi_n_930 ,csa_tree_add_12_51_groupi_n_928);
  not csa_tree_add_12_51_groupi_drc_bufs24241(csa_tree_add_12_51_groupi_n_929 ,csa_tree_add_12_51_groupi_n_928);
  not csa_tree_add_12_51_groupi_drc_bufs24242(csa_tree_add_12_51_groupi_n_928 ,csa_tree_add_12_51_groupi_n_1975);
  not csa_tree_add_12_51_groupi_drc_bufs24244(csa_tree_add_12_51_groupi_n_927 ,csa_tree_add_12_51_groupi_n_925);
  not csa_tree_add_12_51_groupi_drc_bufs24245(csa_tree_add_12_51_groupi_n_926 ,csa_tree_add_12_51_groupi_n_925);
  not csa_tree_add_12_51_groupi_drc_bufs24246(csa_tree_add_12_51_groupi_n_925 ,csa_tree_add_12_51_groupi_n_2064);
  not csa_tree_add_12_51_groupi_drc_bufs24248(csa_tree_add_12_51_groupi_n_924 ,csa_tree_add_12_51_groupi_n_922);
  not csa_tree_add_12_51_groupi_drc_bufs24249(csa_tree_add_12_51_groupi_n_923 ,csa_tree_add_12_51_groupi_n_922);
  not csa_tree_add_12_51_groupi_drc_bufs24250(csa_tree_add_12_51_groupi_n_922 ,csa_tree_add_12_51_groupi_n_2931);
  not csa_tree_add_12_51_groupi_drc_bufs24252(csa_tree_add_12_51_groupi_n_921 ,csa_tree_add_12_51_groupi_n_919);
  not csa_tree_add_12_51_groupi_drc_bufs24253(csa_tree_add_12_51_groupi_n_920 ,csa_tree_add_12_51_groupi_n_919);
  not csa_tree_add_12_51_groupi_drc_bufs24254(csa_tree_add_12_51_groupi_n_919 ,csa_tree_add_12_51_groupi_n_2052);
  not csa_tree_add_12_51_groupi_drc_bufs24256(csa_tree_add_12_51_groupi_n_918 ,csa_tree_add_12_51_groupi_n_916);
  not csa_tree_add_12_51_groupi_drc_bufs24257(csa_tree_add_12_51_groupi_n_917 ,csa_tree_add_12_51_groupi_n_916);
  not csa_tree_add_12_51_groupi_drc_bufs24258(csa_tree_add_12_51_groupi_n_916 ,csa_tree_add_12_51_groupi_n_2050);
  not csa_tree_add_12_51_groupi_drc_bufs24260(csa_tree_add_12_51_groupi_n_915 ,csa_tree_add_12_51_groupi_n_913);
  not csa_tree_add_12_51_groupi_drc_bufs24261(csa_tree_add_12_51_groupi_n_914 ,csa_tree_add_12_51_groupi_n_913);
  not csa_tree_add_12_51_groupi_drc_bufs24262(csa_tree_add_12_51_groupi_n_913 ,csa_tree_add_12_51_groupi_n_2922);
  not csa_tree_add_12_51_groupi_drc_bufs24264(csa_tree_add_12_51_groupi_n_912 ,csa_tree_add_12_51_groupi_n_910);
  not csa_tree_add_12_51_groupi_drc_bufs24265(csa_tree_add_12_51_groupi_n_911 ,csa_tree_add_12_51_groupi_n_910);
  not csa_tree_add_12_51_groupi_drc_bufs24266(csa_tree_add_12_51_groupi_n_910 ,csa_tree_add_12_51_groupi_n_2048);
  not csa_tree_add_12_51_groupi_drc_bufs24268(csa_tree_add_12_51_groupi_n_909 ,csa_tree_add_12_51_groupi_n_907);
  not csa_tree_add_12_51_groupi_drc_bufs24269(csa_tree_add_12_51_groupi_n_908 ,csa_tree_add_12_51_groupi_n_907);
  not csa_tree_add_12_51_groupi_drc_bufs24270(csa_tree_add_12_51_groupi_n_907 ,csa_tree_add_12_51_groupi_n_1999);
  not csa_tree_add_12_51_groupi_drc_bufs24272(csa_tree_add_12_51_groupi_n_906 ,csa_tree_add_12_51_groupi_n_904);
  not csa_tree_add_12_51_groupi_drc_bufs24273(csa_tree_add_12_51_groupi_n_905 ,csa_tree_add_12_51_groupi_n_904);
  not csa_tree_add_12_51_groupi_drc_bufs24274(csa_tree_add_12_51_groupi_n_904 ,csa_tree_add_12_51_groupi_n_2046);
  not csa_tree_add_12_51_groupi_drc_bufs24276(csa_tree_add_12_51_groupi_n_903 ,csa_tree_add_12_51_groupi_n_901);
  not csa_tree_add_12_51_groupi_drc_bufs24277(csa_tree_add_12_51_groupi_n_902 ,csa_tree_add_12_51_groupi_n_901);
  not csa_tree_add_12_51_groupi_drc_bufs24278(csa_tree_add_12_51_groupi_n_901 ,csa_tree_add_12_51_groupi_n_2044);
  not csa_tree_add_12_51_groupi_drc_bufs24280(csa_tree_add_12_51_groupi_n_900 ,csa_tree_add_12_51_groupi_n_898);
  not csa_tree_add_12_51_groupi_drc_bufs24281(csa_tree_add_12_51_groupi_n_899 ,csa_tree_add_12_51_groupi_n_898);
  not csa_tree_add_12_51_groupi_drc_bufs24282(csa_tree_add_12_51_groupi_n_898 ,csa_tree_add_12_51_groupi_n_2005);
  not csa_tree_add_12_51_groupi_drc_bufs24284(csa_tree_add_12_51_groupi_n_897 ,csa_tree_add_12_51_groupi_n_895);
  not csa_tree_add_12_51_groupi_drc_bufs24285(csa_tree_add_12_51_groupi_n_896 ,csa_tree_add_12_51_groupi_n_895);
  not csa_tree_add_12_51_groupi_drc_bufs24286(csa_tree_add_12_51_groupi_n_895 ,csa_tree_add_12_51_groupi_n_2042);
  not csa_tree_add_12_51_groupi_drc_bufs24288(csa_tree_add_12_51_groupi_n_894 ,csa_tree_add_12_51_groupi_n_892);
  not csa_tree_add_12_51_groupi_drc_bufs24289(csa_tree_add_12_51_groupi_n_893 ,csa_tree_add_12_51_groupi_n_892);
  not csa_tree_add_12_51_groupi_drc_bufs24290(csa_tree_add_12_51_groupi_n_892 ,csa_tree_add_12_51_groupi_n_2008);
  not csa_tree_add_12_51_groupi_drc_bufs24292(csa_tree_add_12_51_groupi_n_891 ,csa_tree_add_12_51_groupi_n_889);
  not csa_tree_add_12_51_groupi_drc_bufs24293(csa_tree_add_12_51_groupi_n_890 ,csa_tree_add_12_51_groupi_n_889);
  not csa_tree_add_12_51_groupi_drc_bufs24294(csa_tree_add_12_51_groupi_n_889 ,csa_tree_add_12_51_groupi_n_2040);
  not csa_tree_add_12_51_groupi_drc_bufs24296(csa_tree_add_12_51_groupi_n_888 ,csa_tree_add_12_51_groupi_n_886);
  not csa_tree_add_12_51_groupi_drc_bufs24297(csa_tree_add_12_51_groupi_n_887 ,csa_tree_add_12_51_groupi_n_886);
  not csa_tree_add_12_51_groupi_drc_bufs24298(csa_tree_add_12_51_groupi_n_886 ,csa_tree_add_12_51_groupi_n_2038);
  not csa_tree_add_12_51_groupi_drc_bufs24300(csa_tree_add_12_51_groupi_n_885 ,csa_tree_add_12_51_groupi_n_883);
  not csa_tree_add_12_51_groupi_drc_bufs24301(csa_tree_add_12_51_groupi_n_884 ,csa_tree_add_12_51_groupi_n_883);
  not csa_tree_add_12_51_groupi_drc_bufs24302(csa_tree_add_12_51_groupi_n_883 ,csa_tree_add_12_51_groupi_n_2026);
  not csa_tree_add_12_51_groupi_drc_bufs24304(csa_tree_add_12_51_groupi_n_882 ,csa_tree_add_12_51_groupi_n_880);
  not csa_tree_add_12_51_groupi_drc_bufs24305(csa_tree_add_12_51_groupi_n_881 ,csa_tree_add_12_51_groupi_n_880);
  not csa_tree_add_12_51_groupi_drc_bufs24306(csa_tree_add_12_51_groupi_n_880 ,csa_tree_add_12_51_groupi_n_2036);
  not csa_tree_add_12_51_groupi_drc_bufs24308(csa_tree_add_12_51_groupi_n_879 ,csa_tree_add_12_51_groupi_n_877);
  not csa_tree_add_12_51_groupi_drc_bufs24309(csa_tree_add_12_51_groupi_n_878 ,csa_tree_add_12_51_groupi_n_877);
  not csa_tree_add_12_51_groupi_drc_bufs24310(csa_tree_add_12_51_groupi_n_877 ,csa_tree_add_12_51_groupi_n_2034);
  not csa_tree_add_12_51_groupi_drc_bufs24312(csa_tree_add_12_51_groupi_n_876 ,csa_tree_add_12_51_groupi_n_874);
  not csa_tree_add_12_51_groupi_drc_bufs24313(csa_tree_add_12_51_groupi_n_875 ,csa_tree_add_12_51_groupi_n_874);
  not csa_tree_add_12_51_groupi_drc_bufs24314(csa_tree_add_12_51_groupi_n_874 ,csa_tree_add_12_51_groupi_n_3502);
  not csa_tree_add_12_51_groupi_drc_bufs24316(csa_tree_add_12_51_groupi_n_873 ,csa_tree_add_12_51_groupi_n_871);
  not csa_tree_add_12_51_groupi_drc_bufs24317(csa_tree_add_12_51_groupi_n_872 ,csa_tree_add_12_51_groupi_n_871);
  not csa_tree_add_12_51_groupi_drc_bufs24318(csa_tree_add_12_51_groupi_n_871 ,csa_tree_add_12_51_groupi_n_2032);
  not csa_tree_add_12_51_groupi_drc_bufs24320(csa_tree_add_12_51_groupi_n_870 ,csa_tree_add_12_51_groupi_n_868);
  not csa_tree_add_12_51_groupi_drc_bufs24321(csa_tree_add_12_51_groupi_n_869 ,csa_tree_add_12_51_groupi_n_868);
  not csa_tree_add_12_51_groupi_drc_bufs24322(csa_tree_add_12_51_groupi_n_868 ,csa_tree_add_12_51_groupi_n_2030);
  not csa_tree_add_12_51_groupi_drc_bufs24324(csa_tree_add_12_51_groupi_n_867 ,csa_tree_add_12_51_groupi_n_865);
  not csa_tree_add_12_51_groupi_drc_bufs24325(csa_tree_add_12_51_groupi_n_866 ,csa_tree_add_12_51_groupi_n_865);
  not csa_tree_add_12_51_groupi_drc_bufs24326(csa_tree_add_12_51_groupi_n_865 ,csa_tree_add_12_51_groupi_n_2637);
  not csa_tree_add_12_51_groupi_drc_bufs24328(csa_tree_add_12_51_groupi_n_864 ,csa_tree_add_12_51_groupi_n_862);
  not csa_tree_add_12_51_groupi_drc_bufs24329(csa_tree_add_12_51_groupi_n_863 ,csa_tree_add_12_51_groupi_n_862);
  not csa_tree_add_12_51_groupi_drc_bufs24330(csa_tree_add_12_51_groupi_n_862 ,csa_tree_add_12_51_groupi_n_2024);
  not csa_tree_add_12_51_groupi_drc_bufs24332(csa_tree_add_12_51_groupi_n_861 ,csa_tree_add_12_51_groupi_n_859);
  not csa_tree_add_12_51_groupi_drc_bufs24333(csa_tree_add_12_51_groupi_n_860 ,csa_tree_add_12_51_groupi_n_859);
  not csa_tree_add_12_51_groupi_drc_bufs24334(csa_tree_add_12_51_groupi_n_859 ,csa_tree_add_12_51_groupi_n_2002);
  not csa_tree_add_12_51_groupi_drc_bufs24336(csa_tree_add_12_51_groupi_n_858 ,csa_tree_add_12_51_groupi_n_856);
  not csa_tree_add_12_51_groupi_drc_bufs24337(csa_tree_add_12_51_groupi_n_857 ,csa_tree_add_12_51_groupi_n_856);
  not csa_tree_add_12_51_groupi_drc_bufs24338(csa_tree_add_12_51_groupi_n_856 ,csa_tree_add_12_51_groupi_n_2022);
  not csa_tree_add_12_51_groupi_drc_bufs24340(csa_tree_add_12_51_groupi_n_855 ,csa_tree_add_12_51_groupi_n_853);
  not csa_tree_add_12_51_groupi_drc_bufs24341(csa_tree_add_12_51_groupi_n_854 ,csa_tree_add_12_51_groupi_n_853);
  not csa_tree_add_12_51_groupi_drc_bufs24342(csa_tree_add_12_51_groupi_n_853 ,csa_tree_add_12_51_groupi_n_2022);
  not csa_tree_add_12_51_groupi_drc_bufs24344(csa_tree_add_12_51_groupi_n_852 ,csa_tree_add_12_51_groupi_n_850);
  not csa_tree_add_12_51_groupi_drc_bufs24345(csa_tree_add_12_51_groupi_n_851 ,csa_tree_add_12_51_groupi_n_850);
  not csa_tree_add_12_51_groupi_drc_bufs24346(csa_tree_add_12_51_groupi_n_850 ,csa_tree_add_12_51_groupi_n_1996);
  not csa_tree_add_12_51_groupi_drc_bufs24348(csa_tree_add_12_51_groupi_n_849 ,csa_tree_add_12_51_groupi_n_847);
  not csa_tree_add_12_51_groupi_drc_bufs24349(csa_tree_add_12_51_groupi_n_848 ,csa_tree_add_12_51_groupi_n_847);
  not csa_tree_add_12_51_groupi_drc_bufs24350(csa_tree_add_12_51_groupi_n_847 ,csa_tree_add_12_51_groupi_n_1993);
  not csa_tree_add_12_51_groupi_drc_bufs24352(csa_tree_add_12_51_groupi_n_846 ,csa_tree_add_12_51_groupi_n_844);
  not csa_tree_add_12_51_groupi_drc_bufs24353(csa_tree_add_12_51_groupi_n_845 ,csa_tree_add_12_51_groupi_n_844);
  not csa_tree_add_12_51_groupi_drc_bufs24354(csa_tree_add_12_51_groupi_n_844 ,csa_tree_add_12_51_groupi_n_1990);
  not csa_tree_add_12_51_groupi_drc_bufs24356(csa_tree_add_12_51_groupi_n_843 ,csa_tree_add_12_51_groupi_n_841);
  not csa_tree_add_12_51_groupi_drc_bufs24357(csa_tree_add_12_51_groupi_n_842 ,csa_tree_add_12_51_groupi_n_841);
  not csa_tree_add_12_51_groupi_drc_bufs24358(csa_tree_add_12_51_groupi_n_841 ,csa_tree_add_12_51_groupi_n_1987);
  not csa_tree_add_12_51_groupi_drc_bufs24360(csa_tree_add_12_51_groupi_n_840 ,csa_tree_add_12_51_groupi_n_838);
  not csa_tree_add_12_51_groupi_drc_bufs24361(csa_tree_add_12_51_groupi_n_839 ,csa_tree_add_12_51_groupi_n_838);
  not csa_tree_add_12_51_groupi_drc_bufs24362(csa_tree_add_12_51_groupi_n_838 ,csa_tree_add_12_51_groupi_n_1984);
  not csa_tree_add_12_51_groupi_drc_bufs24364(csa_tree_add_12_51_groupi_n_837 ,csa_tree_add_12_51_groupi_n_835);
  not csa_tree_add_12_51_groupi_drc_bufs24365(csa_tree_add_12_51_groupi_n_836 ,csa_tree_add_12_51_groupi_n_835);
  not csa_tree_add_12_51_groupi_drc_bufs24366(csa_tree_add_12_51_groupi_n_835 ,csa_tree_add_12_51_groupi_n_2643);
  not csa_tree_add_12_51_groupi_drc_bufs24368(csa_tree_add_12_51_groupi_n_834 ,csa_tree_add_12_51_groupi_n_832);
  not csa_tree_add_12_51_groupi_drc_bufs24369(csa_tree_add_12_51_groupi_n_833 ,csa_tree_add_12_51_groupi_n_832);
  not csa_tree_add_12_51_groupi_drc_bufs24370(csa_tree_add_12_51_groupi_n_832 ,csa_tree_add_12_51_groupi_n_2643);
  not csa_tree_add_12_51_groupi_drc_bufs24372(csa_tree_add_12_51_groupi_n_831 ,csa_tree_add_12_51_groupi_n_829);
  not csa_tree_add_12_51_groupi_drc_bufs24373(csa_tree_add_12_51_groupi_n_830 ,csa_tree_add_12_51_groupi_n_829);
  not csa_tree_add_12_51_groupi_drc_bufs24374(csa_tree_add_12_51_groupi_n_829 ,csa_tree_add_12_51_groupi_n_1978);
  not csa_tree_add_12_51_groupi_drc_bufs24376(csa_tree_add_12_51_groupi_n_828 ,csa_tree_add_12_51_groupi_n_826);
  not csa_tree_add_12_51_groupi_drc_bufs24377(csa_tree_add_12_51_groupi_n_827 ,csa_tree_add_12_51_groupi_n_826);
  not csa_tree_add_12_51_groupi_drc_bufs24378(csa_tree_add_12_51_groupi_n_826 ,csa_tree_add_12_51_groupi_n_5175);
  not csa_tree_add_12_51_groupi_drc_bufs24380(csa_tree_add_12_51_groupi_n_825 ,csa_tree_add_12_51_groupi_n_823);
  not csa_tree_add_12_51_groupi_drc_bufs24381(csa_tree_add_12_51_groupi_n_824 ,csa_tree_add_12_51_groupi_n_823);
  not csa_tree_add_12_51_groupi_drc_bufs24382(csa_tree_add_12_51_groupi_n_823 ,csa_tree_add_12_51_groupi_n_5175);
  not csa_tree_add_12_51_groupi_drc_bufs24384(csa_tree_add_12_51_groupi_n_822 ,csa_tree_add_12_51_groupi_n_820);
  not csa_tree_add_12_51_groupi_drc_bufs24385(csa_tree_add_12_51_groupi_n_821 ,csa_tree_add_12_51_groupi_n_820);
  not csa_tree_add_12_51_groupi_drc_bufs24386(csa_tree_add_12_51_groupi_n_820 ,csa_tree_add_12_51_groupi_n_3764);
  not csa_tree_add_12_51_groupi_drc_bufs24388(csa_tree_add_12_51_groupi_n_819 ,csa_tree_add_12_51_groupi_n_817);
  not csa_tree_add_12_51_groupi_drc_bufs24389(csa_tree_add_12_51_groupi_n_818 ,csa_tree_add_12_51_groupi_n_817);
  not csa_tree_add_12_51_groupi_drc_bufs24390(csa_tree_add_12_51_groupi_n_817 ,csa_tree_add_12_51_groupi_n_3764);
  not csa_tree_add_12_51_groupi_drc_bufs24392(csa_tree_add_12_51_groupi_n_816 ,csa_tree_add_12_51_groupi_n_814);
  not csa_tree_add_12_51_groupi_drc_bufs24393(csa_tree_add_12_51_groupi_n_815 ,csa_tree_add_12_51_groupi_n_814);
  not csa_tree_add_12_51_groupi_drc_bufs24394(csa_tree_add_12_51_groupi_n_814 ,csa_tree_add_12_51_groupi_n_1966);
  not csa_tree_add_12_51_groupi_drc_bufs24396(csa_tree_add_12_51_groupi_n_813 ,csa_tree_add_12_51_groupi_n_811);
  not csa_tree_add_12_51_groupi_drc_bufs24397(csa_tree_add_12_51_groupi_n_812 ,csa_tree_add_12_51_groupi_n_811);
  not csa_tree_add_12_51_groupi_drc_bufs24398(csa_tree_add_12_51_groupi_n_811 ,csa_tree_add_12_51_groupi_n_4839);
  not csa_tree_add_12_51_groupi_drc_bufs24400(csa_tree_add_12_51_groupi_n_810 ,csa_tree_add_12_51_groupi_n_808);
  not csa_tree_add_12_51_groupi_drc_bufs24401(csa_tree_add_12_51_groupi_n_809 ,csa_tree_add_12_51_groupi_n_808);
  not csa_tree_add_12_51_groupi_drc_bufs24402(csa_tree_add_12_51_groupi_n_808 ,csa_tree_add_12_51_groupi_n_5842);
  not csa_tree_add_12_51_groupi_drc_bufs24404(csa_tree_add_12_51_groupi_n_807 ,csa_tree_add_12_51_groupi_n_805);
  not csa_tree_add_12_51_groupi_drc_bufs24405(csa_tree_add_12_51_groupi_n_806 ,csa_tree_add_12_51_groupi_n_805);
  not csa_tree_add_12_51_groupi_drc_bufs24406(csa_tree_add_12_51_groupi_n_805 ,csa_tree_add_12_51_groupi_n_5842);
  not csa_tree_add_12_51_groupi_drc_bufs24408(csa_tree_add_12_51_groupi_n_804 ,csa_tree_add_12_51_groupi_n_802);
  not csa_tree_add_12_51_groupi_drc_bufs24409(csa_tree_add_12_51_groupi_n_803 ,csa_tree_add_12_51_groupi_n_802);
  not csa_tree_add_12_51_groupi_drc_bufs24410(csa_tree_add_12_51_groupi_n_802 ,csa_tree_add_12_51_groupi_n_5020);
  not csa_tree_add_12_51_groupi_drc_bufs24412(csa_tree_add_12_51_groupi_n_801 ,csa_tree_add_12_51_groupi_n_799);
  not csa_tree_add_12_51_groupi_drc_bufs24413(csa_tree_add_12_51_groupi_n_800 ,csa_tree_add_12_51_groupi_n_799);
  not csa_tree_add_12_51_groupi_drc_bufs24414(csa_tree_add_12_51_groupi_n_799 ,csa_tree_add_12_51_groupi_n_5020);
  not csa_tree_add_12_51_groupi_drc_bufs24416(csa_tree_add_12_51_groupi_n_798 ,csa_tree_add_12_51_groupi_n_796);
  not csa_tree_add_12_51_groupi_drc_bufs24417(csa_tree_add_12_51_groupi_n_797 ,csa_tree_add_12_51_groupi_n_796);
  not csa_tree_add_12_51_groupi_drc_bufs24418(csa_tree_add_12_51_groupi_n_796 ,csa_tree_add_12_51_groupi_n_5676);
  not csa_tree_add_12_51_groupi_drc_bufs24420(csa_tree_add_12_51_groupi_n_795 ,csa_tree_add_12_51_groupi_n_793);
  not csa_tree_add_12_51_groupi_drc_bufs24421(csa_tree_add_12_51_groupi_n_794 ,csa_tree_add_12_51_groupi_n_793);
  not csa_tree_add_12_51_groupi_drc_bufs24422(csa_tree_add_12_51_groupi_n_793 ,csa_tree_add_12_51_groupi_n_5676);
  not csa_tree_add_12_51_groupi_drc_bufs24424(csa_tree_add_12_51_groupi_n_792 ,csa_tree_add_12_51_groupi_n_2357);
  not csa_tree_add_12_51_groupi_drc_bufs24425(csa_tree_add_12_51_groupi_n_791 ,csa_tree_add_12_51_groupi_n_2357);
  not csa_tree_add_12_51_groupi_drc_bufs24428(csa_tree_add_12_51_groupi_n_790 ,csa_tree_add_12_51_groupi_n_2355);
  not csa_tree_add_12_51_groupi_drc_bufs24429(csa_tree_add_12_51_groupi_n_789 ,csa_tree_add_12_51_groupi_n_2355);
  not csa_tree_add_12_51_groupi_drc_bufs24432(csa_tree_add_12_51_groupi_n_788 ,csa_tree_add_12_51_groupi_n_2388);
  not csa_tree_add_12_51_groupi_drc_bufs24433(csa_tree_add_12_51_groupi_n_787 ,csa_tree_add_12_51_groupi_n_2388);
  not csa_tree_add_12_51_groupi_drc_bufs24436(csa_tree_add_12_51_groupi_n_786 ,csa_tree_add_12_51_groupi_n_2360);
  not csa_tree_add_12_51_groupi_drc_bufs24437(csa_tree_add_12_51_groupi_n_785 ,csa_tree_add_12_51_groupi_n_2360);
  not csa_tree_add_12_51_groupi_drc_bufs24440(csa_tree_add_12_51_groupi_n_784 ,csa_tree_add_12_51_groupi_n_2395);
  not csa_tree_add_12_51_groupi_drc_bufs24441(csa_tree_add_12_51_groupi_n_783 ,csa_tree_add_12_51_groupi_n_2395);
  not csa_tree_add_12_51_groupi_drc_bufs24444(csa_tree_add_12_51_groupi_n_782 ,csa_tree_add_12_51_groupi_n_780);
  not csa_tree_add_12_51_groupi_drc_bufs24445(csa_tree_add_12_51_groupi_n_781 ,csa_tree_add_12_51_groupi_n_780);
  not csa_tree_add_12_51_groupi_drc_bufs24446(csa_tree_add_12_51_groupi_n_780 ,csa_tree_add_12_51_groupi_n_2329);
  not csa_tree_add_12_51_groupi_drc_bufs24448(csa_tree_add_12_51_groupi_n_779 ,csa_tree_add_12_51_groupi_n_2394);
  not csa_tree_add_12_51_groupi_drc_bufs24449(csa_tree_add_12_51_groupi_n_778 ,csa_tree_add_12_51_groupi_n_2394);
  not csa_tree_add_12_51_groupi_drc_bufs24452(csa_tree_add_12_51_groupi_n_777 ,csa_tree_add_12_51_groupi_n_775);
  not csa_tree_add_12_51_groupi_drc_bufs24453(csa_tree_add_12_51_groupi_n_776 ,csa_tree_add_12_51_groupi_n_775);
  not csa_tree_add_12_51_groupi_drc_bufs24454(csa_tree_add_12_51_groupi_n_775 ,csa_tree_add_12_51_groupi_n_2320);
  not csa_tree_add_12_51_groupi_drc_bufs24456(csa_tree_add_12_51_groupi_n_774 ,csa_tree_add_12_51_groupi_n_2393);
  not csa_tree_add_12_51_groupi_drc_bufs24457(csa_tree_add_12_51_groupi_n_773 ,csa_tree_add_12_51_groupi_n_2393);
  not csa_tree_add_12_51_groupi_drc_bufs24460(csa_tree_add_12_51_groupi_n_772 ,csa_tree_add_12_51_groupi_n_770);
  not csa_tree_add_12_51_groupi_drc_bufs24461(csa_tree_add_12_51_groupi_n_771 ,csa_tree_add_12_51_groupi_n_770);
  not csa_tree_add_12_51_groupi_drc_bufs24462(csa_tree_add_12_51_groupi_n_770 ,csa_tree_add_12_51_groupi_n_2311);
  not csa_tree_add_12_51_groupi_drc_bufs24464(csa_tree_add_12_51_groupi_n_769 ,csa_tree_add_12_51_groupi_n_2391);
  not csa_tree_add_12_51_groupi_drc_bufs24465(csa_tree_add_12_51_groupi_n_768 ,csa_tree_add_12_51_groupi_n_2391);
  not csa_tree_add_12_51_groupi_drc_bufs24468(csa_tree_add_12_51_groupi_n_767 ,csa_tree_add_12_51_groupi_n_765);
  not csa_tree_add_12_51_groupi_drc_bufs24469(csa_tree_add_12_51_groupi_n_766 ,csa_tree_add_12_51_groupi_n_765);
  not csa_tree_add_12_51_groupi_drc_bufs24470(csa_tree_add_12_51_groupi_n_765 ,csa_tree_add_12_51_groupi_n_2302);
  not csa_tree_add_12_51_groupi_drc_bufs24472(csa_tree_add_12_51_groupi_n_764 ,csa_tree_add_12_51_groupi_n_2390);
  not csa_tree_add_12_51_groupi_drc_bufs24473(csa_tree_add_12_51_groupi_n_763 ,csa_tree_add_12_51_groupi_n_2390);
  not csa_tree_add_12_51_groupi_drc_bufs24476(csa_tree_add_12_51_groupi_n_762 ,csa_tree_add_12_51_groupi_n_760);
  not csa_tree_add_12_51_groupi_drc_bufs24477(csa_tree_add_12_51_groupi_n_761 ,csa_tree_add_12_51_groupi_n_760);
  not csa_tree_add_12_51_groupi_drc_bufs24478(csa_tree_add_12_51_groupi_n_760 ,csa_tree_add_12_51_groupi_n_2293);
  not csa_tree_add_12_51_groupi_drc_bufs24480(csa_tree_add_12_51_groupi_n_759 ,csa_tree_add_12_51_groupi_n_2389);
  not csa_tree_add_12_51_groupi_drc_bufs24481(csa_tree_add_12_51_groupi_n_758 ,csa_tree_add_12_51_groupi_n_2389);
  not csa_tree_add_12_51_groupi_drc_bufs24484(csa_tree_add_12_51_groupi_n_757 ,csa_tree_add_12_51_groupi_n_2387);
  not csa_tree_add_12_51_groupi_drc_bufs24485(csa_tree_add_12_51_groupi_n_756 ,csa_tree_add_12_51_groupi_n_2387);
  not csa_tree_add_12_51_groupi_drc_bufs24488(csa_tree_add_12_51_groupi_n_755 ,csa_tree_add_12_51_groupi_n_753);
  not csa_tree_add_12_51_groupi_drc_bufs24489(csa_tree_add_12_51_groupi_n_754 ,csa_tree_add_12_51_groupi_n_753);
  not csa_tree_add_12_51_groupi_drc_bufs24490(csa_tree_add_12_51_groupi_n_753 ,csa_tree_add_12_51_groupi_n_2266);
  not csa_tree_add_12_51_groupi_drc_bufs24492(csa_tree_add_12_51_groupi_n_752 ,csa_tree_add_12_51_groupi_n_2359);
  not csa_tree_add_12_51_groupi_drc_bufs24493(csa_tree_add_12_51_groupi_n_751 ,csa_tree_add_12_51_groupi_n_2359);
  not csa_tree_add_12_51_groupi_drc_bufs24496(csa_tree_add_12_51_groupi_n_750 ,csa_tree_add_12_51_groupi_n_2358);
  not csa_tree_add_12_51_groupi_drc_bufs24497(csa_tree_add_12_51_groupi_n_749 ,csa_tree_add_12_51_groupi_n_2358);
  not csa_tree_add_12_51_groupi_drc_bufs24500(csa_tree_add_12_51_groupi_n_748 ,csa_tree_add_12_51_groupi_n_746);
  not csa_tree_add_12_51_groupi_drc_bufs24501(csa_tree_add_12_51_groupi_n_747 ,csa_tree_add_12_51_groupi_n_746);
  not csa_tree_add_12_51_groupi_drc_bufs24502(csa_tree_add_12_51_groupi_n_746 ,csa_tree_add_12_51_groupi_n_2248);
  not csa_tree_add_12_51_groupi_drc_bufs24504(csa_tree_add_12_51_groupi_n_745 ,csa_tree_add_12_51_groupi_n_743);
  not csa_tree_add_12_51_groupi_drc_bufs24505(csa_tree_add_12_51_groupi_n_744 ,csa_tree_add_12_51_groupi_n_743);
  not csa_tree_add_12_51_groupi_drc_bufs24506(csa_tree_add_12_51_groupi_n_743 ,csa_tree_add_12_51_groupi_n_2239);
  not csa_tree_add_12_51_groupi_drc_bufs24508(csa_tree_add_12_51_groupi_n_742 ,csa_tree_add_12_51_groupi_n_2356);
  not csa_tree_add_12_51_groupi_drc_bufs24509(csa_tree_add_12_51_groupi_n_741 ,csa_tree_add_12_51_groupi_n_2356);
  not csa_tree_add_12_51_groupi_drc_bufs24512(csa_tree_add_12_51_groupi_n_740 ,csa_tree_add_12_51_groupi_n_738);
  not csa_tree_add_12_51_groupi_drc_bufs24513(csa_tree_add_12_51_groupi_n_739 ,csa_tree_add_12_51_groupi_n_738);
  not csa_tree_add_12_51_groupi_drc_bufs24514(csa_tree_add_12_51_groupi_n_738 ,csa_tree_add_12_51_groupi_n_2230);
  not csa_tree_add_12_51_groupi_drc_bufs24516(csa_tree_add_12_51_groupi_n_737 ,csa_tree_add_12_51_groupi_n_735);
  not csa_tree_add_12_51_groupi_drc_bufs24517(csa_tree_add_12_51_groupi_n_736 ,csa_tree_add_12_51_groupi_n_735);
  not csa_tree_add_12_51_groupi_drc_bufs24518(csa_tree_add_12_51_groupi_n_735 ,csa_tree_add_12_51_groupi_n_2221);
  not csa_tree_add_12_51_groupi_drc_bufs24520(csa_tree_add_12_51_groupi_n_734 ,csa_tree_add_12_51_groupi_n_2396);
  not csa_tree_add_12_51_groupi_drc_bufs24521(csa_tree_add_12_51_groupi_n_733 ,csa_tree_add_12_51_groupi_n_2396);
  not csa_tree_add_12_51_groupi_drc_bufs24524(csa_tree_add_12_51_groupi_n_732 ,csa_tree_add_12_51_groupi_n_730);
  not csa_tree_add_12_51_groupi_drc_bufs24525(csa_tree_add_12_51_groupi_n_731 ,csa_tree_add_12_51_groupi_n_730);
  not csa_tree_add_12_51_groupi_drc_bufs24526(csa_tree_add_12_51_groupi_n_730 ,csa_tree_add_12_51_groupi_n_2212);
  not csa_tree_add_12_51_groupi_drc_bufs24528(csa_tree_add_12_51_groupi_n_729 ,csa_tree_add_12_51_groupi_n_727);
  not csa_tree_add_12_51_groupi_drc_bufs24529(csa_tree_add_12_51_groupi_n_728 ,csa_tree_add_12_51_groupi_n_727);
  not csa_tree_add_12_51_groupi_drc_bufs24530(csa_tree_add_12_51_groupi_n_727 ,csa_tree_add_12_51_groupi_n_2203);
  not csa_tree_add_12_51_groupi_drc_bufs24532(csa_tree_add_12_51_groupi_n_726 ,csa_tree_add_12_51_groupi_n_2392);
  not csa_tree_add_12_51_groupi_drc_bufs24533(csa_tree_add_12_51_groupi_n_725 ,csa_tree_add_12_51_groupi_n_2392);
  not csa_tree_add_12_51_groupi_drc_bufs24536(csa_tree_add_12_51_groupi_n_724 ,csa_tree_add_12_51_groupi_n_722);
  not csa_tree_add_12_51_groupi_drc_bufs24537(csa_tree_add_12_51_groupi_n_723 ,csa_tree_add_12_51_groupi_n_722);
  not csa_tree_add_12_51_groupi_drc_bufs24538(csa_tree_add_12_51_groupi_n_722 ,csa_tree_add_12_51_groupi_n_2338);
  not csa_tree_add_12_51_groupi_drc_bufs24540(csa_tree_add_12_51_groupi_n_721 ,csa_tree_add_12_51_groupi_n_719);
  not csa_tree_add_12_51_groupi_drc_bufs24541(csa_tree_add_12_51_groupi_n_720 ,csa_tree_add_12_51_groupi_n_719);
  not csa_tree_add_12_51_groupi_drc_bufs24542(csa_tree_add_12_51_groupi_n_719 ,csa_tree_add_12_51_groupi_n_2275);
  not csa_tree_add_12_51_groupi_drc_bufs24544(csa_tree_add_12_51_groupi_n_718 ,csa_tree_add_12_51_groupi_n_716);
  not csa_tree_add_12_51_groupi_drc_bufs24545(csa_tree_add_12_51_groupi_n_717 ,csa_tree_add_12_51_groupi_n_716);
  not csa_tree_add_12_51_groupi_drc_bufs24546(csa_tree_add_12_51_groupi_n_716 ,csa_tree_add_12_51_groupi_n_2257);
  not csa_tree_add_12_51_groupi_drc_bufs24548(csa_tree_add_12_51_groupi_n_715 ,csa_tree_add_12_51_groupi_n_713);
  not csa_tree_add_12_51_groupi_drc_bufs24549(csa_tree_add_12_51_groupi_n_714 ,csa_tree_add_12_51_groupi_n_713);
  not csa_tree_add_12_51_groupi_drc_bufs24550(csa_tree_add_12_51_groupi_n_713 ,csa_tree_add_12_51_groupi_n_2284);
  not csa_tree_add_12_51_groupi_drc_bufs24552(csa_tree_add_12_51_groupi_n_712 ,csa_tree_add_12_51_groupi_n_710);
  not csa_tree_add_12_51_groupi_drc_bufs24553(csa_tree_add_12_51_groupi_n_711 ,csa_tree_add_12_51_groupi_n_710);
  not csa_tree_add_12_51_groupi_drc_bufs24554(csa_tree_add_12_51_groupi_n_710 ,csa_tree_add_12_51_groupi_n_2012);
  not csa_tree_add_12_51_groupi_drc_bufs24556(csa_tree_add_12_51_groupi_n_709 ,csa_tree_add_12_51_groupi_n_707);
  not csa_tree_add_12_51_groupi_drc_bufs24557(csa_tree_add_12_51_groupi_n_708 ,csa_tree_add_12_51_groupi_n_707);
  not csa_tree_add_12_51_groupi_drc_bufs24558(csa_tree_add_12_51_groupi_n_707 ,csa_tree_add_12_51_groupi_n_2010);
  not csa_tree_add_12_51_groupi_drc_bufs24560(csa_tree_add_12_51_groupi_n_706 ,csa_tree_add_12_51_groupi_n_704);
  not csa_tree_add_12_51_groupi_drc_bufs24561(csa_tree_add_12_51_groupi_n_705 ,csa_tree_add_12_51_groupi_n_704);
  not csa_tree_add_12_51_groupi_drc_bufs24562(csa_tree_add_12_51_groupi_n_704 ,csa_tree_add_12_51_groupi_n_2020);
  not csa_tree_add_12_51_groupi_drc_bufs24564(csa_tree_add_12_51_groupi_n_703 ,csa_tree_add_12_51_groupi_n_701);
  not csa_tree_add_12_51_groupi_drc_bufs24565(csa_tree_add_12_51_groupi_n_702 ,csa_tree_add_12_51_groupi_n_701);
  not csa_tree_add_12_51_groupi_drc_bufs24566(csa_tree_add_12_51_groupi_n_701 ,csa_tree_add_12_51_groupi_n_2018);
  not csa_tree_add_12_51_groupi_drc_bufs24568(csa_tree_add_12_51_groupi_n_700 ,csa_tree_add_12_51_groupi_n_698);
  not csa_tree_add_12_51_groupi_drc_bufs24569(csa_tree_add_12_51_groupi_n_699 ,csa_tree_add_12_51_groupi_n_698);
  not csa_tree_add_12_51_groupi_drc_bufs24570(csa_tree_add_12_51_groupi_n_698 ,csa_tree_add_12_51_groupi_n_2208);
  not csa_tree_add_12_51_groupi_drc_bufs24572(csa_tree_add_12_51_groupi_n_697 ,csa_tree_add_12_51_groupi_n_695);
  not csa_tree_add_12_51_groupi_drc_bufs24573(csa_tree_add_12_51_groupi_n_696 ,csa_tree_add_12_51_groupi_n_695);
  not csa_tree_add_12_51_groupi_drc_bufs24574(csa_tree_add_12_51_groupi_n_695 ,csa_tree_add_12_51_groupi_n_2218);
  not csa_tree_add_12_51_groupi_drc_bufs24576(csa_tree_add_12_51_groupi_n_694 ,csa_tree_add_12_51_groupi_n_692);
  not csa_tree_add_12_51_groupi_drc_bufs24577(csa_tree_add_12_51_groupi_n_693 ,csa_tree_add_12_51_groupi_n_692);
  not csa_tree_add_12_51_groupi_drc_bufs24578(csa_tree_add_12_51_groupi_n_692 ,csa_tree_add_12_51_groupi_n_2220);
  not csa_tree_add_12_51_groupi_drc_bufs24580(csa_tree_add_12_51_groupi_n_691 ,csa_tree_add_12_51_groupi_n_689);
  not csa_tree_add_12_51_groupi_drc_bufs24581(csa_tree_add_12_51_groupi_n_690 ,csa_tree_add_12_51_groupi_n_689);
  not csa_tree_add_12_51_groupi_drc_bufs24582(csa_tree_add_12_51_groupi_n_689 ,csa_tree_add_12_51_groupi_n_2252);
  not csa_tree_add_12_51_groupi_drc_bufs24584(csa_tree_add_12_51_groupi_n_688 ,csa_tree_add_12_51_groupi_n_686);
  not csa_tree_add_12_51_groupi_drc_bufs24585(csa_tree_add_12_51_groupi_n_687 ,csa_tree_add_12_51_groupi_n_686);
  not csa_tree_add_12_51_groupi_drc_bufs24586(csa_tree_add_12_51_groupi_n_686 ,csa_tree_add_12_51_groupi_n_2271);
  not csa_tree_add_12_51_groupi_drc_bufs24588(csa_tree_add_12_51_groupi_n_685 ,csa_tree_add_12_51_groupi_n_683);
  not csa_tree_add_12_51_groupi_drc_bufs24589(csa_tree_add_12_51_groupi_n_684 ,csa_tree_add_12_51_groupi_n_683);
  not csa_tree_add_12_51_groupi_drc_bufs24590(csa_tree_add_12_51_groupi_n_683 ,csa_tree_add_12_51_groupi_n_2262);
  not csa_tree_add_12_51_groupi_drc_bufs24592(csa_tree_add_12_51_groupi_n_682 ,csa_tree_add_12_51_groupi_n_680);
  not csa_tree_add_12_51_groupi_drc_bufs24593(csa_tree_add_12_51_groupi_n_681 ,csa_tree_add_12_51_groupi_n_680);
  not csa_tree_add_12_51_groupi_drc_bufs24594(csa_tree_add_12_51_groupi_n_680 ,csa_tree_add_12_51_groupi_n_2270);
  not csa_tree_add_12_51_groupi_drc_bufs24596(csa_tree_add_12_51_groupi_n_679 ,csa_tree_add_12_51_groupi_n_677);
  not csa_tree_add_12_51_groupi_drc_bufs24597(csa_tree_add_12_51_groupi_n_678 ,csa_tree_add_12_51_groupi_n_677);
  not csa_tree_add_12_51_groupi_drc_bufs24598(csa_tree_add_12_51_groupi_n_677 ,csa_tree_add_12_51_groupi_n_2344);
  not csa_tree_add_12_51_groupi_drc_bufs24600(csa_tree_add_12_51_groupi_n_676 ,csa_tree_add_12_51_groupi_n_674);
  not csa_tree_add_12_51_groupi_drc_bufs24601(csa_tree_add_12_51_groupi_n_675 ,csa_tree_add_12_51_groupi_n_674);
  not csa_tree_add_12_51_groupi_drc_bufs24602(csa_tree_add_12_51_groupi_n_674 ,csa_tree_add_12_51_groupi_n_2261);
  not csa_tree_add_12_51_groupi_drc_bufs24604(csa_tree_add_12_51_groupi_n_673 ,csa_tree_add_12_51_groupi_n_671);
  not csa_tree_add_12_51_groupi_drc_bufs24605(csa_tree_add_12_51_groupi_n_672 ,csa_tree_add_12_51_groupi_n_671);
  not csa_tree_add_12_51_groupi_drc_bufs24606(csa_tree_add_12_51_groupi_n_671 ,csa_tree_add_12_51_groupi_n_2246);
  not csa_tree_add_12_51_groupi_drc_bufs24608(csa_tree_add_12_51_groupi_n_670 ,csa_tree_add_12_51_groupi_n_668);
  not csa_tree_add_12_51_groupi_drc_bufs24609(csa_tree_add_12_51_groupi_n_669 ,csa_tree_add_12_51_groupi_n_668);
  not csa_tree_add_12_51_groupi_drc_bufs24610(csa_tree_add_12_51_groupi_n_668 ,csa_tree_add_12_51_groupi_n_2238);
  not csa_tree_add_12_51_groupi_drc_bufs24612(csa_tree_add_12_51_groupi_n_667 ,csa_tree_add_12_51_groupi_n_665);
  not csa_tree_add_12_51_groupi_drc_bufs24613(csa_tree_add_12_51_groupi_n_666 ,csa_tree_add_12_51_groupi_n_665);
  not csa_tree_add_12_51_groupi_drc_bufs24614(csa_tree_add_12_51_groupi_n_665 ,csa_tree_add_12_51_groupi_n_2343);
  not csa_tree_add_12_51_groupi_drc_bufs24616(csa_tree_add_12_51_groupi_n_664 ,csa_tree_add_12_51_groupi_n_662);
  not csa_tree_add_12_51_groupi_drc_bufs24617(csa_tree_add_12_51_groupi_n_663 ,csa_tree_add_12_51_groupi_n_662);
  not csa_tree_add_12_51_groupi_drc_bufs24618(csa_tree_add_12_51_groupi_n_662 ,csa_tree_add_12_51_groupi_n_2337);
  not csa_tree_add_12_51_groupi_drc_bufs24620(csa_tree_add_12_51_groupi_n_661 ,csa_tree_add_12_51_groupi_n_659);
  not csa_tree_add_12_51_groupi_drc_bufs24621(csa_tree_add_12_51_groupi_n_660 ,csa_tree_add_12_51_groupi_n_659);
  not csa_tree_add_12_51_groupi_drc_bufs24622(csa_tree_add_12_51_groupi_n_659 ,csa_tree_add_12_51_groupi_n_2298);
  not csa_tree_add_12_51_groupi_drc_bufs24624(csa_tree_add_12_51_groupi_n_658 ,csa_tree_add_12_51_groupi_n_656);
  not csa_tree_add_12_51_groupi_drc_bufs24625(csa_tree_add_12_51_groupi_n_657 ,csa_tree_add_12_51_groupi_n_656);
  not csa_tree_add_12_51_groupi_drc_bufs24626(csa_tree_add_12_51_groupi_n_656 ,csa_tree_add_12_51_groupi_n_2336);
  not csa_tree_add_12_51_groupi_drc_bufs24628(csa_tree_add_12_51_groupi_n_655 ,csa_tree_add_12_51_groupi_n_653);
  not csa_tree_add_12_51_groupi_drc_bufs24629(csa_tree_add_12_51_groupi_n_654 ,csa_tree_add_12_51_groupi_n_653);
  not csa_tree_add_12_51_groupi_drc_bufs24630(csa_tree_add_12_51_groupi_n_653 ,csa_tree_add_12_51_groupi_n_2328);
  not csa_tree_add_12_51_groupi_drc_bufs24632(csa_tree_add_12_51_groupi_n_652 ,csa_tree_add_12_51_groupi_n_650);
  not csa_tree_add_12_51_groupi_drc_bufs24633(csa_tree_add_12_51_groupi_n_651 ,csa_tree_add_12_51_groupi_n_650);
  not csa_tree_add_12_51_groupi_drc_bufs24634(csa_tree_add_12_51_groupi_n_650 ,csa_tree_add_12_51_groupi_n_2327);
  not csa_tree_add_12_51_groupi_drc_bufs24636(csa_tree_add_12_51_groupi_n_649 ,csa_tree_add_12_51_groupi_n_647);
  not csa_tree_add_12_51_groupi_drc_bufs24637(csa_tree_add_12_51_groupi_n_648 ,csa_tree_add_12_51_groupi_n_647);
  not csa_tree_add_12_51_groupi_drc_bufs24638(csa_tree_add_12_51_groupi_n_647 ,csa_tree_add_12_51_groupi_n_2326);
  not csa_tree_add_12_51_groupi_drc_bufs24640(csa_tree_add_12_51_groupi_n_646 ,csa_tree_add_12_51_groupi_n_644);
  not csa_tree_add_12_51_groupi_drc_bufs24641(csa_tree_add_12_51_groupi_n_645 ,csa_tree_add_12_51_groupi_n_644);
  not csa_tree_add_12_51_groupi_drc_bufs24642(csa_tree_add_12_51_groupi_n_644 ,csa_tree_add_12_51_groupi_n_2346);
  not csa_tree_add_12_51_groupi_drc_bufs24644(csa_tree_add_12_51_groupi_n_643 ,csa_tree_add_12_51_groupi_n_641);
  not csa_tree_add_12_51_groupi_drc_bufs24645(csa_tree_add_12_51_groupi_n_642 ,csa_tree_add_12_51_groupi_n_641);
  not csa_tree_add_12_51_groupi_drc_bufs24646(csa_tree_add_12_51_groupi_n_641 ,csa_tree_add_12_51_groupi_n_2319);
  not csa_tree_add_12_51_groupi_drc_bufs24648(csa_tree_add_12_51_groupi_n_640 ,csa_tree_add_12_51_groupi_n_638);
  not csa_tree_add_12_51_groupi_drc_bufs24649(csa_tree_add_12_51_groupi_n_639 ,csa_tree_add_12_51_groupi_n_638);
  not csa_tree_add_12_51_groupi_drc_bufs24650(csa_tree_add_12_51_groupi_n_638 ,csa_tree_add_12_51_groupi_n_2318);
  not csa_tree_add_12_51_groupi_drc_bufs24652(csa_tree_add_12_51_groupi_n_637 ,csa_tree_add_12_51_groupi_n_635);
  not csa_tree_add_12_51_groupi_drc_bufs24653(csa_tree_add_12_51_groupi_n_636 ,csa_tree_add_12_51_groupi_n_635);
  not csa_tree_add_12_51_groupi_drc_bufs24654(csa_tree_add_12_51_groupi_n_635 ,csa_tree_add_12_51_groupi_n_2317);
  not csa_tree_add_12_51_groupi_drc_bufs24656(csa_tree_add_12_51_groupi_n_634 ,csa_tree_add_12_51_groupi_n_632);
  not csa_tree_add_12_51_groupi_drc_bufs24657(csa_tree_add_12_51_groupi_n_633 ,csa_tree_add_12_51_groupi_n_632);
  not csa_tree_add_12_51_groupi_drc_bufs24658(csa_tree_add_12_51_groupi_n_632 ,csa_tree_add_12_51_groupi_n_2345);
  not csa_tree_add_12_51_groupi_drc_bufs24660(csa_tree_add_12_51_groupi_n_631 ,csa_tree_add_12_51_groupi_n_629);
  not csa_tree_add_12_51_groupi_drc_bufs24661(csa_tree_add_12_51_groupi_n_630 ,csa_tree_add_12_51_groupi_n_629);
  not csa_tree_add_12_51_groupi_drc_bufs24662(csa_tree_add_12_51_groupi_n_629 ,csa_tree_add_12_51_groupi_n_2310);
  not csa_tree_add_12_51_groupi_drc_bufs24664(csa_tree_add_12_51_groupi_n_628 ,csa_tree_add_12_51_groupi_n_626);
  not csa_tree_add_12_51_groupi_drc_bufs24665(csa_tree_add_12_51_groupi_n_627 ,csa_tree_add_12_51_groupi_n_626);
  not csa_tree_add_12_51_groupi_drc_bufs24666(csa_tree_add_12_51_groupi_n_626 ,csa_tree_add_12_51_groupi_n_2253);
  not csa_tree_add_12_51_groupi_drc_bufs24668(csa_tree_add_12_51_groupi_n_625 ,csa_tree_add_12_51_groupi_n_623);
  not csa_tree_add_12_51_groupi_drc_bufs24669(csa_tree_add_12_51_groupi_n_624 ,csa_tree_add_12_51_groupi_n_623);
  not csa_tree_add_12_51_groupi_drc_bufs24670(csa_tree_add_12_51_groupi_n_623 ,csa_tree_add_12_51_groupi_n_2255);
  not csa_tree_add_12_51_groupi_drc_bufs24672(csa_tree_add_12_51_groupi_n_622 ,csa_tree_add_12_51_groupi_n_620);
  not csa_tree_add_12_51_groupi_drc_bufs24673(csa_tree_add_12_51_groupi_n_621 ,csa_tree_add_12_51_groupi_n_620);
  not csa_tree_add_12_51_groupi_drc_bufs24674(csa_tree_add_12_51_groupi_n_620 ,csa_tree_add_12_51_groupi_n_2289);
  not csa_tree_add_12_51_groupi_drc_bufs24676(csa_tree_add_12_51_groupi_n_619 ,csa_tree_add_12_51_groupi_n_617);
  not csa_tree_add_12_51_groupi_drc_bufs24677(csa_tree_add_12_51_groupi_n_618 ,csa_tree_add_12_51_groupi_n_617);
  not csa_tree_add_12_51_groupi_drc_bufs24678(csa_tree_add_12_51_groupi_n_617 ,csa_tree_add_12_51_groupi_n_2309);
  not csa_tree_add_12_51_groupi_drc_bufs24680(csa_tree_add_12_51_groupi_n_616 ,csa_tree_add_12_51_groupi_n_614);
  not csa_tree_add_12_51_groupi_drc_bufs24681(csa_tree_add_12_51_groupi_n_615 ,csa_tree_add_12_51_groupi_n_614);
  not csa_tree_add_12_51_groupi_drc_bufs24682(csa_tree_add_12_51_groupi_n_614 ,csa_tree_add_12_51_groupi_n_2308);
  not csa_tree_add_12_51_groupi_drc_bufs24684(csa_tree_add_12_51_groupi_n_613 ,csa_tree_add_12_51_groupi_n_611);
  not csa_tree_add_12_51_groupi_drc_bufs24685(csa_tree_add_12_51_groupi_n_612 ,csa_tree_add_12_51_groupi_n_611);
  not csa_tree_add_12_51_groupi_drc_bufs24686(csa_tree_add_12_51_groupi_n_611 ,csa_tree_add_12_51_groupi_n_2265);
  not csa_tree_add_12_51_groupi_drc_bufs24688(csa_tree_add_12_51_groupi_n_610 ,csa_tree_add_12_51_groupi_n_608);
  not csa_tree_add_12_51_groupi_drc_bufs24689(csa_tree_add_12_51_groupi_n_609 ,csa_tree_add_12_51_groupi_n_608);
  not csa_tree_add_12_51_groupi_drc_bufs24690(csa_tree_add_12_51_groupi_n_608 ,csa_tree_add_12_51_groupi_n_2300);
  not csa_tree_add_12_51_groupi_drc_bufs24692(csa_tree_add_12_51_groupi_n_607 ,csa_tree_add_12_51_groupi_n_605);
  not csa_tree_add_12_51_groupi_drc_bufs24693(csa_tree_add_12_51_groupi_n_606 ,csa_tree_add_12_51_groupi_n_605);
  not csa_tree_add_12_51_groupi_drc_bufs24694(csa_tree_add_12_51_groupi_n_605 ,csa_tree_add_12_51_groupi_n_2273);
  not csa_tree_add_12_51_groupi_drc_bufs24696(csa_tree_add_12_51_groupi_n_604 ,csa_tree_add_12_51_groupi_n_602);
  not csa_tree_add_12_51_groupi_drc_bufs24697(csa_tree_add_12_51_groupi_n_603 ,csa_tree_add_12_51_groupi_n_602);
  not csa_tree_add_12_51_groupi_drc_bufs24698(csa_tree_add_12_51_groupi_n_602 ,csa_tree_add_12_51_groupi_n_2301);
  not csa_tree_add_12_51_groupi_drc_bufs24700(csa_tree_add_12_51_groupi_n_601 ,csa_tree_add_12_51_groupi_n_599);
  not csa_tree_add_12_51_groupi_drc_bufs24701(csa_tree_add_12_51_groupi_n_600 ,csa_tree_add_12_51_groupi_n_599);
  not csa_tree_add_12_51_groupi_drc_bufs24702(csa_tree_add_12_51_groupi_n_599 ,csa_tree_add_12_51_groupi_n_2256);
  not csa_tree_add_12_51_groupi_drc_bufs24704(csa_tree_add_12_51_groupi_n_598 ,csa_tree_add_12_51_groupi_n_596);
  not csa_tree_add_12_51_groupi_drc_bufs24705(csa_tree_add_12_51_groupi_n_597 ,csa_tree_add_12_51_groupi_n_596);
  not csa_tree_add_12_51_groupi_drc_bufs24706(csa_tree_add_12_51_groupi_n_596 ,csa_tree_add_12_51_groupi_n_2292);
  not csa_tree_add_12_51_groupi_drc_bufs24708(csa_tree_add_12_51_groupi_n_595 ,csa_tree_add_12_51_groupi_n_593);
  not csa_tree_add_12_51_groupi_drc_bufs24709(csa_tree_add_12_51_groupi_n_594 ,csa_tree_add_12_51_groupi_n_593);
  not csa_tree_add_12_51_groupi_drc_bufs24710(csa_tree_add_12_51_groupi_n_593 ,csa_tree_add_12_51_groupi_n_2291);
  not csa_tree_add_12_51_groupi_drc_bufs24712(csa_tree_add_12_51_groupi_n_592 ,csa_tree_add_12_51_groupi_n_590);
  not csa_tree_add_12_51_groupi_drc_bufs24713(csa_tree_add_12_51_groupi_n_591 ,csa_tree_add_12_51_groupi_n_590);
  not csa_tree_add_12_51_groupi_drc_bufs24714(csa_tree_add_12_51_groupi_n_590 ,csa_tree_add_12_51_groupi_n_2283);
  not csa_tree_add_12_51_groupi_drc_bufs24716(csa_tree_add_12_51_groupi_n_589 ,csa_tree_add_12_51_groupi_n_587);
  not csa_tree_add_12_51_groupi_drc_bufs24717(csa_tree_add_12_51_groupi_n_588 ,csa_tree_add_12_51_groupi_n_587);
  not csa_tree_add_12_51_groupi_drc_bufs24718(csa_tree_add_12_51_groupi_n_587 ,csa_tree_add_12_51_groupi_n_2282);
  not csa_tree_add_12_51_groupi_drc_bufs24720(csa_tree_add_12_51_groupi_n_586 ,csa_tree_add_12_51_groupi_n_584);
  not csa_tree_add_12_51_groupi_drc_bufs24721(csa_tree_add_12_51_groupi_n_585 ,csa_tree_add_12_51_groupi_n_584);
  not csa_tree_add_12_51_groupi_drc_bufs24722(csa_tree_add_12_51_groupi_n_584 ,csa_tree_add_12_51_groupi_n_2281);
  not csa_tree_add_12_51_groupi_drc_bufs24724(csa_tree_add_12_51_groupi_n_583 ,csa_tree_add_12_51_groupi_n_581);
  not csa_tree_add_12_51_groupi_drc_bufs24725(csa_tree_add_12_51_groupi_n_582 ,csa_tree_add_12_51_groupi_n_581);
  not csa_tree_add_12_51_groupi_drc_bufs24726(csa_tree_add_12_51_groupi_n_581 ,csa_tree_add_12_51_groupi_n_2288);
  not csa_tree_add_12_51_groupi_drc_bufs24728(csa_tree_add_12_51_groupi_n_580 ,csa_tree_add_12_51_groupi_n_578);
  not csa_tree_add_12_51_groupi_drc_bufs24729(csa_tree_add_12_51_groupi_n_579 ,csa_tree_add_12_51_groupi_n_578);
  not csa_tree_add_12_51_groupi_drc_bufs24730(csa_tree_add_12_51_groupi_n_578 ,csa_tree_add_12_51_groupi_n_2272);
  not csa_tree_add_12_51_groupi_drc_bufs24732(csa_tree_add_12_51_groupi_n_577 ,csa_tree_add_12_51_groupi_n_575);
  not csa_tree_add_12_51_groupi_drc_bufs24733(csa_tree_add_12_51_groupi_n_576 ,csa_tree_add_12_51_groupi_n_575);
  not csa_tree_add_12_51_groupi_drc_bufs24734(csa_tree_add_12_51_groupi_n_575 ,csa_tree_add_12_51_groupi_n_2264);
  not csa_tree_add_12_51_groupi_drc_bufs24736(csa_tree_add_12_51_groupi_n_574 ,csa_tree_add_12_51_groupi_n_572);
  not csa_tree_add_12_51_groupi_drc_bufs24737(csa_tree_add_12_51_groupi_n_573 ,csa_tree_add_12_51_groupi_n_572);
  not csa_tree_add_12_51_groupi_drc_bufs24738(csa_tree_add_12_51_groupi_n_572 ,csa_tree_add_12_51_groupi_n_2263);
  not csa_tree_add_12_51_groupi_drc_bufs24740(csa_tree_add_12_51_groupi_n_571 ,csa_tree_add_12_51_groupi_n_569);
  not csa_tree_add_12_51_groupi_drc_bufs24741(csa_tree_add_12_51_groupi_n_570 ,csa_tree_add_12_51_groupi_n_569);
  not csa_tree_add_12_51_groupi_drc_bufs24742(csa_tree_add_12_51_groupi_n_569 ,csa_tree_add_12_51_groupi_n_2297);
  not csa_tree_add_12_51_groupi_drc_bufs24744(csa_tree_add_12_51_groupi_n_568 ,csa_tree_add_12_51_groupi_n_566);
  not csa_tree_add_12_51_groupi_drc_bufs24745(csa_tree_add_12_51_groupi_n_567 ,csa_tree_add_12_51_groupi_n_566);
  not csa_tree_add_12_51_groupi_drc_bufs24746(csa_tree_add_12_51_groupi_n_566 ,csa_tree_add_12_51_groupi_n_2254);
  not csa_tree_add_12_51_groupi_drc_bufs24748(csa_tree_add_12_51_groupi_n_565 ,csa_tree_add_12_51_groupi_n_563);
  not csa_tree_add_12_51_groupi_drc_bufs24749(csa_tree_add_12_51_groupi_n_564 ,csa_tree_add_12_51_groupi_n_563);
  not csa_tree_add_12_51_groupi_drc_bufs24750(csa_tree_add_12_51_groupi_n_563 ,csa_tree_add_12_51_groupi_n_2274);
  not csa_tree_add_12_51_groupi_drc_bufs24752(csa_tree_add_12_51_groupi_n_562 ,csa_tree_add_12_51_groupi_n_560);
  not csa_tree_add_12_51_groupi_drc_bufs24753(csa_tree_add_12_51_groupi_n_561 ,csa_tree_add_12_51_groupi_n_560);
  not csa_tree_add_12_51_groupi_drc_bufs24754(csa_tree_add_12_51_groupi_n_560 ,csa_tree_add_12_51_groupi_n_2247);
  not csa_tree_add_12_51_groupi_drc_bufs24756(csa_tree_add_12_51_groupi_n_559 ,csa_tree_add_12_51_groupi_n_557);
  not csa_tree_add_12_51_groupi_drc_bufs24757(csa_tree_add_12_51_groupi_n_558 ,csa_tree_add_12_51_groupi_n_557);
  not csa_tree_add_12_51_groupi_drc_bufs24758(csa_tree_add_12_51_groupi_n_557 ,csa_tree_add_12_51_groupi_n_2245);
  not csa_tree_add_12_51_groupi_drc_bufs24760(csa_tree_add_12_51_groupi_n_556 ,csa_tree_add_12_51_groupi_n_554);
  not csa_tree_add_12_51_groupi_drc_bufs24761(csa_tree_add_12_51_groupi_n_555 ,csa_tree_add_12_51_groupi_n_554);
  not csa_tree_add_12_51_groupi_drc_bufs24762(csa_tree_add_12_51_groupi_n_554 ,csa_tree_add_12_51_groupi_n_2237);
  not csa_tree_add_12_51_groupi_drc_bufs24764(csa_tree_add_12_51_groupi_n_553 ,csa_tree_add_12_51_groupi_n_551);
  not csa_tree_add_12_51_groupi_drc_bufs24765(csa_tree_add_12_51_groupi_n_552 ,csa_tree_add_12_51_groupi_n_551);
  not csa_tree_add_12_51_groupi_drc_bufs24766(csa_tree_add_12_51_groupi_n_551 ,csa_tree_add_12_51_groupi_n_2324);
  not csa_tree_add_12_51_groupi_drc_bufs24768(csa_tree_add_12_51_groupi_n_550 ,csa_tree_add_12_51_groupi_n_548);
  not csa_tree_add_12_51_groupi_drc_bufs24769(csa_tree_add_12_51_groupi_n_549 ,csa_tree_add_12_51_groupi_n_548);
  not csa_tree_add_12_51_groupi_drc_bufs24770(csa_tree_add_12_51_groupi_n_548 ,csa_tree_add_12_51_groupi_n_2236);
  not csa_tree_add_12_51_groupi_drc_bufs24772(csa_tree_add_12_51_groupi_n_547 ,csa_tree_add_12_51_groupi_n_545);
  not csa_tree_add_12_51_groupi_drc_bufs24773(csa_tree_add_12_51_groupi_n_546 ,csa_tree_add_12_51_groupi_n_545);
  not csa_tree_add_12_51_groupi_drc_bufs24774(csa_tree_add_12_51_groupi_n_545 ,csa_tree_add_12_51_groupi_n_2307);
  not csa_tree_add_12_51_groupi_drc_bufs24776(csa_tree_add_12_51_groupi_n_544 ,csa_tree_add_12_51_groupi_n_542);
  not csa_tree_add_12_51_groupi_drc_bufs24777(csa_tree_add_12_51_groupi_n_543 ,csa_tree_add_12_51_groupi_n_542);
  not csa_tree_add_12_51_groupi_drc_bufs24778(csa_tree_add_12_51_groupi_n_542 ,csa_tree_add_12_51_groupi_n_2229);
  not csa_tree_add_12_51_groupi_drc_bufs24780(csa_tree_add_12_51_groupi_n_541 ,csa_tree_add_12_51_groupi_n_539);
  not csa_tree_add_12_51_groupi_drc_bufs24781(csa_tree_add_12_51_groupi_n_540 ,csa_tree_add_12_51_groupi_n_539);
  not csa_tree_add_12_51_groupi_drc_bufs24782(csa_tree_add_12_51_groupi_n_539 ,csa_tree_add_12_51_groupi_n_2228);
  not csa_tree_add_12_51_groupi_drc_bufs24784(csa_tree_add_12_51_groupi_n_538 ,csa_tree_add_12_51_groupi_n_536);
  not csa_tree_add_12_51_groupi_drc_bufs24785(csa_tree_add_12_51_groupi_n_537 ,csa_tree_add_12_51_groupi_n_536);
  not csa_tree_add_12_51_groupi_drc_bufs24786(csa_tree_add_12_51_groupi_n_536 ,csa_tree_add_12_51_groupi_n_2227);
  not csa_tree_add_12_51_groupi_drc_bufs24788(csa_tree_add_12_51_groupi_n_535 ,csa_tree_add_12_51_groupi_n_533);
  not csa_tree_add_12_51_groupi_drc_bufs24789(csa_tree_add_12_51_groupi_n_534 ,csa_tree_add_12_51_groupi_n_533);
  not csa_tree_add_12_51_groupi_drc_bufs24790(csa_tree_add_12_51_groupi_n_533 ,csa_tree_add_12_51_groupi_n_2234);
  not csa_tree_add_12_51_groupi_drc_bufs24792(csa_tree_add_12_51_groupi_n_532 ,csa_tree_add_12_51_groupi_n_530);
  not csa_tree_add_12_51_groupi_drc_bufs24793(csa_tree_add_12_51_groupi_n_531 ,csa_tree_add_12_51_groupi_n_530);
  not csa_tree_add_12_51_groupi_drc_bufs24794(csa_tree_add_12_51_groupi_n_530 ,csa_tree_add_12_51_groupi_n_2335);
  not csa_tree_add_12_51_groupi_drc_bufs24796(csa_tree_add_12_51_groupi_n_529 ,csa_tree_add_12_51_groupi_n_527);
  not csa_tree_add_12_51_groupi_drc_bufs24797(csa_tree_add_12_51_groupi_n_528 ,csa_tree_add_12_51_groupi_n_527);
  not csa_tree_add_12_51_groupi_drc_bufs24798(csa_tree_add_12_51_groupi_n_527 ,csa_tree_add_12_51_groupi_n_2290);
  not csa_tree_add_12_51_groupi_drc_bufs24800(csa_tree_add_12_51_groupi_n_526 ,csa_tree_add_12_51_groupi_n_524);
  not csa_tree_add_12_51_groupi_drc_bufs24801(csa_tree_add_12_51_groupi_n_525 ,csa_tree_add_12_51_groupi_n_524);
  not csa_tree_add_12_51_groupi_drc_bufs24802(csa_tree_add_12_51_groupi_n_524 ,csa_tree_add_12_51_groupi_n_2334);
  not csa_tree_add_12_51_groupi_drc_bufs24804(csa_tree_add_12_51_groupi_n_523 ,csa_tree_add_12_51_groupi_n_521);
  not csa_tree_add_12_51_groupi_drc_bufs24805(csa_tree_add_12_51_groupi_n_522 ,csa_tree_add_12_51_groupi_n_521);
  not csa_tree_add_12_51_groupi_drc_bufs24806(csa_tree_add_12_51_groupi_n_521 ,csa_tree_add_12_51_groupi_n_2306);
  not csa_tree_add_12_51_groupi_drc_bufs24808(csa_tree_add_12_51_groupi_n_520 ,csa_tree_add_12_51_groupi_n_518);
  not csa_tree_add_12_51_groupi_drc_bufs24809(csa_tree_add_12_51_groupi_n_519 ,csa_tree_add_12_51_groupi_n_518);
  not csa_tree_add_12_51_groupi_drc_bufs24810(csa_tree_add_12_51_groupi_n_518 ,csa_tree_add_12_51_groupi_n_2316);
  not csa_tree_add_12_51_groupi_drc_bufs24812(csa_tree_add_12_51_groupi_n_517 ,csa_tree_add_12_51_groupi_n_515);
  not csa_tree_add_12_51_groupi_drc_bufs24813(csa_tree_add_12_51_groupi_n_516 ,csa_tree_add_12_51_groupi_n_515);
  not csa_tree_add_12_51_groupi_drc_bufs24814(csa_tree_add_12_51_groupi_n_515 ,csa_tree_add_12_51_groupi_n_2226);
  not csa_tree_add_12_51_groupi_drc_bufs24816(csa_tree_add_12_51_groupi_n_514 ,csa_tree_add_12_51_groupi_n_512);
  not csa_tree_add_12_51_groupi_drc_bufs24817(csa_tree_add_12_51_groupi_n_513 ,csa_tree_add_12_51_groupi_n_512);
  not csa_tree_add_12_51_groupi_drc_bufs24818(csa_tree_add_12_51_groupi_n_512 ,csa_tree_add_12_51_groupi_n_2299);
  not csa_tree_add_12_51_groupi_drc_bufs24820(csa_tree_add_12_51_groupi_n_511 ,csa_tree_add_12_51_groupi_n_509);
  not csa_tree_add_12_51_groupi_drc_bufs24821(csa_tree_add_12_51_groupi_n_510 ,csa_tree_add_12_51_groupi_n_509);
  not csa_tree_add_12_51_groupi_drc_bufs24822(csa_tree_add_12_51_groupi_n_509 ,csa_tree_add_12_51_groupi_n_2280);
  not csa_tree_add_12_51_groupi_drc_bufs24824(csa_tree_add_12_51_groupi_n_508 ,csa_tree_add_12_51_groupi_n_506);
  not csa_tree_add_12_51_groupi_drc_bufs24825(csa_tree_add_12_51_groupi_n_507 ,csa_tree_add_12_51_groupi_n_506);
  not csa_tree_add_12_51_groupi_drc_bufs24826(csa_tree_add_12_51_groupi_n_506 ,csa_tree_add_12_51_groupi_n_2279);
  not csa_tree_add_12_51_groupi_drc_bufs24828(csa_tree_add_12_51_groupi_n_505 ,csa_tree_add_12_51_groupi_n_503);
  not csa_tree_add_12_51_groupi_drc_bufs24829(csa_tree_add_12_51_groupi_n_504 ,csa_tree_add_12_51_groupi_n_503);
  not csa_tree_add_12_51_groupi_drc_bufs24830(csa_tree_add_12_51_groupi_n_503 ,csa_tree_add_12_51_groupi_n_2219);
  not csa_tree_add_12_51_groupi_drc_bufs24832(csa_tree_add_12_51_groupi_n_502 ,csa_tree_add_12_51_groupi_n_500);
  not csa_tree_add_12_51_groupi_drc_bufs24833(csa_tree_add_12_51_groupi_n_501 ,csa_tree_add_12_51_groupi_n_500);
  not csa_tree_add_12_51_groupi_drc_bufs24834(csa_tree_add_12_51_groupi_n_500 ,csa_tree_add_12_51_groupi_n_2315);
  not csa_tree_add_12_51_groupi_drc_bufs24836(csa_tree_add_12_51_groupi_n_499 ,csa_tree_add_12_51_groupi_n_497);
  not csa_tree_add_12_51_groupi_drc_bufs24837(csa_tree_add_12_51_groupi_n_498 ,csa_tree_add_12_51_groupi_n_497);
  not csa_tree_add_12_51_groupi_drc_bufs24838(csa_tree_add_12_51_groupi_n_497 ,csa_tree_add_12_51_groupi_n_2342);
  not csa_tree_add_12_51_groupi_drc_bufs24840(csa_tree_add_12_51_groupi_n_496 ,csa_tree_add_12_51_groupi_n_494);
  not csa_tree_add_12_51_groupi_drc_bufs24841(csa_tree_add_12_51_groupi_n_495 ,csa_tree_add_12_51_groupi_n_494);
  not csa_tree_add_12_51_groupi_drc_bufs24842(csa_tree_add_12_51_groupi_n_494 ,csa_tree_add_12_51_groupi_n_2243);
  not csa_tree_add_12_51_groupi_drc_bufs24844(csa_tree_add_12_51_groupi_n_493 ,csa_tree_add_12_51_groupi_n_491);
  not csa_tree_add_12_51_groupi_drc_bufs24845(csa_tree_add_12_51_groupi_n_492 ,csa_tree_add_12_51_groupi_n_491);
  not csa_tree_add_12_51_groupi_drc_bufs24846(csa_tree_add_12_51_groupi_n_491 ,csa_tree_add_12_51_groupi_n_2225);
  not csa_tree_add_12_51_groupi_drc_bufs24848(csa_tree_add_12_51_groupi_n_490 ,csa_tree_add_12_51_groupi_n_488);
  not csa_tree_add_12_51_groupi_drc_bufs24849(csa_tree_add_12_51_groupi_n_489 ,csa_tree_add_12_51_groupi_n_488);
  not csa_tree_add_12_51_groupi_drc_bufs24850(csa_tree_add_12_51_groupi_n_488 ,csa_tree_add_12_51_groupi_n_2244);
  not csa_tree_add_12_51_groupi_drc_bufs24852(csa_tree_add_12_51_groupi_n_487 ,csa_tree_add_12_51_groupi_n_485);
  not csa_tree_add_12_51_groupi_drc_bufs24853(csa_tree_add_12_51_groupi_n_486 ,csa_tree_add_12_51_groupi_n_485);
  not csa_tree_add_12_51_groupi_drc_bufs24854(csa_tree_add_12_51_groupi_n_485 ,csa_tree_add_12_51_groupi_n_2235);
  not csa_tree_add_12_51_groupi_drc_bufs24856(csa_tree_add_12_51_groupi_n_484 ,csa_tree_add_12_51_groupi_n_482);
  not csa_tree_add_12_51_groupi_drc_bufs24857(csa_tree_add_12_51_groupi_n_483 ,csa_tree_add_12_51_groupi_n_482);
  not csa_tree_add_12_51_groupi_drc_bufs24858(csa_tree_add_12_51_groupi_n_482 ,csa_tree_add_12_51_groupi_n_2325);
  not csa_tree_add_12_51_groupi_drc_bufs24860(csa_tree_add_12_51_groupi_n_481 ,csa_tree_add_12_51_groupi_n_479);
  not csa_tree_add_12_51_groupi_drc_bufs24861(csa_tree_add_12_51_groupi_n_480 ,csa_tree_add_12_51_groupi_n_479);
  not csa_tree_add_12_51_groupi_drc_bufs24862(csa_tree_add_12_51_groupi_n_479 ,csa_tree_add_12_51_groupi_n_2333);
  not csa_tree_add_12_51_groupi_drc_bufs24864(csa_tree_add_12_51_groupi_n_478 ,csa_tree_add_12_51_groupi_n_476);
  not csa_tree_add_12_51_groupi_drc_bufs24865(csa_tree_add_12_51_groupi_n_477 ,csa_tree_add_12_51_groupi_n_476);
  not csa_tree_add_12_51_groupi_drc_bufs24866(csa_tree_add_12_51_groupi_n_476 ,csa_tree_add_12_51_groupi_n_2296);
  not csa_tree_add_12_51_groupi_drc_bufs24868(csa_tree_add_12_51_groupi_n_475 ,csa_tree_add_12_51_groupi_n_473);
  not csa_tree_add_12_51_groupi_drc_bufs24869(csa_tree_add_12_51_groupi_n_474 ,csa_tree_add_12_51_groupi_n_473);
  not csa_tree_add_12_51_groupi_drc_bufs24870(csa_tree_add_12_51_groupi_n_473 ,csa_tree_add_12_51_groupi_n_2295);
  not csa_tree_add_12_51_groupi_drc_bufs24872(csa_tree_add_12_51_groupi_n_472 ,csa_tree_add_12_51_groupi_n_470);
  not csa_tree_add_12_51_groupi_drc_bufs24873(csa_tree_add_12_51_groupi_n_471 ,csa_tree_add_12_51_groupi_n_470);
  not csa_tree_add_12_51_groupi_drc_bufs24874(csa_tree_add_12_51_groupi_n_470 ,csa_tree_add_12_51_groupi_n_2286);
  not csa_tree_add_12_51_groupi_drc_bufs24876(csa_tree_add_12_51_groupi_n_469 ,csa_tree_add_12_51_groupi_n_467);
  not csa_tree_add_12_51_groupi_drc_bufs24877(csa_tree_add_12_51_groupi_n_468 ,csa_tree_add_12_51_groupi_n_467);
  not csa_tree_add_12_51_groupi_drc_bufs24878(csa_tree_add_12_51_groupi_n_467 ,csa_tree_add_12_51_groupi_n_2258);
  not csa_tree_add_12_51_groupi_drc_bufs24880(csa_tree_add_12_51_groupi_n_466 ,csa_tree_add_12_51_groupi_n_464);
  not csa_tree_add_12_51_groupi_drc_bufs24881(csa_tree_add_12_51_groupi_n_465 ,csa_tree_add_12_51_groupi_n_464);
  not csa_tree_add_12_51_groupi_drc_bufs24882(csa_tree_add_12_51_groupi_n_464 ,csa_tree_add_12_51_groupi_n_2249);
  not csa_tree_add_12_51_groupi_drc_bufs24884(csa_tree_add_12_51_groupi_n_463 ,csa_tree_add_12_51_groupi_n_461);
  not csa_tree_add_12_51_groupi_drc_bufs24885(csa_tree_add_12_51_groupi_n_462 ,csa_tree_add_12_51_groupi_n_461);
  not csa_tree_add_12_51_groupi_drc_bufs24886(csa_tree_add_12_51_groupi_n_461 ,csa_tree_add_12_51_groupi_n_2213);
  not csa_tree_add_12_51_groupi_drc_bufs24888(csa_tree_add_12_51_groupi_n_460 ,csa_tree_add_12_51_groupi_n_458);
  not csa_tree_add_12_51_groupi_drc_bufs24889(csa_tree_add_12_51_groupi_n_459 ,csa_tree_add_12_51_groupi_n_458);
  not csa_tree_add_12_51_groupi_drc_bufs24890(csa_tree_add_12_51_groupi_n_458 ,csa_tree_add_12_51_groupi_n_2341);
  not csa_tree_add_12_51_groupi_drc_bufs24892(csa_tree_add_12_51_groupi_n_457 ,csa_tree_add_12_51_groupi_n_455);
  not csa_tree_add_12_51_groupi_drc_bufs24893(csa_tree_add_12_51_groupi_n_456 ,csa_tree_add_12_51_groupi_n_455);
  not csa_tree_add_12_51_groupi_drc_bufs24894(csa_tree_add_12_51_groupi_n_455 ,csa_tree_add_12_51_groupi_n_2210);
  not csa_tree_add_12_51_groupi_drc_bufs24896(csa_tree_add_12_51_groupi_n_454 ,csa_tree_add_12_51_groupi_n_452);
  not csa_tree_add_12_51_groupi_drc_bufs24897(csa_tree_add_12_51_groupi_n_453 ,csa_tree_add_12_51_groupi_n_452);
  not csa_tree_add_12_51_groupi_drc_bufs24898(csa_tree_add_12_51_groupi_n_452 ,csa_tree_add_12_51_groupi_n_2242);
  not csa_tree_add_12_51_groupi_drc_bufs24900(csa_tree_add_12_51_groupi_n_451 ,csa_tree_add_12_51_groupi_n_449);
  not csa_tree_add_12_51_groupi_drc_bufs24901(csa_tree_add_12_51_groupi_n_450 ,csa_tree_add_12_51_groupi_n_449);
  not csa_tree_add_12_51_groupi_drc_bufs24902(csa_tree_add_12_51_groupi_n_449 ,csa_tree_add_12_51_groupi_n_2209);
  not csa_tree_add_12_51_groupi_drc_bufs24904(csa_tree_add_12_51_groupi_n_448 ,csa_tree_add_12_51_groupi_n_446);
  not csa_tree_add_12_51_groupi_drc_bufs24905(csa_tree_add_12_51_groupi_n_447 ,csa_tree_add_12_51_groupi_n_446);
  not csa_tree_add_12_51_groupi_drc_bufs24906(csa_tree_add_12_51_groupi_n_446 ,csa_tree_add_12_51_groupi_n_2321);
  not csa_tree_add_12_51_groupi_drc_bufs24908(csa_tree_add_12_51_groupi_n_445 ,csa_tree_add_12_51_groupi_n_443);
  not csa_tree_add_12_51_groupi_drc_bufs24909(csa_tree_add_12_51_groupi_n_444 ,csa_tree_add_12_51_groupi_n_443);
  not csa_tree_add_12_51_groupi_drc_bufs24910(csa_tree_add_12_51_groupi_n_443 ,csa_tree_add_12_51_groupi_n_2251);
  not csa_tree_add_12_51_groupi_drc_bufs24912(csa_tree_add_12_51_groupi_n_442 ,csa_tree_add_12_51_groupi_n_440);
  not csa_tree_add_12_51_groupi_drc_bufs24913(csa_tree_add_12_51_groupi_n_441 ,csa_tree_add_12_51_groupi_n_440);
  not csa_tree_add_12_51_groupi_drc_bufs24914(csa_tree_add_12_51_groupi_n_440 ,csa_tree_add_12_51_groupi_n_2285);
  not csa_tree_add_12_51_groupi_drc_bufs24916(csa_tree_add_12_51_groupi_n_439 ,csa_tree_add_12_51_groupi_n_437);
  not csa_tree_add_12_51_groupi_drc_bufs24917(csa_tree_add_12_51_groupi_n_438 ,csa_tree_add_12_51_groupi_n_437);
  not csa_tree_add_12_51_groupi_drc_bufs24918(csa_tree_add_12_51_groupi_n_437 ,csa_tree_add_12_51_groupi_n_2305);
  not csa_tree_add_12_51_groupi_drc_bufs24920(csa_tree_add_12_51_groupi_n_436 ,csa_tree_add_12_51_groupi_n_434);
  not csa_tree_add_12_51_groupi_drc_bufs24921(csa_tree_add_12_51_groupi_n_435 ,csa_tree_add_12_51_groupi_n_434);
  not csa_tree_add_12_51_groupi_drc_bufs24922(csa_tree_add_12_51_groupi_n_434 ,csa_tree_add_12_51_groupi_n_2330);
  not csa_tree_add_12_51_groupi_drc_bufs24924(csa_tree_add_12_51_groupi_n_433 ,csa_tree_add_12_51_groupi_n_431);
  not csa_tree_add_12_51_groupi_drc_bufs24925(csa_tree_add_12_51_groupi_n_432 ,csa_tree_add_12_51_groupi_n_431);
  not csa_tree_add_12_51_groupi_drc_bufs24926(csa_tree_add_12_51_groupi_n_431 ,csa_tree_add_12_51_groupi_n_2312);
  not csa_tree_add_12_51_groupi_drc_bufs24928(csa_tree_add_12_51_groupi_n_430 ,csa_tree_add_12_51_groupi_n_428);
  not csa_tree_add_12_51_groupi_drc_bufs24929(csa_tree_add_12_51_groupi_n_429 ,csa_tree_add_12_51_groupi_n_428);
  not csa_tree_add_12_51_groupi_drc_bufs24930(csa_tree_add_12_51_groupi_n_428 ,csa_tree_add_12_51_groupi_n_2304);
  not csa_tree_add_12_51_groupi_drc_bufs24932(csa_tree_add_12_51_groupi_n_427 ,csa_tree_add_12_51_groupi_n_425);
  not csa_tree_add_12_51_groupi_drc_bufs24933(csa_tree_add_12_51_groupi_n_426 ,csa_tree_add_12_51_groupi_n_425);
  not csa_tree_add_12_51_groupi_drc_bufs24934(csa_tree_add_12_51_groupi_n_425 ,csa_tree_add_12_51_groupi_n_2240);
  not csa_tree_add_12_51_groupi_drc_bufs24936(csa_tree_add_12_51_groupi_n_424 ,csa_tree_add_12_51_groupi_n_422);
  not csa_tree_add_12_51_groupi_drc_bufs24937(csa_tree_add_12_51_groupi_n_423 ,csa_tree_add_12_51_groupi_n_422);
  not csa_tree_add_12_51_groupi_drc_bufs24938(csa_tree_add_12_51_groupi_n_422 ,csa_tree_add_12_51_groupi_n_2258);
  not csa_tree_add_12_51_groupi_drc_bufs24940(csa_tree_add_12_51_groupi_n_421 ,csa_tree_add_12_51_groupi_n_419);
  not csa_tree_add_12_51_groupi_drc_bufs24941(csa_tree_add_12_51_groupi_n_420 ,csa_tree_add_12_51_groupi_n_419);
  not csa_tree_add_12_51_groupi_drc_bufs24942(csa_tree_add_12_51_groupi_n_419 ,csa_tree_add_12_51_groupi_n_2332);
  not csa_tree_add_12_51_groupi_drc_bufs24944(csa_tree_add_12_51_groupi_n_418 ,csa_tree_add_12_51_groupi_n_416);
  not csa_tree_add_12_51_groupi_drc_bufs24945(csa_tree_add_12_51_groupi_n_417 ,csa_tree_add_12_51_groupi_n_416);
  not csa_tree_add_12_51_groupi_drc_bufs24946(csa_tree_add_12_51_groupi_n_416 ,csa_tree_add_12_51_groupi_n_2287);
  not csa_tree_add_12_51_groupi_drc_bufs24948(csa_tree_add_12_51_groupi_n_415 ,csa_tree_add_12_51_groupi_n_413);
  not csa_tree_add_12_51_groupi_drc_bufs24949(csa_tree_add_12_51_groupi_n_414 ,csa_tree_add_12_51_groupi_n_413);
  not csa_tree_add_12_51_groupi_drc_bufs24950(csa_tree_add_12_51_groupi_n_413 ,csa_tree_add_12_51_groupi_n_2232);
  not csa_tree_add_12_51_groupi_drc_bufs24952(csa_tree_add_12_51_groupi_n_412 ,csa_tree_add_12_51_groupi_n_410);
  not csa_tree_add_12_51_groupi_drc_bufs24953(csa_tree_add_12_51_groupi_n_411 ,csa_tree_add_12_51_groupi_n_410);
  not csa_tree_add_12_51_groupi_drc_bufs24954(csa_tree_add_12_51_groupi_n_410 ,csa_tree_add_12_51_groupi_n_2231);
  not csa_tree_add_12_51_groupi_drc_bufs24956(csa_tree_add_12_51_groupi_n_409 ,csa_tree_add_12_51_groupi_n_407);
  not csa_tree_add_12_51_groupi_drc_bufs24957(csa_tree_add_12_51_groupi_n_408 ,csa_tree_add_12_51_groupi_n_407);
  not csa_tree_add_12_51_groupi_drc_bufs24958(csa_tree_add_12_51_groupi_n_407 ,csa_tree_add_12_51_groupi_n_2207);
  not csa_tree_add_12_51_groupi_drc_bufs24960(csa_tree_add_12_51_groupi_n_406 ,csa_tree_add_12_51_groupi_n_404);
  not csa_tree_add_12_51_groupi_drc_bufs24961(csa_tree_add_12_51_groupi_n_405 ,csa_tree_add_12_51_groupi_n_404);
  not csa_tree_add_12_51_groupi_drc_bufs24962(csa_tree_add_12_51_groupi_n_404 ,csa_tree_add_12_51_groupi_n_2322);
  not csa_tree_add_12_51_groupi_drc_bufs24964(csa_tree_add_12_51_groupi_n_403 ,csa_tree_add_12_51_groupi_n_401);
  not csa_tree_add_12_51_groupi_drc_bufs24965(csa_tree_add_12_51_groupi_n_402 ,csa_tree_add_12_51_groupi_n_401);
  not csa_tree_add_12_51_groupi_drc_bufs24966(csa_tree_add_12_51_groupi_n_401 ,csa_tree_add_12_51_groupi_n_2294);
  not csa_tree_add_12_51_groupi_drc_bufs24968(csa_tree_add_12_51_groupi_n_400 ,csa_tree_add_12_51_groupi_n_398);
  not csa_tree_add_12_51_groupi_drc_bufs24969(csa_tree_add_12_51_groupi_n_399 ,csa_tree_add_12_51_groupi_n_398);
  not csa_tree_add_12_51_groupi_drc_bufs24970(csa_tree_add_12_51_groupi_n_398 ,csa_tree_add_12_51_groupi_n_2259);
  not csa_tree_add_12_51_groupi_drc_bufs24972(csa_tree_add_12_51_groupi_n_397 ,csa_tree_add_12_51_groupi_n_395);
  not csa_tree_add_12_51_groupi_drc_bufs24973(csa_tree_add_12_51_groupi_n_396 ,csa_tree_add_12_51_groupi_n_395);
  not csa_tree_add_12_51_groupi_drc_bufs24974(csa_tree_add_12_51_groupi_n_395 ,csa_tree_add_12_51_groupi_n_2314);
  not csa_tree_add_12_51_groupi_drc_bufs24976(csa_tree_add_12_51_groupi_n_394 ,csa_tree_add_12_51_groupi_n_392);
  not csa_tree_add_12_51_groupi_drc_bufs24977(csa_tree_add_12_51_groupi_n_393 ,csa_tree_add_12_51_groupi_n_392);
  not csa_tree_add_12_51_groupi_drc_bufs24978(csa_tree_add_12_51_groupi_n_392 ,csa_tree_add_12_51_groupi_n_2223);
  not csa_tree_add_12_51_groupi_drc_bufs24980(csa_tree_add_12_51_groupi_n_391 ,csa_tree_add_12_51_groupi_n_389);
  not csa_tree_add_12_51_groupi_drc_bufs24981(csa_tree_add_12_51_groupi_n_390 ,csa_tree_add_12_51_groupi_n_389);
  not csa_tree_add_12_51_groupi_drc_bufs24982(csa_tree_add_12_51_groupi_n_389 ,csa_tree_add_12_51_groupi_n_2339);
  not csa_tree_add_12_51_groupi_drc_bufs24984(csa_tree_add_12_51_groupi_n_388 ,csa_tree_add_12_51_groupi_n_386);
  not csa_tree_add_12_51_groupi_drc_bufs24985(csa_tree_add_12_51_groupi_n_387 ,csa_tree_add_12_51_groupi_n_386);
  not csa_tree_add_12_51_groupi_drc_bufs24986(csa_tree_add_12_51_groupi_n_386 ,csa_tree_add_12_51_groupi_n_2304);
  not csa_tree_add_12_51_groupi_drc_bufs24988(csa_tree_add_12_51_groupi_n_385 ,csa_tree_add_12_51_groupi_n_383);
  not csa_tree_add_12_51_groupi_drc_bufs24989(csa_tree_add_12_51_groupi_n_384 ,csa_tree_add_12_51_groupi_n_383);
  not csa_tree_add_12_51_groupi_drc_bufs24990(csa_tree_add_12_51_groupi_n_383 ,csa_tree_add_12_51_groupi_n_2287);
  not csa_tree_add_12_51_groupi_drc_bufs24992(csa_tree_add_12_51_groupi_n_382 ,csa_tree_add_12_51_groupi_n_380);
  not csa_tree_add_12_51_groupi_drc_bufs24993(csa_tree_add_12_51_groupi_n_381 ,csa_tree_add_12_51_groupi_n_380);
  not csa_tree_add_12_51_groupi_drc_bufs24994(csa_tree_add_12_51_groupi_n_380 ,csa_tree_add_12_51_groupi_n_2314);
  not csa_tree_add_12_51_groupi_drc_bufs24996(csa_tree_add_12_51_groupi_n_379 ,csa_tree_add_12_51_groupi_n_377);
  not csa_tree_add_12_51_groupi_drc_bufs24997(csa_tree_add_12_51_groupi_n_378 ,csa_tree_add_12_51_groupi_n_377);
  not csa_tree_add_12_51_groupi_drc_bufs24998(csa_tree_add_12_51_groupi_n_377 ,csa_tree_add_12_51_groupi_n_2241);
  not csa_tree_add_12_51_groupi_drc_bufs25000(csa_tree_add_12_51_groupi_n_376 ,csa_tree_add_12_51_groupi_n_374);
  not csa_tree_add_12_51_groupi_drc_bufs25001(csa_tree_add_12_51_groupi_n_375 ,csa_tree_add_12_51_groupi_n_374);
  not csa_tree_add_12_51_groupi_drc_bufs25002(csa_tree_add_12_51_groupi_n_374 ,csa_tree_add_12_51_groupi_n_2250);
  not csa_tree_add_12_51_groupi_drc_bufs25004(csa_tree_add_12_51_groupi_n_373 ,csa_tree_add_12_51_groupi_n_371);
  not csa_tree_add_12_51_groupi_drc_bufs25005(csa_tree_add_12_51_groupi_n_372 ,csa_tree_add_12_51_groupi_n_371);
  not csa_tree_add_12_51_groupi_drc_bufs25006(csa_tree_add_12_51_groupi_n_371 ,csa_tree_add_12_51_groupi_n_2217);
  not csa_tree_add_12_51_groupi_drc_bufs25008(csa_tree_add_12_51_groupi_n_370 ,csa_tree_add_12_51_groupi_n_368);
  not csa_tree_add_12_51_groupi_drc_bufs25009(csa_tree_add_12_51_groupi_n_369 ,csa_tree_add_12_51_groupi_n_368);
  not csa_tree_add_12_51_groupi_drc_bufs25010(csa_tree_add_12_51_groupi_n_368 ,csa_tree_add_12_51_groupi_n_2322);
  not csa_tree_add_12_51_groupi_drc_bufs25012(csa_tree_add_12_51_groupi_n_367 ,csa_tree_add_12_51_groupi_n_365);
  not csa_tree_add_12_51_groupi_drc_bufs25013(csa_tree_add_12_51_groupi_n_366 ,csa_tree_add_12_51_groupi_n_365);
  not csa_tree_add_12_51_groupi_drc_bufs25014(csa_tree_add_12_51_groupi_n_365 ,csa_tree_add_12_51_groupi_n_2303);
  not csa_tree_add_12_51_groupi_drc_bufs25016(csa_tree_add_12_51_groupi_n_364 ,csa_tree_add_12_51_groupi_n_362);
  not csa_tree_add_12_51_groupi_drc_bufs25017(csa_tree_add_12_51_groupi_n_363 ,csa_tree_add_12_51_groupi_n_362);
  not csa_tree_add_12_51_groupi_drc_bufs25018(csa_tree_add_12_51_groupi_n_362 ,csa_tree_add_12_51_groupi_n_2278);
  not csa_tree_add_12_51_groupi_drc_bufs25020(csa_tree_add_12_51_groupi_n_361 ,csa_tree_add_12_51_groupi_n_359);
  not csa_tree_add_12_51_groupi_drc_bufs25021(csa_tree_add_12_51_groupi_n_360 ,csa_tree_add_12_51_groupi_n_359);
  not csa_tree_add_12_51_groupi_drc_bufs25022(csa_tree_add_12_51_groupi_n_359 ,csa_tree_add_12_51_groupi_n_2233);
  not csa_tree_add_12_51_groupi_drc_bufs25024(csa_tree_add_12_51_groupi_n_358 ,csa_tree_add_12_51_groupi_n_356);
  not csa_tree_add_12_51_groupi_drc_bufs25025(csa_tree_add_12_51_groupi_n_357 ,csa_tree_add_12_51_groupi_n_356);
  not csa_tree_add_12_51_groupi_drc_bufs25026(csa_tree_add_12_51_groupi_n_356 ,csa_tree_add_12_51_groupi_n_2232);
  not csa_tree_add_12_51_groupi_drc_bufs25028(csa_tree_add_12_51_groupi_n_355 ,csa_tree_add_12_51_groupi_n_353);
  not csa_tree_add_12_51_groupi_drc_bufs25029(csa_tree_add_12_51_groupi_n_354 ,csa_tree_add_12_51_groupi_n_353);
  not csa_tree_add_12_51_groupi_drc_bufs25030(csa_tree_add_12_51_groupi_n_353 ,csa_tree_add_12_51_groupi_n_2303);
  not csa_tree_add_12_51_groupi_drc_bufs25032(csa_tree_add_12_51_groupi_n_352 ,csa_tree_add_12_51_groupi_n_350);
  not csa_tree_add_12_51_groupi_drc_bufs25033(csa_tree_add_12_51_groupi_n_351 ,csa_tree_add_12_51_groupi_n_350);
  not csa_tree_add_12_51_groupi_drc_bufs25034(csa_tree_add_12_51_groupi_n_350 ,csa_tree_add_12_51_groupi_n_2241);
  not csa_tree_add_12_51_groupi_drc_bufs25036(csa_tree_add_12_51_groupi_n_349 ,csa_tree_add_12_51_groupi_n_347);
  not csa_tree_add_12_51_groupi_drc_bufs25037(csa_tree_add_12_51_groupi_n_348 ,csa_tree_add_12_51_groupi_n_347);
  not csa_tree_add_12_51_groupi_drc_bufs25038(csa_tree_add_12_51_groupi_n_347 ,csa_tree_add_12_51_groupi_n_2269);
  not csa_tree_add_12_51_groupi_drc_bufs25040(csa_tree_add_12_51_groupi_n_346 ,csa_tree_add_12_51_groupi_n_344);
  not csa_tree_add_12_51_groupi_drc_bufs25041(csa_tree_add_12_51_groupi_n_345 ,csa_tree_add_12_51_groupi_n_344);
  not csa_tree_add_12_51_groupi_drc_bufs25042(csa_tree_add_12_51_groupi_n_344 ,csa_tree_add_12_51_groupi_n_2295);
  not csa_tree_add_12_51_groupi_drc_bufs25044(csa_tree_add_12_51_groupi_n_343 ,csa_tree_add_12_51_groupi_n_341);
  not csa_tree_add_12_51_groupi_drc_bufs25045(csa_tree_add_12_51_groupi_n_342 ,csa_tree_add_12_51_groupi_n_341);
  not csa_tree_add_12_51_groupi_drc_bufs25046(csa_tree_add_12_51_groupi_n_341 ,csa_tree_add_12_51_groupi_n_2251);
  not csa_tree_add_12_51_groupi_drc_bufs25048(csa_tree_add_12_51_groupi_n_340 ,csa_tree_add_12_51_groupi_n_338);
  not csa_tree_add_12_51_groupi_drc_bufs25049(csa_tree_add_12_51_groupi_n_339 ,csa_tree_add_12_51_groupi_n_338);
  not csa_tree_add_12_51_groupi_drc_bufs25050(csa_tree_add_12_51_groupi_n_338 ,csa_tree_add_12_51_groupi_n_2233);
  not csa_tree_add_12_51_groupi_drc_bufs25052(csa_tree_add_12_51_groupi_n_337 ,csa_tree_add_12_51_groupi_n_335);
  not csa_tree_add_12_51_groupi_drc_bufs25053(csa_tree_add_12_51_groupi_n_336 ,csa_tree_add_12_51_groupi_n_335);
  not csa_tree_add_12_51_groupi_drc_bufs25054(csa_tree_add_12_51_groupi_n_335 ,csa_tree_add_12_51_groupi_n_2216);
  not csa_tree_add_12_51_groupi_drc_bufs25056(csa_tree_add_12_51_groupi_n_334 ,csa_tree_add_12_51_groupi_n_332);
  not csa_tree_add_12_51_groupi_drc_bufs25057(csa_tree_add_12_51_groupi_n_333 ,csa_tree_add_12_51_groupi_n_332);
  not csa_tree_add_12_51_groupi_drc_bufs25058(csa_tree_add_12_51_groupi_n_332 ,csa_tree_add_12_51_groupi_n_2267);
  not csa_tree_add_12_51_groupi_drc_bufs25060(csa_tree_add_12_51_groupi_n_331 ,csa_tree_add_12_51_groupi_n_329);
  not csa_tree_add_12_51_groupi_drc_bufs25061(csa_tree_add_12_51_groupi_n_330 ,csa_tree_add_12_51_groupi_n_329);
  not csa_tree_add_12_51_groupi_drc_bufs25062(csa_tree_add_12_51_groupi_n_329 ,csa_tree_add_12_51_groupi_n_2276);
  not csa_tree_add_12_51_groupi_drc_bufs25064(csa_tree_add_12_51_groupi_n_328 ,csa_tree_add_12_51_groupi_n_326);
  not csa_tree_add_12_51_groupi_drc_bufs25065(csa_tree_add_12_51_groupi_n_327 ,csa_tree_add_12_51_groupi_n_326);
  not csa_tree_add_12_51_groupi_drc_bufs25066(csa_tree_add_12_51_groupi_n_326 ,csa_tree_add_12_51_groupi_n_2313);
  not csa_tree_add_12_51_groupi_drc_bufs25068(csa_tree_add_12_51_groupi_n_325 ,csa_tree_add_12_51_groupi_n_323);
  not csa_tree_add_12_51_groupi_drc_bufs25069(csa_tree_add_12_51_groupi_n_324 ,csa_tree_add_12_51_groupi_n_323);
  not csa_tree_add_12_51_groupi_drc_bufs25070(csa_tree_add_12_51_groupi_n_323 ,csa_tree_add_12_51_groupi_n_2296);
  not csa_tree_add_12_51_groupi_drc_bufs25072(csa_tree_add_12_51_groupi_n_322 ,csa_tree_add_12_51_groupi_n_320);
  not csa_tree_add_12_51_groupi_drc_bufs25073(csa_tree_add_12_51_groupi_n_321 ,csa_tree_add_12_51_groupi_n_320);
  not csa_tree_add_12_51_groupi_drc_bufs25074(csa_tree_add_12_51_groupi_n_320 ,csa_tree_add_12_51_groupi_n_2214);
  not csa_tree_add_12_51_groupi_drc_bufs25076(csa_tree_add_12_51_groupi_n_319 ,csa_tree_add_12_51_groupi_n_317);
  not csa_tree_add_12_51_groupi_drc_bufs25077(csa_tree_add_12_51_groupi_n_318 ,csa_tree_add_12_51_groupi_n_317);
  not csa_tree_add_12_51_groupi_drc_bufs25078(csa_tree_add_12_51_groupi_n_317 ,csa_tree_add_12_51_groupi_n_2269);
  not csa_tree_add_12_51_groupi_drc_bufs25080(csa_tree_add_12_51_groupi_n_316 ,csa_tree_add_12_51_groupi_n_314);
  not csa_tree_add_12_51_groupi_drc_bufs25081(csa_tree_add_12_51_groupi_n_315 ,csa_tree_add_12_51_groupi_n_314);
  not csa_tree_add_12_51_groupi_drc_bufs25082(csa_tree_add_12_51_groupi_n_314 ,csa_tree_add_12_51_groupi_n_2323);
  not csa_tree_add_12_51_groupi_drc_bufs25084(csa_tree_add_12_51_groupi_n_313 ,csa_tree_add_12_51_groupi_n_311);
  not csa_tree_add_12_51_groupi_drc_bufs25085(csa_tree_add_12_51_groupi_n_312 ,csa_tree_add_12_51_groupi_n_311);
  not csa_tree_add_12_51_groupi_drc_bufs25086(csa_tree_add_12_51_groupi_n_311 ,csa_tree_add_12_51_groupi_n_2277);
  not csa_tree_add_12_51_groupi_drc_bufs25088(csa_tree_add_12_51_groupi_n_310 ,csa_tree_add_12_51_groupi_n_308);
  not csa_tree_add_12_51_groupi_drc_bufs25089(csa_tree_add_12_51_groupi_n_309 ,csa_tree_add_12_51_groupi_n_308);
  not csa_tree_add_12_51_groupi_drc_bufs25090(csa_tree_add_12_51_groupi_n_308 ,csa_tree_add_12_51_groupi_n_2214);
  not csa_tree_add_12_51_groupi_drc_bufs25092(csa_tree_add_12_51_groupi_n_307 ,csa_tree_add_12_51_groupi_n_305);
  not csa_tree_add_12_51_groupi_drc_bufs25093(csa_tree_add_12_51_groupi_n_306 ,csa_tree_add_12_51_groupi_n_305);
  not csa_tree_add_12_51_groupi_drc_bufs25094(csa_tree_add_12_51_groupi_n_305 ,csa_tree_add_12_51_groupi_n_2213);
  not csa_tree_add_12_51_groupi_drc_bufs25096(csa_tree_add_12_51_groupi_n_304 ,csa_tree_add_12_51_groupi_n_302);
  not csa_tree_add_12_51_groupi_drc_bufs25097(csa_tree_add_12_51_groupi_n_303 ,csa_tree_add_12_51_groupi_n_302);
  not csa_tree_add_12_51_groupi_drc_bufs25098(csa_tree_add_12_51_groupi_n_302 ,csa_tree_add_12_51_groupi_n_2215);
  not csa_tree_add_12_51_groupi_drc_bufs25100(csa_tree_add_12_51_groupi_n_301 ,csa_tree_add_12_51_groupi_n_299);
  not csa_tree_add_12_51_groupi_drc_bufs25101(csa_tree_add_12_51_groupi_n_300 ,csa_tree_add_12_51_groupi_n_299);
  not csa_tree_add_12_51_groupi_drc_bufs25102(csa_tree_add_12_51_groupi_n_299 ,csa_tree_add_12_51_groupi_n_2222);
  not csa_tree_add_12_51_groupi_drc_bufs25104(csa_tree_add_12_51_groupi_n_298 ,csa_tree_add_12_51_groupi_n_296);
  not csa_tree_add_12_51_groupi_drc_bufs25105(csa_tree_add_12_51_groupi_n_297 ,csa_tree_add_12_51_groupi_n_296);
  not csa_tree_add_12_51_groupi_drc_bufs25106(csa_tree_add_12_51_groupi_n_296 ,csa_tree_add_12_51_groupi_n_2223);
  not csa_tree_add_12_51_groupi_drc_bufs25108(csa_tree_add_12_51_groupi_n_295 ,csa_tree_add_12_51_groupi_n_293);
  not csa_tree_add_12_51_groupi_drc_bufs25109(csa_tree_add_12_51_groupi_n_294 ,csa_tree_add_12_51_groupi_n_293);
  not csa_tree_add_12_51_groupi_drc_bufs25110(csa_tree_add_12_51_groupi_n_293 ,csa_tree_add_12_51_groupi_n_2211);
  not csa_tree_add_12_51_groupi_drc_bufs25112(csa_tree_add_12_51_groupi_n_292 ,csa_tree_add_12_51_groupi_n_290);
  not csa_tree_add_12_51_groupi_drc_bufs25113(csa_tree_add_12_51_groupi_n_291 ,csa_tree_add_12_51_groupi_n_290);
  not csa_tree_add_12_51_groupi_drc_bufs25114(csa_tree_add_12_51_groupi_n_290 ,csa_tree_add_12_51_groupi_n_2276);
  not csa_tree_add_12_51_groupi_drc_bufs25116(csa_tree_add_12_51_groupi_n_289 ,csa_tree_add_12_51_groupi_n_287);
  not csa_tree_add_12_51_groupi_drc_bufs25117(csa_tree_add_12_51_groupi_n_288 ,csa_tree_add_12_51_groupi_n_287);
  not csa_tree_add_12_51_groupi_drc_bufs25118(csa_tree_add_12_51_groupi_n_287 ,csa_tree_add_12_51_groupi_n_2216);
  not csa_tree_add_12_51_groupi_drc_bufs25120(csa_tree_add_12_51_groupi_n_286 ,csa_tree_add_12_51_groupi_n_284);
  not csa_tree_add_12_51_groupi_drc_bufs25121(csa_tree_add_12_51_groupi_n_285 ,csa_tree_add_12_51_groupi_n_284);
  not csa_tree_add_12_51_groupi_drc_bufs25122(csa_tree_add_12_51_groupi_n_284 ,csa_tree_add_12_51_groupi_n_2268);
  not csa_tree_add_12_51_groupi_drc_bufs25124(csa_tree_add_12_51_groupi_n_283 ,csa_tree_add_12_51_groupi_n_281);
  not csa_tree_add_12_51_groupi_drc_bufs25125(csa_tree_add_12_51_groupi_n_282 ,csa_tree_add_12_51_groupi_n_281);
  not csa_tree_add_12_51_groupi_drc_bufs25126(csa_tree_add_12_51_groupi_n_281 ,csa_tree_add_12_51_groupi_n_2268);
  not csa_tree_add_12_51_groupi_drc_bufs25128(csa_tree_add_12_51_groupi_n_280 ,csa_tree_add_12_51_groupi_n_278);
  not csa_tree_add_12_51_groupi_drc_bufs25129(csa_tree_add_12_51_groupi_n_279 ,csa_tree_add_12_51_groupi_n_278);
  not csa_tree_add_12_51_groupi_drc_bufs25130(csa_tree_add_12_51_groupi_n_278 ,csa_tree_add_12_51_groupi_n_2260);
  not csa_tree_add_12_51_groupi_drc_bufs25132(csa_tree_add_12_51_groupi_n_277 ,csa_tree_add_12_51_groupi_n_275);
  not csa_tree_add_12_51_groupi_drc_bufs25133(csa_tree_add_12_51_groupi_n_276 ,csa_tree_add_12_51_groupi_n_275);
  not csa_tree_add_12_51_groupi_drc_bufs25134(csa_tree_add_12_51_groupi_n_275 ,csa_tree_add_12_51_groupi_n_2242);
  not csa_tree_add_12_51_groupi_drc_bufs25136(csa_tree_add_12_51_groupi_n_274 ,csa_tree_add_12_51_groupi_n_272);
  not csa_tree_add_12_51_groupi_drc_bufs25137(csa_tree_add_12_51_groupi_n_273 ,csa_tree_add_12_51_groupi_n_272);
  not csa_tree_add_12_51_groupi_drc_bufs25138(csa_tree_add_12_51_groupi_n_272 ,csa_tree_add_12_51_groupi_n_2259);
  not csa_tree_add_12_51_groupi_drc_bufs25140(csa_tree_add_12_51_groupi_n_271 ,csa_tree_add_12_51_groupi_n_269);
  not csa_tree_add_12_51_groupi_drc_bufs25141(csa_tree_add_12_51_groupi_n_270 ,csa_tree_add_12_51_groupi_n_269);
  not csa_tree_add_12_51_groupi_drc_bufs25142(csa_tree_add_12_51_groupi_n_269 ,csa_tree_add_12_51_groupi_n_2240);
  not csa_tree_add_12_51_groupi_drc_bufs25144(csa_tree_add_12_51_groupi_n_268 ,csa_tree_add_12_51_groupi_n_266);
  not csa_tree_add_12_51_groupi_drc_bufs25145(csa_tree_add_12_51_groupi_n_267 ,csa_tree_add_12_51_groupi_n_266);
  not csa_tree_add_12_51_groupi_drc_bufs25146(csa_tree_add_12_51_groupi_n_266 ,csa_tree_add_12_51_groupi_n_2267);
  not csa_tree_add_12_51_groupi_drc_bufs25148(csa_tree_add_12_51_groupi_n_265 ,csa_tree_add_12_51_groupi_n_263);
  not csa_tree_add_12_51_groupi_drc_bufs25149(csa_tree_add_12_51_groupi_n_264 ,csa_tree_add_12_51_groupi_n_263);
  not csa_tree_add_12_51_groupi_drc_bufs25150(csa_tree_add_12_51_groupi_n_263 ,csa_tree_add_12_51_groupi_n_2340);
  not csa_tree_add_12_51_groupi_drc_bufs25152(csa_tree_add_12_51_groupi_n_262 ,csa_tree_add_12_51_groupi_n_260);
  not csa_tree_add_12_51_groupi_drc_bufs25153(csa_tree_add_12_51_groupi_n_261 ,csa_tree_add_12_51_groupi_n_260);
  not csa_tree_add_12_51_groupi_drc_bufs25154(csa_tree_add_12_51_groupi_n_260 ,csa_tree_add_12_51_groupi_n_2249);
  not csa_tree_add_12_51_groupi_drc_bufs25156(csa_tree_add_12_51_groupi_n_259 ,csa_tree_add_12_51_groupi_n_257);
  not csa_tree_add_12_51_groupi_drc_bufs25157(csa_tree_add_12_51_groupi_n_258 ,csa_tree_add_12_51_groupi_n_257);
  not csa_tree_add_12_51_groupi_drc_bufs25158(csa_tree_add_12_51_groupi_n_257 ,csa_tree_add_12_51_groupi_n_2331);
  not csa_tree_add_12_51_groupi_drc_bufs25160(csa_tree_add_12_51_groupi_n_256 ,csa_tree_add_12_51_groupi_n_254);
  not csa_tree_add_12_51_groupi_drc_bufs25161(csa_tree_add_12_51_groupi_n_255 ,csa_tree_add_12_51_groupi_n_254);
  not csa_tree_add_12_51_groupi_drc_bufs25162(csa_tree_add_12_51_groupi_n_254 ,csa_tree_add_12_51_groupi_n_2332);
  not csa_tree_add_12_51_groupi_drc_bufs25164(csa_tree_add_12_51_groupi_n_253 ,csa_tree_add_12_51_groupi_n_251);
  not csa_tree_add_12_51_groupi_drc_bufs25165(csa_tree_add_12_51_groupi_n_252 ,csa_tree_add_12_51_groupi_n_251);
  not csa_tree_add_12_51_groupi_drc_bufs25166(csa_tree_add_12_51_groupi_n_251 ,csa_tree_add_12_51_groupi_n_2305);
  not csa_tree_add_12_51_groupi_drc_bufs25168(csa_tree_add_12_51_groupi_n_250 ,csa_tree_add_12_51_groupi_n_248);
  not csa_tree_add_12_51_groupi_drc_bufs25169(csa_tree_add_12_51_groupi_n_249 ,csa_tree_add_12_51_groupi_n_248);
  not csa_tree_add_12_51_groupi_drc_bufs25170(csa_tree_add_12_51_groupi_n_248 ,csa_tree_add_12_51_groupi_n_2339);
  not csa_tree_add_12_51_groupi_drc_bufs25172(csa_tree_add_12_51_groupi_n_247 ,csa_tree_add_12_51_groupi_n_245);
  not csa_tree_add_12_51_groupi_drc_bufs25173(csa_tree_add_12_51_groupi_n_246 ,csa_tree_add_12_51_groupi_n_245);
  not csa_tree_add_12_51_groupi_drc_bufs25174(csa_tree_add_12_51_groupi_n_245 ,csa_tree_add_12_51_groupi_n_2222);
  not csa_tree_add_12_51_groupi_drc_bufs25176(csa_tree_add_12_51_groupi_n_244 ,csa_tree_add_12_51_groupi_n_242);
  not csa_tree_add_12_51_groupi_drc_bufs25177(csa_tree_add_12_51_groupi_n_243 ,csa_tree_add_12_51_groupi_n_242);
  not csa_tree_add_12_51_groupi_drc_bufs25178(csa_tree_add_12_51_groupi_n_242 ,csa_tree_add_12_51_groupi_n_2286);
  not csa_tree_add_12_51_groupi_drc_bufs25180(csa_tree_add_12_51_groupi_n_241 ,csa_tree_add_12_51_groupi_n_239);
  not csa_tree_add_12_51_groupi_drc_bufs25181(csa_tree_add_12_51_groupi_n_240 ,csa_tree_add_12_51_groupi_n_239);
  not csa_tree_add_12_51_groupi_drc_bufs25182(csa_tree_add_12_51_groupi_n_239 ,csa_tree_add_12_51_groupi_n_2278);
  not csa_tree_add_12_51_groupi_drc_bufs25184(csa_tree_add_12_51_groupi_n_238 ,csa_tree_add_12_51_groupi_n_236);
  not csa_tree_add_12_51_groupi_drc_bufs25185(csa_tree_add_12_51_groupi_n_237 ,csa_tree_add_12_51_groupi_n_236);
  not csa_tree_add_12_51_groupi_drc_bufs25186(csa_tree_add_12_51_groupi_n_236 ,csa_tree_add_12_51_groupi_n_2313);
  not csa_tree_add_12_51_groupi_drc_bufs25188(csa_tree_add_12_51_groupi_n_235 ,csa_tree_add_12_51_groupi_n_233);
  not csa_tree_add_12_51_groupi_drc_bufs25189(csa_tree_add_12_51_groupi_n_234 ,csa_tree_add_12_51_groupi_n_233);
  not csa_tree_add_12_51_groupi_drc_bufs25190(csa_tree_add_12_51_groupi_n_233 ,csa_tree_add_12_51_groupi_n_2312);
  not csa_tree_add_12_51_groupi_drc_bufs25192(csa_tree_add_12_51_groupi_n_232 ,csa_tree_add_12_51_groupi_n_230);
  not csa_tree_add_12_51_groupi_drc_bufs25193(csa_tree_add_12_51_groupi_n_231 ,csa_tree_add_12_51_groupi_n_230);
  not csa_tree_add_12_51_groupi_drc_bufs25194(csa_tree_add_12_51_groupi_n_230 ,csa_tree_add_12_51_groupi_n_2330);
  not csa_tree_add_12_51_groupi_drc_bufs25196(csa_tree_add_12_51_groupi_n_229 ,csa_tree_add_12_51_groupi_n_227);
  not csa_tree_add_12_51_groupi_drc_bufs25197(csa_tree_add_12_51_groupi_n_228 ,csa_tree_add_12_51_groupi_n_227);
  not csa_tree_add_12_51_groupi_drc_bufs25198(csa_tree_add_12_51_groupi_n_227 ,csa_tree_add_12_51_groupi_n_2208);
  not csa_tree_add_12_51_groupi_drc_bufs25200(csa_tree_add_12_51_groupi_n_226 ,csa_tree_add_12_51_groupi_n_224);
  not csa_tree_add_12_51_groupi_drc_bufs25201(csa_tree_add_12_51_groupi_n_225 ,csa_tree_add_12_51_groupi_n_224);
  not csa_tree_add_12_51_groupi_drc_bufs25202(csa_tree_add_12_51_groupi_n_224 ,csa_tree_add_12_51_groupi_n_2260);
  not csa_tree_add_12_51_groupi_drc_bufs25204(csa_tree_add_12_51_groupi_n_223 ,csa_tree_add_12_51_groupi_n_221);
  not csa_tree_add_12_51_groupi_drc_bufs25205(csa_tree_add_12_51_groupi_n_222 ,csa_tree_add_12_51_groupi_n_221);
  not csa_tree_add_12_51_groupi_drc_bufs25206(csa_tree_add_12_51_groupi_n_221 ,csa_tree_add_12_51_groupi_n_2250);
  not csa_tree_add_12_51_groupi_drc_bufs25208(csa_tree_add_12_51_groupi_n_220 ,csa_tree_add_12_51_groupi_n_218);
  not csa_tree_add_12_51_groupi_drc_bufs25209(csa_tree_add_12_51_groupi_n_219 ,csa_tree_add_12_51_groupi_n_218);
  not csa_tree_add_12_51_groupi_drc_bufs25210(csa_tree_add_12_51_groupi_n_218 ,csa_tree_add_12_51_groupi_n_2215);
  not csa_tree_add_12_51_groupi_drc_bufs25212(csa_tree_add_12_51_groupi_n_217 ,csa_tree_add_12_51_groupi_n_215);
  not csa_tree_add_12_51_groupi_drc_bufs25213(csa_tree_add_12_51_groupi_n_216 ,csa_tree_add_12_51_groupi_n_215);
  not csa_tree_add_12_51_groupi_drc_bufs25214(csa_tree_add_12_51_groupi_n_215 ,csa_tree_add_12_51_groupi_n_2217);
  not csa_tree_add_12_51_groupi_drc_bufs25216(csa_tree_add_12_51_groupi_n_214 ,csa_tree_add_12_51_groupi_n_212);
  not csa_tree_add_12_51_groupi_drc_bufs25217(csa_tree_add_12_51_groupi_n_213 ,csa_tree_add_12_51_groupi_n_212);
  not csa_tree_add_12_51_groupi_drc_bufs25218(csa_tree_add_12_51_groupi_n_212 ,csa_tree_add_12_51_groupi_n_2231);
  not csa_tree_add_12_51_groupi_drc_bufs25220(csa_tree_add_12_51_groupi_n_211 ,csa_tree_add_12_51_groupi_n_209);
  not csa_tree_add_12_51_groupi_drc_bufs25221(csa_tree_add_12_51_groupi_n_210 ,csa_tree_add_12_51_groupi_n_209);
  not csa_tree_add_12_51_groupi_drc_bufs25222(csa_tree_add_12_51_groupi_n_209 ,csa_tree_add_12_51_groupi_n_2224);
  not csa_tree_add_12_51_groupi_drc_bufs25224(csa_tree_add_12_51_groupi_n_208 ,csa_tree_add_12_51_groupi_n_206);
  not csa_tree_add_12_51_groupi_drc_bufs25225(csa_tree_add_12_51_groupi_n_207 ,csa_tree_add_12_51_groupi_n_206);
  not csa_tree_add_12_51_groupi_drc_bufs25226(csa_tree_add_12_51_groupi_n_206 ,csa_tree_add_12_51_groupi_n_2331);
  not csa_tree_add_12_51_groupi_drc_bufs25228(csa_tree_add_12_51_groupi_n_205 ,csa_tree_add_12_51_groupi_n_203);
  not csa_tree_add_12_51_groupi_drc_bufs25229(csa_tree_add_12_51_groupi_n_204 ,csa_tree_add_12_51_groupi_n_203);
  not csa_tree_add_12_51_groupi_drc_bufs25230(csa_tree_add_12_51_groupi_n_203 ,csa_tree_add_12_51_groupi_n_2323);
  not csa_tree_add_12_51_groupi_drc_bufs25232(csa_tree_add_12_51_groupi_n_202 ,csa_tree_add_12_51_groupi_n_200);
  not csa_tree_add_12_51_groupi_drc_bufs25233(csa_tree_add_12_51_groupi_n_201 ,csa_tree_add_12_51_groupi_n_200);
  not csa_tree_add_12_51_groupi_drc_bufs25234(csa_tree_add_12_51_groupi_n_200 ,csa_tree_add_12_51_groupi_n_2340);
  not csa_tree_add_12_51_groupi_drc_bufs25236(csa_tree_add_12_51_groupi_n_199 ,csa_tree_add_12_51_groupi_n_197);
  not csa_tree_add_12_51_groupi_drc_bufs25237(csa_tree_add_12_51_groupi_n_198 ,csa_tree_add_12_51_groupi_n_197);
  not csa_tree_add_12_51_groupi_drc_bufs25238(csa_tree_add_12_51_groupi_n_197 ,csa_tree_add_12_51_groupi_n_2321);
  not csa_tree_add_12_51_groupi_drc_bufs25240(csa_tree_add_12_51_groupi_n_196 ,csa_tree_add_12_51_groupi_n_194);
  not csa_tree_add_12_51_groupi_drc_bufs25241(csa_tree_add_12_51_groupi_n_195 ,csa_tree_add_12_51_groupi_n_194);
  not csa_tree_add_12_51_groupi_drc_bufs25242(csa_tree_add_12_51_groupi_n_194 ,csa_tree_add_12_51_groupi_n_2294);
  not csa_tree_add_12_51_groupi_drc_bufs25244(csa_tree_add_12_51_groupi_n_193 ,csa_tree_add_12_51_groupi_n_191);
  not csa_tree_add_12_51_groupi_drc_bufs25245(csa_tree_add_12_51_groupi_n_192 ,csa_tree_add_12_51_groupi_n_191);
  not csa_tree_add_12_51_groupi_drc_bufs25246(csa_tree_add_12_51_groupi_n_191 ,csa_tree_add_12_51_groupi_n_2341);
  not csa_tree_add_12_51_groupi_drc_bufs25248(csa_tree_add_12_51_groupi_n_190 ,csa_tree_add_12_51_groupi_n_188);
  not csa_tree_add_12_51_groupi_drc_bufs25249(csa_tree_add_12_51_groupi_n_189 ,csa_tree_add_12_51_groupi_n_188);
  not csa_tree_add_12_51_groupi_drc_bufs25250(csa_tree_add_12_51_groupi_n_188 ,csa_tree_add_12_51_groupi_n_2224);
  not csa_tree_add_12_51_groupi_drc_bufs25252(csa_tree_add_12_51_groupi_n_187 ,csa_tree_add_12_51_groupi_n_185);
  not csa_tree_add_12_51_groupi_drc_bufs25253(csa_tree_add_12_51_groupi_n_186 ,csa_tree_add_12_51_groupi_n_185);
  not csa_tree_add_12_51_groupi_drc_bufs25254(csa_tree_add_12_51_groupi_n_185 ,csa_tree_add_12_51_groupi_n_2285);
  not csa_tree_add_12_51_groupi_drc_bufs25256(csa_tree_add_12_51_groupi_n_184 ,csa_tree_add_12_51_groupi_n_182);
  not csa_tree_add_12_51_groupi_drc_bufs25257(csa_tree_add_12_51_groupi_n_183 ,csa_tree_add_12_51_groupi_n_182);
  not csa_tree_add_12_51_groupi_drc_bufs25258(csa_tree_add_12_51_groupi_n_182 ,csa_tree_add_12_51_groupi_n_2277);
  not csa_tree_add_12_51_groupi_drc_bufs25260(csa_tree_add_12_51_groupi_n_181 ,csa_tree_add_12_51_groupi_n_180);
  not csa_tree_add_12_51_groupi_drc_bufs25262(csa_tree_add_12_51_groupi_n_180 ,csa_tree_add_12_51_groupi_n_2004);
  not csa_tree_add_12_51_groupi_drc_bufs25264(csa_tree_add_12_51_groupi_n_179 ,csa_tree_add_12_51_groupi_n_178);
  not csa_tree_add_12_51_groupi_drc_bufs25266(csa_tree_add_12_51_groupi_n_178 ,csa_tree_add_12_51_groupi_n_1962);
  not csa_tree_add_12_51_groupi_drc_bufs25268(csa_tree_add_12_51_groupi_n_177 ,csa_tree_add_12_51_groupi_n_176);
  not csa_tree_add_12_51_groupi_drc_bufs25270(csa_tree_add_12_51_groupi_n_176 ,csa_tree_add_12_51_groupi_n_1998);
  not csa_tree_add_12_51_groupi_drc_bufs25272(csa_tree_add_12_51_groupi_n_175 ,csa_tree_add_12_51_groupi_n_174);
  not csa_tree_add_12_51_groupi_drc_bufs25274(csa_tree_add_12_51_groupi_n_174 ,csa_tree_add_12_51_groupi_n_1980);
  not csa_tree_add_12_51_groupi_drc_bufs25276(csa_tree_add_12_51_groupi_n_173 ,csa_tree_add_12_51_groupi_n_172);
  not csa_tree_add_12_51_groupi_drc_bufs25278(csa_tree_add_12_51_groupi_n_172 ,csa_tree_add_12_51_groupi_n_1992);
  not csa_tree_add_12_51_groupi_drc_bufs25280(csa_tree_add_12_51_groupi_n_171 ,csa_tree_add_12_51_groupi_n_170);
  not csa_tree_add_12_51_groupi_drc_bufs25282(csa_tree_add_12_51_groupi_n_170 ,csa_tree_add_12_51_groupi_n_1989);
  not csa_tree_add_12_51_groupi_drc_bufs25284(csa_tree_add_12_51_groupi_n_169 ,csa_tree_add_12_51_groupi_n_168);
  not csa_tree_add_12_51_groupi_drc_bufs25286(csa_tree_add_12_51_groupi_n_168 ,csa_tree_add_12_51_groupi_n_2007);
  not csa_tree_add_12_51_groupi_drc_bufs25288(csa_tree_add_12_51_groupi_n_167 ,csa_tree_add_12_51_groupi_n_166);
  not csa_tree_add_12_51_groupi_drc_bufs25290(csa_tree_add_12_51_groupi_n_166 ,csa_tree_add_12_51_groupi_n_1995);
  not csa_tree_add_12_51_groupi_drc_bufs25292(csa_tree_add_12_51_groupi_n_165 ,csa_tree_add_12_51_groupi_n_164);
  not csa_tree_add_12_51_groupi_drc_bufs25294(csa_tree_add_12_51_groupi_n_164 ,csa_tree_add_12_51_groupi_n_1965);
  not csa_tree_add_12_51_groupi_drc_bufs25296(csa_tree_add_12_51_groupi_n_163 ,csa_tree_add_12_51_groupi_n_162);
  not csa_tree_add_12_51_groupi_drc_bufs25298(csa_tree_add_12_51_groupi_n_162 ,csa_tree_add_12_51_groupi_n_2001);
  not csa_tree_add_12_51_groupi_drc_bufs25300(csa_tree_add_12_51_groupi_n_161 ,csa_tree_add_12_51_groupi_n_160);
  not csa_tree_add_12_51_groupi_drc_bufs25302(csa_tree_add_12_51_groupi_n_160 ,csa_tree_add_12_51_groupi_n_1974);
  not csa_tree_add_12_51_groupi_drc_bufs25304(csa_tree_add_12_51_groupi_n_159 ,csa_tree_add_12_51_groupi_n_158);
  not csa_tree_add_12_51_groupi_drc_bufs25306(csa_tree_add_12_51_groupi_n_158 ,csa_tree_add_12_51_groupi_n_1986);
  not csa_tree_add_12_51_groupi_drc_bufs25308(csa_tree_add_12_51_groupi_n_157 ,csa_tree_add_12_51_groupi_n_156);
  not csa_tree_add_12_51_groupi_drc_bufs25310(csa_tree_add_12_51_groupi_n_156 ,csa_tree_add_12_51_groupi_n_1977);
  not csa_tree_add_12_51_groupi_drc_bufs25312(csa_tree_add_12_51_groupi_n_155 ,csa_tree_add_12_51_groupi_n_154);
  not csa_tree_add_12_51_groupi_drc_bufs25314(csa_tree_add_12_51_groupi_n_154 ,csa_tree_add_12_51_groupi_n_1968);
  not csa_tree_add_12_51_groupi_drc_bufs25316(csa_tree_add_12_51_groupi_n_153 ,csa_tree_add_12_51_groupi_n_152);
  not csa_tree_add_12_51_groupi_drc_bufs25318(csa_tree_add_12_51_groupi_n_152 ,csa_tree_add_12_51_groupi_n_1971);
  not csa_tree_add_12_51_groupi_drc_bufs25320(csa_tree_add_12_51_groupi_n_151 ,csa_tree_add_12_51_groupi_n_150);
  not csa_tree_add_12_51_groupi_drc_bufs25322(csa_tree_add_12_51_groupi_n_150 ,csa_tree_add_12_51_groupi_n_1983);
  not csa_tree_add_12_51_groupi_drc_bufs25324(csa_tree_add_12_51_groupi_n_149 ,csa_tree_add_12_51_groupi_n_147);
  not csa_tree_add_12_51_groupi_drc_bufs25325(csa_tree_add_12_51_groupi_n_148 ,csa_tree_add_12_51_groupi_n_147);
  not csa_tree_add_12_51_groupi_drc_bufs25326(csa_tree_add_12_51_groupi_n_147 ,csa_tree_add_12_51_groupi_n_2206);
  not csa_tree_add_12_51_groupi_drc_bufs25328(csa_tree_add_12_51_groupi_n_146 ,csa_tree_add_12_51_groupi_n_144);
  not csa_tree_add_12_51_groupi_drc_bufs25329(csa_tree_add_12_51_groupi_n_145 ,csa_tree_add_12_51_groupi_n_144);
  not csa_tree_add_12_51_groupi_drc_bufs25330(csa_tree_add_12_51_groupi_n_144 ,csa_tree_add_12_51_groupi_n_2207);
  not csa_tree_add_12_51_groupi_drc_bufs25332(csa_tree_add_12_51_groupi_n_143 ,csa_tree_add_12_51_groupi_n_141);
  not csa_tree_add_12_51_groupi_drc_bufs25333(csa_tree_add_12_51_groupi_n_142 ,csa_tree_add_12_51_groupi_n_141);
  not csa_tree_add_12_51_groupi_drc_bufs25334(csa_tree_add_12_51_groupi_n_141 ,csa_tree_add_12_51_groupi_n_2211);
  not csa_tree_add_12_51_groupi_drc_bufs25336(csa_tree_add_12_51_groupi_n_140 ,csa_tree_add_12_51_groupi_n_138);
  not csa_tree_add_12_51_groupi_drc_bufs25337(csa_tree_add_12_51_groupi_n_139 ,csa_tree_add_12_51_groupi_n_138);
  not csa_tree_add_12_51_groupi_drc_bufs25338(csa_tree_add_12_51_groupi_n_138 ,csa_tree_add_12_51_groupi_n_2205);
  not csa_tree_add_12_51_groupi_drc_bufs25340(csa_tree_add_12_51_groupi_n_137 ,csa_tree_add_12_51_groupi_n_135);
  not csa_tree_add_12_51_groupi_drc_bufs25341(csa_tree_add_12_51_groupi_n_136 ,csa_tree_add_12_51_groupi_n_135);
  not csa_tree_add_12_51_groupi_drc_bufs25342(csa_tree_add_12_51_groupi_n_135 ,csa_tree_add_12_51_groupi_n_2204);
  not csa_tree_add_12_51_groupi_drc_bufs25344(csa_tree_add_12_51_groupi_n_134 ,csa_tree_add_12_51_groupi_n_132);
  not csa_tree_add_12_51_groupi_drc_bufs25345(csa_tree_add_12_51_groupi_n_133 ,csa_tree_add_12_51_groupi_n_132);
  not csa_tree_add_12_51_groupi_drc_bufs25346(csa_tree_add_12_51_groupi_n_132 ,csa_tree_add_12_51_groupi_n_2204);
  not csa_tree_add_12_51_groupi_drc_bufs25348(csa_tree_add_12_51_groupi_n_131 ,csa_tree_add_12_51_groupi_n_129);
  not csa_tree_add_12_51_groupi_drc_bufs25349(csa_tree_add_12_51_groupi_n_130 ,csa_tree_add_12_51_groupi_n_129);
  not csa_tree_add_12_51_groupi_drc_bufs25350(csa_tree_add_12_51_groupi_n_129 ,csa_tree_add_12_51_groupi_n_2205);
  not csa_tree_add_12_51_groupi_drc_bufs25352(csa_tree_add_12_51_groupi_n_128 ,csa_tree_add_12_51_groupi_n_126);
  not csa_tree_add_12_51_groupi_drc_bufs25353(csa_tree_add_12_51_groupi_n_127 ,csa_tree_add_12_51_groupi_n_126);
  not csa_tree_add_12_51_groupi_drc_bufs25354(csa_tree_add_12_51_groupi_n_126 ,csa_tree_add_12_51_groupi_n_2206);
  not csa_tree_add_12_51_groupi_drc_bufs25357(csa_tree_add_12_51_groupi_n_125 ,csa_tree_add_12_51_groupi_n_124);
  not csa_tree_add_12_51_groupi_drc_bufs25358(csa_tree_add_12_51_groupi_n_124 ,csa_tree_add_12_51_groupi_n_2398);
  not csa_tree_add_12_51_groupi_drc_bufs25360(csa_tree_add_12_51_groupi_n_123 ,csa_tree_add_12_51_groupi_n_121);
  not csa_tree_add_12_51_groupi_drc_bufs25361(csa_tree_add_12_51_groupi_n_122 ,csa_tree_add_12_51_groupi_n_121);
  not csa_tree_add_12_51_groupi_drc_bufs25362(csa_tree_add_12_51_groupi_n_121 ,csa_tree_add_12_51_groupi_n_2364);
  not csa_tree_add_12_51_groupi_drc_bufs25364(csa_tree_add_12_51_groupi_n_120 ,csa_tree_add_12_51_groupi_n_119);
  not csa_tree_add_12_51_groupi_drc_bufs25366(csa_tree_add_12_51_groupi_n_119 ,csa_tree_add_12_51_groupi_n_2363);
  not csa_tree_add_12_51_groupi_drc_bufs25368(csa_tree_add_12_51_groupi_n_118 ,csa_tree_add_12_51_groupi_n_116);
  not csa_tree_add_12_51_groupi_drc_bufs25369(csa_tree_add_12_51_groupi_n_117 ,csa_tree_add_12_51_groupi_n_116);
  not csa_tree_add_12_51_groupi_drc_bufs25370(csa_tree_add_12_51_groupi_n_116 ,csa_tree_add_12_51_groupi_n_2399);
  not csa_tree_add_12_51_groupi_drc_bufs25372(csa_tree_add_12_51_groupi_n_115 ,csa_tree_add_12_51_groupi_n_113);
  not csa_tree_add_12_51_groupi_drc_bufs25373(csa_tree_add_12_51_groupi_n_114 ,csa_tree_add_12_51_groupi_n_113);
  not csa_tree_add_12_51_groupi_drc_bufs25374(csa_tree_add_12_51_groupi_n_113 ,csa_tree_add_12_51_groupi_n_2397);
  not csa_tree_add_12_51_groupi_drc_bufs25376(csa_tree_add_12_51_groupi_n_112 ,csa_tree_add_12_51_groupi_n_111);
  not csa_tree_add_12_51_groupi_drc_bufs25378(csa_tree_add_12_51_groupi_n_111 ,csa_tree_add_12_51_groupi_n_2403);
  not csa_tree_add_12_51_groupi_drc_bufs25380(csa_tree_add_12_51_groupi_n_110 ,csa_tree_add_12_51_groupi_n_109);
  not csa_tree_add_12_51_groupi_drc_bufs25382(csa_tree_add_12_51_groupi_n_109 ,csa_tree_add_12_51_groupi_n_2399);
  not csa_tree_add_12_51_groupi_drc_bufs25384(csa_tree_add_12_51_groupi_n_108 ,csa_tree_add_12_51_groupi_n_107);
  not csa_tree_add_12_51_groupi_drc_bufs25386(csa_tree_add_12_51_groupi_n_107 ,csa_tree_add_12_51_groupi_n_2404);
  not csa_tree_add_12_51_groupi_drc_bufs25388(csa_tree_add_12_51_groupi_n_106 ,csa_tree_add_12_51_groupi_n_105);
  not csa_tree_add_12_51_groupi_drc_bufs25390(csa_tree_add_12_51_groupi_n_105 ,csa_tree_add_12_51_groupi_n_1959);
  not csa_tree_add_12_51_groupi_drc_bufs25392(csa_tree_add_12_51_groupi_n_104 ,csa_tree_add_12_51_groupi_n_103);
  not csa_tree_add_12_51_groupi_drc_bufs25394(csa_tree_add_12_51_groupi_n_103 ,csa_tree_add_12_51_groupi_n_1942);
  not csa_tree_add_12_51_groupi_drc_bufs25396(csa_tree_add_12_51_groupi_n_102 ,csa_tree_add_12_51_groupi_n_101);
  not csa_tree_add_12_51_groupi_drc_bufs25398(csa_tree_add_12_51_groupi_n_101 ,csa_tree_add_12_51_groupi_n_2364);
  not csa_tree_add_12_51_groupi_drc_bufs25400(csa_tree_add_12_51_groupi_n_100 ,csa_tree_add_12_51_groupi_n_99);
  not csa_tree_add_12_51_groupi_drc_bufs25402(csa_tree_add_12_51_groupi_n_99 ,csa_tree_add_12_51_groupi_n_1960);
  not csa_tree_add_12_51_groupi_drc_bufs25404(csa_tree_add_12_51_groupi_n_98 ,csa_tree_add_12_51_groupi_n_97);
  not csa_tree_add_12_51_groupi_drc_bufs25406(csa_tree_add_12_51_groupi_n_97 ,csa_tree_add_12_51_groupi_n_2400);
  not csa_tree_add_12_51_groupi_drc_bufs25408(csa_tree_add_12_51_groupi_n_96 ,csa_tree_add_12_51_groupi_n_95);
  not csa_tree_add_12_51_groupi_drc_bufs25410(csa_tree_add_12_51_groupi_n_95 ,csa_tree_add_12_51_groupi_n_1945);
  not csa_tree_add_12_51_groupi_drc_bufs25412(csa_tree_add_12_51_groupi_n_94 ,csa_tree_add_12_51_groupi_n_93);
  not csa_tree_add_12_51_groupi_drc_bufs25414(csa_tree_add_12_51_groupi_n_93 ,csa_tree_add_12_51_groupi_n_1890);
  not csa_tree_add_12_51_groupi_drc_bufs25416(csa_tree_add_12_51_groupi_n_92 ,csa_tree_add_12_51_groupi_n_91);
  not csa_tree_add_12_51_groupi_drc_bufs25418(csa_tree_add_12_51_groupi_n_91 ,csa_tree_add_12_51_groupi_n_1887);
  not csa_tree_add_12_51_groupi_drc_bufs25420(csa_tree_add_12_51_groupi_n_90 ,csa_tree_add_12_51_groupi_n_89);
  not csa_tree_add_12_51_groupi_drc_bufs25422(csa_tree_add_12_51_groupi_n_89 ,csa_tree_add_12_51_groupi_n_1881);
  not csa_tree_add_12_51_groupi_drc_bufs25424(csa_tree_add_12_51_groupi_n_88 ,csa_tree_add_12_51_groupi_n_87);
  not csa_tree_add_12_51_groupi_drc_bufs25426(csa_tree_add_12_51_groupi_n_87 ,csa_tree_add_12_51_groupi_n_1869);
  not csa_tree_add_12_51_groupi_drc_bufs25428(csa_tree_add_12_51_groupi_n_86 ,csa_tree_add_12_51_groupi_n_85);
  not csa_tree_add_12_51_groupi_drc_bufs25430(csa_tree_add_12_51_groupi_n_85 ,csa_tree_add_12_51_groupi_n_1866);
  not csa_tree_add_12_51_groupi_drc_bufs25432(csa_tree_add_12_51_groupi_n_84 ,csa_tree_add_12_51_groupi_n_83);
  not csa_tree_add_12_51_groupi_drc_bufs25434(csa_tree_add_12_51_groupi_n_83 ,csa_tree_add_12_51_groupi_n_1878);
  not csa_tree_add_12_51_groupi_drc_bufs25436(csa_tree_add_12_51_groupi_n_82 ,csa_tree_add_12_51_groupi_n_81);
  not csa_tree_add_12_51_groupi_drc_bufs25438(csa_tree_add_12_51_groupi_n_81 ,csa_tree_add_12_51_groupi_n_1863);
  not csa_tree_add_12_51_groupi_drc_bufs25440(csa_tree_add_12_51_groupi_n_80 ,csa_tree_add_12_51_groupi_n_79);
  not csa_tree_add_12_51_groupi_drc_bufs25442(csa_tree_add_12_51_groupi_n_79 ,csa_tree_add_12_51_groupi_n_1860);
  not csa_tree_add_12_51_groupi_drc_bufs25444(csa_tree_add_12_51_groupi_n_78 ,csa_tree_add_12_51_groupi_n_77);
  not csa_tree_add_12_51_groupi_drc_bufs25446(csa_tree_add_12_51_groupi_n_77 ,csa_tree_add_12_51_groupi_n_1884);
  not csa_tree_add_12_51_groupi_drc_bufs25448(csa_tree_add_12_51_groupi_n_76 ,csa_tree_add_12_51_groupi_n_75);
  not csa_tree_add_12_51_groupi_drc_bufs25450(csa_tree_add_12_51_groupi_n_75 ,csa_tree_add_12_51_groupi_n_1875);
  not csa_tree_add_12_51_groupi_drc_bufs25452(csa_tree_add_12_51_groupi_n_74 ,csa_tree_add_12_51_groupi_n_73);
  not csa_tree_add_12_51_groupi_drc_bufs25454(csa_tree_add_12_51_groupi_n_73 ,csa_tree_add_12_51_groupi_n_1857);
  not csa_tree_add_12_51_groupi_drc_bufs25456(csa_tree_add_12_51_groupi_n_72 ,csa_tree_add_12_51_groupi_n_71);
  not csa_tree_add_12_51_groupi_drc_bufs25458(csa_tree_add_12_51_groupi_n_71 ,csa_tree_add_12_51_groupi_n_1854);
  not csa_tree_add_12_51_groupi_drc_bufs25460(csa_tree_add_12_51_groupi_n_70 ,csa_tree_add_12_51_groupi_n_69);
  not csa_tree_add_12_51_groupi_drc_bufs25462(csa_tree_add_12_51_groupi_n_69 ,csa_tree_add_12_51_groupi_n_1872);
  not csa_tree_add_12_51_groupi_drc_bufs25464(csa_tree_add_12_51_groupi_n_68 ,csa_tree_add_12_51_groupi_n_67);
  not csa_tree_add_12_51_groupi_drc_bufs25466(csa_tree_add_12_51_groupi_n_67 ,csa_tree_add_12_51_groupi_n_1851);
  not csa_tree_add_12_51_groupi_drc_bufs25468(csa_tree_add_12_51_groupi_n_66 ,csa_tree_add_12_51_groupi_n_65);
  not csa_tree_add_12_51_groupi_drc_bufs25470(csa_tree_add_12_51_groupi_n_65 ,csa_tree_add_12_51_groupi_n_1848);
  not csa_tree_add_12_51_groupi_drc_bufs25472(csa_tree_add_12_51_groupi_n_64 ,csa_tree_add_12_51_groupi_n_62);
  not csa_tree_add_12_51_groupi_drc_bufs25473(csa_tree_add_12_51_groupi_n_63 ,csa_tree_add_12_51_groupi_n_62);
  not csa_tree_add_12_51_groupi_drc_bufs25474(csa_tree_add_12_51_groupi_n_62 ,csa_tree_add_12_51_groupi_n_2143);
  not csa_tree_add_12_51_groupi_drc_bufs25476(csa_tree_add_12_51_groupi_n_61 ,csa_tree_add_12_51_groupi_n_59);
  not csa_tree_add_12_51_groupi_drc_bufs25477(csa_tree_add_12_51_groupi_n_60 ,csa_tree_add_12_51_groupi_n_59);
  not csa_tree_add_12_51_groupi_drc_bufs25478(csa_tree_add_12_51_groupi_n_59 ,csa_tree_add_12_51_groupi_n_2119);
  not csa_tree_add_12_51_groupi_drc_bufs25480(csa_tree_add_12_51_groupi_n_58 ,csa_tree_add_12_51_groupi_n_56);
  not csa_tree_add_12_51_groupi_drc_bufs25481(csa_tree_add_12_51_groupi_n_57 ,csa_tree_add_12_51_groupi_n_56);
  not csa_tree_add_12_51_groupi_drc_bufs25482(csa_tree_add_12_51_groupi_n_56 ,csa_tree_add_12_51_groupi_n_2134);
  not csa_tree_add_12_51_groupi_drc_bufs25484(csa_tree_add_12_51_groupi_n_55 ,csa_tree_add_12_51_groupi_n_53);
  not csa_tree_add_12_51_groupi_drc_bufs25485(csa_tree_add_12_51_groupi_n_54 ,csa_tree_add_12_51_groupi_n_53);
  not csa_tree_add_12_51_groupi_drc_bufs25486(csa_tree_add_12_51_groupi_n_53 ,csa_tree_add_12_51_groupi_n_2131);
  not csa_tree_add_12_51_groupi_drc_bufs25488(csa_tree_add_12_51_groupi_n_52 ,csa_tree_add_12_51_groupi_n_50);
  not csa_tree_add_12_51_groupi_drc_bufs25489(csa_tree_add_12_51_groupi_n_51 ,csa_tree_add_12_51_groupi_n_50);
  not csa_tree_add_12_51_groupi_drc_bufs25490(csa_tree_add_12_51_groupi_n_50 ,csa_tree_add_12_51_groupi_n_2125);
  not csa_tree_add_12_51_groupi_drc_bufs25492(csa_tree_add_12_51_groupi_n_49 ,csa_tree_add_12_51_groupi_n_47);
  not csa_tree_add_12_51_groupi_drc_bufs25493(csa_tree_add_12_51_groupi_n_48 ,csa_tree_add_12_51_groupi_n_47);
  not csa_tree_add_12_51_groupi_drc_bufs25494(csa_tree_add_12_51_groupi_n_47 ,csa_tree_add_12_51_groupi_n_2122);
  not csa_tree_add_12_51_groupi_drc_bufs25496(csa_tree_add_12_51_groupi_n_46 ,csa_tree_add_12_51_groupi_n_44);
  not csa_tree_add_12_51_groupi_drc_bufs25497(csa_tree_add_12_51_groupi_n_45 ,csa_tree_add_12_51_groupi_n_44);
  not csa_tree_add_12_51_groupi_drc_bufs25498(csa_tree_add_12_51_groupi_n_44 ,csa_tree_add_12_51_groupi_n_2113);
  not csa_tree_add_12_51_groupi_drc_bufs25500(csa_tree_add_12_51_groupi_n_43 ,csa_tree_add_12_51_groupi_n_41);
  not csa_tree_add_12_51_groupi_drc_bufs25501(csa_tree_add_12_51_groupi_n_42 ,csa_tree_add_12_51_groupi_n_41);
  not csa_tree_add_12_51_groupi_drc_bufs25502(csa_tree_add_12_51_groupi_n_41 ,csa_tree_add_12_51_groupi_n_2110);
  not csa_tree_add_12_51_groupi_drc_bufs25504(csa_tree_add_12_51_groupi_n_40 ,csa_tree_add_12_51_groupi_n_38);
  not csa_tree_add_12_51_groupi_drc_bufs25505(csa_tree_add_12_51_groupi_n_39 ,csa_tree_add_12_51_groupi_n_38);
  not csa_tree_add_12_51_groupi_drc_bufs25506(csa_tree_add_12_51_groupi_n_38 ,csa_tree_add_12_51_groupi_n_2149);
  not csa_tree_add_12_51_groupi_drc_bufs25508(csa_tree_add_12_51_groupi_n_37 ,csa_tree_add_12_51_groupi_n_35);
  not csa_tree_add_12_51_groupi_drc_bufs25509(csa_tree_add_12_51_groupi_n_36 ,csa_tree_add_12_51_groupi_n_35);
  not csa_tree_add_12_51_groupi_drc_bufs25510(csa_tree_add_12_51_groupi_n_35 ,csa_tree_add_12_51_groupi_n_2107);
  not csa_tree_add_12_51_groupi_drc_bufs25512(csa_tree_add_12_51_groupi_n_34 ,csa_tree_add_12_51_groupi_n_32);
  not csa_tree_add_12_51_groupi_drc_bufs25513(csa_tree_add_12_51_groupi_n_33 ,csa_tree_add_12_51_groupi_n_32);
  not csa_tree_add_12_51_groupi_drc_bufs25514(csa_tree_add_12_51_groupi_n_32 ,csa_tree_add_12_51_groupi_n_2137);
  not csa_tree_add_12_51_groupi_drc_bufs25516(csa_tree_add_12_51_groupi_n_31 ,csa_tree_add_12_51_groupi_n_29);
  not csa_tree_add_12_51_groupi_drc_bufs25517(csa_tree_add_12_51_groupi_n_30 ,csa_tree_add_12_51_groupi_n_29);
  not csa_tree_add_12_51_groupi_drc_bufs25518(csa_tree_add_12_51_groupi_n_29 ,csa_tree_add_12_51_groupi_n_2128);
  not csa_tree_add_12_51_groupi_drc_bufs25520(csa_tree_add_12_51_groupi_n_28 ,csa_tree_add_12_51_groupi_n_26);
  not csa_tree_add_12_51_groupi_drc_bufs25521(csa_tree_add_12_51_groupi_n_27 ,csa_tree_add_12_51_groupi_n_26);
  not csa_tree_add_12_51_groupi_drc_bufs25522(csa_tree_add_12_51_groupi_n_26 ,csa_tree_add_12_51_groupi_n_2116);
  not csa_tree_add_12_51_groupi_drc_bufs25524(csa_tree_add_12_51_groupi_n_25 ,csa_tree_add_12_51_groupi_n_23);
  not csa_tree_add_12_51_groupi_drc_bufs25525(csa_tree_add_12_51_groupi_n_24 ,csa_tree_add_12_51_groupi_n_23);
  not csa_tree_add_12_51_groupi_drc_bufs25526(csa_tree_add_12_51_groupi_n_23 ,csa_tree_add_12_51_groupi_n_2146);
  not csa_tree_add_12_51_groupi_drc_bufs25528(csa_tree_add_12_51_groupi_n_22 ,csa_tree_add_12_51_groupi_n_20);
  not csa_tree_add_12_51_groupi_drc_bufs25529(csa_tree_add_12_51_groupi_n_21 ,csa_tree_add_12_51_groupi_n_20);
  not csa_tree_add_12_51_groupi_drc_bufs25530(csa_tree_add_12_51_groupi_n_20 ,csa_tree_add_12_51_groupi_n_2140);
  not csa_tree_add_12_51_groupi_drc_bufs25533(csa_tree_add_12_51_groupi_n_19 ,csa_tree_add_12_51_groupi_n_18);
  not csa_tree_add_12_51_groupi_drc_bufs25534(csa_tree_add_12_51_groupi_n_18 ,csa_tree_add_12_51_groupi_n_1814);
  xor csa_tree_add_12_51_groupi_g2(csa_tree_add_12_51_groupi_n_17 ,csa_tree_add_12_51_groupi_n_6756 ,csa_tree_add_12_51_groupi_n_6847);
  xor csa_tree_add_12_51_groupi_g25536(csa_tree_add_12_51_groupi_n_16 ,csa_tree_add_12_51_groupi_n_6749 ,csa_tree_add_12_51_groupi_n_6992);
  xor csa_tree_add_12_51_groupi_g25537(csa_tree_add_12_51_groupi_n_15 ,csa_tree_add_12_51_groupi_n_6447 ,csa_tree_add_12_51_groupi_n_6693);
  xor csa_tree_add_12_51_groupi_g25538(csa_tree_add_12_51_groupi_n_14 ,csa_tree_add_12_51_groupi_n_6063 ,csa_tree_add_12_51_groupi_n_6251);
  xor csa_tree_add_12_51_groupi_g25539(csa_tree_add_12_51_groupi_n_13 ,csa_tree_add_12_51_groupi_n_5755 ,csa_tree_add_12_51_groupi_n_5888);
  xor csa_tree_add_12_51_groupi_g25540(csa_tree_add_12_51_groupi_n_12 ,csa_tree_add_12_51_groupi_n_3530 ,csa_tree_add_12_51_groupi_n_1913);
  xor csa_tree_add_12_51_groupi_g25541(csa_tree_add_12_51_groupi_n_11 ,csa_tree_add_12_51_groupi_n_3247 ,csa_tree_add_12_51_groupi_n_1911);
  xor csa_tree_add_12_51_groupi_g25542(csa_tree_add_12_51_groupi_n_10 ,csa_tree_add_12_51_groupi_n_3529 ,csa_tree_add_12_51_groupi_n_1909);
  xor csa_tree_add_12_51_groupi_g25543(csa_tree_add_12_51_groupi_n_9 ,csa_tree_add_12_51_groupi_n_4782 ,csa_tree_add_12_51_groupi_n_1900);
  xor csa_tree_add_12_51_groupi_g25544(csa_tree_add_12_51_groupi_n_8 ,csa_tree_add_12_51_groupi_n_1893 ,csa_tree_add_12_51_groupi_n_3996);
  xor csa_tree_add_12_51_groupi_g25545(csa_tree_add_12_51_groupi_n_7 ,csa_tree_add_12_51_groupi_n_1891 ,csa_tree_add_12_51_groupi_n_3774);
  xor csa_tree_add_12_51_groupi_g25546(csa_tree_add_12_51_groupi_n_6 ,csa_tree_add_12_51_groupi_n_5117 ,csa_tree_add_12_51_groupi_n_124);
  xor csa_tree_add_12_51_groupi_g25547(csa_tree_add_12_51_groupi_n_5 ,csa_tree_add_12_51_groupi_n_119 ,csa_tree_add_12_51_groupi_n_3998);
  xor csa_tree_add_12_51_groupi_g25548(csa_tree_add_12_51_groupi_n_4 ,csa_tree_add_12_51_groupi_n_111 ,csa_tree_add_12_51_groupi_n_5608);
  xor csa_tree_add_12_51_groupi_g25549(csa_tree_add_12_51_groupi_n_3 ,csa_tree_add_12_51_groupi_n_109 ,csa_tree_add_12_51_groupi_n_4602);
  xor csa_tree_add_12_51_groupi_g25550(csa_tree_add_12_51_groupi_n_2 ,csa_tree_add_12_51_groupi_n_107 ,csa_tree_add_12_51_groupi_n_5120);
  xor csa_tree_add_12_51_groupi_g25551(csa_tree_add_12_51_groupi_n_1 ,csa_tree_add_12_51_groupi_n_101 ,csa_tree_add_12_51_groupi_n_4422);
  xor csa_tree_add_12_51_groupi_g25552(csa_tree_add_12_51_groupi_n_0 ,csa_tree_add_12_51_groupi_n_97 ,csa_tree_add_12_51_groupi_n_5605);
  xnor sub_11_21_g407(out2[16] ,sub_11_21_n_141 ,out1[16]);
  or sub_11_21_g408(sub_11_21_n_141 ,sub_11_21_n_0 ,sub_11_21_n_139);
  xnor sub_11_21_g409(out2[15] ,sub_11_21_n_138 ,sub_11_21_n_85);
  nor sub_11_21_g410(sub_11_21_n_139 ,sub_11_21_n_73 ,sub_11_21_n_138);
  and sub_11_21_g411(sub_11_21_n_138 ,sub_11_21_n_63 ,sub_11_21_n_136);
  xnor sub_11_21_g412(out2[14] ,sub_11_21_n_135 ,sub_11_21_n_84);
  or sub_11_21_g413(sub_11_21_n_136 ,sub_11_21_n_56 ,sub_11_21_n_135);
  and sub_11_21_g414(sub_11_21_n_135 ,sub_11_21_n_74 ,sub_11_21_n_133);
  xnor sub_11_21_g415(out2[13] ,sub_11_21_n_132 ,sub_11_21_n_83);
  or sub_11_21_g416(sub_11_21_n_133 ,sub_11_21_n_65 ,sub_11_21_n_132);
  and sub_11_21_g417(sub_11_21_n_132 ,sub_11_21_n_78 ,sub_11_21_n_130);
  xnor sub_11_21_g418(out2[12] ,sub_11_21_n_129 ,sub_11_21_n_82);
  or sub_11_21_g419(sub_11_21_n_130 ,sub_11_21_n_58 ,sub_11_21_n_129);
  and sub_11_21_g420(sub_11_21_n_129 ,sub_11_21_n_53 ,sub_11_21_n_127);
  xnor sub_11_21_g421(out2[11] ,sub_11_21_n_126 ,sub_11_21_n_89);
  or sub_11_21_g422(sub_11_21_n_127 ,sub_11_21_n_77 ,sub_11_21_n_126);
  and sub_11_21_g423(sub_11_21_n_126 ,sub_11_21_n_71 ,sub_11_21_n_124);
  xnor sub_11_21_g424(out2[10] ,sub_11_21_n_123 ,sub_11_21_n_95);
  or sub_11_21_g425(sub_11_21_n_124 ,sub_11_21_n_67 ,sub_11_21_n_123);
  and sub_11_21_g426(sub_11_21_n_123 ,sub_11_21_n_75 ,sub_11_21_n_121);
  xnor sub_11_21_g427(out2[9] ,sub_11_21_n_120 ,sub_11_21_n_94);
  or sub_11_21_g428(sub_11_21_n_121 ,sub_11_21_n_64 ,sub_11_21_n_120);
  and sub_11_21_g429(sub_11_21_n_120 ,sub_11_21_n_62 ,sub_11_21_n_118);
  xnor sub_11_21_g430(out2[8] ,sub_11_21_n_117 ,sub_11_21_n_93);
  or sub_11_21_g431(sub_11_21_n_118 ,sub_11_21_n_59 ,sub_11_21_n_117);
  and sub_11_21_g432(sub_11_21_n_117 ,sub_11_21_n_57 ,sub_11_21_n_115);
  xnor sub_11_21_g433(out2[7] ,sub_11_21_n_114 ,sub_11_21_n_92);
  or sub_11_21_g434(sub_11_21_n_115 ,sub_11_21_n_55 ,sub_11_21_n_114);
  and sub_11_21_g435(sub_11_21_n_114 ,sub_11_21_n_72 ,sub_11_21_n_112);
  xnor sub_11_21_g436(out2[6] ,sub_11_21_n_111 ,sub_11_21_n_91);
  or sub_11_21_g437(sub_11_21_n_112 ,sub_11_21_n_66 ,sub_11_21_n_111);
  and sub_11_21_g438(sub_11_21_n_111 ,sub_11_21_n_70 ,sub_11_21_n_109);
  xnor sub_11_21_g439(out2[5] ,sub_11_21_n_108 ,sub_11_21_n_90);
  or sub_11_21_g440(sub_11_21_n_109 ,sub_11_21_n_79 ,sub_11_21_n_108);
  and sub_11_21_g441(sub_11_21_n_108 ,sub_11_21_n_68 ,sub_11_21_n_106);
  xnor sub_11_21_g442(out2[4] ,sub_11_21_n_105 ,sub_11_21_n_81);
  or sub_11_21_g443(sub_11_21_n_106 ,sub_11_21_n_69 ,sub_11_21_n_105);
  and sub_11_21_g444(sub_11_21_n_105 ,sub_11_21_n_51 ,sub_11_21_n_103);
  xnor sub_11_21_g445(out2[3] ,sub_11_21_n_102 ,sub_11_21_n_88);
  or sub_11_21_g446(sub_11_21_n_103 ,sub_11_21_n_76 ,sub_11_21_n_102);
  and sub_11_21_g447(sub_11_21_n_102 ,sub_11_21_n_52 ,sub_11_21_n_100);
  xnor sub_11_21_g448(out2[2] ,sub_11_21_n_98 ,sub_11_21_n_87);
  or sub_11_21_g449(sub_11_21_n_100 ,sub_11_21_n_54 ,sub_11_21_n_98);
  xnor sub_11_21_g450(out2[1] ,sub_11_21_n_80 ,sub_11_21_n_86);
  and sub_11_21_g451(sub_11_21_n_98 ,sub_11_21_n_61 ,sub_11_21_n_96);
  xor sub_11_21_g452(out2[0] ,out1[0] ,in3[0]);
  or sub_11_21_g453(sub_11_21_n_96 ,sub_11_21_n_60 ,sub_11_21_n_80);
  xnor sub_11_21_g454(sub_11_21_n_95 ,sub_11_21_n_17 ,in3[10]);
  xnor sub_11_21_g455(sub_11_21_n_94 ,sub_11_21_n_12 ,in3[9]);
  xnor sub_11_21_g456(sub_11_21_n_93 ,sub_11_21_n_16 ,in3[8]);
  xnor sub_11_21_g457(sub_11_21_n_92 ,sub_11_21_n_13 ,in3[7]);
  xnor sub_11_21_g458(sub_11_21_n_91 ,sub_11_21_n_6 ,in3[6]);
  xnor sub_11_21_g459(sub_11_21_n_90 ,sub_11_21_n_15 ,in3[5]);
  xnor sub_11_21_g460(sub_11_21_n_89 ,sub_11_21_n_18 ,in3[11]);
  xnor sub_11_21_g461(sub_11_21_n_88 ,sub_11_21_n_14 ,in3[3]);
  xnor sub_11_21_g462(sub_11_21_n_87 ,sub_11_21_n_20 ,in3[2]);
  xnor sub_11_21_g463(sub_11_21_n_86 ,sub_11_21_n_22 ,in3[1]);
  xnor sub_11_21_g464(sub_11_21_n_85 ,sub_11_21_n_24 ,in3[15]);
  xnor sub_11_21_g465(sub_11_21_n_84 ,sub_11_21_n_21 ,in3[14]);
  xnor sub_11_21_g466(sub_11_21_n_83 ,sub_11_21_n_3 ,in3[13]);
  xnor sub_11_21_g467(sub_11_21_n_82 ,sub_11_21_n_9 ,in3[12]);
  xnor sub_11_21_g468(sub_11_21_n_81 ,sub_11_21_n_19 ,in3[4]);
  nor sub_11_21_g469(sub_11_21_n_79 ,sub_11_21_n_33 ,in3[5]);
  or sub_11_21_g470(sub_11_21_n_78 ,sub_11_21_n_39 ,sub_11_21_n_8);
  nor sub_11_21_g472(sub_11_21_n_77 ,sub_11_21_n_27 ,in3[11]);
  nor sub_11_21_g473(sub_11_21_n_76 ,sub_11_21_n_31 ,in3[3]);
  or sub_11_21_g474(sub_11_21_n_75 ,sub_11_21_n_37 ,sub_11_21_n_11);
  or sub_11_21_g475(sub_11_21_n_74 ,sub_11_21_n_38 ,sub_11_21_n_2);
  nor sub_11_21_g476(sub_11_21_n_73 ,sub_11_21_n_41 ,in3[15]);
  or sub_11_21_g477(sub_11_21_n_72 ,sub_11_21_n_47 ,sub_11_21_n_5);
  or sub_11_21_g478(sub_11_21_n_71 ,sub_11_21_n_49 ,sub_11_21_n_17);
  or sub_11_21_g479(sub_11_21_n_70 ,sub_11_21_n_40 ,sub_11_21_n_15);
  nor sub_11_21_g480(sub_11_21_n_69 ,sub_11_21_n_26 ,in3[4]);
  or sub_11_21_g481(sub_11_21_n_68 ,sub_11_21_n_36 ,sub_11_21_n_19);
  nor sub_11_21_g482(sub_11_21_n_67 ,sub_11_21_n_29 ,in3[10]);
  and sub_11_21_g483(sub_11_21_n_80 ,out1[0] ,sub_11_21_n_50);
  and sub_11_21_g484(sub_11_21_n_66 ,sub_11_21_n_6 ,sub_11_21_n_47);
  and sub_11_21_g485(sub_11_21_n_65 ,sub_11_21_n_3 ,sub_11_21_n_38);
  and sub_11_21_g486(sub_11_21_n_64 ,sub_11_21_n_12 ,sub_11_21_n_37);
  or sub_11_21_g487(sub_11_21_n_63 ,sub_11_21_n_48 ,sub_11_21_n_21);
  or sub_11_21_g488(sub_11_21_n_62 ,sub_11_21_n_43 ,sub_11_21_n_16);
  or sub_11_21_g489(sub_11_21_n_61 ,sub_11_21_n_44 ,sub_11_21_n_22);
  nor sub_11_21_g490(sub_11_21_n_60 ,sub_11_21_n_30 ,in3[1]);
  nor sub_11_21_g491(sub_11_21_n_59 ,sub_11_21_n_28 ,in3[8]);
  and sub_11_21_g492(sub_11_21_n_58 ,sub_11_21_n_9 ,sub_11_21_n_39);
  or sub_11_21_g493(sub_11_21_n_57 ,sub_11_21_n_35 ,sub_11_21_n_13);
  nor sub_11_21_g494(sub_11_21_n_56 ,sub_11_21_n_34 ,in3[14]);
  nor sub_11_21_g495(sub_11_21_n_55 ,sub_11_21_n_32 ,in3[7]);
  nor sub_11_21_g496(sub_11_21_n_54 ,sub_11_21_n_25 ,in3[2]);
  or sub_11_21_g497(sub_11_21_n_53 ,sub_11_21_n_42 ,sub_11_21_n_18);
  or sub_11_21_g498(sub_11_21_n_52 ,sub_11_21_n_46 ,sub_11_21_n_20);
  or sub_11_21_g499(sub_11_21_n_51 ,sub_11_21_n_45 ,sub_11_21_n_14);
  not sub_11_21_g500(sub_11_21_n_50 ,in3[0]);
  not sub_11_21_g501(sub_11_21_n_49 ,in3[10]);
  not sub_11_21_g502(sub_11_21_n_48 ,in3[14]);
  not sub_11_21_g503(sub_11_21_n_47 ,in3[6]);
  not sub_11_21_g504(sub_11_21_n_46 ,in3[2]);
  not sub_11_21_g505(sub_11_21_n_45 ,in3[3]);
  not sub_11_21_g507(sub_11_21_n_44 ,in3[1]);
  not sub_11_21_g509(sub_11_21_n_43 ,in3[8]);
  not sub_11_21_g512(sub_11_21_n_42 ,in3[11]);
  not sub_11_21_g514(sub_11_21_n_41 ,sub_11_21_n_24);
  not sub_11_21_g516(sub_11_21_n_40 ,in3[5]);
  not sub_11_21_g518(sub_11_21_n_39 ,in3[12]);
  not sub_11_21_g520(sub_11_21_n_38 ,in3[13]);
  not sub_11_21_g521(sub_11_21_n_37 ,in3[9]);
  not sub_11_21_g524(sub_11_21_n_36 ,in3[4]);
  not sub_11_21_g526(sub_11_21_n_35 ,in3[7]);
  not sub_11_21_drc_bufs(sub_11_21_n_24 ,sub_11_21_n_23);
  not sub_11_21_drc_bufs528(sub_11_21_n_23 ,out1[15]);
  not sub_11_21_drc_bufs531(sub_11_21_n_22 ,sub_11_21_n_30);
  not sub_11_21_drc_bufs532(sub_11_21_n_30 ,out1[1]);
  not sub_11_21_drc_bufs535(sub_11_21_n_21 ,sub_11_21_n_34);
  not sub_11_21_drc_bufs536(sub_11_21_n_34 ,out1[14]);
  not sub_11_21_drc_bufs539(sub_11_21_n_20 ,sub_11_21_n_25);
  not sub_11_21_drc_bufs540(sub_11_21_n_25 ,out1[2]);
  not sub_11_21_drc_bufs543(sub_11_21_n_19 ,sub_11_21_n_26);
  not sub_11_21_drc_bufs544(sub_11_21_n_26 ,out1[4]);
  not sub_11_21_drc_bufs547(sub_11_21_n_18 ,sub_11_21_n_27);
  not sub_11_21_drc_bufs548(sub_11_21_n_27 ,out1[11]);
  not sub_11_21_drc_bufs551(sub_11_21_n_17 ,sub_11_21_n_29);
  not sub_11_21_drc_bufs552(sub_11_21_n_29 ,out1[10]);
  not sub_11_21_drc_bufs555(sub_11_21_n_16 ,sub_11_21_n_28);
  not sub_11_21_drc_bufs556(sub_11_21_n_28 ,out1[8]);
  not sub_11_21_drc_bufs559(sub_11_21_n_15 ,sub_11_21_n_33);
  not sub_11_21_drc_bufs560(sub_11_21_n_33 ,out1[5]);
  not sub_11_21_drc_bufs563(sub_11_21_n_14 ,sub_11_21_n_31);
  not sub_11_21_drc_bufs564(sub_11_21_n_31 ,out1[3]);
  not sub_11_21_drc_bufs567(sub_11_21_n_13 ,sub_11_21_n_32);
  not sub_11_21_drc_bufs568(sub_11_21_n_32 ,out1[7]);
  not sub_11_21_drc_bufs570(sub_11_21_n_12 ,sub_11_21_n_10);
  not sub_11_21_drc_bufs571(sub_11_21_n_11 ,sub_11_21_n_10);
  not sub_11_21_drc_bufs572(sub_11_21_n_10 ,out1[9]);
  not sub_11_21_drc_bufs574(sub_11_21_n_9 ,sub_11_21_n_7);
  not sub_11_21_drc_bufs575(sub_11_21_n_8 ,sub_11_21_n_7);
  not sub_11_21_drc_bufs576(sub_11_21_n_7 ,out1[12]);
  not sub_11_21_drc_bufs578(sub_11_21_n_6 ,sub_11_21_n_4);
  not sub_11_21_drc_bufs579(sub_11_21_n_5 ,sub_11_21_n_4);
  not sub_11_21_drc_bufs580(sub_11_21_n_4 ,out1[6]);
  not sub_11_21_drc_bufs582(sub_11_21_n_3 ,sub_11_21_n_1);
  not sub_11_21_drc_bufs583(sub_11_21_n_2 ,sub_11_21_n_1);
  not sub_11_21_drc_bufs584(sub_11_21_n_1 ,out1[13]);
  and sub_11_21_g2(sub_11_21_n_0 ,in3[15] ,sub_11_21_n_23);
endmodule
