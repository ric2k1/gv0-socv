module top( n2 , n4 , n6 , n9 , n12 , n18 , n22 , n34 , n35 , 
n42 , n48 , n51 , n56 , n57 , n65 , n67 , n68 , n72 , n75 , 
n77 , n78 , n80 );
    input n2 , n4 , n12 , n18 , n22 , n34 , n35 , n51 , n57 , 
n67 , n72 , n75 , n78 , n80 ;
    output n6 , n9 , n42 , n48 , n56 , n65 , n68 , n77 ;
    wire n0 , n1 , n3 , n5 , n7 , n8 , n10 , n11 , n13 , 
n14 , n15 , n16 , n17 , n19 , n20 , n21 , n23 , n24 , n25 , 
n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n36 , n37 , 
n38 , n39 , n40 , n41 , n43 , n44 , n45 , n46 , n47 , n49 , 
n50 , n52 , n53 , n54 , n55 , n58 , n59 , n60 , n61 , n62 , 
n63 , n64 , n66 , n69 , n70 , n71 , n73 , n74 , n76 , n79 , 
n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 ;
    or g0 ( n77 , n86 , n73 );
    xnor g1 ( n5 , n45 , n53 );
    xor g2 ( n9 , n61 , n30 );
    nor g3 ( n40 , n12 , n27 );
    not g4 ( n16 , n10 );
    not g5 ( n81 , n84 );
    and g6 ( n31 , n34 , n44 );
    or g7 ( n26 , n80 , n2 );
    and g8 ( n58 , n72 , n67 );
    not g9 ( n24 , n2 );
    or g10 ( n14 , n21 , n78 );
    and g11 ( n79 , n39 , n1 );
    or g12 ( n20 , n80 , n67 );
    nor g13 ( n7 , n84 , n76 );
    and g14 ( n52 , n72 , n57 );
    and g15 ( n50 , n28 , n36 );
    not g16 ( n15 , n45 );
    xnor g17 ( n69 , n0 , n50 );
    nand g18 ( n3 , n72 , n4 );
    and g19 ( n43 , n22 , n20 );
    and g20 ( n27 , n53 , n16 );
    not g21 ( n21 , n4 );
    or g22 ( n60 , n37 , n12 );
    and g23 ( n1 , n55 , n70 );
    not g24 ( n88 , n67 );
    and g25 ( n87 , n18 , n26 );
    not g26 ( n48 , n63 );
    not g27 ( n71 , n57 );
    xnor g28 ( n6 , n60 , n5 );
    nor g29 ( n33 , n37 , n77 );
    and g30 ( n59 , n35 , n25 );
    and g31 ( n45 , n54 , n43 );
    or g32 ( n55 , n52 , n64 );
    not g33 ( n29 , n75 );
    nor g34 ( n74 , n29 , n4 );
    or g35 ( n86 , n90 , n11 );
    or g36 ( n73 , n66 , n45 );
    xor g37 ( n42 , n40 , n69 );
    xor g38 ( n65 , n19 , n82 );
    and g39 ( n89 , n9 , n65 );
    not g40 ( n37 , n51 );
    and g41 ( n90 , n14 , n59 );
    or g42 ( n25 , n80 , n4 );
    and g43 ( n49 , n3 , n38 );
    and g44 ( n10 , n51 , n15 );
    nor g45 ( n61 , n12 , n7 );
    or g46 ( n68 , n33 , n63 );
    or g47 ( n70 , n11 , n47 );
    nor g48 ( n36 , n18 , n23 );
    or g49 ( n46 , n71 , n78 );
    nor g50 ( n32 , n90 , n1 );
    or g51 ( n39 , n11 , n81 );
    nor g52 ( n13 , n29 , n57 );
    xor g53 ( n82 , n90 , n49 );
    and g54 ( n56 , n8 , n89 );
    xnor g55 ( n30 , n11 , n55 );
    or g56 ( n41 , n22 , n83 );
    or g57 ( n54 , n88 , n78 );
    not g58 ( n17 , n72 );
    nor g59 ( n19 , n12 , n79 );
    nor g60 ( n38 , n35 , n74 );
    and g61 ( n11 , n46 , n31 );
    nor g62 ( n23 , n29 , n2 );
    or g63 ( n44 , n80 , n57 );
    or g64 ( n76 , n50 , n62 );
    and g65 ( n66 , n85 , n87 );
    or g66 ( n53 , n58 , n41 );
    or g67 ( n85 , n24 , n78 );
    nor g68 ( n83 , n29 , n67 );
    not g69 ( n0 , n66 );
    not g70 ( n47 , n76 );
    or g71 ( n63 , n49 , n32 );
    nor g72 ( n62 , n53 , n66 );
    and g73 ( n8 , n6 , n42 );
    and g74 ( n84 , n0 , n10 );
    or g75 ( n64 , n34 , n13 );
    or g76 ( n28 , n17 , n24 );
endmodule
