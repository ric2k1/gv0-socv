module a;
parameter integer [2:0]x=0;
endmodule
