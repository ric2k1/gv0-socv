module top( n0 , n2 , n17 , n18 , n23 , n24 , n26 , n27 , n29 , n37 , n43 , n58 , n59 , n61 , n66 , n70 , n73 , n75 , n80 , n81 , n84 , n86 , n88 , n89 , n90 , n91 , n94 , n98 , n104 , n107 , n123 , n129 , n130 , n133 , n137 , n145 , n151 , n160 , n164 , n168 , n169 , n174 , n179 , n187 , n194 , n196 , n199 , n210 , n211 , n212 , n213 , n214 , n217 , n221 , n226 , n234 , n237 , n238 , n246 , n249 , n253 , n256 , n260 , n261 , n265 , n272 , n278 , n281 , n286 , n289 , n292 , n304 , n310 );
    input n0 , n2 , n17 , n18 , n23 , n27 , n29 , n37 , n43 , n58 , n59 , n70 , n75 , n84 , n90 , n91 , n107 , n130 , n133 , n137 , n169 , n174 , n179 , n187 , n194 , n196 , n210 , n211 , n214 , n226 , n234 , n237 , n238 , n249 , n256 , n260 , n272 , n278 , n281 , n289 , n292 ;
    output n24 , n26 , n61 , n66 , n73 , n80 , n81 , n86 , n88 , n89 , n94 , n98 , n104 , n123 , n129 , n145 , n151 , n160 , n164 , n168 , n199 , n212 , n213 , n217 , n221 , n246 , n253 , n261 , n265 , n286 , n304 , n310 ;
    wire n1 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n19 , n20 , n21 , n22 , n25 , n28 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n38 , n39 , n40 , n41 , n42 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n60 , n62 , n63 , n64 , n65 , n67 , n68 , n69 , n71 , n72 , n74 , n76 , n77 , n78 , n79 , n82 , n83 , n85 , n87 , n92 , n93 , n95 , n96 , n97 , n99 , n100 , n101 , n102 , n103 , n105 , n106 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n124 , n125 , n126 , n127 , n128 , n131 , n132 , n134 , n135 , n136 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n146 , n147 , n148 , n149 , n150 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n161 , n162 , n163 , n165 , n166 , n167 , n170 , n171 , n172 , n173 , n175 , n176 , n177 , n178 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n188 , n189 , n190 , n191 , n192 , n193 , n195 , n197 , n198 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n215 , n216 , n218 , n219 , n220 , n222 , n223 , n224 , n225 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n235 , n236 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n247 , n248 , n250 , n251 , n252 , n254 , n255 , n257 , n258 , n259 , n262 , n263 , n264 , n266 , n267 , n268 , n269 , n270 , n271 , n273 , n274 , n275 , n276 , n277 , n279 , n280 , n282 , n283 , n284 , n285 , n287 , n288 , n290 , n291 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n305 , n306 , n307 , n308 , n309 , n311 ;
assign n163 = ~(n174 ^ n169);
assign n129 = ~(n153 ^ n210);
assign n53 = n205 | n155;
assign n28 = n279 | n298;
assign n14 = ~(n124 ^ n126);
assign n66 = ~(n30 ^ n29);
assign n143 = n140 | n216;
assign n38 = n301 | n72;
assign n262 = ~(n238 ^ n29);
assign n259 = ~n180;
assign n251 = n96 | n51;
assign n45 = ~(n43 ^ n214);
assign n60 = ~(n8 ^ n114);
assign n19 = n273 | n297;
assign n34 = ~(n70 ^ n174);
assign n209 = n140 | n175;
assign n275 = n53 | n276;
assign n239 = ~(n14 ^ n288);
assign n308 = ~(n70 ^ n2);
assign n255 = n251 | n172;
assign n166 = n305 | n181;
assign n198 = n252 | n173;
assign n86 = ~(n200 ^ n196);
assign n223 = n250 | n46;
assign n5 = n62 | n85;
assign n161 = n178 | n64;
assign n204 = ~n58;
assign n1 = ~(n189 ^ n296);
assign n301 = ~n119;
assign n9 = n283 | n291;
assign n304 = ~(n224 ^ n214);
assign n208 = ~(n225 ^ n83);
assign n21 = n110 | n82;
assign n57 = ~(n135 ^ n197);
assign n296 = ~(n179 ^ n0);
assign n203 = n171 | n103;
assign n243 = n205 | n155;
assign n303 = ~(n237 ^ n210);
assign n191 = ~(n278 ^ n272);
assign n171 = ~n226;
assign n233 = n149 ^ n309;
assign n140 = ~n78;
assign n279 = ~n119;
assign n63 = ~(n130 ^ n107);
assign n220 = n235 | n274;
assign n65 = n128 | n68;
assign n103 = ~n281;
assign n150 = n60;
assign n149 = ~(n32 ^ n141);
assign n270 = n112 | n190;
assign n41 = n155 | n230;
assign n248 = ~(n17 ^ n75);
assign n267 = n56 | n273;
assign n294 = n204 | n103;
assign n85 = n152 | n276;
assign n62 = n140 | n216;
assign n274 = n95 | n76;
assign n311 = ~(n130 ^ n256);
assign n114 = ~(n294 ^ n87);
assign n222 = ~(n77 ^ n191);
assign n69 = n156 | n76;
assign n263 = n162 | n51;
assign n221 = ~(n219 ^ n179);
assign n36 = n258 | n33;
assign n254 = ~(n23 ^ n249);
assign n306 = ~(n290 ^ n10);
assign n297 = ~n279;
assign n286 = ~(n49 ^ n238);
assign n141 = ~(n256 ^ n289);
assign n67 = n167 | n159;
assign n104 = ~(n142 ^ n289);
assign n26 = ~(n115 ^ n169);
assign n92 = n127 | n113;
assign n244 = n243 | n232;
assign n269 = n56 | n72;
assign n142 = n209 | n9;
assign n10 = ~(n234 ^ n196);
assign n215 = n15 | n33;
assign n216 = ~n134;
assign n154 = n263 | n198;
assign n113 = n183 | n230;
assign n186 = n184 | n103;
assign n68 = n206 | n255;
assign n93 = ~n74;
assign n52 = ~(n238 ^ n17);
assign n49 = n28 | n159;
assign n188 = n162 | n106;
assign n250 = n301 | n298;
assign n115 = n105 | n64;
assign n240 = ~(n229 ^ n303);
assign n33 = n267 | n173;
assign n197 = ~(n285 ^ n42);
assign n87 = ~(n278 ^ n234);
assign n88 = ~(n299 ^ n107);
assign n117 = ~(n194 ^ n27);
assign n227 = ~(n242 ^ n240);
assign n89 = ~(n271 ^ n43);
assign n290 = ~(n260 ^ n27);
assign n202 = n101 | n9;
assign n280 = n177 | n297;
assign n155 = ~n60;
assign n46 = n7 | n181;
assign n258 = n301 | n138;
assign n126 = ~(n249 ^ n214);
assign n190 = ~n100;
assign n158 = n112 | n190;
assign n177 = ~n233;
assign n30 = n13 | n274;
assign n175 = ~n134;
assign n232 = n301 | n25;
assign n252 = n96 | n93;
assign n156 = n96 | n93;
assign n160 = ~(n16 ^ n70);
assign n167 = n177 | n51;
assign n159 = n266 | n92;
assign n152 = n150 | n230;
assign n172 = n298 | n93;
assign n287 = ~(n83 ^ n222);
assign n101 = n112 | n231;
assign n235 = n177 | n259;
assign n94 = ~(n223 ^ n137);
assign n310 = ~(n65 ^ n237);
assign n25 = n138 | n106;
assign n299 = n144 | n244;
assign n31 = n38 | n69;
assign n81 = ~(n132 ^ n90);
assign n39 = n301 | n298;
assign n72 = ~n50;
assign n134 = ~n71;
assign n246 = ~(n277 ^ n249);
assign n245 = ~(n136 ^ n108);
assign n11 = n39 | n201;
assign n183 = ~n110;
assign n298 = ~n50;
assign n162 = ~n233;
assign n213 = ~(n220 ^ n75);
assign n305 = n56 | n273;
assign n82 = ~n241;
assign n164 = ~(n161 ^ n2);
assign n131 = ~(n102 ^ n120);
assign n122 = ~(n208 ^ n45);
assign n132 = n158 | n85;
assign n293 = n157 | n103;
assign n95 = n56 | n273;
assign n205 = n57;
assign n257 = ~n91;
assign n148 = n112 | n41;
assign n120 = ~(n187 ^ n211);
assign n283 = n205 | n155;
assign n99 = n307 | n147;
assign n284 = n55 | n46;
assign n6 = ~(n306 ^ n222);
assign n73 = ~(n284 ^ n260);
assign n178 = n112 | n231;
assign n78 = n131 ^ n44;
assign n173 = n140 | n3;
assign n125 = ~(n287 ^ n63);
assign n136 = ~(n163 ^ n195);
assign n195 = ~(n210 ^ n59);
assign n105 = n110 | n175;
assign n7 = n96 | n93;
assign n199 = ~(n36 ^ n187);
assign n277 = n21 | n147;
assign n118 = ~(n293 ^ n34);
assign n145 = ~(n11 ^ n278);
assign n218 = ~(n97 ^ n268);
assign n291 = n297 | n188;
assign n32 = ~(n225 ^ n306);
assign n121 = ~(n137 ^ n260);
assign n48 = n279 | n138;
assign n153 = n143 | n68;
assign n80 = ~(n116 ^ n174);
assign n229 = n257 | n103;
assign n61 = ~(n67 ^ n17);
assign n54 = ~(n2 ^ n169);
assign n200 = n236 | n69;
assign n96 = n227;
assign n193 = n150 | n230;
assign n176 = n280 | n166;
assign n185 = n162 | n297;
assign n128 = n112 | n183;
assign n100 = ~n78;
assign n24 = ~(n5 ^ n59);
assign n77 = ~(n137 ^ n194);
assign n207 = ~(n29 ^ n75);
assign n276 = n269 | n19;
assign n139 = n96 | n93;
assign n212 = ~(n99 ^ n23);
assign n217 = ~(n202 ^ n256);
assign n302 = n185 | n201;
assign n146 = ~(n179 ^ n187);
assign n268 = ~(n90 ^ n59);
assign n206 = n150 | n230;
assign n230 = ~n57;
assign n12 = n241 | n183;
assign n3 = n82 | n41;
assign n109 = n47 | n232;
assign n236 = n162 | n259;
assign n135 = ~(n239 ^ n207);
assign n47 = n150 | n230;
assign n64 = n193 | n291;
assign n4 = n35 | n198;
assign n56 = n74;
assign n264 = n12 | n244;
assign n74 = ~(n122 ^ n218);
assign n168 = ~(n264 ^ n130);
assign n112 = ~n71;
assign n189 = ~(n288 ^ n108);
assign n102 = ~(n14 ^ n136);
assign n8 = ~(n245 ^ n52);
assign n71 = n1 ^ n182;
assign n300 = n155 | n82;
assign n242 = ~(n6 ^ n254);
assign n79 = ~n84;
assign n123 = ~(n215 ^ n211);
assign n151 = ~(n302 ^ n234);
assign n127 = n150 | n175;
assign n266 = n56 | n273;
assign n50 = ~n233;
assign n295 = ~(n23 ^ n43);
assign n22 = n247 | n103;
assign n16 = n270 | n109;
assign n42 = ~(n272 ^ n196);
assign n116 = n20 | n109;
assign n147 = n165 | n255;
assign n181 = n183 | n148;
assign n170 = n241 | n231;
assign n165 = n205 | n155;
assign n225 = ~(n111 ^ n248);
assign n241 = ~n71;
assign n265 = ~(n4 ^ n194);
assign n35 = n301 | n138;
assign n157 = ~n37;
assign n192 = ~n292;
assign n285 = n79 | n103;
assign n184 = ~n18;
assign n55 = n162 | n259;
assign n309 = ~(n186 ^ n54);
assign n119 = n125 ^ n118;
assign n97 = n192 | n103;
assign n13 = n279 | n72;
assign n106 = n273 | n93;
assign n273 = ~n227;
assign n307 = n241 | n190;
assign n231 = ~n100;
assign n51 = ~n180;
assign n76 = n282 | n300;
assign n224 = n228 | n275;
assign n247 = ~n133;
assign n83 = ~(n146 ^ n262);
assign n201 = n139 | n92;
assign n228 = n140 | n82;
assign n182 = ~(n203 ^ n121);
assign n124 = ~(n107 ^ n289);
assign n15 = n162 | n51;
assign n219 = n48 | n166;
assign n253 = ~(n31 ^ n272);
assign n180 = ~n119;
assign n138 = ~n177;
assign n108 = ~(n308 ^ n40);
assign n110 = ~n78;
assign n271 = n170 | n275;
assign n20 = n140 | n175;
assign n98 = ~(n154 ^ n27);
assign n44 = ~(n22 ^ n117);
assign n111 = ~(n0 ^ n211);
assign n282 = n205 | n231;
assign n288 = ~(n311 ^ n295);
assign n40 = ~(n237 ^ n90);
assign n261 = ~(n176 ^ n0);
assign n144 = n110 | n216;
endmodule
