// Benchmark "top" written by ABC on Mon Jun 12 20:58:00 2023

module top ( 
    \1_n1 , \1_n105 , \1_n114 , \1_n117 , \1_n122 , \1_n15 , \1_n152 ,
    \1_n155 , \1_n160 , \1_n162 , \1_n168 , \1_n183 , \1_n187 , \1_n194 ,
    \1_n198 , \1_n206 , \1_n21 , \1_n215 , \1_n218 , \1_n227 , \1_n228 ,
    \1_n23 , \1_n231 , \1_n242 , \1_n269 , \1_n276 , \1_n278 , \1_n28 ,
    \1_n280 , \1_n37 , \1_n38 , \1_n4 , \1_n45 , \1_n52 , \1_n53 , \1_n60 ,
    \1_n75 , \1_n79 , \1_n83 , \1_n87 , \1_n95 , \2_n0 , \2_n107 ,
    \2_n130 , \2_n133 , \2_n137 , \2_n169 , \2_n17 , \2_n174 , \2_n179 ,
    \2_n18 , \2_n187 , \2_n194 , \2_n196 , \2_n2 , \2_n210 , \2_n211 ,
    \2_n214 , \2_n226 , \2_n23 , \2_n234 , \2_n237 , \2_n238 , \2_n249 ,
    \2_n256 , \2_n260 , \2_n27 , \2_n272 , \2_n278 , \2_n281 , \2_n289 ,
    \2_n29 , \2_n292 , \2_n37 , \2_n43 , \2_n58 , \2_n59 , \2_n70 ,
    \2_n75 , \2_n84 , \2_n90 , \2_n91 ,
    \1_n111 , \1_n139 , \1_n154 , \1_n176 , \1_n185 , \1_n191 , \1_n197 ,
    \1_n200 , \1_n205 , \1_n208 , \1_n211 , \1_n214 , \1_n220 , \1_n243 ,
    \1_n248 , \1_n254 , \1_n262 , \1_n265 , \1_n273 , \1_n283 , \1_n3 ,
    \1_n32 , \1_n40 , \1_n47 , \1_n50 , \1_n54 , \1_n72 , \1_n81 , \1_n86 ,
    \1_n91 , \1_n97 , \1_n99 , \2_n104 , \2_n123 , \2_n129 , \2_n145 ,
    \2_n151 , \2_n160 , \2_n164 , \2_n168 , \2_n199 , \2_n212 , \2_n213 ,
    \2_n217 , \2_n221 , \2_n24 , \2_n246 , \2_n253 , \2_n26 , \2_n261 ,
    \2_n265 , \2_n286 , \2_n304 , \2_n310 , \2_n61 , \2_n66 , \2_n73 ,
    \2_n80 , \2_n81 , \2_n86 , \2_n88 , \2_n89 , \2_n94 , \2_n98   );
  input  \1_n1 , \1_n105 , \1_n114 , \1_n117 , \1_n122 , \1_n15 ,
    \1_n152 , \1_n155 , \1_n160 , \1_n162 , \1_n168 , \1_n183 , \1_n187 ,
    \1_n194 , \1_n198 , \1_n206 , \1_n21 , \1_n215 , \1_n218 , \1_n227 ,
    \1_n228 , \1_n23 , \1_n231 , \1_n242 , \1_n269 , \1_n276 , \1_n278 ,
    \1_n28 , \1_n280 , \1_n37 , \1_n38 , \1_n4 , \1_n45 , \1_n52 , \1_n53 ,
    \1_n60 , \1_n75 , \1_n79 , \1_n83 , \1_n87 , \1_n95 , \2_n0 , \2_n107 ,
    \2_n130 , \2_n133 , \2_n137 , \2_n169 , \2_n17 , \2_n174 , \2_n179 ,
    \2_n18 , \2_n187 , \2_n194 , \2_n196 , \2_n2 , \2_n210 , \2_n211 ,
    \2_n214 , \2_n226 , \2_n23 , \2_n234 , \2_n237 , \2_n238 , \2_n249 ,
    \2_n256 , \2_n260 , \2_n27 , \2_n272 , \2_n278 , \2_n281 , \2_n289 ,
    \2_n29 , \2_n292 , \2_n37 , \2_n43 , \2_n58 , \2_n59 , \2_n70 ,
    \2_n75 , \2_n84 , \2_n90 , \2_n91 ;
  output \1_n111 , \1_n139 , \1_n154 , \1_n176 , \1_n185 , \1_n191 , \1_n197 ,
    \1_n200 , \1_n205 , \1_n208 , \1_n211 , \1_n214 , \1_n220 , \1_n243 ,
    \1_n248 , \1_n254 , \1_n262 , \1_n265 , \1_n273 , \1_n283 , \1_n3 ,
    \1_n32 , \1_n40 , \1_n47 , \1_n50 , \1_n54 , \1_n72 , \1_n81 , \1_n86 ,
    \1_n91 , \1_n97 , \1_n99 , \2_n104 , \2_n123 , \2_n129 , \2_n145 ,
    \2_n151 , \2_n160 , \2_n164 , \2_n168 , \2_n199 , \2_n212 , \2_n213 ,
    \2_n217 , \2_n221 , \2_n24 , \2_n246 , \2_n253 , \2_n26 , \2_n261 ,
    \2_n265 , \2_n286 , \2_n304 , \2_n310 , \2_n61 , \2_n66 , \2_n73 ,
    \2_n80 , \2_n81 , \2_n86 , \2_n88 , \2_n89 , \2_n94 , \2_n98 ;
  wire new_n147_, new_n148_, new_n149_, new_n150_, new_n151_, new_n152_,
    new_n153_, new_n154_, new_n155_, new_n156_, new_n157_, new_n158_,
    new_n159_, new_n160_, new_n161_, new_n162_, new_n163_, new_n164_,
    new_n165_, new_n166_, new_n167_, new_n168_, new_n169_, new_n170_,
    new_n171_, new_n172_, new_n173_, new_n174_, new_n175_, new_n176_,
    new_n177_, new_n178_, new_n179_, new_n180_, new_n181_, new_n182_,
    new_n183_, new_n184_, new_n185_, new_n186_, new_n187_, new_n188_,
    new_n189_, new_n190_, new_n191_, new_n192_, new_n193_, new_n194_,
    new_n195_, new_n196_, new_n197_, new_n198_, new_n199_, new_n200_,
    new_n201_, new_n202_, new_n203_, new_n204_, new_n205_, new_n206_,
    new_n207_, new_n208_, new_n209_, new_n210_, new_n211_, new_n212_,
    new_n213_, new_n214_, new_n215_, new_n216_, new_n217_, new_n218_,
    new_n219_, new_n220_, new_n221_, new_n222_, new_n223_, new_n224_,
    new_n225_, new_n226_, new_n227_, new_n228_, new_n229_, new_n230_,
    new_n231_, new_n232_, new_n233_, new_n234_, new_n235_, new_n236_,
    new_n237_, new_n238_, new_n239_, new_n240_, new_n241_, new_n242_,
    new_n243_, new_n244_, new_n245_, new_n246_, new_n247_, new_n248_,
    new_n249_, new_n250_, new_n251_, new_n252_, new_n253_, new_n254_,
    new_n255_, new_n256_, new_n257_, new_n258_, new_n259_, new_n260_,
    new_n261_, new_n262_, new_n263_, new_n264_, new_n265_, new_n266_,
    new_n267_, new_n268_, new_n269_, new_n270_, new_n271_, new_n272_,
    new_n273_, new_n274_, new_n275_, new_n276_, new_n277_, new_n278_,
    new_n279_, new_n280_, new_n281_, new_n282_, new_n283_, new_n284_,
    new_n285_, new_n286_, new_n287_, new_n288_, new_n289_, new_n290_,
    new_n291_, new_n292_, new_n293_, new_n294_, new_n295_, new_n296_,
    new_n297_, new_n298_, new_n299_, new_n300_, new_n301_, new_n302_,
    new_n303_, new_n304_, new_n305_, new_n306_, new_n307_, new_n308_,
    new_n309_, new_n310_, new_n311_, new_n312_, new_n313_, new_n314_,
    new_n315_, new_n316_, new_n317_, new_n318_, new_n319_, new_n320_,
    new_n321_, new_n322_, new_n323_, new_n324_, new_n325_, new_n326_,
    new_n327_, new_n328_, new_n329_, new_n330_, new_n331_, new_n332_,
    new_n333_, new_n334_, new_n335_, new_n336_, new_n337_, new_n338_,
    new_n339_, new_n340_, new_n341_, new_n342_, new_n343_, new_n344_,
    new_n345_, new_n346_, new_n347_, new_n348_, new_n349_, new_n350_,
    new_n351_, new_n352_, new_n353_, new_n354_, new_n355_, new_n356_,
    new_n357_, new_n358_, new_n359_, new_n360_, new_n361_, new_n362_,
    new_n363_, new_n364_, new_n365_, new_n366_, new_n367_, new_n368_,
    new_n369_, new_n370_, new_n371_, new_n372_, new_n373_, new_n374_,
    new_n375_, new_n376_, new_n377_, new_n378_, new_n379_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n388_,
    new_n389_, new_n390_, new_n391_, new_n392_, new_n393_, new_n394_,
    new_n395_, new_n397_, new_n398_, new_n399_, new_n400_, new_n401_,
    new_n403_, new_n404_, new_n405_, new_n406_, new_n407_, new_n409_,
    new_n410_, new_n411_, new_n412_, new_n413_, new_n414_, new_n416_,
    new_n417_, new_n418_, new_n419_, new_n420_, new_n421_, new_n422_,
    new_n423_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n432_, new_n433_, new_n434_, new_n436_, new_n437_,
    new_n438_, new_n439_, new_n441_, new_n442_, new_n443_, new_n444_,
    new_n445_, new_n447_, new_n448_, new_n449_, new_n451_, new_n452_,
    new_n453_, new_n454_, new_n455_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n462_, new_n463_, new_n464_, new_n466_, new_n467_,
    new_n468_, new_n469_, new_n471_, new_n472_, new_n473_, new_n475_,
    new_n476_, new_n477_, new_n478_, new_n480_, new_n481_, new_n482_,
    new_n483_, new_n485_, new_n486_, new_n487_, new_n488_, new_n490_,
    new_n491_, new_n492_, new_n493_, new_n495_, new_n496_, new_n497_,
    new_n499_, new_n500_, new_n501_, new_n503_, new_n504_, new_n505_,
    new_n507_, new_n508_, new_n509_, new_n510_, new_n512_, new_n513_,
    new_n514_, new_n516_, new_n517_, new_n518_, new_n520_, new_n521_,
    new_n522_, new_n524_, new_n525_, new_n526_, new_n528_, new_n529_,
    new_n530_, new_n532_, new_n533_, new_n534_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n541_, new_n542_, new_n543_, new_n544_,
    new_n545_, new_n546_, new_n547_, new_n548_, new_n549_, new_n550_,
    new_n551_, new_n552_, new_n553_, new_n554_, new_n555_, new_n556_,
    new_n557_, new_n558_, new_n559_, new_n560_, new_n561_, new_n562_,
    new_n563_, new_n564_, new_n565_, new_n566_, new_n567_, new_n568_,
    new_n569_, new_n570_, new_n571_, new_n572_, new_n573_, new_n574_,
    new_n575_, new_n576_, new_n577_, new_n578_, new_n579_, new_n580_,
    new_n581_, new_n582_, new_n583_, new_n584_, new_n585_, new_n586_,
    new_n587_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n706_,
    new_n707_, new_n708_, new_n709_, new_n710_, new_n711_, new_n712_,
    new_n713_, new_n714_, new_n715_, new_n716_, new_n717_, new_n718_,
    new_n719_, new_n720_, new_n721_, new_n722_, new_n723_, new_n724_,
    new_n725_, new_n726_, new_n727_, new_n728_, new_n729_, new_n730_,
    new_n731_, new_n732_, new_n733_, new_n734_, new_n735_, new_n736_,
    new_n737_, new_n738_, new_n739_, new_n740_, new_n741_, new_n742_,
    new_n743_, new_n744_, new_n745_, new_n746_, new_n747_, new_n748_,
    new_n749_, new_n750_, new_n751_, new_n752_, new_n753_, new_n754_,
    new_n755_, new_n756_, new_n757_, new_n758_, new_n759_, new_n760_,
    new_n761_, new_n762_, new_n763_, new_n764_, new_n765_, new_n766_,
    new_n767_, new_n768_, new_n769_, new_n770_, new_n771_, new_n772_,
    new_n773_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n804_, new_n805_, new_n806_,
    new_n808_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_,
    new_n814_, new_n816_, new_n817_, new_n818_, new_n819_, new_n821_,
    new_n822_, new_n823_, new_n824_, new_n826_, new_n827_, new_n828_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n843_,
    new_n844_, new_n845_, new_n847_, new_n848_, new_n849_, new_n850_,
    new_n851_, new_n852_, new_n854_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n859_, new_n860_, new_n862_, new_n863_, new_n864_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n871_, new_n872_,
    new_n873_, new_n875_, new_n876_, new_n877_, new_n879_, new_n880_,
    new_n881_, new_n882_, new_n884_, new_n885_, new_n886_, new_n887_,
    new_n889_, new_n890_, new_n891_, new_n892_, new_n894_, new_n895_,
    new_n896_, new_n898_, new_n899_, new_n900_, new_n902_, new_n903_,
    new_n904_, new_n906_, new_n907_, new_n908_, new_n909_, new_n911_,
    new_n912_, new_n913_, new_n915_, new_n916_, new_n917_, new_n919_,
    new_n920_, new_n921_, new_n923_, new_n924_, new_n925_, new_n927_,
    new_n928_, new_n929_, new_n931_, new_n932_, new_n933_, new_n935_,
    new_n936_, new_n937_;
  assign new_n147_ = \1_n87  & ~\1_n242 ;
  assign new_n148_ = ~\1_n87  & \1_n242 ;
  assign new_n149_ = ~new_n147_ & ~new_n148_;
  assign new_n150_ = \1_n52  & ~\1_n278 ;
  assign new_n151_ = ~\1_n52  & \1_n278 ;
  assign new_n152_ = ~new_n150_ & ~new_n151_;
  assign new_n153_ = ~new_n149_ & new_n152_;
  assign new_n154_ = new_n149_ & ~new_n152_;
  assign new_n155_ = ~new_n153_ & ~new_n154_;
  assign new_n156_ = \1_n45  & ~\1_n187 ;
  assign new_n157_ = ~\1_n45  & \1_n187 ;
  assign new_n158_ = ~new_n156_ & ~new_n157_;
  assign new_n159_ = ~new_n155_ & new_n158_;
  assign new_n160_ = new_n155_ & ~new_n158_;
  assign new_n161_ = ~new_n159_ & ~new_n160_;
  assign new_n162_ = \1_n95  & ~\1_n228 ;
  assign new_n163_ = ~\1_n95  & \1_n228 ;
  assign new_n164_ = ~new_n162_ & ~new_n163_;
  assign new_n165_ = ~\1_n53  & \1_n155 ;
  assign new_n166_ = \1_n53  & ~\1_n155 ;
  assign new_n167_ = ~new_n165_ & ~new_n166_;
  assign new_n168_ = ~\1_n23  & \1_n83 ;
  assign new_n169_ = \1_n23  & ~\1_n83 ;
  assign new_n170_ = ~new_n168_ & ~new_n169_;
  assign new_n171_ = ~new_n167_ & new_n170_;
  assign new_n172_ = new_n167_ & ~new_n170_;
  assign new_n173_ = ~new_n171_ & ~new_n172_;
  assign new_n174_ = \1_n4  & \1_n114 ;
  assign new_n175_ = ~new_n173_ & ~new_n174_;
  assign new_n176_ = new_n173_ & new_n174_;
  assign new_n177_ = ~new_n175_ & ~new_n176_;
  assign new_n178_ = ~new_n164_ & new_n177_;
  assign new_n179_ = new_n164_ & ~new_n177_;
  assign new_n180_ = ~new_n178_ & ~new_n179_;
  assign new_n181_ = ~new_n161_ & new_n180_;
  assign new_n182_ = new_n161_ & ~new_n180_;
  assign new_n183_ = ~new_n181_ & ~new_n182_;
  assign new_n184_ = \1_n37  & ~\1_n194 ;
  assign new_n185_ = ~\1_n37  & \1_n194 ;
  assign new_n186_ = ~new_n184_ & ~new_n185_;
  assign new_n187_ = \1_n21  & ~\1_n280 ;
  assign new_n188_ = ~\1_n21  & \1_n280 ;
  assign new_n189_ = ~new_n187_ & ~new_n188_;
  assign new_n190_ = ~new_n186_ & new_n189_;
  assign new_n191_ = new_n186_ & ~new_n189_;
  assign new_n192_ = ~new_n190_ & ~new_n191_;
  assign new_n193_ = \1_n75  & ~\1_n122 ;
  assign new_n194_ = ~\1_n75  & \1_n122 ;
  assign new_n195_ = ~new_n193_ & ~new_n194_;
  assign new_n196_ = ~new_n192_ & new_n195_;
  assign new_n197_ = new_n192_ & ~new_n195_;
  assign new_n198_ = ~new_n196_ & ~new_n197_;
  assign new_n199_ = ~\1_n79  & \1_n276 ;
  assign new_n200_ = \1_n79  & ~\1_n276 ;
  assign new_n201_ = ~new_n199_ & ~new_n200_;
  assign new_n202_ = ~\1_n105  & \1_n160 ;
  assign new_n203_ = \1_n105  & ~\1_n160 ;
  assign new_n204_ = ~new_n202_ & ~new_n203_;
  assign new_n205_ = ~\1_n152  & \1_n227 ;
  assign new_n206_ = \1_n152  & ~\1_n227 ;
  assign new_n207_ = ~new_n205_ & ~new_n206_;
  assign new_n208_ = ~new_n204_ & new_n207_;
  assign new_n209_ = new_n204_ & ~new_n207_;
  assign new_n210_ = ~new_n208_ & ~new_n209_;
  assign new_n211_ = \1_n4  & \1_n60 ;
  assign new_n212_ = ~new_n210_ & ~new_n211_;
  assign new_n213_ = new_n210_ & new_n211_;
  assign new_n214_ = ~new_n212_ & ~new_n213_;
  assign new_n215_ = ~new_n201_ & new_n214_;
  assign new_n216_ = new_n201_ & ~new_n214_;
  assign new_n217_ = ~new_n215_ & ~new_n216_;
  assign new_n218_ = ~new_n198_ & new_n217_;
  assign new_n219_ = new_n198_ & ~new_n217_;
  assign new_n220_ = ~new_n218_ & ~new_n219_;
  assign new_n221_ = \1_n162  & ~\1_n215 ;
  assign new_n222_ = ~\1_n162  & \1_n215 ;
  assign new_n223_ = ~new_n221_ & ~new_n222_;
  assign new_n224_ = ~new_n173_ & new_n223_;
  assign new_n225_ = new_n173_ & ~new_n223_;
  assign new_n226_ = ~new_n224_ & ~new_n225_;
  assign new_n227_ = \1_n15  & ~\1_n28 ;
  assign new_n228_ = ~\1_n15  & \1_n28 ;
  assign new_n229_ = ~new_n227_ & ~new_n228_;
  assign new_n230_ = \1_n4  & \1_n198 ;
  assign new_n231_ = ~new_n210_ & ~new_n230_;
  assign new_n232_ = new_n210_ & new_n230_;
  assign new_n233_ = ~new_n231_ & ~new_n232_;
  assign new_n234_ = ~new_n229_ & new_n233_;
  assign new_n235_ = new_n229_ & ~new_n233_;
  assign new_n236_ = ~new_n234_ & ~new_n235_;
  assign new_n237_ = ~new_n226_ & new_n236_;
  assign new_n238_ = new_n226_ & ~new_n236_;
  assign new_n239_ = ~new_n237_ & ~new_n238_;
  assign new_n240_ = new_n220_ & new_n239_;
  assign new_n241_ = ~new_n183_ & new_n240_;
  assign new_n242_ = ~\1_n122  & \1_n187 ;
  assign new_n243_ = \1_n122  & ~\1_n187 ;
  assign new_n244_ = ~new_n242_ & ~new_n243_;
  assign new_n245_ = \1_n206  & ~\1_n215 ;
  assign new_n246_ = ~\1_n206  & \1_n215 ;
  assign new_n247_ = ~new_n245_ & ~new_n246_;
  assign new_n248_ = ~new_n244_ & new_n247_;
  assign new_n249_ = new_n244_ & ~new_n247_;
  assign new_n250_ = ~new_n248_ & ~new_n249_;
  assign new_n251_ = ~\1_n105  & \1_n194 ;
  assign new_n252_ = \1_n105  & ~\1_n194 ;
  assign new_n253_ = ~new_n251_ & ~new_n252_;
  assign new_n254_ = ~new_n250_ & new_n253_;
  assign new_n255_ = new_n250_ & ~new_n253_;
  assign new_n256_ = ~new_n254_ & ~new_n255_;
  assign new_n257_ = ~\1_n53  & \1_n242 ;
  assign new_n258_ = \1_n53  & ~\1_n242 ;
  assign new_n259_ = ~new_n257_ & ~new_n258_;
  assign new_n260_ = \1_n45  & ~\1_n75 ;
  assign new_n261_ = ~\1_n45  & \1_n75 ;
  assign new_n262_ = ~new_n260_ & ~new_n261_;
  assign new_n263_ = ~\1_n162  & \1_n183 ;
  assign new_n264_ = \1_n162  & ~\1_n183 ;
  assign new_n265_ = ~new_n263_ & ~new_n264_;
  assign new_n266_ = ~new_n262_ & new_n265_;
  assign new_n267_ = new_n262_ & ~new_n265_;
  assign new_n268_ = ~new_n266_ & ~new_n267_;
  assign new_n269_ = \1_n4  & \1_n117 ;
  assign new_n270_ = ~new_n268_ & ~new_n269_;
  assign new_n271_ = new_n268_ & new_n269_;
  assign new_n272_ = ~new_n270_ & ~new_n271_;
  assign new_n273_ = ~new_n259_ & new_n272_;
  assign new_n274_ = new_n259_ & ~new_n272_;
  assign new_n275_ = ~new_n273_ & ~new_n274_;
  assign new_n276_ = ~new_n256_ & new_n275_;
  assign new_n277_ = new_n256_ & ~new_n275_;
  assign new_n278_ = ~new_n276_ & ~new_n277_;
  assign new_n279_ = \1_n183  & ~\1_n206 ;
  assign new_n280_ = ~\1_n183  & \1_n206 ;
  assign new_n281_ = ~new_n279_ & ~new_n280_;
  assign new_n282_ = ~new_n155_ & new_n281_;
  assign new_n283_ = new_n155_ & ~new_n281_;
  assign new_n284_ = ~new_n282_ & ~new_n283_;
  assign new_n285_ = ~\1_n1  & \1_n38 ;
  assign new_n286_ = \1_n1  & ~\1_n38 ;
  assign new_n287_ = ~new_n285_ & ~new_n286_;
  assign new_n288_ = \1_n4  & \1_n269 ;
  assign new_n289_ = ~new_n192_ & ~new_n288_;
  assign new_n290_ = new_n192_ & new_n288_;
  assign new_n291_ = ~new_n289_ & ~new_n290_;
  assign new_n292_ = ~new_n287_ & new_n291_;
  assign new_n293_ = new_n287_ & ~new_n291_;
  assign new_n294_ = ~new_n292_ & ~new_n293_;
  assign new_n295_ = ~new_n284_ & new_n294_;
  assign new_n296_ = new_n284_ & ~new_n294_;
  assign new_n297_ = ~new_n295_ & ~new_n296_;
  assign new_n298_ = new_n278_ & ~new_n297_;
  assign new_n299_ = ~\1_n79  & \1_n228 ;
  assign new_n300_ = \1_n79  & ~\1_n228 ;
  assign new_n301_ = ~new_n299_ & ~new_n300_;
  assign new_n302_ = \1_n1  & ~\1_n28 ;
  assign new_n303_ = ~\1_n1  & \1_n28 ;
  assign new_n304_ = ~new_n302_ & ~new_n303_;
  assign new_n305_ = ~new_n301_ & new_n304_;
  assign new_n306_ = new_n301_ & ~new_n304_;
  assign new_n307_ = ~new_n305_ & ~new_n306_;
  assign new_n308_ = \1_n37  & ~\1_n160 ;
  assign new_n309_ = ~\1_n37  & \1_n160 ;
  assign new_n310_ = ~new_n308_ & ~new_n309_;
  assign new_n311_ = ~new_n307_ & new_n310_;
  assign new_n312_ = new_n307_ & ~new_n310_;
  assign new_n313_ = ~new_n311_ & ~new_n312_;
  assign new_n314_ = \1_n87  & ~\1_n155 ;
  assign new_n315_ = ~\1_n87  & \1_n155 ;
  assign new_n316_ = ~new_n314_ & ~new_n315_;
  assign new_n317_ = \1_n95  & ~\1_n276 ;
  assign new_n318_ = ~\1_n95  & \1_n276 ;
  assign new_n319_ = ~new_n317_ & ~new_n318_;
  assign new_n320_ = ~\1_n15  & \1_n38 ;
  assign new_n321_ = \1_n15  & ~\1_n38 ;
  assign new_n322_ = ~new_n320_ & ~new_n321_;
  assign new_n323_ = ~new_n319_ & new_n322_;
  assign new_n324_ = new_n319_ & ~new_n322_;
  assign new_n325_ = ~new_n323_ & ~new_n324_;
  assign new_n326_ = \1_n4  & \1_n168 ;
  assign new_n327_ = ~new_n325_ & ~new_n326_;
  assign new_n328_ = new_n325_ & new_n326_;
  assign new_n329_ = ~new_n327_ & ~new_n328_;
  assign new_n330_ = ~new_n316_ & new_n329_;
  assign new_n331_ = new_n316_ & ~new_n329_;
  assign new_n332_ = ~new_n330_ & ~new_n331_;
  assign new_n333_ = ~new_n313_ & new_n332_;
  assign new_n334_ = new_n313_ & ~new_n332_;
  assign new_n335_ = ~new_n333_ & ~new_n334_;
  assign new_n336_ = \1_n21  & ~\1_n227 ;
  assign new_n337_ = ~\1_n21  & \1_n227 ;
  assign new_n338_ = ~new_n336_ & ~new_n337_;
  assign new_n339_ = ~new_n268_ & new_n338_;
  assign new_n340_ = new_n268_ & ~new_n338_;
  assign new_n341_ = ~new_n339_ & ~new_n340_;
  assign new_n342_ = \1_n52  & ~\1_n83 ;
  assign new_n343_ = ~\1_n52  & \1_n83 ;
  assign new_n344_ = ~new_n342_ & ~new_n343_;
  assign new_n345_ = \1_n4  & \1_n231 ;
  assign new_n346_ = ~new_n325_ & ~new_n345_;
  assign new_n347_ = new_n325_ & new_n345_;
  assign new_n348_ = ~new_n346_ & ~new_n347_;
  assign new_n349_ = ~new_n344_ & new_n348_;
  assign new_n350_ = new_n344_ & ~new_n348_;
  assign new_n351_ = ~new_n349_ & ~new_n350_;
  assign new_n352_ = ~new_n341_ & new_n351_;
  assign new_n353_ = new_n341_ & ~new_n351_;
  assign new_n354_ = ~new_n352_ & ~new_n353_;
  assign new_n355_ = ~\1_n152  & \1_n280 ;
  assign new_n356_ = \1_n152  & ~\1_n280 ;
  assign new_n357_ = ~new_n355_ & ~new_n356_;
  assign new_n358_ = ~new_n307_ & new_n357_;
  assign new_n359_ = new_n307_ & ~new_n357_;
  assign new_n360_ = ~new_n358_ & ~new_n359_;
  assign new_n361_ = ~\1_n23  & \1_n278 ;
  assign new_n362_ = \1_n23  & ~\1_n278 ;
  assign new_n363_ = ~new_n361_ & ~new_n362_;
  assign new_n364_ = \1_n4  & \1_n218 ;
  assign new_n365_ = ~new_n250_ & ~new_n364_;
  assign new_n366_ = new_n250_ & new_n364_;
  assign new_n367_ = ~new_n365_ & ~new_n366_;
  assign new_n368_ = ~new_n363_ & new_n367_;
  assign new_n369_ = new_n363_ & ~new_n367_;
  assign new_n370_ = ~new_n368_ & ~new_n369_;
  assign new_n371_ = ~new_n360_ & new_n370_;
  assign new_n372_ = new_n360_ & ~new_n370_;
  assign new_n373_ = ~new_n371_ & ~new_n372_;
  assign new_n374_ = new_n354_ & ~new_n373_;
  assign new_n375_ = new_n335_ & new_n374_;
  assign new_n376_ = new_n298_ & new_n375_;
  assign new_n377_ = new_n241_ & new_n376_;
  assign new_n378_ = \1_n278  & new_n377_;
  assign new_n379_ = ~\1_n278  & ~new_n377_;
  assign \1_n3  = ~new_n378_ & ~new_n379_;
  assign new_n381_ = new_n278_ & new_n297_;
  assign new_n382_ = ~new_n335_ & new_n381_;
  assign new_n383_ = new_n374_ & new_n382_;
  assign new_n384_ = new_n241_ & new_n383_;
  assign new_n385_ = \1_n228  & new_n384_;
  assign new_n386_ = ~\1_n228  & ~new_n384_;
  assign \1_n32  = ~new_n385_ & ~new_n386_;
  assign new_n388_ = ~new_n354_ & new_n373_;
  assign new_n389_ = new_n183_ & new_n240_;
  assign new_n390_ = ~new_n278_ & ~new_n297_;
  assign new_n391_ = new_n335_ & new_n390_;
  assign new_n392_ = new_n389_ & new_n391_;
  assign new_n393_ = new_n388_ & new_n392_;
  assign new_n394_ = \1_n183  & new_n393_;
  assign new_n395_ = ~\1_n183  & ~new_n393_;
  assign \1_n40  = ~new_n394_ & ~new_n395_;
  assign new_n397_ = new_n298_ & ~new_n335_;
  assign new_n398_ = new_n389_ & new_n397_;
  assign new_n399_ = new_n388_ & new_n398_;
  assign new_n400_ = \1_n38  & ~new_n399_;
  assign new_n401_ = ~\1_n38  & new_n399_;
  assign \1_n47  = new_n400_ | new_n401_;
  assign new_n403_ = new_n354_ & new_n373_;
  assign new_n404_ = new_n397_ & new_n403_;
  assign new_n405_ = new_n241_ & new_n404_;
  assign new_n406_ = \1_n87  & new_n405_;
  assign new_n407_ = ~\1_n87  & ~new_n405_;
  assign \1_n50  = ~new_n406_ & ~new_n407_;
  assign new_n409_ = ~new_n220_ & ~new_n239_;
  assign new_n410_ = new_n183_ & new_n409_;
  assign new_n411_ = new_n382_ & new_n410_;
  assign new_n412_ = new_n403_ & new_n411_;
  assign new_n413_ = \1_n160  & new_n412_;
  assign new_n414_ = ~\1_n160  & ~new_n412_;
  assign \1_n54  = ~new_n413_ & ~new_n414_;
  assign new_n416_ = new_n220_ & ~new_n239_;
  assign new_n417_ = new_n183_ & new_n416_;
  assign new_n418_ = ~new_n278_ & new_n297_;
  assign new_n419_ = new_n335_ & new_n418_;
  assign new_n420_ = new_n388_ & new_n419_;
  assign new_n421_ = new_n417_ & new_n420_;
  assign new_n422_ = \1_n162  & new_n421_;
  assign new_n423_ = ~\1_n162  & ~new_n421_;
  assign \1_n72  = ~new_n422_ & ~new_n423_;
  assign new_n425_ = ~new_n220_ & new_n239_;
  assign new_n426_ = new_n183_ & new_n425_;
  assign new_n427_ = new_n391_ & new_n426_;
  assign new_n428_ = new_n403_ & new_n427_;
  assign new_n429_ = \1_n194  & new_n428_;
  assign new_n430_ = ~\1_n194  & ~new_n428_;
  assign \1_n81  = ~new_n429_ & ~new_n430_;
  assign new_n432_ = new_n404_ & new_n426_;
  assign new_n433_ = \1_n37  & new_n432_;
  assign new_n434_ = ~\1_n37  & ~new_n432_;
  assign \1_n86  = ~new_n433_ & ~new_n434_;
  assign new_n436_ = new_n375_ & new_n410_;
  assign new_n437_ = new_n381_ & new_n436_;
  assign new_n438_ = \1_n152  & new_n437_;
  assign new_n439_ = ~\1_n152  & ~new_n437_;
  assign \1_n91  = ~new_n438_ & ~new_n439_;
  assign new_n441_ = ~new_n183_ & new_n416_;
  assign new_n442_ = new_n419_ & new_n441_;
  assign new_n443_ = new_n403_ & new_n442_;
  assign new_n444_ = \1_n53  & new_n443_;
  assign new_n445_ = ~\1_n53  & ~new_n443_;
  assign \1_n97  = ~new_n444_ & ~new_n445_;
  assign new_n447_ = new_n376_ & new_n426_;
  assign new_n448_ = \1_n280  & new_n447_;
  assign new_n449_ = ~\1_n280  & ~new_n447_;
  assign \1_n99  = ~new_n448_ & ~new_n449_;
  assign new_n451_ = new_n335_ & new_n388_;
  assign new_n452_ = new_n441_ & new_n451_;
  assign new_n453_ = new_n381_ & new_n452_;
  assign new_n454_ = \1_n83  & new_n453_;
  assign new_n455_ = ~\1_n83  & ~new_n453_;
  assign \1_n111  = ~new_n454_ & ~new_n455_;
  assign new_n457_ = new_n382_ & new_n441_;
  assign new_n458_ = new_n403_ & new_n457_;
  assign new_n459_ = \1_n155  & ~new_n458_;
  assign new_n460_ = ~\1_n155  & new_n458_;
  assign \1_n139  = new_n459_ | new_n460_;
  assign new_n462_ = new_n374_ & new_n392_;
  assign new_n463_ = \1_n206  & new_n462_;
  assign new_n464_ = ~\1_n206  & ~new_n462_;
  assign \1_n154  = ~new_n463_ & ~new_n464_;
  assign new_n466_ = new_n382_ & new_n388_;
  assign new_n467_ = new_n241_ & new_n466_;
  assign new_n468_ = \1_n95  & new_n467_;
  assign new_n469_ = ~\1_n95  & ~new_n467_;
  assign \1_n176  = ~new_n468_ & ~new_n469_;
  assign new_n471_ = new_n426_ & new_n466_;
  assign new_n472_ = \1_n276  & ~new_n471_;
  assign new_n473_ = ~\1_n276  & new_n471_;
  assign \1_n185  = new_n472_ | new_n473_;
  assign new_n475_ = new_n374_ & new_n419_;
  assign new_n476_ = new_n417_ & new_n475_;
  assign new_n477_ = \1_n215  & new_n476_;
  assign new_n478_ = ~\1_n215  & ~new_n476_;
  assign \1_n191  = ~new_n477_ & ~new_n478_;
  assign new_n480_ = new_n241_ & new_n391_;
  assign new_n481_ = new_n403_ & new_n480_;
  assign new_n482_ = \1_n242  & new_n481_;
  assign new_n483_ = ~\1_n242  & ~new_n481_;
  assign \1_n197  = ~new_n482_ & ~new_n483_;
  assign new_n485_ = new_n375_ & new_n441_;
  assign new_n486_ = new_n381_ & new_n485_;
  assign new_n487_ = \1_n23  & new_n486_;
  assign new_n488_ = ~\1_n23  & ~new_n486_;
  assign \1_n200  = ~new_n487_ & ~new_n488_;
  assign new_n490_ = new_n298_ & new_n451_;
  assign new_n491_ = new_n426_ & new_n490_;
  assign new_n492_ = \1_n21  & new_n491_;
  assign new_n493_ = ~\1_n21  & ~new_n491_;
  assign \1_n205  = ~new_n492_ & ~new_n493_;
  assign new_n495_ = new_n241_ & new_n490_;
  assign new_n496_ = \1_n52  & new_n495_;
  assign new_n497_ = ~\1_n52  & ~new_n495_;
  assign \1_n208  = ~new_n496_ & ~new_n497_;
  assign new_n499_ = new_n426_ & new_n475_;
  assign new_n500_ = \1_n122  & new_n499_;
  assign new_n501_ = ~\1_n122  & ~new_n499_;
  assign \1_n211  = ~new_n500_ & ~new_n501_;
  assign new_n503_ = new_n241_ & new_n475_;
  assign new_n504_ = \1_n187  & new_n503_;
  assign new_n505_ = ~\1_n187  & ~new_n503_;
  assign \1_n214  = ~new_n504_ & ~new_n505_;
  assign new_n507_ = new_n410_ & new_n451_;
  assign new_n508_ = new_n381_ & new_n507_;
  assign new_n509_ = \1_n227  & new_n508_;
  assign new_n510_ = ~\1_n227  & ~new_n508_;
  assign \1_n220  = ~new_n509_ & ~new_n510_;
  assign new_n512_ = new_n241_ & new_n420_;
  assign new_n513_ = \1_n45  & new_n512_;
  assign new_n514_ = ~\1_n45  & ~new_n512_;
  assign \1_n243  = ~new_n513_ & ~new_n514_;
  assign new_n516_ = new_n417_ & new_n466_;
  assign new_n517_ = \1_n15  & ~new_n516_;
  assign new_n518_ = ~\1_n15  & new_n516_;
  assign \1_n248  = new_n517_ | new_n518_;
  assign new_n520_ = new_n383_ & new_n417_;
  assign new_n521_ = \1_n28  & ~new_n520_;
  assign new_n522_ = ~\1_n28  & new_n520_;
  assign \1_n254  = new_n521_ | new_n522_;
  assign new_n524_ = new_n374_ & new_n398_;
  assign new_n525_ = \1_n1  & ~new_n524_;
  assign new_n526_ = ~\1_n1  & new_n524_;
  assign \1_n262  = new_n525_ | new_n526_;
  assign new_n528_ = new_n383_ & new_n426_;
  assign new_n529_ = \1_n79  & ~new_n528_;
  assign new_n530_ = ~\1_n79  & new_n528_;
  assign \1_n265  = new_n529_ | new_n530_;
  assign new_n532_ = new_n420_ & new_n426_;
  assign new_n533_ = \1_n75  & new_n532_;
  assign new_n534_ = ~\1_n75  & ~new_n532_;
  assign \1_n273  = ~new_n533_ & ~new_n534_;
  assign new_n536_ = new_n410_ & new_n419_;
  assign new_n537_ = new_n403_ & new_n536_;
  assign new_n538_ = \1_n105  & new_n537_;
  assign new_n539_ = ~\1_n105  & ~new_n537_;
  assign \1_n283  = ~new_n538_ & ~new_n539_;
  assign new_n541_ = ~\2_n107  & \2_n289 ;
  assign new_n542_ = \2_n107  & ~\2_n289 ;
  assign new_n543_ = ~new_n541_ & ~new_n542_;
  assign new_n544_ = \2_n214  & ~\2_n249 ;
  assign new_n545_ = ~\2_n214  & \2_n249 ;
  assign new_n546_ = ~new_n544_ & ~new_n545_;
  assign new_n547_ = ~new_n543_ & new_n546_;
  assign new_n548_ = new_n543_ & ~new_n546_;
  assign new_n549_ = ~new_n547_ & ~new_n548_;
  assign new_n550_ = \2_n169  & ~\2_n174 ;
  assign new_n551_ = ~\2_n169  & \2_n174 ;
  assign new_n552_ = ~new_n550_ & ~new_n551_;
  assign new_n553_ = ~\2_n210  & \2_n59 ;
  assign new_n554_ = \2_n210  & ~\2_n59 ;
  assign new_n555_ = ~new_n553_ & ~new_n554_;
  assign new_n556_ = ~new_n552_ & new_n555_;
  assign new_n557_ = new_n552_ & ~new_n555_;
  assign new_n558_ = ~new_n556_ & ~new_n557_;
  assign new_n559_ = ~new_n549_ & new_n558_;
  assign new_n560_ = new_n549_ & ~new_n558_;
  assign new_n561_ = ~new_n559_ & ~new_n560_;
  assign new_n562_ = ~\2_n187  & \2_n211 ;
  assign new_n563_ = \2_n187  & ~\2_n211 ;
  assign new_n564_ = ~new_n562_ & ~new_n563_;
  assign new_n565_ = ~new_n561_ & new_n564_;
  assign new_n566_ = new_n561_ & ~new_n564_;
  assign new_n567_ = ~new_n565_ & ~new_n566_;
  assign new_n568_ = \2_n133  & \2_n281 ;
  assign new_n569_ = ~\2_n194  & \2_n27 ;
  assign new_n570_ = \2_n194  & ~\2_n27 ;
  assign new_n571_ = ~new_n569_ & ~new_n570_;
  assign new_n572_ = new_n568_ & new_n571_;
  assign new_n573_ = ~new_n568_ & ~new_n571_;
  assign new_n574_ = ~new_n572_ & ~new_n573_;
  assign new_n575_ = ~new_n567_ & new_n574_;
  assign new_n576_ = new_n567_ & ~new_n574_;
  assign new_n577_ = ~new_n575_ & ~new_n576_;
  assign new_n578_ = ~\2_n130  & \2_n256 ;
  assign new_n579_ = \2_n130  & ~\2_n256 ;
  assign new_n580_ = ~new_n578_ & ~new_n579_;
  assign new_n581_ = ~\2_n23  & \2_n43 ;
  assign new_n582_ = \2_n23  & ~\2_n43 ;
  assign new_n583_ = ~new_n581_ & ~new_n582_;
  assign new_n584_ = ~new_n580_ & new_n583_;
  assign new_n585_ = new_n580_ & ~new_n583_;
  assign new_n586_ = ~new_n584_ & ~new_n585_;
  assign new_n587_ = \2_n2  & ~\2_n70 ;
  assign new_n588_ = ~\2_n2  & \2_n70 ;
  assign new_n589_ = ~new_n587_ & ~new_n588_;
  assign new_n590_ = ~\2_n237  & \2_n90 ;
  assign new_n591_ = \2_n237  & ~\2_n90 ;
  assign new_n592_ = ~new_n590_ & ~new_n591_;
  assign new_n593_ = ~new_n589_ & new_n592_;
  assign new_n594_ = new_n589_ & ~new_n592_;
  assign new_n595_ = ~new_n593_ & ~new_n594_;
  assign new_n596_ = ~new_n586_ & new_n595_;
  assign new_n597_ = new_n586_ & ~new_n595_;
  assign new_n598_ = ~new_n596_ & ~new_n597_;
  assign new_n599_ = \2_n0  & ~\2_n179 ;
  assign new_n600_ = ~\2_n0  & \2_n179 ;
  assign new_n601_ = ~new_n599_ & ~new_n600_;
  assign new_n602_ = ~new_n598_ & new_n601_;
  assign new_n603_ = new_n598_ & ~new_n601_;
  assign new_n604_ = ~new_n602_ & ~new_n603_;
  assign new_n605_ = \2_n226  & \2_n281 ;
  assign new_n606_ = ~\2_n137  & \2_n260 ;
  assign new_n607_ = \2_n137  & ~\2_n260 ;
  assign new_n608_ = ~new_n606_ & ~new_n607_;
  assign new_n609_ = new_n605_ & new_n608_;
  assign new_n610_ = ~new_n605_ & ~new_n608_;
  assign new_n611_ = ~new_n609_ & ~new_n610_;
  assign new_n612_ = ~new_n604_ & new_n611_;
  assign new_n613_ = new_n604_ & ~new_n611_;
  assign new_n614_ = ~new_n612_ & ~new_n613_;
  assign new_n615_ = ~new_n577_ & new_n614_;
  assign new_n616_ = ~new_n549_ & new_n586_;
  assign new_n617_ = new_n549_ & ~new_n586_;
  assign new_n618_ = ~new_n616_ & ~new_n617_;
  assign new_n619_ = ~\2_n29  & \2_n75 ;
  assign new_n620_ = \2_n29  & ~\2_n75 ;
  assign new_n621_ = ~new_n619_ & ~new_n620_;
  assign new_n622_ = ~new_n618_ & new_n621_;
  assign new_n623_ = new_n618_ & ~new_n621_;
  assign new_n624_ = ~new_n622_ & ~new_n623_;
  assign new_n625_ = \2_n281  & \2_n84 ;
  assign new_n626_ = \2_n196  & ~\2_n272 ;
  assign new_n627_ = ~\2_n196  & \2_n272 ;
  assign new_n628_ = ~new_n626_ & ~new_n627_;
  assign new_n629_ = new_n625_ & new_n628_;
  assign new_n630_ = ~new_n625_ & ~new_n628_;
  assign new_n631_ = ~new_n629_ & ~new_n630_;
  assign new_n632_ = ~new_n624_ & new_n631_;
  assign new_n633_ = new_n624_ & ~new_n631_;
  assign new_n634_ = ~new_n632_ & ~new_n633_;
  assign new_n635_ = ~new_n558_ & new_n595_;
  assign new_n636_ = new_n558_ & ~new_n595_;
  assign new_n637_ = ~new_n635_ & ~new_n636_;
  assign new_n638_ = \2_n17  & ~\2_n238 ;
  assign new_n639_ = ~\2_n17  & \2_n238 ;
  assign new_n640_ = ~new_n638_ & ~new_n639_;
  assign new_n641_ = ~new_n637_ & new_n640_;
  assign new_n642_ = new_n637_ & ~new_n640_;
  assign new_n643_ = ~new_n641_ & ~new_n642_;
  assign new_n644_ = \2_n281  & \2_n58 ;
  assign new_n645_ = \2_n234  & ~\2_n278 ;
  assign new_n646_ = ~\2_n234  & \2_n278 ;
  assign new_n647_ = ~new_n645_ & ~new_n646_;
  assign new_n648_ = new_n644_ & new_n647_;
  assign new_n649_ = ~new_n644_ & ~new_n647_;
  assign new_n650_ = ~new_n648_ & ~new_n649_;
  assign new_n651_ = ~new_n643_ & new_n650_;
  assign new_n652_ = new_n643_ & ~new_n650_;
  assign new_n653_ = ~new_n651_ & ~new_n652_;
  assign new_n654_ = ~new_n634_ & new_n653_;
  assign new_n655_ = ~\2_n179  & \2_n187 ;
  assign new_n656_ = \2_n179  & ~\2_n187 ;
  assign new_n657_ = ~new_n655_ & ~new_n656_;
  assign new_n658_ = ~\2_n238  & \2_n29 ;
  assign new_n659_ = \2_n238  & ~\2_n29 ;
  assign new_n660_ = ~new_n658_ & ~new_n659_;
  assign new_n661_ = ~new_n657_ & new_n660_;
  assign new_n662_ = new_n657_ & ~new_n660_;
  assign new_n663_ = ~new_n661_ & ~new_n662_;
  assign new_n664_ = ~\2_n137  & \2_n194 ;
  assign new_n665_ = \2_n137  & ~\2_n194 ;
  assign new_n666_ = ~new_n664_ & ~new_n665_;
  assign new_n667_ = \2_n272  & ~\2_n278 ;
  assign new_n668_ = ~\2_n272  & \2_n278 ;
  assign new_n669_ = ~new_n667_ & ~new_n668_;
  assign new_n670_ = ~new_n666_ & new_n669_;
  assign new_n671_ = new_n666_ & ~new_n669_;
  assign new_n672_ = ~new_n670_ & ~new_n671_;
  assign new_n673_ = ~new_n663_ & new_n672_;
  assign new_n674_ = new_n663_ & ~new_n672_;
  assign new_n675_ = ~new_n673_ & ~new_n674_;
  assign new_n676_ = \2_n107  & ~\2_n130 ;
  assign new_n677_ = ~\2_n107  & \2_n130 ;
  assign new_n678_ = ~new_n676_ & ~new_n677_;
  assign new_n679_ = ~new_n675_ & new_n678_;
  assign new_n680_ = new_n675_ & ~new_n678_;
  assign new_n681_ = ~new_n679_ & ~new_n680_;
  assign new_n682_ = \2_n281  & \2_n37 ;
  assign new_n683_ = \2_n174  & ~\2_n70 ;
  assign new_n684_ = ~\2_n174  & \2_n70 ;
  assign new_n685_ = ~new_n683_ & ~new_n684_;
  assign new_n686_ = new_n682_ & new_n685_;
  assign new_n687_ = ~new_n682_ & ~new_n685_;
  assign new_n688_ = ~new_n686_ & ~new_n687_;
  assign new_n689_ = ~new_n681_ & new_n688_;
  assign new_n690_ = new_n681_ & ~new_n688_;
  assign new_n691_ = ~new_n689_ & ~new_n690_;
  assign new_n692_ = ~\2_n0  & \2_n211 ;
  assign new_n693_ = \2_n0  & ~\2_n211 ;
  assign new_n694_ = ~new_n692_ & ~new_n693_;
  assign new_n695_ = ~\2_n17  & \2_n75 ;
  assign new_n696_ = \2_n17  & ~\2_n75 ;
  assign new_n697_ = ~new_n695_ & ~new_n696_;
  assign new_n698_ = ~new_n694_ & new_n697_;
  assign new_n699_ = new_n694_ & ~new_n697_;
  assign new_n700_ = ~new_n698_ & ~new_n699_;
  assign new_n701_ = ~\2_n260  & \2_n27 ;
  assign new_n702_ = \2_n260  & ~\2_n27 ;
  assign new_n703_ = ~new_n701_ & ~new_n702_;
  assign new_n704_ = \2_n196  & ~\2_n234 ;
  assign new_n705_ = ~\2_n196  & \2_n234 ;
  assign new_n706_ = ~new_n704_ & ~new_n705_;
  assign new_n707_ = ~new_n703_ & new_n706_;
  assign new_n708_ = new_n703_ & ~new_n706_;
  assign new_n709_ = ~new_n707_ & ~new_n708_;
  assign new_n710_ = ~new_n700_ & new_n709_;
  assign new_n711_ = new_n700_ & ~new_n709_;
  assign new_n712_ = ~new_n710_ & ~new_n711_;
  assign new_n713_ = ~\2_n256  & \2_n289 ;
  assign new_n714_ = \2_n256  & ~\2_n289 ;
  assign new_n715_ = ~new_n713_ & ~new_n714_;
  assign new_n716_ = ~new_n712_ & new_n715_;
  assign new_n717_ = new_n712_ & ~new_n715_;
  assign new_n718_ = ~new_n716_ & ~new_n717_;
  assign new_n719_ = \2_n18  & \2_n281 ;
  assign new_n720_ = \2_n169  & ~\2_n2 ;
  assign new_n721_ = ~\2_n169  & \2_n2 ;
  assign new_n722_ = ~new_n720_ & ~new_n721_;
  assign new_n723_ = new_n719_ & new_n722_;
  assign new_n724_ = ~new_n719_ & ~new_n722_;
  assign new_n725_ = ~new_n723_ & ~new_n724_;
  assign new_n726_ = ~new_n718_ & new_n725_;
  assign new_n727_ = new_n718_ & ~new_n725_;
  assign new_n728_ = ~new_n726_ & ~new_n727_;
  assign new_n729_ = new_n672_ & ~new_n709_;
  assign new_n730_ = ~new_n672_ & new_n709_;
  assign new_n731_ = ~new_n729_ & ~new_n730_;
  assign new_n732_ = ~\2_n23  & \2_n249 ;
  assign new_n733_ = \2_n23  & ~\2_n249 ;
  assign new_n734_ = ~new_n732_ & ~new_n733_;
  assign new_n735_ = ~new_n731_ & new_n734_;
  assign new_n736_ = new_n731_ & ~new_n734_;
  assign new_n737_ = ~new_n735_ & ~new_n736_;
  assign new_n738_ = \2_n281  & \2_n91 ;
  assign new_n739_ = \2_n210  & ~\2_n237 ;
  assign new_n740_ = ~\2_n210  & \2_n237 ;
  assign new_n741_ = ~new_n739_ & ~new_n740_;
  assign new_n742_ = new_n738_ & new_n741_;
  assign new_n743_ = ~new_n738_ & ~new_n741_;
  assign new_n744_ = ~new_n742_ & ~new_n743_;
  assign new_n745_ = ~new_n737_ & new_n744_;
  assign new_n746_ = new_n737_ & ~new_n744_;
  assign new_n747_ = ~new_n745_ & ~new_n746_;
  assign new_n748_ = new_n663_ & ~new_n700_;
  assign new_n749_ = ~new_n663_ & new_n700_;
  assign new_n750_ = ~new_n748_ & ~new_n749_;
  assign new_n751_ = \2_n214  & ~\2_n43 ;
  assign new_n752_ = ~\2_n214  & \2_n43 ;
  assign new_n753_ = ~new_n751_ & ~new_n752_;
  assign new_n754_ = ~new_n750_ & new_n753_;
  assign new_n755_ = new_n750_ & ~new_n753_;
  assign new_n756_ = ~new_n754_ & ~new_n755_;
  assign new_n757_ = \2_n281  & \2_n292 ;
  assign new_n758_ = \2_n59  & ~\2_n90 ;
  assign new_n759_ = ~\2_n59  & \2_n90 ;
  assign new_n760_ = ~new_n758_ & ~new_n759_;
  assign new_n761_ = new_n757_ & new_n760_;
  assign new_n762_ = ~new_n757_ & ~new_n760_;
  assign new_n763_ = ~new_n761_ & ~new_n762_;
  assign new_n764_ = ~new_n756_ & new_n763_;
  assign new_n765_ = new_n756_ & ~new_n763_;
  assign new_n766_ = ~new_n764_ & ~new_n765_;
  assign new_n767_ = new_n747_ & new_n766_;
  assign new_n768_ = ~new_n728_ & new_n767_;
  assign new_n769_ = new_n691_ & new_n768_;
  assign new_n770_ = new_n654_ & new_n769_;
  assign new_n771_ = new_n615_ & new_n770_;
  assign new_n772_ = \2_n289  & new_n771_;
  assign new_n773_ = ~\2_n289  & ~new_n771_;
  assign \2_n104  = ~new_n772_ & ~new_n773_;
  assign new_n775_ = new_n691_ & ~new_n728_;
  assign new_n776_ = new_n747_ & ~new_n766_;
  assign new_n777_ = new_n634_ & new_n653_;
  assign new_n778_ = new_n614_ & new_n777_;
  assign new_n779_ = ~new_n577_ & new_n778_;
  assign new_n780_ = new_n776_ & new_n779_;
  assign new_n781_ = new_n775_ & new_n780_;
  assign new_n782_ = \2_n211  & new_n781_;
  assign new_n783_ = ~\2_n211  & ~new_n781_;
  assign \2_n123  = ~new_n782_ & ~new_n783_;
  assign new_n785_ = new_n634_ & ~new_n653_;
  assign new_n786_ = new_n691_ & ~new_n747_;
  assign new_n787_ = new_n728_ & new_n766_;
  assign new_n788_ = new_n786_ & new_n787_;
  assign new_n789_ = new_n785_ & new_n788_;
  assign new_n790_ = new_n615_ & new_n789_;
  assign new_n791_ = \2_n210  & new_n790_;
  assign new_n792_ = ~\2_n210  & ~new_n790_;
  assign \2_n129  = ~new_n791_ & ~new_n792_;
  assign new_n794_ = ~new_n691_ & new_n728_;
  assign new_n795_ = ~new_n747_ & new_n766_;
  assign new_n796_ = new_n614_ & ~new_n653_;
  assign new_n797_ = new_n577_ & new_n634_;
  assign new_n798_ = new_n796_ & new_n797_;
  assign new_n799_ = new_n795_ & new_n798_;
  assign new_n800_ = new_n794_ & new_n799_;
  assign new_n801_ = \2_n278  & new_n800_;
  assign new_n802_ = ~\2_n278  & ~new_n800_;
  assign \2_n145  = ~new_n801_ & ~new_n802_;
  assign new_n804_ = new_n775_ & new_n799_;
  assign new_n805_ = \2_n234  & new_n804_;
  assign new_n806_ = ~\2_n234  & ~new_n804_;
  assign \2_n151  = ~new_n805_ & ~new_n806_;
  assign new_n808_ = new_n577_ & ~new_n614_;
  assign new_n809_ = new_n728_ & new_n767_;
  assign new_n810_ = ~new_n691_ & new_n809_;
  assign new_n811_ = new_n785_ & new_n810_;
  assign new_n812_ = new_n808_ & new_n811_;
  assign new_n813_ = \2_n70  & new_n812_;
  assign new_n814_ = ~\2_n70  & ~new_n812_;
  assign \2_n160  = ~new_n813_ & ~new_n814_;
  assign new_n816_ = new_n769_ & new_n785_;
  assign new_n817_ = new_n808_ & new_n816_;
  assign new_n818_ = \2_n2  & new_n817_;
  assign new_n819_ = ~\2_n2  & ~new_n817_;
  assign \2_n164  = ~new_n818_ & ~new_n819_;
  assign new_n821_ = new_n654_ & new_n810_;
  assign new_n822_ = new_n808_ & new_n821_;
  assign new_n823_ = \2_n130  & new_n822_;
  assign new_n824_ = ~\2_n130  & ~new_n822_;
  assign \2_n168  = ~new_n823_ & ~new_n824_;
  assign new_n826_ = new_n780_ & new_n794_;
  assign new_n827_ = \2_n187  & new_n826_;
  assign new_n828_ = ~\2_n187  & ~new_n826_;
  assign \2_n199  = ~new_n827_ & ~new_n828_;
  assign new_n830_ = new_n654_ & new_n788_;
  assign new_n831_ = new_n808_ & new_n830_;
  assign new_n832_ = \2_n23  & new_n831_;
  assign new_n833_ = ~\2_n23  & ~new_n831_;
  assign \2_n212  = ~new_n832_ & ~new_n833_;
  assign new_n835_ = new_n577_ & ~new_n634_;
  assign new_n836_ = new_n614_ & new_n653_;
  assign new_n837_ = new_n835_ & new_n836_;
  assign new_n838_ = new_n776_ & new_n837_;
  assign new_n839_ = new_n775_ & new_n838_;
  assign new_n840_ = \2_n75  & new_n839_;
  assign new_n841_ = ~\2_n75  & ~new_n839_;
  assign \2_n213  = ~new_n840_ & ~new_n841_;
  assign new_n843_ = new_n770_ & new_n808_;
  assign new_n844_ = \2_n256  & new_n843_;
  assign new_n845_ = ~\2_n256  & ~new_n843_;
  assign \2_n217  = ~new_n844_ & ~new_n845_;
  assign new_n847_ = ~new_n614_ & new_n777_;
  assign new_n848_ = new_n577_ & new_n847_;
  assign new_n849_ = new_n776_ & new_n848_;
  assign new_n850_ = new_n794_ & new_n849_;
  assign new_n851_ = \2_n179  & new_n850_;
  assign new_n852_ = ~\2_n179  & ~new_n850_;
  assign \2_n221  = ~new_n851_ & ~new_n852_;
  assign new_n854_ = new_n728_ & ~new_n766_;
  assign new_n855_ = new_n691_ & new_n747_;
  assign new_n856_ = new_n854_ & new_n855_;
  assign new_n857_ = new_n785_ & new_n856_;
  assign new_n858_ = new_n615_ & new_n857_;
  assign new_n859_ = \2_n59  & new_n858_;
  assign new_n860_ = ~\2_n59  & ~new_n858_;
  assign \2_n24  = ~new_n859_ & ~new_n860_;
  assign new_n862_ = new_n615_ & new_n830_;
  assign new_n863_ = \2_n249  & new_n862_;
  assign new_n864_ = ~\2_n249  & ~new_n862_;
  assign \2_n246  = ~new_n863_ & ~new_n864_;
  assign new_n866_ = new_n795_ & new_n837_;
  assign new_n867_ = new_n794_ & new_n866_;
  assign new_n868_ = \2_n272  & new_n867_;
  assign new_n869_ = ~\2_n272  & ~new_n867_;
  assign \2_n253  = ~new_n868_ & ~new_n869_;
  assign new_n871_ = new_n615_ & new_n816_;
  assign new_n872_ = \2_n169  & new_n871_;
  assign new_n873_ = ~\2_n169  & ~new_n871_;
  assign \2_n26  = ~new_n872_ & ~new_n873_;
  assign new_n875_ = new_n775_ & new_n849_;
  assign new_n876_ = \2_n0  & new_n875_;
  assign new_n877_ = ~\2_n0  & ~new_n875_;
  assign \2_n261  = ~new_n876_ & ~new_n877_;
  assign new_n879_ = new_n779_ & new_n795_;
  assign new_n880_ = new_n794_ & new_n879_;
  assign new_n881_ = \2_n194  & new_n880_;
  assign new_n882_ = ~\2_n194  & ~new_n880_;
  assign \2_n265  = ~new_n881_ & ~new_n882_;
  assign new_n884_ = new_n776_ & new_n798_;
  assign new_n885_ = new_n794_ & new_n884_;
  assign new_n886_ = \2_n238  & new_n885_;
  assign new_n887_ = ~\2_n238  & ~new_n885_;
  assign \2_n286  = ~new_n886_ & ~new_n887_;
  assign new_n889_ = new_n654_ & new_n856_;
  assign new_n890_ = new_n615_ & new_n889_;
  assign new_n891_ = \2_n214  & new_n890_;
  assign new_n892_ = ~\2_n214  & ~new_n890_;
  assign \2_n304  = ~new_n891_ & ~new_n892_;
  assign new_n894_ = new_n789_ & new_n808_;
  assign new_n895_ = \2_n237  & new_n894_;
  assign new_n896_ = ~\2_n237  & ~new_n894_;
  assign \2_n310  = ~new_n895_ & ~new_n896_;
  assign new_n898_ = new_n775_ & new_n884_;
  assign new_n899_ = \2_n17  & new_n898_;
  assign new_n900_ = ~\2_n17  & ~new_n898_;
  assign \2_n61  = ~new_n899_ & ~new_n900_;
  assign new_n902_ = new_n794_ & new_n838_;
  assign new_n903_ = \2_n29  & new_n902_;
  assign new_n904_ = ~\2_n29  & ~new_n902_;
  assign \2_n66  = ~new_n903_ & ~new_n904_;
  assign new_n906_ = new_n795_ & new_n848_;
  assign new_n907_ = new_n775_ & new_n906_;
  assign new_n908_ = \2_n260  & new_n907_;
  assign new_n909_ = ~\2_n260  & ~new_n907_;
  assign \2_n73  = ~new_n908_ & ~new_n909_;
  assign new_n911_ = new_n615_ & new_n811_;
  assign new_n912_ = \2_n174  & new_n911_;
  assign new_n913_ = ~\2_n174  & ~new_n911_;
  assign \2_n80  = ~new_n912_ & ~new_n913_;
  assign new_n915_ = new_n808_ & new_n857_;
  assign new_n916_ = \2_n90  & new_n915_;
  assign new_n917_ = ~\2_n90  & ~new_n915_;
  assign \2_n81  = ~new_n916_ & ~new_n917_;
  assign new_n919_ = new_n775_ & new_n866_;
  assign new_n920_ = \2_n196  & new_n919_;
  assign new_n921_ = ~\2_n196  & ~new_n919_;
  assign \2_n86  = ~new_n920_ & ~new_n921_;
  assign new_n923_ = new_n615_ & new_n821_;
  assign new_n924_ = \2_n107  & new_n923_;
  assign new_n925_ = ~\2_n107  & ~new_n923_;
  assign \2_n88  = ~new_n924_ & ~new_n925_;
  assign new_n927_ = new_n808_ & new_n889_;
  assign new_n928_ = \2_n43  & new_n927_;
  assign new_n929_ = ~\2_n43  & ~new_n927_;
  assign \2_n89  = ~new_n928_ & ~new_n929_;
  assign new_n931_ = new_n794_ & new_n906_;
  assign new_n932_ = \2_n137  & new_n931_;
  assign new_n933_ = ~\2_n137  & ~new_n931_;
  assign \2_n94  = ~new_n932_ & ~new_n933_;
  assign new_n935_ = new_n775_ & new_n879_;
  assign new_n936_ = \2_n27  & new_n935_;
  assign new_n937_ = ~\2_n27  & ~new_n935_;
  assign \2_n98  = ~new_n936_ & ~new_n937_;
endmodule


