// Benchmark "top" written by ABC on Sun Jun 11 02:15:05 2023

module top ( 
    \1_n101 , \1_n106 , \1_n107 , \1_n120 , \1_n123 , \1_n136 , \1_n145 ,
    \1_n16 , \1_n165 , \1_n177 , \1_n182 , \1_n216 , \1_n220 , \1_n23 ,
    \1_n24 , \1_n31 , \1_n38 , \1_n41 , \1_n44 , \1_n46 , \1_n53 , \1_n55 ,
    \1_n57 , \1_n62 , \1_n68 , \1_n71 , \1_n72 , \1_n79 , \1_n84 , \1_n92 ,
    \1_n96 , \1_n98 , \2_n100 , \2_n108 , \2_n117 , \2_n123 , \2_n143 ,
    \2_n149 , \2_n151 , \2_n158 , \2_n167 , \2_n189 , \2_n19 , \2_n196 ,
    \2_n197 , \2_n198 , \2_n206 , \2_n209 , \2_n210 , \2_n217 , \2_n218 ,
    \2_n222 , \2_n226 , \2_n233 , \2_n24 , \2_n242 , \2_n258 , \2_n32 ,
    \2_n36 , \2_n49 , \2_n52 , \2_n58 , \2_n59 , \2_n60 , \2_n69 , \2_n73 ,
    \2_n96 , \2_n97 ,
    \1_n126 , \1_n142 , \1_n144 , \1_n153 , \1_n5 , \1_n63 , \1_n78 ,
    \2_n152 , \2_n194 , \2_n224 , \2_n245 , \2_n248 , \2_n29 , \2_n76   );
  input  \1_n101 , \1_n106 , \1_n107 , \1_n120 , \1_n123 , \1_n136 ,
    \1_n145 , \1_n16 , \1_n165 , \1_n177 , \1_n182 , \1_n216 , \1_n220 ,
    \1_n23 , \1_n24 , \1_n31 , \1_n38 , \1_n41 , \1_n44 , \1_n46 , \1_n53 ,
    \1_n55 , \1_n57 , \1_n62 , \1_n68 , \1_n71 , \1_n72 , \1_n79 , \1_n84 ,
    \1_n92 , \1_n96 , \1_n98 , \2_n100 , \2_n108 , \2_n117 , \2_n123 ,
    \2_n143 , \2_n149 , \2_n151 , \2_n158 , \2_n167 , \2_n189 , \2_n19 ,
    \2_n196 , \2_n197 , \2_n198 , \2_n206 , \2_n209 , \2_n210 , \2_n217 ,
    \2_n218 , \2_n222 , \2_n226 , \2_n233 , \2_n24 , \2_n242 , \2_n258 ,
    \2_n32 , \2_n36 , \2_n49 , \2_n52 , \2_n58 , \2_n59 , \2_n60 , \2_n69 ,
    \2_n73 , \2_n96 , \2_n97 ;
  output \1_n126 , \1_n142 , \1_n144 , \1_n153 , \1_n5 , \1_n63 , \1_n78 ,
    \2_n152 , \2_n194 , \2_n224 , \2_n245 , \2_n248 , \2_n29 , \2_n76 ;
  wire new_n83_, new_n84_, new_n85_, new_n86_, new_n87_, new_n88_, new_n89_,
    new_n90_, new_n91_, new_n92_, new_n93_, new_n94_, new_n95_, new_n96_,
    new_n98_, new_n99_, new_n100_, new_n101_, new_n102_, new_n103_,
    new_n104_, new_n105_, new_n106_, new_n107_, new_n108_, new_n109_,
    new_n110_, new_n111_, new_n112_, new_n113_, new_n114_, new_n115_,
    new_n116_, new_n117_, new_n118_, new_n119_, new_n120_, new_n121_,
    new_n122_, new_n123_, new_n124_, new_n125_, new_n126_, new_n127_,
    new_n128_, new_n129_, new_n130_, new_n131_, new_n132_, new_n133_,
    new_n134_, new_n135_, new_n136_, new_n138_, new_n139_, new_n140_,
    new_n141_, new_n142_, new_n143_, new_n144_, new_n145_, new_n146_,
    new_n147_, new_n148_, new_n149_, new_n150_, new_n151_, new_n152_,
    new_n153_, new_n154_, new_n155_, new_n156_, new_n157_, new_n158_,
    new_n159_, new_n160_, new_n161_, new_n162_, new_n163_, new_n164_,
    new_n165_, new_n166_, new_n167_, new_n168_, new_n169_, new_n170_,
    new_n171_, new_n172_, new_n173_, new_n175_, new_n176_, new_n177_,
    new_n178_, new_n179_, new_n180_, new_n181_, new_n182_, new_n183_,
    new_n184_, new_n185_, new_n186_, new_n187_, new_n188_, new_n189_,
    new_n190_, new_n191_, new_n192_, new_n193_, new_n194_, new_n195_,
    new_n196_, new_n197_, new_n198_, new_n199_, new_n200_, new_n201_,
    new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n217_, new_n219_, new_n220_, new_n222_,
    new_n223_, new_n224_, new_n225_, new_n226_, new_n227_, new_n228_,
    new_n229_, new_n230_, new_n232_, new_n233_, new_n234_, new_n235_,
    new_n236_, new_n237_, new_n238_, new_n239_, new_n240_, new_n241_,
    new_n242_, new_n243_, new_n244_, new_n245_, new_n246_, new_n247_,
    new_n249_, new_n250_, new_n251_, new_n252_, new_n253_, new_n254_,
    new_n255_, new_n256_, new_n257_, new_n258_, new_n259_, new_n260_,
    new_n261_, new_n262_, new_n263_, new_n264_, new_n265_, new_n266_,
    new_n267_, new_n268_, new_n269_, new_n270_, new_n271_, new_n272_,
    new_n273_, new_n274_, new_n275_, new_n276_, new_n277_, new_n278_,
    new_n279_, new_n280_, new_n281_, new_n282_, new_n283_, new_n284_,
    new_n285_, new_n286_, new_n287_, new_n288_, new_n289_, new_n290_,
    new_n291_, new_n292_, new_n293_, new_n294_, new_n295_, new_n296_,
    new_n297_, new_n298_, new_n299_, new_n300_, new_n301_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n367_, new_n368_, new_n369_, new_n370_,
    new_n371_, new_n372_, new_n373_, new_n374_, new_n375_, new_n376_,
    new_n377_, new_n378_, new_n379_, new_n380_, new_n381_, new_n382_,
    new_n383_, new_n384_, new_n385_, new_n386_, new_n387_, new_n388_,
    new_n389_, new_n390_, new_n391_, new_n392_, new_n393_, new_n394_,
    new_n395_, new_n396_, new_n397_, new_n398_, new_n399_, new_n400_,
    new_n401_, new_n402_, new_n403_, new_n404_, new_n405_, new_n406_,
    new_n407_, new_n408_, new_n409_, new_n410_, new_n411_, new_n412_,
    new_n413_, new_n415_, new_n416_, new_n417_, new_n418_, new_n420_,
    new_n421_, new_n423_, new_n424_, new_n425_, new_n426_, new_n427_,
    new_n428_, new_n429_, new_n430_, new_n431_, new_n432_, new_n433_,
    new_n434_;
  assign new_n83_ = ~\1_n44  & \1_n53 ;
  assign new_n84_ = ~\1_n41  & \1_n84 ;
  assign new_n85_ = ~new_n83_ & ~new_n84_;
  assign new_n86_ = ~\1_n46  & \1_n182 ;
  assign new_n87_ = new_n85_ & ~new_n86_;
  assign new_n88_ = \1_n38  & ~\1_n71 ;
  assign new_n89_ = new_n87_ & ~new_n88_;
  assign new_n90_ = \1_n96  & ~\1_n98 ;
  assign new_n91_ = new_n89_ & ~new_n90_;
  assign new_n92_ = \1_n55  & ~\1_n165 ;
  assign new_n93_ = new_n91_ & ~new_n92_;
  assign new_n94_ = ~\1_n57  & \1_n68 ;
  assign new_n95_ = new_n93_ & ~new_n94_;
  assign new_n96_ = \1_n84  & ~\1_n101 ;
  assign \1_n5  = ~new_n95_ | new_n96_;
  assign new_n98_ = ~new_n86_ & \1_n5 ;
  assign new_n99_ = ~\1_n220  & ~new_n98_;
  assign new_n100_ = \1_n182  & new_n99_;
  assign new_n101_ = ~\1_n123  & ~new_n98_;
  assign new_n102_ = \1_n182  & new_n101_;
  assign new_n103_ = new_n100_ & new_n102_;
  assign new_n104_ = ~new_n92_ & \1_n5 ;
  assign new_n105_ = ~\1_n16  & ~new_n104_;
  assign new_n106_ = \1_n55  & new_n105_;
  assign new_n107_ = ~\1_n79  & ~new_n104_;
  assign new_n108_ = \1_n55  & new_n107_;
  assign new_n109_ = new_n106_ & new_n108_;
  assign new_n110_ = ~new_n103_ & ~new_n109_;
  assign new_n111_ = ~new_n83_ & \1_n5 ;
  assign new_n112_ = ~\1_n136  & ~new_n111_;
  assign new_n113_ = \1_n53  & new_n112_;
  assign new_n114_ = ~new_n88_ & \1_n5 ;
  assign new_n115_ = ~\1_n23  & ~new_n114_;
  assign new_n116_ = \1_n38  & new_n115_;
  assign new_n117_ = ~new_n96_ & \1_n5 ;
  assign new_n118_ = ~\1_n120  & ~new_n117_;
  assign new_n119_ = \1_n84  & new_n118_;
  assign new_n120_ = ~new_n94_ & \1_n5 ;
  assign new_n121_ = ~\1_n107  & ~new_n120_;
  assign new_n122_ = \1_n68  & new_n121_;
  assign new_n123_ = ~new_n90_ & \1_n5 ;
  assign new_n124_ = ~\1_n72  & ~new_n123_;
  assign new_n125_ = \1_n96  & new_n124_;
  assign new_n126_ = \1_n145  & ~\1_n5 ;
  assign new_n127_ = ~\1_n92  & new_n126_;
  assign new_n128_ = ~new_n125_ & ~new_n127_;
  assign new_n129_ = ~new_n122_ & new_n128_;
  assign new_n130_ = ~new_n108_ & new_n129_;
  assign new_n131_ = ~new_n119_ & new_n130_;
  assign new_n132_ = ~new_n116_ & new_n131_;
  assign new_n133_ = ~new_n113_ & new_n132_;
  assign new_n134_ = ~new_n102_ & new_n133_;
  assign new_n135_ = \1_n84  & ~\1_n5 ;
  assign new_n136_ = ~new_n84_ & ~new_n135_;
  assign \1_n153  = ~new_n134_ | ~new_n136_;
  assign new_n138_ = ~new_n100_ & ~new_n106_;
  assign new_n139_ = ~\1_n153  & ~new_n138_;
  assign new_n140_ = new_n110_ & ~new_n139_;
  assign new_n141_ = \1_n24  & new_n126_;
  assign new_n142_ = new_n127_ & new_n141_;
  assign new_n143_ = ~new_n125_ & \1_n153 ;
  assign new_n144_ = ~new_n123_ & ~new_n143_;
  assign new_n145_ = ~\1_n62  & new_n144_;
  assign new_n146_ = \1_n96  & new_n145_;
  assign new_n147_ = ~new_n142_ & ~new_n146_;
  assign new_n148_ = new_n140_ & new_n147_;
  assign new_n149_ = ~\1_n177  & ~new_n111_;
  assign new_n150_ = \1_n53  & new_n149_;
  assign new_n151_ = new_n113_ & new_n150_;
  assign new_n152_ = ~\1_n216  & ~new_n120_;
  assign new_n153_ = \1_n68  & new_n152_;
  assign new_n154_ = new_n122_ & new_n153_;
  assign new_n155_ = ~new_n151_ & ~new_n154_;
  assign new_n156_ = ~new_n150_ & ~new_n153_;
  assign new_n157_ = ~\1_n153  & ~new_n156_;
  assign new_n158_ = new_n155_ & ~new_n157_;
  assign new_n159_ = \1_n38  & ~new_n114_;
  assign new_n160_ = ~\1_n84  & new_n159_;
  assign new_n161_ = new_n116_ & new_n160_;
  assign new_n162_ = ~\1_n31  & ~new_n117_;
  assign new_n163_ = \1_n84  & new_n162_;
  assign new_n164_ = new_n119_ & new_n163_;
  assign new_n165_ = ~new_n161_ & ~new_n164_;
  assign new_n166_ = ~new_n160_ & ~new_n163_;
  assign new_n167_ = ~\1_n153  & ~new_n166_;
  assign new_n168_ = new_n165_ & ~new_n167_;
  assign new_n169_ = new_n158_ & new_n168_;
  assign new_n170_ = new_n148_ & new_n169_;
  assign new_n171_ = ~\1_n106  & ~new_n136_;
  assign new_n172_ = ~\1_n153  & new_n141_;
  assign new_n173_ = ~new_n171_ & ~new_n172_;
  assign \1_n142  = ~new_n170_ | ~new_n173_;
  assign new_n175_ = \1_n106  & \1_n142 ;
  assign new_n176_ = ~new_n136_ & ~new_n175_;
  assign new_n177_ = \1_n79  & \1_n153 ;
  assign new_n178_ = \1_n165  & \1_n5 ;
  assign new_n179_ = \1_n16  & \1_n142 ;
  assign new_n180_ = ~new_n178_ & ~new_n179_;
  assign new_n181_ = ~new_n177_ & new_n180_;
  assign new_n182_ = \1_n55  & new_n181_;
  assign new_n183_ = \1_n136  & \1_n153 ;
  assign new_n184_ = \1_n44  & \1_n5 ;
  assign new_n185_ = \1_n177  & \1_n142 ;
  assign new_n186_ = ~new_n184_ & ~new_n185_;
  assign new_n187_ = ~new_n183_ & new_n186_;
  assign new_n188_ = \1_n53  & new_n187_;
  assign new_n189_ = new_n182_ & ~new_n188_;
  assign new_n190_ = \1_n107  & \1_n153 ;
  assign new_n191_ = \1_n57  & \1_n5 ;
  assign new_n192_ = \1_n216  & \1_n142 ;
  assign new_n193_ = ~new_n191_ & ~new_n192_;
  assign new_n194_ = ~new_n190_ & new_n193_;
  assign new_n195_ = \1_n68  & new_n194_;
  assign new_n196_ = new_n126_ & ~\1_n142 ;
  assign new_n197_ = ~new_n141_ & ~new_n196_;
  assign new_n198_ = \1_n92  & \1_n153 ;
  assign new_n199_ = ~new_n197_ & ~new_n198_;
  assign new_n200_ = \1_n72  & \1_n153 ;
  assign new_n201_ = \1_n98  & \1_n5 ;
  assign new_n202_ = \1_n62  & \1_n142 ;
  assign new_n203_ = ~new_n201_ & ~new_n202_;
  assign new_n204_ = ~new_n200_ & new_n203_;
  assign new_n205_ = \1_n96  & new_n204_;
  assign new_n206_ = ~new_n199_ & ~new_n205_;
  assign new_n207_ = new_n195_ & new_n206_;
  assign new_n208_ = ~new_n189_ & ~new_n207_;
  assign new_n209_ = ~new_n205_ & new_n208_;
  assign new_n210_ = ~new_n176_ & ~new_n209_;
  assign new_n211_ = ~new_n96_ & ~new_n135_;
  assign new_n212_ = \1_n120  & \1_n153 ;
  assign new_n213_ = ~new_n211_ & ~new_n212_;
  assign new_n214_ = \1_n31  & \1_n142 ;
  assign new_n215_ = new_n213_ & ~new_n214_;
  assign \1_n63  = ~new_n210_ & ~new_n215_;
  assign new_n217_ = ~new_n176_ & ~new_n215_;
  assign \1_n78  = ~new_n206_ | ~new_n217_;
  assign new_n219_ = ~new_n188_ & ~new_n195_;
  assign new_n220_ = new_n206_ & ~new_n219_;
  assign \1_n126  = new_n217_ & ~new_n220_;
  assign new_n222_ = \1_n23  & \1_n153 ;
  assign new_n223_ = \1_n71  & \1_n5 ;
  assign new_n224_ = \1_n84  & \1_n142 ;
  assign new_n225_ = ~new_n223_ & ~new_n224_;
  assign new_n226_ = ~new_n222_ & new_n225_;
  assign new_n227_ = \1_n38  & new_n226_;
  assign new_n228_ = ~new_n182_ & new_n219_;
  assign new_n229_ = ~\1_n78  & new_n228_;
  assign new_n230_ = ~\1_n182  & new_n229_;
  assign \1_n144  = ~new_n227_ & ~new_n230_;
  assign new_n232_ = ~\2_n69  & \2_n73 ;
  assign new_n233_ = ~\2_n151  & \2_n59 ;
  assign new_n234_ = ~\2_n108  & \2_n209 ;
  assign new_n235_ = ~new_n233_ & ~new_n234_;
  assign new_n236_ = ~\2_n210  & \2_n217 ;
  assign new_n237_ = \2_n100  & ~\2_n24 ;
  assign new_n238_ = ~new_n236_ & ~new_n237_;
  assign new_n239_ = new_n235_ & new_n238_;
  assign new_n240_ = ~\2_n218  & \2_n258 ;
  assign new_n241_ = \2_n123  & ~\2_n97 ;
  assign new_n242_ = ~new_n240_ & ~new_n241_;
  assign new_n243_ = \2_n149  & ~\2_n58 ;
  assign new_n244_ = \2_n117  & ~\2_n233 ;
  assign new_n245_ = ~new_n243_ & ~new_n244_;
  assign new_n246_ = new_n242_ & new_n245_;
  assign new_n247_ = new_n239_ & new_n246_;
  assign \2_n29  = new_n232_ | ~new_n247_;
  assign new_n249_ = \2_n151  & \2_n29 ;
  assign new_n250_ = ~new_n232_ & ~\2_n29 ;
  assign new_n251_ = new_n232_ & \2_n29 ;
  assign new_n252_ = ~new_n250_ & ~new_n251_;
  assign new_n253_ = \2_n73  & ~new_n252_;
  assign new_n254_ = ~\2_n242  & new_n253_;
  assign new_n255_ = ~new_n234_ & ~\2_n29 ;
  assign new_n256_ = new_n234_ & \2_n29 ;
  assign new_n257_ = ~new_n255_ & ~new_n256_;
  assign new_n258_ = \2_n209  & ~new_n257_;
  assign new_n259_ = ~\2_n52  & new_n258_;
  assign new_n260_ = ~new_n236_ & ~\2_n29 ;
  assign new_n261_ = new_n236_ & \2_n29 ;
  assign new_n262_ = ~new_n260_ & ~new_n261_;
  assign new_n263_ = \2_n217  & ~new_n262_;
  assign new_n264_ = ~\2_n158  & new_n263_;
  assign new_n265_ = ~new_n259_ & ~new_n264_;
  assign new_n266_ = ~new_n233_ & ~\2_n29 ;
  assign new_n267_ = new_n233_ & \2_n29 ;
  assign new_n268_ = ~new_n266_ & ~new_n267_;
  assign new_n269_ = \2_n59  & ~new_n268_;
  assign new_n270_ = ~\2_n197  & new_n269_;
  assign new_n271_ = ~new_n243_ & ~\2_n29 ;
  assign new_n272_ = new_n243_ & \2_n29 ;
  assign new_n273_ = ~new_n271_ & ~new_n272_;
  assign new_n274_ = \2_n149  & ~new_n273_;
  assign new_n275_ = ~\2_n222  & new_n274_;
  assign new_n276_ = ~new_n270_ & ~new_n275_;
  assign new_n277_ = new_n265_ & new_n276_;
  assign new_n278_ = ~new_n237_ & ~\2_n29 ;
  assign new_n279_ = new_n237_ & \2_n29 ;
  assign new_n280_ = ~new_n278_ & ~new_n279_;
  assign new_n281_ = \2_n100  & ~new_n280_;
  assign new_n282_ = ~\2_n60  & new_n281_;
  assign new_n283_ = ~new_n241_ & ~\2_n29 ;
  assign new_n284_ = new_n241_ & \2_n29 ;
  assign new_n285_ = ~new_n283_ & ~new_n284_;
  assign new_n286_ = \2_n123  & ~new_n285_;
  assign new_n287_ = ~\2_n206  & new_n286_;
  assign new_n288_ = ~new_n282_ & ~new_n287_;
  assign new_n289_ = ~new_n240_ & ~\2_n29 ;
  assign new_n290_ = new_n240_ & \2_n29 ;
  assign new_n291_ = ~new_n289_ & ~new_n290_;
  assign new_n292_ = \2_n258  & ~new_n291_;
  assign new_n293_ = ~\2_n189  & new_n292_;
  assign new_n294_ = ~new_n244_ & ~\2_n29 ;
  assign new_n295_ = new_n244_ & \2_n29 ;
  assign new_n296_ = ~new_n294_ & ~new_n295_;
  assign new_n297_ = \2_n117  & ~new_n296_;
  assign new_n298_ = ~\2_n196  & new_n297_;
  assign new_n299_ = ~new_n293_ & ~new_n298_;
  assign new_n300_ = new_n288_ & new_n299_;
  assign new_n301_ = new_n277_ & new_n300_;
  assign \2_n245  = new_n254_ | ~new_n301_;
  assign new_n303_ = \2_n197  & \2_n245 ;
  assign new_n304_ = ~new_n249_ & ~new_n303_;
  assign new_n305_ = ~\2_n198  & \2_n73 ;
  assign new_n306_ = new_n254_ & ~\2_n245 ;
  assign new_n307_ = ~new_n254_ & \2_n245 ;
  assign new_n308_ = ~new_n306_ & ~new_n307_;
  assign new_n309_ = ~new_n252_ & new_n308_;
  assign new_n310_ = new_n305_ & new_n309_;
  assign new_n311_ = ~\2_n143  & \2_n59 ;
  assign new_n312_ = new_n270_ & ~\2_n245 ;
  assign new_n313_ = ~new_n270_ & \2_n245 ;
  assign new_n314_ = ~new_n312_ & ~new_n313_;
  assign new_n315_ = ~new_n268_ & new_n314_;
  assign new_n316_ = new_n311_ & new_n315_;
  assign new_n317_ = \2_n209  & ~\2_n96 ;
  assign new_n318_ = new_n259_ & ~\2_n245 ;
  assign new_n319_ = ~new_n259_ & \2_n245 ;
  assign new_n320_ = ~new_n318_ & ~new_n319_;
  assign new_n321_ = ~new_n257_ & new_n320_;
  assign new_n322_ = new_n317_ & new_n321_;
  assign new_n323_ = ~new_n316_ & ~new_n322_;
  assign new_n324_ = ~\2_n19  & \2_n217 ;
  assign new_n325_ = new_n264_ & ~\2_n245 ;
  assign new_n326_ = ~new_n264_ & \2_n245 ;
  assign new_n327_ = ~new_n325_ & ~new_n326_;
  assign new_n328_ = ~new_n262_ & new_n327_;
  assign new_n329_ = new_n324_ & new_n328_;
  assign new_n330_ = \2_n100  & ~\2_n167 ;
  assign new_n331_ = new_n282_ & ~\2_n245 ;
  assign new_n332_ = ~new_n282_ & \2_n245 ;
  assign new_n333_ = ~new_n331_ & ~new_n332_;
  assign new_n334_ = ~new_n280_ & new_n333_;
  assign new_n335_ = new_n330_ & new_n334_;
  assign new_n336_ = ~new_n329_ & ~new_n335_;
  assign new_n337_ = new_n323_ & new_n336_;
  assign new_n338_ = \2_n258  & ~\2_n32 ;
  assign new_n339_ = new_n293_ & ~\2_n245 ;
  assign new_n340_ = ~new_n293_ & \2_n245 ;
  assign new_n341_ = ~new_n339_ & ~new_n340_;
  assign new_n342_ = ~new_n291_ & new_n341_;
  assign new_n343_ = new_n338_ & new_n342_;
  assign new_n344_ = \2_n123  & ~\2_n226 ;
  assign new_n345_ = new_n287_ & ~\2_n245 ;
  assign new_n346_ = ~new_n287_ & \2_n245 ;
  assign new_n347_ = ~new_n345_ & ~new_n346_;
  assign new_n348_ = ~new_n285_ & new_n347_;
  assign new_n349_ = new_n344_ & new_n348_;
  assign new_n350_ = ~new_n343_ & ~new_n349_;
  assign new_n351_ = \2_n149  & ~\2_n49 ;
  assign new_n352_ = new_n275_ & ~\2_n245 ;
  assign new_n353_ = ~new_n275_ & \2_n245 ;
  assign new_n354_ = ~new_n352_ & ~new_n353_;
  assign new_n355_ = ~new_n273_ & new_n354_;
  assign new_n356_ = new_n351_ & new_n355_;
  assign new_n357_ = \2_n117  & ~\2_n36 ;
  assign new_n358_ = new_n298_ & ~\2_n245 ;
  assign new_n359_ = ~new_n298_ & \2_n245 ;
  assign new_n360_ = ~new_n358_ & ~new_n359_;
  assign new_n361_ = ~new_n296_ & new_n360_;
  assign new_n362_ = new_n357_ & new_n361_;
  assign new_n363_ = ~new_n356_ & ~new_n362_;
  assign new_n364_ = new_n350_ & new_n363_;
  assign new_n365_ = new_n337_ & new_n364_;
  assign \2_n194  = new_n310_ | ~new_n365_;
  assign new_n367_ = \2_n143  & \2_n194 ;
  assign new_n368_ = \2_n59  & ~new_n367_;
  assign new_n369_ = new_n304_ & new_n368_;
  assign new_n370_ = \2_n108  & \2_n29 ;
  assign new_n371_ = \2_n52  & \2_n245 ;
  assign new_n372_ = ~new_n370_ & ~new_n371_;
  assign new_n373_ = \2_n96  & \2_n194 ;
  assign new_n374_ = \2_n209  & ~new_n373_;
  assign new_n375_ = new_n372_ & new_n374_;
  assign new_n376_ = \2_n210  & \2_n29 ;
  assign new_n377_ = \2_n158  & \2_n245 ;
  assign new_n378_ = ~new_n376_ & ~new_n377_;
  assign new_n379_ = \2_n19  & \2_n194 ;
  assign new_n380_ = \2_n217  & ~new_n379_;
  assign new_n381_ = new_n378_ & new_n380_;
  assign new_n382_ = ~new_n375_ & ~new_n381_;
  assign new_n383_ = \2_n24  & \2_n29 ;
  assign new_n384_ = \2_n60  & \2_n245 ;
  assign new_n385_ = ~new_n383_ & ~new_n384_;
  assign new_n386_ = \2_n167  & \2_n194 ;
  assign new_n387_ = \2_n100  & ~new_n386_;
  assign new_n388_ = new_n385_ & new_n387_;
  assign new_n389_ = \2_n218  & \2_n29 ;
  assign new_n390_ = \2_n189  & \2_n245 ;
  assign new_n391_ = ~new_n389_ & ~new_n390_;
  assign new_n392_ = \2_n32  & \2_n194 ;
  assign new_n393_ = \2_n258  & ~new_n392_;
  assign new_n394_ = new_n391_ & new_n393_;
  assign new_n395_ = ~new_n388_ & new_n394_;
  assign new_n396_ = new_n382_ & new_n395_;
  assign new_n397_ = ~new_n369_ & ~new_n396_;
  assign new_n398_ = ~new_n375_ & new_n381_;
  assign new_n399_ = \2_n97  & \2_n29 ;
  assign new_n400_ = \2_n206  & \2_n245 ;
  assign new_n401_ = ~new_n399_ & ~new_n400_;
  assign new_n402_ = \2_n226  & \2_n194 ;
  assign new_n403_ = \2_n123  & ~new_n402_;
  assign new_n404_ = new_n401_ & new_n403_;
  assign new_n405_ = \2_n58  & \2_n29 ;
  assign new_n406_ = \2_n222  & \2_n245 ;
  assign new_n407_ = ~new_n405_ & ~new_n406_;
  assign new_n408_ = \2_n49  & \2_n194 ;
  assign new_n409_ = \2_n149  & ~new_n408_;
  assign new_n410_ = new_n407_ & new_n409_;
  assign new_n411_ = ~new_n375_ & new_n410_;
  assign new_n412_ = ~new_n404_ & new_n411_;
  assign new_n413_ = ~new_n398_ & ~new_n412_;
  assign \2_n152  = ~new_n397_ | ~new_n413_;
  assign new_n415_ = ~new_n369_ & ~new_n375_;
  assign new_n416_ = ~new_n388_ & new_n404_;
  assign new_n417_ = ~new_n381_ & new_n416_;
  assign new_n418_ = ~new_n396_ & ~new_n417_;
  assign \2_n224  = ~new_n415_ | ~new_n418_;
  assign new_n420_ = ~new_n375_ & ~new_n388_;
  assign new_n421_ = ~new_n369_ & ~new_n398_;
  assign \2_n248  = ~new_n420_ | ~new_n421_;
  assign new_n423_ = ~new_n388_ & ~new_n404_;
  assign new_n424_ = ~new_n394_ & ~new_n410_;
  assign new_n425_ = ~\2_n117  & ~new_n369_;
  assign new_n426_ = new_n424_ & new_n425_;
  assign new_n427_ = new_n423_ & new_n426_;
  assign new_n428_ = new_n382_ & new_n427_;
  assign new_n429_ = \2_n69  & \2_n29 ;
  assign new_n430_ = \2_n242  & \2_n245 ;
  assign new_n431_ = ~new_n429_ & ~new_n430_;
  assign new_n432_ = \2_n198  & \2_n194 ;
  assign new_n433_ = \2_n73  & ~new_n432_;
  assign new_n434_ = new_n431_ & new_n433_;
  assign \2_n76  = ~new_n428_ & ~new_n434_;
endmodule


