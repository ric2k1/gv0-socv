module test(input a, output x, y);
assign x = a, y = a;
endmodule
