module a;
input x[2:0];
endmodule

