module test(input A, output Y, Z);
assign Y = A == A, Z = A != A;
endmodule
