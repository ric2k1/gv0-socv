module top(in1, in2, in3, in4, in5, in6, in7, in8, in9, in10, in11, in12, in13, in14, in15, in16, in17, in18, in19, in20, in21, in22, in23, in24, in25, out1);
  input [8:0] in1, in8, in12, in16, in20, in24;
  input [7:0] in2, in9, in13, in17, in21, in25;
  input in3, in4, in6, in7, in10, in11, in14, in15, in18, in19, in22, in23;
  input [6:0] in5;
  output [16:0] out1;
  wire [8:0] in1, in8, in12, in16, in20, in24;
  wire [7:0] in2, in9, in13, in17, in21, in25;
  wire in3, in4, in6, in7, in10, in11, in14, in15, in18, in19, in22, in23;
  wire [6:0] in5;
  wire [16:0] out1;
  wire w__1, w__2, w__3, w__4, w__5, w__6, w__7, w__8;
  wire w__9, w__10, w__11, w__12, w__13, w__14, w__15, w__16;
  wire w__17, w__18, w__19, w__20, w__21, w__22, w__23, w__24;
  wire w__25, w__26, w__27, w__28, w__29, w__30, w__31, w__32;
  wire w__33, w__34, w__35, w__36, w__37, w__38, w__39, w__40;
  wire w__41, w__42, w__43, w__44, w__45, w__46, w__47, w__48;
  wire w__49, w__50, w__51, w__52, w__53, w__54, w__55, w__56;
  wire w__57, w__58, w__59, w__60, w__61, w__62, w__63, w__64;
  wire w__65, w__66, w__67, w__68, w__69, w__70, w__71, w__72;
  wire w__73, w__74, w__75, w__76, w__77, w__78, w__79, w__80;
  wire w__81, w__82, w__83, w__84, w__85, w__86, w__87, w__88;
  wire w__89, w__90, w__91, w__92, w__93, w__94, w__95, w__96;
  wire w__97, w__98, w__99, w__100, w__101, w__102, w__103, w__104;
  wire w__105, w__106, w__107, w__108, w__109, w__110, w__111, w__112;
  wire w__113, w__114, w__115, w__116, w__117, w__118, w__119, w__120;
  wire w__121, w__122, w__123, w__124, w__125, w__126, w__127, w__128;
  wire w__129, w__130, w__131, w__132, w__133, w__134, w__135, w__136;
  wire w__137, w__138, w__139, w__140, w__141, w__142, w__143, w__144;
  wire w__145, w__146, w__147, w__148, w__149, w__150, w__151, w__152;
  wire w__153, w__154, w__155, w__156, w__157, w__158, w__159, w__160;
  wire w__161, w__162, w__163, w__164, w__165, w__166, w__167, w__168;
  wire w__169, w__170, w__171, w__172, w__173, w__174, w__175, w__176;
  wire w__177, w__178, w__179, w__180, w__181, w__182, w__183, w__184;
  wire w__185, w__186, w__187, w__188, w__189, w__190, w__191, w__192;
  wire w__193, w__194, w__195, w__196, w__197, w__198, w__199, w__200;
  wire w__201, w__202, w__203, w__204, w__205, w__206, w__207, w__208;
  wire w__209, w__210, w__211, w__212, w__213, w__214, w__215, w__216;
  wire w__217, w__218, w__219, w__220, w__221, w__222, w__223, w__224;
  wire w__225, w__226, w__227, w__228, w__229, w__230, w__231, w__232;
  wire w__233, w__234, w__235, w__236, w__237, w__238, w__239, w__240;
  wire w__241, w__242, w__243, w__244, w__245, w__246, w__247, w__248;
  wire w__249, w__250, w__251, w__252, w__253, w__254, w__255, w__256;
  wire w__257, w__258, w__259, w__260, w__261, w__262, w__263, w__264;
  wire w__265, w__266, w__267, w__268, w__269, w__270, w__271, w__272;
  wire w__273, w__274, w__275, w__276, w__277, w__278, w__279, w__280;
  wire w__281, w__282, w__283, w__284, w__285, w__286, w__287, w__288;
  wire w__289, w__290, w__291, w__292, w__293, w__294, w__295, w__296;
  wire w__297, w__298, w__299, w__300, w__301, w__302, w__303, w__304;
  wire w__305, w__306, w__307, w__308, w__309, w__310, w__311, w__312;
  wire w__313, w__314, w__315, w__316, w__317, w__318, w__319, w__320;
  wire w__321, w__322, w__323, w__324, w__325, w__326, w__327, w__328;
  wire w__329, w__330, w__331, w__332, w__333, w__334, w__335, w__336;
  wire w__337, w__338, w__339, w__340, w__341, w__342, w__343, w__344;
  wire w__345, w__346, w__347, w__348, w__349, w__350, w__351, w__352;
  wire w__353, w__354, w__355, w__356, w__357, w__358, w__359, w__360;
  wire w__361, w__362, w__363, w__364, w__365, w__366, w__367, w__368;
  wire w__369, w__370, w__371, w__372, w__373, w__374, w__375, w__376;
  wire w__377, w__378, w__379, w__380, w__381, w__382, w__383, w__384;
  wire w__385, w__386, w__387, w__388, w__389, w__390, w__391, w__392;
  wire w__393, w__394, w__395, w__396, w__397, w__398, w__399, w__400;
  wire w__401, w__402, w__403, w__404, w__405, w__406, w__407, w__408;
  wire w__409, w__410, w__411, w__412, w__413, w__414, w__415, w__416;
  wire w__417, w__418, w__419, w__420, w__421, w__422, w__423, w__424;
  wire w__425, w__426, w__427, w__428, w__429, w__430, w__431, w__432;
  wire w__433, w__434, w__435, w__436, w__437, w__438, w__439, w__440;
  wire w__441, w__442, w__443, w__444, w__445, w__446, w__447, w__448;
  wire w__449, w__450, w__451, w__452, w__453, w__454, w__455, w__456;
  wire w__457, w__458, w__459, w__460, w__461, w__462, w__463, w__464;
  wire w__465, w__466, w__467, w__468, w__469, w__470, w__471, w__472;
  wire w__473, w__474, w__475, w__476, w__477, w__478, w__479, w__480;
  wire w__481, w__482, w__483, w__484, w__485, w__486, w__487, w__488;
  wire w__489, w__490, w__491, w__492, w__493, w__494, w__495, w__496;
  wire w__497, w__498, w__499, w__500, w__501, w__502, w__503, w__504;
  wire w__505, w__506, w__507, w__508, w__509, w__510, w__511, w__512;
  wire w__513, w__514, w__515, w__516, w__517, w__518, w__519, w__520;
  wire w__521, w__522, w__523, w__524, w__525, w__526, w__527, w__528;
  wire w__529, w__530, w__531, w__532, w__533, w__534, w__535, w__536;
  wire w__537, w__538, w__539, w__540, w__541, w__542, w__543, w__544;
  wire w__545, w__546, w__547, w__548, w__549, w__550, w__551, w__552;
  wire w__553, w__554, w__555, w__556, w__557, w__558, w__559, w__560;
  wire w__561, w__562, w__563, w__564, w__565, w__566, w__567, w__568;
  wire w__569, w__570, w__571, w__572, w__573, w__574, w__575, w__576;
  wire w__577, w__578, w__579, w__580, w__581, w__582, w__583, w__584;
  wire w__585, w__586, w__587, w__588, w__589, w__590, w__591, w__592;
  wire w__593, w__594, w__595, w__596, w__597, w__598, w__599, w__600;
  wire w__601, w__602, w__603, w__604, w__605, w__606, w__607, w__608;
  wire w__609, w__610, w__611, w__612, w__613, w__614, w__615, w__616;
  wire w__617, w__618, w__619, w__620, w__621, w__622, w__623, w__624;
  wire w__625, w__626, w__627, w__628, w__629, w__630, w__631, w__632;
  wire w__633, w__634, w__635, w__636, w__637, w__638, w__639, w__640;
  wire w__641, w__642, w__643, w__644, w__645, w__646, w__647, w__648;
  wire w__649, w__650, w__651, w__652, w__653, w__654, w__655, w__656;
  wire w__657, w__658, w__659, w__660, w__661, w__662, w__663, w__664;
  wire w__665, w__666, w__667, w__668, w__669, w__670, w__671, w__672;
  wire w__673, w__674, w__675, w__676, w__677, w__678, w__679, w__680;
  wire w__681, w__682, w__683, w__684, w__685, w__686, w__687, w__688;
  wire w__689, w__690, w__691, w__692, w__693, w__694, w__695, w__696;
  wire w__697, w__698, w__699, w__700, w__701, w__702, w__703, w__704;
  wire w__705, w__706, w__707, w__708, w__709, w__710, w__711, w__712;
  wire w__713, w__714, w__715, w__716, w__717, w__718, w__719, w__720;
  wire w__721, w__722, w__723, w__724, w__725, w__726, w__727, w__728;
  wire w__729, w__730, w__731, w__732, w__733, w__734, w__735, w__736;
  wire w__737, w__738, w__739, w__740, w__741, w__742, w__743, w__744;
  wire w__745, w__746, w__747, w__748, w__749, w__750, w__751, w__752;
  wire w__753, w__754, w__755, w__756, w__757, w__758, w__759, w__760;
  wire w__761, w__762, w__763, w__764, w__765, w__766, w__767, w__768;
  wire w__769, w__770, w__771, w__772, w__773, w__774, w__775, w__776;
  wire w__777, w__778, w__779, w__780, w__781, w__782, w__783, w__784;
  wire w__785, w__786, w__787, w__788, w__789, w__790, w__791, w__792;
  wire w__793, w__794, w__795, w__796, w__797, w__798, w__799, w__800;
  wire w__801, w__802, w__803, w__804, w__805, w__806, w__807, w__808;
  wire w__809, w__810, w__811, w__812, w__813, w__814, w__815, w__816;
  wire w__817, w__818, w__819, w__820, w__821, w__822, w__823, w__824;
  wire w__825, w__826, w__827, w__828, w__829, w__830, w__831, w__832;
  wire w__833, w__834, w__835, w__836, w__837, w__838, w__839, w__840;
  wire w__841, w__842, w__843, w__844, w__845, w__846, w__847, w__848;
  wire w__849, w__850, w__851, w__852, w__853, w__854, w__855, w__856;
  wire w__857, w__858, w__859, w__860, w__861, w__862, w__863, w__864;
  wire w__865, w__866, w__867, w__868, w__869, w__870, w__871, w__872;
  wire w__873, w__874, w__875, w__876, w__877, w__878, w__879, w__880;
  wire w__881, w__882, w__883, w__884, w__885, w__886, w__887, w__888;
  wire w__889, w__890, w__891, w__892, w__893, w__894, w__895, w__896;
  wire w__897, w__898, w__899, w__900, w__901, w__902, w__903, w__904;
  wire w__905, w__906, w__907, w__908, w__909, w__910, w__911, w__912;
  wire w__913, w__914, w__915, w__916, w__917, w__918, w__919, w__920;
  wire w__921, w__922, w__923, w__924, w__925, w__926, w__927, w__928;
  wire w__929, w__930, w__931, w__932, w__933, w__934, w__935, w__936;
  wire w__937, w__938, w__939, w__940, w__941, w__942, w__943, w__944;
  wire w__945, w__946, w__947, w__948, w__949, w__950, w__951, w__952;
  wire w__953, w__954, w__955, w__956, w__957, w__958, w__959, w__960;
  wire w__961, w__962, w__963, w__964, w__965, w__966, w__967, w__968;
  wire w__969, w__970, w__971, w__972, w__973, w__974, w__975, w__976;
  wire w__977, w__978, w__979, w__980, w__981, w__982, w__983, w__984;
  wire w__985, w__986, w__987, w__988, w__989, w__990, w__991, w__992;
  wire w__993, w__994, w__995, w__996, w__997, w__998, w__999, w__1000;
  wire w__1001, w__1002, w__1003, w__1004, w__1005, w__1006, w__1007, w__1008;
  wire w__1009, w__1010, w__1011, w__1012, w__1013, w__1014, w__1015, w__1016;
  wire w__1017, w__1018, w__1019, w__1020, w__1021, w__1022, w__1023, w__1024;
  wire w__1025, w__1026, w__1027, w__1028, w__1029, w__1030, w__1031, w__1032;
  wire w__1033, w__1034, w__1035, w__1036, w__1037, w__1038, w__1039, w__1040;
  wire w__1041, w__1042, w__1043, w__1044, w__1045, w__1046, w__1047, w__1048;
  wire w__1049, w__1050, w__1051, w__1052, w__1053, w__1054, w__1055, w__1056;
  wire w__1057, w__1058, w__1059, w__1060, w__1061, w__1062, w__1063, w__1064;
  wire w__1065, w__1066, w__1067, w__1068, w__1069, w__1070, w__1071, w__1072;
  wire w__1073, w__1074, w__1075, w__1076, w__1077, w__1078, w__1079, w__1080;
  wire w__1081, w__1082, w__1083, w__1084, w__1085, w__1086, w__1087, w__1088;
  wire w__1089, w__1090, w__1091, w__1092, w__1093, w__1094, w__1095, w__1096;
  wire w__1097, w__1098, w__1099, w__1100, w__1101, w__1102, w__1103, w__1104;
  wire w__1105, w__1106, w__1107, w__1108, w__1109, w__1110, w__1111, w__1112;
  wire w__1113, w__1114, w__1115, w__1116, w__1117, w__1118, w__1119, w__1120;
  wire w__1121, w__1122, w__1123, w__1124, w__1125, w__1126, w__1127, w__1128;
  wire w__1129, w__1130, w__1131, w__1132, w__1133, w__1134, w__1135, w__1136;
  wire w__1137, w__1138, w__1139, w__1140, w__1141, w__1142, w__1143, w__1144;
  wire w__1145, w__1146, w__1147, w__1148, w__1149, w__1150, w__1151, w__1152;
  wire w__1153, w__1154, w__1155, w__1156, w__1157, w__1158, w__1159, w__1160;
  wire w__1161, w__1162, w__1163, w__1164, w__1165, w__1166, w__1167, w__1168;
  wire w__1169, w__1170, w__1171, w__1172, w__1173, w__1174, w__1175, w__1176;
  wire w__1177, w__1178, w__1179, w__1180, w__1181, w__1182, w__1183, w__1184;
  wire w__1185, w__1186, w__1187, w__1188, w__1189, w__1190, w__1191, w__1192;
  wire w__1193, w__1194, w__1195, w__1196, w__1197, w__1198, w__1199, w__1200;
  wire w__1201, w__1202, w__1203, w__1204, w__1205, w__1206, w__1207, w__1208;
  wire w__1209, w__1210, w__1211, w__1212, w__1213, w__1214, w__1215, w__1216;
  wire w__1217, w__1218, w__1219, w__1220, w__1221, w__1222, w__1223, w__1224;
  wire w__1225, w__1226, w__1227, w__1228, w__1229, w__1230, w__1231, w__1232;
  wire w__1233, w__1234, w__1235, w__1236, w__1237, w__1238, w__1239, w__1240;
  wire w__1241, w__1242, w__1243, w__1244, w__1245, w__1246, w__1247, w__1248;
  wire w__1249, w__1250, w__1251, w__1252, w__1253, w__1254, w__1255, w__1256;
  wire w__1257, w__1258, w__1259, w__1260, w__1261, w__1262, w__1263, w__1264;
  wire w__1265, w__1266, w__1267, w__1268, w__1269, w__1270, w__1271, w__1272;
  wire w__1273, w__1274, w__1275, w__1276, w__1277, w__1278, w__1279, w__1280;
  wire w__1281, w__1282, w__1283, w__1284, w__1285, w__1286, w__1287, w__1288;
  wire w__1289, w__1290, w__1291, w__1292, w__1293, w__1294, w__1295, w__1296;
  wire w__1297, w__1298, w__1299, w__1300, w__1301, w__1302, w__1303, w__1304;
  wire w__1305, w__1306, w__1307, w__1308, w__1309, w__1310, w__1311, w__1312;
  wire w__1313, w__1314, w__1315, w__1316, w__1317, w__1318, w__1319, w__1320;
  wire w__1321, w__1322, w__1323, w__1324, w__1325, w__1326, w__1327, w__1328;
  wire w__1329, w__1330, w__1331, w__1332, w__1333, w__1334, w__1335, w__1336;
  wire w__1337, w__1338, w__1339, w__1340, w__1341, w__1342, w__1343, w__1344;
  wire w__1345, w__1346, w__1347, w__1348, w__1349, w__1350, w__1351, w__1352;
  wire w__1353, w__1354, w__1355, w__1356, w__1357, w__1358, w__1359, w__1360;
  wire w__1361, w__1362, w__1363, w__1364, w__1365, w__1366, w__1367, w__1368;
  wire w__1369, w__1370, w__1371, w__1372, w__1373, w__1374, w__1375, w__1376;
  wire w__1377, w__1378, w__1379, w__1380, w__1381, w__1382, w__1383, w__1384;
  wire w__1385, w__1386, w__1387, w__1388, w__1389, w__1390, w__1391, w__1392;
  wire w__1393, w__1394, w__1395, w__1396, w__1397, w__1398, w__1399, w__1400;
  wire w__1401, w__1402, w__1403, w__1404, w__1405, w__1406, w__1407, w__1408;
  wire w__1409, w__1410, w__1411, w__1412, w__1413, w__1414, w__1415, w__1416;
  wire w__1417, w__1418, w__1419, w__1420, w__1421, w__1422, w__1423, w__1424;
  wire w__1425, w__1426, w__1427, w__1428, w__1429, w__1430, w__1431, w__1432;
  wire w__1433, w__1434, w__1435, w__1436, w__1437, w__1438, w__1439, w__1440;
  wire w__1441, w__1442, w__1443, w__1444, w__1445, w__1446, w__1447, w__1448;
  wire w__1449, w__1450, w__1451, w__1452, w__1453, w__1454, w__1455, w__1456;
  wire w__1457, w__1458, w__1459, w__1460, w__1461, w__1462, w__1463, w__1464;
  wire w__1465, w__1466, w__1467, w__1468, w__1469, w__1470, w__1471, w__1472;
  wire w__1473, w__1474, w__1475, w__1476, w__1477, w__1478, w__1479, w__1480;
  wire w__1481, w__1482, w__1483, w__1484, w__1485, w__1486, w__1487, w__1488;
  wire w__1489, w__1490, w__1491, w__1492, w__1493, w__1494, w__1495, w__1496;
  wire w__1497, w__1498, w__1499, w__1500, w__1501, w__1502, w__1503, w__1504;
  wire w__1505, w__1506, w__1507, w__1508, w__1509, w__1510, w__1511, w__1512;
  wire w__1513, w__1514, w__1515, w__1516, w__1517, w__1518, w__1519, w__1520;
  wire w__1521, w__1522, w__1523, w__1524, w__1525, w__1526, w__1527, w__1528;
  wire w__1529, w__1530, w__1531, w__1532, w__1533, w__1534, w__1535, w__1536;
  wire w__1537, w__1538, w__1539, w__1540, w__1541, w__1542, w__1543, w__1544;
  wire w__1545, w__1546, w__1547, w__1548, w__1549, w__1550, w__1551, w__1552;
  wire w__1553, w__1554, w__1555, w__1556, w__1557, w__1558, w__1559, w__1560;
  wire w__1561, w__1562, w__1563, w__1564, w__1565, w__1566, w__1567, w__1568;
  wire w__1569, w__1570, w__1571, w__1572, w__1573, w__1574, w__1575, w__1576;
  wire w__1577, w__1578, w__1579, w__1580, w__1581, w__1582, w__1583, w__1584;
  wire w__1585, w__1586, w__1587, w__1588, w__1589, w__1590, w__1591, w__1592;
  wire w__1593, w__1594, w__1595, w__1596, w__1597, w__1598, w__1599, w__1600;
  wire w__1601, w__1602, w__1603, w__1604, w__1605, w__1606, w__1607, w__1608;
  wire w__1609, w__1610, w__1611, w__1612, w__1613, w__1614, w__1615, w__1616;
  wire w__1617, w__1618, w__1619, w__1620, w__1621, w__1622, w__1623, w__1624;
  wire w__1625, w__1626, w__1627, w__1628, w__1629, w__1630, w__1631, w__1632;
  wire w__1633, w__1634, w__1635, w__1636, w__1637, w__1638, w__1639, w__1640;
  wire w__1641, w__1642, w__1643, w__1644, w__1645, w__1646, w__1647, w__1648;
  wire w__1649, w__1650, w__1651, w__1652, w__1653, w__1654, w__1655, w__1656;
  wire w__1657, w__1658, w__1659, w__1660, w__1661, w__1662, w__1663, w__1664;
  wire w__1665, w__1666, w__1667, w__1668, w__1669, w__1670, w__1671, w__1672;
  wire w__1673, w__1674, w__1675, w__1676, w__1677, w__1678, w__1679, w__1680;
  wire w__1681, w__1682, w__1683, w__1684, w__1685, w__1686, w__1687, w__1688;
  wire w__1689, w__1690, w__1691, w__1692, w__1693, w__1694, w__1695, w__1696;
  wire w__1697, w__1698, w__1699, w__1700, w__1701, w__1702, w__1703, w__1704;
  wire w__1705, w__1706, w__1707, w__1708, w__1709, w__1710, w__1711, w__1712;
  wire w__1713, w__1714, w__1715, w__1716, w__1717, w__1718, w__1719, w__1720;
  wire w__1721, w__1722, w__1723, w__1724, w__1725, w__1726, w__1727, w__1728;
  wire w__1729, w__1730, w__1731, w__1732, w__1733, w__1734, w__1735, w__1736;
  wire w__1737, w__1738, w__1739, w__1740, w__1741, w__1742, w__1743, w__1744;
  wire w__1745, w__1746, w__1747, w__1748, w__1749, w__1750, w__1751, w__1752;
  wire w__1753, w__1754, w__1755, w__1756, w__1757, w__1758, w__1759, w__1760;
  wire w__1761, w__1762, w__1763, w__1764, w__1765, w__1766, w__1767, w__1768;
  wire w__1769, w__1770, w__1771, w__1772, w__1773, w__1774, w__1775, w__1776;
  wire w__1777, w__1778, w__1779, w__1780, w__1781, w__1782, w__1783, w__1784;
  wire w__1785, w__1786, w__1787, w__1788, w__1789, w__1790, w__1791, w__1792;
  wire w__1793, w__1794, w__1795, w__1796, w__1797, w__1798, w__1799, w__1800;
  wire w__1801, w__1802, w__1803, w__1804, w__1805, w__1806, w__1807, w__1808;
  wire w__1809, w__1810, w__1811, w__1812, w__1813, w__1814, w__1815, w__1816;
  wire w__1817, w__1818, w__1819, w__1820, w__1821, w__1822, w__1823, w__1824;
  wire w__1825, w__1826, w__1827, w__1828, w__1829, w__1830, w__1831, w__1832;
  wire w__1833, w__1834, w__1835, w__1836, w__1837, w__1838, w__1839, w__1840;
  wire w__1841, w__1842, w__1843, w__1844, w__1845, w__1846, w__1847, w__1848;
  wire w__1849, w__1850, w__1851, w__1852, w__1853, w__1854, w__1855, w__1856;
  wire w__1857, w__1858, w__1859, w__1860, w__1861, w__1862, w__1863, w__1864;
  wire w__1865, w__1866, w__1867, w__1868, w__1869, w__1870, w__1871, w__1872;
  wire w__1873, w__1874, w__1875, w__1876, w__1877, w__1878, w__1879, w__1880;
  wire w__1881, w__1882, w__1883, w__1884, w__1885, w__1886, w__1887, w__1888;
  wire w__1889, w__1890, w__1891, w__1892, w__1893, w__1894, w__1895, w__1896;
  wire w__1897, w__1898, w__1899, w__1900, w__1901, w__1902, w__1903, w__1904;
  wire w__1905, w__1906, w__1907, w__1908, w__1909, w__1910, w__1911, w__1912;
  wire w__1913, w__1914, w__1915, w__1916, w__1917, w__1918, w__1919, w__1920;
  wire w__1921, w__1922, w__1923, w__1924, w__1925, w__1926, w__1927, w__1928;
  wire w__1929, w__1930, w__1931, w__1932, w__1933, w__1934, w__1935, w__1936;
  wire w__1937, w__1938, w__1939, w__1940, w__1941, w__1942, w__1943, w__1944;
  wire w__1945, w__1946, w__1947, w__1948, w__1949, w__1950, w__1951, w__1952;
  wire w__1953, w__1954, w__1955, w__1956, w__1957, w__1958, w__1959, w__1960;
  wire w__1961, w__1962, w__1963, w__1964, w__1965, w__1966, w__1967, w__1968;
  wire w__1969, w__1970, w__1971, w__1972, w__1973, w__1974, w__1975, w__1976;
  wire w__1977, w__1978, w__1979, w__1980, w__1981, w__1982, w__1983, w__1984;
  wire w__1985, w__1986, w__1987, w__1988, w__1989, w__1990, w__1991, w__1992;
  wire w__1993, w__1994, w__1995, w__1996, w__1997, w__1998, w__1999, w__2000;
  wire w__2001, w__2002, w__2003, w__2004, w__2005, w__2006, w__2007, w__2008;
  wire w__2009, w__2010, w__2011, w__2012, w__2013, w__2014, w__2015, w__2016;
  wire w__2017, w__2018, w__2019, w__2020, w__2021, w__2022, w__2023, w__2024;
  wire w__2025, w__2026, w__2027, w__2028, w__2029, w__2030, w__2031, w__2032;
  wire w__2033, w__2034, w__2035, w__2036, w__2037, w__2038, w__2039, w__2040;
  wire w__2041, w__2042, w__2043, w__2044, w__2045, w__2046, w__2047, w__2048;
  wire w__2049, w__2050, w__2051, w__2052, w__2053, w__2054, w__2055, w__2056;
  wire w__2057, w__2058, w__2059, w__2060, w__2061, w__2062, w__2063, w__2064;
  wire w__2065, w__2066, w__2067, w__2068, w__2069, w__2070, w__2071, w__2072;
  wire w__2073, w__2074, w__2075, w__2076, w__2077, w__2078, w__2079, w__2080;
  wire w__2081, w__2082, w__2083, w__2084, w__2085, w__2086, w__2087, w__2088;
  wire w__2089, w__2090, w__2091, w__2092, w__2093, w__2094, w__2095, w__2096;
  wire w__2097, w__2098, w__2099, w__2100, w__2101, w__2102, w__2103, w__2104;
  wire w__2105, w__2106, w__2107, w__2108, w__2109, w__2110, w__2111, w__2112;
  wire w__2113, w__2114, w__2115, w__2116, w__2117, w__2118, w__2119, w__2120;
  wire w__2121, w__2122, w__2123, w__2124, w__2125, w__2126, w__2127, w__2128;
  wire w__2129, w__2130, w__2131, w__2132, w__2133, w__2134, w__2135, w__2136;
  wire w__2137, w__2138, w__2139, w__2140, w__2141, w__2142, w__2143, w__2144;
  wire w__2145, w__2146, w__2147, w__2148, w__2149, w__2150, w__2151, w__2152;
  wire w__2153, w__2154, w__2155, w__2156, w__2157, w__2158, w__2159, w__2160;
  wire w__2161, w__2162, w__2163, w__2164, w__2165, w__2166, w__2167, w__2168;
  wire w__2169, w__2170, w__2171, w__2172, w__2173, w__2174, w__2175, w__2176;
  wire w__2177, w__2178, w__2179, w__2180, w__2181, w__2182, w__2183, w__2184;
  wire w__2185, w__2186, w__2187, w__2188, w__2189, w__2190, w__2191, w__2192;
  wire w__2193, w__2194, w__2195, w__2196, w__2197, w__2198, w__2199, w__2200;
  wire w__2201, w__2202, w__2203, w__2204, w__2205, w__2206, w__2207, w__2208;
  wire w__2209, w__2210, w__2211, w__2212, w__2213, w__2214, w__2215, w__2216;
  wire w__2217, w__2218, w__2219, w__2220, w__2221, w__2222, w__2223, w__2224;
  wire w__2225, w__2226, w__2227, w__2228, w__2229, w__2230, w__2231, w__2232;
  wire w__2233, w__2234, w__2235, w__2236, w__2237, w__2238, w__2239, w__2240;
  wire w__2241, w__2242, w__2243, w__2244, w__2245, w__2246, w__2247, w__2248;
  wire w__2249, w__2250, w__2251, w__2252, w__2253, w__2254, w__2255, w__2256;
  wire w__2257, w__2258, w__2259, w__2260, w__2261, w__2262, w__2263, w__2264;
  wire w__2265, w__2266, w__2267, w__2268, w__2269, w__2270, w__2271, w__2272;
  wire w__2273, w__2274, w__2275, w__2276, w__2277, w__2278, w__2279, w__2280;
  wire w__2281, w__2282, w__2283, w__2284, w__2285, w__2286, w__2287, w__2288;
  wire w__2289, w__2290, w__2291, w__2292, w__2293, w__2294, w__2295, w__2296;
  wire w__2297, w__2298, w__2299, w__2300, w__2301, w__2302, w__2303, w__2304;
  wire w__2305, w__2306, w__2307, w__2308, w__2309, w__2310, w__2311, w__2312;
  wire w__2313, w__2314, w__2315, w__2316, w__2317, w__2318, w__2319, w__2320;
  wire w__2321, w__2322, w__2323, w__2324, w__2325, w__2326, w__2327, w__2328;
  wire w__2329, w__2330, w__2331, w__2332, w__2333, w__2334, w__2335, w__2336;
  wire w__2337, w__2338, w__2339, w__2340, w__2341, w__2342, w__2343, w__2344;
  wire w__2345, w__2346, w__2347, w__2348, w__2349, w__2350, w__2351, w__2352;
  wire w__2353, w__2354, w__2355, w__2356, w__2357, w__2358, w__2359, w__2360;
  wire w__2361, w__2362, w__2363, w__2364, w__2365, w__2366, w__2367, w__2368;
  wire w__2369, w__2370, w__2371, w__2372, w__2373, w__2374, w__2375, w__2376;
  wire w__2377, w__2378, w__2379, w__2380, w__2381, w__2382, w__2383, w__2384;
  wire w__2385, w__2386, w__2387, w__2388, w__2389, w__2390, w__2391, w__2392;
  wire w__2393, w__2394, w__2395, w__2396, w__2397, w__2398, w__2399, w__2400;
  wire w__2401, w__2402, w__2403, w__2404, w__2405, w__2406, w__2407, w__2408;
  wire w__2409, w__2410, w__2411, w__2412, w__2413, w__2414, w__2415, w__2416;
  wire w__2417, w__2418, w__2419, w__2420, w__2421, w__2422, w__2423, w__2424;
  wire w__2425, w__2426, w__2427, w__2428, w__2429, w__2430, w__2431, w__2432;
  wire w__2433, w__2434, w__2435, w__2436, w__2437, w__2438, w__2439, w__2440;
  wire w__2441, w__2442, w__2443, w__2444, w__2445, w__2446, w__2447, w__2448;
  wire w__2449, w__2450, w__2451, w__2452, w__2453, w__2454, w__2455, w__2456;
  wire w__2457, w__2458, w__2459, w__2460, w__2461, w__2462, w__2463, w__2464;
  wire w__2465, w__2466, w__2467, w__2468, w__2469, w__2470, w__2471, w__2472;
  wire w__2473, w__2474, w__2475, w__2476, w__2477, w__2478, w__2479, w__2480;
  wire w__2481, w__2482, w__2483, w__2484, w__2485, w__2486, w__2487, w__2488;
  wire w__2489, w__2490, w__2491, w__2492, w__2493, w__2494, w__2495, w__2496;
  wire w__2497, w__2498, w__2499, w__2500, w__2501, w__2502, w__2503, w__2504;
  wire w__2505, w__2506, w__2507, w__2508, w__2509, w__2510, w__2511, w__2512;
  wire w__2513, w__2514, w__2515, w__2516, w__2517, w__2518, w__2519, w__2520;
  wire w__2521, w__2522, w__2523, w__2524, w__2525, w__2526, w__2527, w__2528;
  wire w__2529, w__2530, w__2531, w__2532, w__2533, w__2534, w__2535, w__2536;
  wire w__2537, w__2538, w__2539, w__2540, w__2541, w__2542, w__2543, w__2544;
  wire w__2545, w__2546, w__2547, w__2548, w__2549, w__2550, w__2551, w__2552;
  wire w__2553, w__2554, w__2555, w__2556, w__2557, w__2558, w__2559, w__2560;
  wire w__2561, w__2562, w__2563, w__2564, w__2565, w__2566, w__2567, w__2568;
  wire w__2569, w__2570, w__2571, w__2572, w__2573, w__2574, w__2575, w__2576;
  wire w__2577, w__2578, w__2579, w__2580, w__2581, w__2582, w__2583, w__2584;
  wire w__2585, w__2586, w__2587, w__2588, w__2589, w__2590, w__2591, w__2592;
  wire w__2593, w__2594, w__2595, w__2596, w__2597, w__2598, w__2599, w__2600;
  wire w__2601, w__2602, w__2603, w__2604, w__2605, w__2606, w__2607, w__2608;
  wire w__2609, w__2610, w__2611, w__2612, w__2613, w__2614, w__2615, w__2616;
  wire w__2617, w__2618, w__2619, w__2620, w__2621, w__2622, w__2623, w__2624;
  wire w__2625, w__2626, w__2627, w__2628, w__2629, w__2630, w__2631, w__2632;
  wire w__2633, w__2634, w__2635, w__2636, w__2637, w__2638, w__2639, w__2640;
  wire w__2641, w__2642, w__2643, w__2644, w__2645, w__2646, w__2647, w__2648;
  wire w__2649, w__2650, w__2651, w__2652, w__2653, w__2654, w__2655, w__2656;
  wire w__2657, w__2658, w__2659, w__2660, w__2661, w__2662, w__2663, w__2664;
  wire w__2665, w__2666, w__2667, w__2668, w__2669, w__2670, w__2671, w__2672;
  wire w__2673, w__2674, w__2675, w__2676, w__2677, w__2678, w__2679, w__2680;
  wire w__2681, w__2682, w__2683, w__2684, w__2685, w__2686, w__2687, w__2688;
  wire w__2689, w__2690, w__2691, w__2692, w__2693, w__2694, w__2695, w__2696;
  wire w__2697, w__2698, w__2699, w__2700, w__2701, w__2702, w__2703, w__2704;
  wire w__2705, w__2706, w__2707, w__2708, w__2709, w__2710, w__2711, w__2712;
  wire w__2713, w__2714, w__2715, w__2716, w__2717, w__2718, w__2719, w__2720;
  wire w__2721, w__2722, w__2723, w__2724, w__2725, w__2726, w__2727, w__2728;
  wire w__2729, w__2730, w__2731, w__2732, w__2733, w__2734, w__2735, w__2736;
  wire w__2737, w__2738, w__2739, w__2740, w__2741, w__2742, w__2743, w__2744;
  wire w__2745, w__2746, w__2747, w__2748, w__2749, w__2750, w__2751, w__2752;
  wire w__2753, w__2754, w__2755, w__2756, w__2757, w__2758, w__2759, w__2760;
  wire w__2761, w__2762, w__2763, w__2764, w__2765, w__2766, w__2767, w__2768;
  wire w__2769, w__2770, w__2771, w__2772, w__2773, w__2774, w__2775, w__2776;
  wire w__2777, w__2778, w__2779, w__2780, w__2781, w__2782, w__2783, w__2784;
  wire w__2785, w__2786, w__2787, w__2788, w__2789, w__2790, w__2791, w__2792;
  wire w__2793, w__2794, w__2795, w__2796, w__2797, w__2798, w__2799, w__2800;
  wire w__2801, w__2802, w__2803, w__2804, w__2805, w__2806, w__2807, w__2808;
  wire w__2809, w__2810, w__2811, w__2812, w__2813, w__2814, w__2815, w__2816;
  wire w__2817, w__2818, w__2819, w__2820, w__2821, w__2822, w__2823, w__2824;
  wire w__2825, w__2826, w__2827, w__2828, w__2829, w__2830, w__2831, w__2832;
  wire w__2833, w__2834, w__2835, w__2836, w__2837, w__2838, w__2839, w__2840;
  wire w__2841, w__2842, w__2843, w__2844, w__2845, w__2846, w__2847, w__2848;
  wire w__2849, w__2850, w__2851, w__2852, w__2853, w__2854, w__2855, w__2856;
  wire w__2857, w__2858, w__2859, w__2860, w__2861, w__2862, w__2863, w__2864;
  wire w__2865, w__2866, w__2867, w__2868, w__2869, w__2870, w__2871, w__2872;
  wire w__2873, w__2874, w__2875, w__2876, w__2877, w__2878, w__2879, w__2880;
  wire w__2881, w__2882, w__2883, w__2884, w__2885, w__2886, w__2887, w__2888;
  wire w__2889, w__2890, w__2891, w__2892, w__2893, w__2894, w__2895, w__2896;
  wire w__2897, w__2898, w__2899, w__2900, w__2901, w__2902, w__2903, w__2904;
  wire w__2905, w__2906, w__2907, w__2908, w__2909, w__2910, w__2911, w__2912;
  wire w__2913, w__2914, w__2915, w__2916, w__2917, w__2918, w__2919, w__2920;
  wire w__2921, w__2922, w__2923, w__2924, w__2925, w__2926, w__2927, w__2928;
  wire w__2929, w__2930, w__2931, w__2932, w__2933, w__2934, w__2935, w__2936;
  wire w__2937, w__2938, w__2939, w__2940, w__2941, w__2942, w__2943, w__2944;
  wire w__2945, w__2946, w__2947, w__2948, w__2949, w__2950, w__2951, w__2952;
  wire w__2953, w__2954, w__2955, w__2956, w__2957, w__2958, w__2959, w__2960;
  wire w__2961, w__2962, w__2963, w__2964, w__2965, w__2966, w__2967, w__2968;
  wire w__2969, w__2970, w__2971, w__2972, w__2973, w__2974, w__2975, w__2976;
  wire w__2977, w__2978, w__2979, w__2980, w__2981, w__2982, w__2983, w__2984;
  wire w__2985, w__2986, w__2987, w__2988, w__2989, w__2990, w__2991, w__2992;
  wire w__2993, w__2994, w__2995, w__2996, w__2997, w__2998, w__2999, w__3000;
  wire w__3001, w__3002, w__3003, w__3004, w__3005, w__3006, w__3007, w__3008;
  wire w__3009, w__3010, w__3011, w__3012, w__3013, w__3014, w__3015, w__3016;
  wire w__3017, w__3018, w__3019, w__3020, w__3021, w__3022, w__3023, w__3024;
  wire w__3025, w__3026, w__3027, w__3028, w__3029, w__3030, w__3031, w__3032;
  wire w__3033, w__3034, w__3035, w__3036, w__3037, w__3038, w__3039, w__3040;
  wire w__3041, w__3042, w__3043, w__3044, w__3045, w__3046, w__3047, w__3048;
  wire w__3049, w__3050, w__3051, w__3052, w__3053, w__3054, w__3055, w__3056;
  wire w__3057, w__3058, w__3059, w__3060, w__3061, w__3062, w__3063, w__3064;
  wire w__3065, w__3066, w__3067, w__3068, w__3069, w__3070, w__3071, w__3072;
  wire w__3073, w__3074, w__3075, w__3076, w__3077, w__3078, w__3079, w__3080;
  wire w__3081, w__3082, w__3083, w__3084, w__3085, w__3086, w__3087, w__3088;
  wire w__3089, w__3090, w__3091, w__3092, w__3093, w__3094, w__3095, w__3096;
  wire w__3097, w__3098, w__3099, w__3100, w__3101, w__3102, w__3103, w__3104;
  wire w__3105, w__3106, w__3107, w__3108, w__3109, w__3110, w__3111, w__3112;
  wire w__3113, w__3114, w__3115, w__3116, w__3117, w__3118, w__3119, w__3120;
  wire w__3121, w__3122, w__3123, w__3124, w__3125, w__3126, w__3127, w__3128;
  wire w__3129, w__3130, w__3131, w__3132, w__3133, w__3134, w__3135, w__3136;
  wire w__3137, w__3138, w__3139, w__3140, w__3141, w__3142, w__3143, w__3144;
  wire w__3145, w__3146, w__3147, w__3148, w__3149, w__3150, w__3151, w__3152;
  wire w__3153, w__3154, w__3155, w__3156, w__3157, w__3158, w__3159, w__3160;
  wire w__3161, w__3162, w__3163, w__3164, w__3165, w__3166, w__3167, w__3168;
  wire w__3169, w__3170, w__3171, w__3172, w__3173, w__3174, w__3175, w__3176;
  wire w__3177, w__3178, w__3179, w__3180, w__3181, w__3182, w__3183, w__3184;
  wire w__3185, w__3186, w__3187, w__3188, w__3189, w__3190, w__3191, w__3192;
  wire w__3193, w__3194, w__3195, w__3196, w__3197, w__3198, w__3199, w__3200;
  wire w__3201, w__3202, w__3203, w__3204, w__3205, w__3206, w__3207, w__3208;
  wire w__3209, w__3210, w__3211, w__3212, w__3213, w__3214, w__3215, w__3216;
  wire w__3217, w__3218, w__3219, w__3220, w__3221, w__3222, w__3223, w__3224;
  wire w__3225, w__3226, w__3227, w__3228, w__3229, w__3230, w__3231, w__3232;
  wire w__3233, w__3234, w__3235, w__3236, w__3237, w__3238, w__3239, w__3240;
  wire w__3241, w__3242, w__3243, w__3244, w__3245, w__3246, w__3247, w__3248;
  wire w__3249, w__3250, w__3251, w__3252, w__3253, w__3254, w__3255, w__3256;
  wire w__3257, w__3258, w__3259, w__3260, w__3261, w__3262, w__3263, w__3264;
  wire w__3265, w__3266, w__3267, w__3268, w__3269, w__3270, w__3271, w__3272;
  wire w__3273, w__3274, w__3275, w__3276, w__3277, w__3278, w__3279, w__3280;
  wire w__3281, w__3282, w__3283, w__3284, w__3285, w__3286, w__3287, w__3288;
  wire w__3289, w__3290, w__3291, w__3292, w__3293, w__3294, w__3295, w__3296;
  wire w__3297, w__3298, w__3299, w__3300, w__3301, w__3302, w__3303, w__3304;
  wire w__3305, w__3306, w__3307, w__3308, w__3309, w__3310, w__3311, w__3312;
  wire w__3313, w__3314, w__3315, w__3316, w__3317, w__3318, w__3319, w__3320;
  wire w__3321, w__3322, w__3323, w__3324, w__3325, w__3326, w__3327, w__3328;
  wire w__3329, w__3330, w__3331, w__3332, w__3333, w__3334, w__3335, w__3336;
  wire w__3337, w__3338, w__3339, w__3340, w__3341, w__3342, w__3343, w__3344;
  wire w__3345, w__3346, w__3347, w__3348, w__3349, w__3350, w__3351, w__3352;
  wire w__3353, w__3354, w__3355, w__3356, w__3357, w__3358, w__3359, w__3360;
  wire w__3361, w__3362, w__3363, w__3364, w__3365, w__3366, w__3367, w__3368;
  wire w__3369, w__3370, w__3371, w__3372, w__3373, w__3374, w__3375, w__3376;
  wire w__3377, w__3378, w__3379, w__3380, w__3381, w__3382, w__3383, w__3384;
  wire w__3385, w__3386, w__3387, w__3388, w__3389, w__3390, w__3391, w__3392;
  wire w__3393, w__3394, w__3395, w__3396, w__3397, w__3398, w__3399, w__3400;
  wire w__3401, w__3402, w__3403, w__3404, w__3405, w__3406, w__3407, w__3408;
  wire w__3409, w__3410, w__3411, w__3412, w__3413, w__3414, w__3415, w__3416;
  wire w__3417, w__3418, w__3419, w__3420, w__3421, w__3422, w__3423, w__3424;
  wire w__3425, w__3426, w__3427, w__3428, w__3429, w__3430, w__3431, w__3432;
  wire w__3433, w__3434, w__3435, w__3436, w__3437, w__3438, w__3439, w__3440;
  wire w__3441, w__3442, w__3443, w__3444, w__3445, w__3446, w__3447, w__3448;
  wire w__3449, w__3450, w__3451, w__3452, w__3453, w__3454, w__3455, w__3456;
  wire w__3457, w__3458, w__3459, w__3460, w__3461, w__3462, w__3463, w__3464;
  wire w__3465, w__3466, w__3467, w__3468, w__3469, w__3470, w__3471, w__3472;
  wire w__3473, w__3474, w__3475, w__3476, w__3477, w__3478, w__3479, w__3480;
  wire w__3481, w__3482, w__3483, w__3484, w__3485, w__3486, w__3487, w__3488;
  wire w__3489, w__3490, w__3491, w__3492, w__3493, w__3494, w__3495, w__3496;
  wire w__3497, w__3498, w__3499, w__3500, w__3501, w__3502, w__3503, w__3504;
  wire w__3505, w__3506, w__3507, w__3508, w__3509, w__3510, w__3511, w__3512;
  wire w__3513, w__3514, w__3515, w__3516, w__3517, w__3518, w__3519, w__3520;
  wire w__3521, w__3522, w__3523, w__3524, w__3525, w__3526, w__3527, w__3528;
  wire w__3529, w__3530, w__3531, w__3532, w__3533, w__3534, w__3535, w__3536;
  wire w__3537, w__3538, w__3539, w__3540, w__3541, w__3542, w__3543, w__3544;
  wire w__3545, w__3546, w__3547, w__3548, w__3549, w__3550, w__3551, w__3552;
  wire w__3553, w__3554, w__3555, w__3556, w__3557, w__3558, w__3559, w__3560;
  wire w__3561, w__3562, w__3563, w__3564, w__3565, w__3566, w__3567, w__3568;
  wire w__3569, w__3570, w__3571, w__3572, w__3573, w__3574, w__3575, w__3576;
  wire w__3577, w__3578, w__3579, w__3580, w__3581, w__3582, w__3583, w__3584;
  wire w__3585, w__3586, w__3587, w__3588, w__3589, w__3590, w__3591, w__3592;
  wire w__3593, w__3594, w__3595, w__3596, w__3597, w__3598, w__3599, w__3600;
  wire w__3601, w__3602, w__3603, w__3604, w__3605, w__3606, w__3607, w__3608;
  wire w__3609, w__3610, w__3611, w__3612, w__3613, w__3614, w__3615, w__3616;
  wire w__3617, w__3618, w__3619, w__3620, w__3621, w__3622, w__3623, w__3624;
  wire w__3625, w__3626, w__3627, w__3628, w__3629, w__3630, w__3631, w__3632;
  wire w__3633, w__3634, w__3635, w__3636, w__3637, w__3638, w__3639, w__3640;
  wire w__3641, w__3642, w__3643, w__3644, w__3645, w__3646, w__3647, w__3648;
  wire w__3649, w__3650, w__3651, w__3652, w__3653, w__3654, w__3655, w__3656;
  wire w__3657, w__3658, w__3659, w__3660, w__3661, w__3662, w__3663, w__3664;
  wire w__3665, w__3666, w__3667, w__3668, w__3669, w__3670, w__3671, w__3672;
  wire w__3673, w__3674, w__3675, w__3676, w__3677, w__3678, w__3679, w__3680;
  wire w__3681, w__3682, w__3683, w__3684, w__3685, w__3686, w__3687, w__3688;
  wire w__3689, w__3690, w__3691, w__3692, w__3693, w__3694, w__3695, w__3696;
  wire w__3697, w__3698, w__3699, w__3700, w__3701, w__3702, w__3703, w__3704;
  wire w__3705, w__3706, w__3707, w__3708, w__3709, w__3710, w__3711, w__3712;
  wire w__3713, w__3714, w__3715, w__3716, w__3717, w__3718, w__3719, w__3720;
  wire w__3721, w__3722, w__3723, w__3724, w__3725, w__3726, w__3727, w__3728;
  wire w__3729, w__3730, w__3731, w__3732, w__3733, w__3734, w__3735, w__3736;
  wire w__3737, w__3738, w__3739, w__3740, w__3741, w__3742, w__3743, w__3744;
  wire w__3745, w__3746, w__3747, w__3748, w__3749, w__3750, w__3751, w__3752;
  wire w__3753, w__3754, w__3755, w__3756, w__3757, w__3758, w__3759, w__3760;
  wire w__3761, w__3762, w__3763, w__3764, w__3765, w__3766, w__3767, w__3768;
  wire w__3769, w__3770, w__3771, w__3772, w__3773, w__3774, w__3775, w__3776;
  wire w__3777, w__3778, w__3779, w__3780, w__3781, w__3782, w__3783, w__3784;
  wire w__3785, w__3786, w__3787, w__3788, w__3789, w__3790, w__3791, w__3792;
  wire w__3793, w__3794, w__3795, w__3796, w__3797, w__3798, w__3799, w__3800;
  wire w__3801, w__3802, w__3803, w__3804, w__3805, w__3806, w__3807, w__3808;
  wire w__3809, w__3810, w__3811, w__3812, w__3813, w__3814, w__3815, w__3816;
  wire w__3817, w__3818, w__3819, w__3820, w__3821, w__3822, w__3823, w__3824;
  wire w__3825, w__3826, w__3827, w__3828, w__3829, w__3830, w__3831, w__3832;
  wire w__3833, w__3834, w__3835, w__3836, w__3837, w__3838, w__3839, w__3840;
  wire w__3841, w__3842, w__3843, w__3844, w__3845, w__3846, w__3847, w__3848;
  wire w__3849, w__3850, w__3851, w__3852, w__3853, w__3854, w__3855, w__3856;
  wire w__3857, w__3858, w__3859, w__3860, w__3861, w__3862, w__3863, w__3864;
  wire w__3865, w__3866, w__3867, w__3868, w__3869, w__3870, w__3871, w__3872;
  wire w__3873, w__3874, w__3875, w__3876, w__3877, w__3878, w__3879, w__3880;
  wire w__3881, w__3882, w__3883, w__3884, w__3885, w__3886, w__3887, w__3888;
  wire w__3889, w__3890, w__3891, w__3892, w__3893, w__3894, w__3895, w__3896;
  wire w__3897, w__3898, w__3899, w__3900, w__3901, w__3902, w__3903, w__3904;
  wire w__3905, w__3906, w__3907, w__3908, w__3909, w__3910, w__3911, w__3912;
  wire w__3913, w__3914, w__3915, w__3916, w__3917, w__3918, w__3919, w__3920;
  wire w__3921, w__3922, w__3923, w__3924, w__3925, w__3926, w__3927, w__3928;
  wire w__3929, w__3930, w__3931, w__3932, w__3933, w__3934, w__3935, w__3936;
  wire w__3937, w__3938, w__3939, w__3940, w__3941, w__3942, w__3943, w__3944;
  wire w__3945, w__3946, w__3947, w__3948, w__3949, w__3950, w__3951, w__3952;
  wire w__3953, w__3954, w__3955, w__3956, w__3957, w__3958, w__3959, w__3960;
  wire w__3961, w__3962, w__3963, w__3964, w__3965, w__3966, w__3967, w__3968;
  wire w__3969, w__3970, w__3971, w__3972, w__3973, w__3974, w__3975, w__3976;
  wire w__3977, w__3978, w__3979, w__3980, w__3981, w__3982, w__3983, w__3984;
  wire w__3985, w__3986, w__3987, w__3988, w__3989, w__3990, w__3991, w__3992;
  wire w__3993, w__3994, w__3995, w__3996, w__3997, w__3998, w__3999, w__4000;
  wire w__4001, w__4002, w__4003, w__4004, w__4005, w__4006, w__4007, w__4008;
  wire w__4009, w__4010, w__4011, w__4012, w__4013, w__4014, w__4015, w__4016;
  wire w__4017, w__4018, w__4019, w__4020, w__4021, w__4022, w__4023, w__4024;
  wire w__4025, w__4026, w__4027, w__4028, w__4029, w__4030, w__4031, w__4032;
  wire w__4033, w__4034, w__4035, w__4036, w__4037, w__4038, w__4039, w__4040;
  wire w__4041, w__4042, w__4043, w__4044, w__4045, w__4046, w__4047, w__4048;
  wire w__4049, w__4050, w__4051, w__4052, w__4053, w__4054, w__4055, w__4056;
  wire w__4057, w__4058, w__4059, w__4060, w__4061, w__4062, w__4063, w__4064;
  wire w__4065, w__4066, w__4067, w__4068, w__4069, w__4070, w__4071, w__4072;
  wire w__4073, w__4074, w__4075, w__4076, w__4077, w__4078, w__4079, w__4080;
  wire w__4081, w__4082, w__4083, w__4084, w__4085, w__4086, w__4087, w__4088;
  wire w__4089, w__4090, w__4091, w__4092, w__4093, w__4094, w__4095, w__4096;
  wire w__4097, w__4098, w__4099, w__4100, w__4101, w__4102, w__4103, w__4104;
  wire w__4105, w__4106, w__4107, w__4108, w__4109, w__4110, w__4111, w__4112;
  wire w__4113, w__4114, w__4115, w__4116, w__4117, w__4118, w__4119, w__4120;
  wire w__4121, w__4122, w__4123, w__4124, w__4125, w__4126, w__4127, w__4128;
  wire w__4129, w__4130, w__4131, w__4132, w__4133, w__4134, w__4135, w__4136;
  wire w__4137, w__4138, w__4139, w__4140, w__4141, w__4142, w__4143, w__4144;
  wire w__4145, w__4146, w__4147, w__4148, w__4149, w__4150, w__4151, w__4152;
  wire w__4153, w__4154, w__4155, w__4156, w__4157, w__4158, w__4159, w__4160;
  wire w__4161, w__4162, w__4163, w__4164, w__4165, w__4166, w__4167, w__4168;
  wire w__4169, w__4170, w__4171, w__4172, w__4173, w__4174, w__4175, w__4176;
  wire w__4177, w__4178, w__4179, w__4180, w__4181, w__4182, w__4183, w__4184;
  wire w__4185, w__4186, w__4187, w__4188, w__4189, w__4190, w__4191, w__4192;
  wire w__4193, w__4194, w__4195, w__4196, w__4197, w__4198, w__4199, w__4200;
  wire w__4201, w__4202, w__4203, w__4204, w__4205, w__4206, w__4207, w__4208;
  wire w__4209, w__4210, w__4211, w__4212, w__4213, w__4214, w__4215, w__4216;
  wire w__4217, w__4218, w__4219, w__4220, w__4221, w__4222, w__4223, w__4224;
  wire w__4225, w__4226, w__4227, w__4228, w__4229, w__4230, w__4231, w__4232;
  wire w__4233, w__4234, w__4235, w__4236, w__4237, w__4238, w__4239, w__4240;
  wire w__4241, w__4242, w__4243, w__4244, w__4245, w__4246, w__4247, w__4248;
  wire w__4249, w__4250, w__4251, w__4252, w__4253, w__4254, w__4255, w__4256;
  wire w__4257, w__4258, w__4259, w__4260, w__4261, w__4262, w__4263, w__4264;
  wire w__4265, w__4266, w__4267, w__4268, w__4269, w__4270, w__4271, w__4272;
  wire w__4273, w__4274, w__4275, w__4276, w__4277, w__4278, w__4279, w__4280;
  wire w__4281, w__4282, w__4283, w__4284, w__4285, w__4286, w__4287, w__4288;
  wire w__4289, w__4290, w__4291, w__4292, w__4293, w__4294, w__4295, w__4296;
  wire w__4297, w__4298, w__4299, w__4300, w__4301, w__4302, w__4303, w__4304;
  wire w__4305, w__4306, w__4307, w__4308, w__4309, w__4310, w__4311, w__4312;
  wire w__4313, w__4314, w__4315, w__4316, w__4317, w__4318, w__4319, w__4320;
  wire w__4321, w__4322, w__4323, w__4324, w__4325, w__4326, w__4327, w__4328;
  wire w__4329, w__4330, w__4331, w__4332, w__4333, w__4334, w__4335, w__4336;
  wire w__4337, w__4338, w__4339, w__4340, w__4341, w__4342, w__4343, w__4344;
  wire w__4345, w__4346, w__4347, w__4348, w__4349, w__4350, w__4351, w__4352;
  wire w__4353, w__4354, w__4355, w__4356, w__4357, w__4358, w__4359, w__4360;
  wire w__4361, w__4362, w__4363, w__4364, w__4365, w__4366, w__4367, w__4368;
  wire w__4369, w__4370, w__4371, w__4372, w__4373, w__4374, w__4375, w__4376;
  wire w__4377, w__4378, w__4379, w__4380, w__4381, w__4382, w__4383, w__4384;
  wire w__4385, w__4386, w__4387, w__4388, w__4389, w__4390, w__4391, w__4392;
  wire w__4393, w__4394, w__4395, w__4396, w__4397, w__4398, w__4399, w__4400;
  wire w__4401, w__4402, w__4403, w__4404, w__4405, w__4406, w__4407, w__4408;
  wire w__4409, w__4410, w__4411, w__4412, w__4413, w__4414, w__4415, w__4416;
  wire w__4417, w__4418, w__4419, w__4420, w__4421, w__4422, w__4423, w__4424;
  wire w__4425, w__4426, w__4427, w__4428, w__4429, w__4430, w__4431, w__4432;
  wire w__4433, w__4434, w__4435, w__4436, w__4437, w__4438, w__4439, w__4440;
  wire w__4441, w__4442, w__4443, w__4444, w__4445, w__4446, w__4447, w__4448;
  wire w__4449, w__4450, w__4451, w__4452, w__4453, w__4454, w__4455, w__4456;
  wire w__4457, w__4458, w__4459, w__4460, w__4461, w__4462, w__4463, w__4464;
  wire w__4465, w__4466, w__4467, w__4468, w__4469, w__4470, w__4471, w__4472;
  wire w__4473, w__4474, w__4475, w__4476, w__4477, w__4478, w__4479, w__4480;
  wire w__4481, w__4482, w__4483, w__4484, w__4485, w__4486, w__4487, w__4488;
  wire w__4489, w__4490, w__4491, w__4492, w__4493, w__4494, w__4495, w__4496;
  wire w__4497, w__4498, w__4499, w__4500, w__4501, w__4502, w__4503, w__4504;
  wire w__4505, w__4506, w__4507, w__4508, w__4509, w__4510, w__4511, w__4512;
  wire w__4513, w__4514, w__4515, w__4516, w__4517, w__4518, w__4519, w__4520;
  wire w__4521, w__4522, w__4523, w__4524, w__4525, w__4526, w__4527, w__4528;
  wire w__4529, w__4530, w__4531, w__4532, w__4533, w__4534, w__4535, w__4536;
  wire w__4537, w__4538, w__4539, w__4540, w__4541, w__4542, w__4543, w__4544;
  wire w__4545, w__4546, w__4547, w__4548, w__4549, w__4550, w__4551, w__4552;
  wire w__4553, w__4554, w__4555, w__4556, w__4557, w__4558, w__4559, w__4560;
  wire w__4561, w__4562, w__4563, w__4564, w__4565, w__4566, w__4567, w__4568;
  wire w__4569, w__4570, w__4571, w__4572, w__4573, w__4574, w__4575, w__4576;
  wire w__4577, w__4578, w__4579, w__4580, w__4581, w__4582, w__4583, w__4584;
  wire w__4585, w__4586, w__4587, w__4588, w__4589, w__4590, w__4591, w__4592;
  wire w__4593, w__4594, w__4595, w__4596, w__4597, w__4598, w__4599, w__4600;
  wire w__4601, w__4602, w__4603, w__4604, w__4605, w__4606, w__4607, w__4608;
  wire w__4609, w__4610, w__4611, w__4612, w__4613, w__4614, w__4615, w__4616;
  wire w__4617, w__4618, w__4619, w__4620, w__4621, w__4622, w__4623, w__4624;
  wire w__4625, w__4626, w__4627, w__4628, w__4629, w__4630, w__4631, w__4632;
  wire w__4633, w__4634, w__4635, w__4636, w__4637, w__4638, w__4639, w__4640;
  wire w__4641, w__4642, w__4643, w__4644, w__4645, w__4646, w__4647, w__4648;
  wire w__4649, w__4650, w__4651, w__4652, w__4653, w__4654, w__4655, w__4656;
  wire w__4657, w__4658, w__4659, w__4660, w__4661, w__4662, w__4663, w__4664;
  wire w__4665, w__4666, w__4667, w__4668, w__4669, w__4670, w__4671, w__4672;
  wire w__4673, w__4674, w__4675, w__4676, w__4677, w__4678, w__4679, w__4680;
  wire w__4681, w__4682, w__4683, w__4684, w__4685, w__4686, w__4687, w__4688;
  wire w__4689, w__4690, w__4691, w__4692, w__4693, w__4694, w__4695, w__4696;
  wire w__4697, w__4698, w__4699, w__4700, w__4701, w__4702, w__4703, w__4704;
  wire w__4705, w__4706, w__4707, w__4708, w__4709, w__4710, w__4711, w__4712;
  wire w__4713, w__4714, w__4715, w__4716, w__4717, w__4718, w__4719, w__4720;
  wire w__4721, w__4722, w__4723, w__4724, w__4725, w__4726, w__4727, w__4728;
  wire w__4729, w__4730, w__4731, w__4732, w__4733, w__4734, w__4735, w__4736;
  wire w__4737, w__4738, w__4739, w__4740, w__4741, w__4742, w__4743, w__4744;
  wire w__4745, w__4746, w__4747, w__4748, w__4749, w__4750, w__4751, w__4752;
  wire w__4753, w__4754, w__4755, w__4756, w__4757, w__4758, w__4759, w__4760;
  wire w__4761, w__4762, w__4763, w__4764, w__4765, w__4766, w__4767, w__4768;
  wire w__4769, w__4770, w__4771, w__4772, w__4773, w__4774, w__4775, w__4776;
  wire w__4777, w__4778, w__4779, w__4780, w__4781, w__4782, w__4783, w__4784;
  wire w__4785, w__4786, w__4787, w__4788, w__4789, w__4790, w__4791, w__4792;
  wire w__4793, w__4794, w__4795, w__4796, w__4797, w__4798, w__4799, w__4800;
  wire w__4801, w__4802, w__4803, w__4804, w__4805, w__4806, w__4807, w__4808;
  wire w__4809, w__4810, w__4811, w__4812, w__4813, w__4814, w__4815, w__4816;
  wire w__4817, w__4818, w__4819;
  buf g__1(w__4198 ,w__4132);
  buf g__2(w__4197 ,w__4131);
  buf g__3(w__4196 ,w__4130);
  buf g__4(w__4179 ,w__4129);
  buf g__5(w__4178 ,w__4127);
  buf g__6(w__4177 ,w__4128);
  buf g__7(w__4176 ,w__4126);
  buf g__8(w__4175 ,w__4125);
  buf g__9(w__4174 ,w__4124);
  buf g__10(w__4173 ,w__4123);
  buf g__11(w__4172 ,w__4122);
  buf g__12(w__4171 ,w__4121);
  buf g__13(w__4170 ,w__4120);
  buf g__14(w__4169 ,w__4119);
  buf g__15(w__4168 ,w__4118);
  buf g__16(w__4167 ,w__4117);
  not g__17(w__4166 ,in22);
  and g__18(w__4102 ,w__4197 ,w__4134);
  and g__19(w__4116 ,w__4167 ,w__4142);
  and g__20(w__4114 ,w__4169 ,w__4143);
  and g__21(w__4110 ,w__4173 ,w__4142);
  and g__22(w__4165 ,w__4198 ,w__4139);
  and g__23(w__4109 ,w__4174 ,w__4140);
  and g__24(w__4113 ,w__4170 ,w__4134);
  and g__25(w__4103 ,w__4196 ,w__4139);
  and g__26(w__4107 ,w__4176 ,w__4136);
  and g__27(w__4115 ,w__4168 ,w__4137);
  and g__28(w__4112 ,w__4171 ,w__4143);
  and g__29(w__4106 ,w__4178 ,w__4136);
  and g__30(w__4105 ,w__4177 ,w__4137);
  and g__31(w__4111 ,w__4172 ,w__4145);
  and g__32(w__4104 ,w__4179 ,w__4140);
  and g__33(w__4108 ,w__4175 ,w__4146);
  not g__34(w__4164 ,w__4162);
  not g__35(w__4163 ,w__4162);
  not g__36(w__4162 ,w__4166);
  buf g__37(w__4101 ,w__4165);
  not g__38(w__4146 ,w__4144);
  not g__39(w__4145 ,w__4144);
  not g__40(w__4144 ,w__4164);
  not g__41(w__4143 ,w__4141);
  not g__42(w__4142 ,w__4141);
  not g__43(w__4141 ,w__4163);
  not g__44(w__4140 ,w__4138);
  not g__45(w__4139 ,w__4138);
  not g__46(w__4138 ,w__4163);
  not g__47(w__4137 ,w__4135);
  not g__48(w__4136 ,w__4135);
  not g__49(w__4135 ,w__4164);
  not g__50(w__4134 ,w__4133);
  not g__51(w__4133 ,w__4146);
  buf g__52(w__4272 ,w__4161);
  buf g__53(w__4271 ,w__4160);
  buf g__54(w__4270 ,w__4159);
  buf g__55(w__4269 ,w__4158);
  buf g__56(w__4268 ,w__4157);
  buf g__57(w__4267 ,w__4156);
  buf g__58(w__4266 ,w__4155);
  buf g__59(w__4265 ,w__4154);
  buf g__60(w__4264 ,w__4153);
  buf g__61(w__4263 ,w__4152);
  buf g__62(w__4262 ,w__4150);
  buf g__63(w__4261 ,w__4149);
  buf g__64(w__4244 ,w__4148);
  buf g__65(w__4243 ,w__4147);
  buf g__66(w__4242 ,w__4151);
  not g__67(w__4241 ,in22);
  and g__68(w__4240 ,w__4272 ,w__4200);
  and g__69(w__4239 ,w__4243 ,w__4208);
  and g__70(w__4238 ,w__4261 ,w__4209);
  and g__71(w__4237 ,w__4264 ,w__4208);
  and g__72(w__4236 ,w__4265 ,w__4206);
  and g__73(w__4097 ,w__4262 ,w__4200);
  and g__74(w__4235 ,w__4271 ,w__4205);
  and g__75(w__4091 ,w__4267 ,w__4202);
  and g__76(w__4099 ,w__4244 ,w__4203);
  and g__77(w__4234 ,w__4242 ,w__4209);
  and g__78(w__4233 ,w__4268 ,w__4202);
  and g__79(w__4089 ,w__4269 ,w__4203);
  and g__80(w__4232 ,w__4263 ,w__4211);
  and g__81(w__4231 ,w__4270 ,w__4206);
  and g__82(w__4092 ,w__4266 ,w__4227);
  not g__83(w__4230 ,w__4228);
  not g__84(w__4229 ,w__4228);
  not g__85(w__4228 ,w__4241);
  buf g__86(w__4096 ,w__4234);
  buf g__87(w__4095 ,w__4232);
  buf g__88(w__4086 ,w__4240);
  buf g__89(w__4094 ,w__4237);
  buf g__90(w__4100 ,w__4239);
  buf g__91(w__4093 ,w__4236);
  buf g__92(w__4090 ,w__4233);
  buf g__93(w__4088 ,w__4231);
  buf g__94(w__4087 ,w__4235);
  buf g__95(w__4098 ,w__4238);
  not g__96(w__4227 ,w__4210);
  not g__97(w__4211 ,w__4210);
  not g__98(w__4210 ,w__4230);
  not g__99(w__4209 ,w__4207);
  not g__100(w__4208 ,w__4207);
  not g__101(w__4207 ,w__4229);
  not g__102(w__4206 ,w__4204);
  not g__103(w__4205 ,w__4204);
  not g__104(w__4204 ,w__4229);
  not g__105(w__4203 ,w__4201);
  not g__106(w__4202 ,w__4201);
  not g__107(w__4201 ,w__4230);
  not g__108(w__4200 ,w__4199);
  not g__109(w__4199 ,w__4227);
  buf g__110(w__4360 ,w__4189);
  buf g__111(w__4359 ,w__4195);
  buf g__112(w__4358 ,w__4194);
  buf g__113(w__4357 ,w__4193);
  buf g__114(w__4341 ,w__4192);
  buf g__115(w__4340 ,w__4191);
  buf g__116(w__4339 ,w__4190);
  buf g__117(w__4338 ,w__4187);
  buf g__118(w__4337 ,w__4188);
  buf g__119(w__4336 ,w__4186);
  buf g__120(w__4335 ,w__4185);
  buf g__121(w__4334 ,w__4184);
  buf g__122(w__4333 ,w__4183);
  buf g__123(w__4332 ,w__4182);
  buf g__124(w__4331 ,w__4181);
  buf g__125(w__4330 ,w__4180);
  not g__126(w__4329 ,in18);
  and g__127(w__4328 ,w__4358 ,w__4274);
  and g__128(w__4085 ,w__4330 ,w__4297);
  and g__129(w__4327 ,w__4332 ,w__4298);
  and g__130(w__4079 ,w__4336 ,w__4297);
  and g__131(w__4326 ,w__4359 ,w__4294);
  and g__132(w__4078 ,w__4338 ,w__4295);
  and g__133(w__4325 ,w__4333 ,w__4274);
  and g__134(w__4072 ,w__4357 ,w__4294);
  and g__135(w__4076 ,w__4360 ,w__4291);
  and g__136(w__4308 ,w__4331 ,w__4292);
  and g__137(w__4081 ,w__4334 ,w__4298);
  and g__138(w__4307 ,w__4339 ,w__4291);
  and g__139(w__4074 ,w__4340 ,w__4292);
  and g__140(w__4306 ,w__4335 ,w__4300);
  and g__141(w__4305 ,w__4341 ,w__4295);
  and g__142(w__4077 ,w__4337 ,w__4301);
  not g__143(w__4304 ,w__4302);
  not g__144(w__4303 ,w__4302);
  not g__145(w__4302 ,w__4329);
  buf g__146(w__4080 ,w__4306);
  buf g__147(w__4070 ,w__4326);
  buf g__148(w__4075 ,w__4307);
  buf g__149(w__4084 ,w__4308);
  buf g__150(w__4082 ,w__4325);
  buf g__151(w__4073 ,w__4305);
  buf g__152(w__4083 ,w__4327);
  buf g__153(w__4071 ,w__4328);
  not g__154(w__4301 ,w__4299);
  not g__155(w__4300 ,w__4299);
  not g__156(w__4299 ,w__4304);
  not g__157(w__4298 ,w__4296);
  not g__158(w__4297 ,w__4296);
  not g__159(w__4296 ,w__4303);
  not g__160(w__4295 ,w__4293);
  not g__161(w__4294 ,w__4293);
  not g__162(w__4293 ,w__4303);
  not g__163(w__4292 ,w__4275);
  not g__164(w__4291 ,w__4275);
  not g__165(w__4275 ,w__4304);
  not g__166(w__4274 ,w__4273);
  not g__167(w__4273 ,w__4301);
  buf g__168(w__4434 ,w__4220);
  buf g__169(w__4433 ,w__4222);
  buf g__170(w__4432 ,w__4221);
  buf g__171(w__4431 ,w__4223);
  buf g__172(w__4430 ,w__4226);
  buf g__173(w__4429 ,w__4225);
  buf g__174(w__4428 ,w__4224);
  buf g__175(w__4427 ,w__4219);
  buf g__176(w__4426 ,w__4218);
  buf g__177(w__4425 ,w__4217);
  buf g__178(w__4424 ,w__4216);
  buf g__179(w__4423 ,w__4215);
  buf g__180(w__4422 ,w__4214);
  buf g__181(w__4406 ,w__4213);
  buf g__182(w__4405 ,w__4212);
  not g__183(w__4404 ,in18);
  and g__184(w__4055 ,w__4430 ,w__4362);
  and g__185(w__4403 ,w__4405 ,w__4370);
  and g__186(w__4067 ,w__4422 ,w__4371);
  and g__187(w__4402 ,w__4426 ,w__4370);
  and g__188(w__4401 ,w__4427 ,w__4368);
  and g__189(w__4066 ,w__4423 ,w__4362);
  and g__190(w__4400 ,w__4429 ,w__4367);
  and g__191(w__4399 ,w__4432 ,w__4364);
  and g__192(w__4398 ,w__4406 ,w__4365);
  and g__193(w__4065 ,w__4424 ,w__4371);
  and g__194(w__4397 ,w__4433 ,w__4364);
  and g__195(w__4396 ,w__4431 ,w__4365);
  and g__196(w__4064 ,w__4425 ,w__4373);
  and g__197(w__4395 ,w__4428 ,w__4368);
  and g__198(w__4394 ,w__4434 ,w__4390);
  not g__199(w__4393 ,w__4391);
  not g__200(w__4392 ,w__4391);
  not g__201(w__4391 ,w__4404);
  buf g__202(w__4062 ,w__4401);
  buf g__203(w__4063 ,w__4402);
  buf g__204(w__4058 ,w__4396);
  buf g__205(w__4059 ,w__4397);
  buf g__206(w__4061 ,w__4394);
  buf g__207(w__4057 ,w__4395);
  buf g__208(w__4068 ,w__4398);
  buf g__209(w__4069 ,w__4403);
  buf g__210(w__4056 ,w__4400);
  buf g__211(w__4060 ,w__4399);
  not g__212(w__4390 ,w__4372);
  not g__213(w__4373 ,w__4372);
  not g__214(w__4372 ,w__4393);
  not g__215(w__4371 ,w__4369);
  not g__216(w__4370 ,w__4369);
  not g__217(w__4369 ,w__4392);
  not g__218(w__4368 ,w__4366);
  not g__219(w__4367 ,w__4366);
  not g__220(w__4366 ,w__4392);
  not g__221(w__4365 ,w__4363);
  not g__222(w__4364 ,w__4363);
  not g__223(w__4363 ,w__4393);
  not g__224(w__4362 ,w__4361);
  not g__225(w__4361 ,w__4390);
  buf g__226(w__4513 ,w__4260);
  buf g__227(w__4512 ,w__4259);
  buf g__228(w__4511 ,w__4258);
  buf g__229(w__4510 ,w__4257);
  buf g__230(w__4509 ,w__4256);
  buf g__231(w__4508 ,w__4255);
  buf g__232(w__4507 ,w__4254);
  buf g__233(w__4506 ,w__4253);
  buf g__234(w__4505 ,w__4252);
  buf g__235(w__4504 ,w__4251);
  buf g__236(w__4503 ,w__4250);
  buf g__237(w__4502 ,w__4249);
  buf g__238(w__4501 ,w__4248);
  buf g__239(w__4500 ,w__4247);
  buf g__240(w__4499 ,w__4246);
  buf g__241(w__4498 ,w__4245);
  not g__242(w__4497 ,in14);
  and g__243(w__4496 ,w__4512 ,w__4436);
  and g__244(w__4495 ,w__4498 ,w__4460);
  and g__245(w__4494 ,w__4500 ,w__4461);
  and g__246(w__4493 ,w__4504 ,w__4460);
  and g__247(w__4492 ,w__4513 ,w__4457);
  and g__248(w__4491 ,w__4505 ,w__4458);
  and g__249(w__4490 ,w__4501 ,w__4436);
  and g__250(w__4489 ,w__4511 ,w__4457);
  and g__251(w__4488 ,w__4507 ,w__4454);
  and g__252(w__4487 ,w__4499 ,w__4455);
  and g__253(w__4486 ,w__4502 ,w__4461);
  and g__254(w__4044 ,w__4508 ,w__4454);
  and g__255(w__4470 ,w__4509 ,w__4455);
  and g__256(w__4469 ,w__4503 ,w__4463);
  and g__257(w__4042 ,w__4510 ,w__4458);
  and g__258(w__4468 ,w__4506 ,w__4464);
  not g__259(w__4467 ,w__4465);
  not g__260(w__4466 ,w__4465);
  not g__261(w__4465 ,w__4497);
  buf g__262(w__4045 ,w__4488);
  buf g__263(w__4039 ,w__4492);
  buf g__264(w__4043 ,w__4470);
  buf g__265(w__4052 ,w__4494);
  buf g__266(w__4053 ,w__4487);
  buf g__267(w__4041 ,w__4489);
  buf g__268(w__4040 ,w__4496);
  buf g__269(w__4054 ,w__4495);
  buf g__270(w__4046 ,w__4468);
  buf g__271(w__4049 ,w__4469);
  buf g__272(w__4048 ,w__4493);
  buf g__273(w__4050 ,w__4486);
  buf g__274(w__4051 ,w__4490);
  buf g__275(w__4047 ,w__4491);
  not g__276(w__4464 ,w__4462);
  not g__277(w__4463 ,w__4462);
  not g__278(w__4462 ,w__4467);
  not g__279(w__4461 ,w__4459);
  not g__280(w__4460 ,w__4459);
  not g__281(w__4459 ,w__4466);
  not g__282(w__4458 ,w__4456);
  not g__283(w__4457 ,w__4456);
  not g__284(w__4456 ,w__4466);
  not g__285(w__4455 ,w__4437);
  not g__286(w__4454 ,w__4437);
  not g__287(w__4437 ,w__4467);
  not g__288(w__4436 ,w__4435);
  not g__289(w__4435 ,w__4464);
  buf g__290(w__4557 ,w__4290);
  buf g__291(w__4556 ,w__4289);
  buf g__292(w__4555 ,w__4288);
  buf g__293(w__4554 ,w__4287);
  buf g__294(w__4553 ,w__4286);
  buf g__295(w__4552 ,w__4285);
  buf g__296(w__4551 ,w__4284);
  buf g__297(w__4550 ,w__4283);
  buf g__298(w__4549 ,w__4282);
  buf g__299(w__4548 ,w__4281);
  buf g__300(w__4547 ,w__4280);
  buf g__301(w__4546 ,w__4279);
  buf g__302(w__4545 ,w__4278);
  buf g__303(w__4544 ,w__4277);
  buf g__304(w__4543 ,w__4276);
  not g__305(w__4542 ,in14);
  and g__306(w__4024 ,w__4557 ,w__4515);
  and g__307(w__4541 ,w__4543 ,w__4523);
  and g__308(w__4540 ,w__4545 ,w__4524);
  and g__309(w__4539 ,w__4549 ,w__4523);
  and g__310(w__4538 ,w__4550 ,w__4521);
  and g__311(w__4537 ,w__4546 ,w__4515);
  and g__312(w__4536 ,w__4556 ,w__4520);
  and g__313(w__4535 ,w__4552 ,w__4517);
  and g__314(w__4534 ,w__4544 ,w__4518);
  and g__315(w__4533 ,w__4547 ,w__4524);
  and g__316(w__4028 ,w__4553 ,w__4517);
  and g__317(w__4532 ,w__4554 ,w__4518);
  and g__318(w__4531 ,w__4548 ,w__4526);
  and g__319(w__4026 ,w__4555 ,w__4521);
  and g__320(w__4030 ,w__4551 ,w__4527);
  not g__321(w__4530 ,w__4528);
  not g__322(w__4529 ,w__4528);
  not g__323(w__4528 ,w__4542);
  buf g__324(w__4031 ,w__4538);
  buf g__325(w__4033 ,w__4531);
  buf g__326(w__4037 ,w__4534);
  buf g__327(w__4038 ,w__4541);
  buf g__328(w__4027 ,w__4532);
  buf g__329(w__4025 ,w__4536);
  buf g__330(w__4032 ,w__4539);
  buf g__331(w__4034 ,w__4533);
  buf g__332(w__4029 ,w__4535);
  buf g__333(w__4035 ,w__4537);
  buf g__334(w__4036 ,w__4540);
  not g__335(w__4527 ,w__4525);
  not g__336(w__4526 ,w__4525);
  not g__337(w__4525 ,w__4530);
  not g__338(w__4524 ,w__4522);
  not g__339(w__4523 ,w__4522);
  not g__340(w__4522 ,w__4529);
  not g__341(w__4521 ,w__4519);
  not g__342(w__4520 ,w__4519);
  not g__343(w__4519 ,w__4529);
  not g__344(w__4518 ,w__4516);
  not g__345(w__4517 ,w__4516);
  not g__346(w__4516 ,w__4530);
  not g__347(w__4515 ,w__4514);
  not g__348(w__4514 ,w__4527);
  buf g__349(w__4607 ,w__4311);
  buf g__350(w__4606 ,w__4324);
  buf g__351(w__4605 ,w__4323);
  buf g__352(w__4604 ,w__4322);
  buf g__353(w__4603 ,w__4321);
  buf g__354(w__4602 ,w__4320);
  buf g__355(w__4601 ,w__4319);
  buf g__356(w__4600 ,w__4318);
  buf g__357(w__4599 ,w__4317);
  buf g__358(w__4598 ,w__4316);
  buf g__359(w__4597 ,w__4315);
  buf g__360(w__4596 ,w__4314);
  buf g__361(w__4595 ,w__4313);
  buf g__362(w__4594 ,w__4312);
  buf g__363(w__4593 ,w__4310);
  buf g__364(w__4592 ,w__4309);
  not g__365(w__4591 ,in10);
  and g__366(w__4590 ,w__4605 ,w__4559);
  and g__367(w__4589 ,w__4592 ,w__4567);
  and g__368(w__4588 ,w__4607 ,w__4568);
  and g__369(w__4587 ,w__4597 ,w__4567);
  and g__370(w__4586 ,w__4606 ,w__4564);
  and g__371(w__4585 ,w__4598 ,w__4565);
  and g__372(w__4584 ,w__4594 ,w__4559);
  and g__373(w__4583 ,w__4604 ,w__4564);
  and g__374(w__4582 ,w__4600 ,w__4561);
  and g__375(w__4581 ,w__4593 ,w__4562);
  and g__376(w__4580 ,w__4595 ,w__4568);
  and g__377(w__4579 ,w__4601 ,w__4561);
  and g__378(w__4578 ,w__4602 ,w__4562);
  and g__379(w__4577 ,w__4596 ,w__4570);
  and g__380(w__4576 ,w__4603 ,w__4565);
  and g__381(w__4575 ,w__4599 ,w__4571);
  not g__382(w__4574 ,w__4572);
  not g__383(w__4573 ,w__4572);
  not g__384(w__4572 ,w__4591);
  buf g__385(w__4017 ,w__4587);
  buf g__386(w__4009 ,w__4590);
  buf g__387(w__4022 ,w__4581);
  buf g__388(w__4023 ,w__4589);
  buf g__389(w__4013 ,w__4579);
  buf g__390(w__4019 ,w__4580);
  buf g__391(w__4015 ,w__4575);
  buf g__392(w__4018 ,w__4577);
  buf g__393(w__4010 ,w__4583);
  buf g__394(w__4021 ,w__4588);
  buf g__395(w__4016 ,w__4585);
  buf g__396(w__4008 ,w__4586);
  buf g__397(w__4014 ,w__4582);
  buf g__398(w__4020 ,w__4584);
  buf g__399(w__4012 ,w__4578);
  buf g__400(w__4011 ,w__4576);
  not g__401(w__4571 ,w__4569);
  not g__402(w__4570 ,w__4569);
  not g__403(w__4569 ,w__4574);
  not g__404(w__4568 ,w__4566);
  not g__405(w__4567 ,w__4566);
  not g__406(w__4566 ,w__4573);
  not g__407(w__4565 ,w__4563);
  not g__408(w__4564 ,w__4563);
  not g__409(w__4563 ,w__4573);
  not g__410(w__4562 ,w__4560);
  not g__411(w__4561 ,w__4560);
  not g__412(w__4560 ,w__4574);
  not g__413(w__4559 ,w__4558);
  not g__414(w__4558 ,w__4571);
  buf g__415(w__4652 ,w__4356);
  buf g__416(w__4651 ,w__4355);
  buf g__417(w__4650 ,w__4354);
  buf g__418(w__4649 ,w__4353);
  buf g__419(w__4648 ,w__4352);
  buf g__420(w__4647 ,w__4351);
  buf g__421(w__4646 ,w__4350);
  buf g__422(w__4645 ,w__4349);
  buf g__423(w__4644 ,w__4348);
  buf g__424(w__4643 ,w__4347);
  buf g__425(w__4642 ,w__4346);
  buf g__426(w__4641 ,w__4345);
  buf g__427(w__4640 ,w__4344);
  buf g__428(w__4639 ,w__4343);
  buf g__429(w__4638 ,w__4342);
  not g__430(w__4637 ,in10);
  and g__431(w__4636 ,w__4652 ,w__4609);
  and g__432(w__4007 ,w__4638 ,w__4617);
  and g__433(w__4635 ,w__4640 ,w__4618);
  and g__434(w__4001 ,w__4644 ,w__4617);
  and g__435(w__4000 ,w__4645 ,w__4615);
  and g__436(w__4634 ,w__4641 ,w__4609);
  and g__437(w__4633 ,w__4651 ,w__4614);
  and g__438(w__4632 ,w__4647 ,w__4611);
  and g__439(w__4631 ,w__4639 ,w__4612);
  and g__440(w__4630 ,w__4642 ,w__4618);
  and g__441(w__4629 ,w__4648 ,w__4611);
  and g__442(w__4628 ,w__4649 ,w__4612);
  and g__443(w__4627 ,w__4643 ,w__4620);
  and g__444(w__4626 ,w__4650 ,w__4615);
  and g__445(w__4625 ,w__4646 ,w__4621);
  not g__446(w__4624 ,w__4622);
  not g__447(w__4623 ,w__4622);
  not g__448(w__4622 ,w__4637);
  buf g__449(w__4002 ,w__4627);
  buf g__450(w__3994 ,w__4633);
  buf g__451(w__3995 ,w__4626);
  buf g__452(w__3996 ,w__4628);
  buf g__453(w__3997 ,w__4629);
  buf g__454(w__4003 ,w__4630);
  buf g__455(w__4006 ,w__4631);
  buf g__456(w__4005 ,w__4635);
  buf g__457(w__3999 ,w__4625);
  buf g__458(w__4004 ,w__4634);
  buf g__459(w__3993 ,w__4636);
  buf g__460(w__3998 ,w__4632);
  not g__461(w__4621 ,w__4619);
  not g__462(w__4620 ,w__4619);
  not g__463(w__4619 ,w__4624);
  not g__464(w__4618 ,w__4616);
  not g__465(w__4617 ,w__4616);
  not g__466(w__4616 ,w__4623);
  not g__467(w__4615 ,w__4613);
  not g__468(w__4614 ,w__4613);
  not g__469(w__4613 ,w__4623);
  not g__470(w__4612 ,w__4610);
  not g__471(w__4611 ,w__4610);
  not g__472(w__4610 ,w__4624);
  not g__473(w__4609 ,w__4608);
  not g__474(w__4608 ,w__4621);
  buf g__475(w__4694 ,w__4389);
  buf g__476(w__4693 ,w__4388);
  buf g__477(w__4692 ,w__4387);
  buf g__478(w__4691 ,w__4386);
  buf g__479(w__4690 ,w__4385);
  buf g__480(w__4689 ,w__4384);
  buf g__481(w__4688 ,w__4383);
  buf g__482(w__4687 ,w__4382);
  buf g__483(w__4686 ,w__4381);
  buf g__484(w__4685 ,w__4380);
  buf g__485(w__4684 ,w__4378);
  buf g__486(w__4683 ,w__4376);
  buf g__487(w__4682 ,w__4375);
  buf g__488(w__4681 ,w__4374);
  buf g__489(w__4680 ,w__4377);
  buf g__490(w__4679 ,w__4379);
  not g__491(w__4678 ,in3);
  and g__492(w__4677 ,w__4693 ,w__4654);
  and g__493(w__3992 ,w__4681 ,w__4662);
  and g__494(w__3990 ,w__4683 ,w__4663);
  and g__495(w__3986 ,w__4685 ,w__4662);
  and g__496(w__4676 ,w__4694 ,w__4659);
  and g__497(w__3985 ,w__4686 ,w__4660);
  and g__498(w__3989 ,w__4680 ,w__4654);
  and g__499(w__3979 ,w__4692 ,w__4659);
  and g__500(w__4675 ,w__4688 ,w__4656);
  and g__501(w__3991 ,w__4682 ,w__4657);
  and g__502(w__4674 ,w__4684 ,w__4663);
  and g__503(w__4673 ,w__4689 ,w__4656);
  and g__504(w__4672 ,w__4690 ,w__4657);
  and g__505(w__4671 ,w__4679 ,w__4665);
  and g__506(w__4670 ,w__4691 ,w__4660);
  and g__507(w__3984 ,w__4687 ,w__4666);
  not g__508(w__4669 ,w__4667);
  not g__509(w__4668 ,w__4667);
  not g__510(w__4667 ,w__4678);
  buf g__511(w__3988 ,w__4674);
  buf g__512(w__3980 ,w__4670);
  buf g__513(w__3981 ,w__4672);
  buf g__514(w__3987 ,w__4671);
  buf g__515(w__3983 ,w__4675);
  buf g__516(w__3982 ,w__4673);
  buf g__517(w__3978 ,w__4677);
  buf g__518(w__3977 ,w__4676);
  not g__519(w__4666 ,w__4664);
  not g__520(w__4665 ,w__4664);
  not g__521(w__4664 ,w__4669);
  not g__522(w__4663 ,w__4661);
  not g__523(w__4662 ,w__4661);
  not g__524(w__4661 ,w__4668);
  not g__525(w__4660 ,w__4658);
  not g__526(w__4659 ,w__4658);
  not g__527(w__4658 ,w__4668);
  not g__528(w__4657 ,w__4655);
  not g__529(w__4656 ,w__4655);
  not g__530(w__4655 ,w__4669);
  not g__531(w__4654 ,w__4653);
  not g__532(w__4653 ,w__4666);
  buf g__533(w__4736 ,w__4421);
  buf g__534(w__4735 ,w__4420);
  buf g__535(w__4734 ,w__4419);
  buf g__536(w__4733 ,w__4418);
  buf g__537(w__4732 ,w__4417);
  buf g__538(w__4731 ,w__4416);
  buf g__539(w__4730 ,w__4415);
  buf g__540(w__4729 ,w__4414);
  buf g__541(w__4728 ,w__4413);
  buf g__542(w__4727 ,w__4412);
  buf g__543(w__4726 ,w__4411);
  buf g__544(w__4725 ,w__4410);
  buf g__545(w__4724 ,w__4409);
  buf g__546(w__4723 ,w__4408);
  buf g__547(w__4722 ,w__4407);
  not g__548(w__4721 ,in3);
  and g__549(w__3962 ,w__4736 ,w__4696);
  and g__550(w__4720 ,w__4722 ,w__4704);
  and g__551(w__3974 ,w__4724 ,w__4705);
  and g__552(w__4719 ,w__4728 ,w__4704);
  and g__553(w__4718 ,w__4729 ,w__4702);
  and g__554(w__4717 ,w__4725 ,w__4696);
  and g__555(w__4716 ,w__4735 ,w__4701);
  and g__556(w__4715 ,w__4731 ,w__4698);
  and g__557(w__4714 ,w__4723 ,w__4699);
  and g__558(w__3972 ,w__4726 ,w__4705);
  and g__559(w__3966 ,w__4732 ,w__4698);
  and g__560(w__4713 ,w__4733 ,w__4699);
  and g__561(w__3971 ,w__4727 ,w__4707);
  and g__562(w__3964 ,w__4734 ,w__4702);
  and g__563(w__4712 ,w__4730 ,w__4708);
  not g__564(w__4711 ,w__4709);
  not g__565(w__4710 ,w__4709);
  not g__566(w__4709 ,w__4721);
  buf g__567(w__3970 ,w__4719);
  buf g__568(w__3965 ,w__4713);
  buf g__569(w__3975 ,w__4714);
  buf g__570(w__3967 ,w__4715);
  buf g__571(w__3976 ,w__4720);
  buf g__572(w__3973 ,w__4717);
  buf g__573(w__3969 ,w__4718);
  buf g__574(w__3968 ,w__4712);
  buf g__575(w__3963 ,w__4716);
  not g__576(w__4708 ,w__4706);
  not g__577(w__4707 ,w__4706);
  not g__578(w__4706 ,w__4711);
  not g__579(w__4705 ,w__4703);
  not g__580(w__4704 ,w__4703);
  not g__581(w__4703 ,w__4710);
  not g__582(w__4702 ,w__4700);
  not g__583(w__4701 ,w__4700);
  not g__584(w__4700 ,w__4710);
  not g__585(w__4699 ,w__4697);
  not g__586(w__4698 ,w__4697);
  not g__587(w__4697 ,w__4711);
  not g__588(w__4696 ,w__4695);
  not g__589(w__4695 ,w__4708);
  buf g__590(w__4780 ,w__4441);
  buf g__591(w__4779 ,w__4453);
  buf g__592(w__4778 ,w__4452);
  buf g__593(w__4777 ,w__4450);
  buf g__594(w__4776 ,w__4449);
  buf g__595(w__4775 ,w__4448);
  buf g__596(w__4774 ,w__4447);
  buf g__597(w__4773 ,w__4446);
  buf g__598(w__4772 ,w__4445);
  buf g__599(w__4771 ,w__4444);
  buf g__600(w__4770 ,w__4443);
  buf g__601(w__4769 ,w__4442);
  buf g__602(w__4768 ,w__4440);
  buf g__603(w__4767 ,w__4439);
  buf g__604(w__4766 ,w__4438);
  buf g__605(w__4765 ,w__4451);
  not g__606(w__4764 ,in6);
  and g__607(w__4763 ,w__4778 ,w__4738);
  and g__608(w__4762 ,w__4766 ,w__4746);
  and g__609(w__3959 ,w__4768 ,w__4747);
  and g__610(w__4761 ,w__4771 ,w__4746);
  and g__611(w__3946 ,w__4779 ,w__4743);
  and g__612(w__4760 ,w__4772 ,w__4744);
  and g__613(w__3958 ,w__4780 ,w__4738);
  and g__614(w__4759 ,w__4765 ,w__4743);
  and g__615(w__4758 ,w__4774 ,w__4740);
  and g__616(w__3960 ,w__4767 ,w__4741);
  and g__617(w__3957 ,w__4769 ,w__4747);
  and g__618(w__4757 ,w__4775 ,w__4740);
  and g__619(w__4756 ,w__4776 ,w__4741);
  and g__620(w__3956 ,w__4770 ,w__4749);
  and g__621(w__4755 ,w__4777 ,w__4744);
  and g__622(w__4754 ,w__4773 ,w__4750);
  not g__623(w__4753 ,w__4751);
  not g__624(w__4752 ,w__4751);
  not g__625(w__4751 ,w__4764);
  buf g__626(w__3954 ,w__4760);
  buf g__627(w__3949 ,w__4755);
  buf g__628(w__3950 ,w__4756);
  buf g__629(w__3951 ,w__4757);
  buf g__630(w__3952 ,w__4758);
  buf g__631(w__3948 ,w__4759);
  buf g__632(w__3947 ,w__4763);
  buf g__633(w__3955 ,w__4761);
  buf g__634(w__3961 ,w__4762);
  buf g__635(w__3953 ,w__4754);
  not g__636(w__4750 ,w__4748);
  not g__637(w__4749 ,w__4748);
  not g__638(w__4748 ,w__4753);
  not g__639(w__4747 ,w__4745);
  not g__640(w__4746 ,w__4745);
  not g__641(w__4745 ,w__4752);
  not g__642(w__4744 ,w__4742);
  not g__643(w__4743 ,w__4742);
  not g__644(w__4742 ,w__4752);
  not g__645(w__4741 ,w__4739);
  not g__646(w__4740 ,w__4739);
  not g__647(w__4739 ,w__4753);
  not g__648(w__4738 ,w__4737);
  not g__649(w__4737 ,w__4750);
  buf g__650(w__4819 ,w__4474);
  buf g__651(w__4818 ,w__4485);
  buf g__652(w__4817 ,w__4484);
  buf g__653(w__4816 ,w__4483);
  buf g__654(w__4815 ,w__4482);
  buf g__655(w__4814 ,w__4481);
  buf g__656(w__4813 ,w__4480);
  buf g__657(w__4812 ,w__4479);
  buf g__658(w__4811 ,w__4478);
  buf g__659(w__4810 ,w__4477);
  buf g__660(w__4809 ,w__4476);
  buf g__661(w__4808 ,w__4475);
  buf g__662(w__4807 ,w__4473);
  buf g__663(w__4806 ,w__4472);
  buf g__664(w__4805 ,w__4471);
  not g__665(w__4804 ,in6);
  and g__666(w__4803 ,w__4818 ,w__4782);
  and g__667(w__4802 ,w__4805 ,w__4790);
  and g__668(w__3943 ,w__4807 ,w__4791);
  and g__669(w__3939 ,w__4810 ,w__4790);
  and g__670(w__3938 ,w__4811 ,w__4788);
  and g__671(w__3942 ,w__4819 ,w__4782);
  and g__672(w__3932 ,w__4817 ,w__4787);
  and g__673(w__3936 ,w__4813 ,w__4784);
  and g__674(w__4801 ,w__4806 ,w__4785);
  and g__675(w__3941 ,w__4808 ,w__4791);
  and g__676(w__4800 ,w__4814 ,w__4784);
  and g__677(w__3934 ,w__4815 ,w__4785);
  and g__678(w__3940 ,w__4809 ,w__4793);
  and g__679(w__4799 ,w__4816 ,w__4788);
  and g__680(w__4798 ,w__4812 ,w__4794);
  not g__681(w__4797 ,w__4795);
  not g__682(w__4796 ,w__4795);
  not g__683(w__4795 ,w__4804);
  buf g__684(w__3933 ,w__4799);
  buf g__685(w__3945 ,w__4802);
  buf g__686(w__3944 ,w__4801);
  buf g__687(w__3937 ,w__4798);
  buf g__688(w__3931 ,w__4803);
  buf g__689(w__3935 ,w__4800);
  not g__690(w__4794 ,w__4792);
  not g__691(w__4793 ,w__4792);
  not g__692(w__4792 ,w__4797);
  not g__693(w__4791 ,w__4789);
  not g__694(w__4790 ,w__4789);
  not g__695(w__4789 ,w__4796);
  not g__696(w__4788 ,w__4786);
  not g__697(w__4787 ,w__4786);
  not g__698(w__4786 ,w__4796);
  not g__699(w__4785 ,w__4783);
  not g__700(w__4784 ,w__4783);
  not g__701(w__4783 ,w__4797);
  not g__702(w__4782 ,w__4781);
  not g__703(w__4781 ,w__4794);
  xnor g__704(out1[16] ,w__1182 ,w__1155);
  nor g__705(w__1182 ,w__1181 ,w__1131);
  xnor g__706(out1[15] ,w__1180 ,w__1156);
  and g__707(w__1181 ,w__1136 ,w__1180);
  or g__708(w__1180 ,w__1134 ,w__1179);
  xnor g__709(out1[14] ,w__1178 ,w__1153);
  nor g__710(w__1179 ,w__1178 ,w__1137);
  and g__711(w__1178 ,w__1138 ,w__1177);
  xnor g__712(out1[13] ,w__1175 ,w__1154);
  or g__713(w__1177 ,w__1132 ,w__1176);
  not g__714(w__1176 ,w__1175);
  or g__715(w__1175 ,w__1145 ,w__1174);
  xnor g__716(out1[12] ,w__1173 ,w__1148);
  nor g__717(w__1174 ,w__1173 ,w__1140);
  and g__718(w__1173 ,w__1123 ,w__1172);
  xnor g__719(out1[11] ,w__1170 ,w__1128);
  or g__720(w__1172 ,w__1121 ,w__1171);
  not g__721(w__1171 ,w__1170);
  or g__722(w__1170 ,w__1139 ,w__1169);
  xnor g__723(out1[10] ,w__1168 ,w__1152);
  nor g__724(w__1169 ,w__1168 ,w__1141);
  and g__725(w__1168 ,w__1147 ,w__1167);
  xnor g__726(out1[9] ,w__1166 ,w__1151);
  or g__727(w__1167 ,w__1146 ,w__1166);
  and g__728(w__1166 ,w__1165 ,w__1122);
  or g__729(w__1165 ,w__1124 ,w__1164);
  and g__730(w__1164 ,w__1144 ,w__1163);
  xnor g__731(out1[7] ,w__1161 ,w__1150);
  or g__732(w__1163 ,w__1143 ,w__1162);
  not g__733(w__1162 ,w__1161);
  or g__734(w__1161 ,w__1160 ,w__1133);
  xnor g__735(out1[6] ,w__1159 ,w__1149);
  and g__736(w__1160 ,w__1135 ,w__1159);
  or g__737(w__1159 ,w__1120 ,w__1158);
  xnor g__738(out1[5] ,w__1157 ,w__1130);
  and g__739(w__1158 ,w__1119 ,w__1157);
  xnor g__740(w__1156 ,w__1102 ,w__1118);
  xnor g__741(w__1155 ,w__1082 ,w__1108);
  xnor g__742(w__1154 ,w__1104 ,w__1117);
  xnor g__743(w__1153 ,w__1085 ,w__1109);
  or g__744(w__1157 ,w__1084 ,w__1142);
  xnor g__745(out1[4] ,w__1127 ,w__1107);
  xnor g__746(w__1152 ,w__1096 ,w__1125);
  xnor g__747(w__1151 ,w__1095 ,w__1112);
  xnor g__748(w__1150 ,w__1113 ,w__1126);
  xnor g__749(w__1149 ,w__1086 ,w__1115);
  xnor g__750(w__1148 ,w__1105 ,w__1114);
  or g__751(w__1147 ,w__1094 ,w__1112);
  nor g__752(w__1146 ,w__1095 ,w__1111);
  nor g__753(w__1145 ,w__1106 ,w__1114);
  or g__754(w__1144 ,w__1126 ,w__1113);
  and g__755(w__1143 ,w__1126 ,w__1113);
  and g__756(w__1142 ,w__1083 ,w__1127);
  and g__757(w__1141 ,w__1097 ,w__1125);
  and g__758(w__1140 ,w__1106 ,w__1114);
  nor g__759(w__1139 ,w__1097 ,w__1125);
  or g__760(w__1138 ,w__1103 ,w__1116);
  and g__761(w__1137 ,w__1085 ,w__1110);
  or g__762(w__1136 ,w__1102 ,w__1118);
  or g__763(w__1135 ,w__1086 ,w__1115);
  nor g__764(w__1134 ,w__1085 ,w__1110);
  and g__765(w__1133 ,w__1086 ,w__1115);
  nor g__766(w__1132 ,w__1104 ,w__1117);
  and g__767(w__1131 ,w__1102 ,w__1118);
  xnor g__768(out1[3] ,w__1080 ,w__1081);
  xnor g__769(w__1130 ,w__1079 ,w__1089);
  xnor g__770(w__1129 ,w__1099 ,w__1088);
  xnor g__771(w__1128 ,w__1101 ,w__1091);
  nor g__772(w__1124 ,w__1099 ,w__1088);
  or g__773(w__1123 ,w__1100 ,w__1090);
  or g__774(w__1122 ,w__1098 ,w__1087);
  nor g__775(w__1121 ,w__1101 ,w__1091);
  and g__776(w__1120 ,w__1079 ,w__1089);
  or g__777(w__1119 ,w__1079 ,w__1089);
  or g__778(w__1127 ,w__1071 ,w__1092);
  and g__779(w__1126 ,w__1076 ,w__1093);
  xnor g__780(w__1125 ,w__997 ,w__1059);
  not g__781(w__1117 ,w__1116);
  not g__782(w__1112 ,w__1111);
  not g__783(w__1110 ,w__1109);
  xnor g__784(w__1108 ,w__1016 ,w__1057);
  xnor g__785(w__1107 ,w__1020 ,w__1067);
  xnor g__786(w__1118 ,w__1019 ,w__1062);
  xnor g__787(w__1116 ,w__988 ,w__1061);
  xnor g__788(w__1115 ,w__1039 ,w__1060);
  xnor g__789(w__1114 ,w__996 ,w__1058);
  xnor g__790(w__1113 ,w__1004 ,w__1056);
  xnor g__791(w__1111 ,w__1027 ,w__1063);
  xnor g__792(w__1109 ,w__1018 ,w__1055);
  not g__793(w__1106 ,w__1105);
  not g__794(w__1103 ,w__1104);
  not g__795(w__1100 ,w__1101);
  not g__796(w__1098 ,w__1099);
  not g__797(w__1097 ,w__1096);
  not g__798(w__1094 ,w__1095);
  or g__799(w__1093 ,w__1025 ,w__1074);
  and g__800(w__1092 ,w__1069 ,w__1080);
  or g__801(w__1105 ,w__1031 ,w__1075);
  or g__802(w__1104 ,w__1054 ,w__1072);
  or g__803(w__1102 ,w__1045 ,w__1073);
  or g__804(w__1101 ,w__1047 ,w__1070);
  or g__805(w__1099 ,w__1051 ,w__1077);
  or g__806(w__1096 ,w__1043 ,w__1068);
  or g__807(w__1095 ,w__1053 ,w__1078);
  not g__808(w__1091 ,w__1090);
  not g__809(w__1087 ,w__1088);
  and g__810(w__1084 ,w__1020 ,w__1067);
  or g__811(w__1083 ,w__1020 ,w__1067);
  nor g__812(w__1082 ,w__1033 ,w__1066);
  xnor g__813(w__1081 ,w__978 ,w__1040);
  xnor g__814(w__1090 ,w__1007 ,w__1028);
  xnor g__815(w__1089 ,w__1010 ,w__1029);
  xnor g__816(w__1088 ,w__1021 ,w__1030);
  or g__817(w__1086 ,w__1037 ,w__1064);
  and g__818(w__1085 ,w__1035 ,w__1065);
  nor g__819(w__1078 ,w__998 ,w__1052);
  and g__820(w__1077 ,w__1024 ,w__1050);
  or g__821(w__1076 ,w__909 ,w__1039);
  and g__822(w__1075 ,w__995 ,w__1034);
  and g__823(w__1074 ,w__909 ,w__1039);
  nor g__824(w__1073 ,w__1049 ,w__1014);
  and g__825(w__1072 ,w__996 ,w__1038);
  and g__826(w__1071 ,w__978 ,w__1040);
  and g__827(w__1070 ,w__997 ,w__1044);
  or g__828(w__1069 ,w__978 ,w__1040);
  and g__829(w__1068 ,w__1027 ,w__1041);
  or g__830(w__1080 ,w__991 ,w__1046);
  or g__831(w__1079 ,w__966 ,w__1048);
  xor g__832(out1[2] ,w__1026 ,w__1017);
  nor g__833(w__1066 ,w__1013 ,w__1032);
  or g__834(w__1065 ,w__989 ,w__1042);
  nor g__835(w__1064 ,w__999 ,w__1036);
  xnor g__836(w__1063 ,w__903 ,w__1005);
  xnor g__837(w__1062 ,w__1011 ,w__1012);
  xnor g__838(w__1061 ,w__900 ,w__1009);
  xor g__839(w__1060 ,w__1025 ,w__909);
  xnor g__840(w__1059 ,w__895 ,w__1023);
  xnor g__841(w__1058 ,w__902 ,w__1002);
  xnor g__842(w__1057 ,w__937 ,w__1000);
  xnor g__843(w__1056 ,w__951 ,w__1024);
  xor g__844(w__1055 ,w__1014 ,w__929);
  xnor g__845(w__1067 ,w__1015 ,w__982);
  nor g__846(w__1054 ,w__902 ,w__1001);
  and g__847(w__1053 ,w__952 ,w__1021);
  nor g__848(w__1052 ,w__952 ,w__1021);
  nor g__849(w__1051 ,w__950 ,w__1004);
  or g__850(w__1050 ,w__951 ,w__1003);
  nor g__851(w__1049 ,w__929 ,w__1018);
  nor g__852(w__1048 ,w__965 ,w__1015);
  nor g__853(w__1047 ,w__895 ,w__1022);
  and g__854(w__1046 ,w__1026 ,w__987);
  and g__855(w__1045 ,w__929 ,w__1018);
  or g__856(w__1044 ,w__894 ,w__1023);
  and g__857(w__1043 ,w__903 ,w__1005);
  nor g__858(w__1042 ,w__899 ,w__1009);
  or g__859(w__1041 ,w__903 ,w__1005);
  or g__860(w__1038 ,w__901 ,w__1002);
  and g__861(w__1037 ,w__898 ,w__1010);
  nor g__862(w__1036 ,w__898 ,w__1010);
  or g__863(w__1035 ,w__900 ,w__1008);
  or g__864(w__1034 ,w__878 ,w__1006);
  nor g__865(w__1033 ,w__1011 ,w__1019);
  and g__866(w__1032 ,w__1011 ,w__1019);
  xnor g__867(out1[1] ,w__880 ,w__979);
  nor g__868(w__1031 ,w__877 ,w__1007);
  xor g__869(w__1030 ,w__952 ,w__998);
  xnor g__870(w__1029 ,w__999 ,w__897);
  xnor g__871(w__1028 ,w__878 ,w__995);
  xnor g__872(w__1040 ,w__957 ,w__980);
  xnor g__873(w__1039 ,w__884 ,w__981);
  not g__874(w__1022 ,w__1023);
  xnor g__875(w__1017 ,w__906 ,w__954);
  nor g__876(w__1016 ,w__958 ,w__986);
  or g__877(w__1027 ,w__888 ,w__984);
  or g__878(w__1026 ,w__960 ,w__990);
  and g__879(w__1025 ,w__970 ,w__993);
  or g__880(w__1024 ,w__975 ,w__992);
  xnor g__881(w__1023 ,w__885 ,w__949);
  xnor g__882(w__1021 ,w__955 ,w__945);
  or g__883(w__1020 ,w__964 ,w__985);
  and g__884(w__1019 ,w__974 ,w__983);
  or g__885(w__1018 ,w__918 ,w__994);
  not g__886(w__1013 ,w__1012);
  not g__887(w__1009 ,w__1008);
  not g__888(w__1007 ,w__1006);
  not g__889(w__1003 ,w__1004);
  not g__890(w__1002 ,w__1001);
  xnor g__891(w__1000 ,w__939 ,w__935);
  xnor g__892(w__1015 ,w__856 ,w__944);
  xnor g__893(w__1014 ,w__893 ,w__943);
  xnor g__894(w__1012 ,w__928 ,w__940);
  xnor g__895(w__1011 ,w__788 ,w__947);
  xnor g__896(w__1010 ,w__908 ,w__941);
  xnor g__897(w__1008 ,w__956 ,w__936);
  xnor g__898(w__1006 ,w__912 ,w__948);
  xnor g__899(w__1005 ,w__913 ,w__938);
  xnor g__900(w__1004 ,w__933 ,w__946);
  xnor g__901(w__1001 ,w__932 ,w__942);
  and g__902(w__994 ,w__921 ,w__956);
  or g__903(w__993 ,w__881 ,w__969);
  and g__904(w__992 ,w__884 ,w__971);
  nor g__905(w__991 ,w__905 ,w__954);
  and g__906(w__990 ,w__880 ,w__959);
  and g__907(w__999 ,w__916 ,w__968);
  and g__908(w__998 ,w__922 ,w__962);
  or g__909(w__997 ,w__889 ,w__961);
  or g__910(w__996 ,w__919 ,w__972);
  or g__911(w__995 ,w__917 ,w__967);
  not g__912(w__989 ,w__988);
  or g__913(w__987 ,w__906 ,w__953);
  nor g__914(w__986 ,w__886 ,w__977);
  nor g__915(w__985 ,w__963 ,w__957);
  and g__916(w__984 ,w__955 ,w__923);
  or g__917(w__983 ,w__865 ,w__973);
  xnor g__918(w__982 ,w__930 ,w__896);
  xnor g__919(w__981 ,w__841 ,w__911);
  xnor g__920(w__980 ,w__875 ,w__892);
  xnor g__921(w__979 ,w__735 ,w__904);
  or g__922(w__988 ,w__891 ,w__976);
  nor g__923(w__977 ,w__853 ,w__928);
  and g__924(w__976 ,w__926 ,w__932);
  nor g__925(w__975 ,w__841 ,w__910);
  or g__926(w__974 ,w__843 ,w__893);
  and g__927(w__973 ,w__843 ,w__893);
  and g__928(w__972 ,w__927 ,w__912);
  or g__929(w__971 ,w__840 ,w__911);
  or g__930(w__970 ,w__754 ,w__907);
  nor g__931(w__969 ,w__753 ,w__908);
  or g__932(w__968 ,w__883 ,w__915);
  and g__933(w__967 ,w__914 ,w__885);
  nor g__934(w__966 ,w__931 ,w__896);
  and g__935(w__965 ,w__931 ,w__896);
  nor g__936(w__964 ,w__876 ,w__892);
  and g__937(w__963 ,w__876 ,w__892);
  or g__938(w__962 ,w__934 ,w__920);
  and g__939(w__961 ,w__890 ,w__913);
  and g__940(w__960 ,w__735 ,w__904);
  or g__941(w__959 ,w__735 ,w__904);
  and g__942(w__958 ,w__853 ,w__928);
  or g__943(w__978 ,w__813 ,w__887);
  not g__944(w__953 ,w__954);
  not g__945(w__950 ,w__951);
  xnor g__946(out1[0] ,w__491 ,w__847);
  xnor g__947(w__949 ,w__842 ,w__859);
  xnor g__948(w__948 ,w__839 ,w__864);
  xnor g__949(w__947 ,w__706 ,w__866);
  xnor g__950(w__946 ,w__751 ,w__858);
  xnor g__951(w__945 ,w__818 ,w__862);
  xnor g__952(w__944 ,w__883 ,w__748);
  xnor g__953(w__943 ,w__865 ,w__843);
  xnor g__954(w__942 ,w__817 ,w__860);
  xnor g__955(w__941 ,w__881 ,w__754);
  xor g__956(w__940 ,w__886 ,w__853);
  or g__957(w__939 ,w__814 ,w__924);
  xnor g__958(w__938 ,w__741 ,w__863);
  xnor g__959(w__937 ,w__629 ,w__848);
  xnor g__960(w__936 ,w__845 ,w__855);
  xnor g__961(w__935 ,w__867 ,w__849);
  xnor g__962(w__957 ,w__747 ,w__852);
  xnor g__963(w__956 ,w__756 ,w__850);
  or g__964(w__955 ,w__779 ,w__925);
  xnor g__965(w__954 ,w__882 ,w__851);
  xnor g__966(w__952 ,w__740 ,w__846);
  xnor g__967(w__951 ,w__879 ,w__799);
  not g__968(w__934 ,w__933);
  not g__969(w__931 ,w__930);
  or g__970(w__927 ,w__839 ,w__864);
  or g__971(w__926 ,w__817 ,w__861);
  and g__972(w__925 ,w__787 ,w__879);
  and g__973(w__924 ,w__831 ,w__866);
  or g__974(w__923 ,w__818 ,w__862);
  or g__975(w__922 ,w__750 ,w__858);
  or g__976(w__921 ,w__845 ,w__854);
  nor g__977(w__920 ,w__751 ,w__857);
  and g__978(w__919 ,w__839 ,w__864);
  nor g__979(w__918 ,w__844 ,w__855);
  and g__980(w__917 ,w__842 ,w__859);
  or g__981(w__916 ,w__748 ,w__856);
  and g__982(w__915 ,w__748 ,w__856);
  or g__983(w__914 ,w__842 ,w__859);
  or g__984(w__933 ,w__834 ,w__871);
  or g__985(w__932 ,w__837 ,w__873);
  or g__986(w__930 ,w__824 ,w__868);
  or g__987(w__929 ,w__829 ,w__872);
  or g__988(w__928 ,w__822 ,w__874);
  not g__989(w__910 ,w__911);
  not g__990(w__907 ,w__908);
  not g__991(w__905 ,w__906);
  not g__992(w__902 ,w__901);
  not g__993(w__900 ,w__899);
  not g__994(w__898 ,w__897);
  not g__995(w__895 ,w__894);
  and g__996(w__891 ,w__817 ,w__861);
  or g__997(w__890 ,w__741 ,w__863);
  and g__998(w__889 ,w__741 ,w__863);
  and g__999(w__888 ,w__818 ,w__862);
  and g__1000(w__887 ,w__812 ,w__882);
  or g__1001(w__913 ,w__827 ,w__870);
  xnor g__1002(w__912 ,w__752 ,w__803);
  xnor g__1003(w__911 ,w__687 ,w__798);
  xor g__1004(w__909 ,w__749 ,w__797);
  xnor g__1005(w__908 ,w__793 ,w__796);
  xnor g__1006(w__906 ,w__691 ,w__807);
  xnor g__1007(w__904 ,w__674 ,w__794);
  xnor g__1008(w__903 ,w__791 ,w__806);
  xnor g__1009(w__901 ,w__744 ,w__804);
  or g__1010(w__899 ,w__815 ,w__869);
  xnor g__1011(w__897 ,w__651 ,w__802);
  xnor g__1012(w__896 ,w__681 ,w__801);
  xnor g__1013(w__894 ,w__2 ,w__795);
  xnor g__1014(w__893 ,w__737 ,w__800);
  xnor g__1015(w__892 ,w__713 ,w__805);
  not g__1016(w__878 ,w__877);
  not g__1017(w__876 ,w__875);
  and g__1018(w__874 ,w__657 ,w__821);
  nor g__1019(w__873 ,w__719 ,w__835);
  nor g__1020(w__872 ,w__715 ,w__823);
  nor g__1021(w__871 ,w__718 ,w__832);
  nor g__1022(w__870 ,w__790 ,w__808);
  nor g__1023(w__869 ,w__692 ,w__809);
  nor g__1024(w__868 ,w__792 ,w__830);
  or g__1025(w__867 ,w__524 ,w__833);
  and g__1026(w__886 ,w__553 ,w__820);
  or g__1027(w__885 ,w__769 ,w__826);
  or g__1028(w__884 ,w__780 ,w__828);
  and g__1029(w__883 ,w__771 ,w__819);
  or g__1030(w__882 ,w__763 ,w__811);
  and g__1031(w__881 ,w__775 ,w__825);
  or g__1032(w__880 ,w__539 ,w__810);
  or g__1033(w__879 ,w__786 ,w__836);
  and g__1034(w__877 ,w__778 ,w__838);
  or g__1035(w__875 ,w__766 ,w__816);
  not g__1036(w__861 ,w__860);
  not g__1037(w__857 ,w__858);
  not g__1038(w__855 ,w__854);
  xor g__1039(w__852 ,w__792 ,w__745);
  xnor g__1040(w__851 ,w__743 ,w__739);
  xor g__1041(w__850 ,w__715 ,w__755);
  xnor g__1042(w__848 ,w__762 ,w__729);
  xnor g__1043(w__847 ,w__424 ,w__759);
  xor g__1044(w__846 ,w__678 ,w__790);
  xnor g__1045(w__866 ,w__399 ,w__733);
  xnor g__1046(w__865 ,w__760 ,w__607);
  xnor g__1047(w__864 ,w__658 ,w__728);
  xnor g__1048(w__863 ,w__619 ,w__734);
  xnor g__1049(w__862 ,w__546 ,w__725);
  xnor g__1050(w__860 ,w__724 ,w__732);
  xnor g__1051(w__859 ,w__618 ,w__726);
  xnor g__1052(w__858 ,w__693 ,w__730);
  xnor g__1053(w__856 ,w__548 ,w__727);
  xnor g__1054(w__854 ,w__721 ,w__731);
  xnor g__1055(w__853 ,w__757 ,w__604);
  not g__1056(w__844 ,w__845);
  not g__1057(w__841 ,w__840);
  or g__1058(w__838 ,w__774 ,w__758);
  nor g__1059(w__837 ,w__670 ,w__752);
  nor g__1060(w__836 ,w__720 ,w__784);
  and g__1061(w__835 ,w__670 ,w__752);
  and g__1062(w__834 ,w__686 ,w__749);
  and g__1063(w__833 ,w__525 ,w__757);
  nor g__1064(w__832 ,w__686 ,w__749);
  or g__1065(w__831 ,w__706 ,w__789);
  and g__1066(w__830 ,w__746 ,w__747);
  and g__1067(w__829 ,w__755 ,w__756);
  and g__1068(w__828 ,w__793 ,w__777);
  and g__1069(w__827 ,w__678 ,w__740);
  and g__1070(w__826 ,w__791 ,w__776);
  or g__1071(w__825 ,w__690 ,w__773);
  nor g__1072(w__824 ,w__746 ,w__747);
  nor g__1073(w__823 ,w__755 ,w__756);
  nor g__1074(w__822 ,w__688 ,w__737);
  or g__1075(w__821 ,w__689 ,w__736);
  or g__1076(w__820 ,w__552 ,w__761);
  or g__1077(w__819 ,w__714 ,w__770);
  or g__1078(w__845 ,w__704 ,w__767);
  and g__1079(w__843 ,w__703 ,w__785);
  or g__1080(w__842 ,w__700 ,w__772);
  or g__1081(w__840 ,w__697 ,w__782);
  or g__1082(w__839 ,w__698 ,w__783);
  and g__1083(w__816 ,w__691 ,w__765);
  and g__1084(w__815 ,w__676 ,w__744);
  and g__1085(w__814 ,w__706 ,w__789);
  nor g__1086(w__813 ,w__742 ,w__739);
  or g__1087(w__812 ,w__743 ,w__738);
  nor g__1088(w__811 ,w__717 ,w__764);
  and g__1089(w__810 ,w__534 ,w__759);
  nor g__1090(w__809 ,w__676 ,w__744);
  nor g__1091(w__808 ,w__678 ,w__740);
  xnor g__1092(w__807 ,w__677 ,w__712);
  xnor g__1093(w__806 ,w__679 ,w__709);
  xnor g__1094(w__805 ,w__654 ,w__673);
  xor g__1095(w__804 ,w__692 ,w__676);
  xor g__1096(w__803 ,w__670 ,w__719);
  xnor g__1097(w__802 ,w__589 ,w__723);
  xnor g__1098(w__801 ,w__711 ,w__690);
  xnor g__1099(w__800 ,w__657 ,w__689);
  xnor g__1100(w__799 ,w__650 ,w__671);
  xor g__1101(w__798 ,w__720 ,w__652);
  xor g__1102(w__797 ,w__718 ,w__686);
  xnor g__1103(w__796 ,w__685 ,w__684);
  xnor g__1104(w__795 ,w__683 ,w__708);
  xnor g__1105(w__794 ,w__716 ,w__675);
  or g__1106(w__818 ,w__665 ,w__768);
  or g__1107(w__817 ,w__664 ,w__781);
  not g__1108(w__789 ,w__788);
  or g__1109(w__787 ,w__650 ,w__671);
  and g__1110(w__786 ,w__652 ,w__687);
  or g__1111(w__785 ,w__702 ,w__722);
  nor g__1112(w__784 ,w__652 ,w__687);
  nor g__1113(w__783 ,w__660 ,w__694);
  nor g__1114(w__782 ,w__695 ,w__723);
  and g__1115(w__781 ,w__658 ,w__705);
  and g__1116(w__780 ,w__685 ,w__684);
  and g__1117(w__779 ,w__650 ,w__671);
  or g__1118(w__778 ,w__682 ,w__707);
  or g__1119(w__777 ,w__685 ,w__684);
  or g__1120(w__776 ,w__679 ,w__709);
  or g__1121(w__775 ,w__710 ,w__680);
  nor g__1122(w__774 ,w__683 ,w__708);
  nor g__1123(w__773 ,w__711 ,w__681);
  nor g__1124(w__772 ,w__659 ,w__701);
  or g__1125(w__771 ,w__653 ,w__673);
  nor g__1126(w__770 ,w__654 ,w__672);
  and g__1127(w__769 ,w__679 ,w__709);
  and g__1128(w__768 ,w__663 ,w__693);
  and g__1129(w__767 ,w__668 ,w__724);
  and g__1130(w__766 ,w__677 ,w__712);
  or g__1131(w__765 ,w__677 ,w__712);
  nor g__1132(w__764 ,w__675 ,w__674);
  and g__1133(w__763 ,w__675 ,w__674);
  nor g__1134(w__762 ,w__527 ,w__666);
  or g__1135(w__793 ,w__643 ,w__699);
  or g__1136(w__791 ,w__631 ,w__669);
  and g__1137(w__790 ,w__536 ,w__667);
  and g__1138(w__788 ,w__569 ,w__696);
  not g__1139(w__761 ,w__760);
  not g__1140(w__758 ,w__2);
  not g__1141(w__754 ,w__753);
  not g__1142(w__750 ,w__751);
  not g__1143(w__746 ,w__745);
  not g__1144(w__742 ,w__743);
  not g__1145(w__738 ,w__739);
  not g__1146(w__736 ,w__737);
  xnor g__1147(w__734 ,w__659 ,w__490);
  xnor g__1148(w__733 ,w__500 ,w__627);
  xnor g__1149(w__732 ,w__479 ,w__624);
  xnor g__1150(w__731 ,w__481 ,w__626);
  xnor g__1151(w__730 ,w__405 ,w__622);
  xnor g__1152(w__729 ,w__611 ,w__603);
  xnor g__1153(w__728 ,w__415 ,w__617);
  xnor g__1154(w__727 ,w__433 ,w__656);
  xor g__1155(w__726 ,w__430 ,w__660);
  xnor g__1156(w__725 ,w__545 ,w__655);
  xnor g__1157(w__760 ,w__381 ,w__600);
  xnor g__1158(w__757 ,w__331 ,w__591);
  xnor g__1159(w__756 ,w__429 ,w__592);
  xnor g__1160(w__755 ,w__327 ,w__598);
  xnor g__1161(w__753 ,w__502 ,w__596);
  xnor g__1162(w__752 ,w__505 ,w__602);
  xnor g__1163(w__751 ,w__661 ,w__601);
  xnor g__1164(w__749 ,w__408 ,w__599);
  xnor g__1165(w__748 ,w__407 ,w__605);
  xnor g__1166(w__747 ,w__397 ,w__606);
  xnor g__1167(w__745 ,w__414 ,w__593);
  xnor g__1168(w__744 ,w__383 ,w__608);
  xnor g__1169(w__743 ,w__423 ,w__595);
  xnor g__1170(w__741 ,w__425 ,w__597);
  xnor g__1171(w__740 ,w__436 ,w__612);
  xnor g__1172(w__737 ,w__628 ,w__613);
  xnor g__1173(w__735 ,w__489 ,w__609);
  not g__1174(w__722 ,w__721);
  not g__1175(w__717 ,w__716);
  not g__1176(w__714 ,w__713);
  not g__1177(w__710 ,w__711);
  not g__1178(w__707 ,w__708);
  or g__1179(w__705 ,w__415 ,w__617);
  nor g__1180(w__704 ,w__479 ,w__623);
  or g__1181(w__703 ,w__480 ,w__625);
  nor g__1182(w__702 ,w__481 ,w__626);
  and g__1183(w__701 ,w__490 ,w__620);
  nor g__1184(w__700 ,w__490 ,w__620);
  and g__1185(w__699 ,w__656 ,w__640);
  and g__1186(w__698 ,w__430 ,w__618);
  and g__1187(w__697 ,w__589 ,w__651);
  or g__1188(w__696 ,w__588 ,w__628);
  nor g__1189(w__695 ,w__589 ,w__651);
  nor g__1190(w__694 ,w__430 ,w__618);
  or g__1191(w__724 ,w__567 ,w__647);
  and g__1192(w__723 ,w__570 ,w__644);
  or g__1193(w__721 ,w__572 ,w__638);
  and g__1194(w__720 ,w__585 ,w__645);
  and g__1195(w__719 ,w__584 ,w__648);
  and g__1196(w__718 ,w__580 ,w__646);
  and g__1197(w__715 ,w__579 ,w__639);
  or g__1198(w__713 ,w__540 ,w__634);
  or g__1199(w__712 ,w__576 ,w__630);
  or g__1200(w__711 ,w__560 ,w__636);
  or g__1201(w__709 ,w__549 ,w__633);
  or g__1202(w__708 ,w__563 ,w__637);
  or g__1203(w__706 ,w__566 ,w__642);
  not g__1204(w__688 ,w__689);
  not g__1205(w__682 ,w__683);
  not g__1206(w__680 ,w__681);
  not g__1207(w__672 ,w__673);
  and g__1208(w__669 ,w__655 ,w__635);
  or g__1209(w__668 ,w__478 ,w__624);
  or g__1210(w__667 ,w__662 ,w__528);
  nor g__1211(w__666 ,w__627 ,w__530);
  nor g__1212(w__665 ,w__404 ,w__622);
  and g__1213(w__664 ,w__415 ,w__617);
  or g__1214(w__663 ,w__405 ,w__621);
  or g__1215(w__693 ,w__538 ,w__649);
  and g__1216(w__692 ,w__557 ,w__641);
  or g__1217(w__691 ,w__542 ,w__632);
  and g__1218(w__690 ,w__558 ,w__616);
  or g__1219(w__689 ,w__535 ,w__615);
  xnor g__1220(w__687 ,w__368 ,w__520);
  xnor g__1221(w__686 ,w__504 ,w__519);
  xnor g__1222(w__685 ,w__387 ,w__518);
  xnor g__1223(w__684 ,w__496 ,w__517);
  xnor g__1224(w__683 ,w__328 ,w__515);
  xnor g__1225(w__681 ,w__446 ,w__513);
  xnor g__1226(w__679 ,w__374 ,w__512);
  xnor g__1227(w__678 ,w__385 ,w__514);
  xnor g__1228(w__677 ,w__323 ,w__511);
  xnor g__1229(w__676 ,w__438 ,w__523);
  xnor g__1230(w__674 ,w__428 ,w__510);
  xnor g__1231(w__673 ,w__364 ,w__516);
  xnor g__1232(w__671 ,w__343 ,w__522);
  xor g__1233(w__670 ,w__494 ,w__521);
  not g__1234(w__662 ,w__661);
  not g__1235(w__653 ,w__654);
  nor g__1236(w__649 ,w__447 ,w__533);
  or g__1237(w__648 ,w__590 ,w__581);
  nor g__1238(w__647 ,w__380 ,w__575);
  or g__1239(w__646 ,w__503 ,w__578);
  or g__1240(w__645 ,w__382 ,w__583);
  or g__1241(w__644 ,w__506 ,w__568);
  nor g__1242(w__643 ,w__432 ,w__548);
  and g__1243(w__642 ,w__381 ,w__565);
  or g__1244(w__641 ,w__505 ,w__529);
  or g__1245(w__640 ,w__433 ,w__547);
  or g__1246(w__639 ,w__384 ,w__551);
  and g__1247(w__638 ,w__383 ,w__556);
  nor g__1248(w__637 ,w__439 ,w__559);
  nor g__1249(w__636 ,w__449 ,w__561);
  or g__1250(w__635 ,w__545 ,w__546);
  nor g__1251(w__634 ,w__443 ,w__550);
  nor g__1252(w__633 ,w__442 ,w__582);
  nor g__1253(w__632 ,w__344 ,w__537);
  and g__1254(w__631 ,w__545 ,w__546);
  nor g__1255(w__630 ,w__440 ,w__543);
  or g__1256(w__629 ,w__459 ,w__532);
  or g__1257(w__661 ,w__467 ,w__531);
  and g__1258(w__660 ,w__469 ,w__571);
  and g__1259(w__659 ,w__457 ,w__555);
  or g__1260(w__658 ,w__462 ,w__577);
  or g__1261(w__657 ,w__460 ,w__544);
  or g__1262(w__656 ,w__463 ,w__564);
  or g__1263(w__655 ,w__458 ,w__541);
  or g__1264(w__654 ,w__456 ,w__554);
  or g__1265(w__652 ,w__475 ,w__586);
  or g__1266(w__651 ,w__468 ,w__573);
  or g__1267(w__650 ,w__472 ,w__587);
  not g__1268(w__625 ,w__626);
  not g__1269(w__623 ,w__624);
  not g__1270(w__621 ,w__622);
  not g__1271(w__620 ,w__619);
  or g__1272(w__616 ,w__508 ,w__1);
  nor g__1273(w__615 ,w__445 ,w__526);
  xnor g__1274(w__614 ,w__426 ,w__4008);
  xnor g__1275(w__613 ,w__370 ,w__420);
  xor g__1276(w__612 ,w__442 ,w__416);
  xnor g__1277(w__610 ,w__435 ,w__396);
  xor g__1278(w__609 ,w__440 ,w__417);
  xnor g__1279(w__608 ,w__409 ,w__431);
  xnor g__1280(w__607 ,w__488 ,w__401);
  xnor g__1281(w__606 ,w__507 ,w__410);
  xnor g__1282(w__605 ,w__506 ,w__413);
  xnor g__1283(w__604 ,w__339 ,w__501);
  xnor g__1284(w__603 ,w__311 ,w__450);
  xnor g__1285(w__602 ,w__337 ,w__403);
  xnor g__1286(w__601 ,w__412 ,w__422);
  xnor g__1287(w__600 ,w__360 ,w__482);
  xor g__1288(w__599 ,w__447 ,w__427);
  xnor g__1289(w__598 ,w__358 ,w__448);
  xor g__1290(w__597 ,w__439 ,w__418);
  xnor g__1291(w__596 ,w__486 ,w__484);
  xor g__1292(w__595 ,w__443 ,w__334);
  xnor g__1293(w__594 ,w__498 ,w__493);
  xor g__1294(w__593 ,w__449 ,w__359);
  xnor g__1295(w__592 ,w__375 ,w__444);
  xnor g__1296(w__591 ,w__335 ,w__441);
  xnor g__1297(w__628 ,w__392 ,w__4037);
  xnor g__1298(w__627 ,w__393 ,w__4038);
  xnor g__1299(w__626 ,w__180 ,w__394);
  xnor g__1300(w__624 ,w__176 ,w__395);
  xnor g__1301(w__622 ,w__342 ,w__389);
  xnor g__1302(w__619 ,w__120 ,w__391);
  xnor g__1303(w__618 ,w__117 ,w__388);
  xnor g__1304(w__617 ,w__179 ,w__390);
  nor g__1305(w__588 ,w__370 ,w__420);
  and g__1306(w__587 ,w__477 ,w__504);
  and g__1307(w__586 ,w__387 ,w__474);
  or g__1308(w__585 ,w__356 ,w__495);
  or g__1309(w__584 ,w__497 ,w__492);
  nor g__1310(w__583 ,w__355 ,w__496);
  nor g__1311(w__582 ,w__436 ,w__416);
  nor g__1312(w__581 ,w__498 ,w__493);
  or g__1313(w__580 ,w__485 ,w__483);
  or g__1314(w__579 ,w__362 ,w__437);
  nor g__1315(w__578 ,w__486 ,w__484);
  nor g__1316(w__577 ,w__378 ,w__476);
  and g__1317(w__576 ,w__417 ,w__489);
  nor g__1318(w__575 ,w__367 ,w__494);
  or g__1319(w__574 ,w__434 ,w__396);
  and g__1320(w__573 ,w__466 ,w__446);
  and g__1321(w__572 ,w__409 ,w__431);
  or g__1322(w__571 ,w__377 ,w__465);
  or g__1323(w__570 ,w__5 ,w__406);
  or g__1324(w__569 ,w__369 ,w__419);
  nor g__1325(w__568 ,w__3 ,w__407);
  and g__1326(w__567 ,w__367 ,w__494);
  and g__1327(w__566 ,w__360 ,w__482);
  or g__1328(w__565 ,w__360 ,w__482);
  and g__1329(w__564 ,w__379 ,w__461);
  and g__1330(w__563 ,w__425 ,w__418);
  and g__1331(w__562 ,w__4008 ,w__426);
  nor g__1332(w__561 ,w__359 ,w__414);
  and g__1333(w__560 ,w__359 ,w__414);
  nor g__1334(w__559 ,w__425 ,w__418);
  or g__1335(w__558 ,w__4 ,w__397);
  or g__1336(w__557 ,w__336 ,w__402);
  or g__1337(w__556 ,w__409 ,w__431);
  or g__1338(w__555 ,w__386 ,w__454);
  nor g__1339(w__554 ,w__341 ,w__455);
  or g__1340(w__553 ,w__487 ,w__401);
  nor g__1341(w__552 ,w__488 ,w__400);
  nor g__1342(w__551 ,w__361 ,w__438);
  nor g__1343(w__550 ,w__334 ,w__423);
  and g__1344(w__549 ,w__436 ,w__416);
  and g__1345(w__590 ,w__353 ,w__471);
  or g__1346(w__589 ,w__303 ,w__451);
  not g__1347(w__547 ,w__548);
  and g__1348(w__544 ,w__464 ,w__448);
  nor g__1349(w__543 ,w__417 ,w__489);
  and g__1350(w__542 ,w__338 ,w__428);
  and g__1351(w__541 ,w__343 ,w__453);
  and g__1352(w__540 ,w__334 ,w__423);
  and g__1353(w__539 ,w__491 ,w__424);
  and g__1354(w__538 ,w__427 ,w__408);
  nor g__1355(w__537 ,w__338 ,w__428);
  or g__1356(w__536 ,w__411 ,w__421);
  and g__1357(w__535 ,w__375 ,w__429);
  or g__1358(w__534 ,w__491 ,w__424);
  nor g__1359(w__533 ,w__427 ,w__408);
  and g__1360(w__532 ,w__470 ,w__441);
  nor g__1361(w__531 ,w__346 ,w__473);
  and g__1362(w__530 ,w__499 ,w__399);
  nor g__1363(w__529 ,w__337 ,w__403);
  nor g__1364(w__528 ,w__412 ,w__422);
  and g__1365(w__527 ,w__500 ,w__398);
  nor g__1366(w__526 ,w__375 ,w__429);
  or g__1367(w__525 ,w__339 ,w__501);
  and g__1368(w__524 ,w__339 ,w__501);
  xnor g__1369(w__523 ,w__384 ,w__362);
  xnor g__1370(w__522 ,w__322 ,w__329);
  xor g__1371(w__521 ,w__380 ,w__367);
  xnor g__1372(w__520 ,w__345 ,w__4045);
  xnor g__1373(w__519 ,w__365 ,w__324);
  xnor g__1374(w__518 ,w__357 ,w__3935);
  xnor g__1375(w__517 ,w__356 ,w__382);
  xnor g__1376(w__516 ,w__178 ,w__379);
  xor g__1377(w__515 ,w__378 ,w__330);
  xnor g__1378(w__514 ,w__326 ,w__333);
  xnor g__1379(w__513 ,w__366 ,w__354);
  xor g__1380(w__512 ,w__377 ,w__372);
  xor g__1381(w__511 ,w__341 ,w__340);
  xor g__1382(w__510 ,w__344 ,w__338);
  xnor g__1383(w__509 ,w__313 ,w__312);
  xnor g__1384(w__548 ,w__376 ,w__315);
  xnor g__1385(w__546 ,w__239 ,w__314);
  or g__1386(w__545 ,w__350 ,w__452);
  not g__1387(w__508 ,w__507);
  not g__1388(w__503 ,w__502);
  not g__1389(w__499 ,w__500);
  not g__1390(w__497 ,w__498);
  not g__1391(w__495 ,w__496);
  not g__1392(w__492 ,w__493);
  not g__1393(w__487 ,w__488);
  not g__1394(w__485 ,w__486);
  not g__1395(w__483 ,w__484);
  not g__1396(w__480 ,w__481);
  not g__1397(w__479 ,w__478);
  or g__1398(w__477 ,w__365 ,w__324);
  nor g__1399(w__476 ,w__328 ,w__330);
  and g__1400(w__475 ,w__3935 ,w__357);
  or g__1401(w__474 ,w__3935 ,w__357);
  nor g__1402(w__473 ,w__4045 ,w__368);
  and g__1403(w__472 ,w__365 ,w__324);
  or g__1404(w__471 ,w__120 ,w__352);
  or g__1405(w__470 ,w__335 ,w__331);
  or g__1406(w__469 ,w__371 ,w__373);
  and g__1407(w__468 ,w__366 ,w__354);
  and g__1408(w__467 ,w__4045 ,w__368);
  or g__1409(w__466 ,w__366 ,w__354);
  nor g__1410(w__465 ,w__372 ,w__374);
  or g__1411(w__464 ,w__358 ,w__327);
  nor g__1412(w__463 ,w__178 ,w__363);
  and g__1413(w__462 ,w__328 ,w__330);
  or g__1414(w__461 ,w__177 ,w__364);
  and g__1415(w__460 ,w__358 ,w__327);
  and g__1416(w__459 ,w__335 ,w__331);
  and g__1417(w__458 ,w__322 ,w__329);
  or g__1418(w__457 ,w__325 ,w__332);
  and g__1419(w__456 ,w__340 ,w__323);
  nor g__1420(w__455 ,w__340 ,w__323);
  nor g__1421(w__454 ,w__326 ,w__333);
  or g__1422(w__453 ,w__322 ,w__329);
  and g__1423(w__452 ,w__342 ,w__351);
  and g__1424(w__451 ,w__266 ,w__376);
  or g__1425(w__450 ,w__126 ,w__319);
  or g__1426(w__507 ,w__105 ,w__321);
  and g__1427(w__506 ,w__72 ,w__349);
  and g__1428(w__505 ,w__285 ,w__348);
  xnor g__1429(w__504 ,w__247 ,w__3998);
  xnor g__1430(w__502 ,w__199 ,w__4059);
  or g__1431(w__501 ,w__65 ,w__318);
  xnor g__1432(w__500 ,w__185 ,w__4100);
  xnor g__1433(w__498 ,w__222 ,w__4002);
  xnor g__1434(w__496 ,w__221 ,w__3982);
  xnor g__1435(w__494 ,w__193 ,w__4003);
  xnor g__1436(w__493 ,w__231 ,w__4018);
  xnor g__1437(w__491 ,w__230 ,w__4101);
  and g__1438(w__490 ,w__310 ,w__320);
  xnor g__1439(w__489 ,w__228 ,w__3993);
  or g__1440(w__488 ,w__305 ,w__347);
  xnor g__1441(w__486 ,w__226 ,w__3951);
  xnor g__1442(w__484 ,w__192 ,w__3997);
  xnor g__1443(w__482 ,w__206 ,w__3960);
  or g__1444(w__481 ,w__267 ,w__317);
  or g__1445(w__478 ,w__262 ,w__316);
  not g__1446(w__445 ,w__444);
  not g__1447(w__437 ,w__438);
  not g__1448(w__434 ,w__435);
  not g__1449(w__432 ,w__433);
  not g__1450(w__421 ,w__422);
  not g__1451(w__419 ,w__420);
  not g__1452(w__411 ,w__412);
  not g__1453(w__406 ,w__407);
  not g__1454(w__404 ,w__405);
  not g__1455(w__402 ,w__403);
  not g__1456(w__400 ,w__401);
  not g__1457(w__398 ,w__399);
  xnor g__1458(w__395 ,w__245 ,w__4066);
  xnor g__1459(w__394 ,w__243 ,w__3943);
  xnor g__1460(w__393 ,w__240 ,w__4023);
  xnor g__1461(w__392 ,w__244 ,w__4022);
  xnor g__1462(w__391 ,w__235 ,w__4063);
  xnor g__1463(w__390 ,w__241 ,w__4081);
  xnor g__1464(w__389 ,w__237 ,w__3937);
  xnor g__1465(w__388 ,w__242 ,w__4080);
  xor g__1466(w__449 ,w__207 ,w__4026);
  xnor g__1467(w__448 ,w__215 ,w__3959);
  xor g__1468(w__447 ,w__213 ,w__3952);
  xnor g__1469(w__446 ,w__184 ,w__3996);
  xnor g__1470(w__444 ,w__224 ,w__3974);
  xor g__1471(w__443 ,w__183 ,w__3979);
  xor g__1472(w__442 ,w__201 ,w__4093);
  xnor g__1473(w__441 ,w__208 ,w__3961);
  xor g__1474(w__440 ,w__203 ,w__4009);
  xor g__1475(w__439 ,w__187 ,w__4017);
  xnor g__1476(w__438 ,w__227 ,w__4020);
  xnor g__1477(w__436 ,w__200 ,w__3954);
  xnor g__1478(w__435 ,w__198 ,w__4072);
  xnor g__1479(w__433 ,w__219 ,w__3950);
  xnor g__1480(w__431 ,w__214 ,w__4097);
  xnor g__1481(w__430 ,w__223 ,w__3987);
  xnor g__1482(w__429 ,w__189 ,w__4067);
  xnor g__1483(w__428 ,w__194 ,w__4024);
  xnor g__1484(w__427 ,w__216 ,w__4014);
  xnor g__1485(w__425 ,w__188 ,w__3955);
  xnor g__1486(w__424 ,w__248 ,w__4039);
  xnor g__1487(w__423 ,w__202 ,w__3932);
  xnor g__1488(w__422 ,w__211 ,w__3968);
  xnor g__1489(w__420 ,w__197 ,w__4099);
  xnor g__1490(w__418 ,w__225 ,w__4094);
  xnor g__1491(w__417 ,w__195 ,w__3962);
  xnor g__1492(w__416 ,w__217 ,w__4016);
  xnor g__1493(w__415 ,w__204 ,w__3988);
  xnor g__1494(w__414 ,w__233 ,w__4042);
  xnor g__1495(w__413 ,w__190 ,w__4012);
  xnor g__1496(w__412 ,w__220 ,w__3953);
  xnor g__1497(w__410 ,w__205 ,w__3964);
  xnor g__1498(w__409 ,w__218 ,w__3958);
  xnor g__1499(w__408 ,w__196 ,w__4029);
  xnor g__1500(w__407 ,w__191 ,w__4027);
  xnor g__1501(w__405 ,w__209 ,w__4061);
  xnor g__1502(w__403 ,w__186 ,w__4019);
  xnor g__1503(w__401 ,w__181 ,w__232);
  xnor g__1504(w__399 ,w__182 ,w__212);
  xnor g__1505(w__397 ,w__238 ,w__210);
  xnor g__1506(w__396 ,w__246 ,w__229);
  not g__1507(w__386 ,w__385);
  not g__1508(w__373 ,w__374);
  not g__1509(w__371 ,w__372);
  not g__1510(w__369 ,w__370);
  not g__1511(w__363 ,w__364);
  not g__1512(w__362 ,w__361);
  not g__1513(w__356 ,w__355);
  or g__1514(w__353 ,w__17 ,w__235);
  nor g__1515(w__352 ,w__4063 ,w__234);
  or g__1516(w__351 ,w__3937 ,w__236);
  nor g__1517(w__350 ,w__10 ,w__237);
  or g__1518(w__349 ,w__155 ,w__238);
  or g__1519(w__348 ,w__260 ,w__242);
  nor g__1520(w__347 ,w__302 ,w__243);
  or g__1521(w__387 ,w__98 ,w__306);
  or g__1522(w__385 ,w__71 ,w__308);
  and g__1523(w__384 ,w__99 ,w__281);
  or g__1524(w__383 ,w__134 ,w__273);
  and g__1525(w__382 ,w__125 ,w__300);
  or g__1526(w__381 ,w__160 ,w__297);
  and g__1527(w__380 ,w__148 ,w__295);
  or g__1528(w__379 ,w__77 ,w__283);
  and g__1529(w__378 ,w__144 ,w__251);
  and g__1530(w__377 ,w__113 ,w__286);
  or g__1531(w__376 ,w__142 ,w__294);
  or g__1532(w__375 ,w__78 ,w__287);
  or g__1533(w__374 ,w__114 ,w__288);
  or g__1534(w__372 ,w__168 ,w__292);
  or g__1535(w__370 ,w__166 ,w__259);
  or g__1536(w__368 ,w__151 ,w__299);
  or g__1537(w__367 ,w__140 ,w__304);
  or g__1538(w__366 ,w__139 ,w__293);
  or g__1539(w__365 ,w__82 ,w__252);
  or g__1540(w__364 ,w__108 ,w__284);
  or g__1541(w__361 ,w__106 ,w__291);
  or g__1542(w__360 ,w__101 ,w__265);
  or g__1543(w__359 ,w__132 ,w__282);
  or g__1544(w__358 ,w__81 ,w__269);
  or g__1545(w__357 ,w__173 ,w__309);
  or g__1546(w__355 ,w__88 ,w__301);
  or g__1547(w__354 ,w__68 ,w__290);
  not g__1548(w__346 ,w__345);
  not g__1549(w__336 ,w__337);
  not g__1550(w__332 ,w__333);
  not g__1551(w__325 ,w__326);
  nor g__1552(w__321 ,w__62 ,w__246);
  or g__1553(w__320 ,w__280 ,w__239);
  nor g__1554(w__319 ,w__73 ,w__240);
  nor g__1555(w__318 ,w__100 ,w__244);
  nor g__1556(w__317 ,w__256 ,w__245);
  nor g__1557(w__316 ,w__261 ,w__241);
  xnor g__1558(w__315 ,w__175 ,w__4043);
  xnor g__1559(w__314 ,w__119 ,w__4062);
  or g__1560(w__313 ,w__115 ,w__298);
  or g__1561(w__312 ,w__141 ,w__249);
  or g__1562(w__311 ,w__107 ,w__258);
  or g__1563(w__345 ,w__85 ,w__296);
  and g__1564(w__344 ,w__111 ,w__268);
  or g__1565(w__343 ,w__91 ,w__263);
  or g__1566(w__342 ,w__94 ,w__278);
  and g__1567(w__341 ,w__149 ,w__274);
  or g__1568(w__340 ,w__109 ,w__277);
  or g__1569(w__339 ,w__152 ,w__250);
  or g__1570(w__337 ,w__95 ,w__253);
  or g__1571(w__335 ,w__167 ,w__264);
  or g__1572(w__334 ,w__136 ,w__289);
  or g__1573(w__333 ,w__161 ,w__276);
  or g__1574(w__331 ,w__92 ,w__270);
  or g__1575(w__330 ,w__84 ,w__254);
  or g__1576(w__329 ,w__102 ,w__272);
  or g__1577(w__328 ,w__63 ,w__255);
  or g__1578(w__327 ,w__66 ,w__307);
  or g__1579(w__326 ,w__110 ,w__271);
  or g__1580(w__324 ,w__147 ,w__279);
  or g__1581(w__323 ,w__138 ,w__275);
  or g__1582(w__322 ,w__163 ,w__257);
  or g__1583(w__310 ,w__39 ,w__119);
  and g__1584(w__309 ,w__4089 ,w__129);
  and g__1585(w__308 ,w__4092 ,w__156);
  and g__1586(w__307 ,w__3989 ,w__150);
  and g__1587(w__306 ,w__4105 ,w__79);
  nor g__1588(w__305 ,w__19 ,w__180);
  and g__1589(w__304 ,w__3956 ,w__97);
  nor g__1590(w__303 ,w__7 ,w__175);
  and g__1591(w__302 ,w__19 ,w__180);
  and g__1592(w__301 ,w__4074 ,w__165);
  or g__1593(w__300 ,w__50 ,w__154);
  and g__1594(w__299 ,w__4106 ,w__162);
  and g__1595(w__298 ,w__4007 ,w__122);
  and g__1596(w__297 ,w__3974 ,w__157);
  and g__1597(w__296 ,w__4044 ,w__143);
  or g__1598(w__295 ,w__31 ,w__86);
  and g__1599(w__294 ,w__4042 ,w__121);
  and g__1600(w__293 ,w__3964 ,w__70);
  and g__1601(w__292 ,w__4000 ,w__135);
  and g__1602(w__291 ,w__4065 ,w__60);
  and g__1603(w__290 ,w__4026 ,w__169);
  and g__1604(w__289 ,w__4024 ,w__103);
  and g__1605(w__288 ,w__3985 ,w__74);
  and g__1606(w__287 ,w__4097 ,w__130);
  or g__1607(w__286 ,w__52 ,w__127);
  or g__1608(w__285 ,w__20 ,w__117);
  and g__1609(w__284 ,w__3979 ,w__90);
  and g__1610(w__283 ,w__3932 ,w__146);
  and g__1611(w__282 ,w__4072 ,w__170);
  or g__1612(w__281 ,w__30 ,w__112);
  nor g__1613(w__280 ,w__4062 ,w__118);
  and g__1614(w__279 ,w__3966 ,w__171);
  and g__1615(w__278 ,w__4107 ,w__158);
  and g__1616(w__277 ,w__3962 ,w__145);
  and g__1617(w__276 ,w__4077 ,w__96);
  and g__1618(w__275 ,w__4055 ,w__93);
  or g__1619(w__274 ,w__42 ,w__153);
  and g__1620(w__273 ,w__3957 ,w__61);
  and g__1621(w__272 ,w__4076 ,w__80);
  and g__1622(w__271 ,w__4030 ,w__128);
  and g__1623(w__270 ,w__4099 ,w__159);
  and g__1624(w__269 ,w__3958 ,w__104);
  or g__1625(w__268 ,w__32 ,w__67);
  nor g__1626(w__267 ,w__14 ,w__176);
  or g__1627(w__266 ,w__4043 ,w__174);
  and g__1628(w__265 ,w__3959 ,w__124);
  and g__1629(w__264 ,w__3960 ,w__76);
  and g__1630(w__263 ,w__4091 ,w__89);
  nor g__1631(w__262 ,w__18 ,w__179);
  and g__1632(w__261 ,w__18 ,w__179);
  nor g__1633(w__260 ,w__4080 ,w__116);
  and g__1634(w__259 ,w__4067 ,w__87);
  and g__1635(w__258 ,w__4085 ,w__75);
  and g__1636(w__257 ,w__3936 ,w__133);
  and g__1637(w__256 ,w__14 ,w__176);
  and g__1638(w__255 ,w__4001 ,w__69);
  and g__1639(w__254 ,w__4079 ,w__164);
  and g__1640(w__253 ,w__4111 ,w__137);
  and g__1641(w__252 ,w__4028 ,w__83);
  or g__1642(w__251 ,w__23 ,w__172);
  nor g__1643(w__250 ,w__181 ,w__123);
  nor g__1644(w__249 ,w__182 ,w__64);
  xnor g__1645(w__248 ,w__4070 ,w__3946);
  xnor g__1646(w__247 ,w__4091 ,w__3967);
  not g__1647(w__236 ,w__237);
  not g__1648(w__234 ,w__235);
  xnor g__1649(w__233 ,w__4011 ,w__3949);
  xnor g__1650(w__232 ,w__3975 ,w__3944);
  xnor g__1651(w__231 ,w__4049 ,w__3956);
  xnor g__1652(w__229 ,w__4041 ,w__3994);
  xnor g__1653(w__228 ,w__4055 ,w__3931);
  xnor g__1654(w__227 ,w__3989 ,w__3973);
  xnor g__1655(w__226 ,w__4106 ,in5[5]);
  xnor g__1656(w__225 ,w__4048 ,w__4001);
  xnor g__1657(w__224 ,w__4098 ,w__4005);
  xnor g__1658(w__223 ,w__4111 ,w__4095);
  xnor g__1659(w__222 ,w__4064 ,w__4033);
  xnor g__1660(w__221 ,w__4044 ,w__4013);
  xnor g__1661(w__220 ,w__4077 ,w__4046);
  xnor g__1662(w__219 ,w__4074 ,w__3981);
  xnor g__1663(w__218 ,w__4082 ,w__4035);
  xnor g__1664(w__217 ,w__3985 ,w__3969);
  xnor g__1665(w__216 ,w__4107 ,in5[6]);
  xnor g__1666(w__215 ,w__4083 ,w__4052);
  xnor g__1667(w__214 ,w__4051 ,w__4004);
  xnor g__1668(w__213 ,w__4076 ,w__3983);
  xnor g__1669(w__212 ,w__3976 ,w__3945);
  xnor g__1670(w__211 ,w__4092 ,w__3999);
  xnor g__1671(w__210 ,w__3995 ,w__3933);
  xnor g__1672(w__209 ,w__4030 ,w__4015);
  xnor g__1673(w__208 ,w__4085 ,w__4054);
  xnor g__1674(w__207 ,w__4073 ,w__3980);
  xnor g__1675(w__206 ,w__4084 ,w__4053);
  xnor g__1676(w__205 ,w__4088 ,w__4057);
  xnor g__1677(w__204 ,w__4112 ,w__4096);
  xnor g__1678(w__203 ,w__4102 ,in5[1]);
  xnor g__1679(w__202 ,w__4056 ,w__4010);
  xnor g__1680(w__201 ,w__4047 ,w__4000);
  xnor g__1681(w__200 ,w__4078 ,w__4031);
  xnor g__1682(w__199 ,w__4075 ,w__4028);
  xnor g__1683(w__198 ,w__3963 ,w__3948);
  xnor g__1684(w__197 ,w__4068 ,w__4006);
  xnor g__1685(w__196 ,w__4060 ,w__3936);
  xnor g__1686(w__195 ,w__3978 ,w__3947);
  xnor g__1687(w__194 ,w__4071 ,w__4040);
  xnor g__1688(w__193 ,w__4065 ,w__4034);
  xnor g__1689(w__192 ,w__4090 ,w__3966);
  xnor g__1690(w__191 ,w__4058 ,w__3934);
  xnor g__1691(w__190 ,w__4105 ,in5[4]);
  xnor g__1692(w__189 ,w__4036 ,w__4021);
  xnor g__1693(w__188 ,w__4079 ,w__4032);
  xnor g__1694(w__187 ,w__3986 ,w__3970);
  xnor g__1695(w__186 ,w__4050 ,w__3957);
  xnor g__1696(w__185 ,w__4069 ,w__4007);
  xnor g__1697(w__184 ,w__4089 ,w__3965);
  xnor g__1698(w__183 ,w__4087 ,w__4025);
  xnor g__1699(w__246 ,w__4103 ,in5[2]);
  xnor g__1700(w__245 ,w__4113 ,w__3942);
  xnor g__1701(w__244 ,w__4115 ,w__3991);
  xnor g__1702(w__243 ,w__4114 ,w__3990);
  xnor g__1703(w__242 ,w__3971 ,w__3940);
  xnor g__1704(w__241 ,w__3972 ,w__3941);
  xnor g__1705(w__240 ,w__4116 ,w__3992);
  xnor g__1706(w__239 ,w__4109 ,w__3938);
  xnor g__1707(w__238 ,w__4104 ,in5[3]);
  xnor g__1708(w__237 ,w__4108 ,w__3984);
  xnor g__1709(w__235 ,w__4110 ,w__3939);
  not g__1710(w__177 ,w__178);
  not g__1711(w__174 ,w__175);
  and g__1712(w__173 ,w__3996 ,w__3965);
  nor g__1713(w__172 ,w__4017 ,w__3970);
  or g__1714(w__171 ,w__4090 ,w__3997);
  or g__1715(w__170 ,w__3963 ,w__3948);
  or g__1716(w__169 ,w__4073 ,w__3980);
  and g__1717(w__168 ,w__4093 ,w__4047);
  and g__1718(w__167 ,w__4084 ,w__4053);
  and g__1719(w__166 ,w__4036 ,w__4021);
  or g__1720(w__165 ,w__3981 ,w__3950);
  or g__1721(w__164 ,w__4032 ,w__3955);
  and g__1722(w__163 ,w__4060 ,w__4029);
  or g__1723(w__162 ,in5[5] ,w__3951);
  and g__1724(w__161 ,w__4046 ,w__3953);
  and g__1725(w__160 ,w__4098 ,w__4005);
  or g__1726(w__159 ,w__4068 ,w__4006);
  or g__1727(w__158 ,in5[6] ,w__4014);
  or g__1728(w__157 ,w__4098 ,w__4005);
  or g__1729(w__156 ,w__3999 ,w__3968);
  nor g__1730(w__155 ,w__3995 ,w__3933);
  nor g__1731(w__154 ,w__4058 ,w__4027);
  nor g__1732(w__153 ,in5[1] ,w__4009);
  and g__1733(w__152 ,w__3975 ,w__3944);
  and g__1734(w__151 ,in5[5] ,w__3951);
  or g__1735(w__150 ,w__4020 ,w__3973);
  or g__1736(w__149 ,w__35 ,w__12);
  or g__1737(w__148 ,w__34 ,w__6);
  and g__1738(w__147 ,w__4090 ,w__3997);
  or g__1739(w__146 ,w__4056 ,w__4010);
  or g__1740(w__145 ,w__3978 ,w__3947);
  or g__1741(w__144 ,w__9 ,w__41);
  or g__1742(w__143 ,w__4013 ,w__3982);
  and g__1743(w__142 ,w__4011 ,w__3949);
  and g__1744(w__141 ,w__3976 ,w__3945);
  and g__1745(w__140 ,w__4049 ,w__4018);
  and g__1746(w__139 ,w__4088 ,w__4057);
  and g__1747(w__138 ,w__3993 ,w__3931);
  or g__1748(w__137 ,w__4095 ,w__3987);
  and g__1749(w__136 ,w__4071 ,w__4040);
  or g__1750(w__135 ,w__4093 ,w__4047);
  and g__1751(w__134 ,w__4050 ,w__4019);
  or g__1752(w__133 ,w__4060 ,w__4029);
  and g__1753(w__132 ,w__3963 ,w__3948);
  and g__1754(w__131 ,w__4101 ,w__3977);
  or g__1755(w__130 ,w__4051 ,w__4004);
  or g__1756(w__129 ,w__3996 ,w__3965);
  or g__1757(w__128 ,w__4061 ,w__4015);
  nor g__1758(w__127 ,w__4031 ,w__3954);
  and g__1759(w__126 ,w__4038 ,w__4023);
  or g__1760(w__125 ,w__36 ,w__40);
  or g__1761(w__124 ,w__4083 ,w__4052);
  nor g__1762(w__123 ,w__3975 ,w__3944);
  or g__1763(w__122 ,w__4100 ,w__4069);
  or g__1764(w__121 ,w__4011 ,w__3949);
  or g__1765(w__182 ,w__28 ,w__29);
  or g__1766(w__181 ,w__56 ,w__46);
  or g__1767(w__180 ,w__43 ,w__53);
  or g__1768(w__179 ,w__48 ,w__58);
  or g__1769(w__178 ,w__24 ,w__27);
  or g__1770(w__176 ,w__22 ,w__49);
  or g__1771(w__175 ,w__26 ,w__54);
  not g__1772(w__118 ,w__119);
  not g__1773(w__116 ,w__117);
  and g__1774(w__115 ,w__4100 ,w__4069);
  and g__1775(w__114 ,w__4016 ,w__3969);
  or g__1776(w__113 ,w__33 ,w__8);
  nor g__1777(w__112 ,w__4096 ,w__3988);
  or g__1778(w__111 ,w__13 ,w__16);
  and g__1779(w__110 ,w__4061 ,w__4015);
  and g__1780(w__109 ,w__3978 ,w__3947);
  and g__1781(w__108 ,w__4087 ,w__4025);
  and g__1782(w__107 ,w__4054 ,w__3961);
  and g__1783(w__106 ,w__4034 ,w__4003);
  and g__1784(w__105 ,w__4041 ,w__3994);
  or g__1785(w__104 ,w__4082 ,w__4035);
  or g__1786(w__103 ,w__4071 ,w__4040);
  and g__1787(w__102 ,w__3983 ,w__3952);
  and g__1788(w__101 ,w__4083 ,w__4052);
  nor g__1789(w__100 ,w__4037 ,w__4022);
  or g__1790(w__99 ,w__38 ,w__37);
  and g__1791(w__98 ,in5[4] ,w__4012);
  or g__1792(w__97 ,w__4049 ,w__4018);
  or g__1793(w__96 ,w__4046 ,w__3953);
  and g__1794(w__95 ,w__4095 ,w__3987);
  and g__1795(w__94 ,in5[6] ,w__4014);
  or g__1796(w__93 ,w__3993 ,w__3931);
  and g__1797(w__92 ,w__4068 ,w__4006);
  and g__1798(w__91 ,w__3998 ,w__3967);
  or g__1799(w__90 ,w__4087 ,w__4025);
  or g__1800(w__89 ,w__3998 ,w__3967);
  and g__1801(w__88 ,w__3981 ,w__3950);
  or g__1802(w__87 ,w__4036 ,w__4021);
  nor g__1803(w__86 ,w__4033 ,w__4002);
  and g__1804(w__85 ,w__4013 ,w__3982);
  and g__1805(w__84 ,w__4032 ,w__3955);
  or g__1806(w__83 ,w__4075 ,w__4059);
  and g__1807(w__82 ,w__4075 ,w__4059);
  and g__1808(w__81 ,w__4082 ,w__4035);
  or g__1809(w__80 ,w__3983 ,w__3952);
  or g__1810(w__79 ,in5[4] ,w__4012);
  and g__1811(w__78 ,w__4051 ,w__4004);
  and g__1812(w__77 ,w__4056 ,w__4010);
  or g__1813(w__76 ,w__4084 ,w__4053);
  or g__1814(w__75 ,w__4054 ,w__3961);
  or g__1815(w__74 ,w__4016 ,w__3969);
  nor g__1816(w__73 ,w__4038 ,w__4023);
  or g__1817(w__72 ,w__11 ,w__15);
  and g__1818(w__71 ,w__3999 ,w__3968);
  or g__1819(w__70 ,w__4088 ,w__4057);
  or g__1820(w__69 ,w__4094 ,w__4048);
  and g__1821(w__68 ,w__4073 ,w__3980);
  nor g__1822(w__67 ,w__4070 ,w__4039);
  and g__1823(w__66 ,w__4020 ,w__3973);
  and g__1824(w__65 ,w__4037 ,w__4022);
  nor g__1825(w__64 ,w__3976 ,w__3945);
  and g__1826(w__63 ,w__4094 ,w__4048);
  nor g__1827(w__62 ,w__4041 ,w__3994);
  or g__1828(w__61 ,w__4050 ,w__4019);
  or g__1829(w__60 ,w__4034 ,w__4003);
  or g__1830(w__59 ,w__57 ,w__25);
  or g__1831(w__120 ,w__45 ,w__55);
  or g__1832(w__119 ,w__44 ,w__47);
  or g__1833(w__117 ,w__51 ,w__21);
  not g__1834(w__58 ,w__3940);
  not g__1835(w__57 ,w__4116);
  not g__1836(w__56 ,w__4114);
  not g__1837(w__55 ,w__3938);
  not g__1838(w__54 ,w__4104);
  not g__1839(w__53 ,w__3942);
  not g__1840(w__52 ,w__4078);
  not g__1841(w__51 ,w__4110);
  not g__1842(w__50 ,w__3934);
  not g__1843(w__49 ,w__3941);
  not g__1844(w__48 ,w__3971);
  not g__1845(w__47 ,w__3984);
  not g__1846(w__46 ,w__3990);
  not g__1847(w__45 ,w__4109);
  not g__1848(w__44 ,w__4108);
  not g__1849(w__43 ,w__4113);
  not g__1850(w__42 ,w__4102);
  not g__1851(w__41 ,w__3970);
  not g__1852(w__40 ,w__4027);
  not g__1853(w__39 ,w__4062);
  not g__1854(w__38 ,w__4096);
  not g__1855(w__37 ,w__3988);
  not g__1856(w__36 ,w__4058);
  not g__1857(w__35 ,in5[1]);
  not g__1858(w__34 ,w__4033);
  not g__1859(w__33 ,w__4031);
  not g__1860(w__32 ,w__3946);
  not g__1861(w__31 ,w__4064);
  not g__1862(w__30 ,w__4112);
  not g__1863(w__29 ,w__3991);
  not g__1864(w__28 ,w__4115);
  not g__1865(w__27 ,w__4103);
  not g__1866(w__26 ,in5[3]);
  not g__1867(w__25 ,w__3992);
  not g__1868(w__24 ,in5[2]);
  not g__1869(w__23 ,w__3986);
  not g__1870(w__22 ,w__3972);
  not g__1871(w__21 ,w__3939);
  not g__1872(w__20 ,w__4080);
  not g__1873(w__19 ,w__3943);
  not g__1874(w__18 ,w__4081);
  not g__1875(w__17 ,w__4063);
  not g__1876(w__16 ,w__4039);
  not g__1877(w__15 ,w__3933);
  not g__1878(w__14 ,w__4066);
  not g__1879(w__13 ,w__4070);
  not g__1880(w__12 ,w__4009);
  not g__1881(w__11 ,w__3995);
  not g__1882(w__10 ,w__3937);
  not g__1883(w__9 ,w__4017);
  not g__1884(w__8 ,w__3954);
  not g__1885(w__7 ,w__4043);
  not g__1886(w__6 ,w__4002);
  not g__1887(w__3 ,w__5);
  not g__1888(w__5 ,w__413);
  not g__1889(w__4 ,w__410);
  xor g__1890(out1[8] ,w__1164 ,w__1129);
  xor g__1891(w__2 ,w__590 ,w__594);
  and g__1892(w__1 ,w__4 ,w__397);
  xnor g__1893(w__4412 ,w__1622 ,w__1639);
  or g__1894(w__4378 ,w__1638 ,w__1640);
  xnor g__1895(w__4411 ,w__1634 ,w__1635);
  nor g__1896(w__1640 ,w__1622 ,w__1637);
  or g__1897(w__4410 ,w__1630 ,w__1636);
  xnor g__1898(w__1639 ,w__1586 ,w__1628);
  xnor g__1899(w__4413 ,w__1613 ,w__1625);
  xnor g__1900(w__4414 ,w__1615 ,w__1624);
  xor g__1901(w__4377 ,w__1621 ,w__1623);
  or g__1902(w__4380 ,w__1619 ,w__1632);
  nor g__1903(w__1638 ,w__1586 ,w__1629);
  or g__1904(w__4409 ,w__1620 ,w__1631);
  and g__1905(w__1637 ,w__1586 ,w__1629);
  and g__1906(w__1636 ,w__1634 ,w__1626);
  or g__1907(w__4379 ,w__1608 ,w__1633);
  or g__1908(w__4381 ,w__1602 ,w__1627);
  xnor g__1909(w__4415 ,w__1614 ,w__1607);
  xnor g__1910(w__1635 ,w__1612 ,w__1588);
  and g__1911(w__1633 ,w__1618 ,w__1613);
  and g__1912(w__1632 ,w__1617 ,w__1615);
  or g__1913(w__4382 ,w__1567 ,w__1616);
  nor g__1914(w__1631 ,w__1610 ,w__1621);
  nor g__1915(w__1630 ,w__1588 ,w__1612);
  or g__1916(w__1634 ,w__1548 ,w__1609);
  not g__1917(w__1629 ,w__1628);
  nor g__1918(w__1627 ,w__1603 ,w__1614);
  or g__1919(w__1626 ,w__1587 ,w__1611);
  xnor g__1920(w__4416 ,w__1599 ,w__1574);
  xnor g__1921(w__1625 ,w__1595 ,w__1592);
  xnor g__1922(w__1624 ,w__1597 ,w__1606);
  xnor g__1923(w__1623 ,w__1593 ,w__1568);
  xnor g__1924(w__1628 ,w__1598 ,w__1572);
  nor g__1925(w__1620 ,w__1568 ,w__1593);
  nor g__1926(w__1619 ,w__1606 ,w__1597);
  or g__1927(w__1618 ,w__1291 ,w__1594);
  or g__1928(w__1617 ,w__1605 ,w__1596);
  or g__1929(w__4408 ,w__1552 ,w__1591);
  nor g__1930(w__1616 ,w__1558 ,w__1599);
  or g__1931(w__4383 ,w__1557 ,w__1600);
  and g__1932(w__1622 ,w__1559 ,w__1601);
  and g__1933(w__1621 ,w__1584 ,w__1604);
  not g__1934(w__1611 ,w__1612);
  and g__1935(w__1610 ,w__1568 ,w__1593);
  and g__1936(w__1609 ,w__1547 ,w__1598);
  nor g__1937(w__1608 ,w__1287 ,w__1595);
  xor g__1938(w__4376 ,w__1589 ,w__1570);
  xnor g__1939(w__4417 ,w__1580 ,w__1576);
  xnor g__1940(w__1607 ,w__1585 ,w__1578);
  xnor g__1941(w__1615 ,w__1569 ,w__1577);
  xnor g__1942(w__1614 ,w__1497 ,w__1571);
  xnor g__1943(w__1613 ,w__1590 ,w__1573);
  xnor g__1944(w__1612 ,w__1554 ,w__1575);
  not g__1945(w__1606 ,w__1605);
  or g__1946(w__1604 ,w__1498 ,w__1581);
  and g__1947(w__1603 ,w__1585 ,w__1579);
  nor g__1948(w__1602 ,w__1585 ,w__1579);
  or g__1949(w__1601 ,w__1555 ,w__1590);
  and g__1950(w__1600 ,w__1556 ,w__1580);
  or g__1951(w__1605 ,w__1563 ,w__1582);
  not g__1952(w__1596 ,w__1597);
  not g__1953(w__1594 ,w__1595);
  nor g__1954(w__1591 ,w__1551 ,w__1589);
  xnor g__1955(w__1599 ,w__1523 ,w__1545);
  xnor g__1956(w__1598 ,w__1519 ,w__1544);
  xnor g__1957(w__1597 ,w__1520 ,w__1546);
  and g__1958(w__1595 ,w__1553 ,w__1583);
  xnor g__1959(w__1593 ,w__1518 ,w__1543);
  xnor g__1960(w__1592 ,w__1521 ,w__1542);
  not g__1961(w__1587 ,w__1588);
  or g__1962(w__1584 ,w__1507 ,w__1554);
  or g__1963(w__1583 ,w__1569 ,w__1565);
  nor g__1964(w__1582 ,w__1497 ,w__1562);
  and g__1965(w__1581 ,w__1507 ,w__1554);
  or g__1966(w__4384 ,w__1478 ,w__1560);
  and g__1967(w__1590 ,w__1530 ,w__1550);
  and g__1968(w__1589 ,w__1528 ,w__1566);
  and g__1969(w__1588 ,w__1526 ,w__1549);
  and g__1970(w__1586 ,w__1537 ,w__1564);
  and g__1971(w__1585 ,w__1534 ,w__1561);
  not g__1972(w__1579 ,w__1578);
  xnor g__1973(w__4418 ,w__1522 ,w__1524);
  xnor g__1974(w__1577 ,w__1506 ,w__1503);
  xnor g__1975(w__1576 ,w__1513 ,w__1484);
  xnor g__1976(w__1575 ,w__1507 ,w__1498);
  xnor g__1977(w__1574 ,w__1539 ,w__1516);
  xnor g__1978(w__1573 ,w__1486 ,w__1511);
  xnor g__1979(w__1572 ,w__1515 ,w__1541);
  xnor g__1980(w__1571 ,w__1509 ,w__1508);
  xnor g__1981(w__1570 ,w__1504 ,w__1481);
  xnor g__1982(w__1580 ,w__1434 ,w__1501);
  xnor g__1983(w__1578 ,w__1499 ,w__1525);
  nor g__1984(w__1567 ,w__1539 ,w__1517);
  or g__1985(w__1566 ,w__1532 ,w__1518);
  nor g__1986(w__1565 ,w__1505 ,w__1503);
  or g__1987(w__1564 ,w__1521 ,w__1536);
  nor g__1988(w__1563 ,w__1508 ,w__1509);
  and g__1989(w__1562 ,w__1508 ,w__1509);
  or g__1990(w__1561 ,w__1533 ,w__1523);
  nor g__1991(w__1560 ,w__1489 ,w__1522);
  or g__1992(w__1559 ,w__1485 ,w__1511);
  and g__1993(w__1558 ,w__1539 ,w__1517);
  nor g__1994(w__1557 ,w__1484 ,w__1513);
  or g__1995(w__1556 ,w__1483 ,w__1512);
  nor g__1996(w__1555 ,w__1486 ,w__1510);
  and g__1997(w__1569 ,w__1477 ,w__1529);
  and g__1998(w__1568 ,w__1430 ,w__1538);
  or g__1999(w__1553 ,w__1506 ,w__1502);
  nor g__2000(w__1552 ,w__1481 ,w__1504);
  and g__2001(w__1551 ,w__1481 ,w__1504);
  or g__2002(w__1550 ,w__1520 ,w__1535);
  or g__2003(w__1549 ,w__1531 ,w__1519);
  nor g__2004(w__1548 ,w__1541 ,w__1515);
  or g__2005(w__1547 ,w__1540 ,w__1514);
  or g__2006(w__4407 ,w__1394 ,w__1527);
  xor g__2007(w__4375 ,w__1488 ,w__1448);
  xnor g__2008(w__1546 ,w__1487 ,w__1479);
  xnor g__2009(w__1545 ,w__1494 ,w__1192);
  xnor g__2010(w__1544 ,w__1410 ,w__1496);
  xnor g__2011(w__1543 ,w__1349 ,w__1482);
  xnor g__2012(w__1542 ,w__1493 ,w__1480);
  xnor g__2013(w__1554 ,w__1500 ,w__1449);
  not g__2014(w__1540 ,w__1541);
  or g__2015(w__1538 ,w__1392 ,w__1500);
  or g__2016(w__1537 ,w__1480 ,w__1493);
  and g__2017(w__1536 ,w__1480 ,w__1493);
  and g__2018(w__1535 ,w__1479 ,w__1487);
  or g__2019(w__1534 ,w__1192 ,w__1494);
  and g__2020(w__1533 ,w__1192 ,w__1494);
  and g__2021(w__1532 ,w__1349 ,w__1482);
  nor g__2022(w__1531 ,w__1410 ,w__1495);
  or g__2023(w__1530 ,w__1479 ,w__1487);
  or g__2024(w__1529 ,w__1499 ,w__1490);
  or g__2025(w__4385 ,w__1393 ,w__1476);
  or g__2026(w__1528 ,w__1349 ,w__1482);
  nor g__2027(w__1527 ,w__1408 ,w__1488);
  or g__2028(w__1526 ,w__1409 ,w__1496);
  xnor g__2029(w__1525 ,w__1432 ,w__1475);
  xnor g__2030(w__1524 ,w__1411 ,w__1193);
  and g__2031(w__1541 ,w__1415 ,w__1491);
  and g__2032(w__1539 ,w__1466 ,w__1492);
  not g__2033(w__1517 ,w__1516);
  not g__2034(w__1514 ,w__1515);
  not g__2035(w__1512 ,w__1513);
  not g__2036(w__1510 ,w__1511);
  not g__2037(w__1505 ,w__1506);
  not g__2038(w__1502 ,w__1503);
  xor g__2039(w__4419 ,w__1195 ,w__1455);
  xnor g__2040(w__1501 ,w__1328 ,w__1196);
  xnor g__2041(w__1523 ,w__1373 ,w__1456);
  xnor g__2042(w__1522 ,w__1379 ,w__1438);
  xnor g__2043(w__1521 ,w__1381 ,w__1452);
  xnor g__2044(w__1520 ,w__1362 ,w__1447);
  xnor g__2045(w__1519 ,w__1355 ,w__1445);
  xnor g__2046(w__1518 ,w__1352 ,w__1444);
  xnor g__2047(w__1516 ,w__1435 ,w__1441);
  xnor g__2048(w__1515 ,w__1330 ,w__1454);
  xnor g__2049(w__1513 ,w__1335 ,w__1440);
  xnor g__2050(w__1511 ,w__1194 ,w__1439);
  xnor g__2051(w__1509 ,w__1325 ,w__1450);
  xnor g__2052(w__1508 ,w__1315 ,w__1451);
  xnor g__2053(w__1507 ,w__1350 ,w__1453);
  xnor g__2054(w__1506 ,w__1380 ,w__1446);
  xnor g__2055(w__1504 ,w__1354 ,w__1442);
  xnor g__2056(w__1503 ,w__1437 ,w__1443);
  not g__2057(w__1495 ,w__1496);
  or g__2058(w__1492 ,w__1473 ,w__1196);
  or g__2059(w__1491 ,w__1422 ,w__1194);
  nor g__2060(w__1490 ,w__1432 ,w__1474);
  and g__2061(w__1489 ,w__1412 ,w__1193);
  and g__2062(w__1500 ,w__1420 ,w__1472);
  and g__2063(w__1499 ,w__1427 ,w__1464);
  and g__2064(w__1498 ,w__1421 ,w__1462);
  and g__2065(w__1497 ,w__1407 ,w__1470);
  and g__2066(w__1496 ,w__1402 ,w__1465);
  and g__2067(w__1494 ,w__1404 ,w__1468);
  and g__2068(w__1493 ,w__1425 ,w__1457);
  not g__2069(w__1485 ,w__1486);
  not g__2070(w__1483 ,w__1484);
  nor g__2071(w__1478 ,w__1412 ,w__1193);
  or g__2072(w__1477 ,w__1431 ,w__1475);
  nor g__2073(w__1476 ,w__1418 ,w__1195);
  and g__2074(w__1488 ,w__1395 ,w__1469);
  and g__2075(w__1487 ,w__1390 ,w__1463);
  or g__2076(w__1486 ,w__1414 ,w__1461);
  and g__2077(w__1484 ,w__1400 ,w__1460);
  and g__2078(w__1482 ,w__1399 ,w__1471);
  and g__2079(w__1481 ,w__1391 ,w__1458);
  and g__2080(w__1480 ,w__1416 ,w__1467);
  and g__2081(w__1479 ,w__1423 ,w__1459);
  not g__2082(w__1474 ,w__1475);
  nor g__2083(w__1473 ,w__1327 ,w__1434);
  or g__2084(w__1472 ,w__1346 ,w__1405);
  or g__2085(w__1471 ,w__1345 ,w__1417);
  or g__2086(w__1470 ,w__1428 ,w__1436);
  or g__2087(w__1469 ,w__1338 ,w__1401);
  or g__2088(w__1468 ,w__1335 ,w__1406);
  or g__2089(w__1467 ,w__1380 ,w__1403);
  or g__2090(w__1466 ,w__1328 ,w__1433);
  or g__2091(w__1465 ,w__1381 ,w__1429);
  or g__2092(w__1464 ,w__1373 ,w__1424);
  or g__2093(w__1463 ,w__1343 ,w__1413);
  or g__2094(w__1462 ,w__1336 ,w__1397);
  and g__2095(w__1461 ,w__1419 ,w__1437);
  or g__2096(w__1460 ,w__1379 ,w__1396);
  or g__2097(w__1459 ,w__1382 ,w__1398);
  or g__2098(w__1458 ,w__1337 ,w__1389);
  xor g__2099(w__4420 ,w__1347 ,w__1387);
  or g__2100(w__1457 ,w__1376 ,w__1426);
  xnor g__2101(w__1456 ,w__1366 ,w__1369);
  xnor g__2102(w__1455 ,w__1351 ,w__1363);
  xnor g__2103(w__1475 ,w__1383 ,w__1371);
  xnor g__2104(w__1454 ,w__1324 ,w__1336);
  xnor g__2105(w__1453 ,w__1329 ,w__1345);
  xnor g__2106(w__1452 ,w__1326 ,w__1357);
  xnor g__2107(w__1451 ,w__1323 ,w__1343);
  xnor g__2108(w__1450 ,w__1318 ,w__1382);
  xnor g__2109(w__1449 ,w__1316 ,w__1321);
  xnor g__2110(w__1448 ,w__1370 ,w__1364);
  xnor g__2111(w__1447 ,w__1322 ,w__1376);
  xnor g__2112(w__1446 ,w__1320 ,w__1358);
  xnor g__2113(w__1445 ,w__1368 ,w__1346);
  xnor g__2114(w__1444 ,w__1367 ,w__1337);
  xnor g__2115(w__1443 ,w__1314 ,w__1332);
  xnor g__2116(w__1442 ,w__1319 ,w__1338);
  xnor g__2117(w__1441 ,w__1348 ,w__1356);
  xnor g__2118(w__1440 ,w__1353 ,w__1361);
  xnor g__2119(w__1439 ,w__1317 ,w__1360);
  xnor g__2120(w__1438 ,w__1365 ,w__1359);
  not g__2121(w__1436 ,w__1435);
  not g__2122(w__1433 ,w__1434);
  not g__2123(w__1431 ,w__1432);
  or g__2124(w__1430 ,w__1316 ,w__1321);
  and g__2125(w__1429 ,w__1326 ,w__1357);
  and g__2126(w__1428 ,w__1348 ,w__1356);
  or g__2127(w__1427 ,w__1366 ,w__1369);
  and g__2128(w__1426 ,w__1362 ,w__1322);
  or g__2129(w__1425 ,w__1362 ,w__1322);
  and g__2130(w__1424 ,w__1366 ,w__1369);
  or g__2131(w__1423 ,w__1325 ,w__1318);
  and g__2132(w__1422 ,w__1317 ,w__1360);
  or g__2133(w__1421 ,w__1330 ,w__1324);
  or g__2134(w__1420 ,w__1355 ,w__1368);
  or g__2135(w__1419 ,w__1313 ,w__1331);
  and g__2136(w__1418 ,w__1351 ,w__1363);
  and g__2137(w__1417 ,w__1350 ,w__1329);
  or g__2138(w__1416 ,w__1320 ,w__1358);
  or g__2139(w__1415 ,w__1317 ,w__1360);
  nor g__2140(w__1414 ,w__1314 ,w__1332);
  and g__2141(w__1413 ,w__1323 ,w__1315);
  and g__2142(w__1437 ,w__1384 ,w__1372);
  and g__2143(w__1435 ,w__1333 ,w__1344);
  and g__2144(w__1434 ,w__1378 ,w__1340);
  and g__2145(w__1432 ,w__1375 ,w__1334);
  not g__2146(w__1412 ,w__1411);
  not g__2147(w__1409 ,w__1410);
  and g__2148(w__1408 ,w__1370 ,w__1364);
  or g__2149(w__1407 ,w__1348 ,w__1356);
  and g__2150(w__1406 ,w__1353 ,w__1361);
  and g__2151(w__1405 ,w__1355 ,w__1368);
  or g__2152(w__1404 ,w__1353 ,w__1361);
  and g__2153(w__1403 ,w__1320 ,w__1358);
  or g__2154(w__1402 ,w__1326 ,w__1357);
  and g__2155(w__1401 ,w__1354 ,w__1319);
  or g__2156(w__1400 ,w__1365 ,w__1359);
  or g__2157(w__1399 ,w__1350 ,w__1329);
  and g__2158(w__1398 ,w__1325 ,w__1318);
  and g__2159(w__1397 ,w__1330 ,w__1324);
  and g__2160(w__1396 ,w__1365 ,w__1359);
  or g__2161(w__1395 ,w__1354 ,w__1319);
  nor g__2162(w__1394 ,w__1370 ,w__1364);
  nor g__2163(w__1393 ,w__1351 ,w__1363);
  and g__2164(w__1392 ,w__1316 ,w__1321);
  or g__2165(w__1391 ,w__1352 ,w__1367);
  or g__2166(w__1390 ,w__1323 ,w__1315);
  and g__2167(w__1389 ,w__1352 ,w__1367);
  nor g__2168(w__1388 ,w__1387 ,w__1347);
  and g__2169(w__1411 ,w__1386 ,w__1342);
  and g__2170(w__1410 ,w__1341 ,w__1339);
  not g__2171(w__1386 ,w__1385);
  not g__2172(w__1384 ,w__1383);
  not g__2173(w__1378 ,w__1377);
  not g__2174(w__1375 ,w__1374);
  not g__2175(w__1372 ,w__1371);
  and g__2176(w__4374 ,in1[8] ,in2[7]);
  or g__2177(w__1387 ,w__1209 ,w__1302);
  or g__2178(w__1385 ,w__1249 ,w__1229);
  or g__2179(w__1383 ,w__1204 ,w__1272);
  or g__2180(w__1382 ,w__1211 ,w__1239);
  or g__2181(w__1381 ,w__1243 ,w__1254);
  or g__2182(w__1380 ,w__1243 ,w__1233);
  or g__2183(w__1379 ,w__1249 ,w__1234);
  or g__2184(w__1377 ,w__1223 ,w__1272);
  or g__2185(w__1376 ,w__1219 ,w__1230);
  or g__2186(w__1374 ,w__1261 ,w__1229);
  or g__2187(w__1373 ,w__1221 ,w__1240);
  or g__2188(w__1371 ,w__1225 ,w__1230);
  or g__2189(w__1370 ,w__1258 ,w__1269);
  or g__2190(w__1369 ,w__1214 ,w__1201);
  or g__2191(w__1368 ,w__1217 ,w__1251);
  or g__2192(w__1367 ,w__1258 ,w__1227);
  or g__2193(w__1366 ,w__1307 ,w__1263);
  or g__2194(w__1365 ,w__1231 ,w__1198);
  or g__2195(w__1364 ,w__1207 ,w__1245);
  or g__2196(w__1363 ,w__1279 ,w__1233);
  or g__2197(w__1362 ,w__1261 ,w__1286);
  or g__2198(w__1361 ,w__1248 ,w__1255);
  or g__2199(w__1360 ,w__1213 ,w__1246);
  or g__2200(w__1359 ,w__1276 ,w__1202);
  or g__2201(w__1358 ,w__1216 ,w__1284);
  or g__2202(w__1357 ,w__1300 ,w__1264);
  or g__2203(w__1356 ,w__1275 ,w__1237);
  or g__2204(w__1355 ,w__1299 ,w__1266);
  or g__2205(w__1354 ,w__1308 ,w__1267);
  or g__2206(w__1353 ,w__1278 ,w__1199);
  or g__2207(w__1352 ,w__1260 ,w__1270);
  or g__2208(w__1351 ,w__1281 ,w__1254);
  or g__2209(w__1350 ,w__1211 ,w__1252);
  or g__2210(w__1349 ,w__1242 ,w__1245);
  or g__2211(w__1348 ,w__1281 ,w__1251);
  not g__2212(w__1332 ,w__1331);
  not g__2213(w__1328 ,w__1327);
  not g__2214(w__1314 ,w__1313);
  nor g__2215(w__1312 ,w__1276 ,w__1184);
  nor g__2216(w__1311 ,w__1279 ,w__1186);
  nor g__2217(w__1310 ,w__1302 ,w__1188);
  nor g__2218(w__1309 ,w__1282 ,w__1273);
  or g__2219(w__1347 ,w__1231 ,w__1239);
  or g__2220(w__1346 ,w__1204 ,w__1263);
  or g__2221(w__1345 ,w__1206 ,w__1286);
  and g__2222(w__1344 ,in1[5] ,in2[0]);
  or g__2223(w__1343 ,w__1305 ,w__1255);
  and g__2224(w__1342 ,in1[3] ,in2[0]);
  and g__2225(w__1341 ,in1[7] ,in2[2]);
  and g__2226(w__1340 ,in1[4] ,in2[0]);
  and g__2227(w__1339 ,in1[8] ,in2[1]);
  or g__2228(w__1338 ,w__1304 ,w__1237);
  or g__2229(w__1337 ,w__1207 ,w__1284);
  or g__2230(w__1336 ,w__1219 ,w__1234);
  or g__2231(w__1335 ,w__1214 ,w__1240);
  and g__2232(w__1334 ,in1[6] ,in2[0]);
  and g__2233(w__1333 ,in1[4] ,in2[1]);
  and g__2234(w__1331 ,in1[3] ,in2[5]);
  or g__2235(w__1330 ,w__1260 ,w__1294);
  or g__2236(w__1329 ,w__1297 ,w__1264);
  and g__2237(w__1327 ,in1[0] ,in2[5]);
  or g__2238(w__1326 ,w__1217 ,w__1236);
  or g__2239(w__1325 ,w__1275 ,w__1246);
  or g__2240(w__1324 ,w__1257 ,w__1202);
  or g__2241(w__1323 ,w__1282 ,w__1266);
  or g__2242(w__1322 ,w__1225 ,w__1273);
  or g__2243(w__1321 ,w__1242 ,w__1227);
  or g__2244(w__1320 ,w__1278 ,w__1269);
  or g__2245(w__1319 ,w__1257 ,w__1252);
  or g__2246(w__1318 ,w__1209 ,w__1236);
  or g__2247(w__1317 ,w__1248 ,w__1267);
  or g__2248(w__1316 ,w__1221 ,w__1270);
  or g__2249(w__1315 ,w__1223 ,w__1199);
  and g__2250(w__1313 ,in1[2] ,in2[6]);
  not g__2251(w__1308 ,in1[6]);
  not g__2252(w__1307 ,in1[2]);
  not g__2253(w__1306 ,in1[1]);
  not g__2254(w__1305 ,in1[4]);
  not g__2255(w__1304 ,in1[8]);
  not g__2256(w__1303 ,in2[3]);
  not g__2257(w__1302 ,in2[0]);
  not g__2258(w__1301 ,in2[1]);
  not g__2259(w__1300 ,in1[5]);
  not g__2260(w__1299 ,in1[3]);
  not g__2261(w__1298 ,in1[0]);
  not g__2262(w__1297 ,in1[7]);
  not g__2263(w__1296 ,in2[4]);
  not g__2264(w__1295 ,in2[2]);
  not g__2265(w__1294 ,in2[5]);
  not g__2266(w__1293 ,in2[7]);
  not g__2267(w__1292 ,in2[6]);
  not g__2268(w__1191 ,w__1290);
  not g__2269(w__1290 ,w__1298);
  not g__2270(w__1190 ,w__1289);
  not g__2271(w__1183 ,w__1289);
  not g__2272(w__1289 ,w__1301);
  not g__2273(w__1189 ,w__1288);
  not g__2274(w__1288 ,w__1302);
  buf g__2275(w__4387 ,w__1312);
  buf g__2276(w__4421 ,w__1309);
  buf g__2277(w__4389 ,w__1310);
  buf g__2278(w__4388 ,w__1311);
  buf g__2279(w__4386 ,w__1388);
  not g__2280(w__1287 ,w__1291);
  not g__2281(w__1291 ,w__1592);
  not g__2282(w__1286 ,w__1285);
  not g__2283(w__1285 ,w__1303);
  not g__2284(w__1284 ,w__1283);
  not g__2285(w__1283 ,w__1296);
  not g__2286(w__1282 ,w__1280);
  not g__2287(w__1281 ,w__1280);
  not g__2288(w__1280 ,w__1298);
  not g__2289(w__1279 ,w__1277);
  not g__2290(w__1278 ,w__1277);
  not g__2291(w__1277 ,w__1306);
  not g__2292(w__1276 ,w__1274);
  not g__2293(w__1275 ,w__1274);
  not g__2294(w__1274 ,w__1306);
  not g__2295(w__1273 ,w__1271);
  not g__2296(w__1272 ,w__1271);
  not g__2297(w__1271 ,w__1190);
  not g__2298(w__1270 ,w__1268);
  not g__2299(w__1269 ,w__1268);
  not g__2300(w__1268 ,w__1293);
  not g__2301(w__1267 ,w__1265);
  not g__2302(w__1266 ,w__1265);
  not g__2303(w__1265 ,w__1293);
  not g__2304(w__1264 ,w__1262);
  not g__2305(w__1263 ,w__1262);
  not g__2306(w__1262 ,w__1296);
  not g__2307(w__1261 ,w__1259);
  not g__2308(w__1260 ,w__1259);
  not g__2309(w__1259 ,w__1300);
  not g__2310(w__1258 ,w__1256);
  not g__2311(w__1257 ,w__1256);
  not g__2312(w__1256 ,w__1297);
  not g__2313(w__1255 ,w__1253);
  not g__2314(w__1254 ,w__1253);
  not g__2315(w__1253 ,w__1303);
  not g__2316(w__1252 ,w__1250);
  not g__2317(w__1251 ,w__1250);
  not g__2318(w__1250 ,w__1292);
  not g__2319(w__1249 ,w__1247);
  not g__2320(w__1248 ,w__1247);
  not g__2321(w__1247 ,w__1307);
  not g__2322(w__1246 ,w__1244);
  not g__2323(w__1245 ,w__1244);
  not g__2324(w__1244 ,w__1292);
  not g__2325(w__1243 ,w__1241);
  not g__2326(w__1242 ,w__1241);
  not g__2327(w__1241 ,w__1308);
  not g__2328(w__1240 ,w__1238);
  not g__2329(w__1239 ,w__1238);
  not g__2330(w__1238 ,w__1295);
  not g__2331(w__1237 ,w__1235);
  not g__2332(w__1236 ,w__1235);
  not g__2333(w__1235 ,w__1294);
  not g__2334(w__1234 ,w__1232);
  not g__2335(w__1233 ,w__1232);
  not g__2336(w__1232 ,w__1295);
  not g__2337(w__1188 ,w__1187);
  not g__2338(w__1231 ,w__1187);
  not g__2339(w__1187 ,w__1191);
  not g__2340(w__1186 ,w__1185);
  not g__2341(w__1230 ,w__1185);
  not g__2342(w__1185 ,w__1189);
  not g__2343(w__1184 ,w__1228);
  not g__2344(w__1229 ,w__1228);
  not g__2345(w__1228 ,w__1183);
  not g__2346(w__1227 ,w__1226);
  not g__2347(w__1226 ,w__1294);
  not g__2348(w__1225 ,w__1224);
  not g__2349(w__1224 ,w__1297);
  not g__2350(w__1223 ,w__1222);
  not g__2351(w__1222 ,w__1299);
  not g__2352(w__1221 ,w__1220);
  not g__2353(w__1220 ,w__1305);
  not g__2354(w__1219 ,w__1218);
  not g__2355(w__1218 ,w__1304);
  not g__2356(w__1217 ,w__1215);
  not g__2357(w__1216 ,w__1215);
  not g__2358(w__1215 ,w__1305);
  not g__2359(w__1214 ,w__1212);
  not g__2360(w__1213 ,w__1212);
  not g__2361(w__1212 ,w__1299);
  not g__2362(w__1211 ,w__1210);
  not g__2363(w__1210 ,w__1300);
  not g__2364(w__1209 ,w__1208);
  not g__2365(w__1208 ,w__1307);
  not g__2366(w__1207 ,w__1205);
  not g__2367(w__1206 ,w__1205);
  not g__2368(w__1205 ,w__1304);
  not g__2369(w__1204 ,w__1203);
  not g__2370(w__1203 ,w__1308);
  not g__2371(w__1202 ,w__1200);
  not g__2372(w__1201 ,w__1200);
  not g__2373(w__1200 ,w__1303);
  not g__2374(w__1199 ,w__1197);
  not g__2375(w__1198 ,w__1197);
  not g__2376(w__1197 ,w__1296);
  xnor g__2377(w__1196 ,w__1333 ,w__1344);
  xor g__2378(w__1195 ,w__1385 ,w__1342);
  xnor g__2379(w__1194 ,w__1341 ,w__1339);
  xor g__2380(w__1193 ,w__1377 ,w__1340);
  xor g__2381(w__1192 ,w__1374 ,w__1334);
  xnor g__2382(w__4476 ,w__2080 ,w__2097);
  or g__2383(w__4442 ,w__2096 ,w__2098);
  xnor g__2384(w__4475 ,w__2092 ,w__2093);
  nor g__2385(w__2098 ,w__2080 ,w__2095);
  or g__2386(w__4474 ,w__2088 ,w__2094);
  xnor g__2387(w__2097 ,w__2044 ,w__2086);
  xnor g__2388(w__4477 ,w__2071 ,w__2083);
  xnor g__2389(w__4478 ,w__2073 ,w__2082);
  xor g__2390(w__4441 ,w__2079 ,w__2081);
  or g__2391(w__4444 ,w__2077 ,w__2090);
  nor g__2392(w__2096 ,w__2044 ,w__2087);
  or g__2393(w__4473 ,w__2078 ,w__2089);
  and g__2394(w__2095 ,w__2044 ,w__2087);
  and g__2395(w__2094 ,w__2092 ,w__2084);
  or g__2396(w__4443 ,w__2066 ,w__2091);
  or g__2397(w__4445 ,w__2060 ,w__2085);
  xnor g__2398(w__4479 ,w__2072 ,w__2065);
  xnor g__2399(w__2093 ,w__2070 ,w__2046);
  and g__2400(w__2091 ,w__2076 ,w__2071);
  and g__2401(w__2090 ,w__2075 ,w__2073);
  or g__2402(w__4446 ,w__2025 ,w__2074);
  nor g__2403(w__2089 ,w__2068 ,w__2079);
  nor g__2404(w__2088 ,w__2046 ,w__2070);
  or g__2405(w__2092 ,w__2006 ,w__2067);
  not g__2406(w__2087 ,w__2086);
  nor g__2407(w__2085 ,w__2061 ,w__2072);
  or g__2408(w__2084 ,w__2045 ,w__2069);
  xnor g__2409(w__4480 ,w__2057 ,w__2032);
  xnor g__2410(w__2083 ,w__2053 ,w__2050);
  xnor g__2411(w__2082 ,w__2055 ,w__2064);
  xnor g__2412(w__2081 ,w__2051 ,w__2026);
  xnor g__2413(w__2086 ,w__2056 ,w__2030);
  nor g__2414(w__2078 ,w__2026 ,w__2051);
  nor g__2415(w__2077 ,w__2064 ,w__2055);
  or g__2416(w__2076 ,w__1749 ,w__2052);
  or g__2417(w__2075 ,w__2063 ,w__2054);
  or g__2418(w__4472 ,w__2010 ,w__2049);
  nor g__2419(w__2074 ,w__2016 ,w__2057);
  or g__2420(w__4447 ,w__2015 ,w__2058);
  and g__2421(w__2080 ,w__2017 ,w__2059);
  and g__2422(w__2079 ,w__2042 ,w__2062);
  not g__2423(w__2069 ,w__2070);
  and g__2424(w__2068 ,w__2026 ,w__2051);
  and g__2425(w__2067 ,w__2005 ,w__2056);
  nor g__2426(w__2066 ,w__1745 ,w__2053);
  xor g__2427(w__4440 ,w__2047 ,w__2028);
  xnor g__2428(w__4481 ,w__2038 ,w__2034);
  xnor g__2429(w__2065 ,w__2043 ,w__2036);
  xnor g__2430(w__2073 ,w__2027 ,w__2035);
  xnor g__2431(w__2072 ,w__1955 ,w__2029);
  xnor g__2432(w__2071 ,w__2048 ,w__2031);
  xnor g__2433(w__2070 ,w__2012 ,w__2033);
  not g__2434(w__2064 ,w__2063);
  or g__2435(w__2062 ,w__1956 ,w__2039);
  and g__2436(w__2061 ,w__2043 ,w__2037);
  nor g__2437(w__2060 ,w__2043 ,w__2037);
  or g__2438(w__2059 ,w__2013 ,w__2048);
  and g__2439(w__2058 ,w__2014 ,w__2038);
  or g__2440(w__2063 ,w__2021 ,w__2040);
  not g__2441(w__2054 ,w__2055);
  not g__2442(w__2052 ,w__2053);
  nor g__2443(w__2049 ,w__2009 ,w__2047);
  xnor g__2444(w__2057 ,w__1981 ,w__2003);
  xnor g__2445(w__2056 ,w__1977 ,w__2002);
  xnor g__2446(w__2055 ,w__1978 ,w__2004);
  and g__2447(w__2053 ,w__2011 ,w__2041);
  xnor g__2448(w__2051 ,w__1976 ,w__2001);
  xnor g__2449(w__2050 ,w__1979 ,w__2000);
  not g__2450(w__2045 ,w__2046);
  or g__2451(w__2042 ,w__1965 ,w__2012);
  or g__2452(w__2041 ,w__2027 ,w__2023);
  nor g__2453(w__2040 ,w__1955 ,w__2020);
  and g__2454(w__2039 ,w__1965 ,w__2012);
  or g__2455(w__4448 ,w__1936 ,w__2018);
  and g__2456(w__2048 ,w__1988 ,w__2008);
  and g__2457(w__2047 ,w__1986 ,w__2024);
  and g__2458(w__2046 ,w__1984 ,w__2007);
  and g__2459(w__2044 ,w__1995 ,w__2022);
  and g__2460(w__2043 ,w__1992 ,w__2019);
  not g__2461(w__2037 ,w__2036);
  xnor g__2462(w__4482 ,w__1980 ,w__1982);
  xnor g__2463(w__2035 ,w__1964 ,w__1961);
  xnor g__2464(w__2034 ,w__1971 ,w__1942);
  xnor g__2465(w__2033 ,w__1965 ,w__1956);
  xnor g__2466(w__2032 ,w__1997 ,w__1974);
  xnor g__2467(w__2031 ,w__1944 ,w__1969);
  xnor g__2468(w__2030 ,w__1973 ,w__1999);
  xnor g__2469(w__2029 ,w__1967 ,w__1966);
  xnor g__2470(w__2028 ,w__1962 ,w__1939);
  xnor g__2471(w__2038 ,w__1892 ,w__1959);
  xnor g__2472(w__2036 ,w__1957 ,w__1983);
  nor g__2473(w__2025 ,w__1997 ,w__1975);
  or g__2474(w__2024 ,w__1990 ,w__1976);
  nor g__2475(w__2023 ,w__1963 ,w__1961);
  or g__2476(w__2022 ,w__1979 ,w__1994);
  nor g__2477(w__2021 ,w__1966 ,w__1967);
  and g__2478(w__2020 ,w__1966 ,w__1967);
  or g__2479(w__2019 ,w__1991 ,w__1981);
  nor g__2480(w__2018 ,w__1947 ,w__1980);
  or g__2481(w__2017 ,w__1943 ,w__1969);
  and g__2482(w__2016 ,w__1997 ,w__1975);
  nor g__2483(w__2015 ,w__1942 ,w__1971);
  or g__2484(w__2014 ,w__1941 ,w__1970);
  nor g__2485(w__2013 ,w__1944 ,w__1968);
  and g__2486(w__2027 ,w__1935 ,w__1987);
  and g__2487(w__2026 ,w__1888 ,w__1996);
  or g__2488(w__2011 ,w__1964 ,w__1960);
  nor g__2489(w__2010 ,w__1939 ,w__1962);
  and g__2490(w__2009 ,w__1939 ,w__1962);
  or g__2491(w__2008 ,w__1978 ,w__1993);
  or g__2492(w__2007 ,w__1989 ,w__1977);
  nor g__2493(w__2006 ,w__1999 ,w__1973);
  or g__2494(w__2005 ,w__1998 ,w__1972);
  or g__2495(w__4471 ,w__1852 ,w__1985);
  xor g__2496(w__4439 ,w__1946 ,w__1906);
  xnor g__2497(w__2004 ,w__1945 ,w__1937);
  xnor g__2498(w__2003 ,w__1952 ,w__1650);
  xnor g__2499(w__2002 ,w__1868 ,w__1954);
  xnor g__2500(w__2001 ,w__1807 ,w__1940);
  xnor g__2501(w__2000 ,w__1951 ,w__1938);
  xnor g__2502(w__2012 ,w__1958 ,w__1907);
  not g__2503(w__1998 ,w__1999);
  or g__2504(w__1996 ,w__1850 ,w__1958);
  or g__2505(w__1995 ,w__1938 ,w__1951);
  and g__2506(w__1994 ,w__1938 ,w__1951);
  and g__2507(w__1993 ,w__1937 ,w__1945);
  or g__2508(w__1992 ,w__1650 ,w__1952);
  and g__2509(w__1991 ,w__1650 ,w__1952);
  and g__2510(w__1990 ,w__1807 ,w__1940);
  nor g__2511(w__1989 ,w__1868 ,w__1953);
  or g__2512(w__1988 ,w__1937 ,w__1945);
  or g__2513(w__1987 ,w__1957 ,w__1948);
  or g__2514(w__4449 ,w__1851 ,w__1934);
  or g__2515(w__1986 ,w__1807 ,w__1940);
  nor g__2516(w__1985 ,w__1866 ,w__1946);
  or g__2517(w__1984 ,w__1867 ,w__1954);
  xnor g__2518(w__1983 ,w__1890 ,w__1933);
  xnor g__2519(w__1982 ,w__1869 ,w__1651);
  and g__2520(w__1999 ,w__1873 ,w__1949);
  and g__2521(w__1997 ,w__1924 ,w__1950);
  not g__2522(w__1975 ,w__1974);
  not g__2523(w__1972 ,w__1973);
  not g__2524(w__1970 ,w__1971);
  not g__2525(w__1968 ,w__1969);
  not g__2526(w__1963 ,w__1964);
  not g__2527(w__1960 ,w__1961);
  xor g__2528(w__4483 ,w__1653 ,w__1913);
  xnor g__2529(w__1959 ,w__1786 ,w__1654);
  xnor g__2530(w__1981 ,w__1831 ,w__1914);
  xnor g__2531(w__1980 ,w__1837 ,w__1896);
  xnor g__2532(w__1979 ,w__1839 ,w__1910);
  xnor g__2533(w__1978 ,w__1820 ,w__1905);
  xnor g__2534(w__1977 ,w__1813 ,w__1903);
  xnor g__2535(w__1976 ,w__1810 ,w__1902);
  xnor g__2536(w__1974 ,w__1893 ,w__1899);
  xnor g__2537(w__1973 ,w__1788 ,w__1912);
  xnor g__2538(w__1971 ,w__1793 ,w__1898);
  xnor g__2539(w__1969 ,w__1652 ,w__1897);
  xnor g__2540(w__1967 ,w__1783 ,w__1908);
  xnor g__2541(w__1966 ,w__1773 ,w__1909);
  xnor g__2542(w__1965 ,w__1808 ,w__1911);
  xnor g__2543(w__1964 ,w__1838 ,w__1904);
  xnor g__2544(w__1962 ,w__1812 ,w__1900);
  xnor g__2545(w__1961 ,w__1895 ,w__1901);
  not g__2546(w__1953 ,w__1954);
  or g__2547(w__1950 ,w__1931 ,w__1654);
  or g__2548(w__1949 ,w__1880 ,w__1652);
  nor g__2549(w__1948 ,w__1890 ,w__1932);
  and g__2550(w__1947 ,w__1870 ,w__1651);
  and g__2551(w__1958 ,w__1878 ,w__1930);
  and g__2552(w__1957 ,w__1885 ,w__1922);
  and g__2553(w__1956 ,w__1879 ,w__1920);
  and g__2554(w__1955 ,w__1865 ,w__1928);
  and g__2555(w__1954 ,w__1860 ,w__1923);
  and g__2556(w__1952 ,w__1862 ,w__1926);
  and g__2557(w__1951 ,w__1883 ,w__1915);
  not g__2558(w__1943 ,w__1944);
  not g__2559(w__1941 ,w__1942);
  nor g__2560(w__1936 ,w__1870 ,w__1651);
  or g__2561(w__1935 ,w__1889 ,w__1933);
  nor g__2562(w__1934 ,w__1876 ,w__1653);
  and g__2563(w__1946 ,w__1853 ,w__1927);
  and g__2564(w__1945 ,w__1848 ,w__1921);
  or g__2565(w__1944 ,w__1872 ,w__1919);
  and g__2566(w__1942 ,w__1858 ,w__1918);
  and g__2567(w__1940 ,w__1857 ,w__1929);
  and g__2568(w__1939 ,w__1849 ,w__1916);
  and g__2569(w__1938 ,w__1874 ,w__1925);
  and g__2570(w__1937 ,w__1881 ,w__1917);
  not g__2571(w__1932 ,w__1933);
  nor g__2572(w__1931 ,w__1785 ,w__1892);
  or g__2573(w__1930 ,w__1804 ,w__1863);
  or g__2574(w__1929 ,w__1803 ,w__1875);
  or g__2575(w__1928 ,w__1886 ,w__1894);
  or g__2576(w__1927 ,w__1796 ,w__1859);
  or g__2577(w__1926 ,w__1793 ,w__1864);
  or g__2578(w__1925 ,w__1838 ,w__1861);
  or g__2579(w__1924 ,w__1786 ,w__1891);
  or g__2580(w__1923 ,w__1839 ,w__1887);
  or g__2581(w__1922 ,w__1831 ,w__1882);
  or g__2582(w__1921 ,w__1801 ,w__1871);
  or g__2583(w__1920 ,w__1794 ,w__1855);
  and g__2584(w__1919 ,w__1877 ,w__1895);
  or g__2585(w__1918 ,w__1837 ,w__1854);
  or g__2586(w__1917 ,w__1840 ,w__1856);
  or g__2587(w__1916 ,w__1795 ,w__1847);
  xor g__2588(w__4484 ,w__1805 ,w__1845);
  or g__2589(w__1915 ,w__1834 ,w__1884);
  xnor g__2590(w__1914 ,w__1824 ,w__1827);
  xnor g__2591(w__1913 ,w__1809 ,w__1821);
  xnor g__2592(w__1933 ,w__1841 ,w__1829);
  xnor g__2593(w__1912 ,w__1782 ,w__1794);
  xnor g__2594(w__1911 ,w__1787 ,w__1803);
  xnor g__2595(w__1910 ,w__1784 ,w__1815);
  xnor g__2596(w__1909 ,w__1781 ,w__1801);
  xnor g__2597(w__1908 ,w__1776 ,w__1840);
  xnor g__2598(w__1907 ,w__1774 ,w__1779);
  xnor g__2599(w__1906 ,w__1828 ,w__1822);
  xnor g__2600(w__1905 ,w__1780 ,w__1834);
  xnor g__2601(w__1904 ,w__1778 ,w__1816);
  xnor g__2602(w__1903 ,w__1826 ,w__1804);
  xnor g__2603(w__1902 ,w__1825 ,w__1795);
  xnor g__2604(w__1901 ,w__1772 ,w__1790);
  xnor g__2605(w__1900 ,w__1777 ,w__1796);
  xnor g__2606(w__1899 ,w__1806 ,w__1814);
  xnor g__2607(w__1898 ,w__1811 ,w__1819);
  xnor g__2608(w__1897 ,w__1775 ,w__1818);
  xnor g__2609(w__1896 ,w__1823 ,w__1817);
  not g__2610(w__1894 ,w__1893);
  not g__2611(w__1891 ,w__1892);
  not g__2612(w__1889 ,w__1890);
  or g__2613(w__1888 ,w__1774 ,w__1779);
  and g__2614(w__1887 ,w__1784 ,w__1815);
  and g__2615(w__1886 ,w__1806 ,w__1814);
  or g__2616(w__1885 ,w__1824 ,w__1827);
  and g__2617(w__1884 ,w__1820 ,w__1780);
  or g__2618(w__1883 ,w__1820 ,w__1780);
  and g__2619(w__1882 ,w__1824 ,w__1827);
  or g__2620(w__1881 ,w__1783 ,w__1776);
  and g__2621(w__1880 ,w__1775 ,w__1818);
  or g__2622(w__1879 ,w__1788 ,w__1782);
  or g__2623(w__1878 ,w__1813 ,w__1826);
  or g__2624(w__1877 ,w__1771 ,w__1789);
  and g__2625(w__1876 ,w__1809 ,w__1821);
  and g__2626(w__1875 ,w__1808 ,w__1787);
  or g__2627(w__1874 ,w__1778 ,w__1816);
  or g__2628(w__1873 ,w__1775 ,w__1818);
  nor g__2629(w__1872 ,w__1772 ,w__1790);
  and g__2630(w__1871 ,w__1781 ,w__1773);
  and g__2631(w__1895 ,w__1842 ,w__1830);
  and g__2632(w__1893 ,w__1791 ,w__1802);
  and g__2633(w__1892 ,w__1836 ,w__1798);
  and g__2634(w__1890 ,w__1833 ,w__1792);
  not g__2635(w__1870 ,w__1869);
  not g__2636(w__1867 ,w__1868);
  and g__2637(w__1866 ,w__1828 ,w__1822);
  or g__2638(w__1865 ,w__1806 ,w__1814);
  and g__2639(w__1864 ,w__1811 ,w__1819);
  and g__2640(w__1863 ,w__1813 ,w__1826);
  or g__2641(w__1862 ,w__1811 ,w__1819);
  and g__2642(w__1861 ,w__1778 ,w__1816);
  or g__2643(w__1860 ,w__1784 ,w__1815);
  and g__2644(w__1859 ,w__1812 ,w__1777);
  or g__2645(w__1858 ,w__1823 ,w__1817);
  or g__2646(w__1857 ,w__1808 ,w__1787);
  and g__2647(w__1856 ,w__1783 ,w__1776);
  and g__2648(w__1855 ,w__1788 ,w__1782);
  and g__2649(w__1854 ,w__1823 ,w__1817);
  or g__2650(w__1853 ,w__1812 ,w__1777);
  nor g__2651(w__1852 ,w__1828 ,w__1822);
  nor g__2652(w__1851 ,w__1809 ,w__1821);
  and g__2653(w__1850 ,w__1774 ,w__1779);
  or g__2654(w__1849 ,w__1810 ,w__1825);
  or g__2655(w__1848 ,w__1781 ,w__1773);
  and g__2656(w__1847 ,w__1810 ,w__1825);
  nor g__2657(w__1846 ,w__1845 ,w__1805);
  and g__2658(w__1869 ,w__1844 ,w__1800);
  and g__2659(w__1868 ,w__1799 ,w__1797);
  not g__2660(w__1844 ,w__1843);
  not g__2661(w__1842 ,w__1841);
  not g__2662(w__1836 ,w__1835);
  not g__2663(w__1833 ,w__1832);
  not g__2664(w__1830 ,w__1829);
  and g__2665(w__4438 ,in8[8] ,in9[7]);
  or g__2666(w__1845 ,w__1667 ,w__1760);
  or g__2667(w__1843 ,w__1707 ,w__1687);
  or g__2668(w__1841 ,w__1662 ,w__1730);
  or g__2669(w__1840 ,w__1669 ,w__1697);
  or g__2670(w__1839 ,w__1701 ,w__1712);
  or g__2671(w__1838 ,w__1701 ,w__1691);
  or g__2672(w__1837 ,w__1707 ,w__1692);
  or g__2673(w__1835 ,w__1681 ,w__1730);
  or g__2674(w__1834 ,w__1677 ,w__1688);
  or g__2675(w__1832 ,w__1719 ,w__1687);
  or g__2676(w__1831 ,w__1679 ,w__1698);
  or g__2677(w__1829 ,w__1683 ,w__1688);
  or g__2678(w__1828 ,w__1716 ,w__1727);
  or g__2679(w__1827 ,w__1672 ,w__1659);
  or g__2680(w__1826 ,w__1675 ,w__1709);
  or g__2681(w__1825 ,w__1716 ,w__1685);
  or g__2682(w__1824 ,w__1765 ,w__1721);
  or g__2683(w__1823 ,w__1689 ,w__1656);
  or g__2684(w__1822 ,w__1665 ,w__1703);
  or g__2685(w__1821 ,w__1737 ,w__1691);
  or g__2686(w__1820 ,w__1719 ,w__1744);
  or g__2687(w__1819 ,w__1706 ,w__1713);
  or g__2688(w__1818 ,w__1671 ,w__1704);
  or g__2689(w__1817 ,w__1734 ,w__1660);
  or g__2690(w__1816 ,w__1674 ,w__1742);
  or g__2691(w__1815 ,w__1758 ,w__1722);
  or g__2692(w__1814 ,w__1733 ,w__1695);
  or g__2693(w__1813 ,w__1757 ,w__1724);
  or g__2694(w__1812 ,w__1766 ,w__1725);
  or g__2695(w__1811 ,w__1736 ,w__1657);
  or g__2696(w__1810 ,w__1718 ,w__1728);
  or g__2697(w__1809 ,w__1739 ,w__1712);
  or g__2698(w__1808 ,w__1669 ,w__1710);
  or g__2699(w__1807 ,w__1700 ,w__1703);
  or g__2700(w__1806 ,w__1739 ,w__1709);
  not g__2701(w__1790 ,w__1789);
  not g__2702(w__1786 ,w__1785);
  not g__2703(w__1772 ,w__1771);
  nor g__2704(w__1770 ,w__1734 ,w__1642);
  nor g__2705(w__1769 ,w__1737 ,w__1644);
  nor g__2706(w__1768 ,w__1760 ,w__1646);
  nor g__2707(w__1767 ,w__1740 ,w__1731);
  or g__2708(w__1805 ,w__1689 ,w__1697);
  or g__2709(w__1804 ,w__1662 ,w__1721);
  or g__2710(w__1803 ,w__1664 ,w__1744);
  and g__2711(w__1802 ,in8[5] ,in9[0]);
  or g__2712(w__1801 ,w__1763 ,w__1713);
  and g__2713(w__1800 ,in8[3] ,in9[0]);
  and g__2714(w__1799 ,in8[7] ,in9[2]);
  and g__2715(w__1798 ,in8[4] ,in9[0]);
  and g__2716(w__1797 ,in8[8] ,in9[1]);
  or g__2717(w__1796 ,w__1762 ,w__1695);
  or g__2718(w__1795 ,w__1665 ,w__1742);
  or g__2719(w__1794 ,w__1677 ,w__1692);
  or g__2720(w__1793 ,w__1672 ,w__1698);
  and g__2721(w__1792 ,in8[6] ,in9[0]);
  and g__2722(w__1791 ,in8[4] ,in9[1]);
  and g__2723(w__1789 ,in8[3] ,in9[5]);
  or g__2724(w__1788 ,w__1718 ,w__1752);
  or g__2725(w__1787 ,w__1755 ,w__1722);
  and g__2726(w__1785 ,in8[0] ,in9[5]);
  or g__2727(w__1784 ,w__1675 ,w__1694);
  or g__2728(w__1783 ,w__1733 ,w__1704);
  or g__2729(w__1782 ,w__1715 ,w__1660);
  or g__2730(w__1781 ,w__1740 ,w__1724);
  or g__2731(w__1780 ,w__1683 ,w__1731);
  or g__2732(w__1779 ,w__1700 ,w__1685);
  or g__2733(w__1778 ,w__1736 ,w__1727);
  or g__2734(w__1777 ,w__1715 ,w__1710);
  or g__2735(w__1776 ,w__1667 ,w__1694);
  or g__2736(w__1775 ,w__1706 ,w__1725);
  or g__2737(w__1774 ,w__1679 ,w__1728);
  or g__2738(w__1773 ,w__1681 ,w__1657);
  and g__2739(w__1771 ,in8[2] ,in9[6]);
  not g__2740(w__1766 ,in8[6]);
  not g__2741(w__1765 ,in8[2]);
  not g__2742(w__1764 ,in8[1]);
  not g__2743(w__1763 ,in8[4]);
  not g__2744(w__1762 ,in8[8]);
  not g__2745(w__1761 ,in9[3]);
  not g__2746(w__1760 ,in9[0]);
  not g__2747(w__1759 ,in9[1]);
  not g__2748(w__1758 ,in8[5]);
  not g__2749(w__1757 ,in8[3]);
  not g__2750(w__1756 ,in8[0]);
  not g__2751(w__1755 ,in8[7]);
  not g__2752(w__1754 ,in9[4]);
  not g__2753(w__1753 ,in9[2]);
  not g__2754(w__1752 ,in9[5]);
  not g__2755(w__1751 ,in9[7]);
  not g__2756(w__1750 ,in9[6]);
  not g__2757(w__1649 ,w__1748);
  not g__2758(w__1748 ,w__1756);
  not g__2759(w__1648 ,w__1747);
  not g__2760(w__1641 ,w__1747);
  not g__2761(w__1747 ,w__1759);
  not g__2762(w__1647 ,w__1746);
  not g__2763(w__1746 ,w__1760);
  buf g__2764(w__4451 ,w__1770);
  buf g__2765(w__4485 ,w__1767);
  buf g__2766(w__4453 ,w__1768);
  buf g__2767(w__4452 ,w__1769);
  buf g__2768(w__4450 ,w__1846);
  not g__2769(w__1745 ,w__1749);
  not g__2770(w__1749 ,w__2050);
  not g__2771(w__1744 ,w__1743);
  not g__2772(w__1743 ,w__1761);
  not g__2773(w__1742 ,w__1741);
  not g__2774(w__1741 ,w__1754);
  not g__2775(w__1740 ,w__1738);
  not g__2776(w__1739 ,w__1738);
  not g__2777(w__1738 ,w__1756);
  not g__2778(w__1737 ,w__1735);
  not g__2779(w__1736 ,w__1735);
  not g__2780(w__1735 ,w__1764);
  not g__2781(w__1734 ,w__1732);
  not g__2782(w__1733 ,w__1732);
  not g__2783(w__1732 ,w__1764);
  not g__2784(w__1731 ,w__1729);
  not g__2785(w__1730 ,w__1729);
  not g__2786(w__1729 ,w__1648);
  not g__2787(w__1728 ,w__1726);
  not g__2788(w__1727 ,w__1726);
  not g__2789(w__1726 ,w__1751);
  not g__2790(w__1725 ,w__1723);
  not g__2791(w__1724 ,w__1723);
  not g__2792(w__1723 ,w__1751);
  not g__2793(w__1722 ,w__1720);
  not g__2794(w__1721 ,w__1720);
  not g__2795(w__1720 ,w__1754);
  not g__2796(w__1719 ,w__1717);
  not g__2797(w__1718 ,w__1717);
  not g__2798(w__1717 ,w__1758);
  not g__2799(w__1716 ,w__1714);
  not g__2800(w__1715 ,w__1714);
  not g__2801(w__1714 ,w__1755);
  not g__2802(w__1713 ,w__1711);
  not g__2803(w__1712 ,w__1711);
  not g__2804(w__1711 ,w__1761);
  not g__2805(w__1710 ,w__1708);
  not g__2806(w__1709 ,w__1708);
  not g__2807(w__1708 ,w__1750);
  not g__2808(w__1707 ,w__1705);
  not g__2809(w__1706 ,w__1705);
  not g__2810(w__1705 ,w__1765);
  not g__2811(w__1704 ,w__1702);
  not g__2812(w__1703 ,w__1702);
  not g__2813(w__1702 ,w__1750);
  not g__2814(w__1701 ,w__1699);
  not g__2815(w__1700 ,w__1699);
  not g__2816(w__1699 ,w__1766);
  not g__2817(w__1698 ,w__1696);
  not g__2818(w__1697 ,w__1696);
  not g__2819(w__1696 ,w__1753);
  not g__2820(w__1695 ,w__1693);
  not g__2821(w__1694 ,w__1693);
  not g__2822(w__1693 ,w__1752);
  not g__2823(w__1692 ,w__1690);
  not g__2824(w__1691 ,w__1690);
  not g__2825(w__1690 ,w__1753);
  not g__2826(w__1646 ,w__1645);
  not g__2827(w__1689 ,w__1645);
  not g__2828(w__1645 ,w__1649);
  not g__2829(w__1644 ,w__1643);
  not g__2830(w__1688 ,w__1643);
  not g__2831(w__1643 ,w__1647);
  not g__2832(w__1642 ,w__1686);
  not g__2833(w__1687 ,w__1686);
  not g__2834(w__1686 ,w__1641);
  not g__2835(w__1685 ,w__1684);
  not g__2836(w__1684 ,w__1752);
  not g__2837(w__1683 ,w__1682);
  not g__2838(w__1682 ,w__1755);
  not g__2839(w__1681 ,w__1680);
  not g__2840(w__1680 ,w__1757);
  not g__2841(w__1679 ,w__1678);
  not g__2842(w__1678 ,w__1763);
  not g__2843(w__1677 ,w__1676);
  not g__2844(w__1676 ,w__1762);
  not g__2845(w__1675 ,w__1673);
  not g__2846(w__1674 ,w__1673);
  not g__2847(w__1673 ,w__1763);
  not g__2848(w__1672 ,w__1670);
  not g__2849(w__1671 ,w__1670);
  not g__2850(w__1670 ,w__1757);
  not g__2851(w__1669 ,w__1668);
  not g__2852(w__1668 ,w__1758);
  not g__2853(w__1667 ,w__1666);
  not g__2854(w__1666 ,w__1765);
  not g__2855(w__1665 ,w__1663);
  not g__2856(w__1664 ,w__1663);
  not g__2857(w__1663 ,w__1762);
  not g__2858(w__1662 ,w__1661);
  not g__2859(w__1661 ,w__1766);
  not g__2860(w__1660 ,w__1658);
  not g__2861(w__1659 ,w__1658);
  not g__2862(w__1658 ,w__1761);
  not g__2863(w__1657 ,w__1655);
  not g__2864(w__1656 ,w__1655);
  not g__2865(w__1655 ,w__1754);
  xnor g__2866(w__1654 ,w__1791 ,w__1802);
  xor g__2867(w__1653 ,w__1843 ,w__1800);
  xnor g__2868(w__1652 ,w__1799 ,w__1797);
  xor g__2869(w__1651 ,w__1835 ,w__1798);
  xor g__2870(w__1650 ,w__1832 ,w__1792);
  xnor g__2871(w__4347 ,w__2538 ,w__2555);
  or g__2872(w__4313 ,w__2554 ,w__2556);
  xnor g__2873(w__4346 ,w__2550 ,w__2551);
  nor g__2874(w__2556 ,w__2538 ,w__2553);
  or g__2875(w__4345 ,w__2546 ,w__2552);
  xnor g__2876(w__2555 ,w__2502 ,w__2544);
  xnor g__2877(w__4348 ,w__2529 ,w__2541);
  xnor g__2878(w__4349 ,w__2531 ,w__2540);
  xor g__2879(w__4312 ,w__2537 ,w__2539);
  or g__2880(w__4315 ,w__2535 ,w__2548);
  nor g__2881(w__2554 ,w__2502 ,w__2545);
  or g__2882(w__4344 ,w__2536 ,w__2547);
  and g__2883(w__2553 ,w__2502 ,w__2545);
  and g__2884(w__2552 ,w__2550 ,w__2542);
  or g__2885(w__4314 ,w__2524 ,w__2549);
  or g__2886(w__4316 ,w__2518 ,w__2543);
  xnor g__2887(w__4350 ,w__2530 ,w__2523);
  xnor g__2888(w__2551 ,w__2528 ,w__2504);
  and g__2889(w__2549 ,w__2534 ,w__2529);
  and g__2890(w__2548 ,w__2533 ,w__2531);
  or g__2891(w__4317 ,w__2483 ,w__2532);
  nor g__2892(w__2547 ,w__2526 ,w__2537);
  nor g__2893(w__2546 ,w__2504 ,w__2528);
  or g__2894(w__2550 ,w__2464 ,w__2525);
  not g__2895(w__2545 ,w__2544);
  nor g__2896(w__2543 ,w__2519 ,w__2530);
  or g__2897(w__2542 ,w__2503 ,w__2527);
  xnor g__2898(w__4351 ,w__2515 ,w__2490);
  xnor g__2899(w__2541 ,w__2511 ,w__2508);
  xnor g__2900(w__2540 ,w__2513 ,w__2522);
  xnor g__2901(w__2539 ,w__2509 ,w__2484);
  xnor g__2902(w__2544 ,w__2514 ,w__2488);
  nor g__2903(w__2536 ,w__2484 ,w__2509);
  nor g__2904(w__2535 ,w__2522 ,w__2513);
  or g__2905(w__2534 ,w__2207 ,w__2510);
  or g__2906(w__2533 ,w__2521 ,w__2512);
  or g__2907(w__4343 ,w__2468 ,w__2507);
  nor g__2908(w__2532 ,w__2474 ,w__2515);
  or g__2909(w__4318 ,w__2473 ,w__2516);
  and g__2910(w__2538 ,w__2475 ,w__2517);
  and g__2911(w__2537 ,w__2500 ,w__2520);
  not g__2912(w__2527 ,w__2528);
  and g__2913(w__2526 ,w__2484 ,w__2509);
  and g__2914(w__2525 ,w__2463 ,w__2514);
  nor g__2915(w__2524 ,w__2203 ,w__2511);
  xor g__2916(w__4311 ,w__2505 ,w__2486);
  xnor g__2917(w__4352 ,w__2496 ,w__2492);
  xnor g__2918(w__2523 ,w__2501 ,w__2494);
  xnor g__2919(w__2531 ,w__2485 ,w__2493);
  xnor g__2920(w__2530 ,w__2413 ,w__2487);
  xnor g__2921(w__2529 ,w__2506 ,w__2489);
  xnor g__2922(w__2528 ,w__2470 ,w__2491);
  not g__2923(w__2522 ,w__2521);
  or g__2924(w__2520 ,w__2414 ,w__2497);
  and g__2925(w__2519 ,w__2501 ,w__2495);
  nor g__2926(w__2518 ,w__2501 ,w__2495);
  or g__2927(w__2517 ,w__2471 ,w__2506);
  and g__2928(w__2516 ,w__2472 ,w__2496);
  or g__2929(w__2521 ,w__2479 ,w__2498);
  not g__2930(w__2512 ,w__2513);
  not g__2931(w__2510 ,w__2511);
  nor g__2932(w__2507 ,w__2467 ,w__2505);
  xnor g__2933(w__2515 ,w__2439 ,w__2461);
  xnor g__2934(w__2514 ,w__2435 ,w__2460);
  xnor g__2935(w__2513 ,w__2436 ,w__2462);
  and g__2936(w__2511 ,w__2469 ,w__2499);
  xnor g__2937(w__2509 ,w__2434 ,w__2459);
  xnor g__2938(w__2508 ,w__2437 ,w__2458);
  not g__2939(w__2503 ,w__2504);
  or g__2940(w__2500 ,w__2423 ,w__2470);
  or g__2941(w__2499 ,w__2485 ,w__2481);
  nor g__2942(w__2498 ,w__2413 ,w__2478);
  and g__2943(w__2497 ,w__2423 ,w__2470);
  or g__2944(w__4319 ,w__2394 ,w__2476);
  and g__2945(w__2506 ,w__2446 ,w__2466);
  and g__2946(w__2505 ,w__2444 ,w__2482);
  and g__2947(w__2504 ,w__2442 ,w__2465);
  and g__2948(w__2502 ,w__2453 ,w__2480);
  and g__2949(w__2501 ,w__2450 ,w__2477);
  not g__2950(w__2495 ,w__2494);
  xnor g__2951(w__4353 ,w__2438 ,w__2440);
  xnor g__2952(w__2493 ,w__2422 ,w__2419);
  xnor g__2953(w__2492 ,w__2429 ,w__2400);
  xnor g__2954(w__2491 ,w__2423 ,w__2414);
  xnor g__2955(w__2490 ,w__2455 ,w__2432);
  xnor g__2956(w__2489 ,w__2402 ,w__2427);
  xnor g__2957(w__2488 ,w__2431 ,w__2457);
  xnor g__2958(w__2487 ,w__2425 ,w__2424);
  xnor g__2959(w__2486 ,w__2420 ,w__2397);
  xnor g__2960(w__2496 ,w__2350 ,w__2417);
  xnor g__2961(w__2494 ,w__2415 ,w__2441);
  nor g__2962(w__2483 ,w__2455 ,w__2433);
  or g__2963(w__2482 ,w__2448 ,w__2434);
  nor g__2964(w__2481 ,w__2421 ,w__2419);
  or g__2965(w__2480 ,w__2437 ,w__2452);
  nor g__2966(w__2479 ,w__2424 ,w__2425);
  and g__2967(w__2478 ,w__2424 ,w__2425);
  or g__2968(w__2477 ,w__2449 ,w__2439);
  nor g__2969(w__2476 ,w__2405 ,w__2438);
  or g__2970(w__2475 ,w__2401 ,w__2427);
  and g__2971(w__2474 ,w__2455 ,w__2433);
  nor g__2972(w__2473 ,w__2400 ,w__2429);
  or g__2973(w__2472 ,w__2399 ,w__2428);
  nor g__2974(w__2471 ,w__2402 ,w__2426);
  and g__2975(w__2485 ,w__2393 ,w__2445);
  and g__2976(w__2484 ,w__2346 ,w__2454);
  or g__2977(w__2469 ,w__2422 ,w__2418);
  nor g__2978(w__2468 ,w__2397 ,w__2420);
  and g__2979(w__2467 ,w__2397 ,w__2420);
  or g__2980(w__2466 ,w__2436 ,w__2451);
  or g__2981(w__2465 ,w__2447 ,w__2435);
  nor g__2982(w__2464 ,w__2457 ,w__2431);
  or g__2983(w__2463 ,w__2456 ,w__2430);
  or g__2984(w__4342 ,w__2310 ,w__2443);
  xor g__2985(w__4310 ,w__2404 ,w__2364);
  xnor g__2986(w__2462 ,w__2403 ,w__2395);
  xnor g__2987(w__2461 ,w__2410 ,w__2108);
  xnor g__2988(w__2460 ,w__2326 ,w__2412);
  xnor g__2989(w__2459 ,w__2265 ,w__2398);
  xnor g__2990(w__2458 ,w__2409 ,w__2396);
  xnor g__2991(w__2470 ,w__2416 ,w__2365);
  not g__2992(w__2456 ,w__2457);
  or g__2993(w__2454 ,w__2308 ,w__2416);
  or g__2994(w__2453 ,w__2396 ,w__2409);
  and g__2995(w__2452 ,w__2396 ,w__2409);
  and g__2996(w__2451 ,w__2395 ,w__2403);
  or g__2997(w__2450 ,w__2108 ,w__2410);
  and g__2998(w__2449 ,w__2108 ,w__2410);
  and g__2999(w__2448 ,w__2265 ,w__2398);
  nor g__3000(w__2447 ,w__2326 ,w__2411);
  or g__3001(w__2446 ,w__2395 ,w__2403);
  or g__3002(w__2445 ,w__2415 ,w__2406);
  or g__3003(w__4320 ,w__2309 ,w__2392);
  or g__3004(w__2444 ,w__2265 ,w__2398);
  nor g__3005(w__2443 ,w__2324 ,w__2404);
  or g__3006(w__2442 ,w__2325 ,w__2412);
  xnor g__3007(w__2441 ,w__2348 ,w__2391);
  xnor g__3008(w__2440 ,w__2327 ,w__2109);
  and g__3009(w__2457 ,w__2331 ,w__2407);
  and g__3010(w__2455 ,w__2382 ,w__2408);
  not g__3011(w__2433 ,w__2432);
  not g__3012(w__2430 ,w__2431);
  not g__3013(w__2428 ,w__2429);
  not g__3014(w__2426 ,w__2427);
  not g__3015(w__2421 ,w__2422);
  not g__3016(w__2418 ,w__2419);
  xor g__3017(w__4354 ,w__2111 ,w__2371);
  xnor g__3018(w__2417 ,w__2244 ,w__2112);
  xnor g__3019(w__2439 ,w__2289 ,w__2372);
  xnor g__3020(w__2438 ,w__2295 ,w__2354);
  xnor g__3021(w__2437 ,w__2297 ,w__2368);
  xnor g__3022(w__2436 ,w__2278 ,w__2363);
  xnor g__3023(w__2435 ,w__2271 ,w__2361);
  xnor g__3024(w__2434 ,w__2268 ,w__2360);
  xnor g__3025(w__2432 ,w__2351 ,w__2357);
  xnor g__3026(w__2431 ,w__2246 ,w__2370);
  xnor g__3027(w__2429 ,w__2251 ,w__2356);
  xnor g__3028(w__2427 ,w__2110 ,w__2355);
  xnor g__3029(w__2425 ,w__2241 ,w__2366);
  xnor g__3030(w__2424 ,w__2231 ,w__2367);
  xnor g__3031(w__2423 ,w__2266 ,w__2369);
  xnor g__3032(w__2422 ,w__2296 ,w__2362);
  xnor g__3033(w__2420 ,w__2270 ,w__2358);
  xnor g__3034(w__2419 ,w__2353 ,w__2359);
  not g__3035(w__2411 ,w__2412);
  or g__3036(w__2408 ,w__2389 ,w__2112);
  or g__3037(w__2407 ,w__2338 ,w__2110);
  nor g__3038(w__2406 ,w__2348 ,w__2390);
  and g__3039(w__2405 ,w__2328 ,w__2109);
  and g__3040(w__2416 ,w__2336 ,w__2388);
  and g__3041(w__2415 ,w__2343 ,w__2380);
  and g__3042(w__2414 ,w__2337 ,w__2378);
  and g__3043(w__2413 ,w__2323 ,w__2386);
  and g__3044(w__2412 ,w__2318 ,w__2381);
  and g__3045(w__2410 ,w__2320 ,w__2384);
  and g__3046(w__2409 ,w__2341 ,w__2373);
  not g__3047(w__2401 ,w__2402);
  not g__3048(w__2399 ,w__2400);
  nor g__3049(w__2394 ,w__2328 ,w__2109);
  or g__3050(w__2393 ,w__2347 ,w__2391);
  nor g__3051(w__2392 ,w__2334 ,w__2111);
  and g__3052(w__2404 ,w__2311 ,w__2385);
  and g__3053(w__2403 ,w__2306 ,w__2379);
  or g__3054(w__2402 ,w__2330 ,w__2377);
  and g__3055(w__2400 ,w__2316 ,w__2376);
  and g__3056(w__2398 ,w__2315 ,w__2387);
  and g__3057(w__2397 ,w__2307 ,w__2374);
  and g__3058(w__2396 ,w__2332 ,w__2383);
  and g__3059(w__2395 ,w__2339 ,w__2375);
  not g__3060(w__2390 ,w__2391);
  nor g__3061(w__2389 ,w__2243 ,w__2350);
  or g__3062(w__2388 ,w__2262 ,w__2321);
  or g__3063(w__2387 ,w__2261 ,w__2333);
  or g__3064(w__2386 ,w__2344 ,w__2352);
  or g__3065(w__2385 ,w__2254 ,w__2317);
  or g__3066(w__2384 ,w__2251 ,w__2322);
  or g__3067(w__2383 ,w__2296 ,w__2319);
  or g__3068(w__2382 ,w__2244 ,w__2349);
  or g__3069(w__2381 ,w__2297 ,w__2345);
  or g__3070(w__2380 ,w__2289 ,w__2340);
  or g__3071(w__2379 ,w__2259 ,w__2329);
  or g__3072(w__2378 ,w__2252 ,w__2313);
  and g__3073(w__2377 ,w__2335 ,w__2353);
  or g__3074(w__2376 ,w__2295 ,w__2312);
  or g__3075(w__2375 ,w__2298 ,w__2314);
  or g__3076(w__2374 ,w__2253 ,w__2305);
  xor g__3077(w__4355 ,w__2263 ,w__2303);
  or g__3078(w__2373 ,w__2292 ,w__2342);
  xnor g__3079(w__2372 ,w__2282 ,w__2285);
  xnor g__3080(w__2371 ,w__2267 ,w__2279);
  xnor g__3081(w__2391 ,w__2299 ,w__2287);
  xnor g__3082(w__2370 ,w__2240 ,w__2252);
  xnor g__3083(w__2369 ,w__2245 ,w__2261);
  xnor g__3084(w__2368 ,w__2242 ,w__2273);
  xnor g__3085(w__2367 ,w__2239 ,w__2259);
  xnor g__3086(w__2366 ,w__2234 ,w__2298);
  xnor g__3087(w__2365 ,w__2232 ,w__2237);
  xnor g__3088(w__2364 ,w__2286 ,w__2280);
  xnor g__3089(w__2363 ,w__2238 ,w__2292);
  xnor g__3090(w__2362 ,w__2236 ,w__2274);
  xnor g__3091(w__2361 ,w__2284 ,w__2262);
  xnor g__3092(w__2360 ,w__2283 ,w__2253);
  xnor g__3093(w__2359 ,w__2230 ,w__2248);
  xnor g__3094(w__2358 ,w__2235 ,w__2254);
  xnor g__3095(w__2357 ,w__2264 ,w__2272);
  xnor g__3096(w__2356 ,w__2269 ,w__2277);
  xnor g__3097(w__2355 ,w__2233 ,w__2276);
  xnor g__3098(w__2354 ,w__2281 ,w__2275);
  not g__3099(w__2352 ,w__2351);
  not g__3100(w__2349 ,w__2350);
  not g__3101(w__2347 ,w__2348);
  or g__3102(w__2346 ,w__2232 ,w__2237);
  and g__3103(w__2345 ,w__2242 ,w__2273);
  and g__3104(w__2344 ,w__2264 ,w__2272);
  or g__3105(w__2343 ,w__2282 ,w__2285);
  and g__3106(w__2342 ,w__2278 ,w__2238);
  or g__3107(w__2341 ,w__2278 ,w__2238);
  and g__3108(w__2340 ,w__2282 ,w__2285);
  or g__3109(w__2339 ,w__2241 ,w__2234);
  and g__3110(w__2338 ,w__2233 ,w__2276);
  or g__3111(w__2337 ,w__2246 ,w__2240);
  or g__3112(w__2336 ,w__2271 ,w__2284);
  or g__3113(w__2335 ,w__2229 ,w__2247);
  and g__3114(w__2334 ,w__2267 ,w__2279);
  and g__3115(w__2333 ,w__2266 ,w__2245);
  or g__3116(w__2332 ,w__2236 ,w__2274);
  or g__3117(w__2331 ,w__2233 ,w__2276);
  nor g__3118(w__2330 ,w__2230 ,w__2248);
  and g__3119(w__2329 ,w__2239 ,w__2231);
  and g__3120(w__2353 ,w__2300 ,w__2288);
  and g__3121(w__2351 ,w__2249 ,w__2260);
  and g__3122(w__2350 ,w__2294 ,w__2256);
  and g__3123(w__2348 ,w__2291 ,w__2250);
  not g__3124(w__2328 ,w__2327);
  not g__3125(w__2325 ,w__2326);
  and g__3126(w__2324 ,w__2286 ,w__2280);
  or g__3127(w__2323 ,w__2264 ,w__2272);
  and g__3128(w__2322 ,w__2269 ,w__2277);
  and g__3129(w__2321 ,w__2271 ,w__2284);
  or g__3130(w__2320 ,w__2269 ,w__2277);
  and g__3131(w__2319 ,w__2236 ,w__2274);
  or g__3132(w__2318 ,w__2242 ,w__2273);
  and g__3133(w__2317 ,w__2270 ,w__2235);
  or g__3134(w__2316 ,w__2281 ,w__2275);
  or g__3135(w__2315 ,w__2266 ,w__2245);
  and g__3136(w__2314 ,w__2241 ,w__2234);
  and g__3137(w__2313 ,w__2246 ,w__2240);
  and g__3138(w__2312 ,w__2281 ,w__2275);
  or g__3139(w__2311 ,w__2270 ,w__2235);
  nor g__3140(w__2310 ,w__2286 ,w__2280);
  nor g__3141(w__2309 ,w__2267 ,w__2279);
  and g__3142(w__2308 ,w__2232 ,w__2237);
  or g__3143(w__2307 ,w__2268 ,w__2283);
  or g__3144(w__2306 ,w__2239 ,w__2231);
  and g__3145(w__2305 ,w__2268 ,w__2283);
  nor g__3146(w__2304 ,w__2303 ,w__2263);
  and g__3147(w__2327 ,w__2302 ,w__2258);
  and g__3148(w__2326 ,w__2257 ,w__2255);
  not g__3149(w__2302 ,w__2301);
  not g__3150(w__2300 ,w__2299);
  not g__3151(w__2294 ,w__2293);
  not g__3152(w__2291 ,w__2290);
  not g__3153(w__2288 ,w__2287);
  and g__3154(w__4309 ,in12[8] ,in13[7]);
  or g__3155(w__2303 ,w__2125 ,w__2218);
  or g__3156(w__2301 ,w__2165 ,w__2145);
  or g__3157(w__2299 ,w__2120 ,w__2188);
  or g__3158(w__2298 ,w__2127 ,w__2155);
  or g__3159(w__2297 ,w__2159 ,w__2170);
  or g__3160(w__2296 ,w__2159 ,w__2149);
  or g__3161(w__2295 ,w__2165 ,w__2150);
  or g__3162(w__2293 ,w__2139 ,w__2188);
  or g__3163(w__2292 ,w__2135 ,w__2146);
  or g__3164(w__2290 ,w__2177 ,w__2145);
  or g__3165(w__2289 ,w__2137 ,w__2156);
  or g__3166(w__2287 ,w__2141 ,w__2146);
  or g__3167(w__2286 ,w__2174 ,w__2185);
  or g__3168(w__2285 ,w__2130 ,w__2117);
  or g__3169(w__2284 ,w__2133 ,w__2167);
  or g__3170(w__2283 ,w__2174 ,w__2143);
  or g__3171(w__2282 ,w__2223 ,w__2179);
  or g__3172(w__2281 ,w__2147 ,w__2114);
  or g__3173(w__2280 ,w__2123 ,w__2161);
  or g__3174(w__2279 ,w__2195 ,w__2149);
  or g__3175(w__2278 ,w__2177 ,w__2202);
  or g__3176(w__2277 ,w__2164 ,w__2171);
  or g__3177(w__2276 ,w__2129 ,w__2162);
  or g__3178(w__2275 ,w__2192 ,w__2118);
  or g__3179(w__2274 ,w__2132 ,w__2200);
  or g__3180(w__2273 ,w__2216 ,w__2180);
  or g__3181(w__2272 ,w__2191 ,w__2153);
  or g__3182(w__2271 ,w__2215 ,w__2182);
  or g__3183(w__2270 ,w__2224 ,w__2183);
  or g__3184(w__2269 ,w__2194 ,w__2115);
  or g__3185(w__2268 ,w__2176 ,w__2186);
  or g__3186(w__2267 ,w__2197 ,w__2170);
  or g__3187(w__2266 ,w__2127 ,w__2168);
  or g__3188(w__2265 ,w__2158 ,w__2161);
  or g__3189(w__2264 ,w__2197 ,w__2167);
  not g__3190(w__2248 ,w__2247);
  not g__3191(w__2244 ,w__2243);
  not g__3192(w__2230 ,w__2229);
  nor g__3193(w__2228 ,w__2192 ,w__2100);
  nor g__3194(w__2227 ,w__2195 ,w__2102);
  nor g__3195(w__2226 ,w__2218 ,w__2104);
  nor g__3196(w__2225 ,w__2198 ,w__2189);
  or g__3197(w__2263 ,w__2147 ,w__2155);
  or g__3198(w__2262 ,w__2120 ,w__2179);
  or g__3199(w__2261 ,w__2122 ,w__2202);
  and g__3200(w__2260 ,in12[5] ,in13[0]);
  or g__3201(w__2259 ,w__2221 ,w__2171);
  and g__3202(w__2258 ,in12[3] ,in13[0]);
  and g__3203(w__2257 ,in12[7] ,in13[2]);
  and g__3204(w__2256 ,in12[4] ,in13[0]);
  and g__3205(w__2255 ,in12[8] ,in13[1]);
  or g__3206(w__2254 ,w__2220 ,w__2153);
  or g__3207(w__2253 ,w__2123 ,w__2200);
  or g__3208(w__2252 ,w__2135 ,w__2150);
  or g__3209(w__2251 ,w__2130 ,w__2156);
  and g__3210(w__2250 ,in12[6] ,in13[0]);
  and g__3211(w__2249 ,in12[4] ,in13[1]);
  and g__3212(w__2247 ,in12[3] ,in13[5]);
  or g__3213(w__2246 ,w__2176 ,w__2210);
  or g__3214(w__2245 ,w__2213 ,w__2180);
  and g__3215(w__2243 ,in12[0] ,in13[5]);
  or g__3216(w__2242 ,w__2133 ,w__2152);
  or g__3217(w__2241 ,w__2191 ,w__2162);
  or g__3218(w__2240 ,w__2173 ,w__2118);
  or g__3219(w__2239 ,w__2198 ,w__2182);
  or g__3220(w__2238 ,w__2141 ,w__2189);
  or g__3221(w__2237 ,w__2158 ,w__2143);
  or g__3222(w__2236 ,w__2194 ,w__2185);
  or g__3223(w__2235 ,w__2173 ,w__2168);
  or g__3224(w__2234 ,w__2125 ,w__2152);
  or g__3225(w__2233 ,w__2164 ,w__2183);
  or g__3226(w__2232 ,w__2137 ,w__2186);
  or g__3227(w__2231 ,w__2139 ,w__2115);
  and g__3228(w__2229 ,in12[2] ,in13[6]);
  not g__3229(w__2224 ,in12[6]);
  not g__3230(w__2223 ,in12[2]);
  not g__3231(w__2222 ,in12[1]);
  not g__3232(w__2221 ,in12[4]);
  not g__3233(w__2220 ,in12[8]);
  not g__3234(w__2219 ,in13[3]);
  not g__3235(w__2218 ,in13[0]);
  not g__3236(w__2217 ,in13[1]);
  not g__3237(w__2216 ,in12[5]);
  not g__3238(w__2215 ,in12[3]);
  not g__3239(w__2214 ,in12[0]);
  not g__3240(w__2213 ,in12[7]);
  not g__3241(w__2212 ,in13[4]);
  not g__3242(w__2211 ,in13[2]);
  not g__3243(w__2210 ,in13[5]);
  not g__3244(w__2209 ,in13[7]);
  not g__3245(w__2208 ,in13[6]);
  not g__3246(w__2107 ,w__2206);
  not g__3247(w__2206 ,w__2214);
  not g__3248(w__2106 ,w__2205);
  not g__3249(w__2099 ,w__2205);
  not g__3250(w__2205 ,w__2217);
  not g__3251(w__2105 ,w__2204);
  not g__3252(w__2204 ,w__2218);
  buf g__3253(w__4322 ,w__2228);
  buf g__3254(w__4356 ,w__2225);
  buf g__3255(w__4324 ,w__2226);
  buf g__3256(w__4323 ,w__2227);
  buf g__3257(w__4321 ,w__2304);
  not g__3258(w__2203 ,w__2207);
  not g__3259(w__2207 ,w__2508);
  not g__3260(w__2202 ,w__2201);
  not g__3261(w__2201 ,w__2219);
  not g__3262(w__2200 ,w__2199);
  not g__3263(w__2199 ,w__2212);
  not g__3264(w__2198 ,w__2196);
  not g__3265(w__2197 ,w__2196);
  not g__3266(w__2196 ,w__2214);
  not g__3267(w__2195 ,w__2193);
  not g__3268(w__2194 ,w__2193);
  not g__3269(w__2193 ,w__2222);
  not g__3270(w__2192 ,w__2190);
  not g__3271(w__2191 ,w__2190);
  not g__3272(w__2190 ,w__2222);
  not g__3273(w__2189 ,w__2187);
  not g__3274(w__2188 ,w__2187);
  not g__3275(w__2187 ,w__2106);
  not g__3276(w__2186 ,w__2184);
  not g__3277(w__2185 ,w__2184);
  not g__3278(w__2184 ,w__2209);
  not g__3279(w__2183 ,w__2181);
  not g__3280(w__2182 ,w__2181);
  not g__3281(w__2181 ,w__2209);
  not g__3282(w__2180 ,w__2178);
  not g__3283(w__2179 ,w__2178);
  not g__3284(w__2178 ,w__2212);
  not g__3285(w__2177 ,w__2175);
  not g__3286(w__2176 ,w__2175);
  not g__3287(w__2175 ,w__2216);
  not g__3288(w__2174 ,w__2172);
  not g__3289(w__2173 ,w__2172);
  not g__3290(w__2172 ,w__2213);
  not g__3291(w__2171 ,w__2169);
  not g__3292(w__2170 ,w__2169);
  not g__3293(w__2169 ,w__2219);
  not g__3294(w__2168 ,w__2166);
  not g__3295(w__2167 ,w__2166);
  not g__3296(w__2166 ,w__2208);
  not g__3297(w__2165 ,w__2163);
  not g__3298(w__2164 ,w__2163);
  not g__3299(w__2163 ,w__2223);
  not g__3300(w__2162 ,w__2160);
  not g__3301(w__2161 ,w__2160);
  not g__3302(w__2160 ,w__2208);
  not g__3303(w__2159 ,w__2157);
  not g__3304(w__2158 ,w__2157);
  not g__3305(w__2157 ,w__2224);
  not g__3306(w__2156 ,w__2154);
  not g__3307(w__2155 ,w__2154);
  not g__3308(w__2154 ,w__2211);
  not g__3309(w__2153 ,w__2151);
  not g__3310(w__2152 ,w__2151);
  not g__3311(w__2151 ,w__2210);
  not g__3312(w__2150 ,w__2148);
  not g__3313(w__2149 ,w__2148);
  not g__3314(w__2148 ,w__2211);
  not g__3315(w__2104 ,w__2103);
  not g__3316(w__2147 ,w__2103);
  not g__3317(w__2103 ,w__2107);
  not g__3318(w__2102 ,w__2101);
  not g__3319(w__2146 ,w__2101);
  not g__3320(w__2101 ,w__2105);
  not g__3321(w__2100 ,w__2144);
  not g__3322(w__2145 ,w__2144);
  not g__3323(w__2144 ,w__2099);
  not g__3324(w__2143 ,w__2142);
  not g__3325(w__2142 ,w__2210);
  not g__3326(w__2141 ,w__2140);
  not g__3327(w__2140 ,w__2213);
  not g__3328(w__2139 ,w__2138);
  not g__3329(w__2138 ,w__2215);
  not g__3330(w__2137 ,w__2136);
  not g__3331(w__2136 ,w__2221);
  not g__3332(w__2135 ,w__2134);
  not g__3333(w__2134 ,w__2220);
  not g__3334(w__2133 ,w__2131);
  not g__3335(w__2132 ,w__2131);
  not g__3336(w__2131 ,w__2221);
  not g__3337(w__2130 ,w__2128);
  not g__3338(w__2129 ,w__2128);
  not g__3339(w__2128 ,w__2215);
  not g__3340(w__2127 ,w__2126);
  not g__3341(w__2126 ,w__2216);
  not g__3342(w__2125 ,w__2124);
  not g__3343(w__2124 ,w__2223);
  not g__3344(w__2123 ,w__2121);
  not g__3345(w__2122 ,w__2121);
  not g__3346(w__2121 ,w__2220);
  not g__3347(w__2120 ,w__2119);
  not g__3348(w__2119 ,w__2224);
  not g__3349(w__2118 ,w__2116);
  not g__3350(w__2117 ,w__2116);
  not g__3351(w__2116 ,w__2219);
  not g__3352(w__2115 ,w__2113);
  not g__3353(w__2114 ,w__2113);
  not g__3354(w__2113 ,w__2212);
  xnor g__3355(w__2112 ,w__2249 ,w__2260);
  xor g__3356(w__2111 ,w__2301 ,w__2258);
  xnor g__3357(w__2110 ,w__2257 ,w__2255);
  xor g__3358(w__2109 ,w__2293 ,w__2256);
  xor g__3359(w__2108 ,w__2290 ,w__2250);
  xnor g__3360(w__4281 ,w__2996 ,w__3013);
  or g__3361(w__4249 ,w__3012 ,w__3014);
  xnor g__3362(w__4280 ,w__3008 ,w__3009);
  nor g__3363(w__3014 ,w__2996 ,w__3011);
  or g__3364(w__4279 ,w__3004 ,w__3010);
  xnor g__3365(w__3013 ,w__2960 ,w__3002);
  xnor g__3366(w__4282 ,w__2987 ,w__2999);
  xnor g__3367(w__4283 ,w__2989 ,w__2998);
  xor g__3368(w__4248 ,w__2995 ,w__2997);
  or g__3369(w__4251 ,w__2993 ,w__3006);
  nor g__3370(w__3012 ,w__2960 ,w__3003);
  or g__3371(w__4278 ,w__2994 ,w__3005);
  and g__3372(w__3011 ,w__2960 ,w__3003);
  and g__3373(w__3010 ,w__3008 ,w__3000);
  or g__3374(w__4250 ,w__2982 ,w__3007);
  or g__3375(w__4252 ,w__2976 ,w__3001);
  xnor g__3376(w__4284 ,w__2988 ,w__2981);
  xnor g__3377(w__3009 ,w__2986 ,w__2962);
  and g__3378(w__3007 ,w__2992 ,w__2987);
  and g__3379(w__3006 ,w__2991 ,w__2989);
  or g__3380(w__4253 ,w__2941 ,w__2990);
  nor g__3381(w__3005 ,w__2984 ,w__2995);
  nor g__3382(w__3004 ,w__2962 ,w__2986);
  or g__3383(w__3008 ,w__2922 ,w__2983);
  not g__3384(w__3003 ,w__3002);
  nor g__3385(w__3001 ,w__2977 ,w__2988);
  or g__3386(w__3000 ,w__2961 ,w__2985);
  xnor g__3387(w__4285 ,w__2973 ,w__2948);
  xnor g__3388(w__2999 ,w__2969 ,w__2966);
  xnor g__3389(w__2998 ,w__2971 ,w__2980);
  xnor g__3390(w__2997 ,w__2967 ,w__2942);
  xnor g__3391(w__3002 ,w__2972 ,w__2946);
  nor g__3392(w__2994 ,w__2942 ,w__2967);
  nor g__3393(w__2993 ,w__2980 ,w__2971);
  or g__3394(w__2992 ,w__2665 ,w__2968);
  or g__3395(w__2991 ,w__2979 ,w__2970);
  or g__3396(w__4277 ,w__2926 ,w__2965);
  nor g__3397(w__2990 ,w__2932 ,w__2973);
  or g__3398(w__4254 ,w__2931 ,w__2974);
  and g__3399(w__2996 ,w__2933 ,w__2975);
  and g__3400(w__2995 ,w__2958 ,w__2978);
  not g__3401(w__2985 ,w__2986);
  and g__3402(w__2984 ,w__2942 ,w__2967);
  and g__3403(w__2983 ,w__2921 ,w__2972);
  nor g__3404(w__2982 ,w__2661 ,w__2969);
  xor g__3405(w__4247 ,w__2963 ,w__2944);
  xnor g__3406(w__4286 ,w__2954 ,w__2950);
  xnor g__3407(w__2981 ,w__2959 ,w__2952);
  xnor g__3408(w__2989 ,w__2943 ,w__2951);
  xnor g__3409(w__2988 ,w__2871 ,w__2945);
  xnor g__3410(w__2987 ,w__2964 ,w__2947);
  xnor g__3411(w__2986 ,w__2928 ,w__2949);
  not g__3412(w__2980 ,w__2979);
  or g__3413(w__2978 ,w__2872 ,w__2955);
  and g__3414(w__2977 ,w__2959 ,w__2953);
  nor g__3415(w__2976 ,w__2959 ,w__2953);
  or g__3416(w__2975 ,w__2929 ,w__2964);
  and g__3417(w__2974 ,w__2930 ,w__2954);
  or g__3418(w__2979 ,w__2937 ,w__2956);
  not g__3419(w__2970 ,w__2971);
  not g__3420(w__2968 ,w__2969);
  nor g__3421(w__2965 ,w__2925 ,w__2963);
  xnor g__3422(w__2973 ,w__2897 ,w__2919);
  xnor g__3423(w__2972 ,w__2893 ,w__2918);
  xnor g__3424(w__2971 ,w__2894 ,w__2920);
  and g__3425(w__2969 ,w__2927 ,w__2957);
  xnor g__3426(w__2967 ,w__2892 ,w__2917);
  xnor g__3427(w__2966 ,w__2895 ,w__2916);
  not g__3428(w__2961 ,w__2962);
  or g__3429(w__2958 ,w__2881 ,w__2928);
  or g__3430(w__2957 ,w__2943 ,w__2939);
  nor g__3431(w__2956 ,w__2871 ,w__2936);
  and g__3432(w__2955 ,w__2881 ,w__2928);
  or g__3433(w__4255 ,w__2852 ,w__2934);
  and g__3434(w__2964 ,w__2904 ,w__2924);
  and g__3435(w__2963 ,w__2902 ,w__2940);
  and g__3436(w__2962 ,w__2900 ,w__2923);
  and g__3437(w__2960 ,w__2911 ,w__2938);
  and g__3438(w__2959 ,w__2908 ,w__2935);
  not g__3439(w__2953 ,w__2952);
  xnor g__3440(w__4287 ,w__2896 ,w__2898);
  xnor g__3441(w__2951 ,w__2880 ,w__2877);
  xnor g__3442(w__2950 ,w__2887 ,w__2858);
  xnor g__3443(w__2949 ,w__2881 ,w__2872);
  xnor g__3444(w__2948 ,w__2913 ,w__2890);
  xnor g__3445(w__2947 ,w__2860 ,w__2885);
  xnor g__3446(w__2946 ,w__2889 ,w__2915);
  xnor g__3447(w__2945 ,w__2883 ,w__2882);
  xnor g__3448(w__2944 ,w__2878 ,w__2855);
  xnor g__3449(w__2954 ,w__2808 ,w__2875);
  xnor g__3450(w__2952 ,w__2873 ,w__2899);
  nor g__3451(w__2941 ,w__2913 ,w__2891);
  or g__3452(w__2940 ,w__2906 ,w__2892);
  nor g__3453(w__2939 ,w__2879 ,w__2877);
  or g__3454(w__2938 ,w__2895 ,w__2910);
  nor g__3455(w__2937 ,w__2882 ,w__2883);
  and g__3456(w__2936 ,w__2882 ,w__2883);
  or g__3457(w__2935 ,w__2907 ,w__2897);
  nor g__3458(w__2934 ,w__2863 ,w__2896);
  or g__3459(w__2933 ,w__2859 ,w__2885);
  and g__3460(w__2932 ,w__2913 ,w__2891);
  nor g__3461(w__2931 ,w__2858 ,w__2887);
  or g__3462(w__2930 ,w__2857 ,w__2886);
  nor g__3463(w__2929 ,w__2860 ,w__2884);
  and g__3464(w__2943 ,w__2851 ,w__2903);
  and g__3465(w__2942 ,w__2804 ,w__2912);
  or g__3466(w__2927 ,w__2880 ,w__2876);
  nor g__3467(w__2926 ,w__2855 ,w__2878);
  and g__3468(w__2925 ,w__2855 ,w__2878);
  or g__3469(w__2924 ,w__2894 ,w__2909);
  or g__3470(w__2923 ,w__2905 ,w__2893);
  nor g__3471(w__2922 ,w__2915 ,w__2889);
  or g__3472(w__2921 ,w__2914 ,w__2888);
  or g__3473(w__4276 ,w__2768 ,w__2901);
  xor g__3474(w__4246 ,w__2862 ,w__2822);
  xnor g__3475(w__2920 ,w__2861 ,w__2853);
  xnor g__3476(w__2919 ,w__2868 ,w__2566);
  xnor g__3477(w__2918 ,w__2784 ,w__2870);
  xnor g__3478(w__2917 ,w__2723 ,w__2856);
  xnor g__3479(w__2916 ,w__2867 ,w__2854);
  xnor g__3480(w__2928 ,w__2874 ,w__2823);
  not g__3481(w__2914 ,w__2915);
  or g__3482(w__2912 ,w__2766 ,w__2874);
  or g__3483(w__2911 ,w__2854 ,w__2867);
  and g__3484(w__2910 ,w__2854 ,w__2867);
  and g__3485(w__2909 ,w__2853 ,w__2861);
  or g__3486(w__2908 ,w__2566 ,w__2868);
  and g__3487(w__2907 ,w__2566 ,w__2868);
  and g__3488(w__2906 ,w__2723 ,w__2856);
  nor g__3489(w__2905 ,w__2784 ,w__2869);
  or g__3490(w__2904 ,w__2853 ,w__2861);
  or g__3491(w__2903 ,w__2873 ,w__2864);
  or g__3492(w__4256 ,w__2767 ,w__2850);
  or g__3493(w__2902 ,w__2723 ,w__2856);
  nor g__3494(w__2901 ,w__2782 ,w__2862);
  or g__3495(w__2900 ,w__2783 ,w__2870);
  xnor g__3496(w__2899 ,w__2806 ,w__2849);
  xnor g__3497(w__2898 ,w__2785 ,w__2567);
  and g__3498(w__2915 ,w__2789 ,w__2865);
  and g__3499(w__2913 ,w__2840 ,w__2866);
  not g__3500(w__2891 ,w__2890);
  not g__3501(w__2888 ,w__2889);
  not g__3502(w__2886 ,w__2887);
  not g__3503(w__2884 ,w__2885);
  not g__3504(w__2879 ,w__2880);
  not g__3505(w__2876 ,w__2877);
  xor g__3506(w__4288 ,w__2569 ,w__2829);
  xnor g__3507(w__2875 ,w__2702 ,w__2570);
  xnor g__3508(w__2897 ,w__2747 ,w__2830);
  xnor g__3509(w__2896 ,w__2753 ,w__2812);
  xnor g__3510(w__2895 ,w__2755 ,w__2826);
  xnor g__3511(w__2894 ,w__2736 ,w__2821);
  xnor g__3512(w__2893 ,w__2729 ,w__2819);
  xnor g__3513(w__2892 ,w__2726 ,w__2818);
  xnor g__3514(w__2890 ,w__2809 ,w__2815);
  xnor g__3515(w__2889 ,w__2704 ,w__2828);
  xnor g__3516(w__2887 ,w__2709 ,w__2814);
  xnor g__3517(w__2885 ,w__2568 ,w__2813);
  xnor g__3518(w__2883 ,w__2699 ,w__2824);
  xnor g__3519(w__2882 ,w__2689 ,w__2825);
  xnor g__3520(w__2881 ,w__2724 ,w__2827);
  xnor g__3521(w__2880 ,w__2754 ,w__2820);
  xnor g__3522(w__2878 ,w__2728 ,w__2816);
  xnor g__3523(w__2877 ,w__2811 ,w__2817);
  not g__3524(w__2869 ,w__2870);
  or g__3525(w__2866 ,w__2847 ,w__2570);
  or g__3526(w__2865 ,w__2796 ,w__2568);
  nor g__3527(w__2864 ,w__2806 ,w__2848);
  and g__3528(w__2863 ,w__2786 ,w__2567);
  and g__3529(w__2874 ,w__2794 ,w__2846);
  and g__3530(w__2873 ,w__2801 ,w__2838);
  and g__3531(w__2872 ,w__2795 ,w__2836);
  and g__3532(w__2871 ,w__2781 ,w__2844);
  and g__3533(w__2870 ,w__2776 ,w__2839);
  and g__3534(w__2868 ,w__2778 ,w__2842);
  and g__3535(w__2867 ,w__2799 ,w__2831);
  not g__3536(w__2859 ,w__2860);
  not g__3537(w__2857 ,w__2858);
  nor g__3538(w__2852 ,w__2786 ,w__2567);
  or g__3539(w__2851 ,w__2805 ,w__2849);
  nor g__3540(w__2850 ,w__2792 ,w__2569);
  and g__3541(w__2862 ,w__2769 ,w__2843);
  and g__3542(w__2861 ,w__2764 ,w__2837);
  or g__3543(w__2860 ,w__2788 ,w__2835);
  and g__3544(w__2858 ,w__2774 ,w__2834);
  and g__3545(w__2856 ,w__2773 ,w__2845);
  and g__3546(w__2855 ,w__2765 ,w__2832);
  and g__3547(w__2854 ,w__2790 ,w__2841);
  and g__3548(w__2853 ,w__2797 ,w__2833);
  not g__3549(w__2848 ,w__2849);
  nor g__3550(w__2847 ,w__2701 ,w__2808);
  or g__3551(w__2846 ,w__2720 ,w__2779);
  or g__3552(w__2845 ,w__2719 ,w__2791);
  or g__3553(w__2844 ,w__2802 ,w__2810);
  or g__3554(w__2843 ,w__2712 ,w__2775);
  or g__3555(w__2842 ,w__2709 ,w__2780);
  or g__3556(w__2841 ,w__2754 ,w__2777);
  or g__3557(w__2840 ,w__2702 ,w__2807);
  or g__3558(w__2839 ,w__2755 ,w__2803);
  or g__3559(w__2838 ,w__2747 ,w__2798);
  or g__3560(w__2837 ,w__2717 ,w__2787);
  or g__3561(w__2836 ,w__2710 ,w__2771);
  and g__3562(w__2835 ,w__2793 ,w__2811);
  or g__3563(w__2834 ,w__2753 ,w__2770);
  or g__3564(w__2833 ,w__2756 ,w__2772);
  or g__3565(w__2832 ,w__2711 ,w__2763);
  xor g__3566(w__4289 ,w__2721 ,w__2761);
  or g__3567(w__2831 ,w__2750 ,w__2800);
  xnor g__3568(w__2830 ,w__2740 ,w__2743);
  xnor g__3569(w__2829 ,w__2725 ,w__2737);
  xnor g__3570(w__2849 ,w__2757 ,w__2745);
  xnor g__3571(w__2828 ,w__2698 ,w__2710);
  xnor g__3572(w__2827 ,w__2703 ,w__2719);
  xnor g__3573(w__2826 ,w__2700 ,w__2731);
  xnor g__3574(w__2825 ,w__2697 ,w__2717);
  xnor g__3575(w__2824 ,w__2692 ,w__2756);
  xnor g__3576(w__2823 ,w__2690 ,w__2695);
  xnor g__3577(w__2822 ,w__2744 ,w__2738);
  xnor g__3578(w__2821 ,w__2696 ,w__2750);
  xnor g__3579(w__2820 ,w__2694 ,w__2732);
  xnor g__3580(w__2819 ,w__2742 ,w__2720);
  xnor g__3581(w__2818 ,w__2741 ,w__2711);
  xnor g__3582(w__2817 ,w__2688 ,w__2706);
  xnor g__3583(w__2816 ,w__2693 ,w__2712);
  xnor g__3584(w__2815 ,w__2722 ,w__2730);
  xnor g__3585(w__2814 ,w__2727 ,w__2735);
  xnor g__3586(w__2813 ,w__2691 ,w__2734);
  xnor g__3587(w__2812 ,w__2739 ,w__2733);
  not g__3588(w__2810 ,w__2809);
  not g__3589(w__2807 ,w__2808);
  not g__3590(w__2805 ,w__2806);
  or g__3591(w__2804 ,w__2690 ,w__2695);
  and g__3592(w__2803 ,w__2700 ,w__2731);
  and g__3593(w__2802 ,w__2722 ,w__2730);
  or g__3594(w__2801 ,w__2740 ,w__2743);
  and g__3595(w__2800 ,w__2736 ,w__2696);
  or g__3596(w__2799 ,w__2736 ,w__2696);
  and g__3597(w__2798 ,w__2740 ,w__2743);
  or g__3598(w__2797 ,w__2699 ,w__2692);
  and g__3599(w__2796 ,w__2691 ,w__2734);
  or g__3600(w__2795 ,w__2704 ,w__2698);
  or g__3601(w__2794 ,w__2729 ,w__2742);
  or g__3602(w__2793 ,w__2687 ,w__2705);
  and g__3603(w__2792 ,w__2725 ,w__2737);
  and g__3604(w__2791 ,w__2724 ,w__2703);
  or g__3605(w__2790 ,w__2694 ,w__2732);
  or g__3606(w__2789 ,w__2691 ,w__2734);
  nor g__3607(w__2788 ,w__2688 ,w__2706);
  and g__3608(w__2787 ,w__2697 ,w__2689);
  and g__3609(w__2811 ,w__2758 ,w__2746);
  and g__3610(w__2809 ,w__2707 ,w__2718);
  and g__3611(w__2808 ,w__2752 ,w__2714);
  and g__3612(w__2806 ,w__2749 ,w__2708);
  not g__3613(w__2786 ,w__2785);
  not g__3614(w__2783 ,w__2784);
  and g__3615(w__2782 ,w__2744 ,w__2738);
  or g__3616(w__2781 ,w__2722 ,w__2730);
  and g__3617(w__2780 ,w__2727 ,w__2735);
  and g__3618(w__2779 ,w__2729 ,w__2742);
  or g__3619(w__2778 ,w__2727 ,w__2735);
  and g__3620(w__2777 ,w__2694 ,w__2732);
  or g__3621(w__2776 ,w__2700 ,w__2731);
  and g__3622(w__2775 ,w__2728 ,w__2693);
  or g__3623(w__2774 ,w__2739 ,w__2733);
  or g__3624(w__2773 ,w__2724 ,w__2703);
  and g__3625(w__2772 ,w__2699 ,w__2692);
  and g__3626(w__2771 ,w__2704 ,w__2698);
  and g__3627(w__2770 ,w__2739 ,w__2733);
  or g__3628(w__2769 ,w__2728 ,w__2693);
  nor g__3629(w__2768 ,w__2744 ,w__2738);
  nor g__3630(w__2767 ,w__2725 ,w__2737);
  and g__3631(w__2766 ,w__2690 ,w__2695);
  or g__3632(w__2765 ,w__2726 ,w__2741);
  or g__3633(w__2764 ,w__2697 ,w__2689);
  and g__3634(w__2763 ,w__2726 ,w__2741);
  nor g__3635(w__2762 ,w__2761 ,w__2721);
  and g__3636(w__2785 ,w__2760 ,w__2716);
  and g__3637(w__2784 ,w__2715 ,w__2713);
  not g__3638(w__2760 ,w__2759);
  not g__3639(w__2758 ,w__2757);
  not g__3640(w__2752 ,w__2751);
  not g__3641(w__2749 ,w__2748);
  not g__3642(w__2746 ,w__2745);
  and g__3643(w__4245 ,in16[8] ,in17[7]);
  or g__3644(w__2761 ,w__2583 ,w__2676);
  or g__3645(w__2759 ,w__2623 ,w__2603);
  or g__3646(w__2757 ,w__2578 ,w__2646);
  or g__3647(w__2756 ,w__2585 ,w__2613);
  or g__3648(w__2755 ,w__2617 ,w__2628);
  or g__3649(w__2754 ,w__2617 ,w__2607);
  or g__3650(w__2753 ,w__2623 ,w__2608);
  or g__3651(w__2751 ,w__2597 ,w__2646);
  or g__3652(w__2750 ,w__2593 ,w__2604);
  or g__3653(w__2748 ,w__2635 ,w__2603);
  or g__3654(w__2747 ,w__2595 ,w__2614);
  or g__3655(w__2745 ,w__2599 ,w__2604);
  or g__3656(w__2744 ,w__2632 ,w__2643);
  or g__3657(w__2743 ,w__2588 ,w__2575);
  or g__3658(w__2742 ,w__2591 ,w__2625);
  or g__3659(w__2741 ,w__2632 ,w__2601);
  or g__3660(w__2740 ,w__2681 ,w__2637);
  or g__3661(w__2739 ,w__2605 ,w__2572);
  or g__3662(w__2738 ,w__2581 ,w__2619);
  or g__3663(w__2737 ,w__2653 ,w__2607);
  or g__3664(w__2736 ,w__2635 ,w__2660);
  or g__3665(w__2735 ,w__2622 ,w__2629);
  or g__3666(w__2734 ,w__2587 ,w__2620);
  or g__3667(w__2733 ,w__2650 ,w__2576);
  or g__3668(w__2732 ,w__2590 ,w__2658);
  or g__3669(w__2731 ,w__2674 ,w__2638);
  or g__3670(w__2730 ,w__2649 ,w__2611);
  or g__3671(w__2729 ,w__2673 ,w__2640);
  or g__3672(w__2728 ,w__2682 ,w__2641);
  or g__3673(w__2727 ,w__2652 ,w__2573);
  or g__3674(w__2726 ,w__2634 ,w__2644);
  or g__3675(w__2725 ,w__2655 ,w__2628);
  or g__3676(w__2724 ,w__2585 ,w__2626);
  or g__3677(w__2723 ,w__2616 ,w__2619);
  or g__3678(w__2722 ,w__2655 ,w__2625);
  not g__3679(w__2706 ,w__2705);
  not g__3680(w__2702 ,w__2701);
  not g__3681(w__2688 ,w__2687);
  nor g__3682(w__2686 ,w__2650 ,w__2558);
  nor g__3683(w__2685 ,w__2653 ,w__2560);
  nor g__3684(w__2684 ,w__2676 ,w__2562);
  nor g__3685(w__2683 ,w__2656 ,w__2647);
  or g__3686(w__2721 ,w__2605 ,w__2613);
  or g__3687(w__2720 ,w__2578 ,w__2637);
  or g__3688(w__2719 ,w__2580 ,w__2660);
  and g__3689(w__2718 ,in16[5] ,in17[0]);
  or g__3690(w__2717 ,w__2679 ,w__2629);
  and g__3691(w__2716 ,in16[3] ,in17[0]);
  and g__3692(w__2715 ,in16[7] ,in17[2]);
  and g__3693(w__2714 ,in16[4] ,in17[0]);
  and g__3694(w__2713 ,in16[8] ,in17[1]);
  or g__3695(w__2712 ,w__2678 ,w__2611);
  or g__3696(w__2711 ,w__2581 ,w__2658);
  or g__3697(w__2710 ,w__2593 ,w__2608);
  or g__3698(w__2709 ,w__2588 ,w__2614);
  and g__3699(w__2708 ,in16[6] ,in17[0]);
  and g__3700(w__2707 ,in16[4] ,in17[1]);
  and g__3701(w__2705 ,in16[3] ,in17[5]);
  or g__3702(w__2704 ,w__2634 ,w__2668);
  or g__3703(w__2703 ,w__2671 ,w__2638);
  and g__3704(w__2701 ,in16[0] ,in17[5]);
  or g__3705(w__2700 ,w__2591 ,w__2610);
  or g__3706(w__2699 ,w__2649 ,w__2620);
  or g__3707(w__2698 ,w__2631 ,w__2576);
  or g__3708(w__2697 ,w__2656 ,w__2640);
  or g__3709(w__2696 ,w__2599 ,w__2647);
  or g__3710(w__2695 ,w__2616 ,w__2601);
  or g__3711(w__2694 ,w__2652 ,w__2643);
  or g__3712(w__2693 ,w__2631 ,w__2626);
  or g__3713(w__2692 ,w__2583 ,w__2610);
  or g__3714(w__2691 ,w__2622 ,w__2641);
  or g__3715(w__2690 ,w__2595 ,w__2644);
  or g__3716(w__2689 ,w__2597 ,w__2573);
  and g__3717(w__2687 ,in16[2] ,in17[6]);
  not g__3718(w__2682 ,in16[6]);
  not g__3719(w__2681 ,in16[2]);
  not g__3720(w__2680 ,in16[1]);
  not g__3721(w__2679 ,in16[4]);
  not g__3722(w__2678 ,in16[8]);
  not g__3723(w__2677 ,in17[3]);
  not g__3724(w__2676 ,in17[0]);
  not g__3725(w__2675 ,in17[1]);
  not g__3726(w__2674 ,in16[5]);
  not g__3727(w__2673 ,in16[3]);
  not g__3728(w__2672 ,in16[0]);
  not g__3729(w__2671 ,in16[7]);
  not g__3730(w__2670 ,in17[4]);
  not g__3731(w__2669 ,in17[2]);
  not g__3732(w__2668 ,in17[5]);
  not g__3733(w__2667 ,in17[7]);
  not g__3734(w__2666 ,in17[6]);
  not g__3735(w__2565 ,w__2664);
  not g__3736(w__2664 ,w__2672);
  not g__3737(w__2564 ,w__2663);
  not g__3738(w__2557 ,w__2663);
  not g__3739(w__2663 ,w__2675);
  not g__3740(w__2563 ,w__2662);
  not g__3741(w__2662 ,w__2676);
  buf g__3742(w__4258 ,w__2686);
  buf g__3743(w__4290 ,w__2683);
  buf g__3744(w__4260 ,w__2684);
  buf g__3745(w__4259 ,w__2685);
  buf g__3746(w__4257 ,w__2762);
  not g__3747(w__2661 ,w__2665);
  not g__3748(w__2665 ,w__2966);
  not g__3749(w__2660 ,w__2659);
  not g__3750(w__2659 ,w__2677);
  not g__3751(w__2658 ,w__2657);
  not g__3752(w__2657 ,w__2670);
  not g__3753(w__2656 ,w__2654);
  not g__3754(w__2655 ,w__2654);
  not g__3755(w__2654 ,w__2672);
  not g__3756(w__2653 ,w__2651);
  not g__3757(w__2652 ,w__2651);
  not g__3758(w__2651 ,w__2680);
  not g__3759(w__2650 ,w__2648);
  not g__3760(w__2649 ,w__2648);
  not g__3761(w__2648 ,w__2680);
  not g__3762(w__2647 ,w__2645);
  not g__3763(w__2646 ,w__2645);
  not g__3764(w__2645 ,w__2564);
  not g__3765(w__2644 ,w__2642);
  not g__3766(w__2643 ,w__2642);
  not g__3767(w__2642 ,w__2667);
  not g__3768(w__2641 ,w__2639);
  not g__3769(w__2640 ,w__2639);
  not g__3770(w__2639 ,w__2667);
  not g__3771(w__2638 ,w__2636);
  not g__3772(w__2637 ,w__2636);
  not g__3773(w__2636 ,w__2670);
  not g__3774(w__2635 ,w__2633);
  not g__3775(w__2634 ,w__2633);
  not g__3776(w__2633 ,w__2674);
  not g__3777(w__2632 ,w__2630);
  not g__3778(w__2631 ,w__2630);
  not g__3779(w__2630 ,w__2671);
  not g__3780(w__2629 ,w__2627);
  not g__3781(w__2628 ,w__2627);
  not g__3782(w__2627 ,w__2677);
  not g__3783(w__2626 ,w__2624);
  not g__3784(w__2625 ,w__2624);
  not g__3785(w__2624 ,w__2666);
  not g__3786(w__2623 ,w__2621);
  not g__3787(w__2622 ,w__2621);
  not g__3788(w__2621 ,w__2681);
  not g__3789(w__2620 ,w__2618);
  not g__3790(w__2619 ,w__2618);
  not g__3791(w__2618 ,w__2666);
  not g__3792(w__2617 ,w__2615);
  not g__3793(w__2616 ,w__2615);
  not g__3794(w__2615 ,w__2682);
  not g__3795(w__2614 ,w__2612);
  not g__3796(w__2613 ,w__2612);
  not g__3797(w__2612 ,w__2669);
  not g__3798(w__2611 ,w__2609);
  not g__3799(w__2610 ,w__2609);
  not g__3800(w__2609 ,w__2668);
  not g__3801(w__2608 ,w__2606);
  not g__3802(w__2607 ,w__2606);
  not g__3803(w__2606 ,w__2669);
  not g__3804(w__2562 ,w__2561);
  not g__3805(w__2605 ,w__2561);
  not g__3806(w__2561 ,w__2565);
  not g__3807(w__2560 ,w__2559);
  not g__3808(w__2604 ,w__2559);
  not g__3809(w__2559 ,w__2563);
  not g__3810(w__2558 ,w__2602);
  not g__3811(w__2603 ,w__2602);
  not g__3812(w__2602 ,w__2557);
  not g__3813(w__2601 ,w__2600);
  not g__3814(w__2600 ,w__2668);
  not g__3815(w__2599 ,w__2598);
  not g__3816(w__2598 ,w__2671);
  not g__3817(w__2597 ,w__2596);
  not g__3818(w__2596 ,w__2673);
  not g__3819(w__2595 ,w__2594);
  not g__3820(w__2594 ,w__2679);
  not g__3821(w__2593 ,w__2592);
  not g__3822(w__2592 ,w__2678);
  not g__3823(w__2591 ,w__2589);
  not g__3824(w__2590 ,w__2589);
  not g__3825(w__2589 ,w__2679);
  not g__3826(w__2588 ,w__2586);
  not g__3827(w__2587 ,w__2586);
  not g__3828(w__2586 ,w__2673);
  not g__3829(w__2585 ,w__2584);
  not g__3830(w__2584 ,w__2674);
  not g__3831(w__2583 ,w__2582);
  not g__3832(w__2582 ,w__2681);
  not g__3833(w__2581 ,w__2579);
  not g__3834(w__2580 ,w__2579);
  not g__3835(w__2579 ,w__2678);
  not g__3836(w__2578 ,w__2577);
  not g__3837(w__2577 ,w__2682);
  not g__3838(w__2576 ,w__2574);
  not g__3839(w__2575 ,w__2574);
  not g__3840(w__2574 ,w__2677);
  not g__3841(w__2573 ,w__2571);
  not g__3842(w__2572 ,w__2571);
  not g__3843(w__2571 ,w__2670);
  xnor g__3844(w__2570 ,w__2707 ,w__2718);
  xor g__3845(w__2569 ,w__2759 ,w__2716);
  xnor g__3846(w__2568 ,w__2715 ,w__2713);
  xor g__3847(w__2567 ,w__2751 ,w__2714);
  xor g__3848(w__2566 ,w__2748 ,w__2708);
  xnor g__3849(w__4217 ,w__3454 ,w__3471);
  or g__3850(w__4184 ,w__3470 ,w__3472);
  xnor g__3851(w__4216 ,w__3466 ,w__3467);
  nor g__3852(w__3472 ,w__3454 ,w__3469);
  or g__3853(w__4215 ,w__3462 ,w__3468);
  xnor g__3854(w__3471 ,w__3418 ,w__3460);
  xnor g__3855(w__4218 ,w__3445 ,w__3457);
  xnor g__3856(w__4219 ,w__3447 ,w__3456);
  xor g__3857(w__4183 ,w__3453 ,w__3455);
  or g__3858(w__4186 ,w__3451 ,w__3464);
  nor g__3859(w__3470 ,w__3418 ,w__3461);
  or g__3860(w__4214 ,w__3452 ,w__3463);
  and g__3861(w__3469 ,w__3418 ,w__3461);
  and g__3862(w__3468 ,w__3466 ,w__3458);
  or g__3863(w__4185 ,w__3440 ,w__3465);
  or g__3864(w__4187 ,w__3434 ,w__3459);
  xnor g__3865(w__4220 ,w__3446 ,w__3439);
  xnor g__3866(w__3467 ,w__3444 ,w__3420);
  and g__3867(w__3465 ,w__3450 ,w__3445);
  and g__3868(w__3464 ,w__3449 ,w__3447);
  or g__3869(w__4188 ,w__3399 ,w__3448);
  nor g__3870(w__3463 ,w__3442 ,w__3453);
  nor g__3871(w__3462 ,w__3420 ,w__3444);
  or g__3872(w__3466 ,w__3380 ,w__3441);
  not g__3873(w__3461 ,w__3460);
  nor g__3874(w__3459 ,w__3435 ,w__3446);
  or g__3875(w__3458 ,w__3419 ,w__3443);
  xnor g__3876(w__4221 ,w__3431 ,w__3406);
  xnor g__3877(w__3457 ,w__3427 ,w__3424);
  xnor g__3878(w__3456 ,w__3429 ,w__3438);
  xnor g__3879(w__3455 ,w__3425 ,w__3400);
  xnor g__3880(w__3460 ,w__3430 ,w__3404);
  nor g__3881(w__3452 ,w__3400 ,w__3425);
  nor g__3882(w__3451 ,w__3438 ,w__3429);
  or g__3883(w__3450 ,w__3123 ,w__3426);
  or g__3884(w__3449 ,w__3437 ,w__3428);
  or g__3885(w__4213 ,w__3384 ,w__3423);
  nor g__3886(w__3448 ,w__3390 ,w__3431);
  or g__3887(w__4189 ,w__3389 ,w__3432);
  and g__3888(w__3454 ,w__3391 ,w__3433);
  and g__3889(w__3453 ,w__3416 ,w__3436);
  not g__3890(w__3443 ,w__3444);
  and g__3891(w__3442 ,w__3400 ,w__3425);
  and g__3892(w__3441 ,w__3379 ,w__3430);
  nor g__3893(w__3440 ,w__3119 ,w__3427);
  xor g__3894(w__4182 ,w__3421 ,w__3402);
  xnor g__3895(w__4222 ,w__3412 ,w__3408);
  xnor g__3896(w__3439 ,w__3417 ,w__3410);
  xnor g__3897(w__3447 ,w__3401 ,w__3409);
  xnor g__3898(w__3446 ,w__3329 ,w__3403);
  xnor g__3899(w__3445 ,w__3422 ,w__3405);
  xnor g__3900(w__3444 ,w__3386 ,w__3407);
  not g__3901(w__3438 ,w__3437);
  or g__3902(w__3436 ,w__3330 ,w__3413);
  and g__3903(w__3435 ,w__3417 ,w__3411);
  nor g__3904(w__3434 ,w__3417 ,w__3411);
  or g__3905(w__3433 ,w__3387 ,w__3422);
  and g__3906(w__3432 ,w__3388 ,w__3412);
  or g__3907(w__3437 ,w__3395 ,w__3414);
  not g__3908(w__3428 ,w__3429);
  not g__3909(w__3426 ,w__3427);
  nor g__3910(w__3423 ,w__3383 ,w__3421);
  xnor g__3911(w__3431 ,w__3355 ,w__3377);
  xnor g__3912(w__3430 ,w__3351 ,w__3376);
  xnor g__3913(w__3429 ,w__3352 ,w__3378);
  and g__3914(w__3427 ,w__3385 ,w__3415);
  xnor g__3915(w__3425 ,w__3350 ,w__3375);
  xnor g__3916(w__3424 ,w__3353 ,w__3374);
  not g__3917(w__3419 ,w__3420);
  or g__3918(w__3416 ,w__3339 ,w__3386);
  or g__3919(w__3415 ,w__3401 ,w__3397);
  nor g__3920(w__3414 ,w__3329 ,w__3394);
  and g__3921(w__3413 ,w__3339 ,w__3386);
  or g__3922(w__4190 ,w__3310 ,w__3392);
  and g__3923(w__3422 ,w__3362 ,w__3382);
  and g__3924(w__3421 ,w__3360 ,w__3398);
  and g__3925(w__3420 ,w__3358 ,w__3381);
  and g__3926(w__3418 ,w__3369 ,w__3396);
  and g__3927(w__3417 ,w__3366 ,w__3393);
  not g__3928(w__3411 ,w__3410);
  xnor g__3929(w__4223 ,w__3354 ,w__3356);
  xnor g__3930(w__3409 ,w__3338 ,w__3335);
  xnor g__3931(w__3408 ,w__3345 ,w__3316);
  xnor g__3932(w__3407 ,w__3339 ,w__3330);
  xnor g__3933(w__3406 ,w__3371 ,w__3348);
  xnor g__3934(w__3405 ,w__3318 ,w__3343);
  xnor g__3935(w__3404 ,w__3347 ,w__3373);
  xnor g__3936(w__3403 ,w__3341 ,w__3340);
  xnor g__3937(w__3402 ,w__3336 ,w__3313);
  xnor g__3938(w__3412 ,w__3266 ,w__3333);
  xnor g__3939(w__3410 ,w__3331 ,w__3357);
  nor g__3940(w__3399 ,w__3371 ,w__3349);
  or g__3941(w__3398 ,w__3364 ,w__3350);
  nor g__3942(w__3397 ,w__3337 ,w__3335);
  or g__3943(w__3396 ,w__3353 ,w__3368);
  nor g__3944(w__3395 ,w__3340 ,w__3341);
  and g__3945(w__3394 ,w__3340 ,w__3341);
  or g__3946(w__3393 ,w__3365 ,w__3355);
  nor g__3947(w__3392 ,w__3321 ,w__3354);
  or g__3948(w__3391 ,w__3317 ,w__3343);
  and g__3949(w__3390 ,w__3371 ,w__3349);
  nor g__3950(w__3389 ,w__3316 ,w__3345);
  or g__3951(w__3388 ,w__3315 ,w__3344);
  nor g__3952(w__3387 ,w__3318 ,w__3342);
  and g__3953(w__3401 ,w__3309 ,w__3361);
  and g__3954(w__3400 ,w__3262 ,w__3370);
  or g__3955(w__3385 ,w__3338 ,w__3334);
  nor g__3956(w__3384 ,w__3313 ,w__3336);
  and g__3957(w__3383 ,w__3313 ,w__3336);
  or g__3958(w__3382 ,w__3352 ,w__3367);
  or g__3959(w__3381 ,w__3363 ,w__3351);
  nor g__3960(w__3380 ,w__3373 ,w__3347);
  or g__3961(w__3379 ,w__3372 ,w__3346);
  or g__3962(w__4212 ,w__3226 ,w__3359);
  xor g__3963(w__4181 ,w__3320 ,w__3280);
  xnor g__3964(w__3378 ,w__3319 ,w__3311);
  xnor g__3965(w__3377 ,w__3326 ,w__3024);
  xnor g__3966(w__3376 ,w__3242 ,w__3328);
  xnor g__3967(w__3375 ,w__3181 ,w__3314);
  xnor g__3968(w__3374 ,w__3325 ,w__3312);
  xnor g__3969(w__3386 ,w__3332 ,w__3281);
  not g__3970(w__3372 ,w__3373);
  or g__3971(w__3370 ,w__3224 ,w__3332);
  or g__3972(w__3369 ,w__3312 ,w__3325);
  and g__3973(w__3368 ,w__3312 ,w__3325);
  and g__3974(w__3367 ,w__3311 ,w__3319);
  or g__3975(w__3366 ,w__3024 ,w__3326);
  and g__3976(w__3365 ,w__3024 ,w__3326);
  and g__3977(w__3364 ,w__3181 ,w__3314);
  nor g__3978(w__3363 ,w__3242 ,w__3327);
  or g__3979(w__3362 ,w__3311 ,w__3319);
  or g__3980(w__3361 ,w__3331 ,w__3322);
  or g__3981(w__4191 ,w__3225 ,w__3308);
  or g__3982(w__3360 ,w__3181 ,w__3314);
  nor g__3983(w__3359 ,w__3240 ,w__3320);
  or g__3984(w__3358 ,w__3241 ,w__3328);
  xnor g__3985(w__3357 ,w__3264 ,w__3307);
  xnor g__3986(w__3356 ,w__3243 ,w__3025);
  and g__3987(w__3373 ,w__3247 ,w__3323);
  and g__3988(w__3371 ,w__3298 ,w__3324);
  not g__3989(w__3349 ,w__3348);
  not g__3990(w__3346 ,w__3347);
  not g__3991(w__3344 ,w__3345);
  not g__3992(w__3342 ,w__3343);
  not g__3993(w__3337 ,w__3338);
  not g__3994(w__3334 ,w__3335);
  xor g__3995(w__4224 ,w__3027 ,w__3287);
  xnor g__3996(w__3333 ,w__3160 ,w__3028);
  xnor g__3997(w__3355 ,w__3205 ,w__3288);
  xnor g__3998(w__3354 ,w__3211 ,w__3270);
  xnor g__3999(w__3353 ,w__3213 ,w__3284);
  xnor g__4000(w__3352 ,w__3194 ,w__3279);
  xnor g__4001(w__3351 ,w__3187 ,w__3277);
  xnor g__4002(w__3350 ,w__3184 ,w__3276);
  xnor g__4003(w__3348 ,w__3267 ,w__3273);
  xnor g__4004(w__3347 ,w__3162 ,w__3286);
  xnor g__4005(w__3345 ,w__3167 ,w__3272);
  xnor g__4006(w__3343 ,w__3026 ,w__3271);
  xnor g__4007(w__3341 ,w__3157 ,w__3282);
  xnor g__4008(w__3340 ,w__3147 ,w__3283);
  xnor g__4009(w__3339 ,w__3182 ,w__3285);
  xnor g__4010(w__3338 ,w__3212 ,w__3278);
  xnor g__4011(w__3336 ,w__3186 ,w__3274);
  xnor g__4012(w__3335 ,w__3269 ,w__3275);
  not g__4013(w__3327 ,w__3328);
  or g__4014(w__3324 ,w__3305 ,w__3028);
  or g__4015(w__3323 ,w__3254 ,w__3026);
  nor g__4016(w__3322 ,w__3264 ,w__3306);
  and g__4017(w__3321 ,w__3244 ,w__3025);
  and g__4018(w__3332 ,w__3252 ,w__3304);
  and g__4019(w__3331 ,w__3259 ,w__3296);
  and g__4020(w__3330 ,w__3253 ,w__3294);
  and g__4021(w__3329 ,w__3239 ,w__3302);
  and g__4022(w__3328 ,w__3234 ,w__3297);
  and g__4023(w__3326 ,w__3236 ,w__3300);
  and g__4024(w__3325 ,w__3257 ,w__3289);
  not g__4025(w__3317 ,w__3318);
  not g__4026(w__3315 ,w__3316);
  nor g__4027(w__3310 ,w__3244 ,w__3025);
  or g__4028(w__3309 ,w__3263 ,w__3307);
  nor g__4029(w__3308 ,w__3250 ,w__3027);
  and g__4030(w__3320 ,w__3227 ,w__3301);
  and g__4031(w__3319 ,w__3222 ,w__3295);
  or g__4032(w__3318 ,w__3246 ,w__3293);
  and g__4033(w__3316 ,w__3232 ,w__3292);
  and g__4034(w__3314 ,w__3231 ,w__3303);
  and g__4035(w__3313 ,w__3223 ,w__3290);
  and g__4036(w__3312 ,w__3248 ,w__3299);
  and g__4037(w__3311 ,w__3255 ,w__3291);
  not g__4038(w__3306 ,w__3307);
  nor g__4039(w__3305 ,w__3159 ,w__3266);
  or g__4040(w__3304 ,w__3178 ,w__3237);
  or g__4041(w__3303 ,w__3177 ,w__3249);
  or g__4042(w__3302 ,w__3260 ,w__3268);
  or g__4043(w__3301 ,w__3170 ,w__3233);
  or g__4044(w__3300 ,w__3167 ,w__3238);
  or g__4045(w__3299 ,w__3212 ,w__3235);
  or g__4046(w__3298 ,w__3160 ,w__3265);
  or g__4047(w__3297 ,w__3213 ,w__3261);
  or g__4048(w__3296 ,w__3205 ,w__3256);
  or g__4049(w__3295 ,w__3175 ,w__3245);
  or g__4050(w__3294 ,w__3168 ,w__3229);
  and g__4051(w__3293 ,w__3251 ,w__3269);
  or g__4052(w__3292 ,w__3211 ,w__3228);
  or g__4053(w__3291 ,w__3214 ,w__3230);
  or g__4054(w__3290 ,w__3169 ,w__3221);
  xor g__4055(w__4225 ,w__3179 ,w__3219);
  or g__4056(w__3289 ,w__3208 ,w__3258);
  xnor g__4057(w__3288 ,w__3198 ,w__3201);
  xnor g__4058(w__3287 ,w__3183 ,w__3195);
  xnor g__4059(w__3307 ,w__3215 ,w__3203);
  xnor g__4060(w__3286 ,w__3156 ,w__3168);
  xnor g__4061(w__3285 ,w__3161 ,w__3177);
  xnor g__4062(w__3284 ,w__3158 ,w__3189);
  xnor g__4063(w__3283 ,w__3155 ,w__3175);
  xnor g__4064(w__3282 ,w__3150 ,w__3214);
  xnor g__4065(w__3281 ,w__3148 ,w__3153);
  xnor g__4066(w__3280 ,w__3202 ,w__3196);
  xnor g__4067(w__3279 ,w__3154 ,w__3208);
  xnor g__4068(w__3278 ,w__3152 ,w__3190);
  xnor g__4069(w__3277 ,w__3200 ,w__3178);
  xnor g__4070(w__3276 ,w__3199 ,w__3169);
  xnor g__4071(w__3275 ,w__3146 ,w__3164);
  xnor g__4072(w__3274 ,w__3151 ,w__3170);
  xnor g__4073(w__3273 ,w__3180 ,w__3188);
  xnor g__4074(w__3272 ,w__3185 ,w__3193);
  xnor g__4075(w__3271 ,w__3149 ,w__3192);
  xnor g__4076(w__3270 ,w__3197 ,w__3191);
  not g__4077(w__3268 ,w__3267);
  not g__4078(w__3265 ,w__3266);
  not g__4079(w__3263 ,w__3264);
  or g__4080(w__3262 ,w__3148 ,w__3153);
  and g__4081(w__3261 ,w__3158 ,w__3189);
  and g__4082(w__3260 ,w__3180 ,w__3188);
  or g__4083(w__3259 ,w__3198 ,w__3201);
  and g__4084(w__3258 ,w__3194 ,w__3154);
  or g__4085(w__3257 ,w__3194 ,w__3154);
  and g__4086(w__3256 ,w__3198 ,w__3201);
  or g__4087(w__3255 ,w__3157 ,w__3150);
  and g__4088(w__3254 ,w__3149 ,w__3192);
  or g__4089(w__3253 ,w__3162 ,w__3156);
  or g__4090(w__3252 ,w__3187 ,w__3200);
  or g__4091(w__3251 ,w__3145 ,w__3163);
  and g__4092(w__3250 ,w__3183 ,w__3195);
  and g__4093(w__3249 ,w__3182 ,w__3161);
  or g__4094(w__3248 ,w__3152 ,w__3190);
  or g__4095(w__3247 ,w__3149 ,w__3192);
  nor g__4096(w__3246 ,w__3146 ,w__3164);
  and g__4097(w__3245 ,w__3155 ,w__3147);
  and g__4098(w__3269 ,w__3216 ,w__3204);
  and g__4099(w__3267 ,w__3165 ,w__3176);
  and g__4100(w__3266 ,w__3210 ,w__3172);
  and g__4101(w__3264 ,w__3207 ,w__3166);
  not g__4102(w__3244 ,w__3243);
  not g__4103(w__3241 ,w__3242);
  and g__4104(w__3240 ,w__3202 ,w__3196);
  or g__4105(w__3239 ,w__3180 ,w__3188);
  and g__4106(w__3238 ,w__3185 ,w__3193);
  and g__4107(w__3237 ,w__3187 ,w__3200);
  or g__4108(w__3236 ,w__3185 ,w__3193);
  and g__4109(w__3235 ,w__3152 ,w__3190);
  or g__4110(w__3234 ,w__3158 ,w__3189);
  and g__4111(w__3233 ,w__3186 ,w__3151);
  or g__4112(w__3232 ,w__3197 ,w__3191);
  or g__4113(w__3231 ,w__3182 ,w__3161);
  and g__4114(w__3230 ,w__3157 ,w__3150);
  and g__4115(w__3229 ,w__3162 ,w__3156);
  and g__4116(w__3228 ,w__3197 ,w__3191);
  or g__4117(w__3227 ,w__3186 ,w__3151);
  nor g__4118(w__3226 ,w__3202 ,w__3196);
  nor g__4119(w__3225 ,w__3183 ,w__3195);
  and g__4120(w__3224 ,w__3148 ,w__3153);
  or g__4121(w__3223 ,w__3184 ,w__3199);
  or g__4122(w__3222 ,w__3155 ,w__3147);
  and g__4123(w__3221 ,w__3184 ,w__3199);
  nor g__4124(w__3220 ,w__3219 ,w__3179);
  and g__4125(w__3243 ,w__3218 ,w__3174);
  and g__4126(w__3242 ,w__3173 ,w__3171);
  not g__4127(w__3218 ,w__3217);
  not g__4128(w__3216 ,w__3215);
  not g__4129(w__3210 ,w__3209);
  not g__4130(w__3207 ,w__3206);
  not g__4131(w__3204 ,w__3203);
  and g__4132(w__4180 ,in20[8] ,in21[7]);
  or g__4133(w__3219 ,w__3041 ,w__3134);
  or g__4134(w__3217 ,w__3081 ,w__3061);
  or g__4135(w__3215 ,w__3036 ,w__3104);
  or g__4136(w__3214 ,w__3043 ,w__3071);
  or g__4137(w__3213 ,w__3075 ,w__3086);
  or g__4138(w__3212 ,w__3075 ,w__3065);
  or g__4139(w__3211 ,w__3081 ,w__3066);
  or g__4140(w__3209 ,w__3055 ,w__3104);
  or g__4141(w__3208 ,w__3051 ,w__3062);
  or g__4142(w__3206 ,w__3093 ,w__3061);
  or g__4143(w__3205 ,w__3053 ,w__3072);
  or g__4144(w__3203 ,w__3057 ,w__3062);
  or g__4145(w__3202 ,w__3090 ,w__3101);
  or g__4146(w__3201 ,w__3046 ,w__3033);
  or g__4147(w__3200 ,w__3049 ,w__3083);
  or g__4148(w__3199 ,w__3090 ,w__3059);
  or g__4149(w__3198 ,w__3139 ,w__3095);
  or g__4150(w__3197 ,w__3063 ,w__3030);
  or g__4151(w__3196 ,w__3039 ,w__3077);
  or g__4152(w__3195 ,w__3111 ,w__3065);
  or g__4153(w__3194 ,w__3093 ,w__3118);
  or g__4154(w__3193 ,w__3080 ,w__3087);
  or g__4155(w__3192 ,w__3045 ,w__3078);
  or g__4156(w__3191 ,w__3108 ,w__3034);
  or g__4157(w__3190 ,w__3048 ,w__3116);
  or g__4158(w__3189 ,w__3132 ,w__3096);
  or g__4159(w__3188 ,w__3107 ,w__3069);
  or g__4160(w__3187 ,w__3131 ,w__3098);
  or g__4161(w__3186 ,w__3140 ,w__3099);
  or g__4162(w__3185 ,w__3110 ,w__3031);
  or g__4163(w__3184 ,w__3092 ,w__3102);
  or g__4164(w__3183 ,w__3113 ,w__3086);
  or g__4165(w__3182 ,w__3043 ,w__3084);
  or g__4166(w__3181 ,w__3074 ,w__3077);
  or g__4167(w__3180 ,w__3113 ,w__3083);
  not g__4168(w__3164 ,w__3163);
  not g__4169(w__3160 ,w__3159);
  not g__4170(w__3146 ,w__3145);
  nor g__4171(w__3144 ,w__3108 ,w__3016);
  nor g__4172(w__3143 ,w__3111 ,w__3018);
  nor g__4173(w__3142 ,w__3134 ,w__3020);
  nor g__4174(w__3141 ,w__3114 ,w__3105);
  or g__4175(w__3179 ,w__3063 ,w__3071);
  or g__4176(w__3178 ,w__3036 ,w__3095);
  or g__4177(w__3177 ,w__3038 ,w__3118);
  and g__4178(w__3176 ,in20[5] ,in21[0]);
  or g__4179(w__3175 ,w__3137 ,w__3087);
  and g__4180(w__3174 ,in20[3] ,in21[0]);
  and g__4181(w__3173 ,in20[7] ,in21[2]);
  and g__4182(w__3172 ,in20[4] ,in21[0]);
  and g__4183(w__3171 ,in20[8] ,in21[1]);
  or g__4184(w__3170 ,w__3136 ,w__3069);
  or g__4185(w__3169 ,w__3039 ,w__3116);
  or g__4186(w__3168 ,w__3051 ,w__3066);
  or g__4187(w__3167 ,w__3046 ,w__3072);
  and g__4188(w__3166 ,in20[6] ,in21[0]);
  and g__4189(w__3165 ,in20[4] ,in21[1]);
  and g__4190(w__3163 ,in20[3] ,in21[5]);
  or g__4191(w__3162 ,w__3092 ,w__3126);
  or g__4192(w__3161 ,w__3129 ,w__3096);
  and g__4193(w__3159 ,in20[0] ,in21[5]);
  or g__4194(w__3158 ,w__3049 ,w__3068);
  or g__4195(w__3157 ,w__3107 ,w__3078);
  or g__4196(w__3156 ,w__3089 ,w__3034);
  or g__4197(w__3155 ,w__3114 ,w__3098);
  or g__4198(w__3154 ,w__3057 ,w__3105);
  or g__4199(w__3153 ,w__3074 ,w__3059);
  or g__4200(w__3152 ,w__3110 ,w__3101);
  or g__4201(w__3151 ,w__3089 ,w__3084);
  or g__4202(w__3150 ,w__3041 ,w__3068);
  or g__4203(w__3149 ,w__3080 ,w__3099);
  or g__4204(w__3148 ,w__3053 ,w__3102);
  or g__4205(w__3147 ,w__3055 ,w__3031);
  and g__4206(w__3145 ,in20[2] ,in21[6]);
  not g__4207(w__3140 ,in20[6]);
  not g__4208(w__3139 ,in20[2]);
  not g__4209(w__3138 ,in20[1]);
  not g__4210(w__3137 ,in20[4]);
  not g__4211(w__3136 ,in20[8]);
  not g__4212(w__3135 ,in21[3]);
  not g__4213(w__3134 ,in21[0]);
  not g__4214(w__3133 ,in21[1]);
  not g__4215(w__3132 ,in20[5]);
  not g__4216(w__3131 ,in20[3]);
  not g__4217(w__3130 ,in20[0]);
  not g__4218(w__3129 ,in20[7]);
  not g__4219(w__3128 ,in21[4]);
  not g__4220(w__3127 ,in21[2]);
  not g__4221(w__3126 ,in21[5]);
  not g__4222(w__3125 ,in21[7]);
  not g__4223(w__3124 ,in21[6]);
  not g__4224(w__3023 ,w__3122);
  not g__4225(w__3122 ,w__3130);
  not g__4226(w__3022 ,w__3121);
  not g__4227(w__3015 ,w__3121);
  not g__4228(w__3121 ,w__3133);
  not g__4229(w__3021 ,w__3120);
  not g__4230(w__3120 ,w__3134);
  buf g__4231(w__4193 ,w__3144);
  buf g__4232(w__4226 ,w__3141);
  buf g__4233(w__4195 ,w__3142);
  buf g__4234(w__4194 ,w__3143);
  buf g__4235(w__4192 ,w__3220);
  not g__4236(w__3119 ,w__3123);
  not g__4237(w__3123 ,w__3424);
  not g__4238(w__3118 ,w__3117);
  not g__4239(w__3117 ,w__3135);
  not g__4240(w__3116 ,w__3115);
  not g__4241(w__3115 ,w__3128);
  not g__4242(w__3114 ,w__3112);
  not g__4243(w__3113 ,w__3112);
  not g__4244(w__3112 ,w__3130);
  not g__4245(w__3111 ,w__3109);
  not g__4246(w__3110 ,w__3109);
  not g__4247(w__3109 ,w__3138);
  not g__4248(w__3108 ,w__3106);
  not g__4249(w__3107 ,w__3106);
  not g__4250(w__3106 ,w__3138);
  not g__4251(w__3105 ,w__3103);
  not g__4252(w__3104 ,w__3103);
  not g__4253(w__3103 ,w__3022);
  not g__4254(w__3102 ,w__3100);
  not g__4255(w__3101 ,w__3100);
  not g__4256(w__3100 ,w__3125);
  not g__4257(w__3099 ,w__3097);
  not g__4258(w__3098 ,w__3097);
  not g__4259(w__3097 ,w__3125);
  not g__4260(w__3096 ,w__3094);
  not g__4261(w__3095 ,w__3094);
  not g__4262(w__3094 ,w__3128);
  not g__4263(w__3093 ,w__3091);
  not g__4264(w__3092 ,w__3091);
  not g__4265(w__3091 ,w__3132);
  not g__4266(w__3090 ,w__3088);
  not g__4267(w__3089 ,w__3088);
  not g__4268(w__3088 ,w__3129);
  not g__4269(w__3087 ,w__3085);
  not g__4270(w__3086 ,w__3085);
  not g__4271(w__3085 ,w__3135);
  not g__4272(w__3084 ,w__3082);
  not g__4273(w__3083 ,w__3082);
  not g__4274(w__3082 ,w__3124);
  not g__4275(w__3081 ,w__3079);
  not g__4276(w__3080 ,w__3079);
  not g__4277(w__3079 ,w__3139);
  not g__4278(w__3078 ,w__3076);
  not g__4279(w__3077 ,w__3076);
  not g__4280(w__3076 ,w__3124);
  not g__4281(w__3075 ,w__3073);
  not g__4282(w__3074 ,w__3073);
  not g__4283(w__3073 ,w__3140);
  not g__4284(w__3072 ,w__3070);
  not g__4285(w__3071 ,w__3070);
  not g__4286(w__3070 ,w__3127);
  not g__4287(w__3069 ,w__3067);
  not g__4288(w__3068 ,w__3067);
  not g__4289(w__3067 ,w__3126);
  not g__4290(w__3066 ,w__3064);
  not g__4291(w__3065 ,w__3064);
  not g__4292(w__3064 ,w__3127);
  not g__4293(w__3020 ,w__3019);
  not g__4294(w__3063 ,w__3019);
  not g__4295(w__3019 ,w__3023);
  not g__4296(w__3018 ,w__3017);
  not g__4297(w__3062 ,w__3017);
  not g__4298(w__3017 ,w__3021);
  not g__4299(w__3016 ,w__3060);
  not g__4300(w__3061 ,w__3060);
  not g__4301(w__3060 ,w__3015);
  not g__4302(w__3059 ,w__3058);
  not g__4303(w__3058 ,w__3126);
  not g__4304(w__3057 ,w__3056);
  not g__4305(w__3056 ,w__3129);
  not g__4306(w__3055 ,w__3054);
  not g__4307(w__3054 ,w__3131);
  not g__4308(w__3053 ,w__3052);
  not g__4309(w__3052 ,w__3137);
  not g__4310(w__3051 ,w__3050);
  not g__4311(w__3050 ,w__3136);
  not g__4312(w__3049 ,w__3047);
  not g__4313(w__3048 ,w__3047);
  not g__4314(w__3047 ,w__3137);
  not g__4315(w__3046 ,w__3044);
  not g__4316(w__3045 ,w__3044);
  not g__4317(w__3044 ,w__3131);
  not g__4318(w__3043 ,w__3042);
  not g__4319(w__3042 ,w__3132);
  not g__4320(w__3041 ,w__3040);
  not g__4321(w__3040 ,w__3139);
  not g__4322(w__3039 ,w__3037);
  not g__4323(w__3038 ,w__3037);
  not g__4324(w__3037 ,w__3136);
  not g__4325(w__3036 ,w__3035);
  not g__4326(w__3035 ,w__3140);
  not g__4327(w__3034 ,w__3032);
  not g__4328(w__3033 ,w__3032);
  not g__4329(w__3032 ,w__3135);
  not g__4330(w__3031 ,w__3029);
  not g__4331(w__3030 ,w__3029);
  not g__4332(w__3029 ,w__3128);
  xnor g__4333(w__3028 ,w__3165 ,w__3176);
  xor g__4334(w__3027 ,w__3217 ,w__3174);
  xnor g__4335(w__3026 ,w__3173 ,w__3171);
  xor g__4336(w__3025 ,w__3209 ,w__3172);
  xor g__4337(w__3024 ,w__3206 ,w__3166);
  xnor g__4338(w__4152 ,w__3912 ,w__3929);
  or g__4339(w__4121 ,w__3928 ,w__3930);
  xnor g__4340(w__4151 ,w__3924 ,w__3925);
  nor g__4341(w__3930 ,w__3912 ,w__3927);
  or g__4342(w__4150 ,w__3920 ,w__3926);
  xnor g__4343(w__3929 ,w__3876 ,w__3918);
  xnor g__4344(w__4153 ,w__3903 ,w__3915);
  xnor g__4345(w__4154 ,w__3905 ,w__3914);
  xor g__4346(w__4120 ,w__3911 ,w__3913);
  or g__4347(w__4123 ,w__3909 ,w__3922);
  nor g__4348(w__3928 ,w__3876 ,w__3919);
  or g__4349(w__4149 ,w__3910 ,w__3921);
  and g__4350(w__3927 ,w__3876 ,w__3919);
  and g__4351(w__3926 ,w__3924 ,w__3916);
  or g__4352(w__4122 ,w__3898 ,w__3923);
  or g__4353(w__4124 ,w__3892 ,w__3917);
  xnor g__4354(w__4155 ,w__3904 ,w__3897);
  xnor g__4355(w__3925 ,w__3902 ,w__3878);
  and g__4356(w__3923 ,w__3908 ,w__3903);
  and g__4357(w__3922 ,w__3907 ,w__3905);
  or g__4358(w__4125 ,w__3857 ,w__3906);
  nor g__4359(w__3921 ,w__3900 ,w__3911);
  nor g__4360(w__3920 ,w__3878 ,w__3902);
  or g__4361(w__3924 ,w__3838 ,w__3899);
  not g__4362(w__3919 ,w__3918);
  nor g__4363(w__3917 ,w__3893 ,w__3904);
  or g__4364(w__3916 ,w__3877 ,w__3901);
  xnor g__4365(w__4156 ,w__3889 ,w__3864);
  xnor g__4366(w__3915 ,w__3885 ,w__3882);
  xnor g__4367(w__3914 ,w__3887 ,w__3896);
  xnor g__4368(w__3913 ,w__3883 ,w__3858);
  xnor g__4369(w__3918 ,w__3888 ,w__3862);
  nor g__4370(w__3910 ,w__3858 ,w__3883);
  nor g__4371(w__3909 ,w__3896 ,w__3887);
  or g__4372(w__3908 ,w__3581 ,w__3884);
  or g__4373(w__3907 ,w__3895 ,w__3886);
  or g__4374(w__4148 ,w__3842 ,w__3881);
  nor g__4375(w__3906 ,w__3848 ,w__3889);
  or g__4376(w__4126 ,w__3847 ,w__3890);
  and g__4377(w__3912 ,w__3849 ,w__3891);
  and g__4378(w__3911 ,w__3874 ,w__3894);
  not g__4379(w__3901 ,w__3902);
  and g__4380(w__3900 ,w__3858 ,w__3883);
  and g__4381(w__3899 ,w__3837 ,w__3888);
  nor g__4382(w__3898 ,w__3577 ,w__3885);
  xor g__4383(w__4119 ,w__3879 ,w__3860);
  xnor g__4384(w__4157 ,w__3870 ,w__3866);
  xnor g__4385(w__3897 ,w__3875 ,w__3868);
  xnor g__4386(w__3905 ,w__3859 ,w__3867);
  xnor g__4387(w__3904 ,w__3787 ,w__3861);
  xnor g__4388(w__3903 ,w__3880 ,w__3863);
  xnor g__4389(w__3902 ,w__3844 ,w__3865);
  not g__4390(w__3896 ,w__3895);
  or g__4391(w__3894 ,w__3788 ,w__3871);
  and g__4392(w__3893 ,w__3875 ,w__3869);
  nor g__4393(w__3892 ,w__3875 ,w__3869);
  or g__4394(w__3891 ,w__3845 ,w__3880);
  and g__4395(w__3890 ,w__3846 ,w__3870);
  or g__4396(w__3895 ,w__3853 ,w__3872);
  not g__4397(w__3886 ,w__3887);
  not g__4398(w__3884 ,w__3885);
  nor g__4399(w__3881 ,w__3841 ,w__3879);
  xnor g__4400(w__3889 ,w__3813 ,w__3835);
  xnor g__4401(w__3888 ,w__3809 ,w__3834);
  xnor g__4402(w__3887 ,w__3810 ,w__3836);
  and g__4403(w__3885 ,w__3843 ,w__3873);
  xnor g__4404(w__3883 ,w__3808 ,w__3833);
  xnor g__4405(w__3882 ,w__3811 ,w__3832);
  not g__4406(w__3877 ,w__3878);
  or g__4407(w__3874 ,w__3797 ,w__3844);
  or g__4408(w__3873 ,w__3859 ,w__3855);
  nor g__4409(w__3872 ,w__3787 ,w__3852);
  and g__4410(w__3871 ,w__3797 ,w__3844);
  or g__4411(w__4127 ,w__3768 ,w__3850);
  and g__4412(w__3880 ,w__3820 ,w__3840);
  and g__4413(w__3879 ,w__3818 ,w__3856);
  and g__4414(w__3878 ,w__3816 ,w__3839);
  and g__4415(w__3876 ,w__3827 ,w__3854);
  and g__4416(w__3875 ,w__3824 ,w__3851);
  not g__4417(w__3869 ,w__3868);
  xnor g__4418(w__4158 ,w__3812 ,w__3814);
  xnor g__4419(w__3867 ,w__3796 ,w__3793);
  xnor g__4420(w__3866 ,w__3803 ,w__3774);
  xnor g__4421(w__3865 ,w__3797 ,w__3788);
  xnor g__4422(w__3864 ,w__3829 ,w__3806);
  xnor g__4423(w__3863 ,w__3776 ,w__3801);
  xnor g__4424(w__3862 ,w__3805 ,w__3831);
  xnor g__4425(w__3861 ,w__3799 ,w__3798);
  xnor g__4426(w__3860 ,w__3794 ,w__3771);
  xnor g__4427(w__3870 ,w__3724 ,w__3791);
  xnor g__4428(w__3868 ,w__3789 ,w__3815);
  nor g__4429(w__3857 ,w__3829 ,w__3807);
  or g__4430(w__3856 ,w__3822 ,w__3808);
  nor g__4431(w__3855 ,w__3795 ,w__3793);
  or g__4432(w__3854 ,w__3811 ,w__3826);
  nor g__4433(w__3853 ,w__3798 ,w__3799);
  and g__4434(w__3852 ,w__3798 ,w__3799);
  or g__4435(w__3851 ,w__3823 ,w__3813);
  nor g__4436(w__3850 ,w__3779 ,w__3812);
  or g__4437(w__3849 ,w__3775 ,w__3801);
  and g__4438(w__3848 ,w__3829 ,w__3807);
  nor g__4439(w__3847 ,w__3774 ,w__3803);
  or g__4440(w__3846 ,w__3773 ,w__3802);
  nor g__4441(w__3845 ,w__3776 ,w__3800);
  and g__4442(w__3859 ,w__3767 ,w__3819);
  and g__4443(w__3858 ,w__3720 ,w__3828);
  or g__4444(w__3843 ,w__3796 ,w__3792);
  nor g__4445(w__3842 ,w__3771 ,w__3794);
  and g__4446(w__3841 ,w__3771 ,w__3794);
  or g__4447(w__3840 ,w__3810 ,w__3825);
  or g__4448(w__3839 ,w__3821 ,w__3809);
  nor g__4449(w__3838 ,w__3831 ,w__3805);
  or g__4450(w__3837 ,w__3830 ,w__3804);
  or g__4451(w__4147 ,w__3684 ,w__3817);
  xor g__4452(w__4118 ,w__3778 ,w__3738);
  xnor g__4453(w__3836 ,w__3777 ,w__3769);
  xnor g__4454(w__3835 ,w__3784 ,w__3482);
  xnor g__4455(w__3834 ,w__3700 ,w__3786);
  xnor g__4456(w__3833 ,w__3639 ,w__3772);
  xnor g__4457(w__3832 ,w__3783 ,w__3770);
  xnor g__4458(w__3844 ,w__3790 ,w__3739);
  not g__4459(w__3830 ,w__3831);
  or g__4460(w__3828 ,w__3682 ,w__3790);
  or g__4461(w__3827 ,w__3770 ,w__3783);
  and g__4462(w__3826 ,w__3770 ,w__3783);
  and g__4463(w__3825 ,w__3769 ,w__3777);
  or g__4464(w__3824 ,w__3482 ,w__3784);
  and g__4465(w__3823 ,w__3482 ,w__3784);
  and g__4466(w__3822 ,w__3639 ,w__3772);
  nor g__4467(w__3821 ,w__3700 ,w__3785);
  or g__4468(w__3820 ,w__3769 ,w__3777);
  or g__4469(w__3819 ,w__3789 ,w__3780);
  or g__4470(w__4128 ,w__3683 ,w__3766);
  or g__4471(w__3818 ,w__3639 ,w__3772);
  nor g__4472(w__3817 ,w__3698 ,w__3778);
  or g__4473(w__3816 ,w__3699 ,w__3786);
  xnor g__4474(w__3815 ,w__3722 ,w__3765);
  xnor g__4475(w__3814 ,w__3701 ,w__3483);
  and g__4476(w__3831 ,w__3705 ,w__3781);
  and g__4477(w__3829 ,w__3756 ,w__3782);
  not g__4478(w__3807 ,w__3806);
  not g__4479(w__3804 ,w__3805);
  not g__4480(w__3802 ,w__3803);
  not g__4481(w__3800 ,w__3801);
  not g__4482(w__3795 ,w__3796);
  not g__4483(w__3792 ,w__3793);
  xor g__4484(w__4159 ,w__3485 ,w__3745);
  xnor g__4485(w__3791 ,w__3618 ,w__3486);
  xnor g__4486(w__3813 ,w__3663 ,w__3746);
  xnor g__4487(w__3812 ,w__3669 ,w__3728);
  xnor g__4488(w__3811 ,w__3671 ,w__3742);
  xnor g__4489(w__3810 ,w__3652 ,w__3737);
  xnor g__4490(w__3809 ,w__3645 ,w__3735);
  xnor g__4491(w__3808 ,w__3642 ,w__3734);
  xnor g__4492(w__3806 ,w__3725 ,w__3731);
  xnor g__4493(w__3805 ,w__3620 ,w__3744);
  xnor g__4494(w__3803 ,w__3625 ,w__3730);
  xnor g__4495(w__3801 ,w__3484 ,w__3729);
  xnor g__4496(w__3799 ,w__3615 ,w__3740);
  xnor g__4497(w__3798 ,w__3605 ,w__3741);
  xnor g__4498(w__3797 ,w__3640 ,w__3743);
  xnor g__4499(w__3796 ,w__3670 ,w__3736);
  xnor g__4500(w__3794 ,w__3644 ,w__3732);
  xnor g__4501(w__3793 ,w__3727 ,w__3733);
  not g__4502(w__3785 ,w__3786);
  or g__4503(w__3782 ,w__3763 ,w__3486);
  or g__4504(w__3781 ,w__3712 ,w__3484);
  nor g__4505(w__3780 ,w__3722 ,w__3764);
  and g__4506(w__3779 ,w__3702 ,w__3483);
  and g__4507(w__3790 ,w__3710 ,w__3762);
  and g__4508(w__3789 ,w__3717 ,w__3754);
  and g__4509(w__3788 ,w__3711 ,w__3752);
  and g__4510(w__3787 ,w__3697 ,w__3760);
  and g__4511(w__3786 ,w__3692 ,w__3755);
  and g__4512(w__3784 ,w__3694 ,w__3758);
  and g__4513(w__3783 ,w__3715 ,w__3747);
  not g__4514(w__3775 ,w__3776);
  not g__4515(w__3773 ,w__3774);
  nor g__4516(w__3768 ,w__3702 ,w__3483);
  or g__4517(w__3767 ,w__3721 ,w__3765);
  nor g__4518(w__3766 ,w__3708 ,w__3485);
  and g__4519(w__3778 ,w__3685 ,w__3759);
  and g__4520(w__3777 ,w__3680 ,w__3753);
  or g__4521(w__3776 ,w__3704 ,w__3751);
  and g__4522(w__3774 ,w__3690 ,w__3750);
  and g__4523(w__3772 ,w__3689 ,w__3761);
  and g__4524(w__3771 ,w__3681 ,w__3748);
  and g__4525(w__3770 ,w__3706 ,w__3757);
  and g__4526(w__3769 ,w__3713 ,w__3749);
  not g__4527(w__3764 ,w__3765);
  nor g__4528(w__3763 ,w__3617 ,w__3724);
  or g__4529(w__3762 ,w__3636 ,w__3695);
  or g__4530(w__3761 ,w__3635 ,w__3707);
  or g__4531(w__3760 ,w__3718 ,w__3726);
  or g__4532(w__3759 ,w__3628 ,w__3691);
  or g__4533(w__3758 ,w__3625 ,w__3696);
  or g__4534(w__3757 ,w__3670 ,w__3693);
  or g__4535(w__3756 ,w__3618 ,w__3723);
  or g__4536(w__3755 ,w__3671 ,w__3719);
  or g__4537(w__3754 ,w__3663 ,w__3714);
  or g__4538(w__3753 ,w__3633 ,w__3703);
  or g__4539(w__3752 ,w__3626 ,w__3687);
  and g__4540(w__3751 ,w__3709 ,w__3727);
  or g__4541(w__3750 ,w__3669 ,w__3686);
  or g__4542(w__3749 ,w__3672 ,w__3688);
  or g__4543(w__3748 ,w__3627 ,w__3679);
  xor g__4544(w__4160 ,w__3637 ,w__3677);
  or g__4545(w__3747 ,w__3666 ,w__3716);
  xnor g__4546(w__3746 ,w__3656 ,w__3659);
  xnor g__4547(w__3745 ,w__3641 ,w__3653);
  xnor g__4548(w__3765 ,w__3673 ,w__3661);
  xnor g__4549(w__3744 ,w__3614 ,w__3626);
  xnor g__4550(w__3743 ,w__3619 ,w__3635);
  xnor g__4551(w__3742 ,w__3616 ,w__3647);
  xnor g__4552(w__3741 ,w__3613 ,w__3633);
  xnor g__4553(w__3740 ,w__3608 ,w__3672);
  xnor g__4554(w__3739 ,w__3606 ,w__3611);
  xnor g__4555(w__3738 ,w__3660 ,w__3654);
  xnor g__4556(w__3737 ,w__3612 ,w__3666);
  xnor g__4557(w__3736 ,w__3610 ,w__3648);
  xnor g__4558(w__3735 ,w__3658 ,w__3636);
  xnor g__4559(w__3734 ,w__3657 ,w__3627);
  xnor g__4560(w__3733 ,w__3604 ,w__3622);
  xnor g__4561(w__3732 ,w__3609 ,w__3628);
  xnor g__4562(w__3731 ,w__3638 ,w__3646);
  xnor g__4563(w__3730 ,w__3643 ,w__3651);
  xnor g__4564(w__3729 ,w__3607 ,w__3650);
  xnor g__4565(w__3728 ,w__3655 ,w__3649);
  not g__4566(w__3726 ,w__3725);
  not g__4567(w__3723 ,w__3724);
  not g__4568(w__3721 ,w__3722);
  or g__4569(w__3720 ,w__3606 ,w__3611);
  and g__4570(w__3719 ,w__3616 ,w__3647);
  and g__4571(w__3718 ,w__3638 ,w__3646);
  or g__4572(w__3717 ,w__3656 ,w__3659);
  and g__4573(w__3716 ,w__3652 ,w__3612);
  or g__4574(w__3715 ,w__3652 ,w__3612);
  and g__4575(w__3714 ,w__3656 ,w__3659);
  or g__4576(w__3713 ,w__3615 ,w__3608);
  and g__4577(w__3712 ,w__3607 ,w__3650);
  or g__4578(w__3711 ,w__3620 ,w__3614);
  or g__4579(w__3710 ,w__3645 ,w__3658);
  or g__4580(w__3709 ,w__3603 ,w__3621);
  and g__4581(w__3708 ,w__3641 ,w__3653);
  and g__4582(w__3707 ,w__3640 ,w__3619);
  or g__4583(w__3706 ,w__3610 ,w__3648);
  or g__4584(w__3705 ,w__3607 ,w__3650);
  nor g__4585(w__3704 ,w__3604 ,w__3622);
  and g__4586(w__3703 ,w__3613 ,w__3605);
  and g__4587(w__3727 ,w__3674 ,w__3662);
  and g__4588(w__3725 ,w__3623 ,w__3634);
  and g__4589(w__3724 ,w__3668 ,w__3630);
  and g__4590(w__3722 ,w__3665 ,w__3624);
  not g__4591(w__3702 ,w__3701);
  not g__4592(w__3699 ,w__3700);
  and g__4593(w__3698 ,w__3660 ,w__3654);
  or g__4594(w__3697 ,w__3638 ,w__3646);
  and g__4595(w__3696 ,w__3643 ,w__3651);
  and g__4596(w__3695 ,w__3645 ,w__3658);
  or g__4597(w__3694 ,w__3643 ,w__3651);
  and g__4598(w__3693 ,w__3610 ,w__3648);
  or g__4599(w__3692 ,w__3616 ,w__3647);
  and g__4600(w__3691 ,w__3644 ,w__3609);
  or g__4601(w__3690 ,w__3655 ,w__3649);
  or g__4602(w__3689 ,w__3640 ,w__3619);
  and g__4603(w__3688 ,w__3615 ,w__3608);
  and g__4604(w__3687 ,w__3620 ,w__3614);
  and g__4605(w__3686 ,w__3655 ,w__3649);
  or g__4606(w__3685 ,w__3644 ,w__3609);
  nor g__4607(w__3684 ,w__3660 ,w__3654);
  nor g__4608(w__3683 ,w__3641 ,w__3653);
  and g__4609(w__3682 ,w__3606 ,w__3611);
  or g__4610(w__3681 ,w__3642 ,w__3657);
  or g__4611(w__3680 ,w__3613 ,w__3605);
  and g__4612(w__3679 ,w__3642 ,w__3657);
  nor g__4613(w__3678 ,w__3677 ,w__3637);
  and g__4614(w__3701 ,w__3676 ,w__3632);
  and g__4615(w__3700 ,w__3631 ,w__3629);
  not g__4616(w__3676 ,w__3675);
  not g__4617(w__3674 ,w__3673);
  not g__4618(w__3668 ,w__3667);
  not g__4619(w__3665 ,w__3664);
  not g__4620(w__3662 ,w__3661);
  and g__4621(w__4117 ,in24[8] ,in25[7]);
  or g__4622(w__3677 ,w__3499 ,w__3592);
  or g__4623(w__3675 ,w__3539 ,w__3519);
  or g__4624(w__3673 ,w__3494 ,w__3562);
  or g__4625(w__3672 ,w__3501 ,w__3529);
  or g__4626(w__3671 ,w__3533 ,w__3544);
  or g__4627(w__3670 ,w__3533 ,w__3523);
  or g__4628(w__3669 ,w__3539 ,w__3524);
  or g__4629(w__3667 ,w__3513 ,w__3562);
  or g__4630(w__3666 ,w__3509 ,w__3520);
  or g__4631(w__3664 ,w__3551 ,w__3519);
  or g__4632(w__3663 ,w__3511 ,w__3530);
  or g__4633(w__3661 ,w__3515 ,w__3520);
  or g__4634(w__3660 ,w__3548 ,w__3559);
  or g__4635(w__3659 ,w__3504 ,w__3491);
  or g__4636(w__3658 ,w__3507 ,w__3541);
  or g__4637(w__3657 ,w__3548 ,w__3517);
  or g__4638(w__3656 ,w__3597 ,w__3553);
  or g__4639(w__3655 ,w__3521 ,w__3488);
  or g__4640(w__3654 ,w__3497 ,w__3535);
  or g__4641(w__3653 ,w__3569 ,w__3523);
  or g__4642(w__3652 ,w__3551 ,w__3576);
  or g__4643(w__3651 ,w__3538 ,w__3545);
  or g__4644(w__3650 ,w__3503 ,w__3536);
  or g__4645(w__3649 ,w__3566 ,w__3492);
  or g__4646(w__3648 ,w__3506 ,w__3574);
  or g__4647(w__3647 ,w__3590 ,w__3554);
  or g__4648(w__3646 ,w__3565 ,w__3527);
  or g__4649(w__3645 ,w__3589 ,w__3556);
  or g__4650(w__3644 ,w__3598 ,w__3557);
  or g__4651(w__3643 ,w__3568 ,w__3489);
  or g__4652(w__3642 ,w__3550 ,w__3560);
  or g__4653(w__3641 ,w__3571 ,w__3544);
  or g__4654(w__3640 ,w__3501 ,w__3542);
  or g__4655(w__3639 ,w__3532 ,w__3535);
  or g__4656(w__3638 ,w__3571 ,w__3541);
  not g__4657(w__3622 ,w__3621);
  not g__4658(w__3618 ,w__3617);
  not g__4659(w__3604 ,w__3603);
  nor g__4660(w__3602 ,w__3566 ,w__3474);
  nor g__4661(w__3601 ,w__3569 ,w__3476);
  nor g__4662(w__3600 ,w__3592 ,w__3478);
  nor g__4663(w__3599 ,w__3572 ,w__3563);
  or g__4664(w__3637 ,w__3521 ,w__3529);
  or g__4665(w__3636 ,w__3494 ,w__3553);
  or g__4666(w__3635 ,w__3496 ,w__3576);
  and g__4667(w__3634 ,in24[5] ,in25[0]);
  or g__4668(w__3633 ,w__3595 ,w__3545);
  and g__4669(w__3632 ,in24[3] ,in25[0]);
  and g__4670(w__3631 ,in24[7] ,in25[2]);
  and g__4671(w__3630 ,in24[4] ,in25[0]);
  and g__4672(w__3629 ,in24[8] ,in25[1]);
  or g__4673(w__3628 ,w__3594 ,w__3527);
  or g__4674(w__3627 ,w__3497 ,w__3574);
  or g__4675(w__3626 ,w__3509 ,w__3524);
  or g__4676(w__3625 ,w__3504 ,w__3530);
  and g__4677(w__3624 ,in24[6] ,in25[0]);
  and g__4678(w__3623 ,in24[4] ,in25[1]);
  and g__4679(w__3621 ,in24[3] ,in25[5]);
  or g__4680(w__3620 ,w__3550 ,w__3584);
  or g__4681(w__3619 ,w__3587 ,w__3554);
  and g__4682(w__3617 ,in24[0] ,in25[5]);
  or g__4683(w__3616 ,w__3507 ,w__3526);
  or g__4684(w__3615 ,w__3565 ,w__3536);
  or g__4685(w__3614 ,w__3547 ,w__3492);
  or g__4686(w__3613 ,w__3572 ,w__3556);
  or g__4687(w__3612 ,w__3515 ,w__3563);
  or g__4688(w__3611 ,w__3532 ,w__3517);
  or g__4689(w__3610 ,w__3568 ,w__3559);
  or g__4690(w__3609 ,w__3547 ,w__3542);
  or g__4691(w__3608 ,w__3499 ,w__3526);
  or g__4692(w__3607 ,w__3538 ,w__3557);
  or g__4693(w__3606 ,w__3511 ,w__3560);
  or g__4694(w__3605 ,w__3513 ,w__3489);
  and g__4695(w__3603 ,in24[2] ,in25[6]);
  not g__4696(w__3598 ,in24[6]);
  not g__4697(w__3597 ,in24[2]);
  not g__4698(w__3596 ,in24[1]);
  not g__4699(w__3595 ,in24[4]);
  not g__4700(w__3594 ,in24[8]);
  not g__4701(w__3593 ,in25[3]);
  not g__4702(w__3592 ,in25[0]);
  not g__4703(w__3591 ,in25[1]);
  not g__4704(w__3590 ,in24[5]);
  not g__4705(w__3589 ,in24[3]);
  not g__4706(w__3588 ,in24[0]);
  not g__4707(w__3587 ,in24[7]);
  not g__4708(w__3586 ,in25[4]);
  not g__4709(w__3585 ,in25[2]);
  not g__4710(w__3584 ,in25[5]);
  not g__4711(w__3583 ,in25[7]);
  not g__4712(w__3582 ,in25[6]);
  not g__4713(w__3481 ,w__3580);
  not g__4714(w__3580 ,w__3588);
  not g__4715(w__3480 ,w__3579);
  not g__4716(w__3473 ,w__3579);
  not g__4717(w__3579 ,w__3591);
  not g__4718(w__3479 ,w__3578);
  not g__4719(w__3578 ,w__3592);
  buf g__4720(w__4130 ,w__3602);
  buf g__4721(w__4161 ,w__3599);
  buf g__4722(w__4132 ,w__3600);
  buf g__4723(w__4131 ,w__3601);
  buf g__4724(w__4129 ,w__3678);
  not g__4725(w__3577 ,w__3581);
  not g__4726(w__3581 ,w__3882);
  not g__4727(w__3576 ,w__3575);
  not g__4728(w__3575 ,w__3593);
  not g__4729(w__3574 ,w__3573);
  not g__4730(w__3573 ,w__3586);
  not g__4731(w__3572 ,w__3570);
  not g__4732(w__3571 ,w__3570);
  not g__4733(w__3570 ,w__3588);
  not g__4734(w__3569 ,w__3567);
  not g__4735(w__3568 ,w__3567);
  not g__4736(w__3567 ,w__3596);
  not g__4737(w__3566 ,w__3564);
  not g__4738(w__3565 ,w__3564);
  not g__4739(w__3564 ,w__3596);
  not g__4740(w__3563 ,w__3561);
  not g__4741(w__3562 ,w__3561);
  not g__4742(w__3561 ,w__3480);
  not g__4743(w__3560 ,w__3558);
  not g__4744(w__3559 ,w__3558);
  not g__4745(w__3558 ,w__3583);
  not g__4746(w__3557 ,w__3555);
  not g__4747(w__3556 ,w__3555);
  not g__4748(w__3555 ,w__3583);
  not g__4749(w__3554 ,w__3552);
  not g__4750(w__3553 ,w__3552);
  not g__4751(w__3552 ,w__3586);
  not g__4752(w__3551 ,w__3549);
  not g__4753(w__3550 ,w__3549);
  not g__4754(w__3549 ,w__3590);
  not g__4755(w__3548 ,w__3546);
  not g__4756(w__3547 ,w__3546);
  not g__4757(w__3546 ,w__3587);
  not g__4758(w__3545 ,w__3543);
  not g__4759(w__3544 ,w__3543);
  not g__4760(w__3543 ,w__3593);
  not g__4761(w__3542 ,w__3540);
  not g__4762(w__3541 ,w__3540);
  not g__4763(w__3540 ,w__3582);
  not g__4764(w__3539 ,w__3537);
  not g__4765(w__3538 ,w__3537);
  not g__4766(w__3537 ,w__3597);
  not g__4767(w__3536 ,w__3534);
  not g__4768(w__3535 ,w__3534);
  not g__4769(w__3534 ,w__3582);
  not g__4770(w__3533 ,w__3531);
  not g__4771(w__3532 ,w__3531);
  not g__4772(w__3531 ,w__3598);
  not g__4773(w__3530 ,w__3528);
  not g__4774(w__3529 ,w__3528);
  not g__4775(w__3528 ,w__3585);
  not g__4776(w__3527 ,w__3525);
  not g__4777(w__3526 ,w__3525);
  not g__4778(w__3525 ,w__3584);
  not g__4779(w__3524 ,w__3522);
  not g__4780(w__3523 ,w__3522);
  not g__4781(w__3522 ,w__3585);
  not g__4782(w__3478 ,w__3477);
  not g__4783(w__3521 ,w__3477);
  not g__4784(w__3477 ,w__3481);
  not g__4785(w__3476 ,w__3475);
  not g__4786(w__3520 ,w__3475);
  not g__4787(w__3475 ,w__3479);
  not g__4788(w__3474 ,w__3518);
  not g__4789(w__3519 ,w__3518);
  not g__4790(w__3518 ,w__3473);
  not g__4791(w__3517 ,w__3516);
  not g__4792(w__3516 ,w__3584);
  not g__4793(w__3515 ,w__3514);
  not g__4794(w__3514 ,w__3587);
  not g__4795(w__3513 ,w__3512);
  not g__4796(w__3512 ,w__3589);
  not g__4797(w__3511 ,w__3510);
  not g__4798(w__3510 ,w__3595);
  not g__4799(w__3509 ,w__3508);
  not g__4800(w__3508 ,w__3594);
  not g__4801(w__3507 ,w__3505);
  not g__4802(w__3506 ,w__3505);
  not g__4803(w__3505 ,w__3595);
  not g__4804(w__3504 ,w__3502);
  not g__4805(w__3503 ,w__3502);
  not g__4806(w__3502 ,w__3589);
  not g__4807(w__3501 ,w__3500);
  not g__4808(w__3500 ,w__3590);
  not g__4809(w__3499 ,w__3498);
  not g__4810(w__3498 ,w__3597);
  not g__4811(w__3497 ,w__3495);
  not g__4812(w__3496 ,w__3495);
  not g__4813(w__3495 ,w__3594);
  not g__4814(w__3494 ,w__3493);
  not g__4815(w__3493 ,w__3598);
  not g__4816(w__3492 ,w__3490);
  not g__4817(w__3491 ,w__3490);
  not g__4818(w__3490 ,w__3593);
  not g__4819(w__3489 ,w__3487);
  not g__4820(w__3488 ,w__3487);
  not g__4821(w__3487 ,w__3586);
  xnor g__4822(w__3486 ,w__3623 ,w__3634);
  xor g__4823(w__3485 ,w__3675 ,w__3632);
  xnor g__4824(w__3484 ,w__3631 ,w__3629);
  xor g__4825(w__3483 ,w__3667 ,w__3630);
  xor g__4826(w__3482 ,w__3664 ,w__3624);
  buf g__4827(w__426 ,in5[0]);
  not g__4828(w__611 ,w__59);
  not g__4829(w__230 ,w__3977);
  buf g__4830(w__338 ,w__131);
  buf g__4831(w__675 ,w__4086);
  not g__4832(w__759 ,w__614);
  buf g__4833(w__716 ,w__562);
  not g__4834(w__739 ,w__610);
  buf g__4835(w__792 ,w__574);
  not g__4836(w__849 ,w__509);
endmodule
