module top( 1_n1 , 1_n4 , 1_n10 , 1_n13 , 1_n26 , 1_n27 , 1_n32 , 1_n34 , 1_n46 , 1_n52 , 1_n54 , 1_n58 , 1_n61 , 1_n64 , 1_n65 , 1_n66 );
    input 1_n1 , 1_n4 , 1_n10 , 1_n13 , 1_n27 , 1_n32 , 1_n46 , 1_n58 , 1_n61 , 1_n64 , 1_n65 , 1_n66 ;
    output 1_n26 , 1_n34 , 1_n52 , 1_n54 ;
    wire 1_n0 , 1_n2 , 1_n3 , 1_n5 , 1_n6 , 1_n7 , 1_n8 , 1_n9 , 1_n11 , 1_n12 , 1_n14 , 1_n15 , 1_n16 , 1_n17 , 1_n18 , 1_n19 , 1_n20 , 1_n21 , 1_n22 , 1_n23 , 1_n24 , 1_n25 , 1_n28 , 1_n29 , 1_n30 , 1_n31 , 1_n33 , 1_n35 , 1_n36 , 1_n37 , 1_n38 , 1_n39 , 1_n40 , 1_n41 , 1_n42 , 1_n43 , 1_n44 , 1_n45 , 1_n47 , 1_n48 , 1_n49 , 1_n50 , 1_n51 , 1_n53 , 1_n55 , 1_n56 , 1_n57 , 1_n59 , 1_n60 , 1_n62 , 1_n63 , 1_n67 , 1_n68 , 1_n69 , 1_n70 ;
assign 1_n33 = ~1_n46;
assign 1_n17 = 1_n8 & 1_n40;
assign 1_n23 = ~(1_n14 ^ 1_n64);
assign 1_n47 = ~(1_n17 | 1_n49);
assign 1_n29 = 1_n61 | 1_n33;
assign 1_n69 = ~(1_n19 | 1_n36);
assign 1_n34 = ~(1_n49 ^ 1_n0);
assign 1_n18 = ~(1_n40 | 1_n8);
assign 1_n7 = ~1_n58;
assign 1_n16 = ~(1_n20 ^ 1_n1);
assign 1_n37 = ~1_n70;
assign 1_n8 = ~(1_n70 ^ 1_n44);
assign 1_n53 = ~1_n24;
assign 1_n40 = ~1_n27;
assign 1_n14 = ~(1_n18 | 1_n47);
assign 1_n24 = 1_n41 & 1_n2;
assign 1_n12 = ~(1_n48 | 1_n69);
assign 1_n35 = ~(1_n29 ^ 1_n63);
assign 1_n60 = ~1_n55;
assign 1_n63 = 1_n66 | 1_n7;
assign 1_n55 = 1_n67 & 1_n11;
assign 1_n68 = 1_n11 | 1_n67;
assign 1_n22 = 1_n1 | 1_n60;
assign 1_n25 = ~(1_n57 | 1_n12);
assign 1_n19 = ~1_n53;
assign 1_n51 = ~(1_n13 | 1_n66);
assign 1_n39 = ~(1_n25 ^ 1_n50);
assign 1_n41 = ~1_n13;
assign 1_n50 = ~(1_n70 | 1_n44);
assign 1_n43 = ~(1_n39 ^ 1_n23);
assign 1_n38 = ~(1_n24 ^ 1_n48);
assign 1_n20 = 1_n9 | 1_n37;
assign 1_n70 = 1_n53 | 1_n28;
assign 1_n28 = ~1_n67;
assign 1_n11 = ~1_n4;
assign 1_n31 = ~1_n55;
assign 1_n44 = ~(1_n36 ^ 1_n38);
assign 1_n9 = ~(1_n56 | 1_n51);
assign 1_n15 = 1_n42 | 1_n20;
assign 1_n67 = 1_n62 & 1_n3;
assign 1_n21 = 1_n13 | 1_n30;
assign 1_n49 = 1_n15 & 1_n22;
assign 1_n30 = ~1_n10;
assign 1_n48 = 1_n66 | 1_n5;
assign 1_n52 = ~(1_n59 ^ 1_n43);
assign 1_n0 = ~(1_n8 ^ 1_n27);
assign 1_n45 = ~(1_n6 ^ 1_n21);
assign 1_n54 = 1_n60 & 1_n68;
assign 1_n57 = 1_n36 & 1_n19;
assign 1_n5 = ~1_n65;
assign 1_n62 = ~1_n61;
assign 1_n3 = ~1_n66;
assign 1_n2 = ~1_n32;
assign 1_n56 = ~(1_n61 | 1_n32);
assign 1_n59 = ~(1_n35 ^ 1_n45);
assign 1_n26 = ~(1_n55 ^ 1_n16);
assign 1_n36 = 1_n62 & 1_n10;
assign 1_n42 = 1_n31 & 1_n1;
assign 1_n6 = ~(1_n32 | 1_n5);
endmodule
