interface iface;
endinterface

module a (
  iface x = 1'b0
);
endmodule
