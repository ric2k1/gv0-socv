module top(in1, in2, in3, out2);
  input [31:0] in1, in2, in3;
  output [40:0] out2;
  wire [31:0] in1, in2, in3;
  wire [40:0] out2;
  wire csa_tree_add_7_25_groupi_n_0, csa_tree_add_7_25_groupi_n_1, csa_tree_add_7_25_groupi_n_2, csa_tree_add_7_25_groupi_n_7, csa_tree_add_7_25_groupi_n_8, csa_tree_add_7_25_groupi_n_9, csa_tree_add_7_25_groupi_n_10, csa_tree_add_7_25_groupi_n_11;
  wire csa_tree_add_7_25_groupi_n_12, csa_tree_add_7_25_groupi_n_13, csa_tree_add_7_25_groupi_n_14, csa_tree_add_7_25_groupi_n_15, csa_tree_add_7_25_groupi_n_16, csa_tree_add_7_25_groupi_n_17, csa_tree_add_7_25_groupi_n_18, csa_tree_add_7_25_groupi_n_19;
  wire csa_tree_add_7_25_groupi_n_20, csa_tree_add_7_25_groupi_n_21, csa_tree_add_7_25_groupi_n_22, csa_tree_add_7_25_groupi_n_23, csa_tree_add_7_25_groupi_n_24, csa_tree_add_7_25_groupi_n_25, csa_tree_add_7_25_groupi_n_26, csa_tree_add_7_25_groupi_n_27;
  wire csa_tree_add_7_25_groupi_n_28, csa_tree_add_7_25_groupi_n_29, csa_tree_add_7_25_groupi_n_30, csa_tree_add_7_25_groupi_n_31, csa_tree_add_7_25_groupi_n_32, csa_tree_add_7_25_groupi_n_33, csa_tree_add_7_25_groupi_n_34, csa_tree_add_7_25_groupi_n_35;
  wire csa_tree_add_7_25_groupi_n_36, csa_tree_add_7_25_groupi_n_37, csa_tree_add_7_25_groupi_n_38, csa_tree_add_7_25_groupi_n_39, csa_tree_add_7_25_groupi_n_40, csa_tree_add_7_25_groupi_n_41, csa_tree_add_7_25_groupi_n_42, csa_tree_add_7_25_groupi_n_43;
  wire csa_tree_add_7_25_groupi_n_44, csa_tree_add_7_25_groupi_n_45, csa_tree_add_7_25_groupi_n_46, csa_tree_add_7_25_groupi_n_47, csa_tree_add_7_25_groupi_n_48, csa_tree_add_7_25_groupi_n_49, csa_tree_add_7_25_groupi_n_50, csa_tree_add_7_25_groupi_n_51;
  wire csa_tree_add_7_25_groupi_n_52, csa_tree_add_7_25_groupi_n_53, csa_tree_add_7_25_groupi_n_54, csa_tree_add_7_25_groupi_n_55, csa_tree_add_7_25_groupi_n_56, csa_tree_add_7_25_groupi_n_57, csa_tree_add_7_25_groupi_n_58, csa_tree_add_7_25_groupi_n_59;
  wire csa_tree_add_7_25_groupi_n_60, csa_tree_add_7_25_groupi_n_61, csa_tree_add_7_25_groupi_n_62, csa_tree_add_7_25_groupi_n_63, csa_tree_add_7_25_groupi_n_64, csa_tree_add_7_25_groupi_n_65, csa_tree_add_7_25_groupi_n_66, csa_tree_add_7_25_groupi_n_67;
  wire csa_tree_add_7_25_groupi_n_68, csa_tree_add_7_25_groupi_n_69, csa_tree_add_7_25_groupi_n_70, csa_tree_add_7_25_groupi_n_71, csa_tree_add_7_25_groupi_n_72, csa_tree_add_7_25_groupi_n_73, csa_tree_add_7_25_groupi_n_74, csa_tree_add_7_25_groupi_n_75;
  wire csa_tree_add_7_25_groupi_n_76, csa_tree_add_7_25_groupi_n_77, csa_tree_add_7_25_groupi_n_78, csa_tree_add_7_25_groupi_n_79, csa_tree_add_7_25_groupi_n_80, csa_tree_add_7_25_groupi_n_81, csa_tree_add_7_25_groupi_n_82, csa_tree_add_7_25_groupi_n_83;
  wire csa_tree_add_7_25_groupi_n_84, csa_tree_add_7_25_groupi_n_85, csa_tree_add_7_25_groupi_n_86, csa_tree_add_7_25_groupi_n_87, csa_tree_add_7_25_groupi_n_88, csa_tree_add_7_25_groupi_n_89, csa_tree_add_7_25_groupi_n_90, csa_tree_add_7_25_groupi_n_91;
  wire csa_tree_add_7_25_groupi_n_92, csa_tree_add_7_25_groupi_n_93, csa_tree_add_7_25_groupi_n_94, csa_tree_add_7_25_groupi_n_95, csa_tree_add_7_25_groupi_n_96, csa_tree_add_7_25_groupi_n_97, csa_tree_add_7_25_groupi_n_98, csa_tree_add_7_25_groupi_n_99;
  wire csa_tree_add_7_25_groupi_n_100, csa_tree_add_7_25_groupi_n_101, csa_tree_add_7_25_groupi_n_102, csa_tree_add_7_25_groupi_n_103, csa_tree_add_7_25_groupi_n_104, csa_tree_add_7_25_groupi_n_105, csa_tree_add_7_25_groupi_n_106, csa_tree_add_7_25_groupi_n_107;
  wire csa_tree_add_7_25_groupi_n_108, csa_tree_add_7_25_groupi_n_109, csa_tree_add_7_25_groupi_n_110, csa_tree_add_7_25_groupi_n_111, csa_tree_add_7_25_groupi_n_112, csa_tree_add_7_25_groupi_n_113, csa_tree_add_7_25_groupi_n_114, csa_tree_add_7_25_groupi_n_115;
  wire csa_tree_add_7_25_groupi_n_116, csa_tree_add_7_25_groupi_n_117, csa_tree_add_7_25_groupi_n_118, csa_tree_add_7_25_groupi_n_119, csa_tree_add_7_25_groupi_n_120, csa_tree_add_7_25_groupi_n_121, csa_tree_add_7_25_groupi_n_122, csa_tree_add_7_25_groupi_n_123;
  wire csa_tree_add_7_25_groupi_n_124, csa_tree_add_7_25_groupi_n_125, csa_tree_add_7_25_groupi_n_126, csa_tree_add_7_25_groupi_n_127, csa_tree_add_7_25_groupi_n_128, csa_tree_add_7_25_groupi_n_129, csa_tree_add_7_25_groupi_n_130, csa_tree_add_7_25_groupi_n_131;
  wire csa_tree_add_7_25_groupi_n_132, csa_tree_add_7_25_groupi_n_133, csa_tree_add_7_25_groupi_n_134, csa_tree_add_7_25_groupi_n_135, csa_tree_add_7_25_groupi_n_136, csa_tree_add_7_25_groupi_n_137, csa_tree_add_7_25_groupi_n_138, csa_tree_add_7_25_groupi_n_139;
  wire csa_tree_add_7_25_groupi_n_140, csa_tree_add_7_25_groupi_n_141, csa_tree_add_7_25_groupi_n_142, csa_tree_add_7_25_groupi_n_143, csa_tree_add_7_25_groupi_n_144, csa_tree_add_7_25_groupi_n_145, csa_tree_add_7_25_groupi_n_146, csa_tree_add_7_25_groupi_n_147;
  wire csa_tree_add_7_25_groupi_n_148, csa_tree_add_7_25_groupi_n_149, csa_tree_add_7_25_groupi_n_150, csa_tree_add_7_25_groupi_n_151, csa_tree_add_7_25_groupi_n_152, csa_tree_add_7_25_groupi_n_153, csa_tree_add_7_25_groupi_n_154, csa_tree_add_7_25_groupi_n_155;
  wire csa_tree_add_7_25_groupi_n_156, csa_tree_add_7_25_groupi_n_157, csa_tree_add_7_25_groupi_n_158, csa_tree_add_7_25_groupi_n_159, csa_tree_add_7_25_groupi_n_160, csa_tree_add_7_25_groupi_n_161, csa_tree_add_7_25_groupi_n_162, csa_tree_add_7_25_groupi_n_163;
  wire csa_tree_add_7_25_groupi_n_164, csa_tree_add_7_25_groupi_n_165, csa_tree_add_7_25_groupi_n_166, csa_tree_add_7_25_groupi_n_167, csa_tree_add_7_25_groupi_n_168, csa_tree_add_7_25_groupi_n_169, csa_tree_add_7_25_groupi_n_170, csa_tree_add_7_25_groupi_n_171;
  wire csa_tree_add_7_25_groupi_n_172, csa_tree_add_7_25_groupi_n_173, csa_tree_add_7_25_groupi_n_174, csa_tree_add_7_25_groupi_n_175, csa_tree_add_7_25_groupi_n_176, csa_tree_add_7_25_groupi_n_177, csa_tree_add_7_25_groupi_n_178, csa_tree_add_7_25_groupi_n_179;
  wire csa_tree_add_7_25_groupi_n_180, csa_tree_add_7_25_groupi_n_181, csa_tree_add_7_25_groupi_n_182, csa_tree_add_7_25_groupi_n_183, csa_tree_add_7_25_groupi_n_184, csa_tree_add_7_25_groupi_n_185, csa_tree_add_7_25_groupi_n_186, csa_tree_add_7_25_groupi_n_187;
  wire csa_tree_add_7_25_groupi_n_188, csa_tree_add_7_25_groupi_n_189, csa_tree_add_7_25_groupi_n_190, csa_tree_add_7_25_groupi_n_191, csa_tree_add_7_25_groupi_n_192, csa_tree_add_7_25_groupi_n_193, csa_tree_add_7_25_groupi_n_194, csa_tree_add_7_25_groupi_n_195;
  wire csa_tree_add_7_25_groupi_n_196, csa_tree_add_7_25_groupi_n_197, csa_tree_add_7_25_groupi_n_198, csa_tree_add_7_25_groupi_n_199, csa_tree_add_7_25_groupi_n_200, csa_tree_add_7_25_groupi_n_201, csa_tree_add_7_25_groupi_n_202, csa_tree_add_7_25_groupi_n_203;
  wire csa_tree_add_7_25_groupi_n_204, csa_tree_add_7_25_groupi_n_205, csa_tree_add_7_25_groupi_n_206, csa_tree_add_7_25_groupi_n_207, csa_tree_add_7_25_groupi_n_208, csa_tree_add_7_25_groupi_n_209, csa_tree_add_7_25_groupi_n_210, csa_tree_add_7_25_groupi_n_211;
  wire csa_tree_add_7_25_groupi_n_212, csa_tree_add_7_25_groupi_n_213, csa_tree_add_7_25_groupi_n_214, csa_tree_add_7_25_groupi_n_215, csa_tree_add_7_25_groupi_n_216, csa_tree_add_7_25_groupi_n_217, csa_tree_add_7_25_groupi_n_218, csa_tree_add_7_25_groupi_n_219;
  wire csa_tree_add_7_25_groupi_n_220, csa_tree_add_7_25_groupi_n_221, csa_tree_add_7_25_groupi_n_222, csa_tree_add_7_25_groupi_n_223, csa_tree_add_7_25_groupi_n_224, csa_tree_add_7_25_groupi_n_225, csa_tree_add_7_25_groupi_n_226, csa_tree_add_7_25_groupi_n_227;
  wire csa_tree_add_7_25_groupi_n_228, csa_tree_add_7_25_groupi_n_229, csa_tree_add_7_25_groupi_n_230, csa_tree_add_7_25_groupi_n_231, csa_tree_add_7_25_groupi_n_232, csa_tree_add_7_25_groupi_n_233, csa_tree_add_7_25_groupi_n_234, csa_tree_add_7_25_groupi_n_235;
  wire csa_tree_add_7_25_groupi_n_236, csa_tree_add_7_25_groupi_n_237, csa_tree_add_7_25_groupi_n_238, csa_tree_add_7_25_groupi_n_239, csa_tree_add_7_25_groupi_n_240, csa_tree_add_7_25_groupi_n_241, csa_tree_add_7_25_groupi_n_242, csa_tree_add_7_25_groupi_n_243;
  wire csa_tree_add_7_25_groupi_n_244, csa_tree_add_7_25_groupi_n_245, csa_tree_add_7_25_groupi_n_246, csa_tree_add_7_25_groupi_n_247, csa_tree_add_7_25_groupi_n_248, csa_tree_add_7_25_groupi_n_249, csa_tree_add_7_25_groupi_n_250, csa_tree_add_7_25_groupi_n_251;
  wire csa_tree_add_7_25_groupi_n_252, csa_tree_add_7_25_groupi_n_253, csa_tree_add_7_25_groupi_n_254, csa_tree_add_7_25_groupi_n_255, csa_tree_add_7_25_groupi_n_256, csa_tree_add_7_25_groupi_n_257, csa_tree_add_7_25_groupi_n_258, csa_tree_add_7_25_groupi_n_259;
  wire csa_tree_add_7_25_groupi_n_260, csa_tree_add_7_25_groupi_n_261, csa_tree_add_7_25_groupi_n_262, csa_tree_add_7_25_groupi_n_263, csa_tree_add_7_25_groupi_n_264, csa_tree_add_7_25_groupi_n_265, csa_tree_add_7_25_groupi_n_266, csa_tree_add_7_25_groupi_n_267;
  wire csa_tree_add_7_25_groupi_n_268, csa_tree_add_7_25_groupi_n_269, csa_tree_add_7_25_groupi_n_270, csa_tree_add_7_25_groupi_n_271, csa_tree_add_7_25_groupi_n_272, csa_tree_add_7_25_groupi_n_273, csa_tree_add_7_25_groupi_n_274, csa_tree_add_7_25_groupi_n_275;
  wire csa_tree_add_7_25_groupi_n_276, csa_tree_add_7_25_groupi_n_277, csa_tree_add_7_25_groupi_n_278, csa_tree_add_7_25_groupi_n_279, csa_tree_add_7_25_groupi_n_280, csa_tree_add_7_25_groupi_n_281, csa_tree_add_7_25_groupi_n_282, csa_tree_add_7_25_groupi_n_283;
  wire csa_tree_add_7_25_groupi_n_284, csa_tree_add_7_25_groupi_n_285, csa_tree_add_7_25_groupi_n_286, csa_tree_add_7_25_groupi_n_287, csa_tree_add_7_25_groupi_n_288, csa_tree_add_7_25_groupi_n_289, csa_tree_add_7_25_groupi_n_290, csa_tree_add_7_25_groupi_n_291;
  wire csa_tree_add_7_25_groupi_n_292, csa_tree_add_7_25_groupi_n_293, csa_tree_add_7_25_groupi_n_294, csa_tree_add_7_25_groupi_n_295, csa_tree_add_7_25_groupi_n_296, csa_tree_add_7_25_groupi_n_297, csa_tree_add_7_25_groupi_n_298, csa_tree_add_7_25_groupi_n_299;
  wire csa_tree_add_7_25_groupi_n_300, csa_tree_add_7_25_groupi_n_301, csa_tree_add_7_25_groupi_n_302, csa_tree_add_7_25_groupi_n_303, csa_tree_add_7_25_groupi_n_304, csa_tree_add_7_25_groupi_n_305, csa_tree_add_7_25_groupi_n_306, csa_tree_add_7_25_groupi_n_307;
  wire csa_tree_add_7_25_groupi_n_308, csa_tree_add_7_25_groupi_n_309, csa_tree_add_7_25_groupi_n_310, csa_tree_add_7_25_groupi_n_311, csa_tree_add_7_25_groupi_n_312, csa_tree_add_7_25_groupi_n_313, csa_tree_add_7_25_groupi_n_314, csa_tree_add_7_25_groupi_n_315;
  wire csa_tree_add_7_25_groupi_n_316, csa_tree_add_7_25_groupi_n_317, csa_tree_add_7_25_groupi_n_318, csa_tree_add_7_25_groupi_n_319, csa_tree_add_7_25_groupi_n_320, csa_tree_add_7_25_groupi_n_321, csa_tree_add_7_25_groupi_n_322, csa_tree_add_7_25_groupi_n_323;
  wire csa_tree_add_7_25_groupi_n_324, csa_tree_add_7_25_groupi_n_325, csa_tree_add_7_25_groupi_n_326, csa_tree_add_7_25_groupi_n_327, csa_tree_add_7_25_groupi_n_328, csa_tree_add_7_25_groupi_n_329, csa_tree_add_7_25_groupi_n_330, csa_tree_add_7_25_groupi_n_331;
  wire csa_tree_add_7_25_groupi_n_332, csa_tree_add_7_25_groupi_n_333, csa_tree_add_7_25_groupi_n_334, csa_tree_add_7_25_groupi_n_335, csa_tree_add_7_25_groupi_n_336, csa_tree_add_7_25_groupi_n_337, csa_tree_add_7_25_groupi_n_338, csa_tree_add_7_25_groupi_n_339;
  wire csa_tree_add_7_25_groupi_n_340, csa_tree_add_7_25_groupi_n_341, csa_tree_add_7_25_groupi_n_342, csa_tree_add_7_25_groupi_n_343, csa_tree_add_7_25_groupi_n_344, csa_tree_add_7_25_groupi_n_345, csa_tree_add_7_25_groupi_n_346, csa_tree_add_7_25_groupi_n_347;
  wire csa_tree_add_7_25_groupi_n_348, csa_tree_add_7_25_groupi_n_349, csa_tree_add_7_25_groupi_n_350, csa_tree_add_7_25_groupi_n_351, csa_tree_add_7_25_groupi_n_352, csa_tree_add_7_25_groupi_n_353, csa_tree_add_7_25_groupi_n_354, csa_tree_add_7_25_groupi_n_355;
  wire csa_tree_add_7_25_groupi_n_356, csa_tree_add_7_25_groupi_n_357, csa_tree_add_7_25_groupi_n_358, csa_tree_add_7_25_groupi_n_359, csa_tree_add_7_25_groupi_n_360, csa_tree_add_7_25_groupi_n_361, csa_tree_add_7_25_groupi_n_362, csa_tree_add_7_25_groupi_n_363;
  wire csa_tree_add_7_25_groupi_n_364, csa_tree_add_7_25_groupi_n_365, csa_tree_add_7_25_groupi_n_366, csa_tree_add_7_25_groupi_n_367, csa_tree_add_7_25_groupi_n_368, csa_tree_add_7_25_groupi_n_369, csa_tree_add_7_25_groupi_n_370, csa_tree_add_7_25_groupi_n_371;
  wire csa_tree_add_7_25_groupi_n_372, csa_tree_add_7_25_groupi_n_373, csa_tree_add_7_25_groupi_n_374, csa_tree_add_7_25_groupi_n_375, csa_tree_add_7_25_groupi_n_376, csa_tree_add_7_25_groupi_n_377, csa_tree_add_7_25_groupi_n_378, csa_tree_add_7_25_groupi_n_379;
  wire csa_tree_add_7_25_groupi_n_380, csa_tree_add_7_25_groupi_n_381, csa_tree_add_7_25_groupi_n_382, csa_tree_add_7_25_groupi_n_383, csa_tree_add_7_25_groupi_n_384, csa_tree_add_7_25_groupi_n_385, csa_tree_add_7_25_groupi_n_386, csa_tree_add_7_25_groupi_n_387;
  wire csa_tree_add_7_25_groupi_n_388, csa_tree_add_7_25_groupi_n_389, csa_tree_add_7_25_groupi_n_390, csa_tree_add_7_25_groupi_n_391, csa_tree_add_7_25_groupi_n_392, csa_tree_add_7_25_groupi_n_393, csa_tree_add_7_25_groupi_n_394, csa_tree_add_7_25_groupi_n_395;
  wire csa_tree_add_7_25_groupi_n_396, csa_tree_add_7_25_groupi_n_397, csa_tree_add_7_25_groupi_n_398, csa_tree_add_7_25_groupi_n_399, csa_tree_add_7_25_groupi_n_400, csa_tree_add_7_25_groupi_n_401, csa_tree_add_7_25_groupi_n_402, csa_tree_add_7_25_groupi_n_403;
  wire csa_tree_add_7_25_groupi_n_404, csa_tree_add_7_25_groupi_n_405, csa_tree_add_7_25_groupi_n_406, csa_tree_add_7_25_groupi_n_407, csa_tree_add_7_25_groupi_n_408, csa_tree_add_7_25_groupi_n_409, csa_tree_add_7_25_groupi_n_410, csa_tree_add_7_25_groupi_n_411;
  wire csa_tree_add_7_25_groupi_n_412, csa_tree_add_7_25_groupi_n_413, csa_tree_add_7_25_groupi_n_414, csa_tree_add_7_25_groupi_n_415, csa_tree_add_7_25_groupi_n_416, csa_tree_add_7_25_groupi_n_417, csa_tree_add_7_25_groupi_n_418, csa_tree_add_7_25_groupi_n_419;
  wire csa_tree_add_7_25_groupi_n_420, csa_tree_add_7_25_groupi_n_421, csa_tree_add_7_25_groupi_n_422, csa_tree_add_7_25_groupi_n_423, csa_tree_add_7_25_groupi_n_424, csa_tree_add_7_25_groupi_n_425, csa_tree_add_7_25_groupi_n_426, csa_tree_add_7_25_groupi_n_427;
  wire csa_tree_add_7_25_groupi_n_428, csa_tree_add_7_25_groupi_n_429, csa_tree_add_7_25_groupi_n_430, csa_tree_add_7_25_groupi_n_431, csa_tree_add_7_25_groupi_n_432, csa_tree_add_7_25_groupi_n_433, csa_tree_add_7_25_groupi_n_434, csa_tree_add_7_25_groupi_n_435;
  wire csa_tree_add_7_25_groupi_n_436, csa_tree_add_7_25_groupi_n_437, csa_tree_add_7_25_groupi_n_438, csa_tree_add_7_25_groupi_n_439, csa_tree_add_7_25_groupi_n_440, csa_tree_add_7_25_groupi_n_441, csa_tree_add_7_25_groupi_n_442, csa_tree_add_7_25_groupi_n_443;
  wire csa_tree_add_7_25_groupi_n_444, csa_tree_add_7_25_groupi_n_445, csa_tree_add_7_25_groupi_n_446, csa_tree_add_7_25_groupi_n_447, csa_tree_add_7_25_groupi_n_448, csa_tree_add_7_25_groupi_n_449, csa_tree_add_7_25_groupi_n_450, csa_tree_add_7_25_groupi_n_451;
  wire csa_tree_add_7_25_groupi_n_452, csa_tree_add_7_25_groupi_n_453, csa_tree_add_7_25_groupi_n_454, csa_tree_add_7_25_groupi_n_455, csa_tree_add_7_25_groupi_n_456, csa_tree_add_7_25_groupi_n_457, csa_tree_add_7_25_groupi_n_458, csa_tree_add_7_25_groupi_n_459;
  wire csa_tree_add_7_25_groupi_n_460, csa_tree_add_7_25_groupi_n_461, csa_tree_add_7_25_groupi_n_462, csa_tree_add_7_25_groupi_n_463, csa_tree_add_7_25_groupi_n_464, csa_tree_add_7_25_groupi_n_465, csa_tree_add_7_25_groupi_n_466, csa_tree_add_7_25_groupi_n_467;
  wire csa_tree_add_7_25_groupi_n_468, csa_tree_add_7_25_groupi_n_469, csa_tree_add_7_25_groupi_n_470, csa_tree_add_7_25_groupi_n_471, csa_tree_add_7_25_groupi_n_472, csa_tree_add_7_25_groupi_n_473, csa_tree_add_7_25_groupi_n_474, csa_tree_add_7_25_groupi_n_475;
  wire csa_tree_add_7_25_groupi_n_476, csa_tree_add_7_25_groupi_n_477, csa_tree_add_7_25_groupi_n_478, csa_tree_add_7_25_groupi_n_479, csa_tree_add_7_25_groupi_n_480, csa_tree_add_7_25_groupi_n_481, csa_tree_add_7_25_groupi_n_482, csa_tree_add_7_25_groupi_n_483;
  wire csa_tree_add_7_25_groupi_n_484, csa_tree_add_7_25_groupi_n_485, csa_tree_add_7_25_groupi_n_486, csa_tree_add_7_25_groupi_n_487, csa_tree_add_7_25_groupi_n_488, csa_tree_add_7_25_groupi_n_489, csa_tree_add_7_25_groupi_n_490, csa_tree_add_7_25_groupi_n_491;
  wire csa_tree_add_7_25_groupi_n_492, csa_tree_add_7_25_groupi_n_493, csa_tree_add_7_25_groupi_n_494, csa_tree_add_7_25_groupi_n_495, csa_tree_add_7_25_groupi_n_496, csa_tree_add_7_25_groupi_n_497, csa_tree_add_7_25_groupi_n_498, csa_tree_add_7_25_groupi_n_499;
  wire csa_tree_add_7_25_groupi_n_500, csa_tree_add_7_25_groupi_n_501, csa_tree_add_7_25_groupi_n_502, csa_tree_add_7_25_groupi_n_503, csa_tree_add_7_25_groupi_n_504, csa_tree_add_7_25_groupi_n_505, csa_tree_add_7_25_groupi_n_506, csa_tree_add_7_25_groupi_n_507;
  wire csa_tree_add_7_25_groupi_n_508, csa_tree_add_7_25_groupi_n_509, csa_tree_add_7_25_groupi_n_510, csa_tree_add_7_25_groupi_n_511, csa_tree_add_7_25_groupi_n_512, csa_tree_add_7_25_groupi_n_513, csa_tree_add_7_25_groupi_n_514, csa_tree_add_7_25_groupi_n_515;
  wire csa_tree_add_7_25_groupi_n_516, csa_tree_add_7_25_groupi_n_517, csa_tree_add_7_25_groupi_n_518, csa_tree_add_7_25_groupi_n_519, csa_tree_add_7_25_groupi_n_520, csa_tree_add_7_25_groupi_n_521, csa_tree_add_7_25_groupi_n_522, csa_tree_add_7_25_groupi_n_523;
  wire csa_tree_add_7_25_groupi_n_524, csa_tree_add_7_25_groupi_n_525, csa_tree_add_7_25_groupi_n_526, csa_tree_add_7_25_groupi_n_527, csa_tree_add_7_25_groupi_n_528, csa_tree_add_7_25_groupi_n_529, csa_tree_add_7_25_groupi_n_530, csa_tree_add_7_25_groupi_n_531;
  wire csa_tree_add_7_25_groupi_n_532, csa_tree_add_7_25_groupi_n_533, csa_tree_add_7_25_groupi_n_534, csa_tree_add_7_25_groupi_n_535, csa_tree_add_7_25_groupi_n_536, csa_tree_add_7_25_groupi_n_537, csa_tree_add_7_25_groupi_n_538, csa_tree_add_7_25_groupi_n_539;
  wire csa_tree_add_7_25_groupi_n_540, csa_tree_add_7_25_groupi_n_541, csa_tree_add_7_25_groupi_n_542, csa_tree_add_7_25_groupi_n_543, csa_tree_add_7_25_groupi_n_544, csa_tree_add_7_25_groupi_n_545, csa_tree_add_7_25_groupi_n_546, csa_tree_add_7_25_groupi_n_547;
  wire csa_tree_add_7_25_groupi_n_548, csa_tree_add_7_25_groupi_n_549, csa_tree_add_7_25_groupi_n_550, csa_tree_add_7_25_groupi_n_551, csa_tree_add_7_25_groupi_n_552, csa_tree_add_7_25_groupi_n_553, csa_tree_add_7_25_groupi_n_554, csa_tree_add_7_25_groupi_n_555;
  wire csa_tree_add_7_25_groupi_n_556, csa_tree_add_7_25_groupi_n_557, csa_tree_add_7_25_groupi_n_558, csa_tree_add_7_25_groupi_n_559, csa_tree_add_7_25_groupi_n_560, csa_tree_add_7_25_groupi_n_561, csa_tree_add_7_25_groupi_n_562, csa_tree_add_7_25_groupi_n_563;
  wire csa_tree_add_7_25_groupi_n_564, csa_tree_add_7_25_groupi_n_565, csa_tree_add_7_25_groupi_n_566, csa_tree_add_7_25_groupi_n_567, csa_tree_add_7_25_groupi_n_568, csa_tree_add_7_25_groupi_n_569, csa_tree_add_7_25_groupi_n_570, csa_tree_add_7_25_groupi_n_571;
  wire csa_tree_add_7_25_groupi_n_572, csa_tree_add_7_25_groupi_n_573, csa_tree_add_7_25_groupi_n_574, csa_tree_add_7_25_groupi_n_575, csa_tree_add_7_25_groupi_n_576, csa_tree_add_7_25_groupi_n_577, csa_tree_add_7_25_groupi_n_578, csa_tree_add_7_25_groupi_n_579;
  wire csa_tree_add_7_25_groupi_n_580, csa_tree_add_7_25_groupi_n_581, csa_tree_add_7_25_groupi_n_582, csa_tree_add_7_25_groupi_n_583, csa_tree_add_7_25_groupi_n_584, csa_tree_add_7_25_groupi_n_585, csa_tree_add_7_25_groupi_n_586, csa_tree_add_7_25_groupi_n_587;
  wire csa_tree_add_7_25_groupi_n_588, csa_tree_add_7_25_groupi_n_589, csa_tree_add_7_25_groupi_n_590, csa_tree_add_7_25_groupi_n_591, csa_tree_add_7_25_groupi_n_592, csa_tree_add_7_25_groupi_n_593, csa_tree_add_7_25_groupi_n_594, csa_tree_add_7_25_groupi_n_595;
  wire csa_tree_add_7_25_groupi_n_596, csa_tree_add_7_25_groupi_n_597, csa_tree_add_7_25_groupi_n_598, csa_tree_add_7_25_groupi_n_599, csa_tree_add_7_25_groupi_n_600, csa_tree_add_7_25_groupi_n_601, csa_tree_add_7_25_groupi_n_602, csa_tree_add_7_25_groupi_n_603;
  wire csa_tree_add_7_25_groupi_n_604, csa_tree_add_7_25_groupi_n_605, csa_tree_add_7_25_groupi_n_606, csa_tree_add_7_25_groupi_n_607, csa_tree_add_7_25_groupi_n_608, csa_tree_add_7_25_groupi_n_609, csa_tree_add_7_25_groupi_n_610, csa_tree_add_7_25_groupi_n_611;
  wire csa_tree_add_7_25_groupi_n_612, csa_tree_add_7_25_groupi_n_613, csa_tree_add_7_25_groupi_n_614, csa_tree_add_7_25_groupi_n_615, csa_tree_add_7_25_groupi_n_616, csa_tree_add_7_25_groupi_n_617, csa_tree_add_7_25_groupi_n_618, csa_tree_add_7_25_groupi_n_619;
  wire csa_tree_add_7_25_groupi_n_620, csa_tree_add_7_25_groupi_n_621, csa_tree_add_7_25_groupi_n_622, csa_tree_add_7_25_groupi_n_623, csa_tree_add_7_25_groupi_n_624, csa_tree_add_7_25_groupi_n_625, csa_tree_add_7_25_groupi_n_626, csa_tree_add_7_25_groupi_n_627;
  wire csa_tree_add_7_25_groupi_n_628, csa_tree_add_7_25_groupi_n_629, csa_tree_add_7_25_groupi_n_630, csa_tree_add_7_25_groupi_n_631, csa_tree_add_7_25_groupi_n_632, csa_tree_add_7_25_groupi_n_633, csa_tree_add_7_25_groupi_n_634, csa_tree_add_7_25_groupi_n_635;
  wire csa_tree_add_7_25_groupi_n_636, csa_tree_add_7_25_groupi_n_637, csa_tree_add_7_25_groupi_n_638, csa_tree_add_7_25_groupi_n_639, csa_tree_add_7_25_groupi_n_640, csa_tree_add_7_25_groupi_n_641, csa_tree_add_7_25_groupi_n_642, csa_tree_add_7_25_groupi_n_643;
  wire csa_tree_add_7_25_groupi_n_644, csa_tree_add_7_25_groupi_n_645, csa_tree_add_7_25_groupi_n_646, csa_tree_add_7_25_groupi_n_647, csa_tree_add_7_25_groupi_n_648, csa_tree_add_7_25_groupi_n_649, csa_tree_add_7_25_groupi_n_650, csa_tree_add_7_25_groupi_n_651;
  wire csa_tree_add_7_25_groupi_n_652, csa_tree_add_7_25_groupi_n_653, csa_tree_add_7_25_groupi_n_654, csa_tree_add_7_25_groupi_n_655, csa_tree_add_7_25_groupi_n_656, csa_tree_add_7_25_groupi_n_657, csa_tree_add_7_25_groupi_n_658, csa_tree_add_7_25_groupi_n_659;
  wire csa_tree_add_7_25_groupi_n_660, csa_tree_add_7_25_groupi_n_661, csa_tree_add_7_25_groupi_n_662, csa_tree_add_7_25_groupi_n_663, csa_tree_add_7_25_groupi_n_664, csa_tree_add_7_25_groupi_n_665, csa_tree_add_7_25_groupi_n_666, csa_tree_add_7_25_groupi_n_667;
  wire csa_tree_add_7_25_groupi_n_668, csa_tree_add_7_25_groupi_n_669, csa_tree_add_7_25_groupi_n_670, csa_tree_add_7_25_groupi_n_671, csa_tree_add_7_25_groupi_n_672, csa_tree_add_7_25_groupi_n_673, csa_tree_add_7_25_groupi_n_674, csa_tree_add_7_25_groupi_n_675;
  wire csa_tree_add_7_25_groupi_n_676, csa_tree_add_7_25_groupi_n_677, csa_tree_add_7_25_groupi_n_678, csa_tree_add_7_25_groupi_n_679, csa_tree_add_7_25_groupi_n_680, csa_tree_add_7_25_groupi_n_681, csa_tree_add_7_25_groupi_n_682, csa_tree_add_7_25_groupi_n_683;
  wire csa_tree_add_7_25_groupi_n_684, csa_tree_add_7_25_groupi_n_685, csa_tree_add_7_25_groupi_n_686, csa_tree_add_7_25_groupi_n_687, csa_tree_add_7_25_groupi_n_688, csa_tree_add_7_25_groupi_n_689, csa_tree_add_7_25_groupi_n_690, csa_tree_add_7_25_groupi_n_691;
  wire csa_tree_add_7_25_groupi_n_692, csa_tree_add_7_25_groupi_n_693, csa_tree_add_7_25_groupi_n_694, csa_tree_add_7_25_groupi_n_695, csa_tree_add_7_25_groupi_n_696, csa_tree_add_7_25_groupi_n_697, csa_tree_add_7_25_groupi_n_698, csa_tree_add_7_25_groupi_n_699;
  wire csa_tree_add_7_25_groupi_n_700, csa_tree_add_7_25_groupi_n_701, csa_tree_add_7_25_groupi_n_702, csa_tree_add_7_25_groupi_n_703, csa_tree_add_7_25_groupi_n_704, csa_tree_add_7_25_groupi_n_705, csa_tree_add_7_25_groupi_n_706, csa_tree_add_7_25_groupi_n_707;
  wire csa_tree_add_7_25_groupi_n_708, csa_tree_add_7_25_groupi_n_709, csa_tree_add_7_25_groupi_n_710, csa_tree_add_7_25_groupi_n_711, csa_tree_add_7_25_groupi_n_712, csa_tree_add_7_25_groupi_n_713, csa_tree_add_7_25_groupi_n_714, csa_tree_add_7_25_groupi_n_715;
  wire csa_tree_add_7_25_groupi_n_716, csa_tree_add_7_25_groupi_n_717, csa_tree_add_7_25_groupi_n_718, csa_tree_add_7_25_groupi_n_719, csa_tree_add_7_25_groupi_n_720, csa_tree_add_7_25_groupi_n_721, csa_tree_add_7_25_groupi_n_722, csa_tree_add_7_25_groupi_n_723;
  wire csa_tree_add_7_25_groupi_n_724, csa_tree_add_7_25_groupi_n_725, csa_tree_add_7_25_groupi_n_726, csa_tree_add_7_25_groupi_n_727, csa_tree_add_7_25_groupi_n_728, csa_tree_add_7_25_groupi_n_729, csa_tree_add_7_25_groupi_n_730, csa_tree_add_7_25_groupi_n_731;
  wire csa_tree_add_7_25_groupi_n_732, csa_tree_add_7_25_groupi_n_733, csa_tree_add_7_25_groupi_n_734, csa_tree_add_7_25_groupi_n_735, csa_tree_add_7_25_groupi_n_736, csa_tree_add_7_25_groupi_n_737, csa_tree_add_7_25_groupi_n_738, csa_tree_add_7_25_groupi_n_739;
  wire csa_tree_add_7_25_groupi_n_740, csa_tree_add_7_25_groupi_n_741, csa_tree_add_7_25_groupi_n_742, csa_tree_add_7_25_groupi_n_743, csa_tree_add_7_25_groupi_n_744, csa_tree_add_7_25_groupi_n_745, csa_tree_add_7_25_groupi_n_746, csa_tree_add_7_25_groupi_n_747;
  wire csa_tree_add_7_25_groupi_n_748, csa_tree_add_7_25_groupi_n_749, csa_tree_add_7_25_groupi_n_750, csa_tree_add_7_25_groupi_n_751, csa_tree_add_7_25_groupi_n_752, csa_tree_add_7_25_groupi_n_753, csa_tree_add_7_25_groupi_n_754, csa_tree_add_7_25_groupi_n_755;
  wire csa_tree_add_7_25_groupi_n_756, csa_tree_add_7_25_groupi_n_757, csa_tree_add_7_25_groupi_n_758, csa_tree_add_7_25_groupi_n_759, csa_tree_add_7_25_groupi_n_760, csa_tree_add_7_25_groupi_n_761, csa_tree_add_7_25_groupi_n_762, csa_tree_add_7_25_groupi_n_763;
  wire csa_tree_add_7_25_groupi_n_764, csa_tree_add_7_25_groupi_n_765, csa_tree_add_7_25_groupi_n_766, csa_tree_add_7_25_groupi_n_767, csa_tree_add_7_25_groupi_n_768, csa_tree_add_7_25_groupi_n_769, csa_tree_add_7_25_groupi_n_770, csa_tree_add_7_25_groupi_n_771;
  wire csa_tree_add_7_25_groupi_n_772, csa_tree_add_7_25_groupi_n_773, csa_tree_add_7_25_groupi_n_774, csa_tree_add_7_25_groupi_n_775, csa_tree_add_7_25_groupi_n_776, csa_tree_add_7_25_groupi_n_777, csa_tree_add_7_25_groupi_n_778, csa_tree_add_7_25_groupi_n_779;
  wire csa_tree_add_7_25_groupi_n_780, csa_tree_add_7_25_groupi_n_781, csa_tree_add_7_25_groupi_n_782, csa_tree_add_7_25_groupi_n_783, csa_tree_add_7_25_groupi_n_784, csa_tree_add_7_25_groupi_n_785, csa_tree_add_7_25_groupi_n_786, csa_tree_add_7_25_groupi_n_787;
  wire csa_tree_add_7_25_groupi_n_788, csa_tree_add_7_25_groupi_n_789, csa_tree_add_7_25_groupi_n_790, csa_tree_add_7_25_groupi_n_791, csa_tree_add_7_25_groupi_n_792, csa_tree_add_7_25_groupi_n_793, csa_tree_add_7_25_groupi_n_794, csa_tree_add_7_25_groupi_n_795;
  wire csa_tree_add_7_25_groupi_n_796, csa_tree_add_7_25_groupi_n_797, csa_tree_add_7_25_groupi_n_798, csa_tree_add_7_25_groupi_n_799, csa_tree_add_7_25_groupi_n_800, csa_tree_add_7_25_groupi_n_801, csa_tree_add_7_25_groupi_n_802, csa_tree_add_7_25_groupi_n_803;
  wire csa_tree_add_7_25_groupi_n_804, csa_tree_add_7_25_groupi_n_805, csa_tree_add_7_25_groupi_n_806, csa_tree_add_7_25_groupi_n_807, csa_tree_add_7_25_groupi_n_808, csa_tree_add_7_25_groupi_n_809, csa_tree_add_7_25_groupi_n_810, csa_tree_add_7_25_groupi_n_811;
  wire csa_tree_add_7_25_groupi_n_812, csa_tree_add_7_25_groupi_n_813, csa_tree_add_7_25_groupi_n_814, csa_tree_add_7_25_groupi_n_815, csa_tree_add_7_25_groupi_n_816, csa_tree_add_7_25_groupi_n_817, csa_tree_add_7_25_groupi_n_818, csa_tree_add_7_25_groupi_n_819;
  wire csa_tree_add_7_25_groupi_n_820, csa_tree_add_7_25_groupi_n_821, csa_tree_add_7_25_groupi_n_822, csa_tree_add_7_25_groupi_n_823, csa_tree_add_7_25_groupi_n_824, csa_tree_add_7_25_groupi_n_825, csa_tree_add_7_25_groupi_n_826, csa_tree_add_7_25_groupi_n_827;
  wire csa_tree_add_7_25_groupi_n_828, csa_tree_add_7_25_groupi_n_829, csa_tree_add_7_25_groupi_n_830, csa_tree_add_7_25_groupi_n_831, csa_tree_add_7_25_groupi_n_832, csa_tree_add_7_25_groupi_n_833, csa_tree_add_7_25_groupi_n_834, csa_tree_add_7_25_groupi_n_835;
  wire csa_tree_add_7_25_groupi_n_836, csa_tree_add_7_25_groupi_n_837, csa_tree_add_7_25_groupi_n_838, csa_tree_add_7_25_groupi_n_839, csa_tree_add_7_25_groupi_n_840, csa_tree_add_7_25_groupi_n_841, csa_tree_add_7_25_groupi_n_842, csa_tree_add_7_25_groupi_n_843;
  wire csa_tree_add_7_25_groupi_n_844, csa_tree_add_7_25_groupi_n_845, csa_tree_add_7_25_groupi_n_846, csa_tree_add_7_25_groupi_n_847, csa_tree_add_7_25_groupi_n_848, csa_tree_add_7_25_groupi_n_849, csa_tree_add_7_25_groupi_n_850, csa_tree_add_7_25_groupi_n_851;
  wire csa_tree_add_7_25_groupi_n_852, csa_tree_add_7_25_groupi_n_853, csa_tree_add_7_25_groupi_n_854, csa_tree_add_7_25_groupi_n_855, csa_tree_add_7_25_groupi_n_856, csa_tree_add_7_25_groupi_n_857, csa_tree_add_7_25_groupi_n_858, csa_tree_add_7_25_groupi_n_859;
  wire csa_tree_add_7_25_groupi_n_860, csa_tree_add_7_25_groupi_n_861, csa_tree_add_7_25_groupi_n_862, csa_tree_add_7_25_groupi_n_863, csa_tree_add_7_25_groupi_n_864, csa_tree_add_7_25_groupi_n_865, csa_tree_add_7_25_groupi_n_866, csa_tree_add_7_25_groupi_n_867;
  wire csa_tree_add_7_25_groupi_n_868, csa_tree_add_7_25_groupi_n_869, csa_tree_add_7_25_groupi_n_870, csa_tree_add_7_25_groupi_n_871, csa_tree_add_7_25_groupi_n_872, csa_tree_add_7_25_groupi_n_873, csa_tree_add_7_25_groupi_n_874, csa_tree_add_7_25_groupi_n_875;
  wire csa_tree_add_7_25_groupi_n_876, csa_tree_add_7_25_groupi_n_877, csa_tree_add_7_25_groupi_n_878, csa_tree_add_7_25_groupi_n_879, csa_tree_add_7_25_groupi_n_880, csa_tree_add_7_25_groupi_n_881, csa_tree_add_7_25_groupi_n_882, csa_tree_add_7_25_groupi_n_883;
  wire csa_tree_add_7_25_groupi_n_884, csa_tree_add_7_25_groupi_n_885, csa_tree_add_7_25_groupi_n_886, csa_tree_add_7_25_groupi_n_887, csa_tree_add_7_25_groupi_n_888, csa_tree_add_7_25_groupi_n_889, csa_tree_add_7_25_groupi_n_890, csa_tree_add_7_25_groupi_n_891;
  wire csa_tree_add_7_25_groupi_n_892, csa_tree_add_7_25_groupi_n_893, csa_tree_add_7_25_groupi_n_894, csa_tree_add_7_25_groupi_n_895, csa_tree_add_7_25_groupi_n_896, csa_tree_add_7_25_groupi_n_897, csa_tree_add_7_25_groupi_n_898, csa_tree_add_7_25_groupi_n_899;
  wire csa_tree_add_7_25_groupi_n_900, csa_tree_add_7_25_groupi_n_901, csa_tree_add_7_25_groupi_n_902, csa_tree_add_7_25_groupi_n_903, csa_tree_add_7_25_groupi_n_904, csa_tree_add_7_25_groupi_n_905, csa_tree_add_7_25_groupi_n_906, csa_tree_add_7_25_groupi_n_907;
  wire csa_tree_add_7_25_groupi_n_908, csa_tree_add_7_25_groupi_n_909, csa_tree_add_7_25_groupi_n_910, csa_tree_add_7_25_groupi_n_911, csa_tree_add_7_25_groupi_n_912, csa_tree_add_7_25_groupi_n_913, csa_tree_add_7_25_groupi_n_914, csa_tree_add_7_25_groupi_n_915;
  wire csa_tree_add_7_25_groupi_n_916, csa_tree_add_7_25_groupi_n_917, csa_tree_add_7_25_groupi_n_918, csa_tree_add_7_25_groupi_n_919, csa_tree_add_7_25_groupi_n_920, csa_tree_add_7_25_groupi_n_921, csa_tree_add_7_25_groupi_n_922, csa_tree_add_7_25_groupi_n_923;
  wire csa_tree_add_7_25_groupi_n_924, csa_tree_add_7_25_groupi_n_925, csa_tree_add_7_25_groupi_n_926, csa_tree_add_7_25_groupi_n_927, csa_tree_add_7_25_groupi_n_928, csa_tree_add_7_25_groupi_n_929, csa_tree_add_7_25_groupi_n_930, csa_tree_add_7_25_groupi_n_931;
  wire csa_tree_add_7_25_groupi_n_932, csa_tree_add_7_25_groupi_n_933, csa_tree_add_7_25_groupi_n_934, csa_tree_add_7_25_groupi_n_935, csa_tree_add_7_25_groupi_n_936, csa_tree_add_7_25_groupi_n_937, csa_tree_add_7_25_groupi_n_938, csa_tree_add_7_25_groupi_n_939;
  wire csa_tree_add_7_25_groupi_n_940, csa_tree_add_7_25_groupi_n_941, csa_tree_add_7_25_groupi_n_942, csa_tree_add_7_25_groupi_n_943, csa_tree_add_7_25_groupi_n_944, csa_tree_add_7_25_groupi_n_945, csa_tree_add_7_25_groupi_n_946, csa_tree_add_7_25_groupi_n_947;
  wire csa_tree_add_7_25_groupi_n_948, csa_tree_add_7_25_groupi_n_949, csa_tree_add_7_25_groupi_n_950, csa_tree_add_7_25_groupi_n_951, csa_tree_add_7_25_groupi_n_952, csa_tree_add_7_25_groupi_n_953, csa_tree_add_7_25_groupi_n_954, csa_tree_add_7_25_groupi_n_955;
  wire csa_tree_add_7_25_groupi_n_956, csa_tree_add_7_25_groupi_n_957, csa_tree_add_7_25_groupi_n_958, csa_tree_add_7_25_groupi_n_959, csa_tree_add_7_25_groupi_n_960, csa_tree_add_7_25_groupi_n_961, csa_tree_add_7_25_groupi_n_962, csa_tree_add_7_25_groupi_n_963;
  wire csa_tree_add_7_25_groupi_n_964, csa_tree_add_7_25_groupi_n_965, csa_tree_add_7_25_groupi_n_966, csa_tree_add_7_25_groupi_n_967, csa_tree_add_7_25_groupi_n_968, csa_tree_add_7_25_groupi_n_969, csa_tree_add_7_25_groupi_n_970, csa_tree_add_7_25_groupi_n_971;
  wire csa_tree_add_7_25_groupi_n_972, csa_tree_add_7_25_groupi_n_973, csa_tree_add_7_25_groupi_n_974, csa_tree_add_7_25_groupi_n_975, csa_tree_add_7_25_groupi_n_976, csa_tree_add_7_25_groupi_n_977, csa_tree_add_7_25_groupi_n_978, csa_tree_add_7_25_groupi_n_979;
  wire csa_tree_add_7_25_groupi_n_980, csa_tree_add_7_25_groupi_n_981, csa_tree_add_7_25_groupi_n_982, csa_tree_add_7_25_groupi_n_983, csa_tree_add_7_25_groupi_n_984, csa_tree_add_7_25_groupi_n_985, csa_tree_add_7_25_groupi_n_986, csa_tree_add_7_25_groupi_n_987;
  wire csa_tree_add_7_25_groupi_n_988, csa_tree_add_7_25_groupi_n_989, csa_tree_add_7_25_groupi_n_990, csa_tree_add_7_25_groupi_n_991, csa_tree_add_7_25_groupi_n_992, csa_tree_add_7_25_groupi_n_993, csa_tree_add_7_25_groupi_n_994, csa_tree_add_7_25_groupi_n_995;
  wire csa_tree_add_7_25_groupi_n_996, csa_tree_add_7_25_groupi_n_997, csa_tree_add_7_25_groupi_n_998, csa_tree_add_7_25_groupi_n_999, csa_tree_add_7_25_groupi_n_1000, csa_tree_add_7_25_groupi_n_1001, csa_tree_add_7_25_groupi_n_1002, csa_tree_add_7_25_groupi_n_1003;
  wire csa_tree_add_7_25_groupi_n_1004, csa_tree_add_7_25_groupi_n_1005, csa_tree_add_7_25_groupi_n_1006, csa_tree_add_7_25_groupi_n_1007, csa_tree_add_7_25_groupi_n_1008, csa_tree_add_7_25_groupi_n_1009, csa_tree_add_7_25_groupi_n_1010, csa_tree_add_7_25_groupi_n_1011;
  wire csa_tree_add_7_25_groupi_n_1012, csa_tree_add_7_25_groupi_n_1013, csa_tree_add_7_25_groupi_n_1014, csa_tree_add_7_25_groupi_n_1015, csa_tree_add_7_25_groupi_n_1016, csa_tree_add_7_25_groupi_n_1017, csa_tree_add_7_25_groupi_n_1018, csa_tree_add_7_25_groupi_n_1019;
  wire csa_tree_add_7_25_groupi_n_1020, csa_tree_add_7_25_groupi_n_1021, csa_tree_add_7_25_groupi_n_1022, csa_tree_add_7_25_groupi_n_1023, csa_tree_add_7_25_groupi_n_1024, csa_tree_add_7_25_groupi_n_1025, csa_tree_add_7_25_groupi_n_1026, csa_tree_add_7_25_groupi_n_1027;
  wire csa_tree_add_7_25_groupi_n_1028, csa_tree_add_7_25_groupi_n_1029, csa_tree_add_7_25_groupi_n_1030, csa_tree_add_7_25_groupi_n_1031, csa_tree_add_7_25_groupi_n_1032, csa_tree_add_7_25_groupi_n_1033, csa_tree_add_7_25_groupi_n_1034, csa_tree_add_7_25_groupi_n_1035;
  wire csa_tree_add_7_25_groupi_n_1036, csa_tree_add_7_25_groupi_n_1037, csa_tree_add_7_25_groupi_n_1038, csa_tree_add_7_25_groupi_n_1039, csa_tree_add_7_25_groupi_n_1040, csa_tree_add_7_25_groupi_n_1041, csa_tree_add_7_25_groupi_n_1042, csa_tree_add_7_25_groupi_n_1043;
  wire csa_tree_add_7_25_groupi_n_1044, csa_tree_add_7_25_groupi_n_1045, csa_tree_add_7_25_groupi_n_1046, csa_tree_add_7_25_groupi_n_1047, csa_tree_add_7_25_groupi_n_1048, csa_tree_add_7_25_groupi_n_1049, csa_tree_add_7_25_groupi_n_1050, csa_tree_add_7_25_groupi_n_1051;
  wire csa_tree_add_7_25_groupi_n_1052, csa_tree_add_7_25_groupi_n_1053, csa_tree_add_7_25_groupi_n_1054, csa_tree_add_7_25_groupi_n_1055, csa_tree_add_7_25_groupi_n_1056, csa_tree_add_7_25_groupi_n_1057, csa_tree_add_7_25_groupi_n_1058, csa_tree_add_7_25_groupi_n_1059;
  wire csa_tree_add_7_25_groupi_n_1060, csa_tree_add_7_25_groupi_n_1061, csa_tree_add_7_25_groupi_n_1062, csa_tree_add_7_25_groupi_n_1063, csa_tree_add_7_25_groupi_n_1064, csa_tree_add_7_25_groupi_n_1065, csa_tree_add_7_25_groupi_n_1066, csa_tree_add_7_25_groupi_n_1067;
  wire csa_tree_add_7_25_groupi_n_1068, csa_tree_add_7_25_groupi_n_1069, csa_tree_add_7_25_groupi_n_1070, csa_tree_add_7_25_groupi_n_1071, csa_tree_add_7_25_groupi_n_1072, csa_tree_add_7_25_groupi_n_1073, csa_tree_add_7_25_groupi_n_1074, csa_tree_add_7_25_groupi_n_1075;
  wire csa_tree_add_7_25_groupi_n_1076, csa_tree_add_7_25_groupi_n_1077, csa_tree_add_7_25_groupi_n_1078, csa_tree_add_7_25_groupi_n_1079, csa_tree_add_7_25_groupi_n_1080, csa_tree_add_7_25_groupi_n_1081, csa_tree_add_7_25_groupi_n_1082, csa_tree_add_7_25_groupi_n_1083;
  wire csa_tree_add_7_25_groupi_n_1084, csa_tree_add_7_25_groupi_n_1085, csa_tree_add_7_25_groupi_n_1086, csa_tree_add_7_25_groupi_n_1087, csa_tree_add_7_25_groupi_n_1088, csa_tree_add_7_25_groupi_n_1089, csa_tree_add_7_25_groupi_n_1090, csa_tree_add_7_25_groupi_n_1091;
  wire csa_tree_add_7_25_groupi_n_1092, csa_tree_add_7_25_groupi_n_1093, csa_tree_add_7_25_groupi_n_1094, csa_tree_add_7_25_groupi_n_1095, csa_tree_add_7_25_groupi_n_1096, csa_tree_add_7_25_groupi_n_1097, csa_tree_add_7_25_groupi_n_1098, csa_tree_add_7_25_groupi_n_1099;
  wire csa_tree_add_7_25_groupi_n_1100, csa_tree_add_7_25_groupi_n_1101, csa_tree_add_7_25_groupi_n_1102, csa_tree_add_7_25_groupi_n_1103, csa_tree_add_7_25_groupi_n_1104, csa_tree_add_7_25_groupi_n_1105, csa_tree_add_7_25_groupi_n_1106, csa_tree_add_7_25_groupi_n_1107;
  wire csa_tree_add_7_25_groupi_n_1108, csa_tree_add_7_25_groupi_n_1109, csa_tree_add_7_25_groupi_n_1110, csa_tree_add_7_25_groupi_n_1111, csa_tree_add_7_25_groupi_n_1112, csa_tree_add_7_25_groupi_n_1113, csa_tree_add_7_25_groupi_n_1114, csa_tree_add_7_25_groupi_n_1115;
  wire csa_tree_add_7_25_groupi_n_1116, csa_tree_add_7_25_groupi_n_1117, csa_tree_add_7_25_groupi_n_1118, csa_tree_add_7_25_groupi_n_1119, csa_tree_add_7_25_groupi_n_1120, csa_tree_add_7_25_groupi_n_1121, csa_tree_add_7_25_groupi_n_1122, csa_tree_add_7_25_groupi_n_1123;
  wire csa_tree_add_7_25_groupi_n_1124, csa_tree_add_7_25_groupi_n_1125, csa_tree_add_7_25_groupi_n_1126, csa_tree_add_7_25_groupi_n_1127, csa_tree_add_7_25_groupi_n_1128, csa_tree_add_7_25_groupi_n_1129, csa_tree_add_7_25_groupi_n_1130, csa_tree_add_7_25_groupi_n_1131;
  wire csa_tree_add_7_25_groupi_n_1132, csa_tree_add_7_25_groupi_n_1133, csa_tree_add_7_25_groupi_n_1134, csa_tree_add_7_25_groupi_n_1135, csa_tree_add_7_25_groupi_n_1136, csa_tree_add_7_25_groupi_n_1137, csa_tree_add_7_25_groupi_n_1138, csa_tree_add_7_25_groupi_n_1139;
  wire csa_tree_add_7_25_groupi_n_1140, csa_tree_add_7_25_groupi_n_1141, csa_tree_add_7_25_groupi_n_1142, csa_tree_add_7_25_groupi_n_1143, csa_tree_add_7_25_groupi_n_1144, csa_tree_add_7_25_groupi_n_1145, csa_tree_add_7_25_groupi_n_1146, csa_tree_add_7_25_groupi_n_1147;
  wire csa_tree_add_7_25_groupi_n_1148, csa_tree_add_7_25_groupi_n_1149, csa_tree_add_7_25_groupi_n_1150, csa_tree_add_7_25_groupi_n_1151, csa_tree_add_7_25_groupi_n_1152, csa_tree_add_7_25_groupi_n_1153, csa_tree_add_7_25_groupi_n_1154, csa_tree_add_7_25_groupi_n_1155;
  wire csa_tree_add_7_25_groupi_n_1156, csa_tree_add_7_25_groupi_n_1157, csa_tree_add_7_25_groupi_n_1158, csa_tree_add_7_25_groupi_n_1159, csa_tree_add_7_25_groupi_n_1160, csa_tree_add_7_25_groupi_n_1161, csa_tree_add_7_25_groupi_n_1162, csa_tree_add_7_25_groupi_n_1163;
  wire csa_tree_add_7_25_groupi_n_1164, csa_tree_add_7_25_groupi_n_1165, csa_tree_add_7_25_groupi_n_1166, csa_tree_add_7_25_groupi_n_1167, csa_tree_add_7_25_groupi_n_1168, csa_tree_add_7_25_groupi_n_1169, csa_tree_add_7_25_groupi_n_1170, csa_tree_add_7_25_groupi_n_1171;
  wire csa_tree_add_7_25_groupi_n_1172, csa_tree_add_7_25_groupi_n_1173, csa_tree_add_7_25_groupi_n_1174, csa_tree_add_7_25_groupi_n_1175, csa_tree_add_7_25_groupi_n_1176, csa_tree_add_7_25_groupi_n_1177, csa_tree_add_7_25_groupi_n_1178, csa_tree_add_7_25_groupi_n_1179;
  wire csa_tree_add_7_25_groupi_n_1180, csa_tree_add_7_25_groupi_n_1181, csa_tree_add_7_25_groupi_n_1182, csa_tree_add_7_25_groupi_n_1183, csa_tree_add_7_25_groupi_n_1184, csa_tree_add_7_25_groupi_n_1185, csa_tree_add_7_25_groupi_n_1186, csa_tree_add_7_25_groupi_n_1187;
  wire csa_tree_add_7_25_groupi_n_1188, csa_tree_add_7_25_groupi_n_1189, csa_tree_add_7_25_groupi_n_1190, csa_tree_add_7_25_groupi_n_1191, csa_tree_add_7_25_groupi_n_1192, csa_tree_add_7_25_groupi_n_1193, csa_tree_add_7_25_groupi_n_1194, csa_tree_add_7_25_groupi_n_1195;
  wire csa_tree_add_7_25_groupi_n_1196, csa_tree_add_7_25_groupi_n_1197, csa_tree_add_7_25_groupi_n_1198, csa_tree_add_7_25_groupi_n_1199, csa_tree_add_7_25_groupi_n_1200, csa_tree_add_7_25_groupi_n_1201, csa_tree_add_7_25_groupi_n_1202, csa_tree_add_7_25_groupi_n_1203;
  wire csa_tree_add_7_25_groupi_n_1204, csa_tree_add_7_25_groupi_n_1205, csa_tree_add_7_25_groupi_n_1206, csa_tree_add_7_25_groupi_n_1207, csa_tree_add_7_25_groupi_n_1208, csa_tree_add_7_25_groupi_n_1209, csa_tree_add_7_25_groupi_n_1210, csa_tree_add_7_25_groupi_n_1211;
  wire csa_tree_add_7_25_groupi_n_1212, csa_tree_add_7_25_groupi_n_1213, csa_tree_add_7_25_groupi_n_1214, csa_tree_add_7_25_groupi_n_1215, csa_tree_add_7_25_groupi_n_1216, csa_tree_add_7_25_groupi_n_1217, csa_tree_add_7_25_groupi_n_1218, csa_tree_add_7_25_groupi_n_1219;
  wire csa_tree_add_7_25_groupi_n_1220, csa_tree_add_7_25_groupi_n_1221, csa_tree_add_7_25_groupi_n_1222, csa_tree_add_7_25_groupi_n_1223, csa_tree_add_7_25_groupi_n_1224, csa_tree_add_7_25_groupi_n_1225, csa_tree_add_7_25_groupi_n_1226, csa_tree_add_7_25_groupi_n_1227;
  wire csa_tree_add_7_25_groupi_n_1228, csa_tree_add_7_25_groupi_n_1229, csa_tree_add_7_25_groupi_n_1230, csa_tree_add_7_25_groupi_n_1231, csa_tree_add_7_25_groupi_n_1232, csa_tree_add_7_25_groupi_n_1233, csa_tree_add_7_25_groupi_n_1234, csa_tree_add_7_25_groupi_n_1235;
  wire csa_tree_add_7_25_groupi_n_1236, csa_tree_add_7_25_groupi_n_1237, csa_tree_add_7_25_groupi_n_1238, csa_tree_add_7_25_groupi_n_1239, csa_tree_add_7_25_groupi_n_1240, csa_tree_add_7_25_groupi_n_1241, csa_tree_add_7_25_groupi_n_1242, csa_tree_add_7_25_groupi_n_1243;
  wire csa_tree_add_7_25_groupi_n_1244, csa_tree_add_7_25_groupi_n_1245, csa_tree_add_7_25_groupi_n_1246, csa_tree_add_7_25_groupi_n_1247, csa_tree_add_7_25_groupi_n_1248, csa_tree_add_7_25_groupi_n_1249, csa_tree_add_7_25_groupi_n_1250, csa_tree_add_7_25_groupi_n_1251;
  wire csa_tree_add_7_25_groupi_n_1252, csa_tree_add_7_25_groupi_n_1253, csa_tree_add_7_25_groupi_n_1254, csa_tree_add_7_25_groupi_n_1255, csa_tree_add_7_25_groupi_n_1256, csa_tree_add_7_25_groupi_n_1257, csa_tree_add_7_25_groupi_n_1258, csa_tree_add_7_25_groupi_n_1259;
  wire csa_tree_add_7_25_groupi_n_1260, csa_tree_add_7_25_groupi_n_1261, csa_tree_add_7_25_groupi_n_1262, csa_tree_add_7_25_groupi_n_1263, csa_tree_add_7_25_groupi_n_1264, csa_tree_add_7_25_groupi_n_1265, csa_tree_add_7_25_groupi_n_1266, csa_tree_add_7_25_groupi_n_1267;
  wire csa_tree_add_7_25_groupi_n_1268, csa_tree_add_7_25_groupi_n_1269, csa_tree_add_7_25_groupi_n_1270, csa_tree_add_7_25_groupi_n_1271, csa_tree_add_7_25_groupi_n_1272, csa_tree_add_7_25_groupi_n_1273, csa_tree_add_7_25_groupi_n_1274, csa_tree_add_7_25_groupi_n_1275;
  wire csa_tree_add_7_25_groupi_n_1276, csa_tree_add_7_25_groupi_n_1277, csa_tree_add_7_25_groupi_n_1278, csa_tree_add_7_25_groupi_n_1279, csa_tree_add_7_25_groupi_n_1280, csa_tree_add_7_25_groupi_n_1281, csa_tree_add_7_25_groupi_n_1282, csa_tree_add_7_25_groupi_n_1283;
  wire csa_tree_add_7_25_groupi_n_1284, csa_tree_add_7_25_groupi_n_1285, csa_tree_add_7_25_groupi_n_1286, csa_tree_add_7_25_groupi_n_1287, csa_tree_add_7_25_groupi_n_1288, csa_tree_add_7_25_groupi_n_1289, csa_tree_add_7_25_groupi_n_1290, csa_tree_add_7_25_groupi_n_1291;
  wire csa_tree_add_7_25_groupi_n_1292, csa_tree_add_7_25_groupi_n_1293, csa_tree_add_7_25_groupi_n_1294, csa_tree_add_7_25_groupi_n_1295, csa_tree_add_7_25_groupi_n_1296, csa_tree_add_7_25_groupi_n_1297, csa_tree_add_7_25_groupi_n_1298, csa_tree_add_7_25_groupi_n_1299;
  wire csa_tree_add_7_25_groupi_n_1300, csa_tree_add_7_25_groupi_n_1301, csa_tree_add_7_25_groupi_n_1302, csa_tree_add_7_25_groupi_n_1303, csa_tree_add_7_25_groupi_n_1304, csa_tree_add_7_25_groupi_n_1305, csa_tree_add_7_25_groupi_n_1306, csa_tree_add_7_25_groupi_n_1307;
  wire csa_tree_add_7_25_groupi_n_1308, csa_tree_add_7_25_groupi_n_1309, csa_tree_add_7_25_groupi_n_1310, csa_tree_add_7_25_groupi_n_1311, csa_tree_add_7_25_groupi_n_1312, csa_tree_add_7_25_groupi_n_1313, csa_tree_add_7_25_groupi_n_1314, csa_tree_add_7_25_groupi_n_1315;
  wire csa_tree_add_7_25_groupi_n_1316, csa_tree_add_7_25_groupi_n_1317, csa_tree_add_7_25_groupi_n_1318, csa_tree_add_7_25_groupi_n_1319, csa_tree_add_7_25_groupi_n_1320, csa_tree_add_7_25_groupi_n_1321, csa_tree_add_7_25_groupi_n_1322, csa_tree_add_7_25_groupi_n_1323;
  wire csa_tree_add_7_25_groupi_n_1324, csa_tree_add_7_25_groupi_n_1325, csa_tree_add_7_25_groupi_n_1326, csa_tree_add_7_25_groupi_n_1327, csa_tree_add_7_25_groupi_n_1328, csa_tree_add_7_25_groupi_n_1329, csa_tree_add_7_25_groupi_n_1330, csa_tree_add_7_25_groupi_n_1331;
  wire csa_tree_add_7_25_groupi_n_1332, csa_tree_add_7_25_groupi_n_1333, csa_tree_add_7_25_groupi_n_1334, csa_tree_add_7_25_groupi_n_1335, csa_tree_add_7_25_groupi_n_1336, csa_tree_add_7_25_groupi_n_1337, csa_tree_add_7_25_groupi_n_1338, csa_tree_add_7_25_groupi_n_1339;
  wire csa_tree_add_7_25_groupi_n_1340, csa_tree_add_7_25_groupi_n_1341, csa_tree_add_7_25_groupi_n_1342, csa_tree_add_7_25_groupi_n_1343, csa_tree_add_7_25_groupi_n_1344, csa_tree_add_7_25_groupi_n_1345, csa_tree_add_7_25_groupi_n_1346, csa_tree_add_7_25_groupi_n_1347;
  wire csa_tree_add_7_25_groupi_n_1348, csa_tree_add_7_25_groupi_n_1349, csa_tree_add_7_25_groupi_n_1350, csa_tree_add_7_25_groupi_n_1351, csa_tree_add_7_25_groupi_n_1352, csa_tree_add_7_25_groupi_n_1353, csa_tree_add_7_25_groupi_n_1354, csa_tree_add_7_25_groupi_n_1355;
  wire csa_tree_add_7_25_groupi_n_1356, csa_tree_add_7_25_groupi_n_1357, csa_tree_add_7_25_groupi_n_1358, csa_tree_add_7_25_groupi_n_1359, csa_tree_add_7_25_groupi_n_1360, csa_tree_add_7_25_groupi_n_1361, csa_tree_add_7_25_groupi_n_1362, csa_tree_add_7_25_groupi_n_1363;
  wire csa_tree_add_7_25_groupi_n_1364, csa_tree_add_7_25_groupi_n_1365, csa_tree_add_7_25_groupi_n_1366, csa_tree_add_7_25_groupi_n_1367, csa_tree_add_7_25_groupi_n_1368, csa_tree_add_7_25_groupi_n_1369, csa_tree_add_7_25_groupi_n_1370, csa_tree_add_7_25_groupi_n_1371;
  wire csa_tree_add_7_25_groupi_n_1372, csa_tree_add_7_25_groupi_n_1373, csa_tree_add_7_25_groupi_n_1374, csa_tree_add_7_25_groupi_n_1375, csa_tree_add_7_25_groupi_n_1376, csa_tree_add_7_25_groupi_n_1377, csa_tree_add_7_25_groupi_n_1378, csa_tree_add_7_25_groupi_n_1379;
  wire csa_tree_add_7_25_groupi_n_1380, csa_tree_add_7_25_groupi_n_1381, csa_tree_add_7_25_groupi_n_1382, csa_tree_add_7_25_groupi_n_1383, csa_tree_add_7_25_groupi_n_1384, csa_tree_add_7_25_groupi_n_1385, csa_tree_add_7_25_groupi_n_1386, csa_tree_add_7_25_groupi_n_1387;
  wire csa_tree_add_7_25_groupi_n_1388, csa_tree_add_7_25_groupi_n_1389, csa_tree_add_7_25_groupi_n_1390, csa_tree_add_7_25_groupi_n_1391, csa_tree_add_7_25_groupi_n_1392, csa_tree_add_7_25_groupi_n_1393, csa_tree_add_7_25_groupi_n_1394, csa_tree_add_7_25_groupi_n_1395;
  wire csa_tree_add_7_25_groupi_n_1396, csa_tree_add_7_25_groupi_n_1397, csa_tree_add_7_25_groupi_n_1398, csa_tree_add_7_25_groupi_n_1399, csa_tree_add_7_25_groupi_n_1400, csa_tree_add_7_25_groupi_n_1401, csa_tree_add_7_25_groupi_n_1402, csa_tree_add_7_25_groupi_n_1403;
  wire csa_tree_add_7_25_groupi_n_1404, csa_tree_add_7_25_groupi_n_1405, csa_tree_add_7_25_groupi_n_1406, csa_tree_add_7_25_groupi_n_1407, csa_tree_add_7_25_groupi_n_1408, csa_tree_add_7_25_groupi_n_1409, csa_tree_add_7_25_groupi_n_1410, csa_tree_add_7_25_groupi_n_1411;
  wire csa_tree_add_7_25_groupi_n_1412, csa_tree_add_7_25_groupi_n_1413, csa_tree_add_7_25_groupi_n_1414, csa_tree_add_7_25_groupi_n_1415, csa_tree_add_7_25_groupi_n_1416, csa_tree_add_7_25_groupi_n_1417, csa_tree_add_7_25_groupi_n_1418, csa_tree_add_7_25_groupi_n_1419;
  wire csa_tree_add_7_25_groupi_n_1420, csa_tree_add_7_25_groupi_n_1421, csa_tree_add_7_25_groupi_n_1422, csa_tree_add_7_25_groupi_n_1423, csa_tree_add_7_25_groupi_n_1424, csa_tree_add_7_25_groupi_n_1425, csa_tree_add_7_25_groupi_n_1426, csa_tree_add_7_25_groupi_n_1427;
  wire csa_tree_add_7_25_groupi_n_1428, csa_tree_add_7_25_groupi_n_1429, csa_tree_add_7_25_groupi_n_1430, csa_tree_add_7_25_groupi_n_1431, csa_tree_add_7_25_groupi_n_1432, csa_tree_add_7_25_groupi_n_1433, csa_tree_add_7_25_groupi_n_1434, csa_tree_add_7_25_groupi_n_1435;
  wire csa_tree_add_7_25_groupi_n_1436, csa_tree_add_7_25_groupi_n_1437, csa_tree_add_7_25_groupi_n_1438, csa_tree_add_7_25_groupi_n_1439, csa_tree_add_7_25_groupi_n_1440, csa_tree_add_7_25_groupi_n_1441, csa_tree_add_7_25_groupi_n_1442, csa_tree_add_7_25_groupi_n_1443;
  wire csa_tree_add_7_25_groupi_n_1444, csa_tree_add_7_25_groupi_n_1445, csa_tree_add_7_25_groupi_n_1446, csa_tree_add_7_25_groupi_n_1447, csa_tree_add_7_25_groupi_n_1448, csa_tree_add_7_25_groupi_n_1449, csa_tree_add_7_25_groupi_n_1450, csa_tree_add_7_25_groupi_n_1451;
  wire csa_tree_add_7_25_groupi_n_1452, csa_tree_add_7_25_groupi_n_1453, csa_tree_add_7_25_groupi_n_1454, csa_tree_add_7_25_groupi_n_1455, csa_tree_add_7_25_groupi_n_1456, csa_tree_add_7_25_groupi_n_1457, csa_tree_add_7_25_groupi_n_1458, csa_tree_add_7_25_groupi_n_1459;
  wire csa_tree_add_7_25_groupi_n_1460, csa_tree_add_7_25_groupi_n_1461, csa_tree_add_7_25_groupi_n_1462, csa_tree_add_7_25_groupi_n_1463, csa_tree_add_7_25_groupi_n_1464, csa_tree_add_7_25_groupi_n_1465, csa_tree_add_7_25_groupi_n_1466, csa_tree_add_7_25_groupi_n_1467;
  wire csa_tree_add_7_25_groupi_n_1468, csa_tree_add_7_25_groupi_n_1469, csa_tree_add_7_25_groupi_n_1470, csa_tree_add_7_25_groupi_n_1471, csa_tree_add_7_25_groupi_n_1472, csa_tree_add_7_25_groupi_n_1473, csa_tree_add_7_25_groupi_n_1474, csa_tree_add_7_25_groupi_n_1475;
  wire csa_tree_add_7_25_groupi_n_1476, csa_tree_add_7_25_groupi_n_1477, csa_tree_add_7_25_groupi_n_1478, csa_tree_add_7_25_groupi_n_1479, csa_tree_add_7_25_groupi_n_1480, csa_tree_add_7_25_groupi_n_1481, csa_tree_add_7_25_groupi_n_1482, csa_tree_add_7_25_groupi_n_1483;
  wire csa_tree_add_7_25_groupi_n_1484, csa_tree_add_7_25_groupi_n_1485, csa_tree_add_7_25_groupi_n_1486, csa_tree_add_7_25_groupi_n_1487, csa_tree_add_7_25_groupi_n_1488, csa_tree_add_7_25_groupi_n_1489, csa_tree_add_7_25_groupi_n_1490, csa_tree_add_7_25_groupi_n_1491;
  wire csa_tree_add_7_25_groupi_n_1492, csa_tree_add_7_25_groupi_n_1493, csa_tree_add_7_25_groupi_n_1494, csa_tree_add_7_25_groupi_n_1495, csa_tree_add_7_25_groupi_n_1496, csa_tree_add_7_25_groupi_n_1497, csa_tree_add_7_25_groupi_n_1498, csa_tree_add_7_25_groupi_n_1499;
  wire csa_tree_add_7_25_groupi_n_1500, csa_tree_add_7_25_groupi_n_1501, csa_tree_add_7_25_groupi_n_1502, csa_tree_add_7_25_groupi_n_1503, csa_tree_add_7_25_groupi_n_1504, csa_tree_add_7_25_groupi_n_1505, csa_tree_add_7_25_groupi_n_1506, csa_tree_add_7_25_groupi_n_1507;
  wire csa_tree_add_7_25_groupi_n_1508, csa_tree_add_7_25_groupi_n_1509, csa_tree_add_7_25_groupi_n_1510, csa_tree_add_7_25_groupi_n_1511, csa_tree_add_7_25_groupi_n_1512, csa_tree_add_7_25_groupi_n_1513, csa_tree_add_7_25_groupi_n_1514, csa_tree_add_7_25_groupi_n_1515;
  wire csa_tree_add_7_25_groupi_n_1516, csa_tree_add_7_25_groupi_n_1517, csa_tree_add_7_25_groupi_n_1518, csa_tree_add_7_25_groupi_n_1519, csa_tree_add_7_25_groupi_n_1520, csa_tree_add_7_25_groupi_n_1521, csa_tree_add_7_25_groupi_n_1522, csa_tree_add_7_25_groupi_n_1523;
  wire csa_tree_add_7_25_groupi_n_1524, csa_tree_add_7_25_groupi_n_1525, csa_tree_add_7_25_groupi_n_1526, csa_tree_add_7_25_groupi_n_1527, csa_tree_add_7_25_groupi_n_1528, csa_tree_add_7_25_groupi_n_1529, csa_tree_add_7_25_groupi_n_1530, csa_tree_add_7_25_groupi_n_1531;
  wire csa_tree_add_7_25_groupi_n_1532, csa_tree_add_7_25_groupi_n_1533, csa_tree_add_7_25_groupi_n_1534, csa_tree_add_7_25_groupi_n_1535, csa_tree_add_7_25_groupi_n_1536, csa_tree_add_7_25_groupi_n_1537, csa_tree_add_7_25_groupi_n_1538, csa_tree_add_7_25_groupi_n_1539;
  wire csa_tree_add_7_25_groupi_n_1540, csa_tree_add_7_25_groupi_n_1541, csa_tree_add_7_25_groupi_n_1542, csa_tree_add_7_25_groupi_n_1543, csa_tree_add_7_25_groupi_n_1544, csa_tree_add_7_25_groupi_n_1545, csa_tree_add_7_25_groupi_n_1546, csa_tree_add_7_25_groupi_n_1547;
  wire csa_tree_add_7_25_groupi_n_1548, csa_tree_add_7_25_groupi_n_1549, csa_tree_add_7_25_groupi_n_1550, csa_tree_add_7_25_groupi_n_1551, csa_tree_add_7_25_groupi_n_1552, csa_tree_add_7_25_groupi_n_1553, csa_tree_add_7_25_groupi_n_1554, csa_tree_add_7_25_groupi_n_1555;
  wire csa_tree_add_7_25_groupi_n_1556, csa_tree_add_7_25_groupi_n_1557, csa_tree_add_7_25_groupi_n_1558, csa_tree_add_7_25_groupi_n_1559, csa_tree_add_7_25_groupi_n_1560, csa_tree_add_7_25_groupi_n_1561, csa_tree_add_7_25_groupi_n_1562, csa_tree_add_7_25_groupi_n_1563;
  wire csa_tree_add_7_25_groupi_n_1564, csa_tree_add_7_25_groupi_n_1565, csa_tree_add_7_25_groupi_n_1566, csa_tree_add_7_25_groupi_n_1567, csa_tree_add_7_25_groupi_n_1568, csa_tree_add_7_25_groupi_n_1569, csa_tree_add_7_25_groupi_n_1570, csa_tree_add_7_25_groupi_n_1571;
  wire csa_tree_add_7_25_groupi_n_1572, csa_tree_add_7_25_groupi_n_1573, csa_tree_add_7_25_groupi_n_1574, csa_tree_add_7_25_groupi_n_1575, csa_tree_add_7_25_groupi_n_1576, csa_tree_add_7_25_groupi_n_1577, csa_tree_add_7_25_groupi_n_1578, csa_tree_add_7_25_groupi_n_1579;
  wire csa_tree_add_7_25_groupi_n_1580, csa_tree_add_7_25_groupi_n_1581, csa_tree_add_7_25_groupi_n_1582, csa_tree_add_7_25_groupi_n_1583, csa_tree_add_7_25_groupi_n_1584, csa_tree_add_7_25_groupi_n_1585, csa_tree_add_7_25_groupi_n_1586, csa_tree_add_7_25_groupi_n_1587;
  wire csa_tree_add_7_25_groupi_n_1588, csa_tree_add_7_25_groupi_n_1589, csa_tree_add_7_25_groupi_n_1590, csa_tree_add_7_25_groupi_n_1591, csa_tree_add_7_25_groupi_n_1592, csa_tree_add_7_25_groupi_n_1593, csa_tree_add_7_25_groupi_n_1594, csa_tree_add_7_25_groupi_n_1595;
  wire csa_tree_add_7_25_groupi_n_1596, csa_tree_add_7_25_groupi_n_1597, csa_tree_add_7_25_groupi_n_1598, csa_tree_add_7_25_groupi_n_1599, csa_tree_add_7_25_groupi_n_1600, csa_tree_add_7_25_groupi_n_1601, csa_tree_add_7_25_groupi_n_1602, csa_tree_add_7_25_groupi_n_1603;
  wire csa_tree_add_7_25_groupi_n_1604, csa_tree_add_7_25_groupi_n_1605, csa_tree_add_7_25_groupi_n_1606, csa_tree_add_7_25_groupi_n_1607, csa_tree_add_7_25_groupi_n_1608, csa_tree_add_7_25_groupi_n_1609, csa_tree_add_7_25_groupi_n_1610, csa_tree_add_7_25_groupi_n_1611;
  wire csa_tree_add_7_25_groupi_n_1612, csa_tree_add_7_25_groupi_n_1613, csa_tree_add_7_25_groupi_n_1614, csa_tree_add_7_25_groupi_n_1615, csa_tree_add_7_25_groupi_n_1616, csa_tree_add_7_25_groupi_n_1617, csa_tree_add_7_25_groupi_n_1618, csa_tree_add_7_25_groupi_n_1619;
  wire csa_tree_add_7_25_groupi_n_1620, csa_tree_add_7_25_groupi_n_1621, csa_tree_add_7_25_groupi_n_1622, csa_tree_add_7_25_groupi_n_1623, csa_tree_add_7_25_groupi_n_1624, csa_tree_add_7_25_groupi_n_1625, csa_tree_add_7_25_groupi_n_1626, csa_tree_add_7_25_groupi_n_1627;
  wire csa_tree_add_7_25_groupi_n_1628, csa_tree_add_7_25_groupi_n_1629, csa_tree_add_7_25_groupi_n_1630, csa_tree_add_7_25_groupi_n_1631, csa_tree_add_7_25_groupi_n_1632, csa_tree_add_7_25_groupi_n_1633, csa_tree_add_7_25_groupi_n_1634, csa_tree_add_7_25_groupi_n_1635;
  wire csa_tree_add_7_25_groupi_n_1636, csa_tree_add_7_25_groupi_n_1637, csa_tree_add_7_25_groupi_n_1638, csa_tree_add_7_25_groupi_n_1639, csa_tree_add_7_25_groupi_n_1640, csa_tree_add_7_25_groupi_n_1641, csa_tree_add_7_25_groupi_n_1642, csa_tree_add_7_25_groupi_n_1643;
  wire csa_tree_add_7_25_groupi_n_1644, csa_tree_add_7_25_groupi_n_1645, csa_tree_add_7_25_groupi_n_1646, csa_tree_add_7_25_groupi_n_1647, csa_tree_add_7_25_groupi_n_1648, csa_tree_add_7_25_groupi_n_1649, csa_tree_add_7_25_groupi_n_1650, csa_tree_add_7_25_groupi_n_1651;
  wire csa_tree_add_7_25_groupi_n_1652, csa_tree_add_7_25_groupi_n_1653, csa_tree_add_7_25_groupi_n_1654, csa_tree_add_7_25_groupi_n_1655, csa_tree_add_7_25_groupi_n_1656, csa_tree_add_7_25_groupi_n_1657, csa_tree_add_7_25_groupi_n_1658, csa_tree_add_7_25_groupi_n_1659;
  wire csa_tree_add_7_25_groupi_n_1660, csa_tree_add_7_25_groupi_n_1661, csa_tree_add_7_25_groupi_n_1662, csa_tree_add_7_25_groupi_n_1663, csa_tree_add_7_25_groupi_n_1664, csa_tree_add_7_25_groupi_n_1665, csa_tree_add_7_25_groupi_n_1666, csa_tree_add_7_25_groupi_n_1667;
  wire csa_tree_add_7_25_groupi_n_1668, csa_tree_add_7_25_groupi_n_1669, csa_tree_add_7_25_groupi_n_1670, csa_tree_add_7_25_groupi_n_1671, csa_tree_add_7_25_groupi_n_1672, csa_tree_add_7_25_groupi_n_1673, csa_tree_add_7_25_groupi_n_1674, csa_tree_add_7_25_groupi_n_1675;
  wire csa_tree_add_7_25_groupi_n_1676, csa_tree_add_7_25_groupi_n_1677, csa_tree_add_7_25_groupi_n_1678, csa_tree_add_7_25_groupi_n_1679, csa_tree_add_7_25_groupi_n_1680, csa_tree_add_7_25_groupi_n_1681, csa_tree_add_7_25_groupi_n_1682, csa_tree_add_7_25_groupi_n_1683;
  wire csa_tree_add_7_25_groupi_n_1684, csa_tree_add_7_25_groupi_n_1685, csa_tree_add_7_25_groupi_n_1686, csa_tree_add_7_25_groupi_n_1687, csa_tree_add_7_25_groupi_n_1688, csa_tree_add_7_25_groupi_n_1689, csa_tree_add_7_25_groupi_n_1690, csa_tree_add_7_25_groupi_n_1691;
  wire csa_tree_add_7_25_groupi_n_1692, csa_tree_add_7_25_groupi_n_1693, csa_tree_add_7_25_groupi_n_1694, csa_tree_add_7_25_groupi_n_1695, csa_tree_add_7_25_groupi_n_1696, csa_tree_add_7_25_groupi_n_1697, csa_tree_add_7_25_groupi_n_1698, csa_tree_add_7_25_groupi_n_1699;
  wire csa_tree_add_7_25_groupi_n_1700, csa_tree_add_7_25_groupi_n_1701, csa_tree_add_7_25_groupi_n_1702, csa_tree_add_7_25_groupi_n_1703, csa_tree_add_7_25_groupi_n_1704, csa_tree_add_7_25_groupi_n_1705, csa_tree_add_7_25_groupi_n_1706, csa_tree_add_7_25_groupi_n_1707;
  wire csa_tree_add_7_25_groupi_n_1708, csa_tree_add_7_25_groupi_n_1709, csa_tree_add_7_25_groupi_n_1710, csa_tree_add_7_25_groupi_n_1711, csa_tree_add_7_25_groupi_n_1712, csa_tree_add_7_25_groupi_n_1713, csa_tree_add_7_25_groupi_n_1714, csa_tree_add_7_25_groupi_n_1715;
  wire csa_tree_add_7_25_groupi_n_1716, csa_tree_add_7_25_groupi_n_1717, csa_tree_add_7_25_groupi_n_1718, csa_tree_add_7_25_groupi_n_1719, csa_tree_add_7_25_groupi_n_1720, csa_tree_add_7_25_groupi_n_1721, csa_tree_add_7_25_groupi_n_1722, csa_tree_add_7_25_groupi_n_1723;
  wire csa_tree_add_7_25_groupi_n_1724, csa_tree_add_7_25_groupi_n_1725, csa_tree_add_7_25_groupi_n_1726, csa_tree_add_7_25_groupi_n_1727, csa_tree_add_7_25_groupi_n_1728, csa_tree_add_7_25_groupi_n_1729, csa_tree_add_7_25_groupi_n_1730, csa_tree_add_7_25_groupi_n_1731;
  wire csa_tree_add_7_25_groupi_n_1732, csa_tree_add_7_25_groupi_n_1733, csa_tree_add_7_25_groupi_n_1734, csa_tree_add_7_25_groupi_n_1735, csa_tree_add_7_25_groupi_n_1736, csa_tree_add_7_25_groupi_n_1737, csa_tree_add_7_25_groupi_n_1738, csa_tree_add_7_25_groupi_n_1739;
  wire csa_tree_add_7_25_groupi_n_1740, csa_tree_add_7_25_groupi_n_1741, csa_tree_add_7_25_groupi_n_1742, csa_tree_add_7_25_groupi_n_1743, csa_tree_add_7_25_groupi_n_1744, csa_tree_add_7_25_groupi_n_1745, csa_tree_add_7_25_groupi_n_1746, csa_tree_add_7_25_groupi_n_1747;
  wire csa_tree_add_7_25_groupi_n_1748, csa_tree_add_7_25_groupi_n_1749, csa_tree_add_7_25_groupi_n_1750, csa_tree_add_7_25_groupi_n_1751, csa_tree_add_7_25_groupi_n_1752, csa_tree_add_7_25_groupi_n_1753, csa_tree_add_7_25_groupi_n_1754, csa_tree_add_7_25_groupi_n_1755;
  wire csa_tree_add_7_25_groupi_n_1756, csa_tree_add_7_25_groupi_n_1757, csa_tree_add_7_25_groupi_n_1758, csa_tree_add_7_25_groupi_n_1759, csa_tree_add_7_25_groupi_n_1760, csa_tree_add_7_25_groupi_n_1761, csa_tree_add_7_25_groupi_n_1762, csa_tree_add_7_25_groupi_n_1763;
  wire csa_tree_add_7_25_groupi_n_1764, csa_tree_add_7_25_groupi_n_1765, csa_tree_add_7_25_groupi_n_1766, csa_tree_add_7_25_groupi_n_1767, csa_tree_add_7_25_groupi_n_1768, csa_tree_add_7_25_groupi_n_1769, csa_tree_add_7_25_groupi_n_1770, csa_tree_add_7_25_groupi_n_1771;
  wire csa_tree_add_7_25_groupi_n_1772, csa_tree_add_7_25_groupi_n_1773, csa_tree_add_7_25_groupi_n_1774, csa_tree_add_7_25_groupi_n_1775, csa_tree_add_7_25_groupi_n_1776, csa_tree_add_7_25_groupi_n_1777, csa_tree_add_7_25_groupi_n_1778, csa_tree_add_7_25_groupi_n_1779;
  wire csa_tree_add_7_25_groupi_n_1780, csa_tree_add_7_25_groupi_n_1781, csa_tree_add_7_25_groupi_n_1782, csa_tree_add_7_25_groupi_n_1783, csa_tree_add_7_25_groupi_n_1784, csa_tree_add_7_25_groupi_n_1785, csa_tree_add_7_25_groupi_n_1786, csa_tree_add_7_25_groupi_n_1787;
  wire csa_tree_add_7_25_groupi_n_1788, csa_tree_add_7_25_groupi_n_1789, csa_tree_add_7_25_groupi_n_1790, csa_tree_add_7_25_groupi_n_1791, csa_tree_add_7_25_groupi_n_1792, csa_tree_add_7_25_groupi_n_1793, csa_tree_add_7_25_groupi_n_1794, csa_tree_add_7_25_groupi_n_1795;
  wire csa_tree_add_7_25_groupi_n_1796, csa_tree_add_7_25_groupi_n_1797, csa_tree_add_7_25_groupi_n_1798, csa_tree_add_7_25_groupi_n_1799, csa_tree_add_7_25_groupi_n_1800, csa_tree_add_7_25_groupi_n_1801, csa_tree_add_7_25_groupi_n_1802, csa_tree_add_7_25_groupi_n_1803;
  wire csa_tree_add_7_25_groupi_n_1804, csa_tree_add_7_25_groupi_n_1805, csa_tree_add_7_25_groupi_n_1806, csa_tree_add_7_25_groupi_n_1807, csa_tree_add_7_25_groupi_n_1808, csa_tree_add_7_25_groupi_n_1809, csa_tree_add_7_25_groupi_n_1810, csa_tree_add_7_25_groupi_n_1811;
  wire csa_tree_add_7_25_groupi_n_1812, csa_tree_add_7_25_groupi_n_1813, csa_tree_add_7_25_groupi_n_1814, csa_tree_add_7_25_groupi_n_1815, csa_tree_add_7_25_groupi_n_1816, csa_tree_add_7_25_groupi_n_1817, csa_tree_add_7_25_groupi_n_1818, csa_tree_add_7_25_groupi_n_1819;
  wire csa_tree_add_7_25_groupi_n_1820, csa_tree_add_7_25_groupi_n_1821, csa_tree_add_7_25_groupi_n_1822, csa_tree_add_7_25_groupi_n_1823, csa_tree_add_7_25_groupi_n_1824, csa_tree_add_7_25_groupi_n_1825, csa_tree_add_7_25_groupi_n_1826, csa_tree_add_7_25_groupi_n_1827;
  wire csa_tree_add_7_25_groupi_n_1828, csa_tree_add_7_25_groupi_n_1829, csa_tree_add_7_25_groupi_n_1830, csa_tree_add_7_25_groupi_n_1831, csa_tree_add_7_25_groupi_n_1832, csa_tree_add_7_25_groupi_n_1833, csa_tree_add_7_25_groupi_n_1834, csa_tree_add_7_25_groupi_n_1835;
  wire csa_tree_add_7_25_groupi_n_1836, csa_tree_add_7_25_groupi_n_1837, csa_tree_add_7_25_groupi_n_1838, csa_tree_add_7_25_groupi_n_1839, csa_tree_add_7_25_groupi_n_1840, csa_tree_add_7_25_groupi_n_1841, csa_tree_add_7_25_groupi_n_1842, csa_tree_add_7_25_groupi_n_1843;
  wire csa_tree_add_7_25_groupi_n_1844, csa_tree_add_7_25_groupi_n_1845, csa_tree_add_7_25_groupi_n_1846, csa_tree_add_7_25_groupi_n_1847, csa_tree_add_7_25_groupi_n_1848, csa_tree_add_7_25_groupi_n_1849, csa_tree_add_7_25_groupi_n_1850, csa_tree_add_7_25_groupi_n_1851;
  wire csa_tree_add_7_25_groupi_n_1852, csa_tree_add_7_25_groupi_n_1853, csa_tree_add_7_25_groupi_n_1854, csa_tree_add_7_25_groupi_n_1855, csa_tree_add_7_25_groupi_n_1856, csa_tree_add_7_25_groupi_n_1857, csa_tree_add_7_25_groupi_n_1858, csa_tree_add_7_25_groupi_n_1859;
  wire csa_tree_add_7_25_groupi_n_1860, csa_tree_add_7_25_groupi_n_1861, csa_tree_add_7_25_groupi_n_1862, csa_tree_add_7_25_groupi_n_1863, csa_tree_add_7_25_groupi_n_1864, csa_tree_add_7_25_groupi_n_1865, csa_tree_add_7_25_groupi_n_1866, csa_tree_add_7_25_groupi_n_1867;
  wire csa_tree_add_7_25_groupi_n_1868, csa_tree_add_7_25_groupi_n_1869, csa_tree_add_7_25_groupi_n_1870, csa_tree_add_7_25_groupi_n_1871, csa_tree_add_7_25_groupi_n_1872, csa_tree_add_7_25_groupi_n_1873, csa_tree_add_7_25_groupi_n_1874, csa_tree_add_7_25_groupi_n_1875;
  wire csa_tree_add_7_25_groupi_n_1876, csa_tree_add_7_25_groupi_n_1877, csa_tree_add_7_25_groupi_n_1878, csa_tree_add_7_25_groupi_n_1879, csa_tree_add_7_25_groupi_n_1880, csa_tree_add_7_25_groupi_n_1881, csa_tree_add_7_25_groupi_n_1882, csa_tree_add_7_25_groupi_n_1883;
  wire csa_tree_add_7_25_groupi_n_1884, csa_tree_add_7_25_groupi_n_1885, csa_tree_add_7_25_groupi_n_1886, csa_tree_add_7_25_groupi_n_1887, csa_tree_add_7_25_groupi_n_1888, csa_tree_add_7_25_groupi_n_1889, csa_tree_add_7_25_groupi_n_1890, csa_tree_add_7_25_groupi_n_1891;
  wire csa_tree_add_7_25_groupi_n_1892, csa_tree_add_7_25_groupi_n_1893, csa_tree_add_7_25_groupi_n_1894, csa_tree_add_7_25_groupi_n_1895, csa_tree_add_7_25_groupi_n_1896, csa_tree_add_7_25_groupi_n_1897, csa_tree_add_7_25_groupi_n_1898, csa_tree_add_7_25_groupi_n_1899;
  wire csa_tree_add_7_25_groupi_n_1900, csa_tree_add_7_25_groupi_n_1901, csa_tree_add_7_25_groupi_n_1902, csa_tree_add_7_25_groupi_n_1903, csa_tree_add_7_25_groupi_n_1904, csa_tree_add_7_25_groupi_n_1905, csa_tree_add_7_25_groupi_n_1906, csa_tree_add_7_25_groupi_n_1907;
  wire csa_tree_add_7_25_groupi_n_1908, csa_tree_add_7_25_groupi_n_1909, csa_tree_add_7_25_groupi_n_1910, csa_tree_add_7_25_groupi_n_1911, csa_tree_add_7_25_groupi_n_1912, csa_tree_add_7_25_groupi_n_1913, csa_tree_add_7_25_groupi_n_1914, csa_tree_add_7_25_groupi_n_1915;
  wire csa_tree_add_7_25_groupi_n_1916, csa_tree_add_7_25_groupi_n_1917, csa_tree_add_7_25_groupi_n_1918, csa_tree_add_7_25_groupi_n_1919, csa_tree_add_7_25_groupi_n_1920, csa_tree_add_7_25_groupi_n_1921, csa_tree_add_7_25_groupi_n_1922, csa_tree_add_7_25_groupi_n_1923;
  wire csa_tree_add_7_25_groupi_n_1924, csa_tree_add_7_25_groupi_n_1925, csa_tree_add_7_25_groupi_n_1926, csa_tree_add_7_25_groupi_n_1927, csa_tree_add_7_25_groupi_n_1928, csa_tree_add_7_25_groupi_n_1929, csa_tree_add_7_25_groupi_n_1930, csa_tree_add_7_25_groupi_n_1931;
  wire csa_tree_add_7_25_groupi_n_1932, csa_tree_add_7_25_groupi_n_1933, csa_tree_add_7_25_groupi_n_1934, csa_tree_add_7_25_groupi_n_1935, csa_tree_add_7_25_groupi_n_1936, csa_tree_add_7_25_groupi_n_1937, csa_tree_add_7_25_groupi_n_1938, csa_tree_add_7_25_groupi_n_1939;
  wire csa_tree_add_7_25_groupi_n_1940, csa_tree_add_7_25_groupi_n_1941, csa_tree_add_7_25_groupi_n_1942, csa_tree_add_7_25_groupi_n_1943, csa_tree_add_7_25_groupi_n_1944, csa_tree_add_7_25_groupi_n_1945, csa_tree_add_7_25_groupi_n_1946, csa_tree_add_7_25_groupi_n_1947;
  wire csa_tree_add_7_25_groupi_n_1948, csa_tree_add_7_25_groupi_n_1949, csa_tree_add_7_25_groupi_n_1950, csa_tree_add_7_25_groupi_n_1951, csa_tree_add_7_25_groupi_n_1952, csa_tree_add_7_25_groupi_n_1953, csa_tree_add_7_25_groupi_n_1954, csa_tree_add_7_25_groupi_n_1955;
  wire csa_tree_add_7_25_groupi_n_1956, csa_tree_add_7_25_groupi_n_1957, csa_tree_add_7_25_groupi_n_1958, csa_tree_add_7_25_groupi_n_1959, csa_tree_add_7_25_groupi_n_1960, csa_tree_add_7_25_groupi_n_1961, csa_tree_add_7_25_groupi_n_1962, csa_tree_add_7_25_groupi_n_1963;
  wire csa_tree_add_7_25_groupi_n_1964, csa_tree_add_7_25_groupi_n_1965, csa_tree_add_7_25_groupi_n_1966, csa_tree_add_7_25_groupi_n_1967, csa_tree_add_7_25_groupi_n_1968, csa_tree_add_7_25_groupi_n_1969, csa_tree_add_7_25_groupi_n_1970, csa_tree_add_7_25_groupi_n_1971;
  wire csa_tree_add_7_25_groupi_n_1972, csa_tree_add_7_25_groupi_n_1973, csa_tree_add_7_25_groupi_n_1974, csa_tree_add_7_25_groupi_n_1975, csa_tree_add_7_25_groupi_n_1976, csa_tree_add_7_25_groupi_n_1977, csa_tree_add_7_25_groupi_n_1978, csa_tree_add_7_25_groupi_n_1979;
  wire csa_tree_add_7_25_groupi_n_1980, csa_tree_add_7_25_groupi_n_1981, csa_tree_add_7_25_groupi_n_1982, csa_tree_add_7_25_groupi_n_1983, csa_tree_add_7_25_groupi_n_1984, csa_tree_add_7_25_groupi_n_1985, csa_tree_add_7_25_groupi_n_1986, csa_tree_add_7_25_groupi_n_1987;
  wire csa_tree_add_7_25_groupi_n_1988, csa_tree_add_7_25_groupi_n_1989, csa_tree_add_7_25_groupi_n_1990, csa_tree_add_7_25_groupi_n_1991, csa_tree_add_7_25_groupi_n_1992, csa_tree_add_7_25_groupi_n_1993, csa_tree_add_7_25_groupi_n_1994, csa_tree_add_7_25_groupi_n_1995;
  wire csa_tree_add_7_25_groupi_n_1996, csa_tree_add_7_25_groupi_n_1997, csa_tree_add_7_25_groupi_n_1998, csa_tree_add_7_25_groupi_n_1999, csa_tree_add_7_25_groupi_n_2000, csa_tree_add_7_25_groupi_n_2001, csa_tree_add_7_25_groupi_n_2002, csa_tree_add_7_25_groupi_n_2003;
  wire csa_tree_add_7_25_groupi_n_2004, csa_tree_add_7_25_groupi_n_2005, csa_tree_add_7_25_groupi_n_2006, csa_tree_add_7_25_groupi_n_2007, csa_tree_add_7_25_groupi_n_2008, csa_tree_add_7_25_groupi_n_2009, csa_tree_add_7_25_groupi_n_2010, csa_tree_add_7_25_groupi_n_2011;
  wire csa_tree_add_7_25_groupi_n_2012, csa_tree_add_7_25_groupi_n_2013, csa_tree_add_7_25_groupi_n_2014, csa_tree_add_7_25_groupi_n_2015, csa_tree_add_7_25_groupi_n_2016, csa_tree_add_7_25_groupi_n_2017, csa_tree_add_7_25_groupi_n_2018, csa_tree_add_7_25_groupi_n_2019;
  wire csa_tree_add_7_25_groupi_n_2020, csa_tree_add_7_25_groupi_n_2021, csa_tree_add_7_25_groupi_n_2022, csa_tree_add_7_25_groupi_n_2023, csa_tree_add_7_25_groupi_n_2024, csa_tree_add_7_25_groupi_n_2025, csa_tree_add_7_25_groupi_n_2026, csa_tree_add_7_25_groupi_n_2027;
  wire csa_tree_add_7_25_groupi_n_2028, csa_tree_add_7_25_groupi_n_2029, csa_tree_add_7_25_groupi_n_2030, csa_tree_add_7_25_groupi_n_2031, csa_tree_add_7_25_groupi_n_2032, csa_tree_add_7_25_groupi_n_2033, csa_tree_add_7_25_groupi_n_2034, csa_tree_add_7_25_groupi_n_2035;
  wire csa_tree_add_7_25_groupi_n_2036, csa_tree_add_7_25_groupi_n_2037, csa_tree_add_7_25_groupi_n_2038, csa_tree_add_7_25_groupi_n_2039, csa_tree_add_7_25_groupi_n_2040, csa_tree_add_7_25_groupi_n_2041, csa_tree_add_7_25_groupi_n_2042, csa_tree_add_7_25_groupi_n_2043;
  wire csa_tree_add_7_25_groupi_n_2044, csa_tree_add_7_25_groupi_n_2045, csa_tree_add_7_25_groupi_n_2046, csa_tree_add_7_25_groupi_n_2047, csa_tree_add_7_25_groupi_n_2048, csa_tree_add_7_25_groupi_n_2049, csa_tree_add_7_25_groupi_n_2050, csa_tree_add_7_25_groupi_n_2051;
  wire csa_tree_add_7_25_groupi_n_2052, csa_tree_add_7_25_groupi_n_2053, csa_tree_add_7_25_groupi_n_2054, csa_tree_add_7_25_groupi_n_2055, csa_tree_add_7_25_groupi_n_2056, csa_tree_add_7_25_groupi_n_2057, csa_tree_add_7_25_groupi_n_2058, csa_tree_add_7_25_groupi_n_2059;
  wire csa_tree_add_7_25_groupi_n_2060, csa_tree_add_7_25_groupi_n_2061, csa_tree_add_7_25_groupi_n_2062, csa_tree_add_7_25_groupi_n_2063, csa_tree_add_7_25_groupi_n_2064, csa_tree_add_7_25_groupi_n_2065, csa_tree_add_7_25_groupi_n_2066, csa_tree_add_7_25_groupi_n_2067;
  wire csa_tree_add_7_25_groupi_n_2068, csa_tree_add_7_25_groupi_n_2069, csa_tree_add_7_25_groupi_n_2070, csa_tree_add_7_25_groupi_n_2071, csa_tree_add_7_25_groupi_n_2072, csa_tree_add_7_25_groupi_n_2073, csa_tree_add_7_25_groupi_n_2074, csa_tree_add_7_25_groupi_n_2075;
  wire csa_tree_add_7_25_groupi_n_2076, csa_tree_add_7_25_groupi_n_2077, csa_tree_add_7_25_groupi_n_2078, csa_tree_add_7_25_groupi_n_2079, csa_tree_add_7_25_groupi_n_2080, csa_tree_add_7_25_groupi_n_2081, csa_tree_add_7_25_groupi_n_2082, csa_tree_add_7_25_groupi_n_2083;
  wire csa_tree_add_7_25_groupi_n_2084, csa_tree_add_7_25_groupi_n_2085, csa_tree_add_7_25_groupi_n_2086, csa_tree_add_7_25_groupi_n_2087, csa_tree_add_7_25_groupi_n_2088, csa_tree_add_7_25_groupi_n_2089, csa_tree_add_7_25_groupi_n_2090, csa_tree_add_7_25_groupi_n_2091;
  wire csa_tree_add_7_25_groupi_n_2092, csa_tree_add_7_25_groupi_n_2093, csa_tree_add_7_25_groupi_n_2094, csa_tree_add_7_25_groupi_n_2095, csa_tree_add_7_25_groupi_n_2096, csa_tree_add_7_25_groupi_n_2097, csa_tree_add_7_25_groupi_n_2098, csa_tree_add_7_25_groupi_n_2099;
  wire csa_tree_add_7_25_groupi_n_2100, csa_tree_add_7_25_groupi_n_2101, csa_tree_add_7_25_groupi_n_2102, csa_tree_add_7_25_groupi_n_2103, csa_tree_add_7_25_groupi_n_2104, csa_tree_add_7_25_groupi_n_2105, csa_tree_add_7_25_groupi_n_2106, csa_tree_add_7_25_groupi_n_2107;
  wire csa_tree_add_7_25_groupi_n_2108, csa_tree_add_7_25_groupi_n_2109, csa_tree_add_7_25_groupi_n_2110, csa_tree_add_7_25_groupi_n_2111, csa_tree_add_7_25_groupi_n_2112, csa_tree_add_7_25_groupi_n_2113, csa_tree_add_7_25_groupi_n_2114, csa_tree_add_7_25_groupi_n_2115;
  wire csa_tree_add_7_25_groupi_n_2116, csa_tree_add_7_25_groupi_n_2117, csa_tree_add_7_25_groupi_n_2118, csa_tree_add_7_25_groupi_n_2119, csa_tree_add_7_25_groupi_n_2120, csa_tree_add_7_25_groupi_n_2121, csa_tree_add_7_25_groupi_n_2122, csa_tree_add_7_25_groupi_n_2123;
  wire csa_tree_add_7_25_groupi_n_2124, csa_tree_add_7_25_groupi_n_2125, csa_tree_add_7_25_groupi_n_2126, csa_tree_add_7_25_groupi_n_2127, csa_tree_add_7_25_groupi_n_2128, csa_tree_add_7_25_groupi_n_2129, csa_tree_add_7_25_groupi_n_2130, csa_tree_add_7_25_groupi_n_2131;
  wire csa_tree_add_7_25_groupi_n_2132, csa_tree_add_7_25_groupi_n_2133, csa_tree_add_7_25_groupi_n_2134, csa_tree_add_7_25_groupi_n_2135, csa_tree_add_7_25_groupi_n_2136, csa_tree_add_7_25_groupi_n_2137, csa_tree_add_7_25_groupi_n_2138, csa_tree_add_7_25_groupi_n_2139;
  wire csa_tree_add_7_25_groupi_n_2140, csa_tree_add_7_25_groupi_n_2141, csa_tree_add_7_25_groupi_n_2142, csa_tree_add_7_25_groupi_n_2143, csa_tree_add_7_25_groupi_n_2144, csa_tree_add_7_25_groupi_n_2145, csa_tree_add_7_25_groupi_n_2146, csa_tree_add_7_25_groupi_n_2147;
  wire csa_tree_add_7_25_groupi_n_2148, csa_tree_add_7_25_groupi_n_2149, csa_tree_add_7_25_groupi_n_2150, csa_tree_add_7_25_groupi_n_2151, csa_tree_add_7_25_groupi_n_2152, csa_tree_add_7_25_groupi_n_2153, csa_tree_add_7_25_groupi_n_2154, csa_tree_add_7_25_groupi_n_2155;
  wire csa_tree_add_7_25_groupi_n_2156, csa_tree_add_7_25_groupi_n_2157, csa_tree_add_7_25_groupi_n_2158, csa_tree_add_7_25_groupi_n_2159, csa_tree_add_7_25_groupi_n_2160, csa_tree_add_7_25_groupi_n_2161, csa_tree_add_7_25_groupi_n_2162, csa_tree_add_7_25_groupi_n_2163;
  wire csa_tree_add_7_25_groupi_n_2164, csa_tree_add_7_25_groupi_n_2165, csa_tree_add_7_25_groupi_n_2166, csa_tree_add_7_25_groupi_n_2167, csa_tree_add_7_25_groupi_n_2168, csa_tree_add_7_25_groupi_n_2169, csa_tree_add_7_25_groupi_n_2170, csa_tree_add_7_25_groupi_n_2171;
  wire csa_tree_add_7_25_groupi_n_2172, csa_tree_add_7_25_groupi_n_2173, csa_tree_add_7_25_groupi_n_2174, csa_tree_add_7_25_groupi_n_2175, csa_tree_add_7_25_groupi_n_2176, csa_tree_add_7_25_groupi_n_2177, csa_tree_add_7_25_groupi_n_2178, csa_tree_add_7_25_groupi_n_2179;
  wire csa_tree_add_7_25_groupi_n_2180, csa_tree_add_7_25_groupi_n_2181, csa_tree_add_7_25_groupi_n_2182, csa_tree_add_7_25_groupi_n_2183, csa_tree_add_7_25_groupi_n_2184, csa_tree_add_7_25_groupi_n_2185, csa_tree_add_7_25_groupi_n_2186, csa_tree_add_7_25_groupi_n_2187;
  wire csa_tree_add_7_25_groupi_n_2188, csa_tree_add_7_25_groupi_n_2189, csa_tree_add_7_25_groupi_n_2190, csa_tree_add_7_25_groupi_n_2191, csa_tree_add_7_25_groupi_n_2192, csa_tree_add_7_25_groupi_n_2193, csa_tree_add_7_25_groupi_n_2194, csa_tree_add_7_25_groupi_n_2195;
  wire csa_tree_add_7_25_groupi_n_2196, csa_tree_add_7_25_groupi_n_2197, csa_tree_add_7_25_groupi_n_2198, csa_tree_add_7_25_groupi_n_2199, csa_tree_add_7_25_groupi_n_2200, csa_tree_add_7_25_groupi_n_2201, csa_tree_add_7_25_groupi_n_2202, csa_tree_add_7_25_groupi_n_2203;
  wire csa_tree_add_7_25_groupi_n_2204, csa_tree_add_7_25_groupi_n_2205, csa_tree_add_7_25_groupi_n_2206, csa_tree_add_7_25_groupi_n_2207, csa_tree_add_7_25_groupi_n_2208, csa_tree_add_7_25_groupi_n_2209, csa_tree_add_7_25_groupi_n_2210, csa_tree_add_7_25_groupi_n_2211;
  wire csa_tree_add_7_25_groupi_n_2212, csa_tree_add_7_25_groupi_n_2213, csa_tree_add_7_25_groupi_n_2214, csa_tree_add_7_25_groupi_n_2215, csa_tree_add_7_25_groupi_n_2216, csa_tree_add_7_25_groupi_n_2217, csa_tree_add_7_25_groupi_n_2218, csa_tree_add_7_25_groupi_n_2219;
  wire csa_tree_add_7_25_groupi_n_2220, csa_tree_add_7_25_groupi_n_2221, csa_tree_add_7_25_groupi_n_2222, csa_tree_add_7_25_groupi_n_2223, csa_tree_add_7_25_groupi_n_2224, csa_tree_add_7_25_groupi_n_2225, csa_tree_add_7_25_groupi_n_2226, csa_tree_add_7_25_groupi_n_2227;
  wire csa_tree_add_7_25_groupi_n_2228, csa_tree_add_7_25_groupi_n_2229, csa_tree_add_7_25_groupi_n_2230, csa_tree_add_7_25_groupi_n_2231, csa_tree_add_7_25_groupi_n_2232, csa_tree_add_7_25_groupi_n_2233, csa_tree_add_7_25_groupi_n_2234, csa_tree_add_7_25_groupi_n_2235;
  wire csa_tree_add_7_25_groupi_n_2236, csa_tree_add_7_25_groupi_n_2237, csa_tree_add_7_25_groupi_n_2238, csa_tree_add_7_25_groupi_n_2239, csa_tree_add_7_25_groupi_n_2240, csa_tree_add_7_25_groupi_n_2241, csa_tree_add_7_25_groupi_n_2242, csa_tree_add_7_25_groupi_n_2243;
  wire csa_tree_add_7_25_groupi_n_2244, csa_tree_add_7_25_groupi_n_2245, csa_tree_add_7_25_groupi_n_2246, csa_tree_add_7_25_groupi_n_2247, csa_tree_add_7_25_groupi_n_2248, csa_tree_add_7_25_groupi_n_2249, csa_tree_add_7_25_groupi_n_2250, csa_tree_add_7_25_groupi_n_2251;
  wire csa_tree_add_7_25_groupi_n_2252, csa_tree_add_7_25_groupi_n_2253, csa_tree_add_7_25_groupi_n_2254, csa_tree_add_7_25_groupi_n_2255, csa_tree_add_7_25_groupi_n_2256, csa_tree_add_7_25_groupi_n_2257, csa_tree_add_7_25_groupi_n_2258, csa_tree_add_7_25_groupi_n_2259;
  wire csa_tree_add_7_25_groupi_n_2260, csa_tree_add_7_25_groupi_n_2261, csa_tree_add_7_25_groupi_n_2262, csa_tree_add_7_25_groupi_n_2263, csa_tree_add_7_25_groupi_n_2264, csa_tree_add_7_25_groupi_n_2265, csa_tree_add_7_25_groupi_n_2266, csa_tree_add_7_25_groupi_n_2267;
  wire csa_tree_add_7_25_groupi_n_2268, csa_tree_add_7_25_groupi_n_2269, csa_tree_add_7_25_groupi_n_2270, csa_tree_add_7_25_groupi_n_2271, csa_tree_add_7_25_groupi_n_2272, csa_tree_add_7_25_groupi_n_2273, csa_tree_add_7_25_groupi_n_2274, csa_tree_add_7_25_groupi_n_2275;
  wire csa_tree_add_7_25_groupi_n_2276, csa_tree_add_7_25_groupi_n_2277, csa_tree_add_7_25_groupi_n_2278, csa_tree_add_7_25_groupi_n_2279, csa_tree_add_7_25_groupi_n_2280, csa_tree_add_7_25_groupi_n_2281, csa_tree_add_7_25_groupi_n_2282, csa_tree_add_7_25_groupi_n_2283;
  wire csa_tree_add_7_25_groupi_n_2284, csa_tree_add_7_25_groupi_n_2285, csa_tree_add_7_25_groupi_n_2286, csa_tree_add_7_25_groupi_n_2287, csa_tree_add_7_25_groupi_n_2288, csa_tree_add_7_25_groupi_n_2289, csa_tree_add_7_25_groupi_n_2290, csa_tree_add_7_25_groupi_n_2291;
  wire csa_tree_add_7_25_groupi_n_2292, csa_tree_add_7_25_groupi_n_2293, csa_tree_add_7_25_groupi_n_2294, csa_tree_add_7_25_groupi_n_2295, csa_tree_add_7_25_groupi_n_2296, csa_tree_add_7_25_groupi_n_2297, csa_tree_add_7_25_groupi_n_2298, csa_tree_add_7_25_groupi_n_2299;
  wire csa_tree_add_7_25_groupi_n_2300, csa_tree_add_7_25_groupi_n_2301, csa_tree_add_7_25_groupi_n_2302, csa_tree_add_7_25_groupi_n_2303, csa_tree_add_7_25_groupi_n_2304, csa_tree_add_7_25_groupi_n_2305, csa_tree_add_7_25_groupi_n_2306, csa_tree_add_7_25_groupi_n_2307;
  wire csa_tree_add_7_25_groupi_n_2308, csa_tree_add_7_25_groupi_n_2309, csa_tree_add_7_25_groupi_n_2310, csa_tree_add_7_25_groupi_n_2311, csa_tree_add_7_25_groupi_n_2312, csa_tree_add_7_25_groupi_n_2313, csa_tree_add_7_25_groupi_n_2314, csa_tree_add_7_25_groupi_n_2315;
  wire csa_tree_add_7_25_groupi_n_2316, csa_tree_add_7_25_groupi_n_2317, csa_tree_add_7_25_groupi_n_2318, csa_tree_add_7_25_groupi_n_2319, csa_tree_add_7_25_groupi_n_2320, csa_tree_add_7_25_groupi_n_2321, csa_tree_add_7_25_groupi_n_2322, csa_tree_add_7_25_groupi_n_2323;
  wire csa_tree_add_7_25_groupi_n_2324, csa_tree_add_7_25_groupi_n_2325, csa_tree_add_7_25_groupi_n_2326, csa_tree_add_7_25_groupi_n_2327, csa_tree_add_7_25_groupi_n_2328, csa_tree_add_7_25_groupi_n_2329, csa_tree_add_7_25_groupi_n_2330, csa_tree_add_7_25_groupi_n_2331;
  wire csa_tree_add_7_25_groupi_n_2332, csa_tree_add_7_25_groupi_n_2333, csa_tree_add_7_25_groupi_n_2334, csa_tree_add_7_25_groupi_n_2335, csa_tree_add_7_25_groupi_n_2336, csa_tree_add_7_25_groupi_n_2337, csa_tree_add_7_25_groupi_n_2338, csa_tree_add_7_25_groupi_n_2339;
  wire csa_tree_add_7_25_groupi_n_2340, csa_tree_add_7_25_groupi_n_2341, csa_tree_add_7_25_groupi_n_2342, csa_tree_add_7_25_groupi_n_2343, csa_tree_add_7_25_groupi_n_2344, csa_tree_add_7_25_groupi_n_2345, csa_tree_add_7_25_groupi_n_2346, csa_tree_add_7_25_groupi_n_2347;
  wire csa_tree_add_7_25_groupi_n_2349, csa_tree_add_7_25_groupi_n_2350, csa_tree_add_7_25_groupi_n_2351, csa_tree_add_7_25_groupi_n_2352, csa_tree_add_7_25_groupi_n_2353, csa_tree_add_7_25_groupi_n_2354, csa_tree_add_7_25_groupi_n_2355, csa_tree_add_7_25_groupi_n_2356;
  wire csa_tree_add_7_25_groupi_n_2357, csa_tree_add_7_25_groupi_n_2358, csa_tree_add_7_25_groupi_n_2359, csa_tree_add_7_25_groupi_n_2360, csa_tree_add_7_25_groupi_n_2361, csa_tree_add_7_25_groupi_n_2362, csa_tree_add_7_25_groupi_n_2363, csa_tree_add_7_25_groupi_n_2364;
  wire csa_tree_add_7_25_groupi_n_2365, csa_tree_add_7_25_groupi_n_2366, csa_tree_add_7_25_groupi_n_2367, csa_tree_add_7_25_groupi_n_2368, csa_tree_add_7_25_groupi_n_2369, csa_tree_add_7_25_groupi_n_2370, csa_tree_add_7_25_groupi_n_2371, csa_tree_add_7_25_groupi_n_2372;
  wire csa_tree_add_7_25_groupi_n_2373, csa_tree_add_7_25_groupi_n_2374, csa_tree_add_7_25_groupi_n_2375, csa_tree_add_7_25_groupi_n_2376, csa_tree_add_7_25_groupi_n_2377, csa_tree_add_7_25_groupi_n_2378, csa_tree_add_7_25_groupi_n_2379, csa_tree_add_7_25_groupi_n_2380;
  wire csa_tree_add_7_25_groupi_n_2381, csa_tree_add_7_25_groupi_n_2382, csa_tree_add_7_25_groupi_n_2383, csa_tree_add_7_25_groupi_n_2384, csa_tree_add_7_25_groupi_n_2385, csa_tree_add_7_25_groupi_n_2386, csa_tree_add_7_25_groupi_n_2387, csa_tree_add_7_25_groupi_n_2388;
  wire csa_tree_add_7_25_groupi_n_2389, csa_tree_add_7_25_groupi_n_2390, csa_tree_add_7_25_groupi_n_2391, csa_tree_add_7_25_groupi_n_2392, csa_tree_add_7_25_groupi_n_2393, csa_tree_add_7_25_groupi_n_2394, csa_tree_add_7_25_groupi_n_2395, csa_tree_add_7_25_groupi_n_2396;
  wire csa_tree_add_7_25_groupi_n_2397, csa_tree_add_7_25_groupi_n_2398, csa_tree_add_7_25_groupi_n_2399, csa_tree_add_7_25_groupi_n_2400, csa_tree_add_7_25_groupi_n_2401, csa_tree_add_7_25_groupi_n_2402, csa_tree_add_7_25_groupi_n_2403, csa_tree_add_7_25_groupi_n_2404;
  wire csa_tree_add_7_25_groupi_n_2405, csa_tree_add_7_25_groupi_n_2406, csa_tree_add_7_25_groupi_n_2407, csa_tree_add_7_25_groupi_n_2408, csa_tree_add_7_25_groupi_n_2409, csa_tree_add_7_25_groupi_n_2410, csa_tree_add_7_25_groupi_n_2411, csa_tree_add_7_25_groupi_n_2412;
  wire csa_tree_add_7_25_groupi_n_2413, csa_tree_add_7_25_groupi_n_2414, csa_tree_add_7_25_groupi_n_2415, csa_tree_add_7_25_groupi_n_2416, csa_tree_add_7_25_groupi_n_2417, csa_tree_add_7_25_groupi_n_2418, csa_tree_add_7_25_groupi_n_2419, csa_tree_add_7_25_groupi_n_2420;
  wire csa_tree_add_7_25_groupi_n_2421, csa_tree_add_7_25_groupi_n_2422, csa_tree_add_7_25_groupi_n_2423, csa_tree_add_7_25_groupi_n_2424, csa_tree_add_7_25_groupi_n_2425, csa_tree_add_7_25_groupi_n_2426, csa_tree_add_7_25_groupi_n_2427, csa_tree_add_7_25_groupi_n_2428;
  wire csa_tree_add_7_25_groupi_n_2429, csa_tree_add_7_25_groupi_n_2430, csa_tree_add_7_25_groupi_n_2431, csa_tree_add_7_25_groupi_n_2432, csa_tree_add_7_25_groupi_n_2433, csa_tree_add_7_25_groupi_n_2434, csa_tree_add_7_25_groupi_n_2435, csa_tree_add_7_25_groupi_n_2436;
  wire csa_tree_add_7_25_groupi_n_2437, csa_tree_add_7_25_groupi_n_2438, csa_tree_add_7_25_groupi_n_2439, csa_tree_add_7_25_groupi_n_2440, csa_tree_add_7_25_groupi_n_2441, csa_tree_add_7_25_groupi_n_2442, csa_tree_add_7_25_groupi_n_2443, csa_tree_add_7_25_groupi_n_2444;
  wire csa_tree_add_7_25_groupi_n_2445, csa_tree_add_7_25_groupi_n_2446, csa_tree_add_7_25_groupi_n_2447, csa_tree_add_7_25_groupi_n_2448, csa_tree_add_7_25_groupi_n_2449, csa_tree_add_7_25_groupi_n_2450, csa_tree_add_7_25_groupi_n_2451, csa_tree_add_7_25_groupi_n_2452;
  wire csa_tree_add_7_25_groupi_n_2453, csa_tree_add_7_25_groupi_n_2454, csa_tree_add_7_25_groupi_n_2455, csa_tree_add_7_25_groupi_n_2456, csa_tree_add_7_25_groupi_n_2457, csa_tree_add_7_25_groupi_n_2458, csa_tree_add_7_25_groupi_n_2459, csa_tree_add_7_25_groupi_n_2460;
  wire csa_tree_add_7_25_groupi_n_2461, csa_tree_add_7_25_groupi_n_2462, csa_tree_add_7_25_groupi_n_2463, csa_tree_add_7_25_groupi_n_2464, csa_tree_add_7_25_groupi_n_2465, csa_tree_add_7_25_groupi_n_2466, csa_tree_add_7_25_groupi_n_2467, csa_tree_add_7_25_groupi_n_2468;
  wire csa_tree_add_7_25_groupi_n_2469, csa_tree_add_7_25_groupi_n_2470, csa_tree_add_7_25_groupi_n_2471, csa_tree_add_7_25_groupi_n_2472, csa_tree_add_7_25_groupi_n_2473, csa_tree_add_7_25_groupi_n_2474, csa_tree_add_7_25_groupi_n_2475, csa_tree_add_7_25_groupi_n_2476;
  wire csa_tree_add_7_25_groupi_n_2477, csa_tree_add_7_25_groupi_n_2478, csa_tree_add_7_25_groupi_n_2479, csa_tree_add_7_25_groupi_n_2480, csa_tree_add_7_25_groupi_n_2481, csa_tree_add_7_25_groupi_n_2482, csa_tree_add_7_25_groupi_n_2483, csa_tree_add_7_25_groupi_n_2484;
  wire csa_tree_add_7_25_groupi_n_2485, csa_tree_add_7_25_groupi_n_2486, csa_tree_add_7_25_groupi_n_2487, csa_tree_add_7_25_groupi_n_2488, csa_tree_add_7_25_groupi_n_2489, csa_tree_add_7_25_groupi_n_2490, csa_tree_add_7_25_groupi_n_2491, csa_tree_add_7_25_groupi_n_2492;
  wire csa_tree_add_7_25_groupi_n_2494, csa_tree_add_7_25_groupi_n_2495, csa_tree_add_7_25_groupi_n_2496, csa_tree_add_7_25_groupi_n_2497, csa_tree_add_7_25_groupi_n_2498, csa_tree_add_7_25_groupi_n_2499, csa_tree_add_7_25_groupi_n_2500, csa_tree_add_7_25_groupi_n_2501;
  wire csa_tree_add_7_25_groupi_n_2502, csa_tree_add_7_25_groupi_n_2503, csa_tree_add_7_25_groupi_n_2504, csa_tree_add_7_25_groupi_n_2505, csa_tree_add_7_25_groupi_n_2506, csa_tree_add_7_25_groupi_n_2507, csa_tree_add_7_25_groupi_n_2508, csa_tree_add_7_25_groupi_n_2509;
  wire csa_tree_add_7_25_groupi_n_2510, csa_tree_add_7_25_groupi_n_2511, csa_tree_add_7_25_groupi_n_2512, csa_tree_add_7_25_groupi_n_2513, csa_tree_add_7_25_groupi_n_2514, csa_tree_add_7_25_groupi_n_2515, csa_tree_add_7_25_groupi_n_2516, csa_tree_add_7_25_groupi_n_2517;
  wire csa_tree_add_7_25_groupi_n_2518, csa_tree_add_7_25_groupi_n_2519, csa_tree_add_7_25_groupi_n_2520, csa_tree_add_7_25_groupi_n_2521, csa_tree_add_7_25_groupi_n_2522, csa_tree_add_7_25_groupi_n_2523, csa_tree_add_7_25_groupi_n_2524, csa_tree_add_7_25_groupi_n_2525;
  wire csa_tree_add_7_25_groupi_n_2526, csa_tree_add_7_25_groupi_n_2527, csa_tree_add_7_25_groupi_n_2528, csa_tree_add_7_25_groupi_n_2529, csa_tree_add_7_25_groupi_n_2530, csa_tree_add_7_25_groupi_n_2531, csa_tree_add_7_25_groupi_n_2532, csa_tree_add_7_25_groupi_n_2533;
  wire csa_tree_add_7_25_groupi_n_2534, csa_tree_add_7_25_groupi_n_2535, csa_tree_add_7_25_groupi_n_2536, csa_tree_add_7_25_groupi_n_2537, csa_tree_add_7_25_groupi_n_2538, csa_tree_add_7_25_groupi_n_2539, csa_tree_add_7_25_groupi_n_2540, csa_tree_add_7_25_groupi_n_2541;
  wire csa_tree_add_7_25_groupi_n_2542, csa_tree_add_7_25_groupi_n_2543, csa_tree_add_7_25_groupi_n_2544, csa_tree_add_7_25_groupi_n_2545, csa_tree_add_7_25_groupi_n_2546, csa_tree_add_7_25_groupi_n_2547, csa_tree_add_7_25_groupi_n_2548, csa_tree_add_7_25_groupi_n_2549;
  wire csa_tree_add_7_25_groupi_n_2550, csa_tree_add_7_25_groupi_n_2551, csa_tree_add_7_25_groupi_n_2552, csa_tree_add_7_25_groupi_n_2553, csa_tree_add_7_25_groupi_n_2554, csa_tree_add_7_25_groupi_n_2555, csa_tree_add_7_25_groupi_n_2556, csa_tree_add_7_25_groupi_n_2557;
  wire csa_tree_add_7_25_groupi_n_2558, csa_tree_add_7_25_groupi_n_2559, csa_tree_add_7_25_groupi_n_2560, csa_tree_add_7_25_groupi_n_2561, csa_tree_add_7_25_groupi_n_2562, csa_tree_add_7_25_groupi_n_2563, csa_tree_add_7_25_groupi_n_2564, csa_tree_add_7_25_groupi_n_2565;
  wire csa_tree_add_7_25_groupi_n_2566, csa_tree_add_7_25_groupi_n_2567, csa_tree_add_7_25_groupi_n_2568, csa_tree_add_7_25_groupi_n_2569, csa_tree_add_7_25_groupi_n_2570, csa_tree_add_7_25_groupi_n_2571, csa_tree_add_7_25_groupi_n_2572, csa_tree_add_7_25_groupi_n_2573;
  wire csa_tree_add_7_25_groupi_n_2574, csa_tree_add_7_25_groupi_n_2575, csa_tree_add_7_25_groupi_n_2576, csa_tree_add_7_25_groupi_n_2577, csa_tree_add_7_25_groupi_n_2578, csa_tree_add_7_25_groupi_n_2579, csa_tree_add_7_25_groupi_n_2580, csa_tree_add_7_25_groupi_n_2581;
  wire csa_tree_add_7_25_groupi_n_2582, csa_tree_add_7_25_groupi_n_2583, csa_tree_add_7_25_groupi_n_2584, csa_tree_add_7_25_groupi_n_2585, csa_tree_add_7_25_groupi_n_2586, csa_tree_add_7_25_groupi_n_2587, csa_tree_add_7_25_groupi_n_2588, csa_tree_add_7_25_groupi_n_2589;
  wire csa_tree_add_7_25_groupi_n_2590, csa_tree_add_7_25_groupi_n_2591, csa_tree_add_7_25_groupi_n_2592, csa_tree_add_7_25_groupi_n_2593, csa_tree_add_7_25_groupi_n_2594, csa_tree_add_7_25_groupi_n_2595, csa_tree_add_7_25_groupi_n_2596, csa_tree_add_7_25_groupi_n_2597;
  wire csa_tree_add_7_25_groupi_n_2598, csa_tree_add_7_25_groupi_n_2599, csa_tree_add_7_25_groupi_n_2600, csa_tree_add_7_25_groupi_n_2601, csa_tree_add_7_25_groupi_n_2602, csa_tree_add_7_25_groupi_n_2603, csa_tree_add_7_25_groupi_n_2604, csa_tree_add_7_25_groupi_n_2605;
  wire csa_tree_add_7_25_groupi_n_2606, csa_tree_add_7_25_groupi_n_2607, csa_tree_add_7_25_groupi_n_2608, csa_tree_add_7_25_groupi_n_2609, csa_tree_add_7_25_groupi_n_2610, csa_tree_add_7_25_groupi_n_2611, csa_tree_add_7_25_groupi_n_2612, csa_tree_add_7_25_groupi_n_2613;
  wire csa_tree_add_7_25_groupi_n_2614, csa_tree_add_7_25_groupi_n_2615, csa_tree_add_7_25_groupi_n_2616, csa_tree_add_7_25_groupi_n_2617, csa_tree_add_7_25_groupi_n_2618, csa_tree_add_7_25_groupi_n_2619, csa_tree_add_7_25_groupi_n_2620, csa_tree_add_7_25_groupi_n_2621;
  wire csa_tree_add_7_25_groupi_n_2622, csa_tree_add_7_25_groupi_n_2623, csa_tree_add_7_25_groupi_n_2624, csa_tree_add_7_25_groupi_n_2625, csa_tree_add_7_25_groupi_n_2626, csa_tree_add_7_25_groupi_n_2627, csa_tree_add_7_25_groupi_n_2628, csa_tree_add_7_25_groupi_n_2629;
  wire csa_tree_add_7_25_groupi_n_2630, csa_tree_add_7_25_groupi_n_2631, csa_tree_add_7_25_groupi_n_2632, csa_tree_add_7_25_groupi_n_2633, csa_tree_add_7_25_groupi_n_2634, csa_tree_add_7_25_groupi_n_2635, csa_tree_add_7_25_groupi_n_2636, csa_tree_add_7_25_groupi_n_2637;
  wire csa_tree_add_7_25_groupi_n_2638, csa_tree_add_7_25_groupi_n_2639, csa_tree_add_7_25_groupi_n_2640, csa_tree_add_7_25_groupi_n_2641, csa_tree_add_7_25_groupi_n_2642, csa_tree_add_7_25_groupi_n_2643, csa_tree_add_7_25_groupi_n_2644, csa_tree_add_7_25_groupi_n_2645;
  wire csa_tree_add_7_25_groupi_n_2646, csa_tree_add_7_25_groupi_n_2647, csa_tree_add_7_25_groupi_n_2648, csa_tree_add_7_25_groupi_n_2649, csa_tree_add_7_25_groupi_n_2650, csa_tree_add_7_25_groupi_n_2651, csa_tree_add_7_25_groupi_n_2652, csa_tree_add_7_25_groupi_n_2653;
  wire csa_tree_add_7_25_groupi_n_2654, csa_tree_add_7_25_groupi_n_2655, csa_tree_add_7_25_groupi_n_2656, csa_tree_add_7_25_groupi_n_2657, csa_tree_add_7_25_groupi_n_2658, csa_tree_add_7_25_groupi_n_2659, csa_tree_add_7_25_groupi_n_2660, csa_tree_add_7_25_groupi_n_2661;
  wire csa_tree_add_7_25_groupi_n_2662, csa_tree_add_7_25_groupi_n_2663, csa_tree_add_7_25_groupi_n_2664, csa_tree_add_7_25_groupi_n_2665, csa_tree_add_7_25_groupi_n_2666, csa_tree_add_7_25_groupi_n_2667, csa_tree_add_7_25_groupi_n_2668, csa_tree_add_7_25_groupi_n_2669;
  wire csa_tree_add_7_25_groupi_n_2670, csa_tree_add_7_25_groupi_n_2671, csa_tree_add_7_25_groupi_n_2672, csa_tree_add_7_25_groupi_n_2673, csa_tree_add_7_25_groupi_n_2674, csa_tree_add_7_25_groupi_n_2675, csa_tree_add_7_25_groupi_n_2676, csa_tree_add_7_25_groupi_n_2677;
  wire csa_tree_add_7_25_groupi_n_2678, csa_tree_add_7_25_groupi_n_2679, csa_tree_add_7_25_groupi_n_2680, csa_tree_add_7_25_groupi_n_2681, csa_tree_add_7_25_groupi_n_2682, csa_tree_add_7_25_groupi_n_2683, csa_tree_add_7_25_groupi_n_2684, csa_tree_add_7_25_groupi_n_2685;
  wire csa_tree_add_7_25_groupi_n_2686, csa_tree_add_7_25_groupi_n_2687, csa_tree_add_7_25_groupi_n_2688, csa_tree_add_7_25_groupi_n_2689, csa_tree_add_7_25_groupi_n_2690, csa_tree_add_7_25_groupi_n_2691, csa_tree_add_7_25_groupi_n_2692, csa_tree_add_7_25_groupi_n_2693;
  wire csa_tree_add_7_25_groupi_n_2694, csa_tree_add_7_25_groupi_n_2695, csa_tree_add_7_25_groupi_n_2696, csa_tree_add_7_25_groupi_n_2697, csa_tree_add_7_25_groupi_n_2698, csa_tree_add_7_25_groupi_n_2699, csa_tree_add_7_25_groupi_n_2700, csa_tree_add_7_25_groupi_n_2701;
  wire csa_tree_add_7_25_groupi_n_2702, csa_tree_add_7_25_groupi_n_2703, csa_tree_add_7_25_groupi_n_2704, csa_tree_add_7_25_groupi_n_2705, csa_tree_add_7_25_groupi_n_2706, csa_tree_add_7_25_groupi_n_2707, csa_tree_add_7_25_groupi_n_2708, csa_tree_add_7_25_groupi_n_2709;
  wire csa_tree_add_7_25_groupi_n_2710, csa_tree_add_7_25_groupi_n_2711, csa_tree_add_7_25_groupi_n_2712, csa_tree_add_7_25_groupi_n_2713, csa_tree_add_7_25_groupi_n_2714, csa_tree_add_7_25_groupi_n_2715, csa_tree_add_7_25_groupi_n_2716, csa_tree_add_7_25_groupi_n_2717;
  wire csa_tree_add_7_25_groupi_n_2718, csa_tree_add_7_25_groupi_n_2719, csa_tree_add_7_25_groupi_n_2720, csa_tree_add_7_25_groupi_n_2721, csa_tree_add_7_25_groupi_n_2722, csa_tree_add_7_25_groupi_n_2723, csa_tree_add_7_25_groupi_n_2724, csa_tree_add_7_25_groupi_n_2725;
  wire csa_tree_add_7_25_groupi_n_2726, csa_tree_add_7_25_groupi_n_2727, csa_tree_add_7_25_groupi_n_2728, csa_tree_add_7_25_groupi_n_2729, csa_tree_add_7_25_groupi_n_2730, csa_tree_add_7_25_groupi_n_2731, csa_tree_add_7_25_groupi_n_2732, csa_tree_add_7_25_groupi_n_2733;
  wire csa_tree_add_7_25_groupi_n_2734, csa_tree_add_7_25_groupi_n_2735, csa_tree_add_7_25_groupi_n_2736, csa_tree_add_7_25_groupi_n_2737, csa_tree_add_7_25_groupi_n_2738, csa_tree_add_7_25_groupi_n_2739, csa_tree_add_7_25_groupi_n_2740, csa_tree_add_7_25_groupi_n_2741;
  wire csa_tree_add_7_25_groupi_n_2742, csa_tree_add_7_25_groupi_n_2743, csa_tree_add_7_25_groupi_n_2744, csa_tree_add_7_25_groupi_n_2745, csa_tree_add_7_25_groupi_n_2746, csa_tree_add_7_25_groupi_n_2747, csa_tree_add_7_25_groupi_n_2748, csa_tree_add_7_25_groupi_n_2749;
  wire csa_tree_add_7_25_groupi_n_2750, csa_tree_add_7_25_groupi_n_2751, csa_tree_add_7_25_groupi_n_2752, csa_tree_add_7_25_groupi_n_2753, csa_tree_add_7_25_groupi_n_2754, csa_tree_add_7_25_groupi_n_2755, csa_tree_add_7_25_groupi_n_2756, csa_tree_add_7_25_groupi_n_2757;
  wire csa_tree_add_7_25_groupi_n_2758, csa_tree_add_7_25_groupi_n_2759, csa_tree_add_7_25_groupi_n_2760, csa_tree_add_7_25_groupi_n_2761, csa_tree_add_7_25_groupi_n_2762, csa_tree_add_7_25_groupi_n_2763, csa_tree_add_7_25_groupi_n_2764, csa_tree_add_7_25_groupi_n_2765;
  wire csa_tree_add_7_25_groupi_n_2766, csa_tree_add_7_25_groupi_n_2767, csa_tree_add_7_25_groupi_n_2768, csa_tree_add_7_25_groupi_n_2769, csa_tree_add_7_25_groupi_n_2770, csa_tree_add_7_25_groupi_n_2771, csa_tree_add_7_25_groupi_n_2772, csa_tree_add_7_25_groupi_n_2773;
  wire csa_tree_add_7_25_groupi_n_2774, csa_tree_add_7_25_groupi_n_2775, csa_tree_add_7_25_groupi_n_2776, csa_tree_add_7_25_groupi_n_2777, csa_tree_add_7_25_groupi_n_2778, csa_tree_add_7_25_groupi_n_2779, csa_tree_add_7_25_groupi_n_2780, csa_tree_add_7_25_groupi_n_2781;
  wire csa_tree_add_7_25_groupi_n_2782, csa_tree_add_7_25_groupi_n_2783, csa_tree_add_7_25_groupi_n_2784, csa_tree_add_7_25_groupi_n_2785, csa_tree_add_7_25_groupi_n_2786, csa_tree_add_7_25_groupi_n_2787, csa_tree_add_7_25_groupi_n_2788, csa_tree_add_7_25_groupi_n_2789;
  wire csa_tree_add_7_25_groupi_n_2790, csa_tree_add_7_25_groupi_n_2791, csa_tree_add_7_25_groupi_n_2792, csa_tree_add_7_25_groupi_n_2793, csa_tree_add_7_25_groupi_n_2794, csa_tree_add_7_25_groupi_n_2795, csa_tree_add_7_25_groupi_n_2796, csa_tree_add_7_25_groupi_n_2797;
  wire csa_tree_add_7_25_groupi_n_2798, csa_tree_add_7_25_groupi_n_2799, csa_tree_add_7_25_groupi_n_2800, csa_tree_add_7_25_groupi_n_2801, csa_tree_add_7_25_groupi_n_2802, csa_tree_add_7_25_groupi_n_2803, csa_tree_add_7_25_groupi_n_2804, csa_tree_add_7_25_groupi_n_2805;
  wire csa_tree_add_7_25_groupi_n_2806, csa_tree_add_7_25_groupi_n_2807, csa_tree_add_7_25_groupi_n_2808, csa_tree_add_7_25_groupi_n_2809, csa_tree_add_7_25_groupi_n_2810, csa_tree_add_7_25_groupi_n_2811, csa_tree_add_7_25_groupi_n_2812, csa_tree_add_7_25_groupi_n_2813;
  wire csa_tree_add_7_25_groupi_n_2814, csa_tree_add_7_25_groupi_n_2815, csa_tree_add_7_25_groupi_n_2816, csa_tree_add_7_25_groupi_n_2817, csa_tree_add_7_25_groupi_n_2818, csa_tree_add_7_25_groupi_n_2819, csa_tree_add_7_25_groupi_n_2820, csa_tree_add_7_25_groupi_n_2821;
  wire csa_tree_add_7_25_groupi_n_2822, csa_tree_add_7_25_groupi_n_2823, csa_tree_add_7_25_groupi_n_2824, csa_tree_add_7_25_groupi_n_2825, csa_tree_add_7_25_groupi_n_2826, csa_tree_add_7_25_groupi_n_2827, csa_tree_add_7_25_groupi_n_2828, csa_tree_add_7_25_groupi_n_2829;
  wire csa_tree_add_7_25_groupi_n_2830, csa_tree_add_7_25_groupi_n_2831, csa_tree_add_7_25_groupi_n_2832, csa_tree_add_7_25_groupi_n_2833, csa_tree_add_7_25_groupi_n_2834, csa_tree_add_7_25_groupi_n_2835, csa_tree_add_7_25_groupi_n_2836, csa_tree_add_7_25_groupi_n_2837;
  wire csa_tree_add_7_25_groupi_n_2838, csa_tree_add_7_25_groupi_n_2839, csa_tree_add_7_25_groupi_n_2840, csa_tree_add_7_25_groupi_n_2841, csa_tree_add_7_25_groupi_n_2842, csa_tree_add_7_25_groupi_n_2843, csa_tree_add_7_25_groupi_n_2844, csa_tree_add_7_25_groupi_n_2845;
  wire csa_tree_add_7_25_groupi_n_2846, csa_tree_add_7_25_groupi_n_2847, csa_tree_add_7_25_groupi_n_2848, csa_tree_add_7_25_groupi_n_2849, csa_tree_add_7_25_groupi_n_2850, csa_tree_add_7_25_groupi_n_2851, csa_tree_add_7_25_groupi_n_2852, csa_tree_add_7_25_groupi_n_2853;
  wire csa_tree_add_7_25_groupi_n_2854, csa_tree_add_7_25_groupi_n_2855, csa_tree_add_7_25_groupi_n_2856, csa_tree_add_7_25_groupi_n_2857, csa_tree_add_7_25_groupi_n_2858, csa_tree_add_7_25_groupi_n_2859, csa_tree_add_7_25_groupi_n_2860, csa_tree_add_7_25_groupi_n_2861;
  wire csa_tree_add_7_25_groupi_n_2862, csa_tree_add_7_25_groupi_n_2863, csa_tree_add_7_25_groupi_n_2864, csa_tree_add_7_25_groupi_n_2865, csa_tree_add_7_25_groupi_n_2866, csa_tree_add_7_25_groupi_n_2867, csa_tree_add_7_25_groupi_n_2868, csa_tree_add_7_25_groupi_n_2869;
  wire csa_tree_add_7_25_groupi_n_2870, csa_tree_add_7_25_groupi_n_2871, csa_tree_add_7_25_groupi_n_2872, csa_tree_add_7_25_groupi_n_2873, csa_tree_add_7_25_groupi_n_2874, csa_tree_add_7_25_groupi_n_2875, csa_tree_add_7_25_groupi_n_2876, csa_tree_add_7_25_groupi_n_2877;
  wire csa_tree_add_7_25_groupi_n_2878, csa_tree_add_7_25_groupi_n_2879, csa_tree_add_7_25_groupi_n_2880, csa_tree_add_7_25_groupi_n_2881, csa_tree_add_7_25_groupi_n_2882, csa_tree_add_7_25_groupi_n_2883, csa_tree_add_7_25_groupi_n_2884, csa_tree_add_7_25_groupi_n_2885;
  wire csa_tree_add_7_25_groupi_n_2886, csa_tree_add_7_25_groupi_n_2887, csa_tree_add_7_25_groupi_n_2888, csa_tree_add_7_25_groupi_n_2889, csa_tree_add_7_25_groupi_n_2890, csa_tree_add_7_25_groupi_n_2891, csa_tree_add_7_25_groupi_n_2892, csa_tree_add_7_25_groupi_n_2893;
  wire csa_tree_add_7_25_groupi_n_2894, csa_tree_add_7_25_groupi_n_2895, csa_tree_add_7_25_groupi_n_2896, csa_tree_add_7_25_groupi_n_2897, csa_tree_add_7_25_groupi_n_2898, csa_tree_add_7_25_groupi_n_2899, csa_tree_add_7_25_groupi_n_2900, csa_tree_add_7_25_groupi_n_2901;
  wire csa_tree_add_7_25_groupi_n_2902, csa_tree_add_7_25_groupi_n_2903, csa_tree_add_7_25_groupi_n_2904, csa_tree_add_7_25_groupi_n_2905, csa_tree_add_7_25_groupi_n_2906, csa_tree_add_7_25_groupi_n_2907, csa_tree_add_7_25_groupi_n_2908, csa_tree_add_7_25_groupi_n_2909;
  wire csa_tree_add_7_25_groupi_n_2910, csa_tree_add_7_25_groupi_n_2911, csa_tree_add_7_25_groupi_n_2912, csa_tree_add_7_25_groupi_n_2913, csa_tree_add_7_25_groupi_n_2914, csa_tree_add_7_25_groupi_n_2915, csa_tree_add_7_25_groupi_n_2916, csa_tree_add_7_25_groupi_n_2917;
  wire csa_tree_add_7_25_groupi_n_2918, csa_tree_add_7_25_groupi_n_2919, csa_tree_add_7_25_groupi_n_2920, csa_tree_add_7_25_groupi_n_2921, csa_tree_add_7_25_groupi_n_2922, csa_tree_add_7_25_groupi_n_2923, csa_tree_add_7_25_groupi_n_2924, csa_tree_add_7_25_groupi_n_2925;
  wire csa_tree_add_7_25_groupi_n_2926, csa_tree_add_7_25_groupi_n_2927, csa_tree_add_7_25_groupi_n_2928, csa_tree_add_7_25_groupi_n_2929, csa_tree_add_7_25_groupi_n_2930, csa_tree_add_7_25_groupi_n_2931, csa_tree_add_7_25_groupi_n_2932, csa_tree_add_7_25_groupi_n_2933;
  wire csa_tree_add_7_25_groupi_n_2934, csa_tree_add_7_25_groupi_n_2935, csa_tree_add_7_25_groupi_n_2936, csa_tree_add_7_25_groupi_n_2937, csa_tree_add_7_25_groupi_n_2938, csa_tree_add_7_25_groupi_n_2939, csa_tree_add_7_25_groupi_n_2940, csa_tree_add_7_25_groupi_n_2941;
  wire csa_tree_add_7_25_groupi_n_2942, csa_tree_add_7_25_groupi_n_2943, csa_tree_add_7_25_groupi_n_2944, csa_tree_add_7_25_groupi_n_2945, csa_tree_add_7_25_groupi_n_2946, csa_tree_add_7_25_groupi_n_2947, csa_tree_add_7_25_groupi_n_2948, csa_tree_add_7_25_groupi_n_2949;
  wire csa_tree_add_7_25_groupi_n_2950, csa_tree_add_7_25_groupi_n_2951, csa_tree_add_7_25_groupi_n_2952, csa_tree_add_7_25_groupi_n_2953, csa_tree_add_7_25_groupi_n_2954, csa_tree_add_7_25_groupi_n_2955, csa_tree_add_7_25_groupi_n_2956, csa_tree_add_7_25_groupi_n_2957;
  wire csa_tree_add_7_25_groupi_n_2958, csa_tree_add_7_25_groupi_n_2959, csa_tree_add_7_25_groupi_n_2960, csa_tree_add_7_25_groupi_n_2961, csa_tree_add_7_25_groupi_n_2962, csa_tree_add_7_25_groupi_n_2963, csa_tree_add_7_25_groupi_n_2964, csa_tree_add_7_25_groupi_n_2965;
  wire csa_tree_add_7_25_groupi_n_2966, csa_tree_add_7_25_groupi_n_2967, csa_tree_add_7_25_groupi_n_2968, csa_tree_add_7_25_groupi_n_2969, csa_tree_add_7_25_groupi_n_2970, csa_tree_add_7_25_groupi_n_2971, csa_tree_add_7_25_groupi_n_2972, csa_tree_add_7_25_groupi_n_2973;
  wire csa_tree_add_7_25_groupi_n_2974, csa_tree_add_7_25_groupi_n_2975, csa_tree_add_7_25_groupi_n_2976, csa_tree_add_7_25_groupi_n_2977, csa_tree_add_7_25_groupi_n_2978, csa_tree_add_7_25_groupi_n_2979, csa_tree_add_7_25_groupi_n_2980, csa_tree_add_7_25_groupi_n_2981;
  wire csa_tree_add_7_25_groupi_n_2982, csa_tree_add_7_25_groupi_n_2983, csa_tree_add_7_25_groupi_n_2984, csa_tree_add_7_25_groupi_n_2985, csa_tree_add_7_25_groupi_n_2986, csa_tree_add_7_25_groupi_n_2987, csa_tree_add_7_25_groupi_n_2988, csa_tree_add_7_25_groupi_n_2989;
  wire csa_tree_add_7_25_groupi_n_2990, csa_tree_add_7_25_groupi_n_2991, csa_tree_add_7_25_groupi_n_2992, csa_tree_add_7_25_groupi_n_2993, csa_tree_add_7_25_groupi_n_2994, csa_tree_add_7_25_groupi_n_2995, csa_tree_add_7_25_groupi_n_2996, csa_tree_add_7_25_groupi_n_2997;
  wire csa_tree_add_7_25_groupi_n_2998, csa_tree_add_7_25_groupi_n_2999, csa_tree_add_7_25_groupi_n_3000, csa_tree_add_7_25_groupi_n_3001, csa_tree_add_7_25_groupi_n_3002, csa_tree_add_7_25_groupi_n_3003, csa_tree_add_7_25_groupi_n_3004, csa_tree_add_7_25_groupi_n_3005;
  wire csa_tree_add_7_25_groupi_n_3006, csa_tree_add_7_25_groupi_n_3007, csa_tree_add_7_25_groupi_n_3008, csa_tree_add_7_25_groupi_n_3009, csa_tree_add_7_25_groupi_n_3010, csa_tree_add_7_25_groupi_n_3011, csa_tree_add_7_25_groupi_n_3012, csa_tree_add_7_25_groupi_n_3013;
  wire csa_tree_add_7_25_groupi_n_3014, csa_tree_add_7_25_groupi_n_3015, csa_tree_add_7_25_groupi_n_3016, csa_tree_add_7_25_groupi_n_3017, csa_tree_add_7_25_groupi_n_3018, csa_tree_add_7_25_groupi_n_3019, csa_tree_add_7_25_groupi_n_3020, csa_tree_add_7_25_groupi_n_3021;
  wire csa_tree_add_7_25_groupi_n_3022, csa_tree_add_7_25_groupi_n_3023, csa_tree_add_7_25_groupi_n_3024, csa_tree_add_7_25_groupi_n_3025, csa_tree_add_7_25_groupi_n_3026, csa_tree_add_7_25_groupi_n_3027, csa_tree_add_7_25_groupi_n_3028, csa_tree_add_7_25_groupi_n_3029;
  wire csa_tree_add_7_25_groupi_n_3030, csa_tree_add_7_25_groupi_n_3031, csa_tree_add_7_25_groupi_n_3032, csa_tree_add_7_25_groupi_n_3033, csa_tree_add_7_25_groupi_n_3034, csa_tree_add_7_25_groupi_n_3035, csa_tree_add_7_25_groupi_n_3036, csa_tree_add_7_25_groupi_n_3037;
  wire csa_tree_add_7_25_groupi_n_3038, csa_tree_add_7_25_groupi_n_3039, csa_tree_add_7_25_groupi_n_3040, csa_tree_add_7_25_groupi_n_3041, csa_tree_add_7_25_groupi_n_3042, csa_tree_add_7_25_groupi_n_3043, csa_tree_add_7_25_groupi_n_3044, csa_tree_add_7_25_groupi_n_3045;
  wire csa_tree_add_7_25_groupi_n_3046, csa_tree_add_7_25_groupi_n_3047, csa_tree_add_7_25_groupi_n_3048, csa_tree_add_7_25_groupi_n_3049, csa_tree_add_7_25_groupi_n_3050, csa_tree_add_7_25_groupi_n_3051, csa_tree_add_7_25_groupi_n_3052, csa_tree_add_7_25_groupi_n_3053;
  wire csa_tree_add_7_25_groupi_n_3054, csa_tree_add_7_25_groupi_n_3055, csa_tree_add_7_25_groupi_n_3056, csa_tree_add_7_25_groupi_n_3057, csa_tree_add_7_25_groupi_n_3058, csa_tree_add_7_25_groupi_n_3059, csa_tree_add_7_25_groupi_n_3060, csa_tree_add_7_25_groupi_n_3061;
  wire csa_tree_add_7_25_groupi_n_3062, csa_tree_add_7_25_groupi_n_3063, csa_tree_add_7_25_groupi_n_3064, csa_tree_add_7_25_groupi_n_3065, csa_tree_add_7_25_groupi_n_3066, csa_tree_add_7_25_groupi_n_3067, csa_tree_add_7_25_groupi_n_3068, csa_tree_add_7_25_groupi_n_3069;
  wire csa_tree_add_7_25_groupi_n_3070, csa_tree_add_7_25_groupi_n_3071, csa_tree_add_7_25_groupi_n_3072, csa_tree_add_7_25_groupi_n_3073, csa_tree_add_7_25_groupi_n_3074, csa_tree_add_7_25_groupi_n_3075, csa_tree_add_7_25_groupi_n_3076, csa_tree_add_7_25_groupi_n_3077;
  wire csa_tree_add_7_25_groupi_n_3078, csa_tree_add_7_25_groupi_n_3079, csa_tree_add_7_25_groupi_n_3080, csa_tree_add_7_25_groupi_n_3081, csa_tree_add_7_25_groupi_n_3082, csa_tree_add_7_25_groupi_n_3083, csa_tree_add_7_25_groupi_n_3084, csa_tree_add_7_25_groupi_n_3085;
  wire csa_tree_add_7_25_groupi_n_3086, csa_tree_add_7_25_groupi_n_3087, csa_tree_add_7_25_groupi_n_3088, csa_tree_add_7_25_groupi_n_3089, csa_tree_add_7_25_groupi_n_3090, csa_tree_add_7_25_groupi_n_3091, csa_tree_add_7_25_groupi_n_3092, csa_tree_add_7_25_groupi_n_3093;
  wire csa_tree_add_7_25_groupi_n_3094, csa_tree_add_7_25_groupi_n_3095, csa_tree_add_7_25_groupi_n_3096, csa_tree_add_7_25_groupi_n_3097, csa_tree_add_7_25_groupi_n_3098, csa_tree_add_7_25_groupi_n_3099, csa_tree_add_7_25_groupi_n_3100, csa_tree_add_7_25_groupi_n_3101;
  wire csa_tree_add_7_25_groupi_n_3102, csa_tree_add_7_25_groupi_n_3103, csa_tree_add_7_25_groupi_n_3104, csa_tree_add_7_25_groupi_n_3105, csa_tree_add_7_25_groupi_n_3106, csa_tree_add_7_25_groupi_n_3107, csa_tree_add_7_25_groupi_n_3108, csa_tree_add_7_25_groupi_n_3109;
  wire csa_tree_add_7_25_groupi_n_3110, csa_tree_add_7_25_groupi_n_3111, csa_tree_add_7_25_groupi_n_3112, csa_tree_add_7_25_groupi_n_3113, csa_tree_add_7_25_groupi_n_3114, csa_tree_add_7_25_groupi_n_3115, csa_tree_add_7_25_groupi_n_3116, csa_tree_add_7_25_groupi_n_3117;
  wire csa_tree_add_7_25_groupi_n_3118, csa_tree_add_7_25_groupi_n_3119, csa_tree_add_7_25_groupi_n_3120, csa_tree_add_7_25_groupi_n_3121, csa_tree_add_7_25_groupi_n_3122, csa_tree_add_7_25_groupi_n_3123, csa_tree_add_7_25_groupi_n_3124, csa_tree_add_7_25_groupi_n_3125;
  wire csa_tree_add_7_25_groupi_n_3126, csa_tree_add_7_25_groupi_n_3127, csa_tree_add_7_25_groupi_n_3128, csa_tree_add_7_25_groupi_n_3129, csa_tree_add_7_25_groupi_n_3130, csa_tree_add_7_25_groupi_n_3131, csa_tree_add_7_25_groupi_n_3132, csa_tree_add_7_25_groupi_n_3133;
  wire csa_tree_add_7_25_groupi_n_3134, csa_tree_add_7_25_groupi_n_3135, csa_tree_add_7_25_groupi_n_3136, csa_tree_add_7_25_groupi_n_3137, csa_tree_add_7_25_groupi_n_3138, csa_tree_add_7_25_groupi_n_3139, csa_tree_add_7_25_groupi_n_3140, csa_tree_add_7_25_groupi_n_3141;
  wire csa_tree_add_7_25_groupi_n_3142, csa_tree_add_7_25_groupi_n_3143, csa_tree_add_7_25_groupi_n_3144, csa_tree_add_7_25_groupi_n_3145, csa_tree_add_7_25_groupi_n_3146, csa_tree_add_7_25_groupi_n_3147, csa_tree_add_7_25_groupi_n_3148, csa_tree_add_7_25_groupi_n_3149;
  wire csa_tree_add_7_25_groupi_n_3150, csa_tree_add_7_25_groupi_n_3151, csa_tree_add_7_25_groupi_n_3152, csa_tree_add_7_25_groupi_n_3153, csa_tree_add_7_25_groupi_n_3154, csa_tree_add_7_25_groupi_n_3155, csa_tree_add_7_25_groupi_n_3156, csa_tree_add_7_25_groupi_n_3157;
  wire csa_tree_add_7_25_groupi_n_3158, csa_tree_add_7_25_groupi_n_3159, csa_tree_add_7_25_groupi_n_3160, csa_tree_add_7_25_groupi_n_3161, csa_tree_add_7_25_groupi_n_3162, csa_tree_add_7_25_groupi_n_3163, csa_tree_add_7_25_groupi_n_3164, csa_tree_add_7_25_groupi_n_3165;
  wire csa_tree_add_7_25_groupi_n_3166, csa_tree_add_7_25_groupi_n_3167, csa_tree_add_7_25_groupi_n_3168, csa_tree_add_7_25_groupi_n_3169, csa_tree_add_7_25_groupi_n_3170, csa_tree_add_7_25_groupi_n_3171, csa_tree_add_7_25_groupi_n_3172, csa_tree_add_7_25_groupi_n_3173;
  wire csa_tree_add_7_25_groupi_n_3174, csa_tree_add_7_25_groupi_n_3175, csa_tree_add_7_25_groupi_n_3176, csa_tree_add_7_25_groupi_n_3177, csa_tree_add_7_25_groupi_n_3178, csa_tree_add_7_25_groupi_n_3179, csa_tree_add_7_25_groupi_n_3180, csa_tree_add_7_25_groupi_n_3181;
  wire csa_tree_add_7_25_groupi_n_3182, csa_tree_add_7_25_groupi_n_3183, csa_tree_add_7_25_groupi_n_3184, csa_tree_add_7_25_groupi_n_3185, csa_tree_add_7_25_groupi_n_3186, csa_tree_add_7_25_groupi_n_3187, csa_tree_add_7_25_groupi_n_3188, csa_tree_add_7_25_groupi_n_3189;
  wire csa_tree_add_7_25_groupi_n_3190, csa_tree_add_7_25_groupi_n_3191, csa_tree_add_7_25_groupi_n_3192, csa_tree_add_7_25_groupi_n_3193, csa_tree_add_7_25_groupi_n_3194, csa_tree_add_7_25_groupi_n_3195, csa_tree_add_7_25_groupi_n_3196, csa_tree_add_7_25_groupi_n_3197;
  wire csa_tree_add_7_25_groupi_n_3198, csa_tree_add_7_25_groupi_n_3199, csa_tree_add_7_25_groupi_n_3200, csa_tree_add_7_25_groupi_n_3201, csa_tree_add_7_25_groupi_n_3202, csa_tree_add_7_25_groupi_n_3203, csa_tree_add_7_25_groupi_n_3204, csa_tree_add_7_25_groupi_n_3205;
  wire csa_tree_add_7_25_groupi_n_3206, csa_tree_add_7_25_groupi_n_3207, csa_tree_add_7_25_groupi_n_3208, csa_tree_add_7_25_groupi_n_3209, csa_tree_add_7_25_groupi_n_3210, csa_tree_add_7_25_groupi_n_3211, csa_tree_add_7_25_groupi_n_3212, csa_tree_add_7_25_groupi_n_3213;
  wire csa_tree_add_7_25_groupi_n_3214, csa_tree_add_7_25_groupi_n_3215, csa_tree_add_7_25_groupi_n_3216, csa_tree_add_7_25_groupi_n_3217, csa_tree_add_7_25_groupi_n_3218, csa_tree_add_7_25_groupi_n_3219, csa_tree_add_7_25_groupi_n_3220, csa_tree_add_7_25_groupi_n_3221;
  wire csa_tree_add_7_25_groupi_n_3222, csa_tree_add_7_25_groupi_n_3223, csa_tree_add_7_25_groupi_n_3224, csa_tree_add_7_25_groupi_n_3225, csa_tree_add_7_25_groupi_n_3226, csa_tree_add_7_25_groupi_n_3227, csa_tree_add_7_25_groupi_n_3228, csa_tree_add_7_25_groupi_n_3229;
  wire csa_tree_add_7_25_groupi_n_3230, csa_tree_add_7_25_groupi_n_3231, csa_tree_add_7_25_groupi_n_3232, csa_tree_add_7_25_groupi_n_3233, csa_tree_add_7_25_groupi_n_3234, csa_tree_add_7_25_groupi_n_3235, csa_tree_add_7_25_groupi_n_3236, csa_tree_add_7_25_groupi_n_3237;
  wire csa_tree_add_7_25_groupi_n_3238, csa_tree_add_7_25_groupi_n_3239, csa_tree_add_7_25_groupi_n_3240, csa_tree_add_7_25_groupi_n_3241, csa_tree_add_7_25_groupi_n_3242, csa_tree_add_7_25_groupi_n_3243, csa_tree_add_7_25_groupi_n_3244, csa_tree_add_7_25_groupi_n_3245;
  wire csa_tree_add_7_25_groupi_n_3246, csa_tree_add_7_25_groupi_n_3247, csa_tree_add_7_25_groupi_n_3248, csa_tree_add_7_25_groupi_n_3249, csa_tree_add_7_25_groupi_n_3250, csa_tree_add_7_25_groupi_n_3251, csa_tree_add_7_25_groupi_n_3252, csa_tree_add_7_25_groupi_n_3253;
  wire csa_tree_add_7_25_groupi_n_3254, csa_tree_add_7_25_groupi_n_3255, csa_tree_add_7_25_groupi_n_3256, csa_tree_add_7_25_groupi_n_3257, csa_tree_add_7_25_groupi_n_3258, csa_tree_add_7_25_groupi_n_3259, csa_tree_add_7_25_groupi_n_3260, csa_tree_add_7_25_groupi_n_3261;
  wire csa_tree_add_7_25_groupi_n_3262, csa_tree_add_7_25_groupi_n_3263, csa_tree_add_7_25_groupi_n_3264, csa_tree_add_7_25_groupi_n_3265, csa_tree_add_7_25_groupi_n_3266, csa_tree_add_7_25_groupi_n_3267, csa_tree_add_7_25_groupi_n_3268, csa_tree_add_7_25_groupi_n_3269;
  wire csa_tree_add_7_25_groupi_n_3270, csa_tree_add_7_25_groupi_n_3271, csa_tree_add_7_25_groupi_n_3272, csa_tree_add_7_25_groupi_n_3273, csa_tree_add_7_25_groupi_n_3274, csa_tree_add_7_25_groupi_n_3275, csa_tree_add_7_25_groupi_n_3276, csa_tree_add_7_25_groupi_n_3277;
  wire csa_tree_add_7_25_groupi_n_3278, csa_tree_add_7_25_groupi_n_3279, csa_tree_add_7_25_groupi_n_3280, csa_tree_add_7_25_groupi_n_3281, csa_tree_add_7_25_groupi_n_3282, csa_tree_add_7_25_groupi_n_3283, csa_tree_add_7_25_groupi_n_3284, csa_tree_add_7_25_groupi_n_3285;
  wire csa_tree_add_7_25_groupi_n_3286, csa_tree_add_7_25_groupi_n_3287, csa_tree_add_7_25_groupi_n_3288, csa_tree_add_7_25_groupi_n_3289, csa_tree_add_7_25_groupi_n_3290, csa_tree_add_7_25_groupi_n_3291, csa_tree_add_7_25_groupi_n_3292, csa_tree_add_7_25_groupi_n_3293;
  wire csa_tree_add_7_25_groupi_n_3294, csa_tree_add_7_25_groupi_n_3295, csa_tree_add_7_25_groupi_n_3296, csa_tree_add_7_25_groupi_n_3297, csa_tree_add_7_25_groupi_n_3298, csa_tree_add_7_25_groupi_n_3299, csa_tree_add_7_25_groupi_n_3300, csa_tree_add_7_25_groupi_n_3301;
  wire csa_tree_add_7_25_groupi_n_3302, csa_tree_add_7_25_groupi_n_3303, csa_tree_add_7_25_groupi_n_3304, csa_tree_add_7_25_groupi_n_3305, csa_tree_add_7_25_groupi_n_3306, csa_tree_add_7_25_groupi_n_3307, csa_tree_add_7_25_groupi_n_3308, csa_tree_add_7_25_groupi_n_3309;
  wire csa_tree_add_7_25_groupi_n_3310, csa_tree_add_7_25_groupi_n_3311, csa_tree_add_7_25_groupi_n_3312, csa_tree_add_7_25_groupi_n_3313, csa_tree_add_7_25_groupi_n_3314, csa_tree_add_7_25_groupi_n_3315, csa_tree_add_7_25_groupi_n_3316, csa_tree_add_7_25_groupi_n_3317;
  wire csa_tree_add_7_25_groupi_n_3318, csa_tree_add_7_25_groupi_n_3319, csa_tree_add_7_25_groupi_n_3320, csa_tree_add_7_25_groupi_n_3321, csa_tree_add_7_25_groupi_n_3322, csa_tree_add_7_25_groupi_n_3323, csa_tree_add_7_25_groupi_n_3324, csa_tree_add_7_25_groupi_n_3325;
  wire csa_tree_add_7_25_groupi_n_3326, csa_tree_add_7_25_groupi_n_3327, csa_tree_add_7_25_groupi_n_3328, csa_tree_add_7_25_groupi_n_3329, csa_tree_add_7_25_groupi_n_3330, csa_tree_add_7_25_groupi_n_3331, csa_tree_add_7_25_groupi_n_3332, csa_tree_add_7_25_groupi_n_3333;
  wire csa_tree_add_7_25_groupi_n_3334, csa_tree_add_7_25_groupi_n_3335, csa_tree_add_7_25_groupi_n_3336, csa_tree_add_7_25_groupi_n_3337, csa_tree_add_7_25_groupi_n_3338, csa_tree_add_7_25_groupi_n_3339, csa_tree_add_7_25_groupi_n_3340, csa_tree_add_7_25_groupi_n_3341;
  wire csa_tree_add_7_25_groupi_n_3342, csa_tree_add_7_25_groupi_n_3343, csa_tree_add_7_25_groupi_n_3344, csa_tree_add_7_25_groupi_n_3345, csa_tree_add_7_25_groupi_n_3346, csa_tree_add_7_25_groupi_n_3347, csa_tree_add_7_25_groupi_n_3348, csa_tree_add_7_25_groupi_n_3349;
  wire csa_tree_add_7_25_groupi_n_3350, csa_tree_add_7_25_groupi_n_3351, csa_tree_add_7_25_groupi_n_3352, csa_tree_add_7_25_groupi_n_3353, csa_tree_add_7_25_groupi_n_3354, csa_tree_add_7_25_groupi_n_3355, csa_tree_add_7_25_groupi_n_3356, csa_tree_add_7_25_groupi_n_3357;
  wire csa_tree_add_7_25_groupi_n_3358, csa_tree_add_7_25_groupi_n_3359, csa_tree_add_7_25_groupi_n_3360, csa_tree_add_7_25_groupi_n_3361, csa_tree_add_7_25_groupi_n_3362, csa_tree_add_7_25_groupi_n_3363, csa_tree_add_7_25_groupi_n_3364, csa_tree_add_7_25_groupi_n_3365;
  wire csa_tree_add_7_25_groupi_n_3366, csa_tree_add_7_25_groupi_n_3367, csa_tree_add_7_25_groupi_n_3368, csa_tree_add_7_25_groupi_n_3369, csa_tree_add_7_25_groupi_n_3370, csa_tree_add_7_25_groupi_n_3371, csa_tree_add_7_25_groupi_n_3372, csa_tree_add_7_25_groupi_n_3373;
  wire csa_tree_add_7_25_groupi_n_3374, csa_tree_add_7_25_groupi_n_3375, csa_tree_add_7_25_groupi_n_3376, csa_tree_add_7_25_groupi_n_3377, csa_tree_add_7_25_groupi_n_3378, csa_tree_add_7_25_groupi_n_3379, csa_tree_add_7_25_groupi_n_3380, csa_tree_add_7_25_groupi_n_3381;
  wire csa_tree_add_7_25_groupi_n_3382, csa_tree_add_7_25_groupi_n_3383, csa_tree_add_7_25_groupi_n_3384, csa_tree_add_7_25_groupi_n_3385, csa_tree_add_7_25_groupi_n_3386, csa_tree_add_7_25_groupi_n_3387, csa_tree_add_7_25_groupi_n_3388, csa_tree_add_7_25_groupi_n_3389;
  wire csa_tree_add_7_25_groupi_n_3390, csa_tree_add_7_25_groupi_n_3391, csa_tree_add_7_25_groupi_n_3392, csa_tree_add_7_25_groupi_n_3393, csa_tree_add_7_25_groupi_n_3394, csa_tree_add_7_25_groupi_n_3395, csa_tree_add_7_25_groupi_n_3396, csa_tree_add_7_25_groupi_n_3397;
  wire csa_tree_add_7_25_groupi_n_3398, csa_tree_add_7_25_groupi_n_3399, csa_tree_add_7_25_groupi_n_3400, csa_tree_add_7_25_groupi_n_3401, csa_tree_add_7_25_groupi_n_3402, csa_tree_add_7_25_groupi_n_3403, csa_tree_add_7_25_groupi_n_3404, csa_tree_add_7_25_groupi_n_3405;
  wire csa_tree_add_7_25_groupi_n_3406, csa_tree_add_7_25_groupi_n_3407, csa_tree_add_7_25_groupi_n_3408, csa_tree_add_7_25_groupi_n_3409, csa_tree_add_7_25_groupi_n_3410, csa_tree_add_7_25_groupi_n_3411, csa_tree_add_7_25_groupi_n_3412, csa_tree_add_7_25_groupi_n_3413;
  wire csa_tree_add_7_25_groupi_n_3414, csa_tree_add_7_25_groupi_n_3415, csa_tree_add_7_25_groupi_n_3416, csa_tree_add_7_25_groupi_n_3417, csa_tree_add_7_25_groupi_n_3418, csa_tree_add_7_25_groupi_n_3419, csa_tree_add_7_25_groupi_n_3420, csa_tree_add_7_25_groupi_n_3421;
  wire csa_tree_add_7_25_groupi_n_3422, csa_tree_add_7_25_groupi_n_3423, csa_tree_add_7_25_groupi_n_3424, csa_tree_add_7_25_groupi_n_3425, csa_tree_add_7_25_groupi_n_3426, csa_tree_add_7_25_groupi_n_3427, csa_tree_add_7_25_groupi_n_3428, csa_tree_add_7_25_groupi_n_3429;
  wire csa_tree_add_7_25_groupi_n_3430, csa_tree_add_7_25_groupi_n_3431, csa_tree_add_7_25_groupi_n_3432, csa_tree_add_7_25_groupi_n_3433, csa_tree_add_7_25_groupi_n_3434, csa_tree_add_7_25_groupi_n_3435, csa_tree_add_7_25_groupi_n_3436, csa_tree_add_7_25_groupi_n_3437;
  wire csa_tree_add_7_25_groupi_n_3438, csa_tree_add_7_25_groupi_n_3439, csa_tree_add_7_25_groupi_n_3440, csa_tree_add_7_25_groupi_n_3441, csa_tree_add_7_25_groupi_n_3442, csa_tree_add_7_25_groupi_n_3443, csa_tree_add_7_25_groupi_n_3444, csa_tree_add_7_25_groupi_n_3445;
  wire csa_tree_add_7_25_groupi_n_3446, csa_tree_add_7_25_groupi_n_3447, csa_tree_add_7_25_groupi_n_3448, csa_tree_add_7_25_groupi_n_3449, csa_tree_add_7_25_groupi_n_3450, csa_tree_add_7_25_groupi_n_3451, csa_tree_add_7_25_groupi_n_3452, csa_tree_add_7_25_groupi_n_3453;
  wire csa_tree_add_7_25_groupi_n_3454, csa_tree_add_7_25_groupi_n_3455, csa_tree_add_7_25_groupi_n_3456, csa_tree_add_7_25_groupi_n_3457, csa_tree_add_7_25_groupi_n_3458, csa_tree_add_7_25_groupi_n_3459, csa_tree_add_7_25_groupi_n_3460, csa_tree_add_7_25_groupi_n_3461;
  wire csa_tree_add_7_25_groupi_n_3462, csa_tree_add_7_25_groupi_n_3463, csa_tree_add_7_25_groupi_n_3464, csa_tree_add_7_25_groupi_n_3465, csa_tree_add_7_25_groupi_n_3466, csa_tree_add_7_25_groupi_n_3467, csa_tree_add_7_25_groupi_n_3468, csa_tree_add_7_25_groupi_n_3469;
  wire csa_tree_add_7_25_groupi_n_3470, csa_tree_add_7_25_groupi_n_3471, csa_tree_add_7_25_groupi_n_3472, csa_tree_add_7_25_groupi_n_3473, csa_tree_add_7_25_groupi_n_3474, csa_tree_add_7_25_groupi_n_3475, csa_tree_add_7_25_groupi_n_3476, csa_tree_add_7_25_groupi_n_3477;
  wire csa_tree_add_7_25_groupi_n_3478, csa_tree_add_7_25_groupi_n_3479, csa_tree_add_7_25_groupi_n_3480, csa_tree_add_7_25_groupi_n_3481, csa_tree_add_7_25_groupi_n_3482, csa_tree_add_7_25_groupi_n_3483, csa_tree_add_7_25_groupi_n_3484, csa_tree_add_7_25_groupi_n_3485;
  wire csa_tree_add_7_25_groupi_n_3486, csa_tree_add_7_25_groupi_n_3487, csa_tree_add_7_25_groupi_n_3488, csa_tree_add_7_25_groupi_n_3489, csa_tree_add_7_25_groupi_n_3490, csa_tree_add_7_25_groupi_n_3491, csa_tree_add_7_25_groupi_n_3492, csa_tree_add_7_25_groupi_n_3493;
  wire csa_tree_add_7_25_groupi_n_3494, csa_tree_add_7_25_groupi_n_3495, csa_tree_add_7_25_groupi_n_3496, csa_tree_add_7_25_groupi_n_3497, csa_tree_add_7_25_groupi_n_3498, csa_tree_add_7_25_groupi_n_3499, csa_tree_add_7_25_groupi_n_3500, csa_tree_add_7_25_groupi_n_3501;
  wire csa_tree_add_7_25_groupi_n_3502, csa_tree_add_7_25_groupi_n_3503, csa_tree_add_7_25_groupi_n_3504, csa_tree_add_7_25_groupi_n_3505, csa_tree_add_7_25_groupi_n_3506, csa_tree_add_7_25_groupi_n_3507, csa_tree_add_7_25_groupi_n_3508, csa_tree_add_7_25_groupi_n_3509;
  wire csa_tree_add_7_25_groupi_n_3510, csa_tree_add_7_25_groupi_n_3511, csa_tree_add_7_25_groupi_n_3512, csa_tree_add_7_25_groupi_n_3513, csa_tree_add_7_25_groupi_n_3514, csa_tree_add_7_25_groupi_n_3515, csa_tree_add_7_25_groupi_n_3516, csa_tree_add_7_25_groupi_n_3517;
  wire csa_tree_add_7_25_groupi_n_3518, csa_tree_add_7_25_groupi_n_3519, csa_tree_add_7_25_groupi_n_3520, csa_tree_add_7_25_groupi_n_3521, csa_tree_add_7_25_groupi_n_3522, csa_tree_add_7_25_groupi_n_3523, csa_tree_add_7_25_groupi_n_3524, csa_tree_add_7_25_groupi_n_3525;
  wire csa_tree_add_7_25_groupi_n_3526, csa_tree_add_7_25_groupi_n_3527, csa_tree_add_7_25_groupi_n_3528, csa_tree_add_7_25_groupi_n_3529, csa_tree_add_7_25_groupi_n_3530, csa_tree_add_7_25_groupi_n_3531, csa_tree_add_7_25_groupi_n_3532, csa_tree_add_7_25_groupi_n_3533;
  wire csa_tree_add_7_25_groupi_n_3534, csa_tree_add_7_25_groupi_n_3535, csa_tree_add_7_25_groupi_n_3536, csa_tree_add_7_25_groupi_n_3537, csa_tree_add_7_25_groupi_n_3538, csa_tree_add_7_25_groupi_n_3539, csa_tree_add_7_25_groupi_n_3540, csa_tree_add_7_25_groupi_n_3541;
  wire csa_tree_add_7_25_groupi_n_3542, csa_tree_add_7_25_groupi_n_3543, csa_tree_add_7_25_groupi_n_3544, csa_tree_add_7_25_groupi_n_3545, csa_tree_add_7_25_groupi_n_3546, csa_tree_add_7_25_groupi_n_3547, csa_tree_add_7_25_groupi_n_3548, csa_tree_add_7_25_groupi_n_3549;
  wire csa_tree_add_7_25_groupi_n_3550, csa_tree_add_7_25_groupi_n_3551, csa_tree_add_7_25_groupi_n_3552, csa_tree_add_7_25_groupi_n_3553, csa_tree_add_7_25_groupi_n_3554, csa_tree_add_7_25_groupi_n_3555, csa_tree_add_7_25_groupi_n_3556, csa_tree_add_7_25_groupi_n_3557;
  wire csa_tree_add_7_25_groupi_n_3558, csa_tree_add_7_25_groupi_n_3559, csa_tree_add_7_25_groupi_n_3560, csa_tree_add_7_25_groupi_n_3561, csa_tree_add_7_25_groupi_n_3562, csa_tree_add_7_25_groupi_n_3563, csa_tree_add_7_25_groupi_n_3564, csa_tree_add_7_25_groupi_n_3565;
  wire csa_tree_add_7_25_groupi_n_3566, csa_tree_add_7_25_groupi_n_3567, csa_tree_add_7_25_groupi_n_3568, csa_tree_add_7_25_groupi_n_3569, csa_tree_add_7_25_groupi_n_3570, csa_tree_add_7_25_groupi_n_3571, csa_tree_add_7_25_groupi_n_3572, csa_tree_add_7_25_groupi_n_3573;
  wire csa_tree_add_7_25_groupi_n_3574, csa_tree_add_7_25_groupi_n_3575, csa_tree_add_7_25_groupi_n_3576, csa_tree_add_7_25_groupi_n_3577, csa_tree_add_7_25_groupi_n_3578, csa_tree_add_7_25_groupi_n_3579, csa_tree_add_7_25_groupi_n_3580, csa_tree_add_7_25_groupi_n_3581;
  wire csa_tree_add_7_25_groupi_n_3582, csa_tree_add_7_25_groupi_n_3583, csa_tree_add_7_25_groupi_n_3584, csa_tree_add_7_25_groupi_n_3585, csa_tree_add_7_25_groupi_n_3586, csa_tree_add_7_25_groupi_n_3587, csa_tree_add_7_25_groupi_n_3588, csa_tree_add_7_25_groupi_n_3589;
  wire csa_tree_add_7_25_groupi_n_3590, csa_tree_add_7_25_groupi_n_3591, csa_tree_add_7_25_groupi_n_3592, csa_tree_add_7_25_groupi_n_3593, csa_tree_add_7_25_groupi_n_3594, csa_tree_add_7_25_groupi_n_3595, csa_tree_add_7_25_groupi_n_3596, csa_tree_add_7_25_groupi_n_3597;
  wire csa_tree_add_7_25_groupi_n_3598, csa_tree_add_7_25_groupi_n_3599, csa_tree_add_7_25_groupi_n_3600, csa_tree_add_7_25_groupi_n_3601, csa_tree_add_7_25_groupi_n_3602, csa_tree_add_7_25_groupi_n_3603, csa_tree_add_7_25_groupi_n_3604, csa_tree_add_7_25_groupi_n_3605;
  wire csa_tree_add_7_25_groupi_n_3606, csa_tree_add_7_25_groupi_n_3607, csa_tree_add_7_25_groupi_n_3608, csa_tree_add_7_25_groupi_n_3609, csa_tree_add_7_25_groupi_n_3610, csa_tree_add_7_25_groupi_n_3611, csa_tree_add_7_25_groupi_n_3612, csa_tree_add_7_25_groupi_n_3613;
  wire csa_tree_add_7_25_groupi_n_3614, csa_tree_add_7_25_groupi_n_3615, csa_tree_add_7_25_groupi_n_3616, csa_tree_add_7_25_groupi_n_3617, csa_tree_add_7_25_groupi_n_3618, csa_tree_add_7_25_groupi_n_3619, csa_tree_add_7_25_groupi_n_3620, csa_tree_add_7_25_groupi_n_3621;
  wire csa_tree_add_7_25_groupi_n_3622, csa_tree_add_7_25_groupi_n_3623, csa_tree_add_7_25_groupi_n_3624, csa_tree_add_7_25_groupi_n_3625, csa_tree_add_7_25_groupi_n_3626, csa_tree_add_7_25_groupi_n_3627, csa_tree_add_7_25_groupi_n_3628, csa_tree_add_7_25_groupi_n_3629;
  wire csa_tree_add_7_25_groupi_n_3630, csa_tree_add_7_25_groupi_n_3631, csa_tree_add_7_25_groupi_n_3632, csa_tree_add_7_25_groupi_n_3633, csa_tree_add_7_25_groupi_n_3634, csa_tree_add_7_25_groupi_n_3635, csa_tree_add_7_25_groupi_n_3636, csa_tree_add_7_25_groupi_n_3637;
  wire csa_tree_add_7_25_groupi_n_3638, csa_tree_add_7_25_groupi_n_3639, csa_tree_add_7_25_groupi_n_3640, csa_tree_add_7_25_groupi_n_3641, csa_tree_add_7_25_groupi_n_3642, csa_tree_add_7_25_groupi_n_3643, csa_tree_add_7_25_groupi_n_3644, csa_tree_add_7_25_groupi_n_3645;
  wire csa_tree_add_7_25_groupi_n_3646, csa_tree_add_7_25_groupi_n_3647, csa_tree_add_7_25_groupi_n_3648, csa_tree_add_7_25_groupi_n_3649, csa_tree_add_7_25_groupi_n_3650, csa_tree_add_7_25_groupi_n_3651, csa_tree_add_7_25_groupi_n_3652, csa_tree_add_7_25_groupi_n_3653;
  wire csa_tree_add_7_25_groupi_n_3654, csa_tree_add_7_25_groupi_n_3655, csa_tree_add_7_25_groupi_n_3656, csa_tree_add_7_25_groupi_n_3657, csa_tree_add_7_25_groupi_n_3658, csa_tree_add_7_25_groupi_n_3659, csa_tree_add_7_25_groupi_n_3660, csa_tree_add_7_25_groupi_n_3661;
  wire csa_tree_add_7_25_groupi_n_3662, csa_tree_add_7_25_groupi_n_3663, csa_tree_add_7_25_groupi_n_3664, csa_tree_add_7_25_groupi_n_3665, csa_tree_add_7_25_groupi_n_3666, csa_tree_add_7_25_groupi_n_3667, csa_tree_add_7_25_groupi_n_3668, csa_tree_add_7_25_groupi_n_3669;
  wire csa_tree_add_7_25_groupi_n_3670, csa_tree_add_7_25_groupi_n_3671, csa_tree_add_7_25_groupi_n_3672, csa_tree_add_7_25_groupi_n_3673, csa_tree_add_7_25_groupi_n_3674, csa_tree_add_7_25_groupi_n_3675, csa_tree_add_7_25_groupi_n_3676, csa_tree_add_7_25_groupi_n_3677;
  wire csa_tree_add_7_25_groupi_n_3678, csa_tree_add_7_25_groupi_n_3679, csa_tree_add_7_25_groupi_n_3680, csa_tree_add_7_25_groupi_n_3681, csa_tree_add_7_25_groupi_n_3682, csa_tree_add_7_25_groupi_n_3683, csa_tree_add_7_25_groupi_n_3684, csa_tree_add_7_25_groupi_n_3685;
  wire csa_tree_add_7_25_groupi_n_3686, csa_tree_add_7_25_groupi_n_3687, csa_tree_add_7_25_groupi_n_3688, csa_tree_add_7_25_groupi_n_3689, csa_tree_add_7_25_groupi_n_3690, csa_tree_add_7_25_groupi_n_3691, csa_tree_add_7_25_groupi_n_3692, csa_tree_add_7_25_groupi_n_3693;
  wire csa_tree_add_7_25_groupi_n_3694, csa_tree_add_7_25_groupi_n_3695, csa_tree_add_7_25_groupi_n_3696, csa_tree_add_7_25_groupi_n_3697, csa_tree_add_7_25_groupi_n_3698, csa_tree_add_7_25_groupi_n_3699, csa_tree_add_7_25_groupi_n_3700, csa_tree_add_7_25_groupi_n_3701;
  wire csa_tree_add_7_25_groupi_n_3702, csa_tree_add_7_25_groupi_n_3703, csa_tree_add_7_25_groupi_n_3704, csa_tree_add_7_25_groupi_n_3705, csa_tree_add_7_25_groupi_n_3706, csa_tree_add_7_25_groupi_n_3707, csa_tree_add_7_25_groupi_n_3708, csa_tree_add_7_25_groupi_n_3709;
  wire csa_tree_add_7_25_groupi_n_3710, csa_tree_add_7_25_groupi_n_3711, csa_tree_add_7_25_groupi_n_3712, csa_tree_add_7_25_groupi_n_3713, csa_tree_add_7_25_groupi_n_3714, csa_tree_add_7_25_groupi_n_3715, csa_tree_add_7_25_groupi_n_3716, csa_tree_add_7_25_groupi_n_3717;
  wire csa_tree_add_7_25_groupi_n_3718, csa_tree_add_7_25_groupi_n_3719, csa_tree_add_7_25_groupi_n_3720, csa_tree_add_7_25_groupi_n_3721, csa_tree_add_7_25_groupi_n_3722, csa_tree_add_7_25_groupi_n_3723, csa_tree_add_7_25_groupi_n_3724, csa_tree_add_7_25_groupi_n_3725;
  wire csa_tree_add_7_25_groupi_n_3726, csa_tree_add_7_25_groupi_n_3727, csa_tree_add_7_25_groupi_n_3728, csa_tree_add_7_25_groupi_n_3729, csa_tree_add_7_25_groupi_n_3730, csa_tree_add_7_25_groupi_n_3731, csa_tree_add_7_25_groupi_n_3732, csa_tree_add_7_25_groupi_n_3733;
  wire csa_tree_add_7_25_groupi_n_3734, csa_tree_add_7_25_groupi_n_3735, csa_tree_add_7_25_groupi_n_3736, csa_tree_add_7_25_groupi_n_3737, csa_tree_add_7_25_groupi_n_3738, csa_tree_add_7_25_groupi_n_3739, csa_tree_add_7_25_groupi_n_3740, csa_tree_add_7_25_groupi_n_3741;
  wire csa_tree_add_7_25_groupi_n_3742, csa_tree_add_7_25_groupi_n_3743, csa_tree_add_7_25_groupi_n_3744, csa_tree_add_7_25_groupi_n_3745, csa_tree_add_7_25_groupi_n_3746, csa_tree_add_7_25_groupi_n_3747, csa_tree_add_7_25_groupi_n_3748, csa_tree_add_7_25_groupi_n_3749;
  wire csa_tree_add_7_25_groupi_n_3750, csa_tree_add_7_25_groupi_n_3751, csa_tree_add_7_25_groupi_n_3752, csa_tree_add_7_25_groupi_n_3753, csa_tree_add_7_25_groupi_n_3754, csa_tree_add_7_25_groupi_n_3755, csa_tree_add_7_25_groupi_n_3756, csa_tree_add_7_25_groupi_n_3757;
  wire csa_tree_add_7_25_groupi_n_3758, csa_tree_add_7_25_groupi_n_3759, csa_tree_add_7_25_groupi_n_3760, csa_tree_add_7_25_groupi_n_3761, csa_tree_add_7_25_groupi_n_3762, csa_tree_add_7_25_groupi_n_3763, csa_tree_add_7_25_groupi_n_3764, csa_tree_add_7_25_groupi_n_3765;
  wire csa_tree_add_7_25_groupi_n_3766, csa_tree_add_7_25_groupi_n_3767, csa_tree_add_7_25_groupi_n_3768, csa_tree_add_7_25_groupi_n_3769, csa_tree_add_7_25_groupi_n_3770, csa_tree_add_7_25_groupi_n_3771, csa_tree_add_7_25_groupi_n_3772, csa_tree_add_7_25_groupi_n_3773;
  wire csa_tree_add_7_25_groupi_n_3774, csa_tree_add_7_25_groupi_n_3775, csa_tree_add_7_25_groupi_n_3776, csa_tree_add_7_25_groupi_n_3777, csa_tree_add_7_25_groupi_n_3778, csa_tree_add_7_25_groupi_n_3779, csa_tree_add_7_25_groupi_n_3780, csa_tree_add_7_25_groupi_n_3781;
  wire csa_tree_add_7_25_groupi_n_3782, csa_tree_add_7_25_groupi_n_3783, csa_tree_add_7_25_groupi_n_3784, csa_tree_add_7_25_groupi_n_3785, csa_tree_add_7_25_groupi_n_3786, csa_tree_add_7_25_groupi_n_3787, csa_tree_add_7_25_groupi_n_3788, csa_tree_add_7_25_groupi_n_3789;
  wire csa_tree_add_7_25_groupi_n_3790, csa_tree_add_7_25_groupi_n_3791, csa_tree_add_7_25_groupi_n_3792, csa_tree_add_7_25_groupi_n_3793, csa_tree_add_7_25_groupi_n_3794, csa_tree_add_7_25_groupi_n_3795, csa_tree_add_7_25_groupi_n_3796, csa_tree_add_7_25_groupi_n_3797;
  wire csa_tree_add_7_25_groupi_n_3798, csa_tree_add_7_25_groupi_n_3799, csa_tree_add_7_25_groupi_n_3800, csa_tree_add_7_25_groupi_n_3801, csa_tree_add_7_25_groupi_n_3802, csa_tree_add_7_25_groupi_n_3803, csa_tree_add_7_25_groupi_n_3804, csa_tree_add_7_25_groupi_n_3805;
  wire csa_tree_add_7_25_groupi_n_3806, csa_tree_add_7_25_groupi_n_3807, csa_tree_add_7_25_groupi_n_3808, csa_tree_add_7_25_groupi_n_3809, csa_tree_add_7_25_groupi_n_3810, csa_tree_add_7_25_groupi_n_3811, csa_tree_add_7_25_groupi_n_3812, csa_tree_add_7_25_groupi_n_3813;
  wire csa_tree_add_7_25_groupi_n_3814, csa_tree_add_7_25_groupi_n_3815, csa_tree_add_7_25_groupi_n_3816, csa_tree_add_7_25_groupi_n_3817, csa_tree_add_7_25_groupi_n_3818, csa_tree_add_7_25_groupi_n_3819, csa_tree_add_7_25_groupi_n_3820, csa_tree_add_7_25_groupi_n_3821;
  wire csa_tree_add_7_25_groupi_n_3822, csa_tree_add_7_25_groupi_n_3823, csa_tree_add_7_25_groupi_n_3824, csa_tree_add_7_25_groupi_n_3825, csa_tree_add_7_25_groupi_n_3826, csa_tree_add_7_25_groupi_n_3827, csa_tree_add_7_25_groupi_n_3828, csa_tree_add_7_25_groupi_n_3829;
  wire csa_tree_add_7_25_groupi_n_3830, csa_tree_add_7_25_groupi_n_3831, csa_tree_add_7_25_groupi_n_3832, csa_tree_add_7_25_groupi_n_3833, csa_tree_add_7_25_groupi_n_3834, csa_tree_add_7_25_groupi_n_3835, csa_tree_add_7_25_groupi_n_3836, csa_tree_add_7_25_groupi_n_3837;
  wire csa_tree_add_7_25_groupi_n_3838, csa_tree_add_7_25_groupi_n_3839, csa_tree_add_7_25_groupi_n_3840, csa_tree_add_7_25_groupi_n_3841, csa_tree_add_7_25_groupi_n_3842, csa_tree_add_7_25_groupi_n_3843, csa_tree_add_7_25_groupi_n_3844, csa_tree_add_7_25_groupi_n_3845;
  wire csa_tree_add_7_25_groupi_n_3846, csa_tree_add_7_25_groupi_n_3847, csa_tree_add_7_25_groupi_n_3848, csa_tree_add_7_25_groupi_n_3849, csa_tree_add_7_25_groupi_n_3850, csa_tree_add_7_25_groupi_n_3851, csa_tree_add_7_25_groupi_n_3852, csa_tree_add_7_25_groupi_n_3853;
  wire csa_tree_add_7_25_groupi_n_3854, csa_tree_add_7_25_groupi_n_3855, csa_tree_add_7_25_groupi_n_3856, csa_tree_add_7_25_groupi_n_3857, csa_tree_add_7_25_groupi_n_3858, csa_tree_add_7_25_groupi_n_3859, csa_tree_add_7_25_groupi_n_3860, csa_tree_add_7_25_groupi_n_3861;
  wire csa_tree_add_7_25_groupi_n_3862, csa_tree_add_7_25_groupi_n_3863, csa_tree_add_7_25_groupi_n_3864, csa_tree_add_7_25_groupi_n_3865, csa_tree_add_7_25_groupi_n_3866, csa_tree_add_7_25_groupi_n_3867, csa_tree_add_7_25_groupi_n_3868, csa_tree_add_7_25_groupi_n_3869;
  wire csa_tree_add_7_25_groupi_n_3870, csa_tree_add_7_25_groupi_n_3871, csa_tree_add_7_25_groupi_n_3872, csa_tree_add_7_25_groupi_n_3873, csa_tree_add_7_25_groupi_n_3874, csa_tree_add_7_25_groupi_n_3875, csa_tree_add_7_25_groupi_n_3876, csa_tree_add_7_25_groupi_n_3877;
  wire csa_tree_add_7_25_groupi_n_3878, csa_tree_add_7_25_groupi_n_3879, csa_tree_add_7_25_groupi_n_3880, csa_tree_add_7_25_groupi_n_3881, csa_tree_add_7_25_groupi_n_3882, csa_tree_add_7_25_groupi_n_3883, csa_tree_add_7_25_groupi_n_3884, csa_tree_add_7_25_groupi_n_3885;
  wire csa_tree_add_7_25_groupi_n_3886, csa_tree_add_7_25_groupi_n_3887, csa_tree_add_7_25_groupi_n_3888, csa_tree_add_7_25_groupi_n_3889, csa_tree_add_7_25_groupi_n_3890, csa_tree_add_7_25_groupi_n_3891, csa_tree_add_7_25_groupi_n_3892, csa_tree_add_7_25_groupi_n_3893;
  wire csa_tree_add_7_25_groupi_n_3894, csa_tree_add_7_25_groupi_n_3895, csa_tree_add_7_25_groupi_n_3896, csa_tree_add_7_25_groupi_n_3897, csa_tree_add_7_25_groupi_n_3898, csa_tree_add_7_25_groupi_n_3899, csa_tree_add_7_25_groupi_n_3900, csa_tree_add_7_25_groupi_n_3901;
  wire csa_tree_add_7_25_groupi_n_3902, csa_tree_add_7_25_groupi_n_3903, csa_tree_add_7_25_groupi_n_3904, csa_tree_add_7_25_groupi_n_3905, csa_tree_add_7_25_groupi_n_3906, csa_tree_add_7_25_groupi_n_3907, csa_tree_add_7_25_groupi_n_3908, csa_tree_add_7_25_groupi_n_3909;
  wire csa_tree_add_7_25_groupi_n_3910, csa_tree_add_7_25_groupi_n_3911, csa_tree_add_7_25_groupi_n_3912, csa_tree_add_7_25_groupi_n_3913, csa_tree_add_7_25_groupi_n_3914, csa_tree_add_7_25_groupi_n_3915, csa_tree_add_7_25_groupi_n_3916, csa_tree_add_7_25_groupi_n_3917;
  wire csa_tree_add_7_25_groupi_n_3918, csa_tree_add_7_25_groupi_n_3919, csa_tree_add_7_25_groupi_n_3920, csa_tree_add_7_25_groupi_n_3921, csa_tree_add_7_25_groupi_n_3922, csa_tree_add_7_25_groupi_n_3923, csa_tree_add_7_25_groupi_n_3924, csa_tree_add_7_25_groupi_n_3925;
  wire csa_tree_add_7_25_groupi_n_3926, csa_tree_add_7_25_groupi_n_3927, csa_tree_add_7_25_groupi_n_3928, csa_tree_add_7_25_groupi_n_3929, csa_tree_add_7_25_groupi_n_3930, csa_tree_add_7_25_groupi_n_3931, csa_tree_add_7_25_groupi_n_3932, csa_tree_add_7_25_groupi_n_3933;
  wire csa_tree_add_7_25_groupi_n_3934, csa_tree_add_7_25_groupi_n_3935, csa_tree_add_7_25_groupi_n_3936, csa_tree_add_7_25_groupi_n_3937, csa_tree_add_7_25_groupi_n_3938, csa_tree_add_7_25_groupi_n_3939, csa_tree_add_7_25_groupi_n_3940, csa_tree_add_7_25_groupi_n_3941;
  wire csa_tree_add_7_25_groupi_n_3942, csa_tree_add_7_25_groupi_n_3943, csa_tree_add_7_25_groupi_n_3944, csa_tree_add_7_25_groupi_n_3945, csa_tree_add_7_25_groupi_n_3946, csa_tree_add_7_25_groupi_n_3947, csa_tree_add_7_25_groupi_n_3948, csa_tree_add_7_25_groupi_n_3949;
  wire csa_tree_add_7_25_groupi_n_3950, csa_tree_add_7_25_groupi_n_3951, csa_tree_add_7_25_groupi_n_3952, csa_tree_add_7_25_groupi_n_3953, csa_tree_add_7_25_groupi_n_3954, csa_tree_add_7_25_groupi_n_3955, csa_tree_add_7_25_groupi_n_3956, csa_tree_add_7_25_groupi_n_3957;
  wire csa_tree_add_7_25_groupi_n_3958, csa_tree_add_7_25_groupi_n_3959, csa_tree_add_7_25_groupi_n_3960, csa_tree_add_7_25_groupi_n_3961, csa_tree_add_7_25_groupi_n_3962, csa_tree_add_7_25_groupi_n_3963, csa_tree_add_7_25_groupi_n_3964, csa_tree_add_7_25_groupi_n_3965;
  wire csa_tree_add_7_25_groupi_n_3966, csa_tree_add_7_25_groupi_n_3967, csa_tree_add_7_25_groupi_n_3968, csa_tree_add_7_25_groupi_n_3969, csa_tree_add_7_25_groupi_n_3970, csa_tree_add_7_25_groupi_n_3971, csa_tree_add_7_25_groupi_n_3972, csa_tree_add_7_25_groupi_n_3973;
  wire csa_tree_add_7_25_groupi_n_3974, csa_tree_add_7_25_groupi_n_3975, csa_tree_add_7_25_groupi_n_3976, csa_tree_add_7_25_groupi_n_3977, csa_tree_add_7_25_groupi_n_3978, csa_tree_add_7_25_groupi_n_3979, csa_tree_add_7_25_groupi_n_3980, csa_tree_add_7_25_groupi_n_3981;
  wire csa_tree_add_7_25_groupi_n_3982, csa_tree_add_7_25_groupi_n_3983, csa_tree_add_7_25_groupi_n_3984, csa_tree_add_7_25_groupi_n_3985, csa_tree_add_7_25_groupi_n_3986, csa_tree_add_7_25_groupi_n_3987, csa_tree_add_7_25_groupi_n_3988, csa_tree_add_7_25_groupi_n_3989;
  wire csa_tree_add_7_25_groupi_n_3990, csa_tree_add_7_25_groupi_n_3991, csa_tree_add_7_25_groupi_n_3992, csa_tree_add_7_25_groupi_n_3993, csa_tree_add_7_25_groupi_n_3994, csa_tree_add_7_25_groupi_n_3995, csa_tree_add_7_25_groupi_n_3996, csa_tree_add_7_25_groupi_n_3997;
  wire csa_tree_add_7_25_groupi_n_3998, csa_tree_add_7_25_groupi_n_3999, csa_tree_add_7_25_groupi_n_4000, csa_tree_add_7_25_groupi_n_4001, csa_tree_add_7_25_groupi_n_4002, csa_tree_add_7_25_groupi_n_4003, csa_tree_add_7_25_groupi_n_4004, csa_tree_add_7_25_groupi_n_4005;
  wire csa_tree_add_7_25_groupi_n_4006, csa_tree_add_7_25_groupi_n_4007, csa_tree_add_7_25_groupi_n_4008, csa_tree_add_7_25_groupi_n_4009, csa_tree_add_7_25_groupi_n_4010, csa_tree_add_7_25_groupi_n_4011, csa_tree_add_7_25_groupi_n_4012, csa_tree_add_7_25_groupi_n_4013;
  wire csa_tree_add_7_25_groupi_n_4014, csa_tree_add_7_25_groupi_n_4015, csa_tree_add_7_25_groupi_n_4016, csa_tree_add_7_25_groupi_n_4017, csa_tree_add_7_25_groupi_n_4018, csa_tree_add_7_25_groupi_n_4019, csa_tree_add_7_25_groupi_n_4020, csa_tree_add_7_25_groupi_n_4021;
  wire csa_tree_add_7_25_groupi_n_4022, csa_tree_add_7_25_groupi_n_4023, csa_tree_add_7_25_groupi_n_4024, csa_tree_add_7_25_groupi_n_4025, csa_tree_add_7_25_groupi_n_4026, csa_tree_add_7_25_groupi_n_4027, csa_tree_add_7_25_groupi_n_4028, csa_tree_add_7_25_groupi_n_4029;
  wire csa_tree_add_7_25_groupi_n_4030, csa_tree_add_7_25_groupi_n_4031, csa_tree_add_7_25_groupi_n_4032, csa_tree_add_7_25_groupi_n_4033, csa_tree_add_7_25_groupi_n_4034, csa_tree_add_7_25_groupi_n_4035, csa_tree_add_7_25_groupi_n_4036, csa_tree_add_7_25_groupi_n_4037;
  wire csa_tree_add_7_25_groupi_n_4038, csa_tree_add_7_25_groupi_n_4039, csa_tree_add_7_25_groupi_n_4040, csa_tree_add_7_25_groupi_n_4041, csa_tree_add_7_25_groupi_n_4042, csa_tree_add_7_25_groupi_n_4043, csa_tree_add_7_25_groupi_n_4044, csa_tree_add_7_25_groupi_n_4045;
  wire csa_tree_add_7_25_groupi_n_4046, csa_tree_add_7_25_groupi_n_4047, csa_tree_add_7_25_groupi_n_4048, csa_tree_add_7_25_groupi_n_4049, csa_tree_add_7_25_groupi_n_4050, csa_tree_add_7_25_groupi_n_4051, csa_tree_add_7_25_groupi_n_4052, csa_tree_add_7_25_groupi_n_4053;
  wire csa_tree_add_7_25_groupi_n_4054, csa_tree_add_7_25_groupi_n_4055, csa_tree_add_7_25_groupi_n_4056, csa_tree_add_7_25_groupi_n_4057, csa_tree_add_7_25_groupi_n_4058, csa_tree_add_7_25_groupi_n_4059, csa_tree_add_7_25_groupi_n_4060, csa_tree_add_7_25_groupi_n_4061;
  wire csa_tree_add_7_25_groupi_n_4062, csa_tree_add_7_25_groupi_n_4063, csa_tree_add_7_25_groupi_n_4064, csa_tree_add_7_25_groupi_n_4065, csa_tree_add_7_25_groupi_n_4066, csa_tree_add_7_25_groupi_n_4067, csa_tree_add_7_25_groupi_n_4068, csa_tree_add_7_25_groupi_n_4069;
  wire csa_tree_add_7_25_groupi_n_4070, csa_tree_add_7_25_groupi_n_4071, csa_tree_add_7_25_groupi_n_4072, csa_tree_add_7_25_groupi_n_4073, csa_tree_add_7_25_groupi_n_4074, csa_tree_add_7_25_groupi_n_4075, csa_tree_add_7_25_groupi_n_4076, csa_tree_add_7_25_groupi_n_4077;
  wire csa_tree_add_7_25_groupi_n_4078, csa_tree_add_7_25_groupi_n_4079, csa_tree_add_7_25_groupi_n_4080, csa_tree_add_7_25_groupi_n_4081, csa_tree_add_7_25_groupi_n_4082, csa_tree_add_7_25_groupi_n_4083, csa_tree_add_7_25_groupi_n_4084, csa_tree_add_7_25_groupi_n_4085;
  wire csa_tree_add_7_25_groupi_n_4086, csa_tree_add_7_25_groupi_n_4087, csa_tree_add_7_25_groupi_n_4088, csa_tree_add_7_25_groupi_n_4089, csa_tree_add_7_25_groupi_n_4090, csa_tree_add_7_25_groupi_n_4091, csa_tree_add_7_25_groupi_n_4092, csa_tree_add_7_25_groupi_n_4093;
  wire csa_tree_add_7_25_groupi_n_4094, csa_tree_add_7_25_groupi_n_4095, csa_tree_add_7_25_groupi_n_4096, csa_tree_add_7_25_groupi_n_4097, csa_tree_add_7_25_groupi_n_4098, csa_tree_add_7_25_groupi_n_4099, csa_tree_add_7_25_groupi_n_4100, csa_tree_add_7_25_groupi_n_4101;
  wire csa_tree_add_7_25_groupi_n_4102, csa_tree_add_7_25_groupi_n_4103, csa_tree_add_7_25_groupi_n_4104, csa_tree_add_7_25_groupi_n_4105, csa_tree_add_7_25_groupi_n_4106, csa_tree_add_7_25_groupi_n_4107, csa_tree_add_7_25_groupi_n_4108, csa_tree_add_7_25_groupi_n_4109;
  wire csa_tree_add_7_25_groupi_n_4110, csa_tree_add_7_25_groupi_n_4111, csa_tree_add_7_25_groupi_n_4112, csa_tree_add_7_25_groupi_n_4113, csa_tree_add_7_25_groupi_n_4114, csa_tree_add_7_25_groupi_n_4115, csa_tree_add_7_25_groupi_n_4116, csa_tree_add_7_25_groupi_n_4117;
  wire csa_tree_add_7_25_groupi_n_4118, csa_tree_add_7_25_groupi_n_4119, csa_tree_add_7_25_groupi_n_4120, csa_tree_add_7_25_groupi_n_4121, csa_tree_add_7_25_groupi_n_4122, csa_tree_add_7_25_groupi_n_4123, csa_tree_add_7_25_groupi_n_4124, csa_tree_add_7_25_groupi_n_4125;
  wire csa_tree_add_7_25_groupi_n_4126, csa_tree_add_7_25_groupi_n_4127, csa_tree_add_7_25_groupi_n_4128, csa_tree_add_7_25_groupi_n_4129, csa_tree_add_7_25_groupi_n_4130, csa_tree_add_7_25_groupi_n_4131, csa_tree_add_7_25_groupi_n_4132, csa_tree_add_7_25_groupi_n_4133;
  wire csa_tree_add_7_25_groupi_n_4134, csa_tree_add_7_25_groupi_n_4135, csa_tree_add_7_25_groupi_n_4136, csa_tree_add_7_25_groupi_n_4137, csa_tree_add_7_25_groupi_n_4138, csa_tree_add_7_25_groupi_n_4139, csa_tree_add_7_25_groupi_n_4140, csa_tree_add_7_25_groupi_n_4141;
  wire csa_tree_add_7_25_groupi_n_4142, csa_tree_add_7_25_groupi_n_4143, csa_tree_add_7_25_groupi_n_4144, csa_tree_add_7_25_groupi_n_4145, csa_tree_add_7_25_groupi_n_4146, csa_tree_add_7_25_groupi_n_4147, csa_tree_add_7_25_groupi_n_4148, csa_tree_add_7_25_groupi_n_4149;
  wire csa_tree_add_7_25_groupi_n_4150, csa_tree_add_7_25_groupi_n_4151, csa_tree_add_7_25_groupi_n_4152, csa_tree_add_7_25_groupi_n_4153, csa_tree_add_7_25_groupi_n_4154, csa_tree_add_7_25_groupi_n_4155, csa_tree_add_7_25_groupi_n_4156, csa_tree_add_7_25_groupi_n_4157;
  wire csa_tree_add_7_25_groupi_n_4158, csa_tree_add_7_25_groupi_n_4159, csa_tree_add_7_25_groupi_n_4160, csa_tree_add_7_25_groupi_n_4161, csa_tree_add_7_25_groupi_n_4162, csa_tree_add_7_25_groupi_n_4163, csa_tree_add_7_25_groupi_n_4164, csa_tree_add_7_25_groupi_n_4165;
  wire csa_tree_add_7_25_groupi_n_4166, csa_tree_add_7_25_groupi_n_4167, csa_tree_add_7_25_groupi_n_4168, csa_tree_add_7_25_groupi_n_4169, csa_tree_add_7_25_groupi_n_4170, csa_tree_add_7_25_groupi_n_4171, csa_tree_add_7_25_groupi_n_4172, csa_tree_add_7_25_groupi_n_4173;
  wire csa_tree_add_7_25_groupi_n_4174, csa_tree_add_7_25_groupi_n_4175, csa_tree_add_7_25_groupi_n_4176, csa_tree_add_7_25_groupi_n_4177, csa_tree_add_7_25_groupi_n_4178, csa_tree_add_7_25_groupi_n_4179, csa_tree_add_7_25_groupi_n_4180, csa_tree_add_7_25_groupi_n_4181;
  wire csa_tree_add_7_25_groupi_n_4182, csa_tree_add_7_25_groupi_n_4183, csa_tree_add_7_25_groupi_n_4184, csa_tree_add_7_25_groupi_n_4185, csa_tree_add_7_25_groupi_n_4186, csa_tree_add_7_25_groupi_n_4187, csa_tree_add_7_25_groupi_n_4188, csa_tree_add_7_25_groupi_n_4189;
  wire csa_tree_add_7_25_groupi_n_4190, csa_tree_add_7_25_groupi_n_4191, csa_tree_add_7_25_groupi_n_4192, csa_tree_add_7_25_groupi_n_4193, csa_tree_add_7_25_groupi_n_4194, csa_tree_add_7_25_groupi_n_4195, csa_tree_add_7_25_groupi_n_4196, csa_tree_add_7_25_groupi_n_4197;
  wire csa_tree_add_7_25_groupi_n_4198, csa_tree_add_7_25_groupi_n_4199, csa_tree_add_7_25_groupi_n_4200, csa_tree_add_7_25_groupi_n_4201, csa_tree_add_7_25_groupi_n_4202, csa_tree_add_7_25_groupi_n_4203, csa_tree_add_7_25_groupi_n_4204, csa_tree_add_7_25_groupi_n_4205;
  wire csa_tree_add_7_25_groupi_n_4206, csa_tree_add_7_25_groupi_n_4207, csa_tree_add_7_25_groupi_n_4208, csa_tree_add_7_25_groupi_n_4209, csa_tree_add_7_25_groupi_n_4210, csa_tree_add_7_25_groupi_n_4211, csa_tree_add_7_25_groupi_n_4212, csa_tree_add_7_25_groupi_n_4213;
  wire csa_tree_add_7_25_groupi_n_4214, csa_tree_add_7_25_groupi_n_4215, csa_tree_add_7_25_groupi_n_4216, csa_tree_add_7_25_groupi_n_4217, csa_tree_add_7_25_groupi_n_4218, csa_tree_add_7_25_groupi_n_4219, csa_tree_add_7_25_groupi_n_4220, csa_tree_add_7_25_groupi_n_4221;
  wire csa_tree_add_7_25_groupi_n_4222, csa_tree_add_7_25_groupi_n_4223, csa_tree_add_7_25_groupi_n_4224, csa_tree_add_7_25_groupi_n_4225, csa_tree_add_7_25_groupi_n_4226, csa_tree_add_7_25_groupi_n_4227, csa_tree_add_7_25_groupi_n_4228, csa_tree_add_7_25_groupi_n_4229;
  wire csa_tree_add_7_25_groupi_n_4230, csa_tree_add_7_25_groupi_n_4231, csa_tree_add_7_25_groupi_n_4232, csa_tree_add_7_25_groupi_n_4233, csa_tree_add_7_25_groupi_n_4234, csa_tree_add_7_25_groupi_n_4235, csa_tree_add_7_25_groupi_n_4236, csa_tree_add_7_25_groupi_n_4237;
  wire csa_tree_add_7_25_groupi_n_4238, csa_tree_add_7_25_groupi_n_4239, csa_tree_add_7_25_groupi_n_4240, csa_tree_add_7_25_groupi_n_4241, csa_tree_add_7_25_groupi_n_4242, csa_tree_add_7_25_groupi_n_4243, csa_tree_add_7_25_groupi_n_4244, csa_tree_add_7_25_groupi_n_4245;
  wire csa_tree_add_7_25_groupi_n_4246, csa_tree_add_7_25_groupi_n_4247, csa_tree_add_7_25_groupi_n_4248, csa_tree_add_7_25_groupi_n_4249, csa_tree_add_7_25_groupi_n_4250, csa_tree_add_7_25_groupi_n_4251, csa_tree_add_7_25_groupi_n_4252, csa_tree_add_7_25_groupi_n_4253;
  wire csa_tree_add_7_25_groupi_n_4254, csa_tree_add_7_25_groupi_n_4255, csa_tree_add_7_25_groupi_n_4256, csa_tree_add_7_25_groupi_n_4257, csa_tree_add_7_25_groupi_n_4258, csa_tree_add_7_25_groupi_n_4259, csa_tree_add_7_25_groupi_n_4260, csa_tree_add_7_25_groupi_n_4261;
  wire csa_tree_add_7_25_groupi_n_4262, csa_tree_add_7_25_groupi_n_4263, csa_tree_add_7_25_groupi_n_4264, csa_tree_add_7_25_groupi_n_4265, csa_tree_add_7_25_groupi_n_4266, csa_tree_add_7_25_groupi_n_4267, csa_tree_add_7_25_groupi_n_4268, csa_tree_add_7_25_groupi_n_4269;
  wire csa_tree_add_7_25_groupi_n_4270, csa_tree_add_7_25_groupi_n_4271, csa_tree_add_7_25_groupi_n_4272, csa_tree_add_7_25_groupi_n_4273, csa_tree_add_7_25_groupi_n_4274, csa_tree_add_7_25_groupi_n_4275, csa_tree_add_7_25_groupi_n_4276, csa_tree_add_7_25_groupi_n_4277;
  wire csa_tree_add_7_25_groupi_n_4278, csa_tree_add_7_25_groupi_n_4279, csa_tree_add_7_25_groupi_n_4280, csa_tree_add_7_25_groupi_n_4281, csa_tree_add_7_25_groupi_n_4282, csa_tree_add_7_25_groupi_n_4283, csa_tree_add_7_25_groupi_n_4284, csa_tree_add_7_25_groupi_n_4285;
  wire csa_tree_add_7_25_groupi_n_4286, csa_tree_add_7_25_groupi_n_4287, csa_tree_add_7_25_groupi_n_4288, csa_tree_add_7_25_groupi_n_4289, csa_tree_add_7_25_groupi_n_4290, csa_tree_add_7_25_groupi_n_4291, csa_tree_add_7_25_groupi_n_4292, csa_tree_add_7_25_groupi_n_4293;
  wire csa_tree_add_7_25_groupi_n_4294, csa_tree_add_7_25_groupi_n_4295, csa_tree_add_7_25_groupi_n_4296, csa_tree_add_7_25_groupi_n_4297, csa_tree_add_7_25_groupi_n_4298, csa_tree_add_7_25_groupi_n_4299, csa_tree_add_7_25_groupi_n_4300, csa_tree_add_7_25_groupi_n_4301;
  wire csa_tree_add_7_25_groupi_n_4302, csa_tree_add_7_25_groupi_n_4303, csa_tree_add_7_25_groupi_n_4304, csa_tree_add_7_25_groupi_n_4305, csa_tree_add_7_25_groupi_n_4306, csa_tree_add_7_25_groupi_n_4307, csa_tree_add_7_25_groupi_n_4308, csa_tree_add_7_25_groupi_n_4309;
  wire csa_tree_add_7_25_groupi_n_4310, csa_tree_add_7_25_groupi_n_4311, csa_tree_add_7_25_groupi_n_4312, csa_tree_add_7_25_groupi_n_4313, csa_tree_add_7_25_groupi_n_4314, csa_tree_add_7_25_groupi_n_4315, csa_tree_add_7_25_groupi_n_4316, csa_tree_add_7_25_groupi_n_4317;
  wire csa_tree_add_7_25_groupi_n_4318, csa_tree_add_7_25_groupi_n_4319, csa_tree_add_7_25_groupi_n_4320, csa_tree_add_7_25_groupi_n_4321, csa_tree_add_7_25_groupi_n_4322, csa_tree_add_7_25_groupi_n_4323, csa_tree_add_7_25_groupi_n_4324, csa_tree_add_7_25_groupi_n_4325;
  wire csa_tree_add_7_25_groupi_n_4326, csa_tree_add_7_25_groupi_n_4327, csa_tree_add_7_25_groupi_n_4328, csa_tree_add_7_25_groupi_n_4329, csa_tree_add_7_25_groupi_n_4330, csa_tree_add_7_25_groupi_n_4331, csa_tree_add_7_25_groupi_n_4332, csa_tree_add_7_25_groupi_n_4333;
  wire csa_tree_add_7_25_groupi_n_4334, csa_tree_add_7_25_groupi_n_4335, csa_tree_add_7_25_groupi_n_4336, csa_tree_add_7_25_groupi_n_4337, csa_tree_add_7_25_groupi_n_4338, csa_tree_add_7_25_groupi_n_4339, csa_tree_add_7_25_groupi_n_4340, csa_tree_add_7_25_groupi_n_4341;
  wire csa_tree_add_7_25_groupi_n_4342, csa_tree_add_7_25_groupi_n_4343, csa_tree_add_7_25_groupi_n_4344, csa_tree_add_7_25_groupi_n_4345, csa_tree_add_7_25_groupi_n_4346, csa_tree_add_7_25_groupi_n_4347, csa_tree_add_7_25_groupi_n_4348, csa_tree_add_7_25_groupi_n_4349;
  wire csa_tree_add_7_25_groupi_n_4350, csa_tree_add_7_25_groupi_n_4351, csa_tree_add_7_25_groupi_n_4352, csa_tree_add_7_25_groupi_n_4353, csa_tree_add_7_25_groupi_n_4354, csa_tree_add_7_25_groupi_n_4355, csa_tree_add_7_25_groupi_n_4356, csa_tree_add_7_25_groupi_n_4357;
  wire csa_tree_add_7_25_groupi_n_4358, csa_tree_add_7_25_groupi_n_4359, csa_tree_add_7_25_groupi_n_4360, csa_tree_add_7_25_groupi_n_4361, csa_tree_add_7_25_groupi_n_4362, csa_tree_add_7_25_groupi_n_4363, csa_tree_add_7_25_groupi_n_4364, csa_tree_add_7_25_groupi_n_4365;
  wire csa_tree_add_7_25_groupi_n_4366, csa_tree_add_7_25_groupi_n_4367, csa_tree_add_7_25_groupi_n_4368, csa_tree_add_7_25_groupi_n_4369, csa_tree_add_7_25_groupi_n_4370, csa_tree_add_7_25_groupi_n_4371, csa_tree_add_7_25_groupi_n_4372, csa_tree_add_7_25_groupi_n_4373;
  wire csa_tree_add_7_25_groupi_n_4374, csa_tree_add_7_25_groupi_n_4375, csa_tree_add_7_25_groupi_n_4376, csa_tree_add_7_25_groupi_n_4377, csa_tree_add_7_25_groupi_n_4378, csa_tree_add_7_25_groupi_n_4379, csa_tree_add_7_25_groupi_n_4380, csa_tree_add_7_25_groupi_n_4381;
  wire csa_tree_add_7_25_groupi_n_4382, csa_tree_add_7_25_groupi_n_4383, csa_tree_add_7_25_groupi_n_4384, csa_tree_add_7_25_groupi_n_4385, csa_tree_add_7_25_groupi_n_4386, csa_tree_add_7_25_groupi_n_4387, csa_tree_add_7_25_groupi_n_4388, csa_tree_add_7_25_groupi_n_4389;
  wire csa_tree_add_7_25_groupi_n_4390, csa_tree_add_7_25_groupi_n_4391, csa_tree_add_7_25_groupi_n_4392, csa_tree_add_7_25_groupi_n_4393, csa_tree_add_7_25_groupi_n_4394, csa_tree_add_7_25_groupi_n_4395, csa_tree_add_7_25_groupi_n_4396, csa_tree_add_7_25_groupi_n_4397;
  wire csa_tree_add_7_25_groupi_n_4398, csa_tree_add_7_25_groupi_n_4399, csa_tree_add_7_25_groupi_n_4400, csa_tree_add_7_25_groupi_n_4401, csa_tree_add_7_25_groupi_n_4402, csa_tree_add_7_25_groupi_n_4403, csa_tree_add_7_25_groupi_n_4404, csa_tree_add_7_25_groupi_n_4405;
  wire csa_tree_add_7_25_groupi_n_4406, csa_tree_add_7_25_groupi_n_4407, csa_tree_add_7_25_groupi_n_4408, csa_tree_add_7_25_groupi_n_4409, csa_tree_add_7_25_groupi_n_4410, csa_tree_add_7_25_groupi_n_4411, csa_tree_add_7_25_groupi_n_4412, csa_tree_add_7_25_groupi_n_4413;
  wire csa_tree_add_7_25_groupi_n_4414, csa_tree_add_7_25_groupi_n_4415, csa_tree_add_7_25_groupi_n_4416, csa_tree_add_7_25_groupi_n_4417, csa_tree_add_7_25_groupi_n_4418, csa_tree_add_7_25_groupi_n_4419, csa_tree_add_7_25_groupi_n_4420, csa_tree_add_7_25_groupi_n_4421;
  wire csa_tree_add_7_25_groupi_n_4422, csa_tree_add_7_25_groupi_n_4423, csa_tree_add_7_25_groupi_n_4424, csa_tree_add_7_25_groupi_n_4425, csa_tree_add_7_25_groupi_n_4426, csa_tree_add_7_25_groupi_n_4427, csa_tree_add_7_25_groupi_n_4428, csa_tree_add_7_25_groupi_n_4429;
  wire csa_tree_add_7_25_groupi_n_4430, csa_tree_add_7_25_groupi_n_4431, csa_tree_add_7_25_groupi_n_4432, csa_tree_add_7_25_groupi_n_4433, csa_tree_add_7_25_groupi_n_4434, csa_tree_add_7_25_groupi_n_4435, csa_tree_add_7_25_groupi_n_4436, csa_tree_add_7_25_groupi_n_4437;
  wire csa_tree_add_7_25_groupi_n_4438, csa_tree_add_7_25_groupi_n_4439, csa_tree_add_7_25_groupi_n_4440, csa_tree_add_7_25_groupi_n_4441, csa_tree_add_7_25_groupi_n_4442, csa_tree_add_7_25_groupi_n_4443, csa_tree_add_7_25_groupi_n_4444, csa_tree_add_7_25_groupi_n_4445;
  wire csa_tree_add_7_25_groupi_n_4446, csa_tree_add_7_25_groupi_n_4447, csa_tree_add_7_25_groupi_n_4448, csa_tree_add_7_25_groupi_n_4449, csa_tree_add_7_25_groupi_n_4450, csa_tree_add_7_25_groupi_n_4451, csa_tree_add_7_25_groupi_n_4452, csa_tree_add_7_25_groupi_n_4453;
  wire csa_tree_add_7_25_groupi_n_4454, csa_tree_add_7_25_groupi_n_4455, csa_tree_add_7_25_groupi_n_4456, csa_tree_add_7_25_groupi_n_4457, csa_tree_add_7_25_groupi_n_4458, csa_tree_add_7_25_groupi_n_4459, csa_tree_add_7_25_groupi_n_4460, csa_tree_add_7_25_groupi_n_4461;
  wire csa_tree_add_7_25_groupi_n_4462, csa_tree_add_7_25_groupi_n_4463, csa_tree_add_7_25_groupi_n_4464, csa_tree_add_7_25_groupi_n_4465, csa_tree_add_7_25_groupi_n_4466, csa_tree_add_7_25_groupi_n_4467, csa_tree_add_7_25_groupi_n_4468, csa_tree_add_7_25_groupi_n_4469;
  wire csa_tree_add_7_25_groupi_n_4470, csa_tree_add_7_25_groupi_n_4471, csa_tree_add_7_25_groupi_n_4472, csa_tree_add_7_25_groupi_n_4473, csa_tree_add_7_25_groupi_n_4474, csa_tree_add_7_25_groupi_n_4475, csa_tree_add_7_25_groupi_n_4476, csa_tree_add_7_25_groupi_n_4477;
  wire csa_tree_add_7_25_groupi_n_4478, csa_tree_add_7_25_groupi_n_4479, csa_tree_add_7_25_groupi_n_4480, csa_tree_add_7_25_groupi_n_4481, csa_tree_add_7_25_groupi_n_4482, csa_tree_add_7_25_groupi_n_4483, csa_tree_add_7_25_groupi_n_4484, csa_tree_add_7_25_groupi_n_4485;
  wire csa_tree_add_7_25_groupi_n_4486, csa_tree_add_7_25_groupi_n_4487, csa_tree_add_7_25_groupi_n_4488, csa_tree_add_7_25_groupi_n_4489, csa_tree_add_7_25_groupi_n_4490, csa_tree_add_7_25_groupi_n_4491, csa_tree_add_7_25_groupi_n_4492, csa_tree_add_7_25_groupi_n_4493;
  wire csa_tree_add_7_25_groupi_n_4494, csa_tree_add_7_25_groupi_n_4495, csa_tree_add_7_25_groupi_n_4496, csa_tree_add_7_25_groupi_n_4497, csa_tree_add_7_25_groupi_n_4498, csa_tree_add_7_25_groupi_n_4499, csa_tree_add_7_25_groupi_n_4500, csa_tree_add_7_25_groupi_n_4501;
  wire csa_tree_add_7_25_groupi_n_4502, csa_tree_add_7_25_groupi_n_4503, csa_tree_add_7_25_groupi_n_4504, csa_tree_add_7_25_groupi_n_4505, csa_tree_add_7_25_groupi_n_4506, csa_tree_add_7_25_groupi_n_4507, csa_tree_add_7_25_groupi_n_4508, csa_tree_add_7_25_groupi_n_4509;
  wire csa_tree_add_7_25_groupi_n_4510, csa_tree_add_7_25_groupi_n_4511, csa_tree_add_7_25_groupi_n_4512, csa_tree_add_7_25_groupi_n_4513, csa_tree_add_7_25_groupi_n_4514, csa_tree_add_7_25_groupi_n_4515, csa_tree_add_7_25_groupi_n_4516, csa_tree_add_7_25_groupi_n_4517;
  wire csa_tree_add_7_25_groupi_n_4518, csa_tree_add_7_25_groupi_n_4519, csa_tree_add_7_25_groupi_n_4520, csa_tree_add_7_25_groupi_n_4521, csa_tree_add_7_25_groupi_n_4522, csa_tree_add_7_25_groupi_n_4523, csa_tree_add_7_25_groupi_n_4524, csa_tree_add_7_25_groupi_n_4525;
  wire csa_tree_add_7_25_groupi_n_4526, csa_tree_add_7_25_groupi_n_4527, csa_tree_add_7_25_groupi_n_4528, csa_tree_add_7_25_groupi_n_4529, csa_tree_add_7_25_groupi_n_4530, csa_tree_add_7_25_groupi_n_4531, csa_tree_add_7_25_groupi_n_4532, csa_tree_add_7_25_groupi_n_4533;
  wire csa_tree_add_7_25_groupi_n_4534, csa_tree_add_7_25_groupi_n_4535, csa_tree_add_7_25_groupi_n_4536, csa_tree_add_7_25_groupi_n_4537, csa_tree_add_7_25_groupi_n_4538, csa_tree_add_7_25_groupi_n_4539, csa_tree_add_7_25_groupi_n_4540, csa_tree_add_7_25_groupi_n_4541;
  wire csa_tree_add_7_25_groupi_n_4542, csa_tree_add_7_25_groupi_n_4543, csa_tree_add_7_25_groupi_n_4544, csa_tree_add_7_25_groupi_n_4545, csa_tree_add_7_25_groupi_n_4546, csa_tree_add_7_25_groupi_n_4547, csa_tree_add_7_25_groupi_n_4548, csa_tree_add_7_25_groupi_n_4549;
  wire csa_tree_add_7_25_groupi_n_4550, csa_tree_add_7_25_groupi_n_4551, csa_tree_add_7_25_groupi_n_4552, csa_tree_add_7_25_groupi_n_4553, csa_tree_add_7_25_groupi_n_4554, csa_tree_add_7_25_groupi_n_4555, csa_tree_add_7_25_groupi_n_4556, csa_tree_add_7_25_groupi_n_4557;
  wire csa_tree_add_7_25_groupi_n_4558, csa_tree_add_7_25_groupi_n_4559, csa_tree_add_7_25_groupi_n_4560, csa_tree_add_7_25_groupi_n_4561, csa_tree_add_7_25_groupi_n_4562, csa_tree_add_7_25_groupi_n_4563, csa_tree_add_7_25_groupi_n_4564, csa_tree_add_7_25_groupi_n_4565;
  wire csa_tree_add_7_25_groupi_n_4566, csa_tree_add_7_25_groupi_n_4567, csa_tree_add_7_25_groupi_n_4568, csa_tree_add_7_25_groupi_n_4569, csa_tree_add_7_25_groupi_n_4570, csa_tree_add_7_25_groupi_n_4571, csa_tree_add_7_25_groupi_n_4572, csa_tree_add_7_25_groupi_n_4573;
  wire csa_tree_add_7_25_groupi_n_4574, csa_tree_add_7_25_groupi_n_4575, csa_tree_add_7_25_groupi_n_4576, csa_tree_add_7_25_groupi_n_4577, csa_tree_add_7_25_groupi_n_4578, csa_tree_add_7_25_groupi_n_4579, csa_tree_add_7_25_groupi_n_4580, csa_tree_add_7_25_groupi_n_4581;
  wire csa_tree_add_7_25_groupi_n_4582, csa_tree_add_7_25_groupi_n_4583, csa_tree_add_7_25_groupi_n_4584, csa_tree_add_7_25_groupi_n_4585, csa_tree_add_7_25_groupi_n_4586, csa_tree_add_7_25_groupi_n_4587, csa_tree_add_7_25_groupi_n_4588, csa_tree_add_7_25_groupi_n_4589;
  wire csa_tree_add_7_25_groupi_n_4590, csa_tree_add_7_25_groupi_n_4591, csa_tree_add_7_25_groupi_n_4592, csa_tree_add_7_25_groupi_n_4593, csa_tree_add_7_25_groupi_n_4594, csa_tree_add_7_25_groupi_n_4595, csa_tree_add_7_25_groupi_n_4596, csa_tree_add_7_25_groupi_n_4597;
  wire csa_tree_add_7_25_groupi_n_4598, csa_tree_add_7_25_groupi_n_4599, csa_tree_add_7_25_groupi_n_4600, csa_tree_add_7_25_groupi_n_4601, csa_tree_add_7_25_groupi_n_4602, csa_tree_add_7_25_groupi_n_4603, csa_tree_add_7_25_groupi_n_4604, csa_tree_add_7_25_groupi_n_4605;
  wire csa_tree_add_7_25_groupi_n_4606, csa_tree_add_7_25_groupi_n_4607, csa_tree_add_7_25_groupi_n_4608, csa_tree_add_7_25_groupi_n_4609, csa_tree_add_7_25_groupi_n_4610, csa_tree_add_7_25_groupi_n_4611, csa_tree_add_7_25_groupi_n_4612, csa_tree_add_7_25_groupi_n_4613;
  wire csa_tree_add_7_25_groupi_n_4614, csa_tree_add_7_25_groupi_n_4615, csa_tree_add_7_25_groupi_n_4616, csa_tree_add_7_25_groupi_n_4617, csa_tree_add_7_25_groupi_n_4618, csa_tree_add_7_25_groupi_n_4619, csa_tree_add_7_25_groupi_n_4620, csa_tree_add_7_25_groupi_n_4621;
  wire csa_tree_add_7_25_groupi_n_4622, csa_tree_add_7_25_groupi_n_4623, csa_tree_add_7_25_groupi_n_4624, csa_tree_add_7_25_groupi_n_4625, csa_tree_add_7_25_groupi_n_4626, csa_tree_add_7_25_groupi_n_4627, csa_tree_add_7_25_groupi_n_4628, csa_tree_add_7_25_groupi_n_4629;
  wire csa_tree_add_7_25_groupi_n_4630, csa_tree_add_7_25_groupi_n_4631, csa_tree_add_7_25_groupi_n_4632, csa_tree_add_7_25_groupi_n_4633, csa_tree_add_7_25_groupi_n_4634, csa_tree_add_7_25_groupi_n_4635, csa_tree_add_7_25_groupi_n_4636, csa_tree_add_7_25_groupi_n_4637;
  wire csa_tree_add_7_25_groupi_n_4638, csa_tree_add_7_25_groupi_n_4639, csa_tree_add_7_25_groupi_n_4640, csa_tree_add_7_25_groupi_n_4641, csa_tree_add_7_25_groupi_n_4642, csa_tree_add_7_25_groupi_n_4643, csa_tree_add_7_25_groupi_n_4644, csa_tree_add_7_25_groupi_n_4645;
  wire csa_tree_add_7_25_groupi_n_4646, csa_tree_add_7_25_groupi_n_4647, csa_tree_add_7_25_groupi_n_4648, csa_tree_add_7_25_groupi_n_4649, csa_tree_add_7_25_groupi_n_4650, csa_tree_add_7_25_groupi_n_4651, csa_tree_add_7_25_groupi_n_4652, csa_tree_add_7_25_groupi_n_4653;
  wire csa_tree_add_7_25_groupi_n_4654, csa_tree_add_7_25_groupi_n_4655, csa_tree_add_7_25_groupi_n_4656, csa_tree_add_7_25_groupi_n_4657, csa_tree_add_7_25_groupi_n_4658, csa_tree_add_7_25_groupi_n_4659, csa_tree_add_7_25_groupi_n_4660, csa_tree_add_7_25_groupi_n_4661;
  wire csa_tree_add_7_25_groupi_n_4662, csa_tree_add_7_25_groupi_n_4663, csa_tree_add_7_25_groupi_n_4664, csa_tree_add_7_25_groupi_n_4665, csa_tree_add_7_25_groupi_n_4666, csa_tree_add_7_25_groupi_n_4667, csa_tree_add_7_25_groupi_n_4668, csa_tree_add_7_25_groupi_n_4669;
  wire csa_tree_add_7_25_groupi_n_4670, csa_tree_add_7_25_groupi_n_4671, csa_tree_add_7_25_groupi_n_4672, csa_tree_add_7_25_groupi_n_4673, csa_tree_add_7_25_groupi_n_4674, csa_tree_add_7_25_groupi_n_4675, csa_tree_add_7_25_groupi_n_4676, csa_tree_add_7_25_groupi_n_4677;
  wire csa_tree_add_7_25_groupi_n_4678, csa_tree_add_7_25_groupi_n_4679, csa_tree_add_7_25_groupi_n_4680, csa_tree_add_7_25_groupi_n_4681, csa_tree_add_7_25_groupi_n_4682, csa_tree_add_7_25_groupi_n_4683, csa_tree_add_7_25_groupi_n_4684, csa_tree_add_7_25_groupi_n_4685;
  wire csa_tree_add_7_25_groupi_n_4686, csa_tree_add_7_25_groupi_n_4687, csa_tree_add_7_25_groupi_n_4688, csa_tree_add_7_25_groupi_n_4689, csa_tree_add_7_25_groupi_n_4690, csa_tree_add_7_25_groupi_n_4691, csa_tree_add_7_25_groupi_n_4692, csa_tree_add_7_25_groupi_n_4693;
  wire csa_tree_add_7_25_groupi_n_4694, csa_tree_add_7_25_groupi_n_4695, csa_tree_add_7_25_groupi_n_4696, csa_tree_add_7_25_groupi_n_4697, csa_tree_add_7_25_groupi_n_4698, csa_tree_add_7_25_groupi_n_4699, csa_tree_add_7_25_groupi_n_4700, csa_tree_add_7_25_groupi_n_4701;
  wire csa_tree_add_7_25_groupi_n_4702, csa_tree_add_7_25_groupi_n_4703, csa_tree_add_7_25_groupi_n_4704, csa_tree_add_7_25_groupi_n_4705, csa_tree_add_7_25_groupi_n_4706, csa_tree_add_7_25_groupi_n_4707, csa_tree_add_7_25_groupi_n_4708, csa_tree_add_7_25_groupi_n_4709;
  wire csa_tree_add_7_25_groupi_n_4710, csa_tree_add_7_25_groupi_n_4711, csa_tree_add_7_25_groupi_n_4712, csa_tree_add_7_25_groupi_n_4713, csa_tree_add_7_25_groupi_n_4714, csa_tree_add_7_25_groupi_n_4715, csa_tree_add_7_25_groupi_n_4716, csa_tree_add_7_25_groupi_n_4717;
  wire csa_tree_add_7_25_groupi_n_4718, csa_tree_add_7_25_groupi_n_4719, csa_tree_add_7_25_groupi_n_4720, csa_tree_add_7_25_groupi_n_4721, csa_tree_add_7_25_groupi_n_4722, csa_tree_add_7_25_groupi_n_4723, csa_tree_add_7_25_groupi_n_4724, csa_tree_add_7_25_groupi_n_4725;
  wire csa_tree_add_7_25_groupi_n_4726, csa_tree_add_7_25_groupi_n_4727, csa_tree_add_7_25_groupi_n_4728, csa_tree_add_7_25_groupi_n_4729, csa_tree_add_7_25_groupi_n_4730, csa_tree_add_7_25_groupi_n_4731, csa_tree_add_7_25_groupi_n_4732, csa_tree_add_7_25_groupi_n_4733;
  wire csa_tree_add_7_25_groupi_n_4734, csa_tree_add_7_25_groupi_n_4735, csa_tree_add_7_25_groupi_n_4736, csa_tree_add_7_25_groupi_n_4737, csa_tree_add_7_25_groupi_n_4738, csa_tree_add_7_25_groupi_n_4739, csa_tree_add_7_25_groupi_n_4740, csa_tree_add_7_25_groupi_n_4741;
  wire csa_tree_add_7_25_groupi_n_4742, csa_tree_add_7_25_groupi_n_4743, csa_tree_add_7_25_groupi_n_4744, csa_tree_add_7_25_groupi_n_4745, csa_tree_add_7_25_groupi_n_4746, csa_tree_add_7_25_groupi_n_4747, csa_tree_add_7_25_groupi_n_4748, csa_tree_add_7_25_groupi_n_4749;
  wire csa_tree_add_7_25_groupi_n_4750, csa_tree_add_7_25_groupi_n_4751, csa_tree_add_7_25_groupi_n_4752, csa_tree_add_7_25_groupi_n_4753, csa_tree_add_7_25_groupi_n_4754, csa_tree_add_7_25_groupi_n_4755, csa_tree_add_7_25_groupi_n_4756, csa_tree_add_7_25_groupi_n_4757;
  wire csa_tree_add_7_25_groupi_n_4758, csa_tree_add_7_25_groupi_n_4759, csa_tree_add_7_25_groupi_n_4760, csa_tree_add_7_25_groupi_n_4761, csa_tree_add_7_25_groupi_n_4762, csa_tree_add_7_25_groupi_n_4763, csa_tree_add_7_25_groupi_n_4764, csa_tree_add_7_25_groupi_n_4765;
  wire csa_tree_add_7_25_groupi_n_4766, csa_tree_add_7_25_groupi_n_4767, csa_tree_add_7_25_groupi_n_4768, csa_tree_add_7_25_groupi_n_4769, csa_tree_add_7_25_groupi_n_4770, csa_tree_add_7_25_groupi_n_4771, csa_tree_add_7_25_groupi_n_4772, csa_tree_add_7_25_groupi_n_4773;
  wire csa_tree_add_7_25_groupi_n_4774, csa_tree_add_7_25_groupi_n_4776, csa_tree_add_7_25_groupi_n_4777, csa_tree_add_7_25_groupi_n_4778, csa_tree_add_7_25_groupi_n_4779, csa_tree_add_7_25_groupi_n_4780, csa_tree_add_7_25_groupi_n_4781, csa_tree_add_7_25_groupi_n_4782;
  wire csa_tree_add_7_25_groupi_n_4783, csa_tree_add_7_25_groupi_n_4784, csa_tree_add_7_25_groupi_n_4785, csa_tree_add_7_25_groupi_n_4786, csa_tree_add_7_25_groupi_n_4787, csa_tree_add_7_25_groupi_n_4788, csa_tree_add_7_25_groupi_n_4789, csa_tree_add_7_25_groupi_n_4790;
  wire csa_tree_add_7_25_groupi_n_4791, csa_tree_add_7_25_groupi_n_4792, csa_tree_add_7_25_groupi_n_4793, csa_tree_add_7_25_groupi_n_4794, csa_tree_add_7_25_groupi_n_4795, csa_tree_add_7_25_groupi_n_4796, csa_tree_add_7_25_groupi_n_4797, csa_tree_add_7_25_groupi_n_4798;
  wire csa_tree_add_7_25_groupi_n_4799, csa_tree_add_7_25_groupi_n_4800, csa_tree_add_7_25_groupi_n_4801, csa_tree_add_7_25_groupi_n_4802, csa_tree_add_7_25_groupi_n_4803, csa_tree_add_7_25_groupi_n_4804, csa_tree_add_7_25_groupi_n_4805, csa_tree_add_7_25_groupi_n_4806;
  wire csa_tree_add_7_25_groupi_n_4807, csa_tree_add_7_25_groupi_n_4808, csa_tree_add_7_25_groupi_n_4809, csa_tree_add_7_25_groupi_n_4810, csa_tree_add_7_25_groupi_n_4811, csa_tree_add_7_25_groupi_n_4812, csa_tree_add_7_25_groupi_n_4813, csa_tree_add_7_25_groupi_n_4814;
  wire csa_tree_add_7_25_groupi_n_4815, csa_tree_add_7_25_groupi_n_4816, csa_tree_add_7_25_groupi_n_4817, csa_tree_add_7_25_groupi_n_4818, csa_tree_add_7_25_groupi_n_4819, csa_tree_add_7_25_groupi_n_4820, csa_tree_add_7_25_groupi_n_4821, csa_tree_add_7_25_groupi_n_4822;
  wire csa_tree_add_7_25_groupi_n_4823, csa_tree_add_7_25_groupi_n_4824, csa_tree_add_7_25_groupi_n_4825, csa_tree_add_7_25_groupi_n_4826, csa_tree_add_7_25_groupi_n_4827, csa_tree_add_7_25_groupi_n_4828, csa_tree_add_7_25_groupi_n_4829, csa_tree_add_7_25_groupi_n_4830;
  wire csa_tree_add_7_25_groupi_n_4831, csa_tree_add_7_25_groupi_n_4832, csa_tree_add_7_25_groupi_n_4833, csa_tree_add_7_25_groupi_n_4834, csa_tree_add_7_25_groupi_n_4835, csa_tree_add_7_25_groupi_n_4836, csa_tree_add_7_25_groupi_n_4837, csa_tree_add_7_25_groupi_n_4838;
  wire csa_tree_add_7_25_groupi_n_4839, csa_tree_add_7_25_groupi_n_4840, csa_tree_add_7_25_groupi_n_4841, csa_tree_add_7_25_groupi_n_4842, csa_tree_add_7_25_groupi_n_4843, csa_tree_add_7_25_groupi_n_4844, csa_tree_add_7_25_groupi_n_4845, csa_tree_add_7_25_groupi_n_4846;
  wire csa_tree_add_7_25_groupi_n_4847, csa_tree_add_7_25_groupi_n_4848, csa_tree_add_7_25_groupi_n_4849, csa_tree_add_7_25_groupi_n_4850, csa_tree_add_7_25_groupi_n_4851, csa_tree_add_7_25_groupi_n_4852, csa_tree_add_7_25_groupi_n_4853, csa_tree_add_7_25_groupi_n_4854;
  wire csa_tree_add_7_25_groupi_n_4855, csa_tree_add_7_25_groupi_n_4856, csa_tree_add_7_25_groupi_n_4857, csa_tree_add_7_25_groupi_n_4858, csa_tree_add_7_25_groupi_n_4859, csa_tree_add_7_25_groupi_n_4860, csa_tree_add_7_25_groupi_n_4861, csa_tree_add_7_25_groupi_n_4862;
  wire csa_tree_add_7_25_groupi_n_4863, csa_tree_add_7_25_groupi_n_4864, csa_tree_add_7_25_groupi_n_4865, csa_tree_add_7_25_groupi_n_4866, csa_tree_add_7_25_groupi_n_4867, csa_tree_add_7_25_groupi_n_4868, csa_tree_add_7_25_groupi_n_4869, csa_tree_add_7_25_groupi_n_4870;
  wire csa_tree_add_7_25_groupi_n_4871, csa_tree_add_7_25_groupi_n_4872, csa_tree_add_7_25_groupi_n_4873, csa_tree_add_7_25_groupi_n_4874, csa_tree_add_7_25_groupi_n_4875, csa_tree_add_7_25_groupi_n_4876, csa_tree_add_7_25_groupi_n_4877, csa_tree_add_7_25_groupi_n_4878;
  wire csa_tree_add_7_25_groupi_n_4879, csa_tree_add_7_25_groupi_n_4880, csa_tree_add_7_25_groupi_n_4881, csa_tree_add_7_25_groupi_n_4882, csa_tree_add_7_25_groupi_n_4883, csa_tree_add_7_25_groupi_n_4884, csa_tree_add_7_25_groupi_n_4886, csa_tree_add_7_25_groupi_n_4887;
  wire csa_tree_add_7_25_groupi_n_4888, csa_tree_add_7_25_groupi_n_4889, csa_tree_add_7_25_groupi_n_4890, csa_tree_add_7_25_groupi_n_4891, csa_tree_add_7_25_groupi_n_4892, csa_tree_add_7_25_groupi_n_4893, csa_tree_add_7_25_groupi_n_4894, csa_tree_add_7_25_groupi_n_4895;
  wire csa_tree_add_7_25_groupi_n_4896, csa_tree_add_7_25_groupi_n_4897, csa_tree_add_7_25_groupi_n_4898, csa_tree_add_7_25_groupi_n_4899, csa_tree_add_7_25_groupi_n_4900, csa_tree_add_7_25_groupi_n_4901, csa_tree_add_7_25_groupi_n_4902, csa_tree_add_7_25_groupi_n_4903;
  wire csa_tree_add_7_25_groupi_n_4904, csa_tree_add_7_25_groupi_n_4905, csa_tree_add_7_25_groupi_n_4906, csa_tree_add_7_25_groupi_n_4907, csa_tree_add_7_25_groupi_n_4908, csa_tree_add_7_25_groupi_n_4909, csa_tree_add_7_25_groupi_n_4910, csa_tree_add_7_25_groupi_n_4911;
  wire csa_tree_add_7_25_groupi_n_4912, csa_tree_add_7_25_groupi_n_4913, csa_tree_add_7_25_groupi_n_4914, csa_tree_add_7_25_groupi_n_4915, csa_tree_add_7_25_groupi_n_4916, csa_tree_add_7_25_groupi_n_4917, csa_tree_add_7_25_groupi_n_4918, csa_tree_add_7_25_groupi_n_4919;
  wire csa_tree_add_7_25_groupi_n_4920, csa_tree_add_7_25_groupi_n_4921, csa_tree_add_7_25_groupi_n_4922, csa_tree_add_7_25_groupi_n_4923, csa_tree_add_7_25_groupi_n_4924, csa_tree_add_7_25_groupi_n_4925, csa_tree_add_7_25_groupi_n_4926, csa_tree_add_7_25_groupi_n_4927;
  wire csa_tree_add_7_25_groupi_n_4928, csa_tree_add_7_25_groupi_n_4929, csa_tree_add_7_25_groupi_n_4930, csa_tree_add_7_25_groupi_n_4931, csa_tree_add_7_25_groupi_n_4932, csa_tree_add_7_25_groupi_n_4933, csa_tree_add_7_25_groupi_n_4934, csa_tree_add_7_25_groupi_n_4935;
  wire csa_tree_add_7_25_groupi_n_4936, csa_tree_add_7_25_groupi_n_4937, csa_tree_add_7_25_groupi_n_4938, csa_tree_add_7_25_groupi_n_4939, csa_tree_add_7_25_groupi_n_4940, csa_tree_add_7_25_groupi_n_4941, csa_tree_add_7_25_groupi_n_4942, csa_tree_add_7_25_groupi_n_4943;
  wire csa_tree_add_7_25_groupi_n_4944, csa_tree_add_7_25_groupi_n_4945, csa_tree_add_7_25_groupi_n_4946, csa_tree_add_7_25_groupi_n_4947, csa_tree_add_7_25_groupi_n_4948, csa_tree_add_7_25_groupi_n_4949, csa_tree_add_7_25_groupi_n_4950, csa_tree_add_7_25_groupi_n_4951;
  wire csa_tree_add_7_25_groupi_n_4952, csa_tree_add_7_25_groupi_n_4953, csa_tree_add_7_25_groupi_n_4954, csa_tree_add_7_25_groupi_n_4955, csa_tree_add_7_25_groupi_n_4956, csa_tree_add_7_25_groupi_n_4957, csa_tree_add_7_25_groupi_n_4958, csa_tree_add_7_25_groupi_n_4959;
  wire csa_tree_add_7_25_groupi_n_4960, csa_tree_add_7_25_groupi_n_4961, csa_tree_add_7_25_groupi_n_4962, csa_tree_add_7_25_groupi_n_4963, csa_tree_add_7_25_groupi_n_4964, csa_tree_add_7_25_groupi_n_4965, csa_tree_add_7_25_groupi_n_4966, csa_tree_add_7_25_groupi_n_4967;
  wire csa_tree_add_7_25_groupi_n_4968, csa_tree_add_7_25_groupi_n_4969, csa_tree_add_7_25_groupi_n_4970, csa_tree_add_7_25_groupi_n_4971, csa_tree_add_7_25_groupi_n_4972, csa_tree_add_7_25_groupi_n_4973, csa_tree_add_7_25_groupi_n_4974, csa_tree_add_7_25_groupi_n_4975;
  wire csa_tree_add_7_25_groupi_n_4976, csa_tree_add_7_25_groupi_n_4977, csa_tree_add_7_25_groupi_n_4978, csa_tree_add_7_25_groupi_n_4979, csa_tree_add_7_25_groupi_n_4980, csa_tree_add_7_25_groupi_n_4981, csa_tree_add_7_25_groupi_n_4982, csa_tree_add_7_25_groupi_n_4983;
  wire csa_tree_add_7_25_groupi_n_4984, csa_tree_add_7_25_groupi_n_4985, csa_tree_add_7_25_groupi_n_4986, csa_tree_add_7_25_groupi_n_4987, csa_tree_add_7_25_groupi_n_4988, csa_tree_add_7_25_groupi_n_4989, csa_tree_add_7_25_groupi_n_4990, csa_tree_add_7_25_groupi_n_4991;
  wire csa_tree_add_7_25_groupi_n_4993, csa_tree_add_7_25_groupi_n_4994, csa_tree_add_7_25_groupi_n_4995, csa_tree_add_7_25_groupi_n_4996, csa_tree_add_7_25_groupi_n_4997, csa_tree_add_7_25_groupi_n_4998, csa_tree_add_7_25_groupi_n_4999, csa_tree_add_7_25_groupi_n_5000;
  wire csa_tree_add_7_25_groupi_n_5001, csa_tree_add_7_25_groupi_n_5002, csa_tree_add_7_25_groupi_n_5003, csa_tree_add_7_25_groupi_n_5004, csa_tree_add_7_25_groupi_n_5005, csa_tree_add_7_25_groupi_n_5006, csa_tree_add_7_25_groupi_n_5007, csa_tree_add_7_25_groupi_n_5008;
  wire csa_tree_add_7_25_groupi_n_5009, csa_tree_add_7_25_groupi_n_5010, csa_tree_add_7_25_groupi_n_5011, csa_tree_add_7_25_groupi_n_5012, csa_tree_add_7_25_groupi_n_5013, csa_tree_add_7_25_groupi_n_5014, csa_tree_add_7_25_groupi_n_5015, csa_tree_add_7_25_groupi_n_5016;
  wire csa_tree_add_7_25_groupi_n_5017, csa_tree_add_7_25_groupi_n_5018, csa_tree_add_7_25_groupi_n_5019, csa_tree_add_7_25_groupi_n_5020, csa_tree_add_7_25_groupi_n_5021, csa_tree_add_7_25_groupi_n_5022, csa_tree_add_7_25_groupi_n_5023, csa_tree_add_7_25_groupi_n_5024;
  wire csa_tree_add_7_25_groupi_n_5025, csa_tree_add_7_25_groupi_n_5026, csa_tree_add_7_25_groupi_n_5027, csa_tree_add_7_25_groupi_n_5028, csa_tree_add_7_25_groupi_n_5029, csa_tree_add_7_25_groupi_n_5030, csa_tree_add_7_25_groupi_n_5031, csa_tree_add_7_25_groupi_n_5032;
  wire csa_tree_add_7_25_groupi_n_5033, csa_tree_add_7_25_groupi_n_5034, csa_tree_add_7_25_groupi_n_5035, csa_tree_add_7_25_groupi_n_5036, csa_tree_add_7_25_groupi_n_5037, csa_tree_add_7_25_groupi_n_5038, csa_tree_add_7_25_groupi_n_5039, csa_tree_add_7_25_groupi_n_5040;
  wire csa_tree_add_7_25_groupi_n_5041, csa_tree_add_7_25_groupi_n_5042, csa_tree_add_7_25_groupi_n_5043, csa_tree_add_7_25_groupi_n_5044, csa_tree_add_7_25_groupi_n_5045, csa_tree_add_7_25_groupi_n_5046, csa_tree_add_7_25_groupi_n_5047, csa_tree_add_7_25_groupi_n_5048;
  wire csa_tree_add_7_25_groupi_n_5049, csa_tree_add_7_25_groupi_n_5050, csa_tree_add_7_25_groupi_n_5051, csa_tree_add_7_25_groupi_n_5052, csa_tree_add_7_25_groupi_n_5053, csa_tree_add_7_25_groupi_n_5054, csa_tree_add_7_25_groupi_n_5055, csa_tree_add_7_25_groupi_n_5056;
  wire csa_tree_add_7_25_groupi_n_5057, csa_tree_add_7_25_groupi_n_5058, csa_tree_add_7_25_groupi_n_5059, csa_tree_add_7_25_groupi_n_5060, csa_tree_add_7_25_groupi_n_5061, csa_tree_add_7_25_groupi_n_5062, csa_tree_add_7_25_groupi_n_5063, csa_tree_add_7_25_groupi_n_5064;
  wire csa_tree_add_7_25_groupi_n_5065, csa_tree_add_7_25_groupi_n_5066, csa_tree_add_7_25_groupi_n_5067, csa_tree_add_7_25_groupi_n_5068, csa_tree_add_7_25_groupi_n_5069, csa_tree_add_7_25_groupi_n_5070, csa_tree_add_7_25_groupi_n_5071, csa_tree_add_7_25_groupi_n_5072;
  wire csa_tree_add_7_25_groupi_n_5073, csa_tree_add_7_25_groupi_n_5074, csa_tree_add_7_25_groupi_n_5075, csa_tree_add_7_25_groupi_n_5076, csa_tree_add_7_25_groupi_n_5077, csa_tree_add_7_25_groupi_n_5078, csa_tree_add_7_25_groupi_n_5080, csa_tree_add_7_25_groupi_n_5081;
  wire csa_tree_add_7_25_groupi_n_5082, csa_tree_add_7_25_groupi_n_5083, csa_tree_add_7_25_groupi_n_5084, csa_tree_add_7_25_groupi_n_5085, csa_tree_add_7_25_groupi_n_5086, csa_tree_add_7_25_groupi_n_5087, csa_tree_add_7_25_groupi_n_5088, csa_tree_add_7_25_groupi_n_5089;
  wire csa_tree_add_7_25_groupi_n_5090, csa_tree_add_7_25_groupi_n_5091, csa_tree_add_7_25_groupi_n_5092, csa_tree_add_7_25_groupi_n_5093, csa_tree_add_7_25_groupi_n_5094, csa_tree_add_7_25_groupi_n_5095, csa_tree_add_7_25_groupi_n_5096, csa_tree_add_7_25_groupi_n_5097;
  wire csa_tree_add_7_25_groupi_n_5098, csa_tree_add_7_25_groupi_n_5099, csa_tree_add_7_25_groupi_n_5100, csa_tree_add_7_25_groupi_n_5101, csa_tree_add_7_25_groupi_n_5102, csa_tree_add_7_25_groupi_n_5103, csa_tree_add_7_25_groupi_n_5104, csa_tree_add_7_25_groupi_n_5105;
  wire csa_tree_add_7_25_groupi_n_5106, csa_tree_add_7_25_groupi_n_5107, csa_tree_add_7_25_groupi_n_5108, csa_tree_add_7_25_groupi_n_5109, csa_tree_add_7_25_groupi_n_5110, csa_tree_add_7_25_groupi_n_5111, csa_tree_add_7_25_groupi_n_5112, csa_tree_add_7_25_groupi_n_5113;
  wire csa_tree_add_7_25_groupi_n_5114, csa_tree_add_7_25_groupi_n_5115, csa_tree_add_7_25_groupi_n_5116, csa_tree_add_7_25_groupi_n_5117, csa_tree_add_7_25_groupi_n_5118, csa_tree_add_7_25_groupi_n_5119, csa_tree_add_7_25_groupi_n_5120, csa_tree_add_7_25_groupi_n_5121;
  wire csa_tree_add_7_25_groupi_n_5122, csa_tree_add_7_25_groupi_n_5123, csa_tree_add_7_25_groupi_n_5124, csa_tree_add_7_25_groupi_n_5125, csa_tree_add_7_25_groupi_n_5126, csa_tree_add_7_25_groupi_n_5127, csa_tree_add_7_25_groupi_n_5128, csa_tree_add_7_25_groupi_n_5129;
  wire csa_tree_add_7_25_groupi_n_5130, csa_tree_add_7_25_groupi_n_5131, csa_tree_add_7_25_groupi_n_5132, csa_tree_add_7_25_groupi_n_5133, csa_tree_add_7_25_groupi_n_5134, csa_tree_add_7_25_groupi_n_5135, csa_tree_add_7_25_groupi_n_5136, csa_tree_add_7_25_groupi_n_5137;
  wire csa_tree_add_7_25_groupi_n_5138, csa_tree_add_7_25_groupi_n_5139, csa_tree_add_7_25_groupi_n_5140, csa_tree_add_7_25_groupi_n_5141, csa_tree_add_7_25_groupi_n_5142, csa_tree_add_7_25_groupi_n_5143, csa_tree_add_7_25_groupi_n_5144, csa_tree_add_7_25_groupi_n_5145;
  wire csa_tree_add_7_25_groupi_n_5146, csa_tree_add_7_25_groupi_n_5147, csa_tree_add_7_25_groupi_n_5148, csa_tree_add_7_25_groupi_n_5149, csa_tree_add_7_25_groupi_n_5150, csa_tree_add_7_25_groupi_n_5151, csa_tree_add_7_25_groupi_n_5152, csa_tree_add_7_25_groupi_n_5153;
  wire csa_tree_add_7_25_groupi_n_5154, csa_tree_add_7_25_groupi_n_5155, csa_tree_add_7_25_groupi_n_5156, csa_tree_add_7_25_groupi_n_5157, csa_tree_add_7_25_groupi_n_5158, csa_tree_add_7_25_groupi_n_5159, csa_tree_add_7_25_groupi_n_5160, csa_tree_add_7_25_groupi_n_5161;
  wire csa_tree_add_7_25_groupi_n_5162, csa_tree_add_7_25_groupi_n_5163, csa_tree_add_7_25_groupi_n_5164, csa_tree_add_7_25_groupi_n_5165, csa_tree_add_7_25_groupi_n_5166, csa_tree_add_7_25_groupi_n_5168, csa_tree_add_7_25_groupi_n_5169, csa_tree_add_7_25_groupi_n_5170;
  wire csa_tree_add_7_25_groupi_n_5171, csa_tree_add_7_25_groupi_n_5172, csa_tree_add_7_25_groupi_n_5173, csa_tree_add_7_25_groupi_n_5174, csa_tree_add_7_25_groupi_n_5175, csa_tree_add_7_25_groupi_n_5176, csa_tree_add_7_25_groupi_n_5177, csa_tree_add_7_25_groupi_n_5178;
  wire csa_tree_add_7_25_groupi_n_5179, csa_tree_add_7_25_groupi_n_5180, csa_tree_add_7_25_groupi_n_5181, csa_tree_add_7_25_groupi_n_5182, csa_tree_add_7_25_groupi_n_5183, csa_tree_add_7_25_groupi_n_5184, csa_tree_add_7_25_groupi_n_5185, csa_tree_add_7_25_groupi_n_5186;
  wire csa_tree_add_7_25_groupi_n_5187, csa_tree_add_7_25_groupi_n_5188, csa_tree_add_7_25_groupi_n_5189, csa_tree_add_7_25_groupi_n_5190, csa_tree_add_7_25_groupi_n_5191, csa_tree_add_7_25_groupi_n_5192, csa_tree_add_7_25_groupi_n_5193, csa_tree_add_7_25_groupi_n_5194;
  wire csa_tree_add_7_25_groupi_n_5195, csa_tree_add_7_25_groupi_n_5196, csa_tree_add_7_25_groupi_n_5197, csa_tree_add_7_25_groupi_n_5198, csa_tree_add_7_25_groupi_n_5199, csa_tree_add_7_25_groupi_n_5200, csa_tree_add_7_25_groupi_n_5201, csa_tree_add_7_25_groupi_n_5202;
  wire csa_tree_add_7_25_groupi_n_5203, csa_tree_add_7_25_groupi_n_5204, csa_tree_add_7_25_groupi_n_5205, csa_tree_add_7_25_groupi_n_5206, csa_tree_add_7_25_groupi_n_5207, csa_tree_add_7_25_groupi_n_5208, csa_tree_add_7_25_groupi_n_5209, csa_tree_add_7_25_groupi_n_5210;
  wire csa_tree_add_7_25_groupi_n_5211, csa_tree_add_7_25_groupi_n_5212, csa_tree_add_7_25_groupi_n_5213, csa_tree_add_7_25_groupi_n_5214, csa_tree_add_7_25_groupi_n_5215, csa_tree_add_7_25_groupi_n_5216, csa_tree_add_7_25_groupi_n_5217, csa_tree_add_7_25_groupi_n_5218;
  wire csa_tree_add_7_25_groupi_n_5219, csa_tree_add_7_25_groupi_n_5220, csa_tree_add_7_25_groupi_n_5221, csa_tree_add_7_25_groupi_n_5222, csa_tree_add_7_25_groupi_n_5223, csa_tree_add_7_25_groupi_n_5224, csa_tree_add_7_25_groupi_n_5225, csa_tree_add_7_25_groupi_n_5226;
  wire csa_tree_add_7_25_groupi_n_5227, csa_tree_add_7_25_groupi_n_5228, csa_tree_add_7_25_groupi_n_5229, csa_tree_add_7_25_groupi_n_5230, csa_tree_add_7_25_groupi_n_5231, csa_tree_add_7_25_groupi_n_5232, csa_tree_add_7_25_groupi_n_5233, csa_tree_add_7_25_groupi_n_5234;
  wire csa_tree_add_7_25_groupi_n_5235, csa_tree_add_7_25_groupi_n_5236, csa_tree_add_7_25_groupi_n_5237, csa_tree_add_7_25_groupi_n_5238, csa_tree_add_7_25_groupi_n_5239, csa_tree_add_7_25_groupi_n_5240, csa_tree_add_7_25_groupi_n_5241, csa_tree_add_7_25_groupi_n_5242;
  wire csa_tree_add_7_25_groupi_n_5243, csa_tree_add_7_25_groupi_n_5244, csa_tree_add_7_25_groupi_n_5245, csa_tree_add_7_25_groupi_n_5246, csa_tree_add_7_25_groupi_n_5247, csa_tree_add_7_25_groupi_n_5248, csa_tree_add_7_25_groupi_n_5249, csa_tree_add_7_25_groupi_n_5250;
  wire csa_tree_add_7_25_groupi_n_5251, csa_tree_add_7_25_groupi_n_5252, csa_tree_add_7_25_groupi_n_5253, csa_tree_add_7_25_groupi_n_5254, csa_tree_add_7_25_groupi_n_5255, csa_tree_add_7_25_groupi_n_5256, csa_tree_add_7_25_groupi_n_5257, csa_tree_add_7_25_groupi_n_5258;
  wire csa_tree_add_7_25_groupi_n_5259, csa_tree_add_7_25_groupi_n_5260, csa_tree_add_7_25_groupi_n_5261, csa_tree_add_7_25_groupi_n_5262, csa_tree_add_7_25_groupi_n_5263, csa_tree_add_7_25_groupi_n_5264, csa_tree_add_7_25_groupi_n_5265, csa_tree_add_7_25_groupi_n_5266;
  wire csa_tree_add_7_25_groupi_n_5267, csa_tree_add_7_25_groupi_n_5268, csa_tree_add_7_25_groupi_n_5269, csa_tree_add_7_25_groupi_n_5270, csa_tree_add_7_25_groupi_n_5271, csa_tree_add_7_25_groupi_n_5272, csa_tree_add_7_25_groupi_n_5273, csa_tree_add_7_25_groupi_n_5274;
  wire csa_tree_add_7_25_groupi_n_5275, csa_tree_add_7_25_groupi_n_5276, csa_tree_add_7_25_groupi_n_5277, csa_tree_add_7_25_groupi_n_5278, csa_tree_add_7_25_groupi_n_5279, csa_tree_add_7_25_groupi_n_5280, csa_tree_add_7_25_groupi_n_5281, csa_tree_add_7_25_groupi_n_5282;
  wire csa_tree_add_7_25_groupi_n_5283, csa_tree_add_7_25_groupi_n_5284, csa_tree_add_7_25_groupi_n_5285, csa_tree_add_7_25_groupi_n_5286, csa_tree_add_7_25_groupi_n_5287, csa_tree_add_7_25_groupi_n_5288, csa_tree_add_7_25_groupi_n_5289, csa_tree_add_7_25_groupi_n_5290;
  wire csa_tree_add_7_25_groupi_n_5291, csa_tree_add_7_25_groupi_n_5292, csa_tree_add_7_25_groupi_n_5293, csa_tree_add_7_25_groupi_n_5294, csa_tree_add_7_25_groupi_n_5295, csa_tree_add_7_25_groupi_n_5296, csa_tree_add_7_25_groupi_n_5297, csa_tree_add_7_25_groupi_n_5298;
  wire csa_tree_add_7_25_groupi_n_5299, csa_tree_add_7_25_groupi_n_5300, csa_tree_add_7_25_groupi_n_5301, csa_tree_add_7_25_groupi_n_5302, csa_tree_add_7_25_groupi_n_5303, csa_tree_add_7_25_groupi_n_5304, csa_tree_add_7_25_groupi_n_5305, csa_tree_add_7_25_groupi_n_5306;
  wire csa_tree_add_7_25_groupi_n_5307, csa_tree_add_7_25_groupi_n_5308, csa_tree_add_7_25_groupi_n_5309, csa_tree_add_7_25_groupi_n_5310, csa_tree_add_7_25_groupi_n_5311, csa_tree_add_7_25_groupi_n_5312, csa_tree_add_7_25_groupi_n_5313, csa_tree_add_7_25_groupi_n_5314;
  wire csa_tree_add_7_25_groupi_n_5315, csa_tree_add_7_25_groupi_n_5316, csa_tree_add_7_25_groupi_n_5317, csa_tree_add_7_25_groupi_n_5318, csa_tree_add_7_25_groupi_n_5319, csa_tree_add_7_25_groupi_n_5320, csa_tree_add_7_25_groupi_n_5321, csa_tree_add_7_25_groupi_n_5322;
  wire csa_tree_add_7_25_groupi_n_5323, csa_tree_add_7_25_groupi_n_5324, csa_tree_add_7_25_groupi_n_5325, csa_tree_add_7_25_groupi_n_5326, csa_tree_add_7_25_groupi_n_5327, csa_tree_add_7_25_groupi_n_5328, csa_tree_add_7_25_groupi_n_5329, csa_tree_add_7_25_groupi_n_5330;
  wire csa_tree_add_7_25_groupi_n_5331, csa_tree_add_7_25_groupi_n_5332, csa_tree_add_7_25_groupi_n_5333, csa_tree_add_7_25_groupi_n_5334, csa_tree_add_7_25_groupi_n_5335, csa_tree_add_7_25_groupi_n_5336, csa_tree_add_7_25_groupi_n_5337, csa_tree_add_7_25_groupi_n_5339;
  wire csa_tree_add_7_25_groupi_n_5340, csa_tree_add_7_25_groupi_n_5341, csa_tree_add_7_25_groupi_n_5342, csa_tree_add_7_25_groupi_n_5343, csa_tree_add_7_25_groupi_n_5344, csa_tree_add_7_25_groupi_n_5345, csa_tree_add_7_25_groupi_n_5346, csa_tree_add_7_25_groupi_n_5347;
  wire csa_tree_add_7_25_groupi_n_5348, csa_tree_add_7_25_groupi_n_5349, csa_tree_add_7_25_groupi_n_5350, csa_tree_add_7_25_groupi_n_5351, csa_tree_add_7_25_groupi_n_5352, csa_tree_add_7_25_groupi_n_5353, csa_tree_add_7_25_groupi_n_5354, csa_tree_add_7_25_groupi_n_5355;
  wire csa_tree_add_7_25_groupi_n_5356, csa_tree_add_7_25_groupi_n_5357, csa_tree_add_7_25_groupi_n_5358, csa_tree_add_7_25_groupi_n_5359, csa_tree_add_7_25_groupi_n_5360, csa_tree_add_7_25_groupi_n_5361, csa_tree_add_7_25_groupi_n_5362, csa_tree_add_7_25_groupi_n_5363;
  wire csa_tree_add_7_25_groupi_n_5364, csa_tree_add_7_25_groupi_n_5365, csa_tree_add_7_25_groupi_n_5366, csa_tree_add_7_25_groupi_n_5367, csa_tree_add_7_25_groupi_n_5368, csa_tree_add_7_25_groupi_n_5369, csa_tree_add_7_25_groupi_n_5370, csa_tree_add_7_25_groupi_n_5371;
  wire csa_tree_add_7_25_groupi_n_5372, csa_tree_add_7_25_groupi_n_5373, csa_tree_add_7_25_groupi_n_5374, csa_tree_add_7_25_groupi_n_5375, csa_tree_add_7_25_groupi_n_5376, csa_tree_add_7_25_groupi_n_5377, csa_tree_add_7_25_groupi_n_5378, csa_tree_add_7_25_groupi_n_5379;
  wire csa_tree_add_7_25_groupi_n_5380, csa_tree_add_7_25_groupi_n_5381, csa_tree_add_7_25_groupi_n_5382, csa_tree_add_7_25_groupi_n_5383, csa_tree_add_7_25_groupi_n_5384, csa_tree_add_7_25_groupi_n_5385, csa_tree_add_7_25_groupi_n_5386, csa_tree_add_7_25_groupi_n_5387;
  wire csa_tree_add_7_25_groupi_n_5388, csa_tree_add_7_25_groupi_n_5389, csa_tree_add_7_25_groupi_n_5390, csa_tree_add_7_25_groupi_n_5391, csa_tree_add_7_25_groupi_n_5392, csa_tree_add_7_25_groupi_n_5393, csa_tree_add_7_25_groupi_n_5394, csa_tree_add_7_25_groupi_n_5395;
  wire csa_tree_add_7_25_groupi_n_5396, csa_tree_add_7_25_groupi_n_5397, csa_tree_add_7_25_groupi_n_5398, csa_tree_add_7_25_groupi_n_5399, csa_tree_add_7_25_groupi_n_5400, csa_tree_add_7_25_groupi_n_5401, csa_tree_add_7_25_groupi_n_5402, csa_tree_add_7_25_groupi_n_5403;
  wire csa_tree_add_7_25_groupi_n_5404, csa_tree_add_7_25_groupi_n_5405, csa_tree_add_7_25_groupi_n_5406, csa_tree_add_7_25_groupi_n_5407, csa_tree_add_7_25_groupi_n_5408, csa_tree_add_7_25_groupi_n_5409, csa_tree_add_7_25_groupi_n_5410, csa_tree_add_7_25_groupi_n_5411;
  wire csa_tree_add_7_25_groupi_n_5412, csa_tree_add_7_25_groupi_n_5413, csa_tree_add_7_25_groupi_n_5414, csa_tree_add_7_25_groupi_n_5415, csa_tree_add_7_25_groupi_n_5416, csa_tree_add_7_25_groupi_n_5417, csa_tree_add_7_25_groupi_n_5418, csa_tree_add_7_25_groupi_n_5419;
  wire csa_tree_add_7_25_groupi_n_5420, csa_tree_add_7_25_groupi_n_5421, csa_tree_add_7_25_groupi_n_5422, csa_tree_add_7_25_groupi_n_5423, csa_tree_add_7_25_groupi_n_5424, csa_tree_add_7_25_groupi_n_5425, csa_tree_add_7_25_groupi_n_5426, csa_tree_add_7_25_groupi_n_5427;
  wire csa_tree_add_7_25_groupi_n_5428, csa_tree_add_7_25_groupi_n_5429, csa_tree_add_7_25_groupi_n_5430, csa_tree_add_7_25_groupi_n_5431, csa_tree_add_7_25_groupi_n_5432, csa_tree_add_7_25_groupi_n_5433, csa_tree_add_7_25_groupi_n_5434, csa_tree_add_7_25_groupi_n_5435;
  wire csa_tree_add_7_25_groupi_n_5436, csa_tree_add_7_25_groupi_n_5437, csa_tree_add_7_25_groupi_n_5438, csa_tree_add_7_25_groupi_n_5439, csa_tree_add_7_25_groupi_n_5440, csa_tree_add_7_25_groupi_n_5441, csa_tree_add_7_25_groupi_n_5442, csa_tree_add_7_25_groupi_n_5443;
  wire csa_tree_add_7_25_groupi_n_5444, csa_tree_add_7_25_groupi_n_5445, csa_tree_add_7_25_groupi_n_5446, csa_tree_add_7_25_groupi_n_5447, csa_tree_add_7_25_groupi_n_5448, csa_tree_add_7_25_groupi_n_5449, csa_tree_add_7_25_groupi_n_5450, csa_tree_add_7_25_groupi_n_5451;
  wire csa_tree_add_7_25_groupi_n_5452, csa_tree_add_7_25_groupi_n_5453, csa_tree_add_7_25_groupi_n_5454, csa_tree_add_7_25_groupi_n_5455, csa_tree_add_7_25_groupi_n_5456, csa_tree_add_7_25_groupi_n_5457, csa_tree_add_7_25_groupi_n_5458, csa_tree_add_7_25_groupi_n_5459;
  wire csa_tree_add_7_25_groupi_n_5460, csa_tree_add_7_25_groupi_n_5461, csa_tree_add_7_25_groupi_n_5463, csa_tree_add_7_25_groupi_n_5464, csa_tree_add_7_25_groupi_n_5465, csa_tree_add_7_25_groupi_n_5466, csa_tree_add_7_25_groupi_n_5467, csa_tree_add_7_25_groupi_n_5468;
  wire csa_tree_add_7_25_groupi_n_5469, csa_tree_add_7_25_groupi_n_5470, csa_tree_add_7_25_groupi_n_5471, csa_tree_add_7_25_groupi_n_5472, csa_tree_add_7_25_groupi_n_5473, csa_tree_add_7_25_groupi_n_5474, csa_tree_add_7_25_groupi_n_5475, csa_tree_add_7_25_groupi_n_5476;
  wire csa_tree_add_7_25_groupi_n_5477, csa_tree_add_7_25_groupi_n_5478, csa_tree_add_7_25_groupi_n_5479, csa_tree_add_7_25_groupi_n_5480, csa_tree_add_7_25_groupi_n_5481, csa_tree_add_7_25_groupi_n_5482, csa_tree_add_7_25_groupi_n_5483, csa_tree_add_7_25_groupi_n_5484;
  wire csa_tree_add_7_25_groupi_n_5485, csa_tree_add_7_25_groupi_n_5486, csa_tree_add_7_25_groupi_n_5487, csa_tree_add_7_25_groupi_n_5488, csa_tree_add_7_25_groupi_n_5489, csa_tree_add_7_25_groupi_n_5490, csa_tree_add_7_25_groupi_n_5491, csa_tree_add_7_25_groupi_n_5492;
  wire csa_tree_add_7_25_groupi_n_5493, csa_tree_add_7_25_groupi_n_5494, csa_tree_add_7_25_groupi_n_5495, csa_tree_add_7_25_groupi_n_5496, csa_tree_add_7_25_groupi_n_5497, csa_tree_add_7_25_groupi_n_5498, csa_tree_add_7_25_groupi_n_5499, csa_tree_add_7_25_groupi_n_5500;
  wire csa_tree_add_7_25_groupi_n_5501, csa_tree_add_7_25_groupi_n_5502, csa_tree_add_7_25_groupi_n_5503, csa_tree_add_7_25_groupi_n_5504, csa_tree_add_7_25_groupi_n_5505, csa_tree_add_7_25_groupi_n_5506, csa_tree_add_7_25_groupi_n_5507, csa_tree_add_7_25_groupi_n_5508;
  wire csa_tree_add_7_25_groupi_n_5509, csa_tree_add_7_25_groupi_n_5510, csa_tree_add_7_25_groupi_n_5511, csa_tree_add_7_25_groupi_n_5512, csa_tree_add_7_25_groupi_n_5513, csa_tree_add_7_25_groupi_n_5514, csa_tree_add_7_25_groupi_n_5515, csa_tree_add_7_25_groupi_n_5516;
  wire csa_tree_add_7_25_groupi_n_5517, csa_tree_add_7_25_groupi_n_5518, csa_tree_add_7_25_groupi_n_5519, csa_tree_add_7_25_groupi_n_5520, csa_tree_add_7_25_groupi_n_5521, csa_tree_add_7_25_groupi_n_5522, csa_tree_add_7_25_groupi_n_5523, csa_tree_add_7_25_groupi_n_5524;
  wire csa_tree_add_7_25_groupi_n_5525, csa_tree_add_7_25_groupi_n_5526, csa_tree_add_7_25_groupi_n_5527, csa_tree_add_7_25_groupi_n_5528, csa_tree_add_7_25_groupi_n_5529, csa_tree_add_7_25_groupi_n_5530, csa_tree_add_7_25_groupi_n_5531, csa_tree_add_7_25_groupi_n_5532;
  wire csa_tree_add_7_25_groupi_n_5533, csa_tree_add_7_25_groupi_n_5534, csa_tree_add_7_25_groupi_n_5535, csa_tree_add_7_25_groupi_n_5536, csa_tree_add_7_25_groupi_n_5537, csa_tree_add_7_25_groupi_n_5538, csa_tree_add_7_25_groupi_n_5539, csa_tree_add_7_25_groupi_n_5540;
  wire csa_tree_add_7_25_groupi_n_5541, csa_tree_add_7_25_groupi_n_5542, csa_tree_add_7_25_groupi_n_5543, csa_tree_add_7_25_groupi_n_5544, csa_tree_add_7_25_groupi_n_5545, csa_tree_add_7_25_groupi_n_5546, csa_tree_add_7_25_groupi_n_5547, csa_tree_add_7_25_groupi_n_5548;
  wire csa_tree_add_7_25_groupi_n_5549, csa_tree_add_7_25_groupi_n_5550, csa_tree_add_7_25_groupi_n_5551, csa_tree_add_7_25_groupi_n_5552, csa_tree_add_7_25_groupi_n_5553, csa_tree_add_7_25_groupi_n_5554, csa_tree_add_7_25_groupi_n_5555, csa_tree_add_7_25_groupi_n_5556;
  wire csa_tree_add_7_25_groupi_n_5557, csa_tree_add_7_25_groupi_n_5558, csa_tree_add_7_25_groupi_n_5559, csa_tree_add_7_25_groupi_n_5560, csa_tree_add_7_25_groupi_n_5561, csa_tree_add_7_25_groupi_n_5562, csa_tree_add_7_25_groupi_n_5563, csa_tree_add_7_25_groupi_n_5564;
  wire csa_tree_add_7_25_groupi_n_5566, csa_tree_add_7_25_groupi_n_5567, csa_tree_add_7_25_groupi_n_5568, csa_tree_add_7_25_groupi_n_5569, csa_tree_add_7_25_groupi_n_5570, csa_tree_add_7_25_groupi_n_5571, csa_tree_add_7_25_groupi_n_5572, csa_tree_add_7_25_groupi_n_5573;
  wire csa_tree_add_7_25_groupi_n_5574, csa_tree_add_7_25_groupi_n_5575, csa_tree_add_7_25_groupi_n_5576, csa_tree_add_7_25_groupi_n_5577, csa_tree_add_7_25_groupi_n_5578, csa_tree_add_7_25_groupi_n_5579, csa_tree_add_7_25_groupi_n_5580, csa_tree_add_7_25_groupi_n_5581;
  wire csa_tree_add_7_25_groupi_n_5582, csa_tree_add_7_25_groupi_n_5583, csa_tree_add_7_25_groupi_n_5584, csa_tree_add_7_25_groupi_n_5585, csa_tree_add_7_25_groupi_n_5586, csa_tree_add_7_25_groupi_n_5587, csa_tree_add_7_25_groupi_n_5588, csa_tree_add_7_25_groupi_n_5589;
  wire csa_tree_add_7_25_groupi_n_5590, csa_tree_add_7_25_groupi_n_5591, csa_tree_add_7_25_groupi_n_5592, csa_tree_add_7_25_groupi_n_5593, csa_tree_add_7_25_groupi_n_5594, csa_tree_add_7_25_groupi_n_5595, csa_tree_add_7_25_groupi_n_5596, csa_tree_add_7_25_groupi_n_5597;
  wire csa_tree_add_7_25_groupi_n_5598, csa_tree_add_7_25_groupi_n_5599, csa_tree_add_7_25_groupi_n_5600, csa_tree_add_7_25_groupi_n_5601, csa_tree_add_7_25_groupi_n_5602, csa_tree_add_7_25_groupi_n_5603, csa_tree_add_7_25_groupi_n_5604, csa_tree_add_7_25_groupi_n_5605;
  wire csa_tree_add_7_25_groupi_n_5606, csa_tree_add_7_25_groupi_n_5607, csa_tree_add_7_25_groupi_n_5608, csa_tree_add_7_25_groupi_n_5609, csa_tree_add_7_25_groupi_n_5610, csa_tree_add_7_25_groupi_n_5611, csa_tree_add_7_25_groupi_n_5612, csa_tree_add_7_25_groupi_n_5613;
  wire csa_tree_add_7_25_groupi_n_5614, csa_tree_add_7_25_groupi_n_5615, csa_tree_add_7_25_groupi_n_5616, csa_tree_add_7_25_groupi_n_5617, csa_tree_add_7_25_groupi_n_5618, csa_tree_add_7_25_groupi_n_5619, csa_tree_add_7_25_groupi_n_5620, csa_tree_add_7_25_groupi_n_5621;
  wire csa_tree_add_7_25_groupi_n_5622, csa_tree_add_7_25_groupi_n_5623, csa_tree_add_7_25_groupi_n_5624, csa_tree_add_7_25_groupi_n_5625, csa_tree_add_7_25_groupi_n_5626, csa_tree_add_7_25_groupi_n_5627, csa_tree_add_7_25_groupi_n_5628, csa_tree_add_7_25_groupi_n_5629;
  wire csa_tree_add_7_25_groupi_n_5630, csa_tree_add_7_25_groupi_n_5631, csa_tree_add_7_25_groupi_n_5632, csa_tree_add_7_25_groupi_n_5633, csa_tree_add_7_25_groupi_n_5634, csa_tree_add_7_25_groupi_n_5635, csa_tree_add_7_25_groupi_n_5636, csa_tree_add_7_25_groupi_n_5637;
  wire csa_tree_add_7_25_groupi_n_5638, csa_tree_add_7_25_groupi_n_5639, csa_tree_add_7_25_groupi_n_5640, csa_tree_add_7_25_groupi_n_5641, csa_tree_add_7_25_groupi_n_5642, csa_tree_add_7_25_groupi_n_5643, csa_tree_add_7_25_groupi_n_5644, csa_tree_add_7_25_groupi_n_5645;
  wire csa_tree_add_7_25_groupi_n_5646, csa_tree_add_7_25_groupi_n_5647, csa_tree_add_7_25_groupi_n_5648, csa_tree_add_7_25_groupi_n_5649, csa_tree_add_7_25_groupi_n_5650, csa_tree_add_7_25_groupi_n_5651, csa_tree_add_7_25_groupi_n_5652, csa_tree_add_7_25_groupi_n_5653;
  wire csa_tree_add_7_25_groupi_n_5654, csa_tree_add_7_25_groupi_n_5655, csa_tree_add_7_25_groupi_n_5656, csa_tree_add_7_25_groupi_n_5657, csa_tree_add_7_25_groupi_n_5658, csa_tree_add_7_25_groupi_n_5659, csa_tree_add_7_25_groupi_n_5660, csa_tree_add_7_25_groupi_n_5661;
  wire csa_tree_add_7_25_groupi_n_5662, csa_tree_add_7_25_groupi_n_5663, csa_tree_add_7_25_groupi_n_5664, csa_tree_add_7_25_groupi_n_5665, csa_tree_add_7_25_groupi_n_5666, csa_tree_add_7_25_groupi_n_5667, csa_tree_add_7_25_groupi_n_5668, csa_tree_add_7_25_groupi_n_5669;
  wire csa_tree_add_7_25_groupi_n_5670, csa_tree_add_7_25_groupi_n_5671, csa_tree_add_7_25_groupi_n_5672, csa_tree_add_7_25_groupi_n_5673, csa_tree_add_7_25_groupi_n_5674, csa_tree_add_7_25_groupi_n_5675, csa_tree_add_7_25_groupi_n_5676, csa_tree_add_7_25_groupi_n_5677;
  wire csa_tree_add_7_25_groupi_n_5678, csa_tree_add_7_25_groupi_n_5679, csa_tree_add_7_25_groupi_n_5680, csa_tree_add_7_25_groupi_n_5682, csa_tree_add_7_25_groupi_n_5683, csa_tree_add_7_25_groupi_n_5684, csa_tree_add_7_25_groupi_n_5685, csa_tree_add_7_25_groupi_n_5686;
  wire csa_tree_add_7_25_groupi_n_5687, csa_tree_add_7_25_groupi_n_5688, csa_tree_add_7_25_groupi_n_5689, csa_tree_add_7_25_groupi_n_5690, csa_tree_add_7_25_groupi_n_5691, csa_tree_add_7_25_groupi_n_5692, csa_tree_add_7_25_groupi_n_5693, csa_tree_add_7_25_groupi_n_5694;
  wire csa_tree_add_7_25_groupi_n_5695, csa_tree_add_7_25_groupi_n_5696, csa_tree_add_7_25_groupi_n_5697, csa_tree_add_7_25_groupi_n_5698, csa_tree_add_7_25_groupi_n_5699, csa_tree_add_7_25_groupi_n_5700, csa_tree_add_7_25_groupi_n_5701, csa_tree_add_7_25_groupi_n_5702;
  wire csa_tree_add_7_25_groupi_n_5703, csa_tree_add_7_25_groupi_n_5704, csa_tree_add_7_25_groupi_n_5705, csa_tree_add_7_25_groupi_n_5706, csa_tree_add_7_25_groupi_n_5707, csa_tree_add_7_25_groupi_n_5708, csa_tree_add_7_25_groupi_n_5709, csa_tree_add_7_25_groupi_n_5710;
  wire csa_tree_add_7_25_groupi_n_5711, csa_tree_add_7_25_groupi_n_5712, csa_tree_add_7_25_groupi_n_5713, csa_tree_add_7_25_groupi_n_5714, csa_tree_add_7_25_groupi_n_5715, csa_tree_add_7_25_groupi_n_5716, csa_tree_add_7_25_groupi_n_5717, csa_tree_add_7_25_groupi_n_5718;
  wire csa_tree_add_7_25_groupi_n_5719, csa_tree_add_7_25_groupi_n_5720, csa_tree_add_7_25_groupi_n_5721, csa_tree_add_7_25_groupi_n_5722, csa_tree_add_7_25_groupi_n_5723, csa_tree_add_7_25_groupi_n_5724, csa_tree_add_7_25_groupi_n_5725, csa_tree_add_7_25_groupi_n_5726;
  wire csa_tree_add_7_25_groupi_n_5727, csa_tree_add_7_25_groupi_n_5728, csa_tree_add_7_25_groupi_n_5729, csa_tree_add_7_25_groupi_n_5730, csa_tree_add_7_25_groupi_n_5731, csa_tree_add_7_25_groupi_n_5732, csa_tree_add_7_25_groupi_n_5733, csa_tree_add_7_25_groupi_n_5734;
  wire csa_tree_add_7_25_groupi_n_5735, csa_tree_add_7_25_groupi_n_5736, csa_tree_add_7_25_groupi_n_5737, csa_tree_add_7_25_groupi_n_5738, csa_tree_add_7_25_groupi_n_5739, csa_tree_add_7_25_groupi_n_5740, csa_tree_add_7_25_groupi_n_5741, csa_tree_add_7_25_groupi_n_5742;
  wire csa_tree_add_7_25_groupi_n_5743, csa_tree_add_7_25_groupi_n_5744, csa_tree_add_7_25_groupi_n_5745, csa_tree_add_7_25_groupi_n_5746, csa_tree_add_7_25_groupi_n_5747, csa_tree_add_7_25_groupi_n_5748, csa_tree_add_7_25_groupi_n_5749, csa_tree_add_7_25_groupi_n_5750;
  wire csa_tree_add_7_25_groupi_n_5751, csa_tree_add_7_25_groupi_n_5752, csa_tree_add_7_25_groupi_n_5753, csa_tree_add_7_25_groupi_n_5754, csa_tree_add_7_25_groupi_n_5755, csa_tree_add_7_25_groupi_n_5756, csa_tree_add_7_25_groupi_n_5757, csa_tree_add_7_25_groupi_n_5758;
  wire csa_tree_add_7_25_groupi_n_5759, csa_tree_add_7_25_groupi_n_5760, csa_tree_add_7_25_groupi_n_5761, csa_tree_add_7_25_groupi_n_5762, csa_tree_add_7_25_groupi_n_5763, csa_tree_add_7_25_groupi_n_5764, csa_tree_add_7_25_groupi_n_5765, csa_tree_add_7_25_groupi_n_5766;
  wire csa_tree_add_7_25_groupi_n_5767, csa_tree_add_7_25_groupi_n_5768, csa_tree_add_7_25_groupi_n_5769, csa_tree_add_7_25_groupi_n_5770, csa_tree_add_7_25_groupi_n_5771, csa_tree_add_7_25_groupi_n_5772, csa_tree_add_7_25_groupi_n_5773, csa_tree_add_7_25_groupi_n_5774;
  wire csa_tree_add_7_25_groupi_n_5775, csa_tree_add_7_25_groupi_n_5776, csa_tree_add_7_25_groupi_n_5777, csa_tree_add_7_25_groupi_n_5778, csa_tree_add_7_25_groupi_n_5779, csa_tree_add_7_25_groupi_n_5780, csa_tree_add_7_25_groupi_n_5781, csa_tree_add_7_25_groupi_n_5782;
  wire csa_tree_add_7_25_groupi_n_5783, csa_tree_add_7_25_groupi_n_5784, csa_tree_add_7_25_groupi_n_5785, csa_tree_add_7_25_groupi_n_5786, csa_tree_add_7_25_groupi_n_5787, csa_tree_add_7_25_groupi_n_5788, csa_tree_add_7_25_groupi_n_5789, csa_tree_add_7_25_groupi_n_5790;
  wire csa_tree_add_7_25_groupi_n_5791, csa_tree_add_7_25_groupi_n_5792, csa_tree_add_7_25_groupi_n_5793, csa_tree_add_7_25_groupi_n_5794, csa_tree_add_7_25_groupi_n_5795, csa_tree_add_7_25_groupi_n_5796, csa_tree_add_7_25_groupi_n_5797, csa_tree_add_7_25_groupi_n_5798;
  wire csa_tree_add_7_25_groupi_n_5799, csa_tree_add_7_25_groupi_n_5800, csa_tree_add_7_25_groupi_n_5802, csa_tree_add_7_25_groupi_n_5803, csa_tree_add_7_25_groupi_n_5804, csa_tree_add_7_25_groupi_n_5805, csa_tree_add_7_25_groupi_n_5806, csa_tree_add_7_25_groupi_n_5807;
  wire csa_tree_add_7_25_groupi_n_5808, csa_tree_add_7_25_groupi_n_5809, csa_tree_add_7_25_groupi_n_5810, csa_tree_add_7_25_groupi_n_5811, csa_tree_add_7_25_groupi_n_5812, csa_tree_add_7_25_groupi_n_5813, csa_tree_add_7_25_groupi_n_5814, csa_tree_add_7_25_groupi_n_5815;
  wire csa_tree_add_7_25_groupi_n_5816, csa_tree_add_7_25_groupi_n_5817, csa_tree_add_7_25_groupi_n_5818, csa_tree_add_7_25_groupi_n_5819, csa_tree_add_7_25_groupi_n_5820, csa_tree_add_7_25_groupi_n_5821, csa_tree_add_7_25_groupi_n_5822, csa_tree_add_7_25_groupi_n_5823;
  wire csa_tree_add_7_25_groupi_n_5824, csa_tree_add_7_25_groupi_n_5825, csa_tree_add_7_25_groupi_n_5826, csa_tree_add_7_25_groupi_n_5827, csa_tree_add_7_25_groupi_n_5828, csa_tree_add_7_25_groupi_n_5829, csa_tree_add_7_25_groupi_n_5830, csa_tree_add_7_25_groupi_n_5831;
  wire csa_tree_add_7_25_groupi_n_5832, csa_tree_add_7_25_groupi_n_5833, csa_tree_add_7_25_groupi_n_5834, csa_tree_add_7_25_groupi_n_5835, csa_tree_add_7_25_groupi_n_5836, csa_tree_add_7_25_groupi_n_5837, csa_tree_add_7_25_groupi_n_5838, csa_tree_add_7_25_groupi_n_5839;
  wire csa_tree_add_7_25_groupi_n_5840, csa_tree_add_7_25_groupi_n_5841, csa_tree_add_7_25_groupi_n_5842, csa_tree_add_7_25_groupi_n_5843, csa_tree_add_7_25_groupi_n_5844, csa_tree_add_7_25_groupi_n_5845, csa_tree_add_7_25_groupi_n_5846, csa_tree_add_7_25_groupi_n_5847;
  wire csa_tree_add_7_25_groupi_n_5848, csa_tree_add_7_25_groupi_n_5849, csa_tree_add_7_25_groupi_n_5850, csa_tree_add_7_25_groupi_n_5851, csa_tree_add_7_25_groupi_n_5852, csa_tree_add_7_25_groupi_n_5853, csa_tree_add_7_25_groupi_n_5854, csa_tree_add_7_25_groupi_n_5855;
  wire csa_tree_add_7_25_groupi_n_5856, csa_tree_add_7_25_groupi_n_5857, csa_tree_add_7_25_groupi_n_5858, csa_tree_add_7_25_groupi_n_5859, csa_tree_add_7_25_groupi_n_5860, csa_tree_add_7_25_groupi_n_5861, csa_tree_add_7_25_groupi_n_5862, csa_tree_add_7_25_groupi_n_5863;
  wire csa_tree_add_7_25_groupi_n_5864, csa_tree_add_7_25_groupi_n_5865, csa_tree_add_7_25_groupi_n_5866, csa_tree_add_7_25_groupi_n_5867, csa_tree_add_7_25_groupi_n_5868, csa_tree_add_7_25_groupi_n_5869, csa_tree_add_7_25_groupi_n_5870, csa_tree_add_7_25_groupi_n_5871;
  wire csa_tree_add_7_25_groupi_n_5872, csa_tree_add_7_25_groupi_n_5873, csa_tree_add_7_25_groupi_n_5874, csa_tree_add_7_25_groupi_n_5875, csa_tree_add_7_25_groupi_n_5876, csa_tree_add_7_25_groupi_n_5877, csa_tree_add_7_25_groupi_n_5878, csa_tree_add_7_25_groupi_n_5879;
  wire csa_tree_add_7_25_groupi_n_5880, csa_tree_add_7_25_groupi_n_5881, csa_tree_add_7_25_groupi_n_5882, csa_tree_add_7_25_groupi_n_5883, csa_tree_add_7_25_groupi_n_5884, csa_tree_add_7_25_groupi_n_5885, csa_tree_add_7_25_groupi_n_5886, csa_tree_add_7_25_groupi_n_5887;
  wire csa_tree_add_7_25_groupi_n_5888, csa_tree_add_7_25_groupi_n_5889, csa_tree_add_7_25_groupi_n_5890, csa_tree_add_7_25_groupi_n_5891, csa_tree_add_7_25_groupi_n_5892, csa_tree_add_7_25_groupi_n_5893, csa_tree_add_7_25_groupi_n_5894, csa_tree_add_7_25_groupi_n_5895;
  wire csa_tree_add_7_25_groupi_n_5896, csa_tree_add_7_25_groupi_n_5898, csa_tree_add_7_25_groupi_n_5899, csa_tree_add_7_25_groupi_n_5900, csa_tree_add_7_25_groupi_n_5901, csa_tree_add_7_25_groupi_n_5902, csa_tree_add_7_25_groupi_n_5903, csa_tree_add_7_25_groupi_n_5904;
  wire csa_tree_add_7_25_groupi_n_5905, csa_tree_add_7_25_groupi_n_5906, csa_tree_add_7_25_groupi_n_5907, csa_tree_add_7_25_groupi_n_5908, csa_tree_add_7_25_groupi_n_5909, csa_tree_add_7_25_groupi_n_5910, csa_tree_add_7_25_groupi_n_5911, csa_tree_add_7_25_groupi_n_5912;
  wire csa_tree_add_7_25_groupi_n_5913, csa_tree_add_7_25_groupi_n_5914, csa_tree_add_7_25_groupi_n_5915, csa_tree_add_7_25_groupi_n_5916, csa_tree_add_7_25_groupi_n_5917, csa_tree_add_7_25_groupi_n_5918, csa_tree_add_7_25_groupi_n_5919, csa_tree_add_7_25_groupi_n_5920;
  wire csa_tree_add_7_25_groupi_n_5921, csa_tree_add_7_25_groupi_n_5922, csa_tree_add_7_25_groupi_n_5923, csa_tree_add_7_25_groupi_n_5924, csa_tree_add_7_25_groupi_n_5925, csa_tree_add_7_25_groupi_n_5926, csa_tree_add_7_25_groupi_n_5927, csa_tree_add_7_25_groupi_n_5928;
  wire csa_tree_add_7_25_groupi_n_5929, csa_tree_add_7_25_groupi_n_5930, csa_tree_add_7_25_groupi_n_5931, csa_tree_add_7_25_groupi_n_5932, csa_tree_add_7_25_groupi_n_5933, csa_tree_add_7_25_groupi_n_5934, csa_tree_add_7_25_groupi_n_5935, csa_tree_add_7_25_groupi_n_5936;
  wire csa_tree_add_7_25_groupi_n_5937, csa_tree_add_7_25_groupi_n_5938, csa_tree_add_7_25_groupi_n_5939, csa_tree_add_7_25_groupi_n_5940, csa_tree_add_7_25_groupi_n_5941, csa_tree_add_7_25_groupi_n_5942, csa_tree_add_7_25_groupi_n_5943, csa_tree_add_7_25_groupi_n_5944;
  wire csa_tree_add_7_25_groupi_n_5945, csa_tree_add_7_25_groupi_n_5946, csa_tree_add_7_25_groupi_n_5947, csa_tree_add_7_25_groupi_n_5948, csa_tree_add_7_25_groupi_n_5949, csa_tree_add_7_25_groupi_n_5950, csa_tree_add_7_25_groupi_n_5951, csa_tree_add_7_25_groupi_n_5952;
  wire csa_tree_add_7_25_groupi_n_5953, csa_tree_add_7_25_groupi_n_5954, csa_tree_add_7_25_groupi_n_5955, csa_tree_add_7_25_groupi_n_5956, csa_tree_add_7_25_groupi_n_5957, csa_tree_add_7_25_groupi_n_5958, csa_tree_add_7_25_groupi_n_5959, csa_tree_add_7_25_groupi_n_5960;
  wire csa_tree_add_7_25_groupi_n_5961, csa_tree_add_7_25_groupi_n_5962, csa_tree_add_7_25_groupi_n_5963, csa_tree_add_7_25_groupi_n_5964, csa_tree_add_7_25_groupi_n_5965, csa_tree_add_7_25_groupi_n_5966, csa_tree_add_7_25_groupi_n_5967, csa_tree_add_7_25_groupi_n_5968;
  wire csa_tree_add_7_25_groupi_n_5969, csa_tree_add_7_25_groupi_n_5970, csa_tree_add_7_25_groupi_n_5971, csa_tree_add_7_25_groupi_n_5972, csa_tree_add_7_25_groupi_n_5973, csa_tree_add_7_25_groupi_n_5974, csa_tree_add_7_25_groupi_n_5975, csa_tree_add_7_25_groupi_n_5976;
  wire csa_tree_add_7_25_groupi_n_5977, csa_tree_add_7_25_groupi_n_5978, csa_tree_add_7_25_groupi_n_5979, csa_tree_add_7_25_groupi_n_5980, csa_tree_add_7_25_groupi_n_5981, csa_tree_add_7_25_groupi_n_5982, csa_tree_add_7_25_groupi_n_5983, csa_tree_add_7_25_groupi_n_5984;
  wire csa_tree_add_7_25_groupi_n_5985, csa_tree_add_7_25_groupi_n_5986, csa_tree_add_7_25_groupi_n_5987, csa_tree_add_7_25_groupi_n_5988, csa_tree_add_7_25_groupi_n_5989, csa_tree_add_7_25_groupi_n_5990, csa_tree_add_7_25_groupi_n_5991, csa_tree_add_7_25_groupi_n_5992;
  wire csa_tree_add_7_25_groupi_n_5993, csa_tree_add_7_25_groupi_n_5994, csa_tree_add_7_25_groupi_n_5995, csa_tree_add_7_25_groupi_n_5996, csa_tree_add_7_25_groupi_n_5997, csa_tree_add_7_25_groupi_n_5998, csa_tree_add_7_25_groupi_n_5999, csa_tree_add_7_25_groupi_n_6000;
  wire csa_tree_add_7_25_groupi_n_6001, csa_tree_add_7_25_groupi_n_6002, csa_tree_add_7_25_groupi_n_6003, csa_tree_add_7_25_groupi_n_6004, csa_tree_add_7_25_groupi_n_6005, csa_tree_add_7_25_groupi_n_6006, csa_tree_add_7_25_groupi_n_6007, csa_tree_add_7_25_groupi_n_6008;
  wire csa_tree_add_7_25_groupi_n_6009, csa_tree_add_7_25_groupi_n_6010, csa_tree_add_7_25_groupi_n_6011, csa_tree_add_7_25_groupi_n_6013, csa_tree_add_7_25_groupi_n_6014, csa_tree_add_7_25_groupi_n_6015, csa_tree_add_7_25_groupi_n_6016, csa_tree_add_7_25_groupi_n_6017;
  wire csa_tree_add_7_25_groupi_n_6018, csa_tree_add_7_25_groupi_n_6019, csa_tree_add_7_25_groupi_n_6020, csa_tree_add_7_25_groupi_n_6021, csa_tree_add_7_25_groupi_n_6022, csa_tree_add_7_25_groupi_n_6023, csa_tree_add_7_25_groupi_n_6024, csa_tree_add_7_25_groupi_n_6025;
  wire csa_tree_add_7_25_groupi_n_6026, csa_tree_add_7_25_groupi_n_6027, csa_tree_add_7_25_groupi_n_6028, csa_tree_add_7_25_groupi_n_6029, csa_tree_add_7_25_groupi_n_6030, csa_tree_add_7_25_groupi_n_6031, csa_tree_add_7_25_groupi_n_6032, csa_tree_add_7_25_groupi_n_6033;
  wire csa_tree_add_7_25_groupi_n_6034, csa_tree_add_7_25_groupi_n_6035, csa_tree_add_7_25_groupi_n_6036, csa_tree_add_7_25_groupi_n_6037, csa_tree_add_7_25_groupi_n_6038, csa_tree_add_7_25_groupi_n_6039, csa_tree_add_7_25_groupi_n_6040, csa_tree_add_7_25_groupi_n_6041;
  wire csa_tree_add_7_25_groupi_n_6042, csa_tree_add_7_25_groupi_n_6043, csa_tree_add_7_25_groupi_n_6044, csa_tree_add_7_25_groupi_n_6045, csa_tree_add_7_25_groupi_n_6046, csa_tree_add_7_25_groupi_n_6047, csa_tree_add_7_25_groupi_n_6048, csa_tree_add_7_25_groupi_n_6049;
  wire csa_tree_add_7_25_groupi_n_6050, csa_tree_add_7_25_groupi_n_6051, csa_tree_add_7_25_groupi_n_6052, csa_tree_add_7_25_groupi_n_6053, csa_tree_add_7_25_groupi_n_6054, csa_tree_add_7_25_groupi_n_6055, csa_tree_add_7_25_groupi_n_6056, csa_tree_add_7_25_groupi_n_6057;
  wire csa_tree_add_7_25_groupi_n_6058, csa_tree_add_7_25_groupi_n_6059, csa_tree_add_7_25_groupi_n_6060, csa_tree_add_7_25_groupi_n_6061, csa_tree_add_7_25_groupi_n_6062, csa_tree_add_7_25_groupi_n_6063, csa_tree_add_7_25_groupi_n_6064, csa_tree_add_7_25_groupi_n_6065;
  wire csa_tree_add_7_25_groupi_n_6066, csa_tree_add_7_25_groupi_n_6067, csa_tree_add_7_25_groupi_n_6068, csa_tree_add_7_25_groupi_n_6069, csa_tree_add_7_25_groupi_n_6070, csa_tree_add_7_25_groupi_n_6071, csa_tree_add_7_25_groupi_n_6072, csa_tree_add_7_25_groupi_n_6073;
  wire csa_tree_add_7_25_groupi_n_6074, csa_tree_add_7_25_groupi_n_6075, csa_tree_add_7_25_groupi_n_6076, csa_tree_add_7_25_groupi_n_6077, csa_tree_add_7_25_groupi_n_6078, csa_tree_add_7_25_groupi_n_6079, csa_tree_add_7_25_groupi_n_6080, csa_tree_add_7_25_groupi_n_6081;
  wire csa_tree_add_7_25_groupi_n_6082, csa_tree_add_7_25_groupi_n_6083, csa_tree_add_7_25_groupi_n_6084, csa_tree_add_7_25_groupi_n_6085, csa_tree_add_7_25_groupi_n_6086, csa_tree_add_7_25_groupi_n_6087, csa_tree_add_7_25_groupi_n_6088, csa_tree_add_7_25_groupi_n_6089;
  wire csa_tree_add_7_25_groupi_n_6090, csa_tree_add_7_25_groupi_n_6091, csa_tree_add_7_25_groupi_n_6092, csa_tree_add_7_25_groupi_n_6093, csa_tree_add_7_25_groupi_n_6094, csa_tree_add_7_25_groupi_n_6095, csa_tree_add_7_25_groupi_n_6096, csa_tree_add_7_25_groupi_n_6097;
  wire csa_tree_add_7_25_groupi_n_6098, csa_tree_add_7_25_groupi_n_6099, csa_tree_add_7_25_groupi_n_6100, csa_tree_add_7_25_groupi_n_6101, csa_tree_add_7_25_groupi_n_6102, csa_tree_add_7_25_groupi_n_6103, csa_tree_add_7_25_groupi_n_6104, csa_tree_add_7_25_groupi_n_6105;
  wire csa_tree_add_7_25_groupi_n_6106, csa_tree_add_7_25_groupi_n_6107, csa_tree_add_7_25_groupi_n_6108, csa_tree_add_7_25_groupi_n_6109, csa_tree_add_7_25_groupi_n_6110, csa_tree_add_7_25_groupi_n_6111, csa_tree_add_7_25_groupi_n_6112, csa_tree_add_7_25_groupi_n_6113;
  wire csa_tree_add_7_25_groupi_n_6114, csa_tree_add_7_25_groupi_n_6115, csa_tree_add_7_25_groupi_n_6116, csa_tree_add_7_25_groupi_n_6117, csa_tree_add_7_25_groupi_n_6118, csa_tree_add_7_25_groupi_n_6119, csa_tree_add_7_25_groupi_n_6120, csa_tree_add_7_25_groupi_n_6121;
  wire csa_tree_add_7_25_groupi_n_6122, csa_tree_add_7_25_groupi_n_6124, csa_tree_add_7_25_groupi_n_6125, csa_tree_add_7_25_groupi_n_6126, csa_tree_add_7_25_groupi_n_6127, csa_tree_add_7_25_groupi_n_6128, csa_tree_add_7_25_groupi_n_6129, csa_tree_add_7_25_groupi_n_6130;
  wire csa_tree_add_7_25_groupi_n_6131, csa_tree_add_7_25_groupi_n_6132, csa_tree_add_7_25_groupi_n_6133, csa_tree_add_7_25_groupi_n_6134, csa_tree_add_7_25_groupi_n_6135, csa_tree_add_7_25_groupi_n_6136, csa_tree_add_7_25_groupi_n_6137, csa_tree_add_7_25_groupi_n_6138;
  wire csa_tree_add_7_25_groupi_n_6139, csa_tree_add_7_25_groupi_n_6140, csa_tree_add_7_25_groupi_n_6141, csa_tree_add_7_25_groupi_n_6142, csa_tree_add_7_25_groupi_n_6143, csa_tree_add_7_25_groupi_n_6144, csa_tree_add_7_25_groupi_n_6145, csa_tree_add_7_25_groupi_n_6146;
  wire csa_tree_add_7_25_groupi_n_6147, csa_tree_add_7_25_groupi_n_6148, csa_tree_add_7_25_groupi_n_6149, csa_tree_add_7_25_groupi_n_6150, csa_tree_add_7_25_groupi_n_6151, csa_tree_add_7_25_groupi_n_6152, csa_tree_add_7_25_groupi_n_6153, csa_tree_add_7_25_groupi_n_6154;
  wire csa_tree_add_7_25_groupi_n_6155, csa_tree_add_7_25_groupi_n_6156, csa_tree_add_7_25_groupi_n_6157, csa_tree_add_7_25_groupi_n_6158, csa_tree_add_7_25_groupi_n_6159, csa_tree_add_7_25_groupi_n_6160, csa_tree_add_7_25_groupi_n_6161, csa_tree_add_7_25_groupi_n_6162;
  wire csa_tree_add_7_25_groupi_n_6163, csa_tree_add_7_25_groupi_n_6164, csa_tree_add_7_25_groupi_n_6165, csa_tree_add_7_25_groupi_n_6166, csa_tree_add_7_25_groupi_n_6167, csa_tree_add_7_25_groupi_n_6168, csa_tree_add_7_25_groupi_n_6169, csa_tree_add_7_25_groupi_n_6170;
  wire csa_tree_add_7_25_groupi_n_6171, csa_tree_add_7_25_groupi_n_6172, csa_tree_add_7_25_groupi_n_6173, csa_tree_add_7_25_groupi_n_6174, csa_tree_add_7_25_groupi_n_6175, csa_tree_add_7_25_groupi_n_6176, csa_tree_add_7_25_groupi_n_6177, csa_tree_add_7_25_groupi_n_6178;
  wire csa_tree_add_7_25_groupi_n_6179, csa_tree_add_7_25_groupi_n_6180, csa_tree_add_7_25_groupi_n_6181, csa_tree_add_7_25_groupi_n_6182, csa_tree_add_7_25_groupi_n_6183, csa_tree_add_7_25_groupi_n_6184, csa_tree_add_7_25_groupi_n_6185, csa_tree_add_7_25_groupi_n_6186;
  wire csa_tree_add_7_25_groupi_n_6187, csa_tree_add_7_25_groupi_n_6188, csa_tree_add_7_25_groupi_n_6189, csa_tree_add_7_25_groupi_n_6190, csa_tree_add_7_25_groupi_n_6191, csa_tree_add_7_25_groupi_n_6192, csa_tree_add_7_25_groupi_n_6193, csa_tree_add_7_25_groupi_n_6194;
  wire csa_tree_add_7_25_groupi_n_6195, csa_tree_add_7_25_groupi_n_6196, csa_tree_add_7_25_groupi_n_6197, csa_tree_add_7_25_groupi_n_6198, csa_tree_add_7_25_groupi_n_6199, csa_tree_add_7_25_groupi_n_6200, csa_tree_add_7_25_groupi_n_6201, csa_tree_add_7_25_groupi_n_6202;
  wire csa_tree_add_7_25_groupi_n_6203, csa_tree_add_7_25_groupi_n_6204, csa_tree_add_7_25_groupi_n_6205, csa_tree_add_7_25_groupi_n_6206, csa_tree_add_7_25_groupi_n_6207, csa_tree_add_7_25_groupi_n_6208, csa_tree_add_7_25_groupi_n_6210, csa_tree_add_7_25_groupi_n_6211;
  wire csa_tree_add_7_25_groupi_n_6212, csa_tree_add_7_25_groupi_n_6213, csa_tree_add_7_25_groupi_n_6214, csa_tree_add_7_25_groupi_n_6215, csa_tree_add_7_25_groupi_n_6216, csa_tree_add_7_25_groupi_n_6217, csa_tree_add_7_25_groupi_n_6218, csa_tree_add_7_25_groupi_n_6219;
  wire csa_tree_add_7_25_groupi_n_6220, csa_tree_add_7_25_groupi_n_6221, csa_tree_add_7_25_groupi_n_6222, csa_tree_add_7_25_groupi_n_6223, csa_tree_add_7_25_groupi_n_6224, csa_tree_add_7_25_groupi_n_6225, csa_tree_add_7_25_groupi_n_6226, csa_tree_add_7_25_groupi_n_6227;
  wire csa_tree_add_7_25_groupi_n_6228, csa_tree_add_7_25_groupi_n_6229, csa_tree_add_7_25_groupi_n_6230, csa_tree_add_7_25_groupi_n_6231, csa_tree_add_7_25_groupi_n_6232, csa_tree_add_7_25_groupi_n_6233, csa_tree_add_7_25_groupi_n_6234, csa_tree_add_7_25_groupi_n_6235;
  wire csa_tree_add_7_25_groupi_n_6236, csa_tree_add_7_25_groupi_n_6237, csa_tree_add_7_25_groupi_n_6238, csa_tree_add_7_25_groupi_n_6239, csa_tree_add_7_25_groupi_n_6240, csa_tree_add_7_25_groupi_n_6241, csa_tree_add_7_25_groupi_n_6242, csa_tree_add_7_25_groupi_n_6243;
  wire csa_tree_add_7_25_groupi_n_6244, csa_tree_add_7_25_groupi_n_6245, csa_tree_add_7_25_groupi_n_6246, csa_tree_add_7_25_groupi_n_6247, csa_tree_add_7_25_groupi_n_6248, csa_tree_add_7_25_groupi_n_6249, csa_tree_add_7_25_groupi_n_6250, csa_tree_add_7_25_groupi_n_6251;
  wire csa_tree_add_7_25_groupi_n_6252, csa_tree_add_7_25_groupi_n_6253, csa_tree_add_7_25_groupi_n_6254, csa_tree_add_7_25_groupi_n_6255, csa_tree_add_7_25_groupi_n_6256, csa_tree_add_7_25_groupi_n_6257, csa_tree_add_7_25_groupi_n_6258, csa_tree_add_7_25_groupi_n_6259;
  wire csa_tree_add_7_25_groupi_n_6260, csa_tree_add_7_25_groupi_n_6261, csa_tree_add_7_25_groupi_n_6262, csa_tree_add_7_25_groupi_n_6263, csa_tree_add_7_25_groupi_n_6264, csa_tree_add_7_25_groupi_n_6265, csa_tree_add_7_25_groupi_n_6266, csa_tree_add_7_25_groupi_n_6267;
  wire csa_tree_add_7_25_groupi_n_6268, csa_tree_add_7_25_groupi_n_6269, csa_tree_add_7_25_groupi_n_6270, csa_tree_add_7_25_groupi_n_6271, csa_tree_add_7_25_groupi_n_6272, csa_tree_add_7_25_groupi_n_6273, csa_tree_add_7_25_groupi_n_6274, csa_tree_add_7_25_groupi_n_6275;
  wire csa_tree_add_7_25_groupi_n_6276, csa_tree_add_7_25_groupi_n_6277, csa_tree_add_7_25_groupi_n_6278, csa_tree_add_7_25_groupi_n_6279, csa_tree_add_7_25_groupi_n_6280, csa_tree_add_7_25_groupi_n_6281, csa_tree_add_7_25_groupi_n_6282, csa_tree_add_7_25_groupi_n_6283;
  wire csa_tree_add_7_25_groupi_n_6284, csa_tree_add_7_25_groupi_n_6285, csa_tree_add_7_25_groupi_n_6286, csa_tree_add_7_25_groupi_n_6287, csa_tree_add_7_25_groupi_n_6288, csa_tree_add_7_25_groupi_n_6289, csa_tree_add_7_25_groupi_n_6290, csa_tree_add_7_25_groupi_n_6291;
  wire csa_tree_add_7_25_groupi_n_6292, csa_tree_add_7_25_groupi_n_6293, csa_tree_add_7_25_groupi_n_6294, csa_tree_add_7_25_groupi_n_6295, csa_tree_add_7_25_groupi_n_6296, csa_tree_add_7_25_groupi_n_6297, csa_tree_add_7_25_groupi_n_6298, csa_tree_add_7_25_groupi_n_6299;
  wire csa_tree_add_7_25_groupi_n_6300, csa_tree_add_7_25_groupi_n_6301, csa_tree_add_7_25_groupi_n_6302, csa_tree_add_7_25_groupi_n_6303, csa_tree_add_7_25_groupi_n_6304, csa_tree_add_7_25_groupi_n_6305, csa_tree_add_7_25_groupi_n_6306, csa_tree_add_7_25_groupi_n_6307;
  wire csa_tree_add_7_25_groupi_n_6308, csa_tree_add_7_25_groupi_n_6309, csa_tree_add_7_25_groupi_n_6310, csa_tree_add_7_25_groupi_n_6311, csa_tree_add_7_25_groupi_n_6312, csa_tree_add_7_25_groupi_n_6313, csa_tree_add_7_25_groupi_n_6315, csa_tree_add_7_25_groupi_n_6316;
  wire csa_tree_add_7_25_groupi_n_6317, csa_tree_add_7_25_groupi_n_6318, csa_tree_add_7_25_groupi_n_6319, csa_tree_add_7_25_groupi_n_6320, csa_tree_add_7_25_groupi_n_6321, csa_tree_add_7_25_groupi_n_6322, csa_tree_add_7_25_groupi_n_6323, csa_tree_add_7_25_groupi_n_6324;
  wire csa_tree_add_7_25_groupi_n_6325, csa_tree_add_7_25_groupi_n_6326, csa_tree_add_7_25_groupi_n_6327, csa_tree_add_7_25_groupi_n_6328, csa_tree_add_7_25_groupi_n_6329, csa_tree_add_7_25_groupi_n_6330, csa_tree_add_7_25_groupi_n_6331, csa_tree_add_7_25_groupi_n_6332;
  wire csa_tree_add_7_25_groupi_n_6333, csa_tree_add_7_25_groupi_n_6334, csa_tree_add_7_25_groupi_n_6335, csa_tree_add_7_25_groupi_n_6336, csa_tree_add_7_25_groupi_n_6337, csa_tree_add_7_25_groupi_n_6338, csa_tree_add_7_25_groupi_n_6339, csa_tree_add_7_25_groupi_n_6340;
  wire csa_tree_add_7_25_groupi_n_6341, csa_tree_add_7_25_groupi_n_6342, csa_tree_add_7_25_groupi_n_6343, csa_tree_add_7_25_groupi_n_6344, csa_tree_add_7_25_groupi_n_6345, csa_tree_add_7_25_groupi_n_6346, csa_tree_add_7_25_groupi_n_6347, csa_tree_add_7_25_groupi_n_6348;
  wire csa_tree_add_7_25_groupi_n_6349, csa_tree_add_7_25_groupi_n_6350, csa_tree_add_7_25_groupi_n_6351, csa_tree_add_7_25_groupi_n_6352, csa_tree_add_7_25_groupi_n_6353, csa_tree_add_7_25_groupi_n_6354, csa_tree_add_7_25_groupi_n_6355, csa_tree_add_7_25_groupi_n_6356;
  wire csa_tree_add_7_25_groupi_n_6357, csa_tree_add_7_25_groupi_n_6358, csa_tree_add_7_25_groupi_n_6359, csa_tree_add_7_25_groupi_n_6360, csa_tree_add_7_25_groupi_n_6361, csa_tree_add_7_25_groupi_n_6362, csa_tree_add_7_25_groupi_n_6363, csa_tree_add_7_25_groupi_n_6364;
  wire csa_tree_add_7_25_groupi_n_6365, csa_tree_add_7_25_groupi_n_6366, csa_tree_add_7_25_groupi_n_6367, csa_tree_add_7_25_groupi_n_6368, csa_tree_add_7_25_groupi_n_6369, csa_tree_add_7_25_groupi_n_6370, csa_tree_add_7_25_groupi_n_6371, csa_tree_add_7_25_groupi_n_6372;
  wire csa_tree_add_7_25_groupi_n_6373, csa_tree_add_7_25_groupi_n_6374, csa_tree_add_7_25_groupi_n_6375, csa_tree_add_7_25_groupi_n_6376, csa_tree_add_7_25_groupi_n_6377, csa_tree_add_7_25_groupi_n_6378, csa_tree_add_7_25_groupi_n_6379, csa_tree_add_7_25_groupi_n_6380;
  wire csa_tree_add_7_25_groupi_n_6381, csa_tree_add_7_25_groupi_n_6382, csa_tree_add_7_25_groupi_n_6383, csa_tree_add_7_25_groupi_n_6384, csa_tree_add_7_25_groupi_n_6385, csa_tree_add_7_25_groupi_n_6386, csa_tree_add_7_25_groupi_n_6387, csa_tree_add_7_25_groupi_n_6388;
  wire csa_tree_add_7_25_groupi_n_6389, csa_tree_add_7_25_groupi_n_6390, csa_tree_add_7_25_groupi_n_6391, csa_tree_add_7_25_groupi_n_6392, csa_tree_add_7_25_groupi_n_6393, csa_tree_add_7_25_groupi_n_6394, csa_tree_add_7_25_groupi_n_6395, csa_tree_add_7_25_groupi_n_6396;
  wire csa_tree_add_7_25_groupi_n_6397, csa_tree_add_7_25_groupi_n_6398, csa_tree_add_7_25_groupi_n_6399, csa_tree_add_7_25_groupi_n_6400, csa_tree_add_7_25_groupi_n_6401, csa_tree_add_7_25_groupi_n_6402, csa_tree_add_7_25_groupi_n_6403, csa_tree_add_7_25_groupi_n_6404;
  wire csa_tree_add_7_25_groupi_n_6405, csa_tree_add_7_25_groupi_n_6406, csa_tree_add_7_25_groupi_n_6407, csa_tree_add_7_25_groupi_n_6408, csa_tree_add_7_25_groupi_n_6409, csa_tree_add_7_25_groupi_n_6410, csa_tree_add_7_25_groupi_n_6411, csa_tree_add_7_25_groupi_n_6412;
  wire csa_tree_add_7_25_groupi_n_6413, csa_tree_add_7_25_groupi_n_6414, csa_tree_add_7_25_groupi_n_6416, csa_tree_add_7_25_groupi_n_6417, csa_tree_add_7_25_groupi_n_6418, csa_tree_add_7_25_groupi_n_6419, csa_tree_add_7_25_groupi_n_6420, csa_tree_add_7_25_groupi_n_6421;
  wire csa_tree_add_7_25_groupi_n_6422, csa_tree_add_7_25_groupi_n_6423, csa_tree_add_7_25_groupi_n_6424, csa_tree_add_7_25_groupi_n_6425, csa_tree_add_7_25_groupi_n_6426, csa_tree_add_7_25_groupi_n_6427, csa_tree_add_7_25_groupi_n_6428, csa_tree_add_7_25_groupi_n_6429;
  wire csa_tree_add_7_25_groupi_n_6430, csa_tree_add_7_25_groupi_n_6431, csa_tree_add_7_25_groupi_n_6432, csa_tree_add_7_25_groupi_n_6433, csa_tree_add_7_25_groupi_n_6434, csa_tree_add_7_25_groupi_n_6435, csa_tree_add_7_25_groupi_n_6436, csa_tree_add_7_25_groupi_n_6437;
  wire csa_tree_add_7_25_groupi_n_6438, csa_tree_add_7_25_groupi_n_6439, csa_tree_add_7_25_groupi_n_6440, csa_tree_add_7_25_groupi_n_6441, csa_tree_add_7_25_groupi_n_6442, csa_tree_add_7_25_groupi_n_6443, csa_tree_add_7_25_groupi_n_6444, csa_tree_add_7_25_groupi_n_6445;
  wire csa_tree_add_7_25_groupi_n_6446, csa_tree_add_7_25_groupi_n_6447, csa_tree_add_7_25_groupi_n_6448, csa_tree_add_7_25_groupi_n_6449, csa_tree_add_7_25_groupi_n_6450, csa_tree_add_7_25_groupi_n_6451, csa_tree_add_7_25_groupi_n_6452, csa_tree_add_7_25_groupi_n_6453;
  wire csa_tree_add_7_25_groupi_n_6454, csa_tree_add_7_25_groupi_n_6455, csa_tree_add_7_25_groupi_n_6456, csa_tree_add_7_25_groupi_n_6457, csa_tree_add_7_25_groupi_n_6458, csa_tree_add_7_25_groupi_n_6459, csa_tree_add_7_25_groupi_n_6460, csa_tree_add_7_25_groupi_n_6461;
  wire csa_tree_add_7_25_groupi_n_6462, csa_tree_add_7_25_groupi_n_6463, csa_tree_add_7_25_groupi_n_6464, csa_tree_add_7_25_groupi_n_6465, csa_tree_add_7_25_groupi_n_6466, csa_tree_add_7_25_groupi_n_6467, csa_tree_add_7_25_groupi_n_6468, csa_tree_add_7_25_groupi_n_6469;
  wire csa_tree_add_7_25_groupi_n_6470, csa_tree_add_7_25_groupi_n_6471, csa_tree_add_7_25_groupi_n_6472, csa_tree_add_7_25_groupi_n_6473, csa_tree_add_7_25_groupi_n_6474, csa_tree_add_7_25_groupi_n_6475, csa_tree_add_7_25_groupi_n_6476, csa_tree_add_7_25_groupi_n_6477;
  wire csa_tree_add_7_25_groupi_n_6478, csa_tree_add_7_25_groupi_n_6479, csa_tree_add_7_25_groupi_n_6480, csa_tree_add_7_25_groupi_n_6481, csa_tree_add_7_25_groupi_n_6482, csa_tree_add_7_25_groupi_n_6483, csa_tree_add_7_25_groupi_n_6484, csa_tree_add_7_25_groupi_n_6485;
  wire csa_tree_add_7_25_groupi_n_6486, csa_tree_add_7_25_groupi_n_6487, csa_tree_add_7_25_groupi_n_6488, csa_tree_add_7_25_groupi_n_6489, csa_tree_add_7_25_groupi_n_6490, csa_tree_add_7_25_groupi_n_6492, csa_tree_add_7_25_groupi_n_6493, csa_tree_add_7_25_groupi_n_6494;
  wire csa_tree_add_7_25_groupi_n_6495, csa_tree_add_7_25_groupi_n_6496, csa_tree_add_7_25_groupi_n_6497, csa_tree_add_7_25_groupi_n_6498, csa_tree_add_7_25_groupi_n_6499, csa_tree_add_7_25_groupi_n_6500, csa_tree_add_7_25_groupi_n_6501, csa_tree_add_7_25_groupi_n_6502;
  wire csa_tree_add_7_25_groupi_n_6503, csa_tree_add_7_25_groupi_n_6504, csa_tree_add_7_25_groupi_n_6505, csa_tree_add_7_25_groupi_n_6506, csa_tree_add_7_25_groupi_n_6507, csa_tree_add_7_25_groupi_n_6508, csa_tree_add_7_25_groupi_n_6509, csa_tree_add_7_25_groupi_n_6510;
  wire csa_tree_add_7_25_groupi_n_6511, csa_tree_add_7_25_groupi_n_6512, csa_tree_add_7_25_groupi_n_6513, csa_tree_add_7_25_groupi_n_6514, csa_tree_add_7_25_groupi_n_6515, csa_tree_add_7_25_groupi_n_6516, csa_tree_add_7_25_groupi_n_6517, csa_tree_add_7_25_groupi_n_6518;
  wire csa_tree_add_7_25_groupi_n_6519, csa_tree_add_7_25_groupi_n_6520, csa_tree_add_7_25_groupi_n_6521, csa_tree_add_7_25_groupi_n_6522, csa_tree_add_7_25_groupi_n_6523, csa_tree_add_7_25_groupi_n_6524, csa_tree_add_7_25_groupi_n_6525, csa_tree_add_7_25_groupi_n_6526;
  wire csa_tree_add_7_25_groupi_n_6527, csa_tree_add_7_25_groupi_n_6528, csa_tree_add_7_25_groupi_n_6529, csa_tree_add_7_25_groupi_n_6530, csa_tree_add_7_25_groupi_n_6531, csa_tree_add_7_25_groupi_n_6532, csa_tree_add_7_25_groupi_n_6533, csa_tree_add_7_25_groupi_n_6534;
  wire csa_tree_add_7_25_groupi_n_6535, csa_tree_add_7_25_groupi_n_6536, csa_tree_add_7_25_groupi_n_6537, csa_tree_add_7_25_groupi_n_6538, csa_tree_add_7_25_groupi_n_6539, csa_tree_add_7_25_groupi_n_6540, csa_tree_add_7_25_groupi_n_6541, csa_tree_add_7_25_groupi_n_6542;
  wire csa_tree_add_7_25_groupi_n_6543, csa_tree_add_7_25_groupi_n_6544, csa_tree_add_7_25_groupi_n_6545, csa_tree_add_7_25_groupi_n_6546, csa_tree_add_7_25_groupi_n_6547, csa_tree_add_7_25_groupi_n_6548, csa_tree_add_7_25_groupi_n_6549, csa_tree_add_7_25_groupi_n_6550;
  wire csa_tree_add_7_25_groupi_n_6551, csa_tree_add_7_25_groupi_n_6552, csa_tree_add_7_25_groupi_n_6553, csa_tree_add_7_25_groupi_n_6554, csa_tree_add_7_25_groupi_n_6555, csa_tree_add_7_25_groupi_n_6556, csa_tree_add_7_25_groupi_n_6557, csa_tree_add_7_25_groupi_n_6558;
  wire csa_tree_add_7_25_groupi_n_6559, csa_tree_add_7_25_groupi_n_6560, csa_tree_add_7_25_groupi_n_6561, csa_tree_add_7_25_groupi_n_6562, csa_tree_add_7_25_groupi_n_6563, csa_tree_add_7_25_groupi_n_6564, csa_tree_add_7_25_groupi_n_6565, csa_tree_add_7_25_groupi_n_6566;
  wire csa_tree_add_7_25_groupi_n_6567, csa_tree_add_7_25_groupi_n_6568, csa_tree_add_7_25_groupi_n_6569, csa_tree_add_7_25_groupi_n_6570, csa_tree_add_7_25_groupi_n_6571, csa_tree_add_7_25_groupi_n_6572, csa_tree_add_7_25_groupi_n_6573, csa_tree_add_7_25_groupi_n_6574;
  wire csa_tree_add_7_25_groupi_n_6575, csa_tree_add_7_25_groupi_n_6576, csa_tree_add_7_25_groupi_n_6577, csa_tree_add_7_25_groupi_n_6578, csa_tree_add_7_25_groupi_n_6579, csa_tree_add_7_25_groupi_n_6580, csa_tree_add_7_25_groupi_n_6581, csa_tree_add_7_25_groupi_n_6582;
  wire csa_tree_add_7_25_groupi_n_6583, csa_tree_add_7_25_groupi_n_6584, csa_tree_add_7_25_groupi_n_6585, csa_tree_add_7_25_groupi_n_6587, csa_tree_add_7_25_groupi_n_6588, csa_tree_add_7_25_groupi_n_6589, csa_tree_add_7_25_groupi_n_6590, csa_tree_add_7_25_groupi_n_6591;
  wire csa_tree_add_7_25_groupi_n_6592, csa_tree_add_7_25_groupi_n_6593, csa_tree_add_7_25_groupi_n_6594, csa_tree_add_7_25_groupi_n_6595, csa_tree_add_7_25_groupi_n_6596, csa_tree_add_7_25_groupi_n_6597, csa_tree_add_7_25_groupi_n_6598, csa_tree_add_7_25_groupi_n_6599;
  wire csa_tree_add_7_25_groupi_n_6600, csa_tree_add_7_25_groupi_n_6601, csa_tree_add_7_25_groupi_n_6602, csa_tree_add_7_25_groupi_n_6603, csa_tree_add_7_25_groupi_n_6604, csa_tree_add_7_25_groupi_n_6605, csa_tree_add_7_25_groupi_n_6606, csa_tree_add_7_25_groupi_n_6607;
  wire csa_tree_add_7_25_groupi_n_6608, csa_tree_add_7_25_groupi_n_6609, csa_tree_add_7_25_groupi_n_6610, csa_tree_add_7_25_groupi_n_6611, csa_tree_add_7_25_groupi_n_6612, csa_tree_add_7_25_groupi_n_6613, csa_tree_add_7_25_groupi_n_6614, csa_tree_add_7_25_groupi_n_6615;
  wire csa_tree_add_7_25_groupi_n_6616, csa_tree_add_7_25_groupi_n_6617, csa_tree_add_7_25_groupi_n_6618, csa_tree_add_7_25_groupi_n_6619, csa_tree_add_7_25_groupi_n_6620, csa_tree_add_7_25_groupi_n_6621, csa_tree_add_7_25_groupi_n_6622, csa_tree_add_7_25_groupi_n_6623;
  wire csa_tree_add_7_25_groupi_n_6624, csa_tree_add_7_25_groupi_n_6625, csa_tree_add_7_25_groupi_n_6626, csa_tree_add_7_25_groupi_n_6627, csa_tree_add_7_25_groupi_n_6628, csa_tree_add_7_25_groupi_n_6629, csa_tree_add_7_25_groupi_n_6630, csa_tree_add_7_25_groupi_n_6631;
  wire csa_tree_add_7_25_groupi_n_6632, csa_tree_add_7_25_groupi_n_6633, csa_tree_add_7_25_groupi_n_6634, csa_tree_add_7_25_groupi_n_6635, csa_tree_add_7_25_groupi_n_6636, csa_tree_add_7_25_groupi_n_6637, csa_tree_add_7_25_groupi_n_6638, csa_tree_add_7_25_groupi_n_6639;
  wire csa_tree_add_7_25_groupi_n_6640, csa_tree_add_7_25_groupi_n_6641, csa_tree_add_7_25_groupi_n_6642, csa_tree_add_7_25_groupi_n_6643, csa_tree_add_7_25_groupi_n_6644, csa_tree_add_7_25_groupi_n_6645, csa_tree_add_7_25_groupi_n_6646, csa_tree_add_7_25_groupi_n_6647;
  wire csa_tree_add_7_25_groupi_n_6648, csa_tree_add_7_25_groupi_n_6649, csa_tree_add_7_25_groupi_n_6650, csa_tree_add_7_25_groupi_n_6651, csa_tree_add_7_25_groupi_n_6652, csa_tree_add_7_25_groupi_n_6653, csa_tree_add_7_25_groupi_n_6654, csa_tree_add_7_25_groupi_n_6655;
  wire csa_tree_add_7_25_groupi_n_6656, csa_tree_add_7_25_groupi_n_6657, csa_tree_add_7_25_groupi_n_6658, csa_tree_add_7_25_groupi_n_6659, csa_tree_add_7_25_groupi_n_6660, csa_tree_add_7_25_groupi_n_6661, csa_tree_add_7_25_groupi_n_6662, csa_tree_add_7_25_groupi_n_6663;
  wire csa_tree_add_7_25_groupi_n_6664, csa_tree_add_7_25_groupi_n_6665, csa_tree_add_7_25_groupi_n_6666, csa_tree_add_7_25_groupi_n_6667, csa_tree_add_7_25_groupi_n_6668, csa_tree_add_7_25_groupi_n_6669, csa_tree_add_7_25_groupi_n_6670, csa_tree_add_7_25_groupi_n_6671;
  wire csa_tree_add_7_25_groupi_n_6672, csa_tree_add_7_25_groupi_n_6673, csa_tree_add_7_25_groupi_n_6674, csa_tree_add_7_25_groupi_n_6675, csa_tree_add_7_25_groupi_n_6676, csa_tree_add_7_25_groupi_n_6678, csa_tree_add_7_25_groupi_n_6679, csa_tree_add_7_25_groupi_n_6680;
  wire csa_tree_add_7_25_groupi_n_6681, csa_tree_add_7_25_groupi_n_6682, csa_tree_add_7_25_groupi_n_6683, csa_tree_add_7_25_groupi_n_6684, csa_tree_add_7_25_groupi_n_6685, csa_tree_add_7_25_groupi_n_6686, csa_tree_add_7_25_groupi_n_6687, csa_tree_add_7_25_groupi_n_6688;
  wire csa_tree_add_7_25_groupi_n_6689, csa_tree_add_7_25_groupi_n_6690, csa_tree_add_7_25_groupi_n_6691, csa_tree_add_7_25_groupi_n_6692, csa_tree_add_7_25_groupi_n_6693, csa_tree_add_7_25_groupi_n_6694, csa_tree_add_7_25_groupi_n_6695, csa_tree_add_7_25_groupi_n_6696;
  wire csa_tree_add_7_25_groupi_n_6697, csa_tree_add_7_25_groupi_n_6698, csa_tree_add_7_25_groupi_n_6699, csa_tree_add_7_25_groupi_n_6700, csa_tree_add_7_25_groupi_n_6701, csa_tree_add_7_25_groupi_n_6702, csa_tree_add_7_25_groupi_n_6703, csa_tree_add_7_25_groupi_n_6704;
  wire csa_tree_add_7_25_groupi_n_6705, csa_tree_add_7_25_groupi_n_6706, csa_tree_add_7_25_groupi_n_6707, csa_tree_add_7_25_groupi_n_6708, csa_tree_add_7_25_groupi_n_6709, csa_tree_add_7_25_groupi_n_6710, csa_tree_add_7_25_groupi_n_6711, csa_tree_add_7_25_groupi_n_6712;
  wire csa_tree_add_7_25_groupi_n_6713, csa_tree_add_7_25_groupi_n_6714, csa_tree_add_7_25_groupi_n_6715, csa_tree_add_7_25_groupi_n_6716, csa_tree_add_7_25_groupi_n_6717, csa_tree_add_7_25_groupi_n_6718, csa_tree_add_7_25_groupi_n_6719, csa_tree_add_7_25_groupi_n_6720;
  wire csa_tree_add_7_25_groupi_n_6721, csa_tree_add_7_25_groupi_n_6722, csa_tree_add_7_25_groupi_n_6723, csa_tree_add_7_25_groupi_n_6724, csa_tree_add_7_25_groupi_n_6725, csa_tree_add_7_25_groupi_n_6726, csa_tree_add_7_25_groupi_n_6727, csa_tree_add_7_25_groupi_n_6728;
  wire csa_tree_add_7_25_groupi_n_6729, csa_tree_add_7_25_groupi_n_6730, csa_tree_add_7_25_groupi_n_6731, csa_tree_add_7_25_groupi_n_6732, csa_tree_add_7_25_groupi_n_6733, csa_tree_add_7_25_groupi_n_6734, csa_tree_add_7_25_groupi_n_6735, csa_tree_add_7_25_groupi_n_6736;
  wire csa_tree_add_7_25_groupi_n_6737, csa_tree_add_7_25_groupi_n_6738, csa_tree_add_7_25_groupi_n_6739, csa_tree_add_7_25_groupi_n_6740, csa_tree_add_7_25_groupi_n_6741, csa_tree_add_7_25_groupi_n_6742, csa_tree_add_7_25_groupi_n_6744, csa_tree_add_7_25_groupi_n_6745;
  wire csa_tree_add_7_25_groupi_n_6746, csa_tree_add_7_25_groupi_n_6747, csa_tree_add_7_25_groupi_n_6748, csa_tree_add_7_25_groupi_n_6749, csa_tree_add_7_25_groupi_n_6750, csa_tree_add_7_25_groupi_n_6751, csa_tree_add_7_25_groupi_n_6752, csa_tree_add_7_25_groupi_n_6753;
  wire csa_tree_add_7_25_groupi_n_6754, csa_tree_add_7_25_groupi_n_6755, csa_tree_add_7_25_groupi_n_6756, csa_tree_add_7_25_groupi_n_6757, csa_tree_add_7_25_groupi_n_6758, csa_tree_add_7_25_groupi_n_6759, csa_tree_add_7_25_groupi_n_6760, csa_tree_add_7_25_groupi_n_6761;
  wire csa_tree_add_7_25_groupi_n_6762, csa_tree_add_7_25_groupi_n_6763, csa_tree_add_7_25_groupi_n_6764, csa_tree_add_7_25_groupi_n_6765, csa_tree_add_7_25_groupi_n_6766, csa_tree_add_7_25_groupi_n_6767, csa_tree_add_7_25_groupi_n_6768, csa_tree_add_7_25_groupi_n_6769;
  wire csa_tree_add_7_25_groupi_n_6770, csa_tree_add_7_25_groupi_n_6771, csa_tree_add_7_25_groupi_n_6772, csa_tree_add_7_25_groupi_n_6773, csa_tree_add_7_25_groupi_n_6774, csa_tree_add_7_25_groupi_n_6775, csa_tree_add_7_25_groupi_n_6776, csa_tree_add_7_25_groupi_n_6777;
  wire csa_tree_add_7_25_groupi_n_6778, csa_tree_add_7_25_groupi_n_6779, csa_tree_add_7_25_groupi_n_6780, csa_tree_add_7_25_groupi_n_6781, csa_tree_add_7_25_groupi_n_6782, csa_tree_add_7_25_groupi_n_6783, csa_tree_add_7_25_groupi_n_6784, csa_tree_add_7_25_groupi_n_6785;
  wire csa_tree_add_7_25_groupi_n_6786, csa_tree_add_7_25_groupi_n_6787, csa_tree_add_7_25_groupi_n_6788, csa_tree_add_7_25_groupi_n_6789, csa_tree_add_7_25_groupi_n_6790, csa_tree_add_7_25_groupi_n_6791, csa_tree_add_7_25_groupi_n_6792, csa_tree_add_7_25_groupi_n_6793;
  wire csa_tree_add_7_25_groupi_n_6794, csa_tree_add_7_25_groupi_n_6795, csa_tree_add_7_25_groupi_n_6796, csa_tree_add_7_25_groupi_n_6797, csa_tree_add_7_25_groupi_n_6798, csa_tree_add_7_25_groupi_n_6799, csa_tree_add_7_25_groupi_n_6800, csa_tree_add_7_25_groupi_n_6801;
  wire csa_tree_add_7_25_groupi_n_6802, csa_tree_add_7_25_groupi_n_6803, csa_tree_add_7_25_groupi_n_6804, csa_tree_add_7_25_groupi_n_6805, csa_tree_add_7_25_groupi_n_6806, csa_tree_add_7_25_groupi_n_6807, csa_tree_add_7_25_groupi_n_6808, csa_tree_add_7_25_groupi_n_6809;
  wire csa_tree_add_7_25_groupi_n_6810, csa_tree_add_7_25_groupi_n_6811, csa_tree_add_7_25_groupi_n_6812, csa_tree_add_7_25_groupi_n_6813, csa_tree_add_7_25_groupi_n_6814, csa_tree_add_7_25_groupi_n_6815, csa_tree_add_7_25_groupi_n_6816, csa_tree_add_7_25_groupi_n_6817;
  wire csa_tree_add_7_25_groupi_n_6818, csa_tree_add_7_25_groupi_n_6819, csa_tree_add_7_25_groupi_n_6820, csa_tree_add_7_25_groupi_n_6821, csa_tree_add_7_25_groupi_n_6822, csa_tree_add_7_25_groupi_n_6823, csa_tree_add_7_25_groupi_n_6824, csa_tree_add_7_25_groupi_n_6825;
  wire csa_tree_add_7_25_groupi_n_6826, csa_tree_add_7_25_groupi_n_6827, csa_tree_add_7_25_groupi_n_6828, csa_tree_add_7_25_groupi_n_6830, csa_tree_add_7_25_groupi_n_6831, csa_tree_add_7_25_groupi_n_6832, csa_tree_add_7_25_groupi_n_6833, csa_tree_add_7_25_groupi_n_6834;
  wire csa_tree_add_7_25_groupi_n_6835, csa_tree_add_7_25_groupi_n_6836, csa_tree_add_7_25_groupi_n_6837, csa_tree_add_7_25_groupi_n_6838, csa_tree_add_7_25_groupi_n_6839, csa_tree_add_7_25_groupi_n_6840, csa_tree_add_7_25_groupi_n_6841, csa_tree_add_7_25_groupi_n_6842;
  wire csa_tree_add_7_25_groupi_n_6843, csa_tree_add_7_25_groupi_n_6844, csa_tree_add_7_25_groupi_n_6845, csa_tree_add_7_25_groupi_n_6846, csa_tree_add_7_25_groupi_n_6847, csa_tree_add_7_25_groupi_n_6848, csa_tree_add_7_25_groupi_n_6849, csa_tree_add_7_25_groupi_n_6850;
  wire csa_tree_add_7_25_groupi_n_6851, csa_tree_add_7_25_groupi_n_6852, csa_tree_add_7_25_groupi_n_6853, csa_tree_add_7_25_groupi_n_6854, csa_tree_add_7_25_groupi_n_6855, csa_tree_add_7_25_groupi_n_6856, csa_tree_add_7_25_groupi_n_6857, csa_tree_add_7_25_groupi_n_6858;
  wire csa_tree_add_7_25_groupi_n_6859, csa_tree_add_7_25_groupi_n_6860, csa_tree_add_7_25_groupi_n_6861, csa_tree_add_7_25_groupi_n_6862, csa_tree_add_7_25_groupi_n_6863, csa_tree_add_7_25_groupi_n_6864, csa_tree_add_7_25_groupi_n_6865, csa_tree_add_7_25_groupi_n_6866;
  wire csa_tree_add_7_25_groupi_n_6867, csa_tree_add_7_25_groupi_n_6868, csa_tree_add_7_25_groupi_n_6869, csa_tree_add_7_25_groupi_n_6870, csa_tree_add_7_25_groupi_n_6871, csa_tree_add_7_25_groupi_n_6872, csa_tree_add_7_25_groupi_n_6873, csa_tree_add_7_25_groupi_n_6874;
  wire csa_tree_add_7_25_groupi_n_6875, csa_tree_add_7_25_groupi_n_6876, csa_tree_add_7_25_groupi_n_6877, csa_tree_add_7_25_groupi_n_6878, csa_tree_add_7_25_groupi_n_6879, csa_tree_add_7_25_groupi_n_6880, csa_tree_add_7_25_groupi_n_6881, csa_tree_add_7_25_groupi_n_6882;
  wire csa_tree_add_7_25_groupi_n_6883, csa_tree_add_7_25_groupi_n_6884, csa_tree_add_7_25_groupi_n_6885, csa_tree_add_7_25_groupi_n_6886, csa_tree_add_7_25_groupi_n_6887, csa_tree_add_7_25_groupi_n_6888, csa_tree_add_7_25_groupi_n_6889, csa_tree_add_7_25_groupi_n_6890;
  wire csa_tree_add_7_25_groupi_n_6891, csa_tree_add_7_25_groupi_n_6892, csa_tree_add_7_25_groupi_n_6893, csa_tree_add_7_25_groupi_n_6894, csa_tree_add_7_25_groupi_n_6895, csa_tree_add_7_25_groupi_n_6896, csa_tree_add_7_25_groupi_n_6897, csa_tree_add_7_25_groupi_n_6898;
  wire csa_tree_add_7_25_groupi_n_6899, csa_tree_add_7_25_groupi_n_6900, csa_tree_add_7_25_groupi_n_6901, csa_tree_add_7_25_groupi_n_6902, csa_tree_add_7_25_groupi_n_6903, csa_tree_add_7_25_groupi_n_6904, csa_tree_add_7_25_groupi_n_6905, csa_tree_add_7_25_groupi_n_6906;
  wire csa_tree_add_7_25_groupi_n_6907, csa_tree_add_7_25_groupi_n_6908, csa_tree_add_7_25_groupi_n_6909, csa_tree_add_7_25_groupi_n_6910, csa_tree_add_7_25_groupi_n_6911, csa_tree_add_7_25_groupi_n_6913, csa_tree_add_7_25_groupi_n_6914, csa_tree_add_7_25_groupi_n_6915;
  wire csa_tree_add_7_25_groupi_n_6916, csa_tree_add_7_25_groupi_n_6917, csa_tree_add_7_25_groupi_n_6918, csa_tree_add_7_25_groupi_n_6919, csa_tree_add_7_25_groupi_n_6920, csa_tree_add_7_25_groupi_n_6921, csa_tree_add_7_25_groupi_n_6922, csa_tree_add_7_25_groupi_n_6923;
  wire csa_tree_add_7_25_groupi_n_6924, csa_tree_add_7_25_groupi_n_6925, csa_tree_add_7_25_groupi_n_6926, csa_tree_add_7_25_groupi_n_6927, csa_tree_add_7_25_groupi_n_6928, csa_tree_add_7_25_groupi_n_6929, csa_tree_add_7_25_groupi_n_6930, csa_tree_add_7_25_groupi_n_6931;
  wire csa_tree_add_7_25_groupi_n_6932, csa_tree_add_7_25_groupi_n_6933, csa_tree_add_7_25_groupi_n_6934, csa_tree_add_7_25_groupi_n_6935, csa_tree_add_7_25_groupi_n_6936, csa_tree_add_7_25_groupi_n_6937, csa_tree_add_7_25_groupi_n_6938, csa_tree_add_7_25_groupi_n_6939;
  wire csa_tree_add_7_25_groupi_n_6940, csa_tree_add_7_25_groupi_n_6941, csa_tree_add_7_25_groupi_n_6942, csa_tree_add_7_25_groupi_n_6943, csa_tree_add_7_25_groupi_n_6944, csa_tree_add_7_25_groupi_n_6945, csa_tree_add_7_25_groupi_n_6946, csa_tree_add_7_25_groupi_n_6947;
  wire csa_tree_add_7_25_groupi_n_6948, csa_tree_add_7_25_groupi_n_6949, csa_tree_add_7_25_groupi_n_6950, csa_tree_add_7_25_groupi_n_6951, csa_tree_add_7_25_groupi_n_6952, csa_tree_add_7_25_groupi_n_6953, csa_tree_add_7_25_groupi_n_6954, csa_tree_add_7_25_groupi_n_6955;
  wire csa_tree_add_7_25_groupi_n_6956, csa_tree_add_7_25_groupi_n_6957, csa_tree_add_7_25_groupi_n_6958, csa_tree_add_7_25_groupi_n_6959, csa_tree_add_7_25_groupi_n_6960, csa_tree_add_7_25_groupi_n_6961, csa_tree_add_7_25_groupi_n_6962, csa_tree_add_7_25_groupi_n_6963;
  wire csa_tree_add_7_25_groupi_n_6964, csa_tree_add_7_25_groupi_n_6965, csa_tree_add_7_25_groupi_n_6966, csa_tree_add_7_25_groupi_n_6967, csa_tree_add_7_25_groupi_n_6968, csa_tree_add_7_25_groupi_n_6969, csa_tree_add_7_25_groupi_n_6970, csa_tree_add_7_25_groupi_n_6971;
  wire csa_tree_add_7_25_groupi_n_6972, csa_tree_add_7_25_groupi_n_6973, csa_tree_add_7_25_groupi_n_6975, csa_tree_add_7_25_groupi_n_6976, csa_tree_add_7_25_groupi_n_6977, csa_tree_add_7_25_groupi_n_6978, csa_tree_add_7_25_groupi_n_6979, csa_tree_add_7_25_groupi_n_6980;
  wire csa_tree_add_7_25_groupi_n_6981, csa_tree_add_7_25_groupi_n_6982, csa_tree_add_7_25_groupi_n_6983, csa_tree_add_7_25_groupi_n_6984, csa_tree_add_7_25_groupi_n_6985, csa_tree_add_7_25_groupi_n_6986, csa_tree_add_7_25_groupi_n_6987, csa_tree_add_7_25_groupi_n_6988;
  wire csa_tree_add_7_25_groupi_n_6989, csa_tree_add_7_25_groupi_n_6990, csa_tree_add_7_25_groupi_n_6991, csa_tree_add_7_25_groupi_n_6992, csa_tree_add_7_25_groupi_n_6993, csa_tree_add_7_25_groupi_n_6994, csa_tree_add_7_25_groupi_n_6995, csa_tree_add_7_25_groupi_n_6996;
  wire csa_tree_add_7_25_groupi_n_6997, csa_tree_add_7_25_groupi_n_6998, csa_tree_add_7_25_groupi_n_6999, csa_tree_add_7_25_groupi_n_7000, csa_tree_add_7_25_groupi_n_7001, csa_tree_add_7_25_groupi_n_7002, csa_tree_add_7_25_groupi_n_7003, csa_tree_add_7_25_groupi_n_7004;
  wire csa_tree_add_7_25_groupi_n_7005, csa_tree_add_7_25_groupi_n_7006, csa_tree_add_7_25_groupi_n_7007, csa_tree_add_7_25_groupi_n_7008, csa_tree_add_7_25_groupi_n_7009, csa_tree_add_7_25_groupi_n_7010, csa_tree_add_7_25_groupi_n_7011, csa_tree_add_7_25_groupi_n_7012;
  wire csa_tree_add_7_25_groupi_n_7013, csa_tree_add_7_25_groupi_n_7014, csa_tree_add_7_25_groupi_n_7015, csa_tree_add_7_25_groupi_n_7016, csa_tree_add_7_25_groupi_n_7017, csa_tree_add_7_25_groupi_n_7018, csa_tree_add_7_25_groupi_n_7019, csa_tree_add_7_25_groupi_n_7020;
  wire csa_tree_add_7_25_groupi_n_7021, csa_tree_add_7_25_groupi_n_7022, csa_tree_add_7_25_groupi_n_7023, csa_tree_add_7_25_groupi_n_7024, csa_tree_add_7_25_groupi_n_7025, csa_tree_add_7_25_groupi_n_7026, csa_tree_add_7_25_groupi_n_7027, csa_tree_add_7_25_groupi_n_7028;
  wire csa_tree_add_7_25_groupi_n_7029, csa_tree_add_7_25_groupi_n_7030, csa_tree_add_7_25_groupi_n_7031, csa_tree_add_7_25_groupi_n_7032, csa_tree_add_7_25_groupi_n_7033, csa_tree_add_7_25_groupi_n_7034, csa_tree_add_7_25_groupi_n_7035, csa_tree_add_7_25_groupi_n_7036;
  wire csa_tree_add_7_25_groupi_n_7037, csa_tree_add_7_25_groupi_n_7038, csa_tree_add_7_25_groupi_n_7039, csa_tree_add_7_25_groupi_n_7040, csa_tree_add_7_25_groupi_n_7041, csa_tree_add_7_25_groupi_n_7042, csa_tree_add_7_25_groupi_n_7043, csa_tree_add_7_25_groupi_n_7044;
  wire csa_tree_add_7_25_groupi_n_7045, csa_tree_add_7_25_groupi_n_7046, csa_tree_add_7_25_groupi_n_7047, csa_tree_add_7_25_groupi_n_7048, csa_tree_add_7_25_groupi_n_7050, csa_tree_add_7_25_groupi_n_7051, csa_tree_add_7_25_groupi_n_7052, csa_tree_add_7_25_groupi_n_7053;
  wire csa_tree_add_7_25_groupi_n_7054, csa_tree_add_7_25_groupi_n_7055, csa_tree_add_7_25_groupi_n_7056, csa_tree_add_7_25_groupi_n_7057, csa_tree_add_7_25_groupi_n_7058, csa_tree_add_7_25_groupi_n_7059, csa_tree_add_7_25_groupi_n_7060, csa_tree_add_7_25_groupi_n_7061;
  wire csa_tree_add_7_25_groupi_n_7062, csa_tree_add_7_25_groupi_n_7063, csa_tree_add_7_25_groupi_n_7064, csa_tree_add_7_25_groupi_n_7065, csa_tree_add_7_25_groupi_n_7066, csa_tree_add_7_25_groupi_n_7067, csa_tree_add_7_25_groupi_n_7068, csa_tree_add_7_25_groupi_n_7069;
  wire csa_tree_add_7_25_groupi_n_7070, csa_tree_add_7_25_groupi_n_7071, csa_tree_add_7_25_groupi_n_7072, csa_tree_add_7_25_groupi_n_7073, csa_tree_add_7_25_groupi_n_7074, csa_tree_add_7_25_groupi_n_7075, csa_tree_add_7_25_groupi_n_7076, csa_tree_add_7_25_groupi_n_7077;
  wire csa_tree_add_7_25_groupi_n_7078, csa_tree_add_7_25_groupi_n_7079, csa_tree_add_7_25_groupi_n_7080, csa_tree_add_7_25_groupi_n_7081, csa_tree_add_7_25_groupi_n_7082, csa_tree_add_7_25_groupi_n_7083, csa_tree_add_7_25_groupi_n_7084, csa_tree_add_7_25_groupi_n_7085;
  wire csa_tree_add_7_25_groupi_n_7086, csa_tree_add_7_25_groupi_n_7087, csa_tree_add_7_25_groupi_n_7088, csa_tree_add_7_25_groupi_n_7089, csa_tree_add_7_25_groupi_n_7090, csa_tree_add_7_25_groupi_n_7091, csa_tree_add_7_25_groupi_n_7092, csa_tree_add_7_25_groupi_n_7093;
  wire csa_tree_add_7_25_groupi_n_7094, csa_tree_add_7_25_groupi_n_7095, csa_tree_add_7_25_groupi_n_7096, csa_tree_add_7_25_groupi_n_7097, csa_tree_add_7_25_groupi_n_7098, csa_tree_add_7_25_groupi_n_7099, csa_tree_add_7_25_groupi_n_7100, csa_tree_add_7_25_groupi_n_7101;
  wire csa_tree_add_7_25_groupi_n_7102, csa_tree_add_7_25_groupi_n_7103, csa_tree_add_7_25_groupi_n_7104, csa_tree_add_7_25_groupi_n_7105, csa_tree_add_7_25_groupi_n_7106, csa_tree_add_7_25_groupi_n_7107, csa_tree_add_7_25_groupi_n_7108, csa_tree_add_7_25_groupi_n_7109;
  wire csa_tree_add_7_25_groupi_n_7110, csa_tree_add_7_25_groupi_n_7111, csa_tree_add_7_25_groupi_n_7112, csa_tree_add_7_25_groupi_n_7113, csa_tree_add_7_25_groupi_n_7114, csa_tree_add_7_25_groupi_n_7116, csa_tree_add_7_25_groupi_n_7117, csa_tree_add_7_25_groupi_n_7118;
  wire csa_tree_add_7_25_groupi_n_7119, csa_tree_add_7_25_groupi_n_7120, csa_tree_add_7_25_groupi_n_7121, csa_tree_add_7_25_groupi_n_7122, csa_tree_add_7_25_groupi_n_7123, csa_tree_add_7_25_groupi_n_7124, csa_tree_add_7_25_groupi_n_7125, csa_tree_add_7_25_groupi_n_7126;
  wire csa_tree_add_7_25_groupi_n_7127, csa_tree_add_7_25_groupi_n_7128, csa_tree_add_7_25_groupi_n_7129, csa_tree_add_7_25_groupi_n_7130, csa_tree_add_7_25_groupi_n_7131, csa_tree_add_7_25_groupi_n_7132, csa_tree_add_7_25_groupi_n_7133, csa_tree_add_7_25_groupi_n_7134;
  wire csa_tree_add_7_25_groupi_n_7135, csa_tree_add_7_25_groupi_n_7136, csa_tree_add_7_25_groupi_n_7137, csa_tree_add_7_25_groupi_n_7138, csa_tree_add_7_25_groupi_n_7139, csa_tree_add_7_25_groupi_n_7140, csa_tree_add_7_25_groupi_n_7141, csa_tree_add_7_25_groupi_n_7142;
  wire csa_tree_add_7_25_groupi_n_7143, csa_tree_add_7_25_groupi_n_7144, csa_tree_add_7_25_groupi_n_7145, csa_tree_add_7_25_groupi_n_7146, csa_tree_add_7_25_groupi_n_7147, csa_tree_add_7_25_groupi_n_7148, csa_tree_add_7_25_groupi_n_7149, csa_tree_add_7_25_groupi_n_7150;
  wire csa_tree_add_7_25_groupi_n_7151, csa_tree_add_7_25_groupi_n_7152, csa_tree_add_7_25_groupi_n_7153, csa_tree_add_7_25_groupi_n_7154, csa_tree_add_7_25_groupi_n_7155, csa_tree_add_7_25_groupi_n_7156, csa_tree_add_7_25_groupi_n_7157, csa_tree_add_7_25_groupi_n_7158;
  wire csa_tree_add_7_25_groupi_n_7159, csa_tree_add_7_25_groupi_n_7160, csa_tree_add_7_25_groupi_n_7162, csa_tree_add_7_25_groupi_n_7163, csa_tree_add_7_25_groupi_n_7164, csa_tree_add_7_25_groupi_n_7165, csa_tree_add_7_25_groupi_n_7166, csa_tree_add_7_25_groupi_n_7167;
  wire csa_tree_add_7_25_groupi_n_7168, csa_tree_add_7_25_groupi_n_7169, csa_tree_add_7_25_groupi_n_7170, csa_tree_add_7_25_groupi_n_7171, csa_tree_add_7_25_groupi_n_7172, csa_tree_add_7_25_groupi_n_7173, csa_tree_add_7_25_groupi_n_7174, csa_tree_add_7_25_groupi_n_7175;
  wire csa_tree_add_7_25_groupi_n_7176, csa_tree_add_7_25_groupi_n_7177, csa_tree_add_7_25_groupi_n_7178, csa_tree_add_7_25_groupi_n_7179, csa_tree_add_7_25_groupi_n_7180, csa_tree_add_7_25_groupi_n_7181, csa_tree_add_7_25_groupi_n_7182, csa_tree_add_7_25_groupi_n_7183;
  wire csa_tree_add_7_25_groupi_n_7184, csa_tree_add_7_25_groupi_n_7185, csa_tree_add_7_25_groupi_n_7186, csa_tree_add_7_25_groupi_n_7187, csa_tree_add_7_25_groupi_n_7188, csa_tree_add_7_25_groupi_n_7189, csa_tree_add_7_25_groupi_n_7190, csa_tree_add_7_25_groupi_n_7191;
  wire csa_tree_add_7_25_groupi_n_7192, csa_tree_add_7_25_groupi_n_7193, csa_tree_add_7_25_groupi_n_7194, csa_tree_add_7_25_groupi_n_7195, csa_tree_add_7_25_groupi_n_7196, csa_tree_add_7_25_groupi_n_7197, csa_tree_add_7_25_groupi_n_7198, csa_tree_add_7_25_groupi_n_7199;
  wire csa_tree_add_7_25_groupi_n_7200, csa_tree_add_7_25_groupi_n_7201, csa_tree_add_7_25_groupi_n_7202, csa_tree_add_7_25_groupi_n_7203, csa_tree_add_7_25_groupi_n_7204, csa_tree_add_7_25_groupi_n_7205, csa_tree_add_7_25_groupi_n_7206, csa_tree_add_7_25_groupi_n_7207;
  wire csa_tree_add_7_25_groupi_n_7208, csa_tree_add_7_25_groupi_n_7209, csa_tree_add_7_25_groupi_n_7210, csa_tree_add_7_25_groupi_n_7211, csa_tree_add_7_25_groupi_n_7212, csa_tree_add_7_25_groupi_n_7213, csa_tree_add_7_25_groupi_n_7214, csa_tree_add_7_25_groupi_n_7217;
  wire csa_tree_add_7_25_groupi_n_7218, csa_tree_add_7_25_groupi_n_7220, csa_tree_add_7_25_groupi_n_7221, csa_tree_add_7_25_groupi_n_7223, csa_tree_add_7_25_groupi_n_7224, csa_tree_add_7_25_groupi_n_7226, csa_tree_add_7_25_groupi_n_7227, csa_tree_add_7_25_groupi_n_7229;
  wire csa_tree_add_7_25_groupi_n_7230, csa_tree_add_7_25_groupi_n_7231, csa_tree_add_7_25_groupi_n_7233, csa_tree_add_7_25_groupi_n_7234, csa_tree_add_7_25_groupi_n_7236, csa_tree_add_7_25_groupi_n_7237, csa_tree_add_7_25_groupi_n_7238, csa_tree_add_7_25_groupi_n_7239;
  wire csa_tree_add_7_25_groupi_n_7240, csa_tree_add_7_25_groupi_n_7241, csa_tree_add_7_25_groupi_n_7243, csa_tree_add_7_25_groupi_n_7244, csa_tree_add_7_25_groupi_n_7245, csa_tree_add_7_25_groupi_n_7246, csa_tree_add_7_25_groupi_n_7247, csa_tree_add_7_25_groupi_n_7248;
  wire csa_tree_add_7_25_groupi_n_7250;
  xnor csa_tree_add_7_25_groupi_g13828__2398(out2[40] ,csa_tree_add_7_25_groupi_n_7250 ,csa_tree_add_7_25_groupi_n_7207);
  or csa_tree_add_7_25_groupi_g13829__5107(csa_tree_add_7_25_groupi_n_7250 ,csa_tree_add_7_25_groupi_n_7248 ,csa_tree_add_7_25_groupi_n_7176);
  xnor csa_tree_add_7_25_groupi_g13830__6260(out2[39] ,csa_tree_add_7_25_groupi_n_7247 ,csa_tree_add_7_25_groupi_n_7187);
  nor csa_tree_add_7_25_groupi_g13831__4319(csa_tree_add_7_25_groupi_n_7248 ,csa_tree_add_7_25_groupi_n_7247 ,csa_tree_add_7_25_groupi_n_7182);
  and csa_tree_add_7_25_groupi_g13832__8428(csa_tree_add_7_25_groupi_n_7247 ,csa_tree_add_7_25_groupi_n_7200 ,csa_tree_add_7_25_groupi_n_7246);
  or csa_tree_add_7_25_groupi_g13834__5526(csa_tree_add_7_25_groupi_n_7246 ,csa_tree_add_7_25_groupi_n_7245 ,csa_tree_add_7_25_groupi_n_7195);
  and csa_tree_add_7_25_groupi_g13836__6783(csa_tree_add_7_25_groupi_n_7245 ,csa_tree_add_7_25_groupi_n_7194 ,csa_tree_add_7_25_groupi_n_7244);
  or csa_tree_add_7_25_groupi_g13838__3680(csa_tree_add_7_25_groupi_n_7244 ,csa_tree_add_7_25_groupi_n_7243 ,csa_tree_add_7_25_groupi_n_7196);
  and csa_tree_add_7_25_groupi_g13840__1617(csa_tree_add_7_25_groupi_n_7243 ,csa_tree_add_7_25_groupi_n_7241 ,csa_tree_add_7_25_groupi_n_7172);
  xnor csa_tree_add_7_25_groupi_g13841__2802(out2[36] ,csa_tree_add_7_25_groupi_n_7240 ,csa_tree_add_7_25_groupi_n_7186);
  or csa_tree_add_7_25_groupi_g13842__1705(csa_tree_add_7_25_groupi_n_7241 ,csa_tree_add_7_25_groupi_n_7240 ,csa_tree_add_7_25_groupi_n_7173);
  and csa_tree_add_7_25_groupi_g13843__5122(csa_tree_add_7_25_groupi_n_7240 ,csa_tree_add_7_25_groupi_n_7239 ,csa_tree_add_7_25_groupi_n_7197);
  or csa_tree_add_7_25_groupi_g13845__8246(csa_tree_add_7_25_groupi_n_7239 ,csa_tree_add_7_25_groupi_n_7238 ,csa_tree_add_7_25_groupi_n_7198);
  and csa_tree_add_7_25_groupi_g13847__7098(csa_tree_add_7_25_groupi_n_7238 ,csa_tree_add_7_25_groupi_n_7191 ,csa_tree_add_7_25_groupi_n_7237);
  or csa_tree_add_7_25_groupi_g13849__6131(csa_tree_add_7_25_groupi_n_7237 ,csa_tree_add_7_25_groupi_n_7204 ,csa_tree_add_7_25_groupi_n_7236);
  and csa_tree_add_7_25_groupi_g13851__1881(csa_tree_add_7_25_groupi_n_7236 ,csa_tree_add_7_25_groupi_n_7175 ,csa_tree_add_7_25_groupi_n_7234);
  xnor csa_tree_add_7_25_groupi_g13852__5115(out2[33] ,csa_tree_add_7_25_groupi_n_7233 ,csa_tree_add_7_25_groupi_n_7185);
  or csa_tree_add_7_25_groupi_g13853__7482(csa_tree_add_7_25_groupi_n_7234 ,csa_tree_add_7_25_groupi_n_7233 ,csa_tree_add_7_25_groupi_n_7174);
  and csa_tree_add_7_25_groupi_g13854__4733(csa_tree_add_7_25_groupi_n_7233 ,csa_tree_add_7_25_groupi_n_7231 ,csa_tree_add_7_25_groupi_n_7202);
  xnor csa_tree_add_7_25_groupi_g13855__6161(out2[32] ,csa_tree_add_7_25_groupi_n_7229 ,csa_tree_add_7_25_groupi_n_7206);
  or csa_tree_add_7_25_groupi_g13856__9315(csa_tree_add_7_25_groupi_n_7231 ,csa_tree_add_7_25_groupi_n_7230 ,csa_tree_add_7_25_groupi_n_7203);
  not csa_tree_add_7_25_groupi_g13857(csa_tree_add_7_25_groupi_n_7230 ,csa_tree_add_7_25_groupi_n_7229);
  or csa_tree_add_7_25_groupi_g13858__9945(csa_tree_add_7_25_groupi_n_7229 ,csa_tree_add_7_25_groupi_n_7227 ,csa_tree_add_7_25_groupi_n_7201);
  xnor csa_tree_add_7_25_groupi_g13859__2883(out2[31] ,csa_tree_add_7_25_groupi_n_7226 ,csa_tree_add_7_25_groupi_n_7205);
  and csa_tree_add_7_25_groupi_g13860__2346(csa_tree_add_7_25_groupi_n_7227 ,csa_tree_add_7_25_groupi_n_7199 ,csa_tree_add_7_25_groupi_n_7226);
  or csa_tree_add_7_25_groupi_g13861__1666(csa_tree_add_7_25_groupi_n_7226 ,csa_tree_add_7_25_groupi_n_7224 ,csa_tree_add_7_25_groupi_n_7181);
  xnor csa_tree_add_7_25_groupi_g13862__7410(out2[30] ,csa_tree_add_7_25_groupi_n_7223 ,csa_tree_add_7_25_groupi_n_7183);
  and csa_tree_add_7_25_groupi_g13863__6417(csa_tree_add_7_25_groupi_n_7224 ,csa_tree_add_7_25_groupi_n_7177 ,csa_tree_add_7_25_groupi_n_7223);
  or csa_tree_add_7_25_groupi_g13864__5477(csa_tree_add_7_25_groupi_n_7223 ,csa_tree_add_7_25_groupi_n_7188 ,csa_tree_add_7_25_groupi_n_7221);
  xnor csa_tree_add_7_25_groupi_g13865__2398(out2[29] ,csa_tree_add_7_25_groupi_n_7220 ,csa_tree_add_7_25_groupi_n_7213);
  and csa_tree_add_7_25_groupi_g13866__5107(csa_tree_add_7_25_groupi_n_7221 ,csa_tree_add_7_25_groupi_n_7220 ,csa_tree_add_7_25_groupi_n_7192);
  or csa_tree_add_7_25_groupi_g13867__6260(csa_tree_add_7_25_groupi_n_7220 ,csa_tree_add_7_25_groupi_n_7190 ,csa_tree_add_7_25_groupi_n_7218);
  xnor csa_tree_add_7_25_groupi_g13868__4319(out2[28] ,csa_tree_add_7_25_groupi_n_7217 ,csa_tree_add_7_25_groupi_n_7211);
  and csa_tree_add_7_25_groupi_g13869__8428(csa_tree_add_7_25_groupi_n_7218 ,csa_tree_add_7_25_groupi_n_7189 ,csa_tree_add_7_25_groupi_n_7217);
  or csa_tree_add_7_25_groupi_g13870__5526(csa_tree_add_7_25_groupi_n_7217 ,csa_tree_add_7_25_groupi_n_7214 ,csa_tree_add_7_25_groupi_n_7178);
  xnor csa_tree_add_7_25_groupi_g13871__6783(out2[27] ,csa_tree_add_7_25_groupi_n_7193 ,csa_tree_add_7_25_groupi_n_7184);
  xnor csa_tree_add_7_25_groupi_g13872__3680(out2[26] ,csa_tree_add_7_25_groupi_n_7158 ,csa_tree_add_7_25_groupi_n_7159);
  and csa_tree_add_7_25_groupi_g13873__1617(csa_tree_add_7_25_groupi_n_7214 ,csa_tree_add_7_25_groupi_n_7193 ,csa_tree_add_7_25_groupi_n_7179);
  xnor csa_tree_add_7_25_groupi_g13874__2802(csa_tree_add_7_25_groupi_n_7213 ,csa_tree_add_7_25_groupi_n_7169 ,csa_tree_add_7_25_groupi_n_7146);
  xnor csa_tree_add_7_25_groupi_g13875__1705(csa_tree_add_7_25_groupi_n_7212 ,csa_tree_add_7_25_groupi_n_7162 ,csa_tree_add_7_25_groupi_n_7141);
  xnor csa_tree_add_7_25_groupi_g13876__5122(csa_tree_add_7_25_groupi_n_7211 ,csa_tree_add_7_25_groupi_n_7154 ,csa_tree_add_7_25_groupi_n_7165);
  xnor csa_tree_add_7_25_groupi_g13877__8246(csa_tree_add_7_25_groupi_n_7210 ,csa_tree_add_7_25_groupi_n_7171 ,csa_tree_add_7_25_groupi_n_7145);
  xnor csa_tree_add_7_25_groupi_g13878__7098(csa_tree_add_7_25_groupi_n_7209 ,csa_tree_add_7_25_groupi_n_7140 ,csa_tree_add_7_25_groupi_n_7163);
  xnor csa_tree_add_7_25_groupi_g13879__6131(csa_tree_add_7_25_groupi_n_7208 ,csa_tree_add_7_25_groupi_n_7143 ,csa_tree_add_7_25_groupi_n_7167);
  xnor csa_tree_add_7_25_groupi_g13880__1881(csa_tree_add_7_25_groupi_n_7207 ,csa_tree_add_7_25_groupi_n_7147 ,csa_tree_add_7_25_groupi_n_7160);
  xnor csa_tree_add_7_25_groupi_g13881__5115(csa_tree_add_7_25_groupi_n_7206 ,csa_tree_add_7_25_groupi_n_7164 ,csa_tree_add_7_25_groupi_n_7150);
  xnor csa_tree_add_7_25_groupi_g13882__7482(csa_tree_add_7_25_groupi_n_7205 ,csa_tree_add_7_25_groupi_n_7157 ,csa_tree_add_7_25_groupi_n_7168);
  nor csa_tree_add_7_25_groupi_g13883__4733(csa_tree_add_7_25_groupi_n_7204 ,csa_tree_add_7_25_groupi_n_7143 ,csa_tree_add_7_25_groupi_n_7167);
  and csa_tree_add_7_25_groupi_g13884__6161(csa_tree_add_7_25_groupi_n_7203 ,csa_tree_add_7_25_groupi_n_7150 ,csa_tree_add_7_25_groupi_n_7164);
  or csa_tree_add_7_25_groupi_g13885__9315(csa_tree_add_7_25_groupi_n_7202 ,csa_tree_add_7_25_groupi_n_7150 ,csa_tree_add_7_25_groupi_n_7164);
  and csa_tree_add_7_25_groupi_g13886__9945(csa_tree_add_7_25_groupi_n_7201 ,csa_tree_add_7_25_groupi_n_7157 ,csa_tree_add_7_25_groupi_n_7168);
  or csa_tree_add_7_25_groupi_g13887__2883(csa_tree_add_7_25_groupi_n_7200 ,csa_tree_add_7_25_groupi_n_7141 ,csa_tree_add_7_25_groupi_n_7162);
  or csa_tree_add_7_25_groupi_g13888__2346(csa_tree_add_7_25_groupi_n_7199 ,csa_tree_add_7_25_groupi_n_7157 ,csa_tree_add_7_25_groupi_n_7168);
  and csa_tree_add_7_25_groupi_g13889__1666(csa_tree_add_7_25_groupi_n_7198 ,csa_tree_add_7_25_groupi_n_7163 ,csa_tree_add_7_25_groupi_n_7140);
  or csa_tree_add_7_25_groupi_g13890__7410(csa_tree_add_7_25_groupi_n_7197 ,csa_tree_add_7_25_groupi_n_7163 ,csa_tree_add_7_25_groupi_n_7140);
  nor csa_tree_add_7_25_groupi_g13891__6417(csa_tree_add_7_25_groupi_n_7196 ,csa_tree_add_7_25_groupi_n_7171 ,csa_tree_add_7_25_groupi_n_7145);
  and csa_tree_add_7_25_groupi_g13892__5477(csa_tree_add_7_25_groupi_n_7195 ,csa_tree_add_7_25_groupi_n_7141 ,csa_tree_add_7_25_groupi_n_7162);
  or csa_tree_add_7_25_groupi_g13893__2398(csa_tree_add_7_25_groupi_n_7194 ,csa_tree_add_7_25_groupi_n_7170 ,csa_tree_add_7_25_groupi_n_7144);
  or csa_tree_add_7_25_groupi_g13894__5107(csa_tree_add_7_25_groupi_n_7192 ,csa_tree_add_7_25_groupi_n_7169 ,csa_tree_add_7_25_groupi_n_7146);
  or csa_tree_add_7_25_groupi_g13895__6260(csa_tree_add_7_25_groupi_n_7191 ,csa_tree_add_7_25_groupi_n_7142 ,csa_tree_add_7_25_groupi_n_7166);
  and csa_tree_add_7_25_groupi_g13896__4319(csa_tree_add_7_25_groupi_n_7190 ,csa_tree_add_7_25_groupi_n_7154 ,csa_tree_add_7_25_groupi_n_7165);
  or csa_tree_add_7_25_groupi_g13897__8428(csa_tree_add_7_25_groupi_n_7189 ,csa_tree_add_7_25_groupi_n_7154 ,csa_tree_add_7_25_groupi_n_7165);
  and csa_tree_add_7_25_groupi_g13898__5526(csa_tree_add_7_25_groupi_n_7188 ,csa_tree_add_7_25_groupi_n_7169 ,csa_tree_add_7_25_groupi_n_7146);
  xnor csa_tree_add_7_25_groupi_g13899__6783(csa_tree_add_7_25_groupi_n_7187 ,csa_tree_add_7_25_groupi_n_7155 ,csa_tree_add_7_25_groupi_n_7131);
  xnor csa_tree_add_7_25_groupi_g13900__3680(csa_tree_add_7_25_groupi_n_7186 ,csa_tree_add_7_25_groupi_n_7133 ,csa_tree_add_7_25_groupi_n_7139);
  xnor csa_tree_add_7_25_groupi_g13901__1617(csa_tree_add_7_25_groupi_n_7185 ,csa_tree_add_7_25_groupi_n_7135 ,csa_tree_add_7_25_groupi_n_7153);
  xnor csa_tree_add_7_25_groupi_g13902__2802(csa_tree_add_7_25_groupi_n_7184 ,csa_tree_add_7_25_groupi_n_7136 ,csa_tree_add_7_25_groupi_n_7130);
  xnor csa_tree_add_7_25_groupi_g13903__1705(csa_tree_add_7_25_groupi_n_7183 ,csa_tree_add_7_25_groupi_n_7151 ,csa_tree_add_7_25_groupi_n_7137);
  or csa_tree_add_7_25_groupi_g13904__5122(csa_tree_add_7_25_groupi_n_7193 ,csa_tree_add_7_25_groupi_n_7148 ,csa_tree_add_7_25_groupi_n_7180);
  and csa_tree_add_7_25_groupi_g13905__8246(csa_tree_add_7_25_groupi_n_7182 ,csa_tree_add_7_25_groupi_n_7156 ,csa_tree_add_7_25_groupi_n_7131);
  and csa_tree_add_7_25_groupi_g13906__7098(csa_tree_add_7_25_groupi_n_7181 ,csa_tree_add_7_25_groupi_n_7151 ,csa_tree_add_7_25_groupi_n_7137);
  and csa_tree_add_7_25_groupi_g13907__6131(csa_tree_add_7_25_groupi_n_7180 ,csa_tree_add_7_25_groupi_n_7149 ,csa_tree_add_7_25_groupi_n_7158);
  or csa_tree_add_7_25_groupi_g13908__1881(csa_tree_add_7_25_groupi_n_7179 ,csa_tree_add_7_25_groupi_n_7136 ,csa_tree_add_7_25_groupi_n_7130);
  and csa_tree_add_7_25_groupi_g13909__5115(csa_tree_add_7_25_groupi_n_7178 ,csa_tree_add_7_25_groupi_n_7136 ,csa_tree_add_7_25_groupi_n_7130);
  or csa_tree_add_7_25_groupi_g13910__7482(csa_tree_add_7_25_groupi_n_7177 ,csa_tree_add_7_25_groupi_n_7151 ,csa_tree_add_7_25_groupi_n_7137);
  nor csa_tree_add_7_25_groupi_g13911__4733(csa_tree_add_7_25_groupi_n_7176 ,csa_tree_add_7_25_groupi_n_7156 ,csa_tree_add_7_25_groupi_n_7131);
  or csa_tree_add_7_25_groupi_g13912__6161(csa_tree_add_7_25_groupi_n_7175 ,csa_tree_add_7_25_groupi_n_7135 ,csa_tree_add_7_25_groupi_n_7152);
  nor csa_tree_add_7_25_groupi_g13913__9315(csa_tree_add_7_25_groupi_n_7174 ,csa_tree_add_7_25_groupi_n_7134 ,csa_tree_add_7_25_groupi_n_7153);
  nor csa_tree_add_7_25_groupi_g13914__9945(csa_tree_add_7_25_groupi_n_7173 ,csa_tree_add_7_25_groupi_n_7132 ,csa_tree_add_7_25_groupi_n_7139);
  or csa_tree_add_7_25_groupi_g13915__2883(csa_tree_add_7_25_groupi_n_7172 ,csa_tree_add_7_25_groupi_n_7133 ,csa_tree_add_7_25_groupi_n_7138);
  not csa_tree_add_7_25_groupi_g13916(csa_tree_add_7_25_groupi_n_7170 ,csa_tree_add_7_25_groupi_n_7171);
  not csa_tree_add_7_25_groupi_g13917(csa_tree_add_7_25_groupi_n_7166 ,csa_tree_add_7_25_groupi_n_7167);
  xnor csa_tree_add_7_25_groupi_g13918__2346(out2[25] ,csa_tree_add_7_25_groupi_n_7103 ,csa_tree_add_7_25_groupi_n_7104);
  xnor csa_tree_add_7_25_groupi_g13919__1666(csa_tree_add_7_25_groupi_n_7160 ,csa_tree_add_7_25_groupi_n_7048 ,csa_tree_add_7_25_groupi_n_7110);
  xnor csa_tree_add_7_25_groupi_g13920__7410(csa_tree_add_7_25_groupi_n_7159 ,csa_tree_add_7_25_groupi_n_7117 ,csa_tree_add_7_25_groupi_n_7073);
  xnor csa_tree_add_7_25_groupi_g13921__6417(csa_tree_add_7_25_groupi_n_7171 ,csa_tree_add_7_25_groupi_n_7053 ,csa_tree_add_7_25_groupi_n_7108);
  xnor csa_tree_add_7_25_groupi_g13922__5477(csa_tree_add_7_25_groupi_n_7169 ,csa_tree_add_7_25_groupi_n_7075 ,csa_tree_add_7_25_groupi_n_7105);
  xnor csa_tree_add_7_25_groupi_g13923__2398(csa_tree_add_7_25_groupi_n_7168 ,csa_tree_add_7_25_groupi_n_7055 ,csa_tree_add_7_25_groupi_n_7106);
  xnor csa_tree_add_7_25_groupi_g13924__5107(csa_tree_add_7_25_groupi_n_7167 ,csa_tree_add_7_25_groupi_n_7057 ,csa_tree_add_7_25_groupi_n_7109);
  xnor csa_tree_add_7_25_groupi_g13925__6260(csa_tree_add_7_25_groupi_n_7165 ,csa_tree_add_7_25_groupi_n_7050 ,csa_tree_add_7_25_groupi_n_7107);
  xnor csa_tree_add_7_25_groupi_g13926__4319(csa_tree_add_7_25_groupi_n_7164 ,csa_tree_add_7_25_groupi_n_7077 ,csa_tree_add_7_25_groupi_n_7113);
  xnor csa_tree_add_7_25_groupi_g13927__8428(csa_tree_add_7_25_groupi_n_7163 ,csa_tree_add_7_25_groupi_n_7078 ,csa_tree_add_7_25_groupi_n_7112);
  xnor csa_tree_add_7_25_groupi_g13928__5526(csa_tree_add_7_25_groupi_n_7162 ,csa_tree_add_7_25_groupi_n_7074 ,csa_tree_add_7_25_groupi_n_7111);
  not csa_tree_add_7_25_groupi_g13929(csa_tree_add_7_25_groupi_n_7156 ,csa_tree_add_7_25_groupi_n_7155);
  not csa_tree_add_7_25_groupi_g13930(csa_tree_add_7_25_groupi_n_7152 ,csa_tree_add_7_25_groupi_n_7153);
  or csa_tree_add_7_25_groupi_g13931__6783(csa_tree_add_7_25_groupi_n_7149 ,csa_tree_add_7_25_groupi_n_7117 ,csa_tree_add_7_25_groupi_n_7073);
  and csa_tree_add_7_25_groupi_g13932__3680(csa_tree_add_7_25_groupi_n_7148 ,csa_tree_add_7_25_groupi_n_7117 ,csa_tree_add_7_25_groupi_n_7073);
  or csa_tree_add_7_25_groupi_g13933__1617(csa_tree_add_7_25_groupi_n_7147 ,csa_tree_add_7_25_groupi_n_7030 ,csa_tree_add_7_25_groupi_n_7126);
  or csa_tree_add_7_25_groupi_g13934__2802(csa_tree_add_7_25_groupi_n_7158 ,csa_tree_add_7_25_groupi_n_7128 ,csa_tree_add_7_25_groupi_n_7101);
  or csa_tree_add_7_25_groupi_g13935__1705(csa_tree_add_7_25_groupi_n_7157 ,csa_tree_add_7_25_groupi_n_7040 ,csa_tree_add_7_25_groupi_n_7129);
  or csa_tree_add_7_25_groupi_g13936__5122(csa_tree_add_7_25_groupi_n_7155 ,csa_tree_add_7_25_groupi_n_7125 ,csa_tree_add_7_25_groupi_n_7102);
  or csa_tree_add_7_25_groupi_g13937__8246(csa_tree_add_7_25_groupi_n_7154 ,csa_tree_add_7_25_groupi_n_7023 ,csa_tree_add_7_25_groupi_n_7124);
  or csa_tree_add_7_25_groupi_g13938__7098(csa_tree_add_7_25_groupi_n_7153 ,csa_tree_add_7_25_groupi_n_7094 ,csa_tree_add_7_25_groupi_n_7122);
  or csa_tree_add_7_25_groupi_g13939__6131(csa_tree_add_7_25_groupi_n_7151 ,csa_tree_add_7_25_groupi_n_7121 ,csa_tree_add_7_25_groupi_n_7083);
  and csa_tree_add_7_25_groupi_g13940__1881(csa_tree_add_7_25_groupi_n_7150 ,csa_tree_add_7_25_groupi_n_7092 ,csa_tree_add_7_25_groupi_n_7120);
  not csa_tree_add_7_25_groupi_g13941(csa_tree_add_7_25_groupi_n_7144 ,csa_tree_add_7_25_groupi_n_7145);
  not csa_tree_add_7_25_groupi_g13942(csa_tree_add_7_25_groupi_n_7142 ,csa_tree_add_7_25_groupi_n_7143);
  not csa_tree_add_7_25_groupi_g13943(csa_tree_add_7_25_groupi_n_7138 ,csa_tree_add_7_25_groupi_n_7139);
  not csa_tree_add_7_25_groupi_g13944(csa_tree_add_7_25_groupi_n_7134 ,csa_tree_add_7_25_groupi_n_7135);
  not csa_tree_add_7_25_groupi_g13945(csa_tree_add_7_25_groupi_n_7132 ,csa_tree_add_7_25_groupi_n_7133);
  or csa_tree_add_7_25_groupi_g13946__5115(csa_tree_add_7_25_groupi_n_7146 ,csa_tree_add_7_25_groupi_n_7080 ,csa_tree_add_7_25_groupi_n_7116);
  or csa_tree_add_7_25_groupi_g13947__7482(csa_tree_add_7_25_groupi_n_7145 ,csa_tree_add_7_25_groupi_n_7028 ,csa_tree_add_7_25_groupi_n_7118);
  or csa_tree_add_7_25_groupi_g13948__4733(csa_tree_add_7_25_groupi_n_7143 ,csa_tree_add_7_25_groupi_n_7021 ,csa_tree_add_7_25_groupi_n_7123);
  and csa_tree_add_7_25_groupi_g13949__6161(csa_tree_add_7_25_groupi_n_7141 ,csa_tree_add_7_25_groupi_n_7098 ,csa_tree_add_7_25_groupi_n_7127);
  and csa_tree_add_7_25_groupi_g13950__9315(csa_tree_add_7_25_groupi_n_7140 ,csa_tree_add_7_25_groupi_n_7114 ,csa_tree_add_7_25_groupi_n_7084);
  or csa_tree_add_7_25_groupi_g13951__9945(csa_tree_add_7_25_groupi_n_7139 ,csa_tree_add_7_25_groupi_n_7082 ,csa_tree_add_7_25_groupi_n_7119);
  xnor csa_tree_add_7_25_groupi_g13952__2883(csa_tree_add_7_25_groupi_n_7137 ,csa_tree_add_7_25_groupi_n_7091 ,csa_tree_add_7_25_groupi_n_7047);
  xnor csa_tree_add_7_25_groupi_g13953__2346(csa_tree_add_7_25_groupi_n_7136 ,csa_tree_add_7_25_groupi_n_7089 ,csa_tree_add_7_25_groupi_n_7046);
  xnor csa_tree_add_7_25_groupi_g13954__1666(csa_tree_add_7_25_groupi_n_7135 ,csa_tree_add_7_25_groupi_n_7090 ,csa_tree_add_7_25_groupi_n_7062);
  xnor csa_tree_add_7_25_groupi_g13955__7410(csa_tree_add_7_25_groupi_n_7133 ,csa_tree_add_7_25_groupi_n_7088 ,csa_tree_add_7_25_groupi_n_7063);
  xnor csa_tree_add_7_25_groupi_g13956__6417(csa_tree_add_7_25_groupi_n_7131 ,csa_tree_add_7_25_groupi_n_7087 ,csa_tree_add_7_25_groupi_n_7064);
  and csa_tree_add_7_25_groupi_g13957__5477(csa_tree_add_7_25_groupi_n_7129 ,csa_tree_add_7_25_groupi_n_7091 ,csa_tree_add_7_25_groupi_n_7041);
  and csa_tree_add_7_25_groupi_g13958__2398(csa_tree_add_7_25_groupi_n_7128 ,csa_tree_add_7_25_groupi_n_7103 ,csa_tree_add_7_25_groupi_n_7096);
  or csa_tree_add_7_25_groupi_g13959__5107(csa_tree_add_7_25_groupi_n_7127 ,csa_tree_add_7_25_groupi_n_7095 ,csa_tree_add_7_25_groupi_n_7059);
  and csa_tree_add_7_25_groupi_g13960__6260(csa_tree_add_7_25_groupi_n_7126 ,csa_tree_add_7_25_groupi_n_7087 ,csa_tree_add_7_25_groupi_n_7031);
  and csa_tree_add_7_25_groupi_g13961__4319(csa_tree_add_7_25_groupi_n_7125 ,csa_tree_add_7_25_groupi_n_7097 ,csa_tree_add_7_25_groupi_n_7074);
  and csa_tree_add_7_25_groupi_g13962__8428(csa_tree_add_7_25_groupi_n_7124 ,csa_tree_add_7_25_groupi_n_7089 ,csa_tree_add_7_25_groupi_n_7022);
  and csa_tree_add_7_25_groupi_g13963__5526(csa_tree_add_7_25_groupi_n_7123 ,csa_tree_add_7_25_groupi_n_7090 ,csa_tree_add_7_25_groupi_n_7032);
  and csa_tree_add_7_25_groupi_g13964__6783(csa_tree_add_7_25_groupi_n_7122 ,csa_tree_add_7_25_groupi_n_7093 ,csa_tree_add_7_25_groupi_n_7077);
  and csa_tree_add_7_25_groupi_g13965__3680(csa_tree_add_7_25_groupi_n_7121 ,csa_tree_add_7_25_groupi_n_7075 ,csa_tree_add_7_25_groupi_n_7086);
  or csa_tree_add_7_25_groupi_g13966__1617(csa_tree_add_7_25_groupi_n_7120 ,csa_tree_add_7_25_groupi_n_7100 ,csa_tree_add_7_25_groupi_n_7060);
  and csa_tree_add_7_25_groupi_g13967__2802(csa_tree_add_7_25_groupi_n_7119 ,csa_tree_add_7_25_groupi_n_7078 ,csa_tree_add_7_25_groupi_n_7081);
  and csa_tree_add_7_25_groupi_g13968__1705(csa_tree_add_7_25_groupi_n_7118 ,csa_tree_add_7_25_groupi_n_7088 ,csa_tree_add_7_25_groupi_n_7027);
  or csa_tree_add_7_25_groupi_g13969__5122(csa_tree_add_7_25_groupi_n_7130 ,csa_tree_add_7_25_groupi_n_6959 ,csa_tree_add_7_25_groupi_n_7099);
  nor csa_tree_add_7_25_groupi_g13970__8246(csa_tree_add_7_25_groupi_n_7116 ,csa_tree_add_7_25_groupi_n_7079 ,csa_tree_add_7_25_groupi_n_7061);
  xnor csa_tree_add_7_25_groupi_g13971__7098(out2[24] ,csa_tree_add_7_25_groupi_n_7043 ,csa_tree_add_7_25_groupi_n_7044);
  or csa_tree_add_7_25_groupi_g13972__6131(csa_tree_add_7_25_groupi_n_7114 ,csa_tree_add_7_25_groupi_n_7085 ,csa_tree_add_7_25_groupi_n_7058);
  xnor csa_tree_add_7_25_groupi_g13973__1881(csa_tree_add_7_25_groupi_n_7113 ,csa_tree_add_7_25_groupi_n_7071 ,csa_tree_add_7_25_groupi_n_6984);
  xnor csa_tree_add_7_25_groupi_g13974__5115(csa_tree_add_7_25_groupi_n_7112 ,csa_tree_add_7_25_groupi_n_7069 ,csa_tree_add_7_25_groupi_n_6982);
  xnor csa_tree_add_7_25_groupi_g13975__7482(csa_tree_add_7_25_groupi_n_7111 ,csa_tree_add_7_25_groupi_n_7067 ,csa_tree_add_7_25_groupi_n_6980);
  xnor csa_tree_add_7_25_groupi_g13976__4733(csa_tree_add_7_25_groupi_n_7110 ,csa_tree_add_7_25_groupi_n_6998 ,csa_tree_add_7_25_groupi_n_7045);
  xnor csa_tree_add_7_25_groupi_g13977__6161(csa_tree_add_7_25_groupi_n_7109 ,csa_tree_add_7_25_groupi_n_7018 ,csa_tree_add_7_25_groupi_n_7058);
  xnor csa_tree_add_7_25_groupi_g13978__9315(csa_tree_add_7_25_groupi_n_7108 ,csa_tree_add_7_25_groupi_n_7020 ,csa_tree_add_7_25_groupi_n_7059);
  xnor csa_tree_add_7_25_groupi_g13979__9945(csa_tree_add_7_25_groupi_n_7107 ,csa_tree_add_7_25_groupi_n_7015 ,csa_tree_add_7_25_groupi_n_7061);
  xnor csa_tree_add_7_25_groupi_g13980__2883(csa_tree_add_7_25_groupi_n_7106 ,csa_tree_add_7_25_groupi_n_7013 ,csa_tree_add_7_25_groupi_n_7060);
  xnor csa_tree_add_7_25_groupi_g13981__2346(csa_tree_add_7_25_groupi_n_7105 ,csa_tree_add_7_25_groupi_n_7072 ,csa_tree_add_7_25_groupi_n_6991);
  xnor csa_tree_add_7_25_groupi_g13982__1666(csa_tree_add_7_25_groupi_n_7104 ,csa_tree_add_7_25_groupi_n_7014 ,csa_tree_add_7_25_groupi_n_7051);
  xnor csa_tree_add_7_25_groupi_g13983__7410(csa_tree_add_7_25_groupi_n_7117 ,csa_tree_add_7_25_groupi_n_7076 ,csa_tree_add_7_25_groupi_n_6971);
  nor csa_tree_add_7_25_groupi_g13984__6417(csa_tree_add_7_25_groupi_n_7102 ,csa_tree_add_7_25_groupi_n_7066 ,csa_tree_add_7_25_groupi_n_6980);
  and csa_tree_add_7_25_groupi_g13985__5477(csa_tree_add_7_25_groupi_n_7101 ,csa_tree_add_7_25_groupi_n_7014 ,csa_tree_add_7_25_groupi_n_7051);
  nor csa_tree_add_7_25_groupi_g13986__2398(csa_tree_add_7_25_groupi_n_7100 ,csa_tree_add_7_25_groupi_n_7054 ,csa_tree_add_7_25_groupi_n_7013);
  and csa_tree_add_7_25_groupi_g13987__5107(csa_tree_add_7_25_groupi_n_7099 ,csa_tree_add_7_25_groupi_n_7076 ,csa_tree_add_7_25_groupi_n_6958);
  or csa_tree_add_7_25_groupi_g13988__6260(csa_tree_add_7_25_groupi_n_7098 ,csa_tree_add_7_25_groupi_n_7053 ,csa_tree_add_7_25_groupi_n_7019);
  or csa_tree_add_7_25_groupi_g13989__4319(csa_tree_add_7_25_groupi_n_7097 ,csa_tree_add_7_25_groupi_n_7067 ,csa_tree_add_7_25_groupi_n_6979);
  or csa_tree_add_7_25_groupi_g13990__8428(csa_tree_add_7_25_groupi_n_7096 ,csa_tree_add_7_25_groupi_n_7014 ,csa_tree_add_7_25_groupi_n_7051);
  nor csa_tree_add_7_25_groupi_g13991__5526(csa_tree_add_7_25_groupi_n_7095 ,csa_tree_add_7_25_groupi_n_7052 ,csa_tree_add_7_25_groupi_n_7020);
  nor csa_tree_add_7_25_groupi_g13992__6783(csa_tree_add_7_25_groupi_n_7094 ,csa_tree_add_7_25_groupi_n_7070 ,csa_tree_add_7_25_groupi_n_6984);
  or csa_tree_add_7_25_groupi_g13993__3680(csa_tree_add_7_25_groupi_n_7093 ,csa_tree_add_7_25_groupi_n_7071 ,csa_tree_add_7_25_groupi_n_6983);
  or csa_tree_add_7_25_groupi_g13994__1617(csa_tree_add_7_25_groupi_n_7092 ,csa_tree_add_7_25_groupi_n_7055 ,csa_tree_add_7_25_groupi_n_7012);
  or csa_tree_add_7_25_groupi_g13995__2802(csa_tree_add_7_25_groupi_n_7103 ,csa_tree_add_7_25_groupi_n_7065 ,csa_tree_add_7_25_groupi_n_7039);
  or csa_tree_add_7_25_groupi_g13996__1705(csa_tree_add_7_25_groupi_n_7086 ,csa_tree_add_7_25_groupi_n_7072 ,csa_tree_add_7_25_groupi_n_6991);
  nor csa_tree_add_7_25_groupi_g13997__5122(csa_tree_add_7_25_groupi_n_7085 ,csa_tree_add_7_25_groupi_n_7056 ,csa_tree_add_7_25_groupi_n_7018);
  or csa_tree_add_7_25_groupi_g13998__8246(csa_tree_add_7_25_groupi_n_7084 ,csa_tree_add_7_25_groupi_n_7057 ,csa_tree_add_7_25_groupi_n_7017);
  and csa_tree_add_7_25_groupi_g13999__7098(csa_tree_add_7_25_groupi_n_7083 ,csa_tree_add_7_25_groupi_n_7072 ,csa_tree_add_7_25_groupi_n_6991);
  nor csa_tree_add_7_25_groupi_g14000__6131(csa_tree_add_7_25_groupi_n_7082 ,csa_tree_add_7_25_groupi_n_7068 ,csa_tree_add_7_25_groupi_n_6982);
  or csa_tree_add_7_25_groupi_g14001__1881(csa_tree_add_7_25_groupi_n_7081 ,csa_tree_add_7_25_groupi_n_7069 ,csa_tree_add_7_25_groupi_n_6981);
  nor csa_tree_add_7_25_groupi_g14002__5115(csa_tree_add_7_25_groupi_n_7080 ,csa_tree_add_7_25_groupi_n_7050 ,csa_tree_add_7_25_groupi_n_7016);
  and csa_tree_add_7_25_groupi_g14003__7482(csa_tree_add_7_25_groupi_n_7079 ,csa_tree_add_7_25_groupi_n_7050 ,csa_tree_add_7_25_groupi_n_7016);
  xnor csa_tree_add_7_25_groupi_g14004__4733(csa_tree_add_7_25_groupi_n_7091 ,csa_tree_add_7_25_groupi_n_7034 ,in3[5]);
  xnor csa_tree_add_7_25_groupi_g14005__6161(csa_tree_add_7_25_groupi_n_7090 ,csa_tree_add_7_25_groupi_n_7033 ,in3[8]);
  xnor csa_tree_add_7_25_groupi_g14006__9315(csa_tree_add_7_25_groupi_n_7089 ,csa_tree_add_7_25_groupi_n_7035 ,in3[2]);
  xnor csa_tree_add_7_25_groupi_g14007__9945(csa_tree_add_7_25_groupi_n_7088 ,csa_tree_add_7_25_groupi_n_7036 ,in3[11]);
  xnor csa_tree_add_7_25_groupi_g14008__2883(csa_tree_add_7_25_groupi_n_7087 ,csa_tree_add_7_25_groupi_n_7037 ,in3[14]);
  not csa_tree_add_7_25_groupi_g14009(csa_tree_add_7_25_groupi_n_7070 ,csa_tree_add_7_25_groupi_n_7071);
  not csa_tree_add_7_25_groupi_g14010(csa_tree_add_7_25_groupi_n_7068 ,csa_tree_add_7_25_groupi_n_7069);
  not csa_tree_add_7_25_groupi_g14011(csa_tree_add_7_25_groupi_n_7066 ,csa_tree_add_7_25_groupi_n_7067);
  and csa_tree_add_7_25_groupi_g14012__2346(csa_tree_add_7_25_groupi_n_7065 ,csa_tree_add_7_25_groupi_n_7043 ,csa_tree_add_7_25_groupi_n_7042);
  xnor csa_tree_add_7_25_groupi_g14013__1666(csa_tree_add_7_25_groupi_n_7064 ,csa_tree_add_7_25_groupi_n_6989 ,csa_tree_add_7_25_groupi_n_6953);
  xnor csa_tree_add_7_25_groupi_g14014__7410(csa_tree_add_7_25_groupi_n_7063 ,csa_tree_add_7_25_groupi_n_6956 ,csa_tree_add_7_25_groupi_n_6978);
  xnor csa_tree_add_7_25_groupi_g14015__6417(csa_tree_add_7_25_groupi_n_7062 ,csa_tree_add_7_25_groupi_n_6951 ,csa_tree_add_7_25_groupi_n_6986);
  or csa_tree_add_7_25_groupi_g14016__5477(csa_tree_add_7_25_groupi_n_7078 ,csa_tree_add_7_25_groupi_n_6879 ,csa_tree_add_7_25_groupi_n_7024);
  or csa_tree_add_7_25_groupi_g14017__2398(csa_tree_add_7_25_groupi_n_7077 ,csa_tree_add_7_25_groupi_n_6874 ,csa_tree_add_7_25_groupi_n_7025);
  xnor csa_tree_add_7_25_groupi_g14018__5107(csa_tree_add_7_25_groupi_n_7076 ,csa_tree_add_7_25_groupi_n_7005 ,in3[2]);
  or csa_tree_add_7_25_groupi_g14019__6260(csa_tree_add_7_25_groupi_n_7075 ,csa_tree_add_7_25_groupi_n_6888 ,csa_tree_add_7_25_groupi_n_7038);
  or csa_tree_add_7_25_groupi_g14020__4319(csa_tree_add_7_25_groupi_n_7074 ,csa_tree_add_7_25_groupi_n_6882 ,csa_tree_add_7_25_groupi_n_7029);
  or csa_tree_add_7_25_groupi_g14021__8428(csa_tree_add_7_25_groupi_n_7073 ,csa_tree_add_7_25_groupi_n_6890 ,csa_tree_add_7_25_groupi_n_7026);
  xnor csa_tree_add_7_25_groupi_g14022__5526(csa_tree_add_7_25_groupi_n_7072 ,csa_tree_add_7_25_groupi_n_6999 ,in3[5]);
  xnor csa_tree_add_7_25_groupi_g14023__6783(csa_tree_add_7_25_groupi_n_7071 ,csa_tree_add_7_25_groupi_n_7000 ,in3[8]);
  xnor csa_tree_add_7_25_groupi_g14024__3680(csa_tree_add_7_25_groupi_n_7069 ,csa_tree_add_7_25_groupi_n_6997 ,in3[11]);
  xnor csa_tree_add_7_25_groupi_g14025__1617(csa_tree_add_7_25_groupi_n_7067 ,csa_tree_add_7_25_groupi_n_7006 ,in3[14]);
  not csa_tree_add_7_25_groupi_g14026(csa_tree_add_7_25_groupi_n_7056 ,csa_tree_add_7_25_groupi_n_7057);
  not csa_tree_add_7_25_groupi_g14027(csa_tree_add_7_25_groupi_n_7054 ,csa_tree_add_7_25_groupi_n_7055);
  not csa_tree_add_7_25_groupi_g14028(csa_tree_add_7_25_groupi_n_7052 ,csa_tree_add_7_25_groupi_n_7053);
  xnor csa_tree_add_7_25_groupi_g14029__2802(out2[23] ,csa_tree_add_7_25_groupi_n_6969 ,csa_tree_add_7_25_groupi_n_6972);
  xnor csa_tree_add_7_25_groupi_g14030__1705(csa_tree_add_7_25_groupi_n_7048 ,csa_tree_add_7_25_groupi_n_7004 ,in3[14]);
  xnor csa_tree_add_7_25_groupi_g14031__5122(csa_tree_add_7_25_groupi_n_7047 ,csa_tree_add_7_25_groupi_n_6954 ,csa_tree_add_7_25_groupi_n_6976);
  xnor csa_tree_add_7_25_groupi_g14032__8246(csa_tree_add_7_25_groupi_n_7046 ,csa_tree_add_7_25_groupi_n_6990 ,csa_tree_add_7_25_groupi_n_6940);
  xnor csa_tree_add_7_25_groupi_g14033__7098(csa_tree_add_7_25_groupi_n_7045 ,csa_tree_add_7_25_groupi_n_6970 ,csa_tree_add_7_25_groupi_n_6908);
  xnor csa_tree_add_7_25_groupi_g14034__6131(csa_tree_add_7_25_groupi_n_7044 ,csa_tree_add_7_25_groupi_n_6987 ,csa_tree_add_7_25_groupi_n_6939);
  xnor csa_tree_add_7_25_groupi_g14035__1881(csa_tree_add_7_25_groupi_n_7061 ,csa_tree_add_7_25_groupi_n_6996 ,csa_tree_add_7_25_groupi_n_6904);
  xnor csa_tree_add_7_25_groupi_g14036__5115(csa_tree_add_7_25_groupi_n_7060 ,csa_tree_add_7_25_groupi_n_6992 ,csa_tree_add_7_25_groupi_n_6911);
  xnor csa_tree_add_7_25_groupi_g14037__7482(csa_tree_add_7_25_groupi_n_7059 ,csa_tree_add_7_25_groupi_n_6995 ,csa_tree_add_7_25_groupi_n_6905);
  xnor csa_tree_add_7_25_groupi_g14038__4733(csa_tree_add_7_25_groupi_n_7058 ,csa_tree_add_7_25_groupi_n_6993 ,csa_tree_add_7_25_groupi_n_6907);
  xnor csa_tree_add_7_25_groupi_g14039__6161(csa_tree_add_7_25_groupi_n_7057 ,csa_tree_add_7_25_groupi_n_7003 ,in3[8]);
  xnor csa_tree_add_7_25_groupi_g14040__9315(csa_tree_add_7_25_groupi_n_7055 ,csa_tree_add_7_25_groupi_n_7001 ,in3[5]);
  xnor csa_tree_add_7_25_groupi_g14041__9945(csa_tree_add_7_25_groupi_n_7053 ,csa_tree_add_7_25_groupi_n_7002 ,in3[11]);
  xnor csa_tree_add_7_25_groupi_g14042__2883(csa_tree_add_7_25_groupi_n_7051 ,csa_tree_add_7_25_groupi_n_6994 ,csa_tree_add_7_25_groupi_n_6901);
  xnor csa_tree_add_7_25_groupi_g14043__2346(csa_tree_add_7_25_groupi_n_7050 ,csa_tree_add_7_25_groupi_n_7007 ,in3[2]);
  or csa_tree_add_7_25_groupi_g14044__1666(csa_tree_add_7_25_groupi_n_7042 ,csa_tree_add_7_25_groupi_n_6987 ,csa_tree_add_7_25_groupi_n_6939);
  or csa_tree_add_7_25_groupi_g14045__7410(csa_tree_add_7_25_groupi_n_7041 ,csa_tree_add_7_25_groupi_n_6954 ,csa_tree_add_7_25_groupi_n_6976);
  and csa_tree_add_7_25_groupi_g14046__6417(csa_tree_add_7_25_groupi_n_7040 ,csa_tree_add_7_25_groupi_n_6954 ,csa_tree_add_7_25_groupi_n_6976);
  and csa_tree_add_7_25_groupi_g14047__5477(csa_tree_add_7_25_groupi_n_7039 ,csa_tree_add_7_25_groupi_n_6987 ,csa_tree_add_7_25_groupi_n_6939);
  and csa_tree_add_7_25_groupi_g14048__2398(csa_tree_add_7_25_groupi_n_7038 ,csa_tree_add_7_25_groupi_n_6996 ,csa_tree_add_7_25_groupi_n_6886);
  nor csa_tree_add_7_25_groupi_g14049__5107(csa_tree_add_7_25_groupi_n_7037 ,csa_tree_add_7_25_groupi_n_4033 ,csa_tree_add_7_25_groupi_n_7009);
  nor csa_tree_add_7_25_groupi_g14050__6260(csa_tree_add_7_25_groupi_n_7036 ,csa_tree_add_7_25_groupi_n_3993 ,csa_tree_add_7_25_groupi_n_6975);
  nor csa_tree_add_7_25_groupi_g14051__4319(csa_tree_add_7_25_groupi_n_7035 ,csa_tree_add_7_25_groupi_n_3475 ,csa_tree_add_7_25_groupi_n_7008);
  nor csa_tree_add_7_25_groupi_g14052__8428(csa_tree_add_7_25_groupi_n_7034 ,csa_tree_add_7_25_groupi_n_3999 ,csa_tree_add_7_25_groupi_n_7011);
  nor csa_tree_add_7_25_groupi_g14053__5526(csa_tree_add_7_25_groupi_n_7033 ,csa_tree_add_7_25_groupi_n_4032 ,csa_tree_add_7_25_groupi_n_6973);
  or csa_tree_add_7_25_groupi_g14054__6783(csa_tree_add_7_25_groupi_n_7043 ,csa_tree_add_7_25_groupi_n_6961 ,csa_tree_add_7_25_groupi_n_7010);
  or csa_tree_add_7_25_groupi_g14055__3680(csa_tree_add_7_25_groupi_n_7032 ,csa_tree_add_7_25_groupi_n_6951 ,csa_tree_add_7_25_groupi_n_6985);
  or csa_tree_add_7_25_groupi_g14056__1617(csa_tree_add_7_25_groupi_n_7031 ,csa_tree_add_7_25_groupi_n_6988 ,csa_tree_add_7_25_groupi_n_6953);
  nor csa_tree_add_7_25_groupi_g14057__2802(csa_tree_add_7_25_groupi_n_7030 ,csa_tree_add_7_25_groupi_n_6989 ,csa_tree_add_7_25_groupi_n_6952);
  and csa_tree_add_7_25_groupi_g14058__1705(csa_tree_add_7_25_groupi_n_7029 ,csa_tree_add_7_25_groupi_n_6995 ,csa_tree_add_7_25_groupi_n_6881);
  nor csa_tree_add_7_25_groupi_g14059__5122(csa_tree_add_7_25_groupi_n_7028 ,csa_tree_add_7_25_groupi_n_6955 ,csa_tree_add_7_25_groupi_n_6978);
  or csa_tree_add_7_25_groupi_g14060__8246(csa_tree_add_7_25_groupi_n_7027 ,csa_tree_add_7_25_groupi_n_6956 ,csa_tree_add_7_25_groupi_n_6977);
  and csa_tree_add_7_25_groupi_g14061__7098(csa_tree_add_7_25_groupi_n_7026 ,csa_tree_add_7_25_groupi_n_6994 ,csa_tree_add_7_25_groupi_n_6896);
  and csa_tree_add_7_25_groupi_g14062__6131(csa_tree_add_7_25_groupi_n_7025 ,csa_tree_add_7_25_groupi_n_6992 ,csa_tree_add_7_25_groupi_n_6873);
  and csa_tree_add_7_25_groupi_g14063__1881(csa_tree_add_7_25_groupi_n_7024 ,csa_tree_add_7_25_groupi_n_6993 ,csa_tree_add_7_25_groupi_n_6878);
  and csa_tree_add_7_25_groupi_g14064__5115(csa_tree_add_7_25_groupi_n_7023 ,csa_tree_add_7_25_groupi_n_6990 ,csa_tree_add_7_25_groupi_n_6940);
  or csa_tree_add_7_25_groupi_g14065__7482(csa_tree_add_7_25_groupi_n_7022 ,csa_tree_add_7_25_groupi_n_6990 ,csa_tree_add_7_25_groupi_n_6940);
  nor csa_tree_add_7_25_groupi_g14066__4733(csa_tree_add_7_25_groupi_n_7021 ,csa_tree_add_7_25_groupi_n_6950 ,csa_tree_add_7_25_groupi_n_6986);
  not csa_tree_add_7_25_groupi_g14067(csa_tree_add_7_25_groupi_n_7019 ,csa_tree_add_7_25_groupi_n_7020);
  not csa_tree_add_7_25_groupi_g14068(csa_tree_add_7_25_groupi_n_7017 ,csa_tree_add_7_25_groupi_n_7018);
  not csa_tree_add_7_25_groupi_g14069(csa_tree_add_7_25_groupi_n_7016 ,csa_tree_add_7_25_groupi_n_7015);
  not csa_tree_add_7_25_groupi_g14070(csa_tree_add_7_25_groupi_n_7012 ,csa_tree_add_7_25_groupi_n_7013);
  nor csa_tree_add_7_25_groupi_g14071__6161(csa_tree_add_7_25_groupi_n_7011 ,csa_tree_add_7_25_groupi_n_2133 ,csa_tree_add_7_25_groupi_n_1115);
  and csa_tree_add_7_25_groupi_g14072__9315(csa_tree_add_7_25_groupi_n_7010 ,csa_tree_add_7_25_groupi_n_6969 ,csa_tree_add_7_25_groupi_n_6962);
  nor csa_tree_add_7_25_groupi_g14073__9945(csa_tree_add_7_25_groupi_n_7009 ,csa_tree_add_7_25_groupi_n_2190 ,csa_tree_add_7_25_groupi_n_6949);
  nor csa_tree_add_7_25_groupi_g14074__2883(csa_tree_add_7_25_groupi_n_7008 ,csa_tree_add_7_25_groupi_n_2175 ,csa_tree_add_7_25_groupi_n_1115);
  or csa_tree_add_7_25_groupi_g14075__2346(csa_tree_add_7_25_groupi_n_7007 ,csa_tree_add_7_25_groupi_n_2811 ,csa_tree_add_7_25_groupi_n_6947);
  nor csa_tree_add_7_25_groupi_g14076__1666(csa_tree_add_7_25_groupi_n_7006 ,csa_tree_add_7_25_groupi_n_4025 ,csa_tree_add_7_25_groupi_n_6967);
  nor csa_tree_add_7_25_groupi_g14077__7410(csa_tree_add_7_25_groupi_n_7005 ,csa_tree_add_7_25_groupi_n_3486 ,csa_tree_add_7_25_groupi_n_6957);
  or csa_tree_add_7_25_groupi_g14078__6417(csa_tree_add_7_25_groupi_n_7004 ,csa_tree_add_7_25_groupi_n_3804 ,csa_tree_add_7_25_groupi_n_6948);
  or csa_tree_add_7_25_groupi_g14079__5477(csa_tree_add_7_25_groupi_n_7003 ,csa_tree_add_7_25_groupi_n_3805 ,csa_tree_add_7_25_groupi_n_6943);
  or csa_tree_add_7_25_groupi_g14080__2398(csa_tree_add_7_25_groupi_n_7002 ,csa_tree_add_7_25_groupi_n_3807 ,csa_tree_add_7_25_groupi_n_6942);
  or csa_tree_add_7_25_groupi_g14081__5107(csa_tree_add_7_25_groupi_n_7001 ,csa_tree_add_7_25_groupi_n_3806 ,csa_tree_add_7_25_groupi_n_6941);
  nor csa_tree_add_7_25_groupi_g14082__6260(csa_tree_add_7_25_groupi_n_7000 ,csa_tree_add_7_25_groupi_n_3916 ,csa_tree_add_7_25_groupi_n_6965);
  nor csa_tree_add_7_25_groupi_g14083__4319(csa_tree_add_7_25_groupi_n_6999 ,csa_tree_add_7_25_groupi_n_3861 ,csa_tree_add_7_25_groupi_n_6966);
  or csa_tree_add_7_25_groupi_g14084__8428(csa_tree_add_7_25_groupi_n_6998 ,csa_tree_add_7_25_groupi_n_6801 ,csa_tree_add_7_25_groupi_n_6963);
  nor csa_tree_add_7_25_groupi_g14085__5526(csa_tree_add_7_25_groupi_n_6997 ,csa_tree_add_7_25_groupi_n_3872 ,csa_tree_add_7_25_groupi_n_6964);
  or csa_tree_add_7_25_groupi_g14086__6783(csa_tree_add_7_25_groupi_n_7020 ,csa_tree_add_7_25_groupi_n_6800 ,csa_tree_add_7_25_groupi_n_6944);
  or csa_tree_add_7_25_groupi_g14087__3680(csa_tree_add_7_25_groupi_n_7018 ,csa_tree_add_7_25_groupi_n_6797 ,csa_tree_add_7_25_groupi_n_6946);
  or csa_tree_add_7_25_groupi_g14088__1617(csa_tree_add_7_25_groupi_n_7015 ,csa_tree_add_7_25_groupi_n_6793 ,csa_tree_add_7_25_groupi_n_6945);
  or csa_tree_add_7_25_groupi_g14089__2802(csa_tree_add_7_25_groupi_n_7014 ,csa_tree_add_7_25_groupi_n_6808 ,csa_tree_add_7_25_groupi_n_6960);
  or csa_tree_add_7_25_groupi_g14090__1705(csa_tree_add_7_25_groupi_n_7013 ,csa_tree_add_7_25_groupi_n_6817 ,csa_tree_add_7_25_groupi_n_6968);
  not csa_tree_add_7_25_groupi_g14091(csa_tree_add_7_25_groupi_n_6988 ,csa_tree_add_7_25_groupi_n_6989);
  not csa_tree_add_7_25_groupi_g14092(csa_tree_add_7_25_groupi_n_6985 ,csa_tree_add_7_25_groupi_n_6986);
  not csa_tree_add_7_25_groupi_g14093(csa_tree_add_7_25_groupi_n_6983 ,csa_tree_add_7_25_groupi_n_6984);
  not csa_tree_add_7_25_groupi_g14094(csa_tree_add_7_25_groupi_n_6981 ,csa_tree_add_7_25_groupi_n_6982);
  not csa_tree_add_7_25_groupi_g14095(csa_tree_add_7_25_groupi_n_6979 ,csa_tree_add_7_25_groupi_n_6980);
  not csa_tree_add_7_25_groupi_g14096(csa_tree_add_7_25_groupi_n_6977 ,csa_tree_add_7_25_groupi_n_6978);
  nor csa_tree_add_7_25_groupi_g14097__5122(csa_tree_add_7_25_groupi_n_6975 ,csa_tree_add_7_25_groupi_n_2097 ,csa_tree_add_7_25_groupi_n_6949);
  xnor csa_tree_add_7_25_groupi_g14098__8246(out2[22] ,csa_tree_add_7_25_groupi_n_6898 ,csa_tree_add_7_25_groupi_n_6903);
  nor csa_tree_add_7_25_groupi_g14099__7098(csa_tree_add_7_25_groupi_n_6973 ,csa_tree_add_7_25_groupi_n_2118 ,csa_tree_add_7_25_groupi_n_1114);
  xnor csa_tree_add_7_25_groupi_g14100__6131(csa_tree_add_7_25_groupi_n_6972 ,csa_tree_add_7_25_groupi_n_6914 ,csa_tree_add_7_25_groupi_n_6863);
  xnor csa_tree_add_7_25_groupi_g14101__1881(csa_tree_add_7_25_groupi_n_6971 ,csa_tree_add_7_25_groupi_n_6913 ,csa_tree_add_7_25_groupi_n_6864);
  xnor csa_tree_add_7_25_groupi_g14102__5115(csa_tree_add_7_25_groupi_n_6970 ,csa_tree_add_7_25_groupi_n_6925 ,in3[17]);
  xnor csa_tree_add_7_25_groupi_g14103__7482(csa_tree_add_7_25_groupi_n_6996 ,csa_tree_add_7_25_groupi_n_6922 ,in3[5]);
  xnor csa_tree_add_7_25_groupi_g14104__4733(csa_tree_add_7_25_groupi_n_6995 ,csa_tree_add_7_25_groupi_n_6921 ,in3[14]);
  xnor csa_tree_add_7_25_groupi_g14105__6161(csa_tree_add_7_25_groupi_n_6994 ,csa_tree_add_7_25_groupi_n_6926 ,in3[2]);
  xnor csa_tree_add_7_25_groupi_g14106__9315(csa_tree_add_7_25_groupi_n_6993 ,csa_tree_add_7_25_groupi_n_6924 ,in3[11]);
  xnor csa_tree_add_7_25_groupi_g14107__9945(csa_tree_add_7_25_groupi_n_6992 ,csa_tree_add_7_25_groupi_n_6923 ,in3[8]);
  xnor csa_tree_add_7_25_groupi_g14108__2883(csa_tree_add_7_25_groupi_n_6991 ,csa_tree_add_7_25_groupi_n_6868 ,csa_tree_add_7_25_groupi_n_6902);
  xnor csa_tree_add_7_25_groupi_g14109__2346(csa_tree_add_7_25_groupi_n_6990 ,csa_tree_add_7_25_groupi_n_6917 ,csa_tree_add_7_25_groupi_n_6822);
  xnor csa_tree_add_7_25_groupi_g14110__1666(csa_tree_add_7_25_groupi_n_6989 ,csa_tree_add_7_25_groupi_n_6916 ,csa_tree_add_7_25_groupi_n_6828);
  xnor csa_tree_add_7_25_groupi_g14111__7410(csa_tree_add_7_25_groupi_n_6987 ,csa_tree_add_7_25_groupi_n_6920 ,csa_tree_add_7_25_groupi_n_6823);
  xnor csa_tree_add_7_25_groupi_g14112__6417(csa_tree_add_7_25_groupi_n_6986 ,csa_tree_add_7_25_groupi_n_6918 ,csa_tree_add_7_25_groupi_n_6826);
  xnor csa_tree_add_7_25_groupi_g14113__5477(csa_tree_add_7_25_groupi_n_6984 ,csa_tree_add_7_25_groupi_n_6866 ,csa_tree_add_7_25_groupi_n_6906);
  xnor csa_tree_add_7_25_groupi_g14114__2398(csa_tree_add_7_25_groupi_n_6982 ,csa_tree_add_7_25_groupi_n_6865 ,csa_tree_add_7_25_groupi_n_6910);
  xnor csa_tree_add_7_25_groupi_g14115__5107(csa_tree_add_7_25_groupi_n_6980 ,csa_tree_add_7_25_groupi_n_6867 ,csa_tree_add_7_25_groupi_n_6909);
  xnor csa_tree_add_7_25_groupi_g14116__6260(csa_tree_add_7_25_groupi_n_6978 ,csa_tree_add_7_25_groupi_n_6919 ,csa_tree_add_7_25_groupi_n_6827);
  xnor csa_tree_add_7_25_groupi_g14117__4319(csa_tree_add_7_25_groupi_n_6976 ,csa_tree_add_7_25_groupi_n_6915 ,csa_tree_add_7_25_groupi_n_6821);
  and csa_tree_add_7_25_groupi_g14118__8428(csa_tree_add_7_25_groupi_n_6968 ,csa_tree_add_7_25_groupi_n_6915 ,csa_tree_add_7_25_groupi_n_6816);
  or csa_tree_add_7_25_groupi_g14119__5526(csa_tree_add_7_25_groupi_n_6967 ,csa_tree_add_7_25_groupi_n_3444 ,csa_tree_add_7_25_groupi_n_6932);
  or csa_tree_add_7_25_groupi_g14120__6783(csa_tree_add_7_25_groupi_n_6966 ,csa_tree_add_7_25_groupi_n_3796 ,csa_tree_add_7_25_groupi_n_6927);
  or csa_tree_add_7_25_groupi_g14121__3680(csa_tree_add_7_25_groupi_n_6965 ,csa_tree_add_7_25_groupi_n_3798 ,csa_tree_add_7_25_groupi_n_6933);
  or csa_tree_add_7_25_groupi_g14122__1617(csa_tree_add_7_25_groupi_n_6964 ,csa_tree_add_7_25_groupi_n_3795 ,csa_tree_add_7_25_groupi_n_6934);
  and csa_tree_add_7_25_groupi_g14123__2802(csa_tree_add_7_25_groupi_n_6963 ,csa_tree_add_7_25_groupi_n_6916 ,csa_tree_add_7_25_groupi_n_6802);
  or csa_tree_add_7_25_groupi_g14124__1705(csa_tree_add_7_25_groupi_n_6962 ,csa_tree_add_7_25_groupi_n_6914 ,csa_tree_add_7_25_groupi_n_6863);
  and csa_tree_add_7_25_groupi_g14125__5122(csa_tree_add_7_25_groupi_n_6961 ,csa_tree_add_7_25_groupi_n_6914 ,csa_tree_add_7_25_groupi_n_6863);
  and csa_tree_add_7_25_groupi_g14126__8246(csa_tree_add_7_25_groupi_n_6960 ,csa_tree_add_7_25_groupi_n_6920 ,csa_tree_add_7_25_groupi_n_6807);
  and csa_tree_add_7_25_groupi_g14127__7098(csa_tree_add_7_25_groupi_n_6959 ,csa_tree_add_7_25_groupi_n_6913 ,csa_tree_add_7_25_groupi_n_6864);
  or csa_tree_add_7_25_groupi_g14128__6131(csa_tree_add_7_25_groupi_n_6958 ,csa_tree_add_7_25_groupi_n_6913 ,csa_tree_add_7_25_groupi_n_6864);
  or csa_tree_add_7_25_groupi_g14129__1881(csa_tree_add_7_25_groupi_n_6957 ,csa_tree_add_7_25_groupi_n_3460 ,csa_tree_add_7_25_groupi_n_6928);
  or csa_tree_add_7_25_groupi_g14130__5115(csa_tree_add_7_25_groupi_n_6969 ,csa_tree_add_7_25_groupi_n_6895 ,csa_tree_add_7_25_groupi_n_6935);
  not csa_tree_add_7_25_groupi_g14131(csa_tree_add_7_25_groupi_n_6955 ,csa_tree_add_7_25_groupi_n_6956);
  not csa_tree_add_7_25_groupi_g14132(csa_tree_add_7_25_groupi_n_6952 ,csa_tree_add_7_25_groupi_n_6953);
  not csa_tree_add_7_25_groupi_g14133(csa_tree_add_7_25_groupi_n_6950 ,csa_tree_add_7_25_groupi_n_6951);
  nor csa_tree_add_7_25_groupi_g14134__7482(csa_tree_add_7_25_groupi_n_6948 ,csa_tree_add_7_25_groupi_n_2189 ,csa_tree_add_7_25_groupi_n_6938);
  nor csa_tree_add_7_25_groupi_g14135__4733(csa_tree_add_7_25_groupi_n_6947 ,csa_tree_add_7_25_groupi_n_2174 ,csa_tree_add_7_25_groupi_n_1123);
  and csa_tree_add_7_25_groupi_g14136__6161(csa_tree_add_7_25_groupi_n_6946 ,csa_tree_add_7_25_groupi_n_6918 ,csa_tree_add_7_25_groupi_n_6796);
  and csa_tree_add_7_25_groupi_g14137__9315(csa_tree_add_7_25_groupi_n_6945 ,csa_tree_add_7_25_groupi_n_6917 ,csa_tree_add_7_25_groupi_n_6792);
  and csa_tree_add_7_25_groupi_g14138__9945(csa_tree_add_7_25_groupi_n_6944 ,csa_tree_add_7_25_groupi_n_6919 ,csa_tree_add_7_25_groupi_n_6799);
  nor csa_tree_add_7_25_groupi_g14139__2883(csa_tree_add_7_25_groupi_n_6943 ,csa_tree_add_7_25_groupi_n_2117 ,csa_tree_add_7_25_groupi_n_1122);
  nor csa_tree_add_7_25_groupi_g14140__2346(csa_tree_add_7_25_groupi_n_6942 ,csa_tree_add_7_25_groupi_n_2096 ,csa_tree_add_7_25_groupi_n_1145);
  nor csa_tree_add_7_25_groupi_g14141__1666(csa_tree_add_7_25_groupi_n_6941 ,csa_tree_add_7_25_groupi_n_2132 ,csa_tree_add_7_25_groupi_n_1123);
  or csa_tree_add_7_25_groupi_g14142__7410(csa_tree_add_7_25_groupi_n_6956 ,csa_tree_add_7_25_groupi_n_6931 ,csa_tree_add_7_25_groupi_n_6883);
  or csa_tree_add_7_25_groupi_g14143__6417(csa_tree_add_7_25_groupi_n_6954 ,csa_tree_add_7_25_groupi_n_6872 ,csa_tree_add_7_25_groupi_n_6929);
  or csa_tree_add_7_25_groupi_g14144__5477(csa_tree_add_7_25_groupi_n_6953 ,csa_tree_add_7_25_groupi_n_6880 ,csa_tree_add_7_25_groupi_n_6937);
  or csa_tree_add_7_25_groupi_g14145__2398(csa_tree_add_7_25_groupi_n_6951 ,csa_tree_add_7_25_groupi_n_6870 ,csa_tree_add_7_25_groupi_n_6930);
  or csa_tree_add_7_25_groupi_g14146__5107(csa_tree_add_7_25_groupi_n_6949 ,csa_tree_add_7_25_groupi_n_2347 ,csa_tree_add_7_25_groupi_n_6936);
  and csa_tree_add_7_25_groupi_g14148__6260(csa_tree_add_7_25_groupi_n_6937 ,csa_tree_add_7_25_groupi_n_6867 ,csa_tree_add_7_25_groupi_n_6876);
  nor csa_tree_add_7_25_groupi_g14149__4319(csa_tree_add_7_25_groupi_n_6936 ,in1[31] ,csa_tree_add_7_25_groupi_n_6900);
  and csa_tree_add_7_25_groupi_g14150__8428(csa_tree_add_7_25_groupi_n_6935 ,csa_tree_add_7_25_groupi_n_6898 ,csa_tree_add_7_25_groupi_n_6894);
  nor csa_tree_add_7_25_groupi_g14151__5526(csa_tree_add_7_25_groupi_n_6934 ,csa_tree_add_7_25_groupi_n_2162 ,csa_tree_add_7_25_groupi_n_1142);
  nor csa_tree_add_7_25_groupi_g14152__6783(csa_tree_add_7_25_groupi_n_6933 ,csa_tree_add_7_25_groupi_n_2108 ,csa_tree_add_7_25_groupi_n_6884);
  nor csa_tree_add_7_25_groupi_g14153__3680(csa_tree_add_7_25_groupi_n_6932 ,csa_tree_add_7_25_groupi_n_2153 ,csa_tree_add_7_25_groupi_n_1142);
  and csa_tree_add_7_25_groupi_g14154__1617(csa_tree_add_7_25_groupi_n_6931 ,csa_tree_add_7_25_groupi_n_6877 ,csa_tree_add_7_25_groupi_n_6865);
  and csa_tree_add_7_25_groupi_g14155__2802(csa_tree_add_7_25_groupi_n_6930 ,csa_tree_add_7_25_groupi_n_6875 ,csa_tree_add_7_25_groupi_n_6866);
  and csa_tree_add_7_25_groupi_g14156__1705(csa_tree_add_7_25_groupi_n_6929 ,csa_tree_add_7_25_groupi_n_6868 ,csa_tree_add_7_25_groupi_n_6871);
  nor csa_tree_add_7_25_groupi_g14157__5122(csa_tree_add_7_25_groupi_n_6928 ,csa_tree_add_7_25_groupi_n_2180 ,csa_tree_add_7_25_groupi_n_6884);
  nor csa_tree_add_7_25_groupi_g14158__8246(csa_tree_add_7_25_groupi_n_6927 ,csa_tree_add_7_25_groupi_n_2192 ,csa_tree_add_7_25_groupi_n_1141);
  nor csa_tree_add_7_25_groupi_g14159__7098(csa_tree_add_7_25_groupi_n_6926 ,csa_tree_add_7_25_groupi_n_3465 ,csa_tree_add_7_25_groupi_n_6869);
  nor csa_tree_add_7_25_groupi_g14160__6131(csa_tree_add_7_25_groupi_n_6925 ,csa_tree_add_7_25_groupi_n_3889 ,csa_tree_add_7_25_groupi_n_6893);
  nor csa_tree_add_7_25_groupi_g14161__1881(csa_tree_add_7_25_groupi_n_6924 ,csa_tree_add_7_25_groupi_n_3905 ,csa_tree_add_7_25_groupi_n_6891);
  nor csa_tree_add_7_25_groupi_g14162__5115(csa_tree_add_7_25_groupi_n_6923 ,csa_tree_add_7_25_groupi_n_3940 ,csa_tree_add_7_25_groupi_n_6889);
  nor csa_tree_add_7_25_groupi_g14163__7482(csa_tree_add_7_25_groupi_n_6922 ,csa_tree_add_7_25_groupi_n_3877 ,csa_tree_add_7_25_groupi_n_6892);
  nor csa_tree_add_7_25_groupi_g14164__4733(csa_tree_add_7_25_groupi_n_6921 ,csa_tree_add_7_25_groupi_n_3832 ,csa_tree_add_7_25_groupi_n_6897);
  or csa_tree_add_7_25_groupi_g14165__6161(csa_tree_add_7_25_groupi_n_6940 ,csa_tree_add_7_25_groupi_n_6729 ,csa_tree_add_7_25_groupi_n_6885);
  or csa_tree_add_7_25_groupi_g14166__9315(csa_tree_add_7_25_groupi_n_6939 ,csa_tree_add_7_25_groupi_n_6730 ,csa_tree_add_7_25_groupi_n_6887);
  or csa_tree_add_7_25_groupi_g14167__9945(csa_tree_add_7_25_groupi_n_6938 ,csa_tree_add_7_25_groupi_n_38 ,csa_tree_add_7_25_groupi_n_6899);
  xnor csa_tree_add_7_25_groupi_g14168__2883(out2[21] ,csa_tree_add_7_25_groupi_n_6819 ,csa_tree_add_7_25_groupi_n_6824);
  xnor csa_tree_add_7_25_groupi_g14169__2346(csa_tree_add_7_25_groupi_n_6911 ,csa_tree_add_7_25_groupi_n_6835 ,csa_tree_add_7_25_groupi_n_6783);
  xnor csa_tree_add_7_25_groupi_g14170__1666(csa_tree_add_7_25_groupi_n_6910 ,csa_tree_add_7_25_groupi_n_6833 ,csa_tree_add_7_25_groupi_n_6755);
  xnor csa_tree_add_7_25_groupi_g14171__7410(csa_tree_add_7_25_groupi_n_6909 ,csa_tree_add_7_25_groupi_n_6831 ,csa_tree_add_7_25_groupi_n_6753);
  xnor csa_tree_add_7_25_groupi_g14172__6417(csa_tree_add_7_25_groupi_n_6908 ,csa_tree_add_7_25_groupi_n_6767 ,csa_tree_add_7_25_groupi_n_6825);
  xnor csa_tree_add_7_25_groupi_g14173__5477(csa_tree_add_7_25_groupi_n_6907 ,csa_tree_add_7_25_groupi_n_6841 ,csa_tree_add_7_25_groupi_n_6788);
  xnor csa_tree_add_7_25_groupi_g14174__2398(csa_tree_add_7_25_groupi_n_6906 ,csa_tree_add_7_25_groupi_n_6845 ,csa_tree_add_7_25_groupi_n_6751);
  xnor csa_tree_add_7_25_groupi_g14175__5107(csa_tree_add_7_25_groupi_n_6905 ,csa_tree_add_7_25_groupi_n_6843 ,csa_tree_add_7_25_groupi_n_6790);
  xnor csa_tree_add_7_25_groupi_g14176__6260(csa_tree_add_7_25_groupi_n_6904 ,csa_tree_add_7_25_groupi_n_6837 ,csa_tree_add_7_25_groupi_n_6786);
  xnor csa_tree_add_7_25_groupi_g14177__4319(csa_tree_add_7_25_groupi_n_6903 ,csa_tree_add_7_25_groupi_n_6791 ,csa_tree_add_7_25_groupi_n_6839);
  xnor csa_tree_add_7_25_groupi_g14178__8428(csa_tree_add_7_25_groupi_n_6902 ,csa_tree_add_7_25_groupi_n_6838 ,csa_tree_add_7_25_groupi_n_6760);
  xnor csa_tree_add_7_25_groupi_g14179__5526(csa_tree_add_7_25_groupi_n_6901 ,csa_tree_add_7_25_groupi_n_6784 ,csa_tree_add_7_25_groupi_n_6846);
  xnor csa_tree_add_7_25_groupi_g14180__6783(csa_tree_add_7_25_groupi_n_6920 ,csa_tree_add_7_25_groupi_n_6849 ,in3[2]);
  xnor csa_tree_add_7_25_groupi_g14181__3680(csa_tree_add_7_25_groupi_n_6919 ,csa_tree_add_7_25_groupi_n_6850 ,in3[14]);
  xnor csa_tree_add_7_25_groupi_g14182__1617(csa_tree_add_7_25_groupi_n_6918 ,csa_tree_add_7_25_groupi_n_6853 ,in3[11]);
  xnor csa_tree_add_7_25_groupi_g14183__2802(csa_tree_add_7_25_groupi_n_6917 ,csa_tree_add_7_25_groupi_n_6854 ,in3[5]);
  xnor csa_tree_add_7_25_groupi_g14184__1705(csa_tree_add_7_25_groupi_n_6916 ,csa_tree_add_7_25_groupi_n_6851 ,in3[17]);
  xnor csa_tree_add_7_25_groupi_g14185__5122(csa_tree_add_7_25_groupi_n_6915 ,csa_tree_add_7_25_groupi_n_6852 ,in3[8]);
  xnor csa_tree_add_7_25_groupi_g14186__8246(csa_tree_add_7_25_groupi_n_6914 ,csa_tree_add_7_25_groupi_n_6847 ,csa_tree_add_7_25_groupi_n_6740);
  xnor csa_tree_add_7_25_groupi_g14187__7098(csa_tree_add_7_25_groupi_n_6913 ,csa_tree_add_7_25_groupi_n_6848 ,csa_tree_add_7_25_groupi_n_6741);
  not csa_tree_add_7_25_groupi_g14188(csa_tree_add_7_25_groupi_n_6900 ,csa_tree_add_7_25_groupi_n_6899);
  or csa_tree_add_7_25_groupi_g14189__6131(csa_tree_add_7_25_groupi_n_6897 ,csa_tree_add_7_25_groupi_n_3790 ,csa_tree_add_7_25_groupi_n_6861);
  or csa_tree_add_7_25_groupi_g14190__1881(csa_tree_add_7_25_groupi_n_6896 ,csa_tree_add_7_25_groupi_n_6784 ,csa_tree_add_7_25_groupi_n_6846);
  and csa_tree_add_7_25_groupi_g14191__5115(csa_tree_add_7_25_groupi_n_6895 ,csa_tree_add_7_25_groupi_n_6791 ,csa_tree_add_7_25_groupi_n_6839);
  or csa_tree_add_7_25_groupi_g14192__7482(csa_tree_add_7_25_groupi_n_6894 ,csa_tree_add_7_25_groupi_n_6791 ,csa_tree_add_7_25_groupi_n_6839);
  or csa_tree_add_7_25_groupi_g14193__4733(csa_tree_add_7_25_groupi_n_6893 ,csa_tree_add_7_25_groupi_n_3792 ,csa_tree_add_7_25_groupi_n_6857);
  or csa_tree_add_7_25_groupi_g14194__6161(csa_tree_add_7_25_groupi_n_6892 ,csa_tree_add_7_25_groupi_n_3791 ,csa_tree_add_7_25_groupi_n_6858);
  or csa_tree_add_7_25_groupi_g14195__9315(csa_tree_add_7_25_groupi_n_6891 ,csa_tree_add_7_25_groupi_n_3794 ,csa_tree_add_7_25_groupi_n_6859);
  and csa_tree_add_7_25_groupi_g14196__9945(csa_tree_add_7_25_groupi_n_6890 ,csa_tree_add_7_25_groupi_n_6784 ,csa_tree_add_7_25_groupi_n_6846);
  or csa_tree_add_7_25_groupi_g14197__2883(csa_tree_add_7_25_groupi_n_6889 ,csa_tree_add_7_25_groupi_n_3793 ,csa_tree_add_7_25_groupi_n_6860);
  nor csa_tree_add_7_25_groupi_g14198__2346(csa_tree_add_7_25_groupi_n_6888 ,csa_tree_add_7_25_groupi_n_6837 ,csa_tree_add_7_25_groupi_n_6785);
  and csa_tree_add_7_25_groupi_g14199__1666(csa_tree_add_7_25_groupi_n_6887 ,csa_tree_add_7_25_groupi_n_6847 ,csa_tree_add_7_25_groupi_n_6736);
  or csa_tree_add_7_25_groupi_g14200__7410(csa_tree_add_7_25_groupi_n_6886 ,csa_tree_add_7_25_groupi_n_6836 ,csa_tree_add_7_25_groupi_n_6786);
  and csa_tree_add_7_25_groupi_g14201__6417(csa_tree_add_7_25_groupi_n_6885 ,csa_tree_add_7_25_groupi_n_6848 ,csa_tree_add_7_25_groupi_n_6728);
  and csa_tree_add_7_25_groupi_g14202__5477(csa_tree_add_7_25_groupi_n_6899 ,csa_tree_add_7_25_groupi_n_2468 ,csa_tree_add_7_25_groupi_n_6862);
  or csa_tree_add_7_25_groupi_g14203__2398(csa_tree_add_7_25_groupi_n_6898 ,csa_tree_add_7_25_groupi_n_6814 ,csa_tree_add_7_25_groupi_n_6855);
  nor csa_tree_add_7_25_groupi_g14204__5107(csa_tree_add_7_25_groupi_n_6883 ,csa_tree_add_7_25_groupi_n_6832 ,csa_tree_add_7_25_groupi_n_6755);
  nor csa_tree_add_7_25_groupi_g14205__6260(csa_tree_add_7_25_groupi_n_6882 ,csa_tree_add_7_25_groupi_n_6843 ,csa_tree_add_7_25_groupi_n_6789);
  or csa_tree_add_7_25_groupi_g14206__4319(csa_tree_add_7_25_groupi_n_6881 ,csa_tree_add_7_25_groupi_n_6842 ,csa_tree_add_7_25_groupi_n_6790);
  nor csa_tree_add_7_25_groupi_g14207__8428(csa_tree_add_7_25_groupi_n_6880 ,csa_tree_add_7_25_groupi_n_6830 ,csa_tree_add_7_25_groupi_n_6753);
  nor csa_tree_add_7_25_groupi_g14208__5526(csa_tree_add_7_25_groupi_n_6879 ,csa_tree_add_7_25_groupi_n_6841 ,csa_tree_add_7_25_groupi_n_6787);
  or csa_tree_add_7_25_groupi_g14209__6783(csa_tree_add_7_25_groupi_n_6878 ,csa_tree_add_7_25_groupi_n_6840 ,csa_tree_add_7_25_groupi_n_6788);
  or csa_tree_add_7_25_groupi_g14210__3680(csa_tree_add_7_25_groupi_n_6877 ,csa_tree_add_7_25_groupi_n_6833 ,csa_tree_add_7_25_groupi_n_6754);
  or csa_tree_add_7_25_groupi_g14211__1617(csa_tree_add_7_25_groupi_n_6876 ,csa_tree_add_7_25_groupi_n_6831 ,csa_tree_add_7_25_groupi_n_6752);
  or csa_tree_add_7_25_groupi_g14212__2802(csa_tree_add_7_25_groupi_n_6875 ,csa_tree_add_7_25_groupi_n_6845 ,csa_tree_add_7_25_groupi_n_6750);
  nor csa_tree_add_7_25_groupi_g14213__1705(csa_tree_add_7_25_groupi_n_6874 ,csa_tree_add_7_25_groupi_n_6835 ,csa_tree_add_7_25_groupi_n_6782);
  or csa_tree_add_7_25_groupi_g14214__5122(csa_tree_add_7_25_groupi_n_6873 ,csa_tree_add_7_25_groupi_n_6834 ,csa_tree_add_7_25_groupi_n_6783);
  and csa_tree_add_7_25_groupi_g14215__8246(csa_tree_add_7_25_groupi_n_6872 ,csa_tree_add_7_25_groupi_n_6838 ,csa_tree_add_7_25_groupi_n_6760);
  or csa_tree_add_7_25_groupi_g14216__7098(csa_tree_add_7_25_groupi_n_6871 ,csa_tree_add_7_25_groupi_n_6838 ,csa_tree_add_7_25_groupi_n_6760);
  nor csa_tree_add_7_25_groupi_g14217__6131(csa_tree_add_7_25_groupi_n_6870 ,csa_tree_add_7_25_groupi_n_6844 ,csa_tree_add_7_25_groupi_n_6751);
  or csa_tree_add_7_25_groupi_g14218__1881(csa_tree_add_7_25_groupi_n_6869 ,csa_tree_add_7_25_groupi_n_3442 ,csa_tree_add_7_25_groupi_n_6856);
  xnor csa_tree_add_7_25_groupi_g14219__5115(csa_tree_add_7_25_groupi_n_6884 ,csa_tree_add_7_25_groupi_n_6820 ,csa_tree_add_7_25_groupi_n_2597);
  or csa_tree_add_7_25_groupi_g14220__7482(csa_tree_add_7_25_groupi_n_6862 ,csa_tree_add_7_25_groupi_n_2464 ,csa_tree_add_7_25_groupi_n_6820);
  nor csa_tree_add_7_25_groupi_g14221__4733(csa_tree_add_7_25_groupi_n_6861 ,csa_tree_add_7_25_groupi_n_2750 ,csa_tree_add_7_25_groupi_n_1131);
  nor csa_tree_add_7_25_groupi_g14222__6161(csa_tree_add_7_25_groupi_n_6860 ,csa_tree_add_7_25_groupi_n_2742 ,csa_tree_add_7_25_groupi_n_1131);
  nor csa_tree_add_7_25_groupi_g14223__9315(csa_tree_add_7_25_groupi_n_6859 ,csa_tree_add_7_25_groupi_n_2738 ,csa_tree_add_7_25_groupi_n_6806);
  nor csa_tree_add_7_25_groupi_g14224__9945(csa_tree_add_7_25_groupi_n_6858 ,csa_tree_add_7_25_groupi_n_2746 ,csa_tree_add_7_25_groupi_n_1130);
  nor csa_tree_add_7_25_groupi_g14225__2883(csa_tree_add_7_25_groupi_n_6857 ,csa_tree_add_7_25_groupi_n_2073 ,csa_tree_add_7_25_groupi_n_1133);
  nor csa_tree_add_7_25_groupi_g14226__2346(csa_tree_add_7_25_groupi_n_6856 ,csa_tree_add_7_25_groupi_n_2836 ,csa_tree_add_7_25_groupi_n_1133);
  and csa_tree_add_7_25_groupi_g14227__1666(csa_tree_add_7_25_groupi_n_6855 ,csa_tree_add_7_25_groupi_n_6819 ,csa_tree_add_7_25_groupi_n_6812);
  nor csa_tree_add_7_25_groupi_g14228__7410(csa_tree_add_7_25_groupi_n_6854 ,csa_tree_add_7_25_groupi_n_4011 ,csa_tree_add_7_25_groupi_n_6815);
  nor csa_tree_add_7_25_groupi_g14229__6417(csa_tree_add_7_25_groupi_n_6853 ,csa_tree_add_7_25_groupi_n_3897 ,csa_tree_add_7_25_groupi_n_6818);
  nor csa_tree_add_7_25_groupi_g14230__5477(csa_tree_add_7_25_groupi_n_6852 ,csa_tree_add_7_25_groupi_n_3878 ,csa_tree_add_7_25_groupi_n_6798);
  nor csa_tree_add_7_25_groupi_g14231__2398(csa_tree_add_7_25_groupi_n_6851 ,csa_tree_add_7_25_groupi_n_4016 ,csa_tree_add_7_25_groupi_n_6811);
  nor csa_tree_add_7_25_groupi_g14232__5107(csa_tree_add_7_25_groupi_n_6850 ,csa_tree_add_7_25_groupi_n_3818 ,csa_tree_add_7_25_groupi_n_6804);
  nor csa_tree_add_7_25_groupi_g14233__6260(csa_tree_add_7_25_groupi_n_6849 ,csa_tree_add_7_25_groupi_n_3479 ,csa_tree_add_7_25_groupi_n_6803);
  or csa_tree_add_7_25_groupi_g14234__4319(csa_tree_add_7_25_groupi_n_6868 ,csa_tree_add_7_25_groupi_n_6662 ,csa_tree_add_7_25_groupi_n_6809);
  or csa_tree_add_7_25_groupi_g14235__8428(csa_tree_add_7_25_groupi_n_6867 ,csa_tree_add_7_25_groupi_n_6640 ,csa_tree_add_7_25_groupi_n_6805);
  or csa_tree_add_7_25_groupi_g14236__5526(csa_tree_add_7_25_groupi_n_6866 ,csa_tree_add_7_25_groupi_n_6635 ,csa_tree_add_7_25_groupi_n_6794);
  or csa_tree_add_7_25_groupi_g14237__6783(csa_tree_add_7_25_groupi_n_6865 ,csa_tree_add_7_25_groupi_n_6646 ,csa_tree_add_7_25_groupi_n_6795);
  or csa_tree_add_7_25_groupi_g14238__3680(csa_tree_add_7_25_groupi_n_6864 ,csa_tree_add_7_25_groupi_n_6652 ,csa_tree_add_7_25_groupi_n_6813);
  or csa_tree_add_7_25_groupi_g14239__1617(csa_tree_add_7_25_groupi_n_6863 ,csa_tree_add_7_25_groupi_n_6657 ,csa_tree_add_7_25_groupi_n_6810);
  not csa_tree_add_7_25_groupi_g14240(csa_tree_add_7_25_groupi_n_6844 ,csa_tree_add_7_25_groupi_n_6845);
  not csa_tree_add_7_25_groupi_g14241(csa_tree_add_7_25_groupi_n_6842 ,csa_tree_add_7_25_groupi_n_6843);
  not csa_tree_add_7_25_groupi_g14242(csa_tree_add_7_25_groupi_n_6840 ,csa_tree_add_7_25_groupi_n_6841);
  not csa_tree_add_7_25_groupi_g14243(csa_tree_add_7_25_groupi_n_6837 ,csa_tree_add_7_25_groupi_n_6836);
  not csa_tree_add_7_25_groupi_g14244(csa_tree_add_7_25_groupi_n_6834 ,csa_tree_add_7_25_groupi_n_6835);
  not csa_tree_add_7_25_groupi_g14245(csa_tree_add_7_25_groupi_n_6832 ,csa_tree_add_7_25_groupi_n_6833);
  not csa_tree_add_7_25_groupi_g14246(csa_tree_add_7_25_groupi_n_6830 ,csa_tree_add_7_25_groupi_n_6831);
  xnor csa_tree_add_7_25_groupi_g14247__2802(out2[20] ,csa_tree_add_7_25_groupi_n_6737 ,csa_tree_add_7_25_groupi_n_6739);
  xnor csa_tree_add_7_25_groupi_g14248__1705(csa_tree_add_7_25_groupi_n_6828 ,csa_tree_add_7_25_groupi_n_6720 ,csa_tree_add_7_25_groupi_n_6745);
  xnor csa_tree_add_7_25_groupi_g14249__5122(csa_tree_add_7_25_groupi_n_6827 ,csa_tree_add_7_25_groupi_n_6747 ,csa_tree_add_7_25_groupi_n_6724);
  xnor csa_tree_add_7_25_groupi_g14250__8246(csa_tree_add_7_25_groupi_n_6826 ,csa_tree_add_7_25_groupi_n_6722 ,csa_tree_add_7_25_groupi_n_6749);
  xnor csa_tree_add_7_25_groupi_g14251__7098(csa_tree_add_7_25_groupi_n_6825 ,csa_tree_add_7_25_groupi_n_6742 ,csa_tree_add_7_25_groupi_n_6666);
  xnor csa_tree_add_7_25_groupi_g14252__6131(csa_tree_add_7_25_groupi_n_6824 ,csa_tree_add_7_25_groupi_n_6707 ,csa_tree_add_7_25_groupi_n_6758);
  xnor csa_tree_add_7_25_groupi_g14253__1881(csa_tree_add_7_25_groupi_n_6823 ,csa_tree_add_7_25_groupi_n_6709 ,csa_tree_add_7_25_groupi_n_6756);
  xnor csa_tree_add_7_25_groupi_g14254__5115(csa_tree_add_7_25_groupi_n_6822 ,csa_tree_add_7_25_groupi_n_6708 ,csa_tree_add_7_25_groupi_n_6759);
  xnor csa_tree_add_7_25_groupi_g14255__7482(csa_tree_add_7_25_groupi_n_6821 ,csa_tree_add_7_25_groupi_n_6757 ,csa_tree_add_7_25_groupi_n_6725);
  xnor csa_tree_add_7_25_groupi_g14256__4733(csa_tree_add_7_25_groupi_n_6848 ,csa_tree_add_7_25_groupi_n_6770 ,in3[5]);
  xnor csa_tree_add_7_25_groupi_g14257__6161(csa_tree_add_7_25_groupi_n_6847 ,csa_tree_add_7_25_groupi_n_6771 ,in3[2]);
  xnor csa_tree_add_7_25_groupi_g14258__9315(csa_tree_add_7_25_groupi_n_6846 ,csa_tree_add_7_25_groupi_n_6765 ,csa_tree_add_7_25_groupi_n_6676);
  xnor csa_tree_add_7_25_groupi_g14259__9945(csa_tree_add_7_25_groupi_n_6845 ,csa_tree_add_7_25_groupi_n_6772 ,in3[11]);
  xnor csa_tree_add_7_25_groupi_g14260__2883(csa_tree_add_7_25_groupi_n_6843 ,csa_tree_add_7_25_groupi_n_6766 ,csa_tree_add_7_25_groupi_n_6670);
  xnor csa_tree_add_7_25_groupi_g14261__2346(csa_tree_add_7_25_groupi_n_6841 ,csa_tree_add_7_25_groupi_n_6763 ,csa_tree_add_7_25_groupi_n_6667);
  xnor csa_tree_add_7_25_groupi_g14262__1666(csa_tree_add_7_25_groupi_n_6839 ,csa_tree_add_7_25_groupi_n_6764 ,csa_tree_add_7_25_groupi_n_6674);
  xnor csa_tree_add_7_25_groupi_g14263__7410(csa_tree_add_7_25_groupi_n_6838 ,csa_tree_add_7_25_groupi_n_6773 ,in3[8]);
  xnor csa_tree_add_7_25_groupi_g14264__6417(csa_tree_add_7_25_groupi_n_6836 ,csa_tree_add_7_25_groupi_n_6761 ,csa_tree_add_7_25_groupi_n_6675);
  xnor csa_tree_add_7_25_groupi_g14265__5477(csa_tree_add_7_25_groupi_n_6835 ,csa_tree_add_7_25_groupi_n_6762 ,csa_tree_add_7_25_groupi_n_6673);
  xnor csa_tree_add_7_25_groupi_g14266__2398(csa_tree_add_7_25_groupi_n_6833 ,csa_tree_add_7_25_groupi_n_6768 ,in3[14]);
  xnor csa_tree_add_7_25_groupi_g14267__5107(csa_tree_add_7_25_groupi_n_6831 ,csa_tree_add_7_25_groupi_n_6769 ,in3[17]);
  or csa_tree_add_7_25_groupi_g14268__6260(csa_tree_add_7_25_groupi_n_6818 ,csa_tree_add_7_25_groupi_n_3789 ,csa_tree_add_7_25_groupi_n_6779);
  and csa_tree_add_7_25_groupi_g14269__4319(csa_tree_add_7_25_groupi_n_6817 ,csa_tree_add_7_25_groupi_n_6757 ,csa_tree_add_7_25_groupi_n_6725);
  or csa_tree_add_7_25_groupi_g14270__8428(csa_tree_add_7_25_groupi_n_6816 ,csa_tree_add_7_25_groupi_n_6757 ,csa_tree_add_7_25_groupi_n_6725);
  or csa_tree_add_7_25_groupi_g14271__5526(csa_tree_add_7_25_groupi_n_6815 ,csa_tree_add_7_25_groupi_n_3451 ,csa_tree_add_7_25_groupi_n_6777);
  and csa_tree_add_7_25_groupi_g14272__6783(csa_tree_add_7_25_groupi_n_6814 ,csa_tree_add_7_25_groupi_n_6707 ,csa_tree_add_7_25_groupi_n_6758);
  and csa_tree_add_7_25_groupi_g14273__3680(csa_tree_add_7_25_groupi_n_6813 ,csa_tree_add_7_25_groupi_n_6765 ,csa_tree_add_7_25_groupi_n_6651);
  or csa_tree_add_7_25_groupi_g14274__1617(csa_tree_add_7_25_groupi_n_6812 ,csa_tree_add_7_25_groupi_n_6707 ,csa_tree_add_7_25_groupi_n_6758);
  or csa_tree_add_7_25_groupi_g14275__2802(csa_tree_add_7_25_groupi_n_6811 ,csa_tree_add_7_25_groupi_n_3417 ,csa_tree_add_7_25_groupi_n_6776);
  and csa_tree_add_7_25_groupi_g14276__1705(csa_tree_add_7_25_groupi_n_6810 ,csa_tree_add_7_25_groupi_n_6764 ,csa_tree_add_7_25_groupi_n_6656);
  and csa_tree_add_7_25_groupi_g14277__5122(csa_tree_add_7_25_groupi_n_6809 ,csa_tree_add_7_25_groupi_n_6761 ,csa_tree_add_7_25_groupi_n_6654);
  and csa_tree_add_7_25_groupi_g14278__8246(csa_tree_add_7_25_groupi_n_6808 ,csa_tree_add_7_25_groupi_n_6709 ,csa_tree_add_7_25_groupi_n_6756);
  or csa_tree_add_7_25_groupi_g14279__7098(csa_tree_add_7_25_groupi_n_6807 ,csa_tree_add_7_25_groupi_n_6709 ,csa_tree_add_7_25_groupi_n_6756);
  and csa_tree_add_7_25_groupi_g14280__6131(csa_tree_add_7_25_groupi_n_6820 ,csa_tree_add_7_25_groupi_n_2432 ,csa_tree_add_7_25_groupi_n_6780);
  or csa_tree_add_7_25_groupi_g14281__1881(csa_tree_add_7_25_groupi_n_6819 ,csa_tree_add_7_25_groupi_n_6774 ,csa_tree_add_7_25_groupi_n_6734);
  and csa_tree_add_7_25_groupi_g14282__5115(csa_tree_add_7_25_groupi_n_6805 ,csa_tree_add_7_25_groupi_n_6766 ,csa_tree_add_7_25_groupi_n_6643);
  or csa_tree_add_7_25_groupi_g14283__7482(csa_tree_add_7_25_groupi_n_6804 ,csa_tree_add_7_25_groupi_n_3785 ,csa_tree_add_7_25_groupi_n_6778);
  or csa_tree_add_7_25_groupi_g14284__4733(csa_tree_add_7_25_groupi_n_6803 ,csa_tree_add_7_25_groupi_n_3429 ,csa_tree_add_7_25_groupi_n_6775);
  or csa_tree_add_7_25_groupi_g14285__6161(csa_tree_add_7_25_groupi_n_6802 ,csa_tree_add_7_25_groupi_n_6720 ,csa_tree_add_7_25_groupi_n_6744);
  nor csa_tree_add_7_25_groupi_g14286__9315(csa_tree_add_7_25_groupi_n_6801 ,csa_tree_add_7_25_groupi_n_6719 ,csa_tree_add_7_25_groupi_n_6745);
  nor csa_tree_add_7_25_groupi_g14287__9945(csa_tree_add_7_25_groupi_n_6800 ,csa_tree_add_7_25_groupi_n_6747 ,csa_tree_add_7_25_groupi_n_6723);
  or csa_tree_add_7_25_groupi_g14288__2883(csa_tree_add_7_25_groupi_n_6799 ,csa_tree_add_7_25_groupi_n_6746 ,csa_tree_add_7_25_groupi_n_6724);
  or csa_tree_add_7_25_groupi_g14289__2346(csa_tree_add_7_25_groupi_n_6798 ,csa_tree_add_7_25_groupi_n_3786 ,csa_tree_add_7_25_groupi_n_6781);
  nor csa_tree_add_7_25_groupi_g14290__1666(csa_tree_add_7_25_groupi_n_6797 ,csa_tree_add_7_25_groupi_n_6721 ,csa_tree_add_7_25_groupi_n_6749);
  or csa_tree_add_7_25_groupi_g14291__7410(csa_tree_add_7_25_groupi_n_6796 ,csa_tree_add_7_25_groupi_n_6722 ,csa_tree_add_7_25_groupi_n_6748);
  and csa_tree_add_7_25_groupi_g14292__6417(csa_tree_add_7_25_groupi_n_6795 ,csa_tree_add_7_25_groupi_n_6763 ,csa_tree_add_7_25_groupi_n_6636);
  and csa_tree_add_7_25_groupi_g14293__5477(csa_tree_add_7_25_groupi_n_6794 ,csa_tree_add_7_25_groupi_n_6762 ,csa_tree_add_7_25_groupi_n_6634);
  and csa_tree_add_7_25_groupi_g14294__2398(csa_tree_add_7_25_groupi_n_6793 ,csa_tree_add_7_25_groupi_n_6708 ,csa_tree_add_7_25_groupi_n_6759);
  or csa_tree_add_7_25_groupi_g14295__5107(csa_tree_add_7_25_groupi_n_6792 ,csa_tree_add_7_25_groupi_n_6708 ,csa_tree_add_7_25_groupi_n_6759);
  xnor csa_tree_add_7_25_groupi_g14296__6260(csa_tree_add_7_25_groupi_n_6806 ,csa_tree_add_7_25_groupi_n_6738 ,csa_tree_add_7_25_groupi_n_2559);
  not csa_tree_add_7_25_groupi_g14297(csa_tree_add_7_25_groupi_n_6789 ,csa_tree_add_7_25_groupi_n_6790);
  not csa_tree_add_7_25_groupi_g14298(csa_tree_add_7_25_groupi_n_6787 ,csa_tree_add_7_25_groupi_n_6788);
  not csa_tree_add_7_25_groupi_g14299(csa_tree_add_7_25_groupi_n_6785 ,csa_tree_add_7_25_groupi_n_6786);
  not csa_tree_add_7_25_groupi_g14300(csa_tree_add_7_25_groupi_n_6782 ,csa_tree_add_7_25_groupi_n_6783);
  nor csa_tree_add_7_25_groupi_g14301__4319(csa_tree_add_7_25_groupi_n_6781 ,csa_tree_add_7_25_groupi_n_2109 ,csa_tree_add_7_25_groupi_n_1128);
  or csa_tree_add_7_25_groupi_g14302__8428(csa_tree_add_7_25_groupi_n_6780 ,csa_tree_add_7_25_groupi_n_2489 ,csa_tree_add_7_25_groupi_n_6738);
  nor csa_tree_add_7_25_groupi_g14303__5526(csa_tree_add_7_25_groupi_n_6779 ,csa_tree_add_7_25_groupi_n_2163 ,csa_tree_add_7_25_groupi_n_1128);
  nor csa_tree_add_7_25_groupi_g14304__6783(csa_tree_add_7_25_groupi_n_6778 ,csa_tree_add_7_25_groupi_n_2154 ,csa_tree_add_7_25_groupi_n_6718);
  nor csa_tree_add_7_25_groupi_g14305__3680(csa_tree_add_7_25_groupi_n_6777 ,csa_tree_add_7_25_groupi_n_2193 ,csa_tree_add_7_25_groupi_n_1127);
  nor csa_tree_add_7_25_groupi_g14306__1617(csa_tree_add_7_25_groupi_n_6776 ,csa_tree_add_7_25_groupi_n_2072 ,csa_tree_add_7_25_groupi_n_1139);
  nor csa_tree_add_7_25_groupi_g14307__2802(csa_tree_add_7_25_groupi_n_6775 ,csa_tree_add_7_25_groupi_n_2181 ,csa_tree_add_7_25_groupi_n_1139);
  and csa_tree_add_7_25_groupi_g14308__1705(csa_tree_add_7_25_groupi_n_6774 ,csa_tree_add_7_25_groupi_n_6737 ,csa_tree_add_7_25_groupi_n_6735);
  nor csa_tree_add_7_25_groupi_g14309__5122(csa_tree_add_7_25_groupi_n_6773 ,csa_tree_add_7_25_groupi_n_3815 ,csa_tree_add_7_25_groupi_n_6717);
  nor csa_tree_add_7_25_groupi_g14310__8246(csa_tree_add_7_25_groupi_n_6772 ,csa_tree_add_7_25_groupi_n_3816 ,csa_tree_add_7_25_groupi_n_6715);
  nor csa_tree_add_7_25_groupi_g14311__7098(csa_tree_add_7_25_groupi_n_6771 ,csa_tree_add_7_25_groupi_n_3468 ,csa_tree_add_7_25_groupi_n_6714);
  nor csa_tree_add_7_25_groupi_g14312__6131(csa_tree_add_7_25_groupi_n_6770 ,csa_tree_add_7_25_groupi_n_4008 ,csa_tree_add_7_25_groupi_n_6733);
  nor csa_tree_add_7_25_groupi_g14313__1881(csa_tree_add_7_25_groupi_n_6769 ,csa_tree_add_7_25_groupi_n_3850 ,csa_tree_add_7_25_groupi_n_6726);
  nor csa_tree_add_7_25_groupi_g14314__5115(csa_tree_add_7_25_groupi_n_6768 ,csa_tree_add_7_25_groupi_n_3922 ,csa_tree_add_7_25_groupi_n_6716);
  or csa_tree_add_7_25_groupi_g14315__7482(csa_tree_add_7_25_groupi_n_6767 ,csa_tree_add_7_25_groupi_n_6555 ,csa_tree_add_7_25_groupi_n_6713);
  or csa_tree_add_7_25_groupi_g14316__4733(csa_tree_add_7_25_groupi_n_6791 ,csa_tree_add_7_25_groupi_n_6568 ,csa_tree_add_7_25_groupi_n_6732);
  or csa_tree_add_7_25_groupi_g14317__6161(csa_tree_add_7_25_groupi_n_6790 ,csa_tree_add_7_25_groupi_n_6551 ,csa_tree_add_7_25_groupi_n_6710);
  or csa_tree_add_7_25_groupi_g14318__9315(csa_tree_add_7_25_groupi_n_6788 ,csa_tree_add_7_25_groupi_n_6549 ,csa_tree_add_7_25_groupi_n_6711);
  or csa_tree_add_7_25_groupi_g14319__9945(csa_tree_add_7_25_groupi_n_6786 ,csa_tree_add_7_25_groupi_n_6545 ,csa_tree_add_7_25_groupi_n_6712);
  or csa_tree_add_7_25_groupi_g14320__2883(csa_tree_add_7_25_groupi_n_6784 ,csa_tree_add_7_25_groupi_n_6561 ,csa_tree_add_7_25_groupi_n_6727);
  or csa_tree_add_7_25_groupi_g14321__2346(csa_tree_add_7_25_groupi_n_6783 ,csa_tree_add_7_25_groupi_n_6572 ,csa_tree_add_7_25_groupi_n_6731);
  not csa_tree_add_7_25_groupi_g14322(csa_tree_add_7_25_groupi_n_6754 ,csa_tree_add_7_25_groupi_n_6755);
  not csa_tree_add_7_25_groupi_g14323(csa_tree_add_7_25_groupi_n_6752 ,csa_tree_add_7_25_groupi_n_6753);
  not csa_tree_add_7_25_groupi_g14324(csa_tree_add_7_25_groupi_n_6750 ,csa_tree_add_7_25_groupi_n_6751);
  not csa_tree_add_7_25_groupi_g14325(csa_tree_add_7_25_groupi_n_6748 ,csa_tree_add_7_25_groupi_n_6749);
  not csa_tree_add_7_25_groupi_g14326(csa_tree_add_7_25_groupi_n_6746 ,csa_tree_add_7_25_groupi_n_6747);
  not csa_tree_add_7_25_groupi_g14327(csa_tree_add_7_25_groupi_n_6744 ,csa_tree_add_7_25_groupi_n_6745);
  xnor csa_tree_add_7_25_groupi_g14328__1666(out2[19] ,csa_tree_add_7_25_groupi_n_6664 ,csa_tree_add_7_25_groupi_n_6665);
  xnor csa_tree_add_7_25_groupi_g14329__7410(csa_tree_add_7_25_groupi_n_6742 ,csa_tree_add_7_25_groupi_n_6694 ,in3[20]);
  xnor csa_tree_add_7_25_groupi_g14330__6417(csa_tree_add_7_25_groupi_n_6741 ,csa_tree_add_7_25_groupi_n_6679 ,csa_tree_add_7_25_groupi_n_6624);
  xnor csa_tree_add_7_25_groupi_g14331__5477(csa_tree_add_7_25_groupi_n_6740 ,csa_tree_add_7_25_groupi_n_6678 ,csa_tree_add_7_25_groupi_n_6625);
  xnor csa_tree_add_7_25_groupi_g14332__2398(csa_tree_add_7_25_groupi_n_6739 ,csa_tree_add_7_25_groupi_n_6680 ,csa_tree_add_7_25_groupi_n_6623);
  xnor csa_tree_add_7_25_groupi_g14333__5107(csa_tree_add_7_25_groupi_n_6766 ,csa_tree_add_7_25_groupi_n_6693 ,in3[17]);
  xnor csa_tree_add_7_25_groupi_g14334__6260(csa_tree_add_7_25_groupi_n_6765 ,csa_tree_add_7_25_groupi_n_6691 ,in3[5]);
  xnor csa_tree_add_7_25_groupi_g14335__4319(csa_tree_add_7_25_groupi_n_6764 ,csa_tree_add_7_25_groupi_n_6688 ,in3[2]);
  xnor csa_tree_add_7_25_groupi_g14336__8428(csa_tree_add_7_25_groupi_n_6763 ,csa_tree_add_7_25_groupi_n_6692 ,in3[14]);
  xnor csa_tree_add_7_25_groupi_g14337__5526(csa_tree_add_7_25_groupi_n_6762 ,csa_tree_add_7_25_groupi_n_6689 ,in3[11]);
  xnor csa_tree_add_7_25_groupi_g14338__6783(csa_tree_add_7_25_groupi_n_6761 ,csa_tree_add_7_25_groupi_n_6690 ,in3[8]);
  xnor csa_tree_add_7_25_groupi_g14339__3680(csa_tree_add_7_25_groupi_n_6760 ,csa_tree_add_7_25_groupi_n_6626 ,csa_tree_add_7_25_groupi_n_6671);
  xnor csa_tree_add_7_25_groupi_g14340__1617(csa_tree_add_7_25_groupi_n_6759 ,csa_tree_add_7_25_groupi_n_6686 ,csa_tree_add_7_25_groupi_n_6578);
  xnor csa_tree_add_7_25_groupi_g14341__2802(csa_tree_add_7_25_groupi_n_6758 ,csa_tree_add_7_25_groupi_n_6683 ,csa_tree_add_7_25_groupi_n_6580);
  xnor csa_tree_add_7_25_groupi_g14342__1705(csa_tree_add_7_25_groupi_n_6757 ,csa_tree_add_7_25_groupi_n_6685 ,csa_tree_add_7_25_groupi_n_6585);
  xnor csa_tree_add_7_25_groupi_g14343__5122(csa_tree_add_7_25_groupi_n_6756 ,csa_tree_add_7_25_groupi_n_6681 ,csa_tree_add_7_25_groupi_n_6579);
  xnor csa_tree_add_7_25_groupi_g14344__8246(csa_tree_add_7_25_groupi_n_6755 ,csa_tree_add_7_25_groupi_n_6628 ,csa_tree_add_7_25_groupi_n_6669);
  xnor csa_tree_add_7_25_groupi_g14345__7098(csa_tree_add_7_25_groupi_n_6753 ,csa_tree_add_7_25_groupi_n_6629 ,csa_tree_add_7_25_groupi_n_6668);
  xnor csa_tree_add_7_25_groupi_g14346__6131(csa_tree_add_7_25_groupi_n_6751 ,csa_tree_add_7_25_groupi_n_6627 ,csa_tree_add_7_25_groupi_n_6672);
  xnor csa_tree_add_7_25_groupi_g14347__1881(csa_tree_add_7_25_groupi_n_6749 ,csa_tree_add_7_25_groupi_n_6684 ,csa_tree_add_7_25_groupi_n_6583);
  xnor csa_tree_add_7_25_groupi_g14348__5115(csa_tree_add_7_25_groupi_n_6747 ,csa_tree_add_7_25_groupi_n_6687 ,csa_tree_add_7_25_groupi_n_6584);
  xnor csa_tree_add_7_25_groupi_g14349__7482(csa_tree_add_7_25_groupi_n_6745 ,csa_tree_add_7_25_groupi_n_6682 ,csa_tree_add_7_25_groupi_n_6577);
  or csa_tree_add_7_25_groupi_g14350__4733(csa_tree_add_7_25_groupi_n_6736 ,csa_tree_add_7_25_groupi_n_6678 ,csa_tree_add_7_25_groupi_n_6625);
  or csa_tree_add_7_25_groupi_g14351__6161(csa_tree_add_7_25_groupi_n_6735 ,csa_tree_add_7_25_groupi_n_6680 ,csa_tree_add_7_25_groupi_n_6623);
  and csa_tree_add_7_25_groupi_g14352__9315(csa_tree_add_7_25_groupi_n_6734 ,csa_tree_add_7_25_groupi_n_6680 ,csa_tree_add_7_25_groupi_n_6623);
  or csa_tree_add_7_25_groupi_g14353__9945(csa_tree_add_7_25_groupi_n_6733 ,csa_tree_add_7_25_groupi_n_3446 ,csa_tree_add_7_25_groupi_n_6702);
  and csa_tree_add_7_25_groupi_g14354__2883(csa_tree_add_7_25_groupi_n_6732 ,csa_tree_add_7_25_groupi_n_6683 ,csa_tree_add_7_25_groupi_n_6567);
  and csa_tree_add_7_25_groupi_g14355__2346(csa_tree_add_7_25_groupi_n_6731 ,csa_tree_add_7_25_groupi_n_6685 ,csa_tree_add_7_25_groupi_n_6573);
  and csa_tree_add_7_25_groupi_g14356__1666(csa_tree_add_7_25_groupi_n_6730 ,csa_tree_add_7_25_groupi_n_6678 ,csa_tree_add_7_25_groupi_n_6625);
  and csa_tree_add_7_25_groupi_g14357__7410(csa_tree_add_7_25_groupi_n_6729 ,csa_tree_add_7_25_groupi_n_6679 ,csa_tree_add_7_25_groupi_n_6624);
  or csa_tree_add_7_25_groupi_g14358__6417(csa_tree_add_7_25_groupi_n_6728 ,csa_tree_add_7_25_groupi_n_6679 ,csa_tree_add_7_25_groupi_n_6624);
  and csa_tree_add_7_25_groupi_g14359__5477(csa_tree_add_7_25_groupi_n_6727 ,csa_tree_add_7_25_groupi_n_6681 ,csa_tree_add_7_25_groupi_n_6570);
  or csa_tree_add_7_25_groupi_g14360__2398(csa_tree_add_7_25_groupi_n_6726 ,csa_tree_add_7_25_groupi_n_3780 ,csa_tree_add_7_25_groupi_n_6701);
  and csa_tree_add_7_25_groupi_g14361__5107(csa_tree_add_7_25_groupi_n_6738 ,csa_tree_add_7_25_groupi_n_2461 ,csa_tree_add_7_25_groupi_n_6697);
  or csa_tree_add_7_25_groupi_g14362__6260(csa_tree_add_7_25_groupi_n_6737 ,csa_tree_add_7_25_groupi_n_6699 ,csa_tree_add_7_25_groupi_n_6661);
  not csa_tree_add_7_25_groupi_g14363(csa_tree_add_7_25_groupi_n_6723 ,csa_tree_add_7_25_groupi_n_6724);
  not csa_tree_add_7_25_groupi_g14364(csa_tree_add_7_25_groupi_n_6721 ,csa_tree_add_7_25_groupi_n_6722);
  not csa_tree_add_7_25_groupi_g14365(csa_tree_add_7_25_groupi_n_6719 ,csa_tree_add_7_25_groupi_n_6720);
  or csa_tree_add_7_25_groupi_g14366__4319(csa_tree_add_7_25_groupi_n_6717 ,csa_tree_add_7_25_groupi_n_3784 ,csa_tree_add_7_25_groupi_n_6703);
  or csa_tree_add_7_25_groupi_g14367__8428(csa_tree_add_7_25_groupi_n_6716 ,csa_tree_add_7_25_groupi_n_3781 ,csa_tree_add_7_25_groupi_n_6704);
  or csa_tree_add_7_25_groupi_g14368__5526(csa_tree_add_7_25_groupi_n_6715 ,csa_tree_add_7_25_groupi_n_3783 ,csa_tree_add_7_25_groupi_n_6705);
  or csa_tree_add_7_25_groupi_g14369__6783(csa_tree_add_7_25_groupi_n_6714 ,csa_tree_add_7_25_groupi_n_3415 ,csa_tree_add_7_25_groupi_n_6700);
  and csa_tree_add_7_25_groupi_g14370__3680(csa_tree_add_7_25_groupi_n_6713 ,csa_tree_add_7_25_groupi_n_6682 ,csa_tree_add_7_25_groupi_n_6554);
  and csa_tree_add_7_25_groupi_g14371__1617(csa_tree_add_7_25_groupi_n_6712 ,csa_tree_add_7_25_groupi_n_6686 ,csa_tree_add_7_25_groupi_n_6544);
  and csa_tree_add_7_25_groupi_g14372__2802(csa_tree_add_7_25_groupi_n_6711 ,csa_tree_add_7_25_groupi_n_6684 ,csa_tree_add_7_25_groupi_n_6548);
  and csa_tree_add_7_25_groupi_g14373__1705(csa_tree_add_7_25_groupi_n_6710 ,csa_tree_add_7_25_groupi_n_6687 ,csa_tree_add_7_25_groupi_n_6550);
  or csa_tree_add_7_25_groupi_g14374__5122(csa_tree_add_7_25_groupi_n_6725 ,csa_tree_add_7_25_groupi_n_6698 ,csa_tree_add_7_25_groupi_n_6630);
  or csa_tree_add_7_25_groupi_g14375__8246(csa_tree_add_7_25_groupi_n_6724 ,csa_tree_add_7_25_groupi_n_6696 ,csa_tree_add_7_25_groupi_n_6638);
  or csa_tree_add_7_25_groupi_g14376__7098(csa_tree_add_7_25_groupi_n_6722 ,csa_tree_add_7_25_groupi_n_6633 ,csa_tree_add_7_25_groupi_n_6695);
  or csa_tree_add_7_25_groupi_g14377__6131(csa_tree_add_7_25_groupi_n_6720 ,csa_tree_add_7_25_groupi_n_6641 ,csa_tree_add_7_25_groupi_n_6706);
  xnor csa_tree_add_7_25_groupi_g14378__1881(csa_tree_add_7_25_groupi_n_6718 ,csa_tree_add_7_25_groupi_n_6663 ,csa_tree_add_7_25_groupi_n_2560);
  and csa_tree_add_7_25_groupi_g14379__5115(csa_tree_add_7_25_groupi_n_6706 ,csa_tree_add_7_25_groupi_n_6642 ,csa_tree_add_7_25_groupi_n_6629);
  nor csa_tree_add_7_25_groupi_g14380__7482(csa_tree_add_7_25_groupi_n_6705 ,csa_tree_add_7_25_groupi_n_2099 ,csa_tree_add_7_25_groupi_n_1120);
  nor csa_tree_add_7_25_groupi_g14381__4733(csa_tree_add_7_25_groupi_n_6704 ,csa_tree_add_7_25_groupi_n_2150 ,csa_tree_add_7_25_groupi_n_1120);
  nor csa_tree_add_7_25_groupi_g14382__6161(csa_tree_add_7_25_groupi_n_6703 ,csa_tree_add_7_25_groupi_n_2120 ,csa_tree_add_7_25_groupi_n_6647);
  nor csa_tree_add_7_25_groupi_g14383__9315(csa_tree_add_7_25_groupi_n_6702 ,csa_tree_add_7_25_groupi_n_2135 ,csa_tree_add_7_25_groupi_n_1119);
  nor csa_tree_add_7_25_groupi_g14384__9945(csa_tree_add_7_25_groupi_n_6701 ,csa_tree_add_7_25_groupi_n_2063 ,csa_tree_add_7_25_groupi_n_1125);
  nor csa_tree_add_7_25_groupi_g14385__2883(csa_tree_add_7_25_groupi_n_6700 ,csa_tree_add_7_25_groupi_n_2177 ,csa_tree_add_7_25_groupi_n_1125);
  and csa_tree_add_7_25_groupi_g14386__2346(csa_tree_add_7_25_groupi_n_6699 ,csa_tree_add_7_25_groupi_n_6655 ,csa_tree_add_7_25_groupi_n_6664);
  and csa_tree_add_7_25_groupi_g14387__1666(csa_tree_add_7_25_groupi_n_6698 ,csa_tree_add_7_25_groupi_n_6631 ,csa_tree_add_7_25_groupi_n_6626);
  or csa_tree_add_7_25_groupi_g14388__7410(csa_tree_add_7_25_groupi_n_6697 ,csa_tree_add_7_25_groupi_n_2441 ,csa_tree_add_7_25_groupi_n_6663);
  and csa_tree_add_7_25_groupi_g14389__6417(csa_tree_add_7_25_groupi_n_6696 ,csa_tree_add_7_25_groupi_n_6628 ,csa_tree_add_7_25_groupi_n_6639);
  and csa_tree_add_7_25_groupi_g14390__5477(csa_tree_add_7_25_groupi_n_6695 ,csa_tree_add_7_25_groupi_n_6627 ,csa_tree_add_7_25_groupi_n_6632);
  nor csa_tree_add_7_25_groupi_g14391__2398(csa_tree_add_7_25_groupi_n_6694 ,csa_tree_add_7_25_groupi_n_3930 ,csa_tree_add_7_25_groupi_n_6649);
  nor csa_tree_add_7_25_groupi_g14392__5107(csa_tree_add_7_25_groupi_n_6693 ,csa_tree_add_7_25_groupi_n_3865 ,csa_tree_add_7_25_groupi_n_6648);
  nor csa_tree_add_7_25_groupi_g14393__6260(csa_tree_add_7_25_groupi_n_6692 ,csa_tree_add_7_25_groupi_n_3819 ,csa_tree_add_7_25_groupi_n_6645);
  nor csa_tree_add_7_25_groupi_g14394__4319(csa_tree_add_7_25_groupi_n_6691 ,csa_tree_add_7_25_groupi_n_4002 ,csa_tree_add_7_25_groupi_n_6659);
  nor csa_tree_add_7_25_groupi_g14395__8428(csa_tree_add_7_25_groupi_n_6690 ,csa_tree_add_7_25_groupi_n_3824 ,csa_tree_add_7_25_groupi_n_6637);
  nor csa_tree_add_7_25_groupi_g14396__5526(csa_tree_add_7_25_groupi_n_6689 ,csa_tree_add_7_25_groupi_n_4071 ,csa_tree_add_7_25_groupi_n_6658);
  nor csa_tree_add_7_25_groupi_g14397__6783(csa_tree_add_7_25_groupi_n_6688 ,csa_tree_add_7_25_groupi_n_3493 ,csa_tree_add_7_25_groupi_n_6644);
  or csa_tree_add_7_25_groupi_g14398__3680(csa_tree_add_7_25_groupi_n_6709 ,csa_tree_add_7_25_groupi_n_6474 ,csa_tree_add_7_25_groupi_n_6650);
  or csa_tree_add_7_25_groupi_g14399__1617(csa_tree_add_7_25_groupi_n_6708 ,csa_tree_add_7_25_groupi_n_6471 ,csa_tree_add_7_25_groupi_n_6653);
  or csa_tree_add_7_25_groupi_g14400__2802(csa_tree_add_7_25_groupi_n_6707 ,csa_tree_add_7_25_groupi_n_6483 ,csa_tree_add_7_25_groupi_n_6660);
  xnor csa_tree_add_7_25_groupi_g14401__1705(out2[18] ,csa_tree_add_7_25_groupi_n_6576 ,csa_tree_add_7_25_groupi_n_6581);
  xnor csa_tree_add_7_25_groupi_g14402__5122(csa_tree_add_7_25_groupi_n_6676 ,csa_tree_add_7_25_groupi_n_6537 ,csa_tree_add_7_25_groupi_n_6603);
  xnor csa_tree_add_7_25_groupi_g14403__8246(csa_tree_add_7_25_groupi_n_6675 ,csa_tree_add_7_25_groupi_n_6534 ,csa_tree_add_7_25_groupi_n_6594);
  xnor csa_tree_add_7_25_groupi_g14404__7098(csa_tree_add_7_25_groupi_n_6674 ,csa_tree_add_7_25_groupi_n_6536 ,csa_tree_add_7_25_groupi_n_6600);
  xnor csa_tree_add_7_25_groupi_g14405__6131(csa_tree_add_7_25_groupi_n_6673 ,csa_tree_add_7_25_groupi_n_6591 ,csa_tree_add_7_25_groupi_n_6543);
  xnor csa_tree_add_7_25_groupi_g14406__1881(csa_tree_add_7_25_groupi_n_6672 ,csa_tree_add_7_25_groupi_n_6593 ,csa_tree_add_7_25_groupi_n_6503);
  xnor csa_tree_add_7_25_groupi_g14407__5115(csa_tree_add_7_25_groupi_n_6671 ,csa_tree_add_7_25_groupi_n_6595 ,csa_tree_add_7_25_groupi_n_6509);
  xnor csa_tree_add_7_25_groupi_g14408__7482(csa_tree_add_7_25_groupi_n_6670 ,csa_tree_add_7_25_groupi_n_6539 ,csa_tree_add_7_25_groupi_n_6597);
  xnor csa_tree_add_7_25_groupi_g14409__4733(csa_tree_add_7_25_groupi_n_6669 ,csa_tree_add_7_25_groupi_n_6589 ,csa_tree_add_7_25_groupi_n_6501);
  xnor csa_tree_add_7_25_groupi_g14410__6161(csa_tree_add_7_25_groupi_n_6668 ,csa_tree_add_7_25_groupi_n_6602 ,csa_tree_add_7_25_groupi_n_6499);
  xnor csa_tree_add_7_25_groupi_g14411__9315(csa_tree_add_7_25_groupi_n_6667 ,csa_tree_add_7_25_groupi_n_6599 ,csa_tree_add_7_25_groupi_n_6541);
  xnor csa_tree_add_7_25_groupi_g14412__9945(csa_tree_add_7_25_groupi_n_6666 ,csa_tree_add_7_25_groupi_n_6520 ,csa_tree_add_7_25_groupi_n_6582);
  xnor csa_tree_add_7_25_groupi_g14413__2883(csa_tree_add_7_25_groupi_n_6665 ,csa_tree_add_7_25_groupi_n_6535 ,csa_tree_add_7_25_groupi_n_6587);
  xnor csa_tree_add_7_25_groupi_g14414__2346(csa_tree_add_7_25_groupi_n_6687 ,csa_tree_add_7_25_groupi_n_6611 ,in3[17]);
  xnor csa_tree_add_7_25_groupi_g14415__1666(csa_tree_add_7_25_groupi_n_6686 ,csa_tree_add_7_25_groupi_n_6607 ,in3[8]);
  xnor csa_tree_add_7_25_groupi_g14416__7410(csa_tree_add_7_25_groupi_n_6685 ,csa_tree_add_7_25_groupi_n_6610 ,in3[11]);
  xnor csa_tree_add_7_25_groupi_g14417__6417(csa_tree_add_7_25_groupi_n_6684 ,csa_tree_add_7_25_groupi_n_6613 ,in3[14]);
  xnor csa_tree_add_7_25_groupi_g14418__5477(csa_tree_add_7_25_groupi_n_6683 ,csa_tree_add_7_25_groupi_n_6612 ,in3[2]);
  xnor csa_tree_add_7_25_groupi_g14419__2398(csa_tree_add_7_25_groupi_n_6682 ,csa_tree_add_7_25_groupi_n_6609 ,in3[20]);
  xnor csa_tree_add_7_25_groupi_g14420__5107(csa_tree_add_7_25_groupi_n_6681 ,csa_tree_add_7_25_groupi_n_6608 ,in3[5]);
  xnor csa_tree_add_7_25_groupi_g14421__6260(csa_tree_add_7_25_groupi_n_6680 ,csa_tree_add_7_25_groupi_n_6604 ,csa_tree_add_7_25_groupi_n_6490);
  xnor csa_tree_add_7_25_groupi_g14422__4319(csa_tree_add_7_25_groupi_n_6679 ,csa_tree_add_7_25_groupi_n_6605 ,csa_tree_add_7_25_groupi_n_6488);
  xnor csa_tree_add_7_25_groupi_g14423__8428(csa_tree_add_7_25_groupi_n_6678 ,csa_tree_add_7_25_groupi_n_6606 ,csa_tree_add_7_25_groupi_n_6489);
  and csa_tree_add_7_25_groupi_g14424__5526(csa_tree_add_7_25_groupi_n_6662 ,csa_tree_add_7_25_groupi_n_6534 ,csa_tree_add_7_25_groupi_n_6594);
  and csa_tree_add_7_25_groupi_g14425__6783(csa_tree_add_7_25_groupi_n_6661 ,csa_tree_add_7_25_groupi_n_6535 ,csa_tree_add_7_25_groupi_n_6587);
  and csa_tree_add_7_25_groupi_g14426__3680(csa_tree_add_7_25_groupi_n_6660 ,csa_tree_add_7_25_groupi_n_6604 ,csa_tree_add_7_25_groupi_n_6475);
  or csa_tree_add_7_25_groupi_g14427__1617(csa_tree_add_7_25_groupi_n_6659 ,csa_tree_add_7_25_groupi_n_3435 ,csa_tree_add_7_25_groupi_n_6619);
  or csa_tree_add_7_25_groupi_g14428__2802(csa_tree_add_7_25_groupi_n_6658 ,csa_tree_add_7_25_groupi_n_3432 ,csa_tree_add_7_25_groupi_n_6620);
  and csa_tree_add_7_25_groupi_g14429__1705(csa_tree_add_7_25_groupi_n_6657 ,csa_tree_add_7_25_groupi_n_6536 ,csa_tree_add_7_25_groupi_n_6600);
  or csa_tree_add_7_25_groupi_g14430__5122(csa_tree_add_7_25_groupi_n_6656 ,csa_tree_add_7_25_groupi_n_6536 ,csa_tree_add_7_25_groupi_n_6600);
  or csa_tree_add_7_25_groupi_g14431__8246(csa_tree_add_7_25_groupi_n_6655 ,csa_tree_add_7_25_groupi_n_6535 ,csa_tree_add_7_25_groupi_n_6587);
  or csa_tree_add_7_25_groupi_g14432__7098(csa_tree_add_7_25_groupi_n_6654 ,csa_tree_add_7_25_groupi_n_6534 ,csa_tree_add_7_25_groupi_n_6594);
  and csa_tree_add_7_25_groupi_g14433__6131(csa_tree_add_7_25_groupi_n_6653 ,csa_tree_add_7_25_groupi_n_6605 ,csa_tree_add_7_25_groupi_n_6472);
  and csa_tree_add_7_25_groupi_g14434__1881(csa_tree_add_7_25_groupi_n_6652 ,csa_tree_add_7_25_groupi_n_6537 ,csa_tree_add_7_25_groupi_n_6603);
  or csa_tree_add_7_25_groupi_g14435__5115(csa_tree_add_7_25_groupi_n_6651 ,csa_tree_add_7_25_groupi_n_6537 ,csa_tree_add_7_25_groupi_n_6603);
  and csa_tree_add_7_25_groupi_g14436__7482(csa_tree_add_7_25_groupi_n_6650 ,csa_tree_add_7_25_groupi_n_6606 ,csa_tree_add_7_25_groupi_n_6473);
  or csa_tree_add_7_25_groupi_g14437__4733(csa_tree_add_7_25_groupi_n_6649 ,csa_tree_add_7_25_groupi_n_3775 ,csa_tree_add_7_25_groupi_n_6616);
  or csa_tree_add_7_25_groupi_g14438__6161(csa_tree_add_7_25_groupi_n_6648 ,csa_tree_add_7_25_groupi_n_3778 ,csa_tree_add_7_25_groupi_n_6618);
  or csa_tree_add_7_25_groupi_g14439__9315(csa_tree_add_7_25_groupi_n_6664 ,csa_tree_add_7_25_groupi_n_6571 ,csa_tree_add_7_25_groupi_n_6614);
  and csa_tree_add_7_25_groupi_g14440__9945(csa_tree_add_7_25_groupi_n_6663 ,csa_tree_add_7_25_groupi_n_2467 ,csa_tree_add_7_25_groupi_n_6617);
  nor csa_tree_add_7_25_groupi_g14441__2883(csa_tree_add_7_25_groupi_n_6646 ,csa_tree_add_7_25_groupi_n_6599 ,csa_tree_add_7_25_groupi_n_6540);
  or csa_tree_add_7_25_groupi_g14442__2346(csa_tree_add_7_25_groupi_n_6645 ,csa_tree_add_7_25_groupi_n_3774 ,csa_tree_add_7_25_groupi_n_6622);
  or csa_tree_add_7_25_groupi_g14443__1666(csa_tree_add_7_25_groupi_n_6644 ,csa_tree_add_7_25_groupi_n_3405 ,csa_tree_add_7_25_groupi_n_6615);
  or csa_tree_add_7_25_groupi_g14444__7410(csa_tree_add_7_25_groupi_n_6643 ,csa_tree_add_7_25_groupi_n_6539 ,csa_tree_add_7_25_groupi_n_6596);
  or csa_tree_add_7_25_groupi_g14445__6417(csa_tree_add_7_25_groupi_n_6642 ,csa_tree_add_7_25_groupi_n_6602 ,csa_tree_add_7_25_groupi_n_6498);
  nor csa_tree_add_7_25_groupi_g14446__5477(csa_tree_add_7_25_groupi_n_6641 ,csa_tree_add_7_25_groupi_n_6601 ,csa_tree_add_7_25_groupi_n_6499);
  nor csa_tree_add_7_25_groupi_g14447__2398(csa_tree_add_7_25_groupi_n_6640 ,csa_tree_add_7_25_groupi_n_6538 ,csa_tree_add_7_25_groupi_n_6597);
  or csa_tree_add_7_25_groupi_g14448__5107(csa_tree_add_7_25_groupi_n_6639 ,csa_tree_add_7_25_groupi_n_6589 ,csa_tree_add_7_25_groupi_n_6500);
  nor csa_tree_add_7_25_groupi_g14449__6260(csa_tree_add_7_25_groupi_n_6638 ,csa_tree_add_7_25_groupi_n_6588 ,csa_tree_add_7_25_groupi_n_6501);
  or csa_tree_add_7_25_groupi_g14450__4319(csa_tree_add_7_25_groupi_n_6637 ,csa_tree_add_7_25_groupi_n_3777 ,csa_tree_add_7_25_groupi_n_6621);
  or csa_tree_add_7_25_groupi_g14451__8428(csa_tree_add_7_25_groupi_n_6636 ,csa_tree_add_7_25_groupi_n_6598 ,csa_tree_add_7_25_groupi_n_6541);
  nor csa_tree_add_7_25_groupi_g14452__5526(csa_tree_add_7_25_groupi_n_6635 ,csa_tree_add_7_25_groupi_n_6591 ,csa_tree_add_7_25_groupi_n_6542);
  or csa_tree_add_7_25_groupi_g14453__6783(csa_tree_add_7_25_groupi_n_6634 ,csa_tree_add_7_25_groupi_n_6590 ,csa_tree_add_7_25_groupi_n_6543);
  nor csa_tree_add_7_25_groupi_g14454__3680(csa_tree_add_7_25_groupi_n_6633 ,csa_tree_add_7_25_groupi_n_6592 ,csa_tree_add_7_25_groupi_n_6503);
  or csa_tree_add_7_25_groupi_g14455__1617(csa_tree_add_7_25_groupi_n_6632 ,csa_tree_add_7_25_groupi_n_6593 ,csa_tree_add_7_25_groupi_n_6502);
  or csa_tree_add_7_25_groupi_g14456__2802(csa_tree_add_7_25_groupi_n_6631 ,csa_tree_add_7_25_groupi_n_6595 ,csa_tree_add_7_25_groupi_n_6509);
  and csa_tree_add_7_25_groupi_g14457__1705(csa_tree_add_7_25_groupi_n_6630 ,csa_tree_add_7_25_groupi_n_6595 ,csa_tree_add_7_25_groupi_n_6509);
  xnor csa_tree_add_7_25_groupi_g14458__5122(csa_tree_add_7_25_groupi_n_6647 ,csa_tree_add_7_25_groupi_n_6575 ,csa_tree_add_7_25_groupi_n_2561);
  nor csa_tree_add_7_25_groupi_g14459__8246(csa_tree_add_7_25_groupi_n_6622 ,csa_tree_add_7_25_groupi_n_2144 ,csa_tree_add_7_25_groupi_n_6560);
  nor csa_tree_add_7_25_groupi_g14460__7098(csa_tree_add_7_25_groupi_n_6621 ,csa_tree_add_7_25_groupi_n_2111 ,csa_tree_add_7_25_groupi_n_1144);
  nor csa_tree_add_7_25_groupi_g14461__6131(csa_tree_add_7_25_groupi_n_6620 ,csa_tree_add_7_25_groupi_n_2090 ,csa_tree_add_7_25_groupi_n_1258);
  nor csa_tree_add_7_25_groupi_g14462__1881(csa_tree_add_7_25_groupi_n_6619 ,csa_tree_add_7_25_groupi_n_2165 ,csa_tree_add_7_25_groupi_n_1144);
  nor csa_tree_add_7_25_groupi_g14463__5115(csa_tree_add_7_25_groupi_n_6618 ,csa_tree_add_7_25_groupi_n_2070 ,csa_tree_add_7_25_groupi_n_1258);
  or csa_tree_add_7_25_groupi_g14464__7482(csa_tree_add_7_25_groupi_n_6617 ,csa_tree_add_7_25_groupi_n_2483 ,csa_tree_add_7_25_groupi_n_6575);
  nor csa_tree_add_7_25_groupi_g14465__4733(csa_tree_add_7_25_groupi_n_6616 ,csa_tree_add_7_25_groupi_n_2037 ,csa_tree_add_7_25_groupi_n_1259);
  nor csa_tree_add_7_25_groupi_g14466__6161(csa_tree_add_7_25_groupi_n_6615 ,csa_tree_add_7_25_groupi_n_2168 ,csa_tree_add_7_25_groupi_n_1259);
  and csa_tree_add_7_25_groupi_g14467__9315(csa_tree_add_7_25_groupi_n_6614 ,csa_tree_add_7_25_groupi_n_6576 ,csa_tree_add_7_25_groupi_n_6569);
  nor csa_tree_add_7_25_groupi_g14468__9945(csa_tree_add_7_25_groupi_n_6613 ,csa_tree_add_7_25_groupi_n_3924 ,csa_tree_add_7_25_groupi_n_6558);
  nor csa_tree_add_7_25_groupi_g14469__2883(csa_tree_add_7_25_groupi_n_6612 ,csa_tree_add_7_25_groupi_n_3473 ,csa_tree_add_7_25_groupi_n_6553);
  nor csa_tree_add_7_25_groupi_g14470__2346(csa_tree_add_7_25_groupi_n_6611 ,csa_tree_add_7_25_groupi_n_3914 ,csa_tree_add_7_25_groupi_n_6559);
  nor csa_tree_add_7_25_groupi_g14471__1666(csa_tree_add_7_25_groupi_n_6610 ,csa_tree_add_7_25_groupi_n_3911 ,csa_tree_add_7_25_groupi_n_6557);
  nor csa_tree_add_7_25_groupi_g14472__7410(csa_tree_add_7_25_groupi_n_6609 ,csa_tree_add_7_25_groupi_n_3942 ,csa_tree_add_7_25_groupi_n_6574);
  nor csa_tree_add_7_25_groupi_g14473__6417(csa_tree_add_7_25_groupi_n_6608 ,csa_tree_add_7_25_groupi_n_3994 ,csa_tree_add_7_25_groupi_n_6564);
  nor csa_tree_add_7_25_groupi_g14474__5477(csa_tree_add_7_25_groupi_n_6607 ,csa_tree_add_7_25_groupi_n_3873 ,csa_tree_add_7_25_groupi_n_6556);
  or csa_tree_add_7_25_groupi_g14475__2398(csa_tree_add_7_25_groupi_n_6629 ,csa_tree_add_7_25_groupi_n_6377 ,csa_tree_add_7_25_groupi_n_6552);
  or csa_tree_add_7_25_groupi_g14476__5107(csa_tree_add_7_25_groupi_n_6628 ,csa_tree_add_7_25_groupi_n_6371 ,csa_tree_add_7_25_groupi_n_6547);
  or csa_tree_add_7_25_groupi_g14477__6260(csa_tree_add_7_25_groupi_n_6627 ,csa_tree_add_7_25_groupi_n_6365 ,csa_tree_add_7_25_groupi_n_6546);
  or csa_tree_add_7_25_groupi_g14478__4319(csa_tree_add_7_25_groupi_n_6626 ,csa_tree_add_7_25_groupi_n_6399 ,csa_tree_add_7_25_groupi_n_6565);
  or csa_tree_add_7_25_groupi_g14479__8428(csa_tree_add_7_25_groupi_n_6625 ,csa_tree_add_7_25_groupi_n_6384 ,csa_tree_add_7_25_groupi_n_6563);
  or csa_tree_add_7_25_groupi_g14480__5526(csa_tree_add_7_25_groupi_n_6624 ,csa_tree_add_7_25_groupi_n_6387 ,csa_tree_add_7_25_groupi_n_6562);
  or csa_tree_add_7_25_groupi_g14481__6783(csa_tree_add_7_25_groupi_n_6623 ,csa_tree_add_7_25_groupi_n_6392 ,csa_tree_add_7_25_groupi_n_6566);
  not csa_tree_add_7_25_groupi_g14482(csa_tree_add_7_25_groupi_n_6601 ,csa_tree_add_7_25_groupi_n_6602);
  not csa_tree_add_7_25_groupi_g14483(csa_tree_add_7_25_groupi_n_6598 ,csa_tree_add_7_25_groupi_n_6599);
  not csa_tree_add_7_25_groupi_g14484(csa_tree_add_7_25_groupi_n_6596 ,csa_tree_add_7_25_groupi_n_6597);
  not csa_tree_add_7_25_groupi_g14485(csa_tree_add_7_25_groupi_n_6592 ,csa_tree_add_7_25_groupi_n_6593);
  not csa_tree_add_7_25_groupi_g14486(csa_tree_add_7_25_groupi_n_6590 ,csa_tree_add_7_25_groupi_n_6591);
  not csa_tree_add_7_25_groupi_g14487(csa_tree_add_7_25_groupi_n_6588 ,csa_tree_add_7_25_groupi_n_6589);
  xnor csa_tree_add_7_25_groupi_g14488__3680(out2[17] ,csa_tree_add_7_25_groupi_n_6485 ,csa_tree_add_7_25_groupi_n_6487);
  xnor csa_tree_add_7_25_groupi_g14489__1617(csa_tree_add_7_25_groupi_n_6585 ,csa_tree_add_7_25_groupi_n_6466 ,csa_tree_add_7_25_groupi_n_6506);
  xnor csa_tree_add_7_25_groupi_g14490__2802(csa_tree_add_7_25_groupi_n_6584 ,csa_tree_add_7_25_groupi_n_6495 ,csa_tree_add_7_25_groupi_n_6465);
  xnor csa_tree_add_7_25_groupi_g14491__1705(csa_tree_add_7_25_groupi_n_6583 ,csa_tree_add_7_25_groupi_n_6470 ,csa_tree_add_7_25_groupi_n_6497);
  xnor csa_tree_add_7_25_groupi_g14492__5122(csa_tree_add_7_25_groupi_n_6582 ,csa_tree_add_7_25_groupi_n_6486 ,csa_tree_add_7_25_groupi_n_6403);
  xnor csa_tree_add_7_25_groupi_g14493__8246(csa_tree_add_7_25_groupi_n_6581 ,csa_tree_add_7_25_groupi_n_6451 ,csa_tree_add_7_25_groupi_n_6507);
  xnor csa_tree_add_7_25_groupi_g14494__7098(csa_tree_add_7_25_groupi_n_6580 ,csa_tree_add_7_25_groupi_n_6450 ,csa_tree_add_7_25_groupi_n_6505);
  xnor csa_tree_add_7_25_groupi_g14495__6131(csa_tree_add_7_25_groupi_n_6579 ,csa_tree_add_7_25_groupi_n_6452 ,csa_tree_add_7_25_groupi_n_6504);
  xnor csa_tree_add_7_25_groupi_g14496__1881(csa_tree_add_7_25_groupi_n_6578 ,csa_tree_add_7_25_groupi_n_6508 ,csa_tree_add_7_25_groupi_n_6449);
  xnor csa_tree_add_7_25_groupi_g14497__5115(csa_tree_add_7_25_groupi_n_6577 ,csa_tree_add_7_25_groupi_n_6493 ,csa_tree_add_7_25_groupi_n_6468);
  xnor csa_tree_add_7_25_groupi_g14498__7482(csa_tree_add_7_25_groupi_n_6606 ,csa_tree_add_7_25_groupi_n_6517 ,in3[5]);
  xnor csa_tree_add_7_25_groupi_g14499__4733(csa_tree_add_7_25_groupi_n_6605 ,csa_tree_add_7_25_groupi_n_6519 ,in3[8]);
  xnor csa_tree_add_7_25_groupi_g14500__6161(csa_tree_add_7_25_groupi_n_6604 ,csa_tree_add_7_25_groupi_n_6524 ,in3[2]);
  xnor csa_tree_add_7_25_groupi_g14501__9315(csa_tree_add_7_25_groupi_n_6603 ,csa_tree_add_7_25_groupi_n_6516 ,csa_tree_add_7_25_groupi_n_6411);
  xnor csa_tree_add_7_25_groupi_g14502__9945(csa_tree_add_7_25_groupi_n_6602 ,csa_tree_add_7_25_groupi_n_6522 ,in3[20]);
  xnor csa_tree_add_7_25_groupi_g14503__2883(csa_tree_add_7_25_groupi_n_6600 ,csa_tree_add_7_25_groupi_n_6511 ,csa_tree_add_7_25_groupi_n_6409);
  xnor csa_tree_add_7_25_groupi_g14504__2346(csa_tree_add_7_25_groupi_n_6599 ,csa_tree_add_7_25_groupi_n_6514 ,csa_tree_add_7_25_groupi_n_6402);
  xnor csa_tree_add_7_25_groupi_g14505__1666(csa_tree_add_7_25_groupi_n_6597 ,csa_tree_add_7_25_groupi_n_6515 ,csa_tree_add_7_25_groupi_n_6404);
  xnor csa_tree_add_7_25_groupi_g14506__7410(csa_tree_add_7_25_groupi_n_6595 ,csa_tree_add_7_25_groupi_n_6523 ,in3[11]);
  xnor csa_tree_add_7_25_groupi_g14507__6417(csa_tree_add_7_25_groupi_n_6594 ,csa_tree_add_7_25_groupi_n_6510 ,csa_tree_add_7_25_groupi_n_6410);
  xnor csa_tree_add_7_25_groupi_g14508__5477(csa_tree_add_7_25_groupi_n_6593 ,csa_tree_add_7_25_groupi_n_6518 ,in3[14]);
  xnor csa_tree_add_7_25_groupi_g14509__2398(csa_tree_add_7_25_groupi_n_6591 ,csa_tree_add_7_25_groupi_n_6513 ,csa_tree_add_7_25_groupi_n_6413);
  xnor csa_tree_add_7_25_groupi_g14510__5107(csa_tree_add_7_25_groupi_n_6589 ,csa_tree_add_7_25_groupi_n_6521 ,in3[17]);
  xnor csa_tree_add_7_25_groupi_g14511__6260(csa_tree_add_7_25_groupi_n_6587 ,csa_tree_add_7_25_groupi_n_6512 ,csa_tree_add_7_25_groupi_n_6412);
  or csa_tree_add_7_25_groupi_g14512__4319(csa_tree_add_7_25_groupi_n_6574 ,csa_tree_add_7_25_groupi_n_3770 ,csa_tree_add_7_25_groupi_n_6526);
  or csa_tree_add_7_25_groupi_g14513__8428(csa_tree_add_7_25_groupi_n_6573 ,csa_tree_add_7_25_groupi_n_6466 ,csa_tree_add_7_25_groupi_n_6506);
  and csa_tree_add_7_25_groupi_g14514__5526(csa_tree_add_7_25_groupi_n_6572 ,csa_tree_add_7_25_groupi_n_6466 ,csa_tree_add_7_25_groupi_n_6506);
  and csa_tree_add_7_25_groupi_g14515__6783(csa_tree_add_7_25_groupi_n_6571 ,csa_tree_add_7_25_groupi_n_6451 ,csa_tree_add_7_25_groupi_n_6507);
  or csa_tree_add_7_25_groupi_g14516__3680(csa_tree_add_7_25_groupi_n_6570 ,csa_tree_add_7_25_groupi_n_6452 ,csa_tree_add_7_25_groupi_n_6504);
  or csa_tree_add_7_25_groupi_g14517__1617(csa_tree_add_7_25_groupi_n_6569 ,csa_tree_add_7_25_groupi_n_6451 ,csa_tree_add_7_25_groupi_n_6507);
  and csa_tree_add_7_25_groupi_g14518__2802(csa_tree_add_7_25_groupi_n_6568 ,csa_tree_add_7_25_groupi_n_6450 ,csa_tree_add_7_25_groupi_n_6505);
  or csa_tree_add_7_25_groupi_g14519__1705(csa_tree_add_7_25_groupi_n_6567 ,csa_tree_add_7_25_groupi_n_6450 ,csa_tree_add_7_25_groupi_n_6505);
  and csa_tree_add_7_25_groupi_g14520__5122(csa_tree_add_7_25_groupi_n_6566 ,csa_tree_add_7_25_groupi_n_6512 ,csa_tree_add_7_25_groupi_n_6393);
  and csa_tree_add_7_25_groupi_g14521__8246(csa_tree_add_7_25_groupi_n_6565 ,csa_tree_add_7_25_groupi_n_6510 ,csa_tree_add_7_25_groupi_n_6389);
  or csa_tree_add_7_25_groupi_g14522__7098(csa_tree_add_7_25_groupi_n_6564 ,csa_tree_add_7_25_groupi_n_3423 ,csa_tree_add_7_25_groupi_n_6528);
  and csa_tree_add_7_25_groupi_g14523__6131(csa_tree_add_7_25_groupi_n_6563 ,csa_tree_add_7_25_groupi_n_6511 ,csa_tree_add_7_25_groupi_n_6388);
  and csa_tree_add_7_25_groupi_g14524__1881(csa_tree_add_7_25_groupi_n_6562 ,csa_tree_add_7_25_groupi_n_6516 ,csa_tree_add_7_25_groupi_n_6386);
  and csa_tree_add_7_25_groupi_g14525__5115(csa_tree_add_7_25_groupi_n_6561 ,csa_tree_add_7_25_groupi_n_6452 ,csa_tree_add_7_25_groupi_n_6504);
  or csa_tree_add_7_25_groupi_g14526__7482(csa_tree_add_7_25_groupi_n_6576 ,csa_tree_add_7_25_groupi_n_6531 ,csa_tree_add_7_25_groupi_n_6479);
  and csa_tree_add_7_25_groupi_g14527__4733(csa_tree_add_7_25_groupi_n_6575 ,csa_tree_add_7_25_groupi_n_2433 ,csa_tree_add_7_25_groupi_n_6532);
  or csa_tree_add_7_25_groupi_g14528__6161(csa_tree_add_7_25_groupi_n_6559 ,csa_tree_add_7_25_groupi_n_3772 ,csa_tree_add_7_25_groupi_n_6527);
  or csa_tree_add_7_25_groupi_g14529__9315(csa_tree_add_7_25_groupi_n_6558 ,csa_tree_add_7_25_groupi_n_3771 ,csa_tree_add_7_25_groupi_n_6529);
  or csa_tree_add_7_25_groupi_g14530__9945(csa_tree_add_7_25_groupi_n_6557 ,csa_tree_add_7_25_groupi_n_3769 ,csa_tree_add_7_25_groupi_n_6530);
  or csa_tree_add_7_25_groupi_g14531__2883(csa_tree_add_7_25_groupi_n_6556 ,csa_tree_add_7_25_groupi_n_3768 ,csa_tree_add_7_25_groupi_n_6525);
  nor csa_tree_add_7_25_groupi_g14532__2346(csa_tree_add_7_25_groupi_n_6555 ,csa_tree_add_7_25_groupi_n_6493 ,csa_tree_add_7_25_groupi_n_6467);
  or csa_tree_add_7_25_groupi_g14533__1666(csa_tree_add_7_25_groupi_n_6554 ,csa_tree_add_7_25_groupi_n_6492 ,csa_tree_add_7_25_groupi_n_6468);
  or csa_tree_add_7_25_groupi_g14534__7410(csa_tree_add_7_25_groupi_n_6553 ,csa_tree_add_7_25_groupi_n_3381 ,csa_tree_add_7_25_groupi_n_6533);
  and csa_tree_add_7_25_groupi_g14535__6417(csa_tree_add_7_25_groupi_n_6552 ,csa_tree_add_7_25_groupi_n_6515 ,csa_tree_add_7_25_groupi_n_6376);
  nor csa_tree_add_7_25_groupi_g14536__5477(csa_tree_add_7_25_groupi_n_6551 ,csa_tree_add_7_25_groupi_n_6495 ,csa_tree_add_7_25_groupi_n_6464);
  or csa_tree_add_7_25_groupi_g14537__2398(csa_tree_add_7_25_groupi_n_6550 ,csa_tree_add_7_25_groupi_n_6494 ,csa_tree_add_7_25_groupi_n_6465);
  nor csa_tree_add_7_25_groupi_g14538__5107(csa_tree_add_7_25_groupi_n_6549 ,csa_tree_add_7_25_groupi_n_6469 ,csa_tree_add_7_25_groupi_n_6497);
  or csa_tree_add_7_25_groupi_g14539__6260(csa_tree_add_7_25_groupi_n_6548 ,csa_tree_add_7_25_groupi_n_6470 ,csa_tree_add_7_25_groupi_n_6496);
  and csa_tree_add_7_25_groupi_g14540__4319(csa_tree_add_7_25_groupi_n_6547 ,csa_tree_add_7_25_groupi_n_6514 ,csa_tree_add_7_25_groupi_n_6370);
  and csa_tree_add_7_25_groupi_g14541__8428(csa_tree_add_7_25_groupi_n_6546 ,csa_tree_add_7_25_groupi_n_6513 ,csa_tree_add_7_25_groupi_n_6368);
  and csa_tree_add_7_25_groupi_g14542__5526(csa_tree_add_7_25_groupi_n_6545 ,csa_tree_add_7_25_groupi_n_6508 ,csa_tree_add_7_25_groupi_n_6449);
  or csa_tree_add_7_25_groupi_g14543__6783(csa_tree_add_7_25_groupi_n_6544 ,csa_tree_add_7_25_groupi_n_6508 ,csa_tree_add_7_25_groupi_n_6449);
  xnor csa_tree_add_7_25_groupi_g14544__3680(csa_tree_add_7_25_groupi_n_6560 ,csa_tree_add_7_25_groupi_n_6484 ,csa_tree_add_7_25_groupi_n_2562);
  not csa_tree_add_7_25_groupi_g14545(csa_tree_add_7_25_groupi_n_6542 ,csa_tree_add_7_25_groupi_n_6543);
  not csa_tree_add_7_25_groupi_g14546(csa_tree_add_7_25_groupi_n_6540 ,csa_tree_add_7_25_groupi_n_6541);
  not csa_tree_add_7_25_groupi_g14547(csa_tree_add_7_25_groupi_n_6538 ,csa_tree_add_7_25_groupi_n_6539);
  nor csa_tree_add_7_25_groupi_g14548__1617(csa_tree_add_7_25_groupi_n_6533 ,csa_tree_add_7_25_groupi_n_2178 ,csa_tree_add_7_25_groupi_n_6463);
  or csa_tree_add_7_25_groupi_g14549__2802(csa_tree_add_7_25_groupi_n_6532 ,csa_tree_add_7_25_groupi_n_2447 ,csa_tree_add_7_25_groupi_n_6484);
  and csa_tree_add_7_25_groupi_g14550__1705(csa_tree_add_7_25_groupi_n_6531 ,csa_tree_add_7_25_groupi_n_6481 ,csa_tree_add_7_25_groupi_n_6485);
  nor csa_tree_add_7_25_groupi_g14551__5122(csa_tree_add_7_25_groupi_n_6530 ,csa_tree_add_7_25_groupi_n_2100 ,csa_tree_add_7_25_groupi_n_1135);
  nor csa_tree_add_7_25_groupi_g14552__8246(csa_tree_add_7_25_groupi_n_6529 ,csa_tree_add_7_25_groupi_n_2151 ,csa_tree_add_7_25_groupi_n_1288);
  nor csa_tree_add_7_25_groupi_g14553__7098(csa_tree_add_7_25_groupi_n_6528 ,csa_tree_add_7_25_groupi_n_2136 ,csa_tree_add_7_25_groupi_n_1135);
  nor csa_tree_add_7_25_groupi_g14554__6131(csa_tree_add_7_25_groupi_n_6527 ,csa_tree_add_7_25_groupi_n_2067 ,csa_tree_add_7_25_groupi_n_1288);
  nor csa_tree_add_7_25_groupi_g14555__1881(csa_tree_add_7_25_groupi_n_6526 ,csa_tree_add_7_25_groupi_n_2036 ,csa_tree_add_7_25_groupi_n_1289);
  nor csa_tree_add_7_25_groupi_g14556__5115(csa_tree_add_7_25_groupi_n_6525 ,csa_tree_add_7_25_groupi_n_2121 ,csa_tree_add_7_25_groupi_n_1289);
  nor csa_tree_add_7_25_groupi_g14557__7482(csa_tree_add_7_25_groupi_n_6524 ,csa_tree_add_7_25_groupi_n_3494 ,csa_tree_add_7_25_groupi_n_6455);
  nor csa_tree_add_7_25_groupi_g14558__4733(csa_tree_add_7_25_groupi_n_6523 ,csa_tree_add_7_25_groupi_n_3945 ,csa_tree_add_7_25_groupi_n_6459);
  nor csa_tree_add_7_25_groupi_g14559__6161(csa_tree_add_7_25_groupi_n_6522 ,csa_tree_add_7_25_groupi_n_3814 ,csa_tree_add_7_25_groupi_n_6461);
  nor csa_tree_add_7_25_groupi_g14560__9315(csa_tree_add_7_25_groupi_n_6521 ,csa_tree_add_7_25_groupi_n_3825 ,csa_tree_add_7_25_groupi_n_6460);
  or csa_tree_add_7_25_groupi_g14561__9945(csa_tree_add_7_25_groupi_n_6520 ,csa_tree_add_7_25_groupi_n_6274 ,csa_tree_add_7_25_groupi_n_6458);
  nor csa_tree_add_7_25_groupi_g14562__2883(csa_tree_add_7_25_groupi_n_6519 ,csa_tree_add_7_25_groupi_n_4012 ,csa_tree_add_7_25_groupi_n_6457);
  nor csa_tree_add_7_25_groupi_g14563__2346(csa_tree_add_7_25_groupi_n_6518 ,csa_tree_add_7_25_groupi_n_4035 ,csa_tree_add_7_25_groupi_n_6462);
  nor csa_tree_add_7_25_groupi_g14564__1666(csa_tree_add_7_25_groupi_n_6517 ,csa_tree_add_7_25_groupi_n_3991 ,csa_tree_add_7_25_groupi_n_6482);
  or csa_tree_add_7_25_groupi_g14565__7410(csa_tree_add_7_25_groupi_n_6543 ,csa_tree_add_7_25_groupi_n_6301 ,csa_tree_add_7_25_groupi_n_6476);
  or csa_tree_add_7_25_groupi_g14566__6417(csa_tree_add_7_25_groupi_n_6541 ,csa_tree_add_7_25_groupi_n_6272 ,csa_tree_add_7_25_groupi_n_6454);
  or csa_tree_add_7_25_groupi_g14567__5477(csa_tree_add_7_25_groupi_n_6539 ,csa_tree_add_7_25_groupi_n_6275 ,csa_tree_add_7_25_groupi_n_6456);
  or csa_tree_add_7_25_groupi_g14568__2398(csa_tree_add_7_25_groupi_n_6537 ,csa_tree_add_7_25_groupi_n_6289 ,csa_tree_add_7_25_groupi_n_6480);
  or csa_tree_add_7_25_groupi_g14569__5107(csa_tree_add_7_25_groupi_n_6536 ,csa_tree_add_7_25_groupi_n_6302 ,csa_tree_add_7_25_groupi_n_6477);
  or csa_tree_add_7_25_groupi_g14570__6260(csa_tree_add_7_25_groupi_n_6535 ,csa_tree_add_7_25_groupi_n_6297 ,csa_tree_add_7_25_groupi_n_6478);
  or csa_tree_add_7_25_groupi_g14571__4319(csa_tree_add_7_25_groupi_n_6534 ,csa_tree_add_7_25_groupi_n_6267 ,csa_tree_add_7_25_groupi_n_6453);
  not csa_tree_add_7_25_groupi_g14572(csa_tree_add_7_25_groupi_n_6502 ,csa_tree_add_7_25_groupi_n_6503);
  not csa_tree_add_7_25_groupi_g14573(csa_tree_add_7_25_groupi_n_6500 ,csa_tree_add_7_25_groupi_n_6501);
  not csa_tree_add_7_25_groupi_g14574(csa_tree_add_7_25_groupi_n_6498 ,csa_tree_add_7_25_groupi_n_6499);
  not csa_tree_add_7_25_groupi_g14575(csa_tree_add_7_25_groupi_n_6496 ,csa_tree_add_7_25_groupi_n_6497);
  not csa_tree_add_7_25_groupi_g14576(csa_tree_add_7_25_groupi_n_6494 ,csa_tree_add_7_25_groupi_n_6495);
  not csa_tree_add_7_25_groupi_g14577(csa_tree_add_7_25_groupi_n_6492 ,csa_tree_add_7_25_groupi_n_6493);
  xnor csa_tree_add_7_25_groupi_g14578__8428(out2[16] ,csa_tree_add_7_25_groupi_n_6400 ,csa_tree_add_7_25_groupi_n_6414);
  xnor csa_tree_add_7_25_groupi_g14579__5526(csa_tree_add_7_25_groupi_n_6490 ,csa_tree_add_7_25_groupi_n_6417 ,csa_tree_add_7_25_groupi_n_6356);
  xnor csa_tree_add_7_25_groupi_g14580__6783(csa_tree_add_7_25_groupi_n_6489 ,csa_tree_add_7_25_groupi_n_6418 ,csa_tree_add_7_25_groupi_n_6358);
  xnor csa_tree_add_7_25_groupi_g14581__3680(csa_tree_add_7_25_groupi_n_6488 ,csa_tree_add_7_25_groupi_n_6357 ,csa_tree_add_7_25_groupi_n_6419);
  xnor csa_tree_add_7_25_groupi_g14582__1617(csa_tree_add_7_25_groupi_n_6487 ,csa_tree_add_7_25_groupi_n_6416 ,csa_tree_add_7_25_groupi_n_6355);
  xnor csa_tree_add_7_25_groupi_g14583__2802(csa_tree_add_7_25_groupi_n_6486 ,csa_tree_add_7_25_groupi_n_6428 ,in3[23]);
  xnor csa_tree_add_7_25_groupi_g14584__1705(csa_tree_add_7_25_groupi_n_6516 ,csa_tree_add_7_25_groupi_n_6434 ,in3[8]);
  xnor csa_tree_add_7_25_groupi_g14585__5122(csa_tree_add_7_25_groupi_n_6515 ,csa_tree_add_7_25_groupi_n_6432 ,in3[20]);
  xnor csa_tree_add_7_25_groupi_g14586__8246(csa_tree_add_7_25_groupi_n_6514 ,csa_tree_add_7_25_groupi_n_6433 ,in3[17]);
  xnor csa_tree_add_7_25_groupi_g14587__7098(csa_tree_add_7_25_groupi_n_6513 ,csa_tree_add_7_25_groupi_n_6429 ,in3[14]);
  xnor csa_tree_add_7_25_groupi_g14588__6131(csa_tree_add_7_25_groupi_n_6512 ,csa_tree_add_7_25_groupi_n_6430 ,in3[2]);
  xnor csa_tree_add_7_25_groupi_g14589__1881(csa_tree_add_7_25_groupi_n_6511 ,csa_tree_add_7_25_groupi_n_6431 ,in3[5]);
  xnor csa_tree_add_7_25_groupi_g14590__5115(csa_tree_add_7_25_groupi_n_6510 ,csa_tree_add_7_25_groupi_n_6435 ,in3[11]);
  xnor csa_tree_add_7_25_groupi_g14591__7482(csa_tree_add_7_25_groupi_n_6509 ,csa_tree_add_7_25_groupi_n_6361 ,csa_tree_add_7_25_groupi_n_6407);
  xnor csa_tree_add_7_25_groupi_g14592__4733(csa_tree_add_7_25_groupi_n_6508 ,csa_tree_add_7_25_groupi_n_6427 ,csa_tree_add_7_25_groupi_n_6306);
  xnor csa_tree_add_7_25_groupi_g14593__6161(csa_tree_add_7_25_groupi_n_6507 ,csa_tree_add_7_25_groupi_n_6421 ,csa_tree_add_7_25_groupi_n_6308);
  xnor csa_tree_add_7_25_groupi_g14594__9315(csa_tree_add_7_25_groupi_n_6506 ,csa_tree_add_7_25_groupi_n_6423 ,csa_tree_add_7_25_groupi_n_6311);
  xnor csa_tree_add_7_25_groupi_g14595__9945(csa_tree_add_7_25_groupi_n_6505 ,csa_tree_add_7_25_groupi_n_6420 ,csa_tree_add_7_25_groupi_n_6304);
  xnor csa_tree_add_7_25_groupi_g14596__2883(csa_tree_add_7_25_groupi_n_6504 ,csa_tree_add_7_25_groupi_n_6422 ,csa_tree_add_7_25_groupi_n_6305);
  xnor csa_tree_add_7_25_groupi_g14597__2346(csa_tree_add_7_25_groupi_n_6503 ,csa_tree_add_7_25_groupi_n_6359 ,csa_tree_add_7_25_groupi_n_6408);
  xnor csa_tree_add_7_25_groupi_g14598__1666(csa_tree_add_7_25_groupi_n_6501 ,csa_tree_add_7_25_groupi_n_6360 ,csa_tree_add_7_25_groupi_n_6406);
  xnor csa_tree_add_7_25_groupi_g14599__7410(csa_tree_add_7_25_groupi_n_6499 ,csa_tree_add_7_25_groupi_n_6362 ,csa_tree_add_7_25_groupi_n_6405);
  xnor csa_tree_add_7_25_groupi_g14600__6417(csa_tree_add_7_25_groupi_n_6497 ,csa_tree_add_7_25_groupi_n_6424 ,csa_tree_add_7_25_groupi_n_6313);
  xnor csa_tree_add_7_25_groupi_g14601__5477(csa_tree_add_7_25_groupi_n_6495 ,csa_tree_add_7_25_groupi_n_6426 ,csa_tree_add_7_25_groupi_n_6312);
  xnor csa_tree_add_7_25_groupi_g14602__2398(csa_tree_add_7_25_groupi_n_6493 ,csa_tree_add_7_25_groupi_n_6425 ,csa_tree_add_7_25_groupi_n_6307);
  and csa_tree_add_7_25_groupi_g14603__5107(csa_tree_add_7_25_groupi_n_6483 ,csa_tree_add_7_25_groupi_n_6417 ,csa_tree_add_7_25_groupi_n_6356);
  or csa_tree_add_7_25_groupi_g14604__6260(csa_tree_add_7_25_groupi_n_6482 ,csa_tree_add_7_25_groupi_n_3410 ,csa_tree_add_7_25_groupi_n_6445);
  or csa_tree_add_7_25_groupi_g14605__4319(csa_tree_add_7_25_groupi_n_6481 ,csa_tree_add_7_25_groupi_n_6416 ,csa_tree_add_7_25_groupi_n_6355);
  and csa_tree_add_7_25_groupi_g14606__8428(csa_tree_add_7_25_groupi_n_6480 ,csa_tree_add_7_25_groupi_n_6422 ,csa_tree_add_7_25_groupi_n_6288);
  and csa_tree_add_7_25_groupi_g14607__5526(csa_tree_add_7_25_groupi_n_6479 ,csa_tree_add_7_25_groupi_n_6416 ,csa_tree_add_7_25_groupi_n_6355);
  and csa_tree_add_7_25_groupi_g14608__6783(csa_tree_add_7_25_groupi_n_6478 ,csa_tree_add_7_25_groupi_n_6421 ,csa_tree_add_7_25_groupi_n_6296);
  and csa_tree_add_7_25_groupi_g14609__3680(csa_tree_add_7_25_groupi_n_6477 ,csa_tree_add_7_25_groupi_n_6420 ,csa_tree_add_7_25_groupi_n_6292);
  and csa_tree_add_7_25_groupi_g14610__1617(csa_tree_add_7_25_groupi_n_6476 ,csa_tree_add_7_25_groupi_n_6423 ,csa_tree_add_7_25_groupi_n_6300);
  or csa_tree_add_7_25_groupi_g14611__2802(csa_tree_add_7_25_groupi_n_6475 ,csa_tree_add_7_25_groupi_n_6417 ,csa_tree_add_7_25_groupi_n_6356);
  and csa_tree_add_7_25_groupi_g14612__1705(csa_tree_add_7_25_groupi_n_6474 ,csa_tree_add_7_25_groupi_n_6418 ,csa_tree_add_7_25_groupi_n_6358);
  or csa_tree_add_7_25_groupi_g14613__5122(csa_tree_add_7_25_groupi_n_6473 ,csa_tree_add_7_25_groupi_n_6418 ,csa_tree_add_7_25_groupi_n_6358);
  or csa_tree_add_7_25_groupi_g14614__8246(csa_tree_add_7_25_groupi_n_6472 ,csa_tree_add_7_25_groupi_n_6357 ,csa_tree_add_7_25_groupi_n_6419);
  and csa_tree_add_7_25_groupi_g14615__7098(csa_tree_add_7_25_groupi_n_6471 ,csa_tree_add_7_25_groupi_n_6357 ,csa_tree_add_7_25_groupi_n_6419);
  or csa_tree_add_7_25_groupi_g14616__6131(csa_tree_add_7_25_groupi_n_6485 ,csa_tree_add_7_25_groupi_n_6397 ,csa_tree_add_7_25_groupi_n_6440);
  and csa_tree_add_7_25_groupi_g14617__1881(csa_tree_add_7_25_groupi_n_6484 ,csa_tree_add_7_25_groupi_n_2449 ,csa_tree_add_7_25_groupi_n_6441);
  not csa_tree_add_7_25_groupi_g14618(csa_tree_add_7_25_groupi_n_6469 ,csa_tree_add_7_25_groupi_n_6470);
  not csa_tree_add_7_25_groupi_g14619(csa_tree_add_7_25_groupi_n_6467 ,csa_tree_add_7_25_groupi_n_6468);
  not csa_tree_add_7_25_groupi_g14620(csa_tree_add_7_25_groupi_n_6464 ,csa_tree_add_7_25_groupi_n_6465);
  or csa_tree_add_7_25_groupi_g14621__5115(csa_tree_add_7_25_groupi_n_6462 ,csa_tree_add_7_25_groupi_n_3325 ,csa_tree_add_7_25_groupi_n_6446);
  or csa_tree_add_7_25_groupi_g14622__7482(csa_tree_add_7_25_groupi_n_6461 ,csa_tree_add_7_25_groupi_n_3762 ,csa_tree_add_7_25_groupi_n_6443);
  or csa_tree_add_7_25_groupi_g14623__4733(csa_tree_add_7_25_groupi_n_6460 ,csa_tree_add_7_25_groupi_n_3765 ,csa_tree_add_7_25_groupi_n_6444);
  or csa_tree_add_7_25_groupi_g14624__6161(csa_tree_add_7_25_groupi_n_6459 ,csa_tree_add_7_25_groupi_n_3767 ,csa_tree_add_7_25_groupi_n_6447);
  and csa_tree_add_7_25_groupi_g14625__9315(csa_tree_add_7_25_groupi_n_6458 ,csa_tree_add_7_25_groupi_n_6425 ,csa_tree_add_7_25_groupi_n_6282);
  or csa_tree_add_7_25_groupi_g14626__9945(csa_tree_add_7_25_groupi_n_6457 ,csa_tree_add_7_25_groupi_n_3407 ,csa_tree_add_7_25_groupi_n_6448);
  and csa_tree_add_7_25_groupi_g14627__2883(csa_tree_add_7_25_groupi_n_6456 ,csa_tree_add_7_25_groupi_n_6426 ,csa_tree_add_7_25_groupi_n_6283);
  or csa_tree_add_7_25_groupi_g14628__2346(csa_tree_add_7_25_groupi_n_6455 ,csa_tree_add_7_25_groupi_n_3348 ,csa_tree_add_7_25_groupi_n_6442);
  and csa_tree_add_7_25_groupi_g14629__1666(csa_tree_add_7_25_groupi_n_6454 ,csa_tree_add_7_25_groupi_n_6424 ,csa_tree_add_7_25_groupi_n_6271);
  and csa_tree_add_7_25_groupi_g14630__7410(csa_tree_add_7_25_groupi_n_6453 ,csa_tree_add_7_25_groupi_n_6427 ,csa_tree_add_7_25_groupi_n_6268);
  or csa_tree_add_7_25_groupi_g14631__6417(csa_tree_add_7_25_groupi_n_6470 ,csa_tree_add_7_25_groupi_n_6367 ,csa_tree_add_7_25_groupi_n_6436);
  or csa_tree_add_7_25_groupi_g14632__5477(csa_tree_add_7_25_groupi_n_6468 ,csa_tree_add_7_25_groupi_n_6438 ,csa_tree_add_7_25_groupi_n_6374);
  or csa_tree_add_7_25_groupi_g14633__2398(csa_tree_add_7_25_groupi_n_6466 ,csa_tree_add_7_25_groupi_n_6439 ,csa_tree_add_7_25_groupi_n_6363);
  or csa_tree_add_7_25_groupi_g14634__5107(csa_tree_add_7_25_groupi_n_6465 ,csa_tree_add_7_25_groupi_n_6437 ,csa_tree_add_7_25_groupi_n_6372);
  xnor csa_tree_add_7_25_groupi_g14635__6260(csa_tree_add_7_25_groupi_n_6463 ,csa_tree_add_7_25_groupi_n_6401 ,csa_tree_add_7_25_groupi_n_2563);
  nor csa_tree_add_7_25_groupi_g14636__4319(csa_tree_add_7_25_groupi_n_6448 ,csa_tree_add_7_25_groupi_n_2108 ,csa_tree_add_7_25_groupi_n_6382);
  nor csa_tree_add_7_25_groupi_g14637__8428(csa_tree_add_7_25_groupi_n_6447 ,csa_tree_add_7_25_groupi_n_2162 ,csa_tree_add_7_25_groupi_n_1137);
  nor csa_tree_add_7_25_groupi_g14638__5526(csa_tree_add_7_25_groupi_n_6446 ,csa_tree_add_7_25_groupi_n_2153 ,csa_tree_add_7_25_groupi_n_1264);
  nor csa_tree_add_7_25_groupi_g14639__6783(csa_tree_add_7_25_groupi_n_6445 ,csa_tree_add_7_25_groupi_n_2192 ,csa_tree_add_7_25_groupi_n_1137);
  nor csa_tree_add_7_25_groupi_g14640__3680(csa_tree_add_7_25_groupi_n_6444 ,csa_tree_add_7_25_groupi_n_2066 ,csa_tree_add_7_25_groupi_n_1264);
  nor csa_tree_add_7_25_groupi_g14641__1617(csa_tree_add_7_25_groupi_n_6443 ,csa_tree_add_7_25_groupi_n_2036 ,csa_tree_add_7_25_groupi_n_1265);
  nor csa_tree_add_7_25_groupi_g14642__2802(csa_tree_add_7_25_groupi_n_6442 ,csa_tree_add_7_25_groupi_n_2180 ,csa_tree_add_7_25_groupi_n_1265);
  or csa_tree_add_7_25_groupi_g14643__1705(csa_tree_add_7_25_groupi_n_6441 ,csa_tree_add_7_25_groupi_n_2436 ,csa_tree_add_7_25_groupi_n_6401);
  and csa_tree_add_7_25_groupi_g14644__5122(csa_tree_add_7_25_groupi_n_6440 ,csa_tree_add_7_25_groupi_n_6396 ,csa_tree_add_7_25_groupi_n_6400);
  and csa_tree_add_7_25_groupi_g14645__8246(csa_tree_add_7_25_groupi_n_6439 ,csa_tree_add_7_25_groupi_n_6364 ,csa_tree_add_7_25_groupi_n_6361);
  and csa_tree_add_7_25_groupi_g14646__7098(csa_tree_add_7_25_groupi_n_6438 ,csa_tree_add_7_25_groupi_n_6375 ,csa_tree_add_7_25_groupi_n_6362);
  and csa_tree_add_7_25_groupi_g14647__6131(csa_tree_add_7_25_groupi_n_6437 ,csa_tree_add_7_25_groupi_n_6360 ,csa_tree_add_7_25_groupi_n_6373);
  and csa_tree_add_7_25_groupi_g14648__1881(csa_tree_add_7_25_groupi_n_6436 ,csa_tree_add_7_25_groupi_n_6366 ,csa_tree_add_7_25_groupi_n_6359);
  nor csa_tree_add_7_25_groupi_g14649__5115(csa_tree_add_7_25_groupi_n_6435 ,csa_tree_add_7_25_groupi_n_3880 ,csa_tree_add_7_25_groupi_n_6378);
  nor csa_tree_add_7_25_groupi_g14650__7482(csa_tree_add_7_25_groupi_n_6434 ,csa_tree_add_7_25_groupi_n_4009 ,csa_tree_add_7_25_groupi_n_6390);
  nor csa_tree_add_7_25_groupi_g14651__4733(csa_tree_add_7_25_groupi_n_6433 ,csa_tree_add_7_25_groupi_n_3912 ,csa_tree_add_7_25_groupi_n_6380);
  nor csa_tree_add_7_25_groupi_g14652__6161(csa_tree_add_7_25_groupi_n_6432 ,csa_tree_add_7_25_groupi_n_3903 ,csa_tree_add_7_25_groupi_n_6381);
  nor csa_tree_add_7_25_groupi_g14653__9315(csa_tree_add_7_25_groupi_n_6431 ,csa_tree_add_7_25_groupi_n_4021 ,csa_tree_add_7_25_groupi_n_6383);
  nor csa_tree_add_7_25_groupi_g14654__9945(csa_tree_add_7_25_groupi_n_6430 ,csa_tree_add_7_25_groupi_n_3491 ,csa_tree_add_7_25_groupi_n_6369);
  nor csa_tree_add_7_25_groupi_g14655__2883(csa_tree_add_7_25_groupi_n_6429 ,csa_tree_add_7_25_groupi_n_3936 ,csa_tree_add_7_25_groupi_n_6379);
  nor csa_tree_add_7_25_groupi_g14656__2346(csa_tree_add_7_25_groupi_n_6428 ,csa_tree_add_7_25_groupi_n_3909 ,csa_tree_add_7_25_groupi_n_6398);
  or csa_tree_add_7_25_groupi_g14657__1666(csa_tree_add_7_25_groupi_n_6452 ,csa_tree_add_7_25_groupi_n_6187 ,csa_tree_add_7_25_groupi_n_6385);
  or csa_tree_add_7_25_groupi_g14658__7410(csa_tree_add_7_25_groupi_n_6451 ,csa_tree_add_7_25_groupi_n_6195 ,csa_tree_add_7_25_groupi_n_6395);
  or csa_tree_add_7_25_groupi_g14659__6417(csa_tree_add_7_25_groupi_n_6450 ,csa_tree_add_7_25_groupi_n_6192 ,csa_tree_add_7_25_groupi_n_6394);
  or csa_tree_add_7_25_groupi_g14660__5477(csa_tree_add_7_25_groupi_n_6449 ,csa_tree_add_7_25_groupi_n_6189 ,csa_tree_add_7_25_groupi_n_6391);
  xnor csa_tree_add_7_25_groupi_g14661__2398(out2[15] ,csa_tree_add_7_25_groupi_n_6285 ,csa_tree_add_7_25_groupi_n_6310);
  xnor csa_tree_add_7_25_groupi_g14662__5107(csa_tree_add_7_25_groupi_n_6414 ,csa_tree_add_7_25_groupi_n_6258 ,csa_tree_add_7_25_groupi_n_6320);
  xnor csa_tree_add_7_25_groupi_g14663__6260(csa_tree_add_7_25_groupi_n_6413 ,csa_tree_add_7_25_groupi_n_6257 ,csa_tree_add_7_25_groupi_n_6317);
  xnor csa_tree_add_7_25_groupi_g14664__4319(csa_tree_add_7_25_groupi_n_6412 ,csa_tree_add_7_25_groupi_n_6259 ,csa_tree_add_7_25_groupi_n_6319);
  xnor csa_tree_add_7_25_groupi_g14665__8428(csa_tree_add_7_25_groupi_n_6411 ,csa_tree_add_7_25_groupi_n_6332 ,csa_tree_add_7_25_groupi_n_6261);
  xnor csa_tree_add_7_25_groupi_g14666__5526(csa_tree_add_7_25_groupi_n_6410 ,csa_tree_add_7_25_groupi_n_6315 ,csa_tree_add_7_25_groupi_n_6260);
  xnor csa_tree_add_7_25_groupi_g14667__6783(csa_tree_add_7_25_groupi_n_6409 ,csa_tree_add_7_25_groupi_n_6266 ,csa_tree_add_7_25_groupi_n_6318);
  xnor csa_tree_add_7_25_groupi_g14668__3680(csa_tree_add_7_25_groupi_n_6408 ,csa_tree_add_7_25_groupi_n_6328 ,csa_tree_add_7_25_groupi_n_6218);
  xnor csa_tree_add_7_25_groupi_g14669__1617(csa_tree_add_7_25_groupi_n_6407 ,csa_tree_add_7_25_groupi_n_6331 ,csa_tree_add_7_25_groupi_n_6226);
  xnor csa_tree_add_7_25_groupi_g14670__2802(csa_tree_add_7_25_groupi_n_6406 ,csa_tree_add_7_25_groupi_n_6330 ,csa_tree_add_7_25_groupi_n_6216);
  xnor csa_tree_add_7_25_groupi_g14671__1705(csa_tree_add_7_25_groupi_n_6405 ,csa_tree_add_7_25_groupi_n_6322 ,csa_tree_add_7_25_groupi_n_6220);
  xnor csa_tree_add_7_25_groupi_g14672__5122(csa_tree_add_7_25_groupi_n_6404 ,csa_tree_add_7_25_groupi_n_6326 ,csa_tree_add_7_25_groupi_n_6263);
  xnor csa_tree_add_7_25_groupi_g14673__8246(csa_tree_add_7_25_groupi_n_6403 ,csa_tree_add_7_25_groupi_n_6241 ,csa_tree_add_7_25_groupi_n_6309);
  xnor csa_tree_add_7_25_groupi_g14674__7098(csa_tree_add_7_25_groupi_n_6402 ,csa_tree_add_7_25_groupi_n_6265 ,csa_tree_add_7_25_groupi_n_6324);
  xnor csa_tree_add_7_25_groupi_g14675__6131(csa_tree_add_7_25_groupi_n_6427 ,csa_tree_add_7_25_groupi_n_6344 ,in3[11]);
  xnor csa_tree_add_7_25_groupi_g14676__1881(csa_tree_add_7_25_groupi_n_6426 ,csa_tree_add_7_25_groupi_n_6340 ,in3[20]);
  xnor csa_tree_add_7_25_groupi_g14677__5115(csa_tree_add_7_25_groupi_n_6425 ,csa_tree_add_7_25_groupi_n_6343 ,in3[23]);
  xnor csa_tree_add_7_25_groupi_g14678__7482(csa_tree_add_7_25_groupi_n_6424 ,csa_tree_add_7_25_groupi_n_6341 ,in3[17]);
  xnor csa_tree_add_7_25_groupi_g14679__4733(csa_tree_add_7_25_groupi_n_6423 ,csa_tree_add_7_25_groupi_n_6337 ,in3[14]);
  xnor csa_tree_add_7_25_groupi_g14680__6161(csa_tree_add_7_25_groupi_n_6422 ,csa_tree_add_7_25_groupi_n_6342 ,in3[8]);
  xnor csa_tree_add_7_25_groupi_g14681__9315(csa_tree_add_7_25_groupi_n_6421 ,csa_tree_add_7_25_groupi_n_6338 ,in3[2]);
  xnor csa_tree_add_7_25_groupi_g14682__9945(csa_tree_add_7_25_groupi_n_6420 ,csa_tree_add_7_25_groupi_n_6339 ,in3[5]);
  xnor csa_tree_add_7_25_groupi_g14683__2883(csa_tree_add_7_25_groupi_n_6419 ,csa_tree_add_7_25_groupi_n_6335 ,csa_tree_add_7_25_groupi_n_6207);
  xnor csa_tree_add_7_25_groupi_g14684__2346(csa_tree_add_7_25_groupi_n_6418 ,csa_tree_add_7_25_groupi_n_6334 ,csa_tree_add_7_25_groupi_n_6206);
  xnor csa_tree_add_7_25_groupi_g14685__1666(csa_tree_add_7_25_groupi_n_6417 ,csa_tree_add_7_25_groupi_n_6336 ,csa_tree_add_7_25_groupi_n_6205);
  xnor csa_tree_add_7_25_groupi_g14686__7410(csa_tree_add_7_25_groupi_n_6416 ,csa_tree_add_7_25_groupi_n_6333 ,csa_tree_add_7_25_groupi_n_6204);
  and csa_tree_add_7_25_groupi_g14687__6417(csa_tree_add_7_25_groupi_n_6399 ,csa_tree_add_7_25_groupi_n_6315 ,csa_tree_add_7_25_groupi_n_6260);
  or csa_tree_add_7_25_groupi_g14688__5477(csa_tree_add_7_25_groupi_n_6398 ,csa_tree_add_7_25_groupi_n_3760 ,csa_tree_add_7_25_groupi_n_6351);
  and csa_tree_add_7_25_groupi_g14689__2398(csa_tree_add_7_25_groupi_n_6397 ,csa_tree_add_7_25_groupi_n_6258 ,csa_tree_add_7_25_groupi_n_6320);
  or csa_tree_add_7_25_groupi_g14690__5107(csa_tree_add_7_25_groupi_n_6396 ,csa_tree_add_7_25_groupi_n_6258 ,csa_tree_add_7_25_groupi_n_6320);
  and csa_tree_add_7_25_groupi_g14691__6260(csa_tree_add_7_25_groupi_n_6395 ,csa_tree_add_7_25_groupi_n_6333 ,csa_tree_add_7_25_groupi_n_6194);
  and csa_tree_add_7_25_groupi_g14692__4319(csa_tree_add_7_25_groupi_n_6394 ,csa_tree_add_7_25_groupi_n_6336 ,csa_tree_add_7_25_groupi_n_6191);
  or csa_tree_add_7_25_groupi_g14693__8428(csa_tree_add_7_25_groupi_n_6393 ,csa_tree_add_7_25_groupi_n_6259 ,csa_tree_add_7_25_groupi_n_6319);
  and csa_tree_add_7_25_groupi_g14694__5526(csa_tree_add_7_25_groupi_n_6392 ,csa_tree_add_7_25_groupi_n_6259 ,csa_tree_add_7_25_groupi_n_6319);
  and csa_tree_add_7_25_groupi_g14695__6783(csa_tree_add_7_25_groupi_n_6391 ,csa_tree_add_7_25_groupi_n_6335 ,csa_tree_add_7_25_groupi_n_6190);
  or csa_tree_add_7_25_groupi_g14696__3680(csa_tree_add_7_25_groupi_n_6390 ,csa_tree_add_7_25_groupi_n_3392 ,csa_tree_add_7_25_groupi_n_6345);
  or csa_tree_add_7_25_groupi_g14697__1617(csa_tree_add_7_25_groupi_n_6389 ,csa_tree_add_7_25_groupi_n_6315 ,csa_tree_add_7_25_groupi_n_6260);
  or csa_tree_add_7_25_groupi_g14698__2802(csa_tree_add_7_25_groupi_n_6388 ,csa_tree_add_7_25_groupi_n_6266 ,csa_tree_add_7_25_groupi_n_6318);
  and csa_tree_add_7_25_groupi_g14699__1705(csa_tree_add_7_25_groupi_n_6387 ,csa_tree_add_7_25_groupi_n_6332 ,csa_tree_add_7_25_groupi_n_6261);
  or csa_tree_add_7_25_groupi_g14700__5122(csa_tree_add_7_25_groupi_n_6386 ,csa_tree_add_7_25_groupi_n_6332 ,csa_tree_add_7_25_groupi_n_6261);
  and csa_tree_add_7_25_groupi_g14701__8246(csa_tree_add_7_25_groupi_n_6385 ,csa_tree_add_7_25_groupi_n_6334 ,csa_tree_add_7_25_groupi_n_6186);
  and csa_tree_add_7_25_groupi_g14702__7098(csa_tree_add_7_25_groupi_n_6384 ,csa_tree_add_7_25_groupi_n_6266 ,csa_tree_add_7_25_groupi_n_6318);
  or csa_tree_add_7_25_groupi_g14703__6131(csa_tree_add_7_25_groupi_n_6383 ,csa_tree_add_7_25_groupi_n_3395 ,csa_tree_add_7_25_groupi_n_6348);
  and csa_tree_add_7_25_groupi_g14704__1881(csa_tree_add_7_25_groupi_n_6401 ,csa_tree_add_7_25_groupi_n_2478 ,csa_tree_add_7_25_groupi_n_6353);
  or csa_tree_add_7_25_groupi_g14705__5115(csa_tree_add_7_25_groupi_n_6400 ,csa_tree_add_7_25_groupi_n_6354 ,csa_tree_add_7_25_groupi_n_6298);
  or csa_tree_add_7_25_groupi_g14706__7482(csa_tree_add_7_25_groupi_n_6381 ,csa_tree_add_7_25_groupi_n_3759 ,csa_tree_add_7_25_groupi_n_6350);
  or csa_tree_add_7_25_groupi_g14707__4733(csa_tree_add_7_25_groupi_n_6380 ,csa_tree_add_7_25_groupi_n_3755 ,csa_tree_add_7_25_groupi_n_6349);
  or csa_tree_add_7_25_groupi_g14708__6161(csa_tree_add_7_25_groupi_n_6379 ,csa_tree_add_7_25_groupi_n_3758 ,csa_tree_add_7_25_groupi_n_6347);
  or csa_tree_add_7_25_groupi_g14709__9315(csa_tree_add_7_25_groupi_n_6378 ,csa_tree_add_7_25_groupi_n_3757 ,csa_tree_add_7_25_groupi_n_6346);
  nor csa_tree_add_7_25_groupi_g14710__9945(csa_tree_add_7_25_groupi_n_6377 ,csa_tree_add_7_25_groupi_n_6326 ,csa_tree_add_7_25_groupi_n_6262);
  or csa_tree_add_7_25_groupi_g14711__2883(csa_tree_add_7_25_groupi_n_6376 ,csa_tree_add_7_25_groupi_n_6325 ,csa_tree_add_7_25_groupi_n_6263);
  or csa_tree_add_7_25_groupi_g14712__2346(csa_tree_add_7_25_groupi_n_6375 ,csa_tree_add_7_25_groupi_n_6322 ,csa_tree_add_7_25_groupi_n_6219);
  nor csa_tree_add_7_25_groupi_g14713__1666(csa_tree_add_7_25_groupi_n_6374 ,csa_tree_add_7_25_groupi_n_6321 ,csa_tree_add_7_25_groupi_n_6220);
  or csa_tree_add_7_25_groupi_g14714__7410(csa_tree_add_7_25_groupi_n_6373 ,csa_tree_add_7_25_groupi_n_6330 ,csa_tree_add_7_25_groupi_n_6215);
  nor csa_tree_add_7_25_groupi_g14715__6417(csa_tree_add_7_25_groupi_n_6372 ,csa_tree_add_7_25_groupi_n_6329 ,csa_tree_add_7_25_groupi_n_6216);
  nor csa_tree_add_7_25_groupi_g14716__5477(csa_tree_add_7_25_groupi_n_6371 ,csa_tree_add_7_25_groupi_n_6264 ,csa_tree_add_7_25_groupi_n_6324);
  or csa_tree_add_7_25_groupi_g14717__2398(csa_tree_add_7_25_groupi_n_6370 ,csa_tree_add_7_25_groupi_n_6265 ,csa_tree_add_7_25_groupi_n_6323);
  or csa_tree_add_7_25_groupi_g14718__5107(csa_tree_add_7_25_groupi_n_6369 ,csa_tree_add_7_25_groupi_n_3330 ,csa_tree_add_7_25_groupi_n_6352);
  or csa_tree_add_7_25_groupi_g14719__6260(csa_tree_add_7_25_groupi_n_6368 ,csa_tree_add_7_25_groupi_n_6257 ,csa_tree_add_7_25_groupi_n_6316);
  nor csa_tree_add_7_25_groupi_g14720__4319(csa_tree_add_7_25_groupi_n_6367 ,csa_tree_add_7_25_groupi_n_6327 ,csa_tree_add_7_25_groupi_n_6218);
  or csa_tree_add_7_25_groupi_g14721__8428(csa_tree_add_7_25_groupi_n_6366 ,csa_tree_add_7_25_groupi_n_6328 ,csa_tree_add_7_25_groupi_n_6217);
  nor csa_tree_add_7_25_groupi_g14722__5526(csa_tree_add_7_25_groupi_n_6365 ,csa_tree_add_7_25_groupi_n_6256 ,csa_tree_add_7_25_groupi_n_6317);
  or csa_tree_add_7_25_groupi_g14723__6783(csa_tree_add_7_25_groupi_n_6364 ,csa_tree_add_7_25_groupi_n_6331 ,csa_tree_add_7_25_groupi_n_6226);
  and csa_tree_add_7_25_groupi_g14724__3680(csa_tree_add_7_25_groupi_n_6363 ,csa_tree_add_7_25_groupi_n_6331 ,csa_tree_add_7_25_groupi_n_6226);
  xnor csa_tree_add_7_25_groupi_g14725__1617(csa_tree_add_7_25_groupi_n_6382 ,csa_tree_add_7_25_groupi_n_6303 ,csa_tree_add_7_25_groupi_n_2564);
  and csa_tree_add_7_25_groupi_g14726__2802(csa_tree_add_7_25_groupi_n_6354 ,csa_tree_add_7_25_groupi_n_6299 ,csa_tree_add_7_25_groupi_n_6285);
  or csa_tree_add_7_25_groupi_g14727__1705(csa_tree_add_7_25_groupi_n_6353 ,csa_tree_add_7_25_groupi_n_2452 ,csa_tree_add_7_25_groupi_n_6303);
  nor csa_tree_add_7_25_groupi_g14728__5122(csa_tree_add_7_25_groupi_n_6352 ,csa_tree_add_7_25_groupi_n_2187 ,csa_tree_add_7_25_groupi_n_1277);
  nor csa_tree_add_7_25_groupi_g14729__8246(csa_tree_add_7_25_groupi_n_6351 ,csa_tree_add_7_25_groupi_n_2030 ,csa_tree_add_7_25_groupi_n_1268);
  nor csa_tree_add_7_25_groupi_g14730__7098(csa_tree_add_7_25_groupi_n_6350 ,csa_tree_add_7_25_groupi_n_2045 ,csa_tree_add_7_25_groupi_n_1267);
  nor csa_tree_add_7_25_groupi_g14731__6131(csa_tree_add_7_25_groupi_n_6349 ,csa_tree_add_7_25_groupi_n_2057 ,csa_tree_add_7_25_groupi_n_1267);
  nor csa_tree_add_7_25_groupi_g14732__1881(csa_tree_add_7_25_groupi_n_6348 ,csa_tree_add_7_25_groupi_n_2139 ,csa_tree_add_7_25_groupi_n_1276);
  nor csa_tree_add_7_25_groupi_g14733__5115(csa_tree_add_7_25_groupi_n_6347 ,csa_tree_add_7_25_groupi_n_2160 ,csa_tree_add_7_25_groupi_n_1276);
  nor csa_tree_add_7_25_groupi_g14734__7482(csa_tree_add_7_25_groupi_n_6346 ,csa_tree_add_7_25_groupi_n_2106 ,csa_tree_add_7_25_groupi_n_1268);
  nor csa_tree_add_7_25_groupi_g14735__4733(csa_tree_add_7_25_groupi_n_6345 ,csa_tree_add_7_25_groupi_n_2127 ,csa_tree_add_7_25_groupi_n_1277);
  nor csa_tree_add_7_25_groupi_g14736__6161(csa_tree_add_7_25_groupi_n_6344 ,csa_tree_add_7_25_groupi_n_3908 ,csa_tree_add_7_25_groupi_n_6277);
  nor csa_tree_add_7_25_groupi_g14737__9315(csa_tree_add_7_25_groupi_n_6343 ,csa_tree_add_7_25_groupi_n_3858 ,csa_tree_add_7_25_groupi_n_6281);
  nor csa_tree_add_7_25_groupi_g14738__9945(csa_tree_add_7_25_groupi_n_6342 ,csa_tree_add_7_25_groupi_n_4003 ,csa_tree_add_7_25_groupi_n_6293);
  nor csa_tree_add_7_25_groupi_g14739__2883(csa_tree_add_7_25_groupi_n_6341 ,csa_tree_add_7_25_groupi_n_3881 ,csa_tree_add_7_25_groupi_n_6279);
  nor csa_tree_add_7_25_groupi_g14740__2346(csa_tree_add_7_25_groupi_n_6340 ,csa_tree_add_7_25_groupi_n_3892 ,csa_tree_add_7_25_groupi_n_6280);
  nor csa_tree_add_7_25_groupi_g14741__1666(csa_tree_add_7_25_groupi_n_6339 ,csa_tree_add_7_25_groupi_n_4092 ,csa_tree_add_7_25_groupi_n_6286);
  nor csa_tree_add_7_25_groupi_g14742__7410(csa_tree_add_7_25_groupi_n_6338 ,csa_tree_add_7_25_groupi_n_3474 ,csa_tree_add_7_25_groupi_n_6269);
  nor csa_tree_add_7_25_groupi_g14743__6417(csa_tree_add_7_25_groupi_n_6337 ,csa_tree_add_7_25_groupi_n_3863 ,csa_tree_add_7_25_groupi_n_6278);
  or csa_tree_add_7_25_groupi_g14744__5477(csa_tree_add_7_25_groupi_n_6362 ,csa_tree_add_7_25_groupi_n_6085 ,csa_tree_add_7_25_groupi_n_6276);
  or csa_tree_add_7_25_groupi_g14745__2398(csa_tree_add_7_25_groupi_n_6361 ,csa_tree_add_7_25_groupi_n_6099 ,csa_tree_add_7_25_groupi_n_6294);
  or csa_tree_add_7_25_groupi_g14746__5107(csa_tree_add_7_25_groupi_n_6360 ,csa_tree_add_7_25_groupi_n_6078 ,csa_tree_add_7_25_groupi_n_6273);
  or csa_tree_add_7_25_groupi_g14747__6260(csa_tree_add_7_25_groupi_n_6359 ,csa_tree_add_7_25_groupi_n_6073 ,csa_tree_add_7_25_groupi_n_6270);
  or csa_tree_add_7_25_groupi_g14748__4319(csa_tree_add_7_25_groupi_n_6358 ,csa_tree_add_7_25_groupi_n_6090 ,csa_tree_add_7_25_groupi_n_6287);
  or csa_tree_add_7_25_groupi_g14749__8428(csa_tree_add_7_25_groupi_n_6357 ,csa_tree_add_7_25_groupi_n_6093 ,csa_tree_add_7_25_groupi_n_6290);
  or csa_tree_add_7_25_groupi_g14750__5526(csa_tree_add_7_25_groupi_n_6356 ,csa_tree_add_7_25_groupi_n_6095 ,csa_tree_add_7_25_groupi_n_6291);
  or csa_tree_add_7_25_groupi_g14751__6783(csa_tree_add_7_25_groupi_n_6355 ,csa_tree_add_7_25_groupi_n_6101 ,csa_tree_add_7_25_groupi_n_6295);
  not csa_tree_add_7_25_groupi_g14752(csa_tree_add_7_25_groupi_n_6329 ,csa_tree_add_7_25_groupi_n_6330);
  not csa_tree_add_7_25_groupi_g14753(csa_tree_add_7_25_groupi_n_6327 ,csa_tree_add_7_25_groupi_n_6328);
  not csa_tree_add_7_25_groupi_g14754(csa_tree_add_7_25_groupi_n_6325 ,csa_tree_add_7_25_groupi_n_6326);
  not csa_tree_add_7_25_groupi_g14755(csa_tree_add_7_25_groupi_n_6323 ,csa_tree_add_7_25_groupi_n_6324);
  not csa_tree_add_7_25_groupi_g14756(csa_tree_add_7_25_groupi_n_6321 ,csa_tree_add_7_25_groupi_n_6322);
  not csa_tree_add_7_25_groupi_g14757(csa_tree_add_7_25_groupi_n_6316 ,csa_tree_add_7_25_groupi_n_6317);
  xnor csa_tree_add_7_25_groupi_g14758__3680(out2[14] ,csa_tree_add_7_25_groupi_n_6202 ,csa_tree_add_7_25_groupi_n_6208);
  xnor csa_tree_add_7_25_groupi_g14759__1617(csa_tree_add_7_25_groupi_n_6313 ,csa_tree_add_7_25_groupi_n_6183 ,csa_tree_add_7_25_groupi_n_6214);
  xnor csa_tree_add_7_25_groupi_g14760__2802(csa_tree_add_7_25_groupi_n_6312 ,csa_tree_add_7_25_groupi_n_6185 ,csa_tree_add_7_25_groupi_n_6212);
  xnor csa_tree_add_7_25_groupi_g14761__1705(csa_tree_add_7_25_groupi_n_6311 ,csa_tree_add_7_25_groupi_n_6223 ,csa_tree_add_7_25_groupi_n_6181);
  xnor csa_tree_add_7_25_groupi_g14762__5122(csa_tree_add_7_25_groupi_n_6310 ,csa_tree_add_7_25_groupi_n_6163 ,csa_tree_add_7_25_groupi_n_6224);
  xnor csa_tree_add_7_25_groupi_g14763__8246(csa_tree_add_7_25_groupi_n_6309 ,csa_tree_add_7_25_groupi_n_6203 ,csa_tree_add_7_25_groupi_n_6110);
  xnor csa_tree_add_7_25_groupi_g14764__7098(csa_tree_add_7_25_groupi_n_6308 ,csa_tree_add_7_25_groupi_n_6164 ,csa_tree_add_7_25_groupi_n_6222);
  xnor csa_tree_add_7_25_groupi_g14765__6131(csa_tree_add_7_25_groupi_n_6307 ,csa_tree_add_7_25_groupi_n_6180 ,csa_tree_add_7_25_groupi_n_6228);
  xnor csa_tree_add_7_25_groupi_g14766__1881(csa_tree_add_7_25_groupi_n_6306 ,csa_tree_add_7_25_groupi_n_6165 ,csa_tree_add_7_25_groupi_n_6225);
  xnor csa_tree_add_7_25_groupi_g14767__5115(csa_tree_add_7_25_groupi_n_6305 ,csa_tree_add_7_25_groupi_n_6162 ,csa_tree_add_7_25_groupi_n_6210);
  xnor csa_tree_add_7_25_groupi_g14768__7482(csa_tree_add_7_25_groupi_n_6304 ,csa_tree_add_7_25_groupi_n_6161 ,csa_tree_add_7_25_groupi_n_6221);
  xnor csa_tree_add_7_25_groupi_g14769__4733(csa_tree_add_7_25_groupi_n_6336 ,csa_tree_add_7_25_groupi_n_6237 ,in3[5]);
  xnor csa_tree_add_7_25_groupi_g14770__6161(csa_tree_add_7_25_groupi_n_6335 ,csa_tree_add_7_25_groupi_n_6243 ,in3[11]);
  xnor csa_tree_add_7_25_groupi_g14771__9315(csa_tree_add_7_25_groupi_n_6334 ,csa_tree_add_7_25_groupi_n_6238 ,in3[8]);
  xnor csa_tree_add_7_25_groupi_g14772__9945(csa_tree_add_7_25_groupi_n_6333 ,csa_tree_add_7_25_groupi_n_6244 ,in3[2]);
  xnor csa_tree_add_7_25_groupi_g14773__2883(csa_tree_add_7_25_groupi_n_6332 ,csa_tree_add_7_25_groupi_n_6229 ,csa_tree_add_7_25_groupi_n_6118);
  xnor csa_tree_add_7_25_groupi_g14774__2346(csa_tree_add_7_25_groupi_n_6331 ,csa_tree_add_7_25_groupi_n_6242 ,in3[14]);
  xnor csa_tree_add_7_25_groupi_g14775__1666(csa_tree_add_7_25_groupi_n_6330 ,csa_tree_add_7_25_groupi_n_6240 ,in3[20]);
  xnor csa_tree_add_7_25_groupi_g14776__7410(csa_tree_add_7_25_groupi_n_6328 ,csa_tree_add_7_25_groupi_n_6245 ,in3[17]);
  xnor csa_tree_add_7_25_groupi_g14777__6417(csa_tree_add_7_25_groupi_n_6326 ,csa_tree_add_7_25_groupi_n_6236 ,csa_tree_add_7_25_groupi_n_6109);
  xnor csa_tree_add_7_25_groupi_g14778__5477(csa_tree_add_7_25_groupi_n_6324 ,csa_tree_add_7_25_groupi_n_6234 ,csa_tree_add_7_25_groupi_n_6112);
  xnor csa_tree_add_7_25_groupi_g14779__2398(csa_tree_add_7_25_groupi_n_6322 ,csa_tree_add_7_25_groupi_n_6239 ,in3[23]);
  xnor csa_tree_add_7_25_groupi_g14780__5107(csa_tree_add_7_25_groupi_n_6320 ,csa_tree_add_7_25_groupi_n_6232 ,csa_tree_add_7_25_groupi_n_6121);
  xnor csa_tree_add_7_25_groupi_g14781__6260(csa_tree_add_7_25_groupi_n_6319 ,csa_tree_add_7_25_groupi_n_6230 ,csa_tree_add_7_25_groupi_n_6119);
  xnor csa_tree_add_7_25_groupi_g14782__4319(csa_tree_add_7_25_groupi_n_6318 ,csa_tree_add_7_25_groupi_n_6235 ,csa_tree_add_7_25_groupi_n_6116);
  xnor csa_tree_add_7_25_groupi_g14783__8428(csa_tree_add_7_25_groupi_n_6317 ,csa_tree_add_7_25_groupi_n_6233 ,csa_tree_add_7_25_groupi_n_6120);
  xnor csa_tree_add_7_25_groupi_g14784__5526(csa_tree_add_7_25_groupi_n_6315 ,csa_tree_add_7_25_groupi_n_6231 ,csa_tree_add_7_25_groupi_n_6117);
  and csa_tree_add_7_25_groupi_g14785__6783(csa_tree_add_7_25_groupi_n_6302 ,csa_tree_add_7_25_groupi_n_6161 ,csa_tree_add_7_25_groupi_n_6221);
  and csa_tree_add_7_25_groupi_g14786__3680(csa_tree_add_7_25_groupi_n_6301 ,csa_tree_add_7_25_groupi_n_6223 ,csa_tree_add_7_25_groupi_n_6181);
  or csa_tree_add_7_25_groupi_g14787__1617(csa_tree_add_7_25_groupi_n_6300 ,csa_tree_add_7_25_groupi_n_6223 ,csa_tree_add_7_25_groupi_n_6181);
  or csa_tree_add_7_25_groupi_g14788__2802(csa_tree_add_7_25_groupi_n_6299 ,csa_tree_add_7_25_groupi_n_6163 ,csa_tree_add_7_25_groupi_n_6224);
  and csa_tree_add_7_25_groupi_g14789__1705(csa_tree_add_7_25_groupi_n_6298 ,csa_tree_add_7_25_groupi_n_6163 ,csa_tree_add_7_25_groupi_n_6224);
  and csa_tree_add_7_25_groupi_g14790__5122(csa_tree_add_7_25_groupi_n_6297 ,csa_tree_add_7_25_groupi_n_6164 ,csa_tree_add_7_25_groupi_n_6222);
  or csa_tree_add_7_25_groupi_g14791__8246(csa_tree_add_7_25_groupi_n_6296 ,csa_tree_add_7_25_groupi_n_6164 ,csa_tree_add_7_25_groupi_n_6222);
  and csa_tree_add_7_25_groupi_g14792__7098(csa_tree_add_7_25_groupi_n_6295 ,csa_tree_add_7_25_groupi_n_6232 ,csa_tree_add_7_25_groupi_n_6100);
  and csa_tree_add_7_25_groupi_g14793__6131(csa_tree_add_7_25_groupi_n_6294 ,csa_tree_add_7_25_groupi_n_6231 ,csa_tree_add_7_25_groupi_n_6098);
  or csa_tree_add_7_25_groupi_g14794__1881(csa_tree_add_7_25_groupi_n_6293 ,csa_tree_add_7_25_groupi_n_3373 ,csa_tree_add_7_25_groupi_n_6254);
  or csa_tree_add_7_25_groupi_g14795__5115(csa_tree_add_7_25_groupi_n_6292 ,csa_tree_add_7_25_groupi_n_6161 ,csa_tree_add_7_25_groupi_n_6221);
  and csa_tree_add_7_25_groupi_g14796__7482(csa_tree_add_7_25_groupi_n_6291 ,csa_tree_add_7_25_groupi_n_6230 ,csa_tree_add_7_25_groupi_n_6094);
  and csa_tree_add_7_25_groupi_g14797__4733(csa_tree_add_7_25_groupi_n_6290 ,csa_tree_add_7_25_groupi_n_6229 ,csa_tree_add_7_25_groupi_n_6092);
  and csa_tree_add_7_25_groupi_g14798__6161(csa_tree_add_7_25_groupi_n_6289 ,csa_tree_add_7_25_groupi_n_6162 ,csa_tree_add_7_25_groupi_n_6210);
  or csa_tree_add_7_25_groupi_g14799__9315(csa_tree_add_7_25_groupi_n_6288 ,csa_tree_add_7_25_groupi_n_6162 ,csa_tree_add_7_25_groupi_n_6210);
  and csa_tree_add_7_25_groupi_g14800__9945(csa_tree_add_7_25_groupi_n_6287 ,csa_tree_add_7_25_groupi_n_6235 ,csa_tree_add_7_25_groupi_n_6089);
  or csa_tree_add_7_25_groupi_g14801__2883(csa_tree_add_7_25_groupi_n_6286 ,csa_tree_add_7_25_groupi_n_3376 ,csa_tree_add_7_25_groupi_n_6251);
  and csa_tree_add_7_25_groupi_g14802__2346(csa_tree_add_7_25_groupi_n_6303 ,csa_tree_add_7_25_groupi_n_2429 ,csa_tree_add_7_25_groupi_n_6255);
  or csa_tree_add_7_25_groupi_g14803__1666(csa_tree_add_7_25_groupi_n_6283 ,csa_tree_add_7_25_groupi_n_6185 ,csa_tree_add_7_25_groupi_n_6211);
  or csa_tree_add_7_25_groupi_g14804__7410(csa_tree_add_7_25_groupi_n_6282 ,csa_tree_add_7_25_groupi_n_6180 ,csa_tree_add_7_25_groupi_n_6227);
  or csa_tree_add_7_25_groupi_g14805__6417(csa_tree_add_7_25_groupi_n_6281 ,csa_tree_add_7_25_groupi_n_3748 ,csa_tree_add_7_25_groupi_n_6248);
  or csa_tree_add_7_25_groupi_g14806__5477(csa_tree_add_7_25_groupi_n_6280 ,csa_tree_add_7_25_groupi_n_3751 ,csa_tree_add_7_25_groupi_n_6249);
  or csa_tree_add_7_25_groupi_g14807__2398(csa_tree_add_7_25_groupi_n_6279 ,csa_tree_add_7_25_groupi_n_3750 ,csa_tree_add_7_25_groupi_n_6250);
  or csa_tree_add_7_25_groupi_g14808__5107(csa_tree_add_7_25_groupi_n_6278 ,csa_tree_add_7_25_groupi_n_3753 ,csa_tree_add_7_25_groupi_n_6252);
  or csa_tree_add_7_25_groupi_g14809__6260(csa_tree_add_7_25_groupi_n_6277 ,csa_tree_add_7_25_groupi_n_3752 ,csa_tree_add_7_25_groupi_n_6253);
  and csa_tree_add_7_25_groupi_g14810__4319(csa_tree_add_7_25_groupi_n_6276 ,csa_tree_add_7_25_groupi_n_6236 ,csa_tree_add_7_25_groupi_n_6084);
  nor csa_tree_add_7_25_groupi_g14811__8428(csa_tree_add_7_25_groupi_n_6275 ,csa_tree_add_7_25_groupi_n_6184 ,csa_tree_add_7_25_groupi_n_6212);
  nor csa_tree_add_7_25_groupi_g14812__5526(csa_tree_add_7_25_groupi_n_6274 ,csa_tree_add_7_25_groupi_n_6179 ,csa_tree_add_7_25_groupi_n_6228);
  and csa_tree_add_7_25_groupi_g14813__6783(csa_tree_add_7_25_groupi_n_6273 ,csa_tree_add_7_25_groupi_n_6234 ,csa_tree_add_7_25_groupi_n_6077);
  nor csa_tree_add_7_25_groupi_g14814__3680(csa_tree_add_7_25_groupi_n_6272 ,csa_tree_add_7_25_groupi_n_6182 ,csa_tree_add_7_25_groupi_n_6214);
  or csa_tree_add_7_25_groupi_g14815__1617(csa_tree_add_7_25_groupi_n_6271 ,csa_tree_add_7_25_groupi_n_6183 ,csa_tree_add_7_25_groupi_n_6213);
  and csa_tree_add_7_25_groupi_g14816__2802(csa_tree_add_7_25_groupi_n_6270 ,csa_tree_add_7_25_groupi_n_6233 ,csa_tree_add_7_25_groupi_n_6072);
  or csa_tree_add_7_25_groupi_g14817__1705(csa_tree_add_7_25_groupi_n_6269 ,csa_tree_add_7_25_groupi_n_3310 ,csa_tree_add_7_25_groupi_n_6247);
  or csa_tree_add_7_25_groupi_g14818__5122(csa_tree_add_7_25_groupi_n_6268 ,csa_tree_add_7_25_groupi_n_6165 ,csa_tree_add_7_25_groupi_n_6225);
  and csa_tree_add_7_25_groupi_g14819__8246(csa_tree_add_7_25_groupi_n_6267 ,csa_tree_add_7_25_groupi_n_6165 ,csa_tree_add_7_25_groupi_n_6225);
  or csa_tree_add_7_25_groupi_g14820__7098(csa_tree_add_7_25_groupi_n_6285 ,csa_tree_add_7_25_groupi_n_6246 ,csa_tree_add_7_25_groupi_n_6176);
  xnor csa_tree_add_7_25_groupi_g14821__6131(csa_tree_add_7_25_groupi_n_6284 ,csa_tree_add_7_25_groupi_n_6201 ,csa_tree_add_7_25_groupi_n_2565);
  not csa_tree_add_7_25_groupi_g14822(csa_tree_add_7_25_groupi_n_6264 ,csa_tree_add_7_25_groupi_n_6265);
  not csa_tree_add_7_25_groupi_g14823(csa_tree_add_7_25_groupi_n_6262 ,csa_tree_add_7_25_groupi_n_6263);
  not csa_tree_add_7_25_groupi_g14824(csa_tree_add_7_25_groupi_n_6256 ,csa_tree_add_7_25_groupi_n_6257);
  or csa_tree_add_7_25_groupi_g14825__1881(csa_tree_add_7_25_groupi_n_6255 ,csa_tree_add_7_25_groupi_n_2473 ,csa_tree_add_7_25_groupi_n_6201);
  nor csa_tree_add_7_25_groupi_g14826__5115(csa_tree_add_7_25_groupi_n_6254 ,csa_tree_add_7_25_groupi_n_2126 ,csa_tree_add_7_25_groupi_n_1271);
  nor csa_tree_add_7_25_groupi_g14827__7482(csa_tree_add_7_25_groupi_n_6253 ,csa_tree_add_7_25_groupi_n_2105 ,csa_tree_add_7_25_groupi_n_1283);
  nor csa_tree_add_7_25_groupi_g14828__4733(csa_tree_add_7_25_groupi_n_6252 ,csa_tree_add_7_25_groupi_n_2159 ,csa_tree_add_7_25_groupi_n_1282);
  nor csa_tree_add_7_25_groupi_g14829__6161(csa_tree_add_7_25_groupi_n_6251 ,csa_tree_add_7_25_groupi_n_2138 ,csa_tree_add_7_25_groupi_n_1282);
  nor csa_tree_add_7_25_groupi_g14830__9315(csa_tree_add_7_25_groupi_n_6250 ,csa_tree_add_7_25_groupi_n_2060 ,csa_tree_add_7_25_groupi_n_1270);
  nor csa_tree_add_7_25_groupi_g14831__9945(csa_tree_add_7_25_groupi_n_6249 ,csa_tree_add_7_25_groupi_n_2043 ,csa_tree_add_7_25_groupi_n_1270);
  nor csa_tree_add_7_25_groupi_g14832__2883(csa_tree_add_7_25_groupi_n_6248 ,csa_tree_add_7_25_groupi_n_2031 ,csa_tree_add_7_25_groupi_n_1283);
  nor csa_tree_add_7_25_groupi_g14833__2346(csa_tree_add_7_25_groupi_n_6247 ,csa_tree_add_7_25_groupi_n_2186 ,csa_tree_add_7_25_groupi_n_1271);
  and csa_tree_add_7_25_groupi_g14834__1666(csa_tree_add_7_25_groupi_n_6246 ,csa_tree_add_7_25_groupi_n_6202 ,csa_tree_add_7_25_groupi_n_6169);
  nor csa_tree_add_7_25_groupi_g14835__7410(csa_tree_add_7_25_groupi_n_6245 ,csa_tree_add_7_25_groupi_n_3907 ,csa_tree_add_7_25_groupi_n_6173);
  nor csa_tree_add_7_25_groupi_g14836__6417(csa_tree_add_7_25_groupi_n_6244 ,csa_tree_add_7_25_groupi_n_3489 ,csa_tree_add_7_25_groupi_n_6167);
  nor csa_tree_add_7_25_groupi_g14837__5477(csa_tree_add_7_25_groupi_n_6243 ,csa_tree_add_7_25_groupi_n_3817 ,csa_tree_add_7_25_groupi_n_6171);
  nor csa_tree_add_7_25_groupi_g14838__2398(csa_tree_add_7_25_groupi_n_6242 ,csa_tree_add_7_25_groupi_n_3913 ,csa_tree_add_7_25_groupi_n_6172);
  or csa_tree_add_7_25_groupi_g14839__5107(csa_tree_add_7_25_groupi_n_6241 ,csa_tree_add_7_25_groupi_n_5961 ,csa_tree_add_7_25_groupi_n_6177);
  nor csa_tree_add_7_25_groupi_g14840__6260(csa_tree_add_7_25_groupi_n_6240 ,csa_tree_add_7_25_groupi_n_3842 ,csa_tree_add_7_25_groupi_n_6174);
  nor csa_tree_add_7_25_groupi_g14841__4319(csa_tree_add_7_25_groupi_n_6239 ,csa_tree_add_7_25_groupi_n_3820 ,csa_tree_add_7_25_groupi_n_6175);
  nor csa_tree_add_7_25_groupi_g14842__8428(csa_tree_add_7_25_groupi_n_6238 ,csa_tree_add_7_25_groupi_n_4099 ,csa_tree_add_7_25_groupi_n_6199);
  nor csa_tree_add_7_25_groupi_g14843__5526(csa_tree_add_7_25_groupi_n_6237 ,csa_tree_add_7_25_groupi_n_4086 ,csa_tree_add_7_25_groupi_n_6198);
  or csa_tree_add_7_25_groupi_g14844__6783(csa_tree_add_7_25_groupi_n_6266 ,csa_tree_add_7_25_groupi_n_5983 ,csa_tree_add_7_25_groupi_n_6193);
  or csa_tree_add_7_25_groupi_g14845__3680(csa_tree_add_7_25_groupi_n_6265 ,csa_tree_add_7_25_groupi_n_5970 ,csa_tree_add_7_25_groupi_n_6168);
  or csa_tree_add_7_25_groupi_g14846__1617(csa_tree_add_7_25_groupi_n_6263 ,csa_tree_add_7_25_groupi_n_5977 ,csa_tree_add_7_25_groupi_n_6170);
  or csa_tree_add_7_25_groupi_g14847__2802(csa_tree_add_7_25_groupi_n_6261 ,csa_tree_add_7_25_groupi_n_5982 ,csa_tree_add_7_25_groupi_n_6188);
  or csa_tree_add_7_25_groupi_g14848__1705(csa_tree_add_7_25_groupi_n_6260 ,csa_tree_add_7_25_groupi_n_5963 ,csa_tree_add_7_25_groupi_n_6166);
  or csa_tree_add_7_25_groupi_g14849__5122(csa_tree_add_7_25_groupi_n_6259 ,csa_tree_add_7_25_groupi_n_5989 ,csa_tree_add_7_25_groupi_n_6196);
  or csa_tree_add_7_25_groupi_g14850__8246(csa_tree_add_7_25_groupi_n_6258 ,csa_tree_add_7_25_groupi_n_5994 ,csa_tree_add_7_25_groupi_n_6197);
  or csa_tree_add_7_25_groupi_g14851__7098(csa_tree_add_7_25_groupi_n_6257 ,csa_tree_add_7_25_groupi_n_5995 ,csa_tree_add_7_25_groupi_n_6200);
  not csa_tree_add_7_25_groupi_g14852(csa_tree_add_7_25_groupi_n_6227 ,csa_tree_add_7_25_groupi_n_6228);
  not csa_tree_add_7_25_groupi_g14853(csa_tree_add_7_25_groupi_n_6219 ,csa_tree_add_7_25_groupi_n_6220);
  not csa_tree_add_7_25_groupi_g14854(csa_tree_add_7_25_groupi_n_6217 ,csa_tree_add_7_25_groupi_n_6218);
  not csa_tree_add_7_25_groupi_g14855(csa_tree_add_7_25_groupi_n_6215 ,csa_tree_add_7_25_groupi_n_6216);
  not csa_tree_add_7_25_groupi_g14856(csa_tree_add_7_25_groupi_n_6213 ,csa_tree_add_7_25_groupi_n_6214);
  not csa_tree_add_7_25_groupi_g14857(csa_tree_add_7_25_groupi_n_6211 ,csa_tree_add_7_25_groupi_n_6212);
  xnor csa_tree_add_7_25_groupi_g14858__6131(out2[13] ,csa_tree_add_7_25_groupi_n_6107 ,csa_tree_add_7_25_groupi_n_6122);
  xnor csa_tree_add_7_25_groupi_g14859__1881(csa_tree_add_7_25_groupi_n_6208 ,csa_tree_add_7_25_groupi_n_6057 ,csa_tree_add_7_25_groupi_n_6126);
  xnor csa_tree_add_7_25_groupi_g14860__5115(csa_tree_add_7_25_groupi_n_6207 ,csa_tree_add_7_25_groupi_n_6128 ,csa_tree_add_7_25_groupi_n_6060);
  xnor csa_tree_add_7_25_groupi_g14861__7482(csa_tree_add_7_25_groupi_n_6206 ,csa_tree_add_7_25_groupi_n_6058 ,csa_tree_add_7_25_groupi_n_6127);
  xnor csa_tree_add_7_25_groupi_g14862__4733(csa_tree_add_7_25_groupi_n_6205 ,csa_tree_add_7_25_groupi_n_6059 ,csa_tree_add_7_25_groupi_n_6125);
  xnor csa_tree_add_7_25_groupi_g14863__6161(csa_tree_add_7_25_groupi_n_6204 ,csa_tree_add_7_25_groupi_n_6061 ,csa_tree_add_7_25_groupi_n_6124);
  xnor csa_tree_add_7_25_groupi_g14864__9315(csa_tree_add_7_25_groupi_n_6203 ,csa_tree_add_7_25_groupi_n_6144 ,in3[26]);
  xnor csa_tree_add_7_25_groupi_g14865__9945(csa_tree_add_7_25_groupi_n_6236 ,csa_tree_add_7_25_groupi_n_6143 ,in3[23]);
  xnor csa_tree_add_7_25_groupi_g14866__2883(csa_tree_add_7_25_groupi_n_6235 ,csa_tree_add_7_25_groupi_n_6141 ,in3[8]);
  xnor csa_tree_add_7_25_groupi_g14867__2346(csa_tree_add_7_25_groupi_n_6234 ,csa_tree_add_7_25_groupi_n_6139 ,in3[20]);
  xnor csa_tree_add_7_25_groupi_g14868__1666(csa_tree_add_7_25_groupi_n_6233 ,csa_tree_add_7_25_groupi_n_6145 ,in3[17]);
  xnor csa_tree_add_7_25_groupi_g14869__7410(csa_tree_add_7_25_groupi_n_6232 ,csa_tree_add_7_25_groupi_n_6142 ,in3[2]);
  xnor csa_tree_add_7_25_groupi_g14870__6417(csa_tree_add_7_25_groupi_n_6231 ,csa_tree_add_7_25_groupi_n_6138 ,in3[14]);
  xnor csa_tree_add_7_25_groupi_g14871__5477(csa_tree_add_7_25_groupi_n_6230 ,csa_tree_add_7_25_groupi_n_6146 ,in3[5]);
  xnor csa_tree_add_7_25_groupi_g14872__2398(csa_tree_add_7_25_groupi_n_6229 ,csa_tree_add_7_25_groupi_n_6140 ,in3[11]);
  xnor csa_tree_add_7_25_groupi_g14873__5107(csa_tree_add_7_25_groupi_n_6228 ,csa_tree_add_7_25_groupi_n_6135 ,csa_tree_add_7_25_groupi_n_6010);
  xnor csa_tree_add_7_25_groupi_g14874__6260(csa_tree_add_7_25_groupi_n_6226 ,csa_tree_add_7_25_groupi_n_6062 ,csa_tree_add_7_25_groupi_n_6114);
  xnor csa_tree_add_7_25_groupi_g14875__4319(csa_tree_add_7_25_groupi_n_6225 ,csa_tree_add_7_25_groupi_n_6131 ,csa_tree_add_7_25_groupi_n_6001);
  xnor csa_tree_add_7_25_groupi_g14876__8428(csa_tree_add_7_25_groupi_n_6224 ,csa_tree_add_7_25_groupi_n_6133 ,csa_tree_add_7_25_groupi_n_6006);
  xnor csa_tree_add_7_25_groupi_g14877__5526(csa_tree_add_7_25_groupi_n_6223 ,csa_tree_add_7_25_groupi_n_6134 ,csa_tree_add_7_25_groupi_n_6011);
  xnor csa_tree_add_7_25_groupi_g14878__6783(csa_tree_add_7_25_groupi_n_6222 ,csa_tree_add_7_25_groupi_n_6130 ,csa_tree_add_7_25_groupi_n_6005);
  xnor csa_tree_add_7_25_groupi_g14879__3680(csa_tree_add_7_25_groupi_n_6221 ,csa_tree_add_7_25_groupi_n_6129 ,csa_tree_add_7_25_groupi_n_6004);
  xnor csa_tree_add_7_25_groupi_g14880__1617(csa_tree_add_7_25_groupi_n_6220 ,csa_tree_add_7_25_groupi_n_6065 ,csa_tree_add_7_25_groupi_n_6111);
  xnor csa_tree_add_7_25_groupi_g14881__2802(csa_tree_add_7_25_groupi_n_6218 ,csa_tree_add_7_25_groupi_n_6063 ,csa_tree_add_7_25_groupi_n_6115);
  xnor csa_tree_add_7_25_groupi_g14882__1705(csa_tree_add_7_25_groupi_n_6216 ,csa_tree_add_7_25_groupi_n_6064 ,csa_tree_add_7_25_groupi_n_6113);
  xnor csa_tree_add_7_25_groupi_g14883__5122(csa_tree_add_7_25_groupi_n_6214 ,csa_tree_add_7_25_groupi_n_6136 ,csa_tree_add_7_25_groupi_n_6008);
  xnor csa_tree_add_7_25_groupi_g14884__8246(csa_tree_add_7_25_groupi_n_6212 ,csa_tree_add_7_25_groupi_n_6137 ,csa_tree_add_7_25_groupi_n_6007);
  xnor csa_tree_add_7_25_groupi_g14885__7098(csa_tree_add_7_25_groupi_n_6210 ,csa_tree_add_7_25_groupi_n_6132 ,csa_tree_add_7_25_groupi_n_6003);
  and csa_tree_add_7_25_groupi_g14886__6131(csa_tree_add_7_25_groupi_n_6200 ,csa_tree_add_7_25_groupi_n_6134 ,csa_tree_add_7_25_groupi_n_5999);
  or csa_tree_add_7_25_groupi_g14887__1881(csa_tree_add_7_25_groupi_n_6199 ,csa_tree_add_7_25_groupi_n_3344 ,csa_tree_add_7_25_groupi_n_6160);
  or csa_tree_add_7_25_groupi_g14888__5115(csa_tree_add_7_25_groupi_n_6198 ,csa_tree_add_7_25_groupi_n_3346 ,csa_tree_add_7_25_groupi_n_6156);
  and csa_tree_add_7_25_groupi_g14889__7482(csa_tree_add_7_25_groupi_n_6197 ,csa_tree_add_7_25_groupi_n_6133 ,csa_tree_add_7_25_groupi_n_5993);
  and csa_tree_add_7_25_groupi_g14890__4733(csa_tree_add_7_25_groupi_n_6196 ,csa_tree_add_7_25_groupi_n_6130 ,csa_tree_add_7_25_groupi_n_5988);
  and csa_tree_add_7_25_groupi_g14891__6161(csa_tree_add_7_25_groupi_n_6195 ,csa_tree_add_7_25_groupi_n_6061 ,csa_tree_add_7_25_groupi_n_6124);
  or csa_tree_add_7_25_groupi_g14892__9315(csa_tree_add_7_25_groupi_n_6194 ,csa_tree_add_7_25_groupi_n_6061 ,csa_tree_add_7_25_groupi_n_6124);
  and csa_tree_add_7_25_groupi_g14893__9945(csa_tree_add_7_25_groupi_n_6193 ,csa_tree_add_7_25_groupi_n_6129 ,csa_tree_add_7_25_groupi_n_5985);
  and csa_tree_add_7_25_groupi_g14894__2883(csa_tree_add_7_25_groupi_n_6192 ,csa_tree_add_7_25_groupi_n_6059 ,csa_tree_add_7_25_groupi_n_6125);
  or csa_tree_add_7_25_groupi_g14895__2346(csa_tree_add_7_25_groupi_n_6191 ,csa_tree_add_7_25_groupi_n_6059 ,csa_tree_add_7_25_groupi_n_6125);
  or csa_tree_add_7_25_groupi_g14896__1666(csa_tree_add_7_25_groupi_n_6190 ,csa_tree_add_7_25_groupi_n_6128 ,csa_tree_add_7_25_groupi_n_6060);
  and csa_tree_add_7_25_groupi_g14897__7410(csa_tree_add_7_25_groupi_n_6189 ,csa_tree_add_7_25_groupi_n_6128 ,csa_tree_add_7_25_groupi_n_6060);
  and csa_tree_add_7_25_groupi_g14898__6417(csa_tree_add_7_25_groupi_n_6188 ,csa_tree_add_7_25_groupi_n_6132 ,csa_tree_add_7_25_groupi_n_5981);
  and csa_tree_add_7_25_groupi_g14899__5477(csa_tree_add_7_25_groupi_n_6187 ,csa_tree_add_7_25_groupi_n_6058 ,csa_tree_add_7_25_groupi_n_6127);
  or csa_tree_add_7_25_groupi_g14900__2398(csa_tree_add_7_25_groupi_n_6186 ,csa_tree_add_7_25_groupi_n_6058 ,csa_tree_add_7_25_groupi_n_6127);
  or csa_tree_add_7_25_groupi_g14901__5107(csa_tree_add_7_25_groupi_n_6202 ,csa_tree_add_7_25_groupi_n_6150 ,csa_tree_add_7_25_groupi_n_6103);
  and csa_tree_add_7_25_groupi_g14902__6260(csa_tree_add_7_25_groupi_n_6201 ,csa_tree_add_7_25_groupi_n_2415 ,csa_tree_add_7_25_groupi_n_6157);
  not csa_tree_add_7_25_groupi_g14903(csa_tree_add_7_25_groupi_n_6184 ,csa_tree_add_7_25_groupi_n_6185);
  not csa_tree_add_7_25_groupi_g14904(csa_tree_add_7_25_groupi_n_6182 ,csa_tree_add_7_25_groupi_n_6183);
  not csa_tree_add_7_25_groupi_g14905(csa_tree_add_7_25_groupi_n_6179 ,csa_tree_add_7_25_groupi_n_6180);
  and csa_tree_add_7_25_groupi_g14906__4319(csa_tree_add_7_25_groupi_n_6177 ,csa_tree_add_7_25_groupi_n_6135 ,csa_tree_add_7_25_groupi_n_5978);
  and csa_tree_add_7_25_groupi_g14907__8428(csa_tree_add_7_25_groupi_n_6176 ,csa_tree_add_7_25_groupi_n_6057 ,csa_tree_add_7_25_groupi_n_6126);
  or csa_tree_add_7_25_groupi_g14908__5526(csa_tree_add_7_25_groupi_n_6175 ,csa_tree_add_7_25_groupi_n_3745 ,csa_tree_add_7_25_groupi_n_6153);
  or csa_tree_add_7_25_groupi_g14909__6783(csa_tree_add_7_25_groupi_n_6174 ,csa_tree_add_7_25_groupi_n_3740 ,csa_tree_add_7_25_groupi_n_6154);
  or csa_tree_add_7_25_groupi_g14910__3680(csa_tree_add_7_25_groupi_n_6173 ,csa_tree_add_7_25_groupi_n_3747 ,csa_tree_add_7_25_groupi_n_6155);
  or csa_tree_add_7_25_groupi_g14911__1617(csa_tree_add_7_25_groupi_n_6172 ,csa_tree_add_7_25_groupi_n_3637 ,csa_tree_add_7_25_groupi_n_6158);
  or csa_tree_add_7_25_groupi_g14912__2802(csa_tree_add_7_25_groupi_n_6171 ,csa_tree_add_7_25_groupi_n_3847 ,csa_tree_add_7_25_groupi_n_6159);
  and csa_tree_add_7_25_groupi_g14913__1705(csa_tree_add_7_25_groupi_n_6170 ,csa_tree_add_7_25_groupi_n_6137 ,csa_tree_add_7_25_groupi_n_5976);
  or csa_tree_add_7_25_groupi_g14914__5122(csa_tree_add_7_25_groupi_n_6169 ,csa_tree_add_7_25_groupi_n_6057 ,csa_tree_add_7_25_groupi_n_6126);
  and csa_tree_add_7_25_groupi_g14915__8246(csa_tree_add_7_25_groupi_n_6168 ,csa_tree_add_7_25_groupi_n_6136 ,csa_tree_add_7_25_groupi_n_5969);
  or csa_tree_add_7_25_groupi_g14916__7098(csa_tree_add_7_25_groupi_n_6167 ,csa_tree_add_7_25_groupi_n_3281 ,csa_tree_add_7_25_groupi_n_6152);
  and csa_tree_add_7_25_groupi_g14917__6131(csa_tree_add_7_25_groupi_n_6166 ,csa_tree_add_7_25_groupi_n_6131 ,csa_tree_add_7_25_groupi_n_5962);
  or csa_tree_add_7_25_groupi_g14918__1881(csa_tree_add_7_25_groupi_n_6185 ,csa_tree_add_7_25_groupi_n_6076 ,csa_tree_add_7_25_groupi_n_6148);
  or csa_tree_add_7_25_groupi_g14919__5115(csa_tree_add_7_25_groupi_n_6183 ,csa_tree_add_7_25_groupi_n_6149 ,csa_tree_add_7_25_groupi_n_6070);
  or csa_tree_add_7_25_groupi_g14920__7482(csa_tree_add_7_25_groupi_n_6181 ,csa_tree_add_7_25_groupi_n_6151 ,csa_tree_add_7_25_groupi_n_6068);
  or csa_tree_add_7_25_groupi_g14921__4733(csa_tree_add_7_25_groupi_n_6180 ,csa_tree_add_7_25_groupi_n_6083 ,csa_tree_add_7_25_groupi_n_6147);
  xnor csa_tree_add_7_25_groupi_g14922__6161(csa_tree_add_7_25_groupi_n_6178 ,csa_tree_add_7_25_groupi_n_6108 ,csa_tree_add_7_25_groupi_n_2566);
  nor csa_tree_add_7_25_groupi_g14923(csa_tree_add_7_25_groupi_n_6160 ,csa_tree_add_7_25_groupi_n_2123 ,csa_tree_add_7_25_groupi_n_1280);
  nor csa_tree_add_7_25_groupi_g14924(csa_tree_add_7_25_groupi_n_6159 ,csa_tree_add_7_25_groupi_n_2102 ,csa_tree_add_7_25_groupi_n_1274);
  nor csa_tree_add_7_25_groupi_g14925(csa_tree_add_7_25_groupi_n_6158 ,csa_tree_add_7_25_groupi_n_2156 ,csa_tree_add_7_25_groupi_n_1273);
  or csa_tree_add_7_25_groupi_g14926(csa_tree_add_7_25_groupi_n_6157 ,csa_tree_add_7_25_groupi_n_2445 ,csa_tree_add_7_25_groupi_n_6108);
  nor csa_tree_add_7_25_groupi_g14927(csa_tree_add_7_25_groupi_n_6156 ,csa_tree_add_7_25_groupi_n_2141 ,csa_tree_add_7_25_groupi_n_1273);
  nor csa_tree_add_7_25_groupi_g14928(csa_tree_add_7_25_groupi_n_6155 ,csa_tree_add_7_25_groupi_n_2064 ,csa_tree_add_7_25_groupi_n_1279);
  nor csa_tree_add_7_25_groupi_g14929(csa_tree_add_7_25_groupi_n_6154 ,csa_tree_add_7_25_groupi_n_2048 ,csa_tree_add_7_25_groupi_n_1279);
  nor csa_tree_add_7_25_groupi_g14930(csa_tree_add_7_25_groupi_n_6153 ,csa_tree_add_7_25_groupi_n_2019 ,csa_tree_add_7_25_groupi_n_1274);
  nor csa_tree_add_7_25_groupi_g14931(csa_tree_add_7_25_groupi_n_6152 ,csa_tree_add_7_25_groupi_n_2183 ,csa_tree_add_7_25_groupi_n_1280);
  and csa_tree_add_7_25_groupi_g14932(csa_tree_add_7_25_groupi_n_6151 ,csa_tree_add_7_25_groupi_n_6062 ,csa_tree_add_7_25_groupi_n_6069);
  and csa_tree_add_7_25_groupi_g14933(csa_tree_add_7_25_groupi_n_6150 ,csa_tree_add_7_25_groupi_n_6107 ,csa_tree_add_7_25_groupi_n_6104);
  and csa_tree_add_7_25_groupi_g14934(csa_tree_add_7_25_groupi_n_6149 ,csa_tree_add_7_25_groupi_n_6071 ,csa_tree_add_7_25_groupi_n_6063);
  and csa_tree_add_7_25_groupi_g14935(csa_tree_add_7_25_groupi_n_6148 ,csa_tree_add_7_25_groupi_n_6086 ,csa_tree_add_7_25_groupi_n_6064);
  and csa_tree_add_7_25_groupi_g14936(csa_tree_add_7_25_groupi_n_6147 ,csa_tree_add_7_25_groupi_n_6065 ,csa_tree_add_7_25_groupi_n_6082);
  nor csa_tree_add_7_25_groupi_g14937(csa_tree_add_7_25_groupi_n_6146 ,csa_tree_add_7_25_groupi_n_4050 ,csa_tree_add_7_25_groupi_n_6105);
  nor csa_tree_add_7_25_groupi_g14938(csa_tree_add_7_25_groupi_n_6145 ,csa_tree_add_7_25_groupi_n_4040 ,csa_tree_add_7_25_groupi_n_6088);
  nor csa_tree_add_7_25_groupi_g14939(csa_tree_add_7_25_groupi_n_6144 ,csa_tree_add_7_25_groupi_n_3926 ,csa_tree_add_7_25_groupi_n_6081);
  nor csa_tree_add_7_25_groupi_g14940(csa_tree_add_7_25_groupi_n_6143 ,csa_tree_add_7_25_groupi_n_3939 ,csa_tree_add_7_25_groupi_n_6080);
  nor csa_tree_add_7_25_groupi_g14941(csa_tree_add_7_25_groupi_n_6142 ,csa_tree_add_7_25_groupi_n_3497 ,csa_tree_add_7_25_groupi_n_6066);
  nor csa_tree_add_7_25_groupi_g14942(csa_tree_add_7_25_groupi_n_6141 ,csa_tree_add_7_25_groupi_n_4039 ,csa_tree_add_7_25_groupi_n_6075);
  nor csa_tree_add_7_25_groupi_g14943(csa_tree_add_7_25_groupi_n_6140 ,csa_tree_add_7_25_groupi_n_4015 ,csa_tree_add_7_25_groupi_n_6106);
  nor csa_tree_add_7_25_groupi_g14944(csa_tree_add_7_25_groupi_n_6139 ,csa_tree_add_7_25_groupi_n_3875 ,csa_tree_add_7_25_groupi_n_6079);
  nor csa_tree_add_7_25_groupi_g14945(csa_tree_add_7_25_groupi_n_6138 ,csa_tree_add_7_25_groupi_n_3823 ,csa_tree_add_7_25_groupi_n_6074);
  or csa_tree_add_7_25_groupi_g14946(csa_tree_add_7_25_groupi_n_6165 ,csa_tree_add_7_25_groupi_n_5875 ,csa_tree_add_7_25_groupi_n_6097);
  or csa_tree_add_7_25_groupi_g14947(csa_tree_add_7_25_groupi_n_6164 ,csa_tree_add_7_25_groupi_n_5878 ,csa_tree_add_7_25_groupi_n_6102);
  or csa_tree_add_7_25_groupi_g14948(csa_tree_add_7_25_groupi_n_6163 ,csa_tree_add_7_25_groupi_n_5851 ,csa_tree_add_7_25_groupi_n_6067);
  or csa_tree_add_7_25_groupi_g14949(csa_tree_add_7_25_groupi_n_6162 ,csa_tree_add_7_25_groupi_n_5870 ,csa_tree_add_7_25_groupi_n_6091);
  or csa_tree_add_7_25_groupi_g14950(csa_tree_add_7_25_groupi_n_6161 ,csa_tree_add_7_25_groupi_n_5872 ,csa_tree_add_7_25_groupi_n_6096);
  xnor csa_tree_add_7_25_groupi_g14951(out2[12] ,csa_tree_add_7_25_groupi_n_5980 ,csa_tree_add_7_25_groupi_n_6009);
  xnor csa_tree_add_7_25_groupi_g14952(csa_tree_add_7_25_groupi_n_6122 ,csa_tree_add_7_25_groupi_n_5948 ,csa_tree_add_7_25_groupi_n_6031);
  xnor csa_tree_add_7_25_groupi_g14953(csa_tree_add_7_25_groupi_n_6121 ,csa_tree_add_7_25_groupi_n_5959 ,csa_tree_add_7_25_groupi_n_6025);
  xnor csa_tree_add_7_25_groupi_g14954(csa_tree_add_7_25_groupi_n_6120 ,csa_tree_add_7_25_groupi_n_5950 ,csa_tree_add_7_25_groupi_n_6020);
  xnor csa_tree_add_7_25_groupi_g14955(csa_tree_add_7_25_groupi_n_6119 ,csa_tree_add_7_25_groupi_n_5951 ,csa_tree_add_7_25_groupi_n_6028);
  xnor csa_tree_add_7_25_groupi_g14956(csa_tree_add_7_25_groupi_n_6118 ,csa_tree_add_7_25_groupi_n_5953 ,csa_tree_add_7_25_groupi_n_6023);
  xnor csa_tree_add_7_25_groupi_g14957(csa_tree_add_7_25_groupi_n_6117 ,csa_tree_add_7_25_groupi_n_5958 ,csa_tree_add_7_25_groupi_n_6024);
  xnor csa_tree_add_7_25_groupi_g14958(csa_tree_add_7_25_groupi_n_6116 ,csa_tree_add_7_25_groupi_n_5952 ,csa_tree_add_7_25_groupi_n_6022);
  xnor csa_tree_add_7_25_groupi_g14959(csa_tree_add_7_25_groupi_n_6115 ,csa_tree_add_7_25_groupi_n_6018 ,csa_tree_add_7_25_groupi_n_5911);
  xnor csa_tree_add_7_25_groupi_g14960(csa_tree_add_7_25_groupi_n_6114 ,csa_tree_add_7_25_groupi_n_6021 ,csa_tree_add_7_25_groupi_n_5898);
  xnor csa_tree_add_7_25_groupi_g14961(csa_tree_add_7_25_groupi_n_6113 ,csa_tree_add_7_25_groupi_n_6014 ,csa_tree_add_7_25_groupi_n_5909);
  xnor csa_tree_add_7_25_groupi_g14962(csa_tree_add_7_25_groupi_n_6112 ,csa_tree_add_7_25_groupi_n_5957 ,csa_tree_add_7_25_groupi_n_6030);
  xnor csa_tree_add_7_25_groupi_g14963(csa_tree_add_7_25_groupi_n_6111 ,csa_tree_add_7_25_groupi_n_6016 ,csa_tree_add_7_25_groupi_n_5907);
  xnor csa_tree_add_7_25_groupi_g14964(csa_tree_add_7_25_groupi_n_6110 ,csa_tree_add_7_25_groupi_n_5933 ,csa_tree_add_7_25_groupi_n_6002);
  xnor csa_tree_add_7_25_groupi_g14965(csa_tree_add_7_25_groupi_n_6109 ,csa_tree_add_7_25_groupi_n_5955 ,csa_tree_add_7_25_groupi_n_6027);
  xnor csa_tree_add_7_25_groupi_g14966(csa_tree_add_7_25_groupi_n_6137 ,csa_tree_add_7_25_groupi_n_6041 ,in3[23]);
  xnor csa_tree_add_7_25_groupi_g14967(csa_tree_add_7_25_groupi_n_6136 ,csa_tree_add_7_25_groupi_n_6040 ,in3[20]);
  xnor csa_tree_add_7_25_groupi_g14968(csa_tree_add_7_25_groupi_n_6135 ,csa_tree_add_7_25_groupi_n_6039 ,in3[26]);
  xnor csa_tree_add_7_25_groupi_g14969(csa_tree_add_7_25_groupi_n_6134 ,csa_tree_add_7_25_groupi_n_6045 ,in3[17]);
  xnor csa_tree_add_7_25_groupi_g14970(csa_tree_add_7_25_groupi_n_6133 ,csa_tree_add_7_25_groupi_n_6037 ,in3[2]);
  xnor csa_tree_add_7_25_groupi_g14971(csa_tree_add_7_25_groupi_n_6132 ,csa_tree_add_7_25_groupi_n_6038 ,in3[11]);
  xnor csa_tree_add_7_25_groupi_g14972(csa_tree_add_7_25_groupi_n_6131 ,csa_tree_add_7_25_groupi_n_6042 ,in3[14]);
  xnor csa_tree_add_7_25_groupi_g14973(csa_tree_add_7_25_groupi_n_6130 ,csa_tree_add_7_25_groupi_n_6043 ,in3[5]);
  xnor csa_tree_add_7_25_groupi_g14974(csa_tree_add_7_25_groupi_n_6129 ,csa_tree_add_7_25_groupi_n_6044 ,in3[8]);
  xnor csa_tree_add_7_25_groupi_g14975(csa_tree_add_7_25_groupi_n_6128 ,csa_tree_add_7_25_groupi_n_6033 ,csa_tree_add_7_25_groupi_n_5893);
  xnor csa_tree_add_7_25_groupi_g14976(csa_tree_add_7_25_groupi_n_6127 ,csa_tree_add_7_25_groupi_n_6034 ,csa_tree_add_7_25_groupi_n_5894);
  xnor csa_tree_add_7_25_groupi_g14977(csa_tree_add_7_25_groupi_n_6126 ,csa_tree_add_7_25_groupi_n_6032 ,csa_tree_add_7_25_groupi_n_5891);
  xnor csa_tree_add_7_25_groupi_g14978(csa_tree_add_7_25_groupi_n_6125 ,csa_tree_add_7_25_groupi_n_6036 ,csa_tree_add_7_25_groupi_n_5895);
  xnor csa_tree_add_7_25_groupi_g14979(csa_tree_add_7_25_groupi_n_6124 ,csa_tree_add_7_25_groupi_n_6035 ,csa_tree_add_7_25_groupi_n_5896);
  or csa_tree_add_7_25_groupi_g14980(csa_tree_add_7_25_groupi_n_6106 ,csa_tree_add_7_25_groupi_n_3332 ,csa_tree_add_7_25_groupi_n_6053);
  or csa_tree_add_7_25_groupi_g14981(csa_tree_add_7_25_groupi_n_6105 ,csa_tree_add_7_25_groupi_n_3336 ,csa_tree_add_7_25_groupi_n_6056);
  or csa_tree_add_7_25_groupi_g14982(csa_tree_add_7_25_groupi_n_6104 ,csa_tree_add_7_25_groupi_n_5948 ,csa_tree_add_7_25_groupi_n_6031);
  and csa_tree_add_7_25_groupi_g14983(csa_tree_add_7_25_groupi_n_6103 ,csa_tree_add_7_25_groupi_n_5948 ,csa_tree_add_7_25_groupi_n_6031);
  and csa_tree_add_7_25_groupi_g14984(csa_tree_add_7_25_groupi_n_6102 ,csa_tree_add_7_25_groupi_n_6035 ,csa_tree_add_7_25_groupi_n_5877);
  and csa_tree_add_7_25_groupi_g14985(csa_tree_add_7_25_groupi_n_6101 ,csa_tree_add_7_25_groupi_n_5959 ,csa_tree_add_7_25_groupi_n_6025);
  or csa_tree_add_7_25_groupi_g14986(csa_tree_add_7_25_groupi_n_6100 ,csa_tree_add_7_25_groupi_n_5959 ,csa_tree_add_7_25_groupi_n_6025);
  and csa_tree_add_7_25_groupi_g14987(csa_tree_add_7_25_groupi_n_6099 ,csa_tree_add_7_25_groupi_n_5958 ,csa_tree_add_7_25_groupi_n_6024);
  or csa_tree_add_7_25_groupi_g14988(csa_tree_add_7_25_groupi_n_6098 ,csa_tree_add_7_25_groupi_n_5958 ,csa_tree_add_7_25_groupi_n_6024);
  and csa_tree_add_7_25_groupi_g14989(csa_tree_add_7_25_groupi_n_6097 ,csa_tree_add_7_25_groupi_n_6033 ,csa_tree_add_7_25_groupi_n_5874);
  and csa_tree_add_7_25_groupi_g14990(csa_tree_add_7_25_groupi_n_6096 ,csa_tree_add_7_25_groupi_n_6036 ,csa_tree_add_7_25_groupi_n_5871);
  and csa_tree_add_7_25_groupi_g14991(csa_tree_add_7_25_groupi_n_6095 ,csa_tree_add_7_25_groupi_n_5951 ,csa_tree_add_7_25_groupi_n_6028);
  or csa_tree_add_7_25_groupi_g14992(csa_tree_add_7_25_groupi_n_6094 ,csa_tree_add_7_25_groupi_n_5951 ,csa_tree_add_7_25_groupi_n_6028);
  and csa_tree_add_7_25_groupi_g14993(csa_tree_add_7_25_groupi_n_6093 ,csa_tree_add_7_25_groupi_n_5953 ,csa_tree_add_7_25_groupi_n_6023);
  or csa_tree_add_7_25_groupi_g14994(csa_tree_add_7_25_groupi_n_6092 ,csa_tree_add_7_25_groupi_n_5953 ,csa_tree_add_7_25_groupi_n_6023);
  and csa_tree_add_7_25_groupi_g14995(csa_tree_add_7_25_groupi_n_6091 ,csa_tree_add_7_25_groupi_n_6034 ,csa_tree_add_7_25_groupi_n_5882);
  and csa_tree_add_7_25_groupi_g14996(csa_tree_add_7_25_groupi_n_6090 ,csa_tree_add_7_25_groupi_n_5952 ,csa_tree_add_7_25_groupi_n_6022);
  or csa_tree_add_7_25_groupi_g14997(csa_tree_add_7_25_groupi_n_6089 ,csa_tree_add_7_25_groupi_n_5952 ,csa_tree_add_7_25_groupi_n_6022);
  or csa_tree_add_7_25_groupi_g14998(csa_tree_add_7_25_groupi_n_6088 ,csa_tree_add_7_25_groupi_n_3337 ,csa_tree_add_7_25_groupi_n_6046);
  and csa_tree_add_7_25_groupi_g14999(csa_tree_add_7_25_groupi_n_6108 ,csa_tree_add_7_25_groupi_n_2426 ,csa_tree_add_7_25_groupi_n_6051);
  or csa_tree_add_7_25_groupi_g15000(csa_tree_add_7_25_groupi_n_6107 ,csa_tree_add_7_25_groupi_n_6055 ,csa_tree_add_7_25_groupi_n_5996);
  or csa_tree_add_7_25_groupi_g15001(csa_tree_add_7_25_groupi_n_6086 ,csa_tree_add_7_25_groupi_n_6014 ,csa_tree_add_7_25_groupi_n_5908);
  nor csa_tree_add_7_25_groupi_g15002(csa_tree_add_7_25_groupi_n_6085 ,csa_tree_add_7_25_groupi_n_5954 ,csa_tree_add_7_25_groupi_n_6027);
  or csa_tree_add_7_25_groupi_g15003(csa_tree_add_7_25_groupi_n_6084 ,csa_tree_add_7_25_groupi_n_5955 ,csa_tree_add_7_25_groupi_n_6026);
  nor csa_tree_add_7_25_groupi_g15004(csa_tree_add_7_25_groupi_n_6083 ,csa_tree_add_7_25_groupi_n_6015 ,csa_tree_add_7_25_groupi_n_5907);
  or csa_tree_add_7_25_groupi_g15005(csa_tree_add_7_25_groupi_n_6082 ,csa_tree_add_7_25_groupi_n_6016 ,csa_tree_add_7_25_groupi_n_5906);
  or csa_tree_add_7_25_groupi_g15006(csa_tree_add_7_25_groupi_n_6081 ,csa_tree_add_7_25_groupi_n_3735 ,csa_tree_add_7_25_groupi_n_6049);
  or csa_tree_add_7_25_groupi_g15007(csa_tree_add_7_25_groupi_n_6080 ,csa_tree_add_7_25_groupi_n_3716 ,csa_tree_add_7_25_groupi_n_6048);
  or csa_tree_add_7_25_groupi_g15008(csa_tree_add_7_25_groupi_n_6079 ,csa_tree_add_7_25_groupi_n_3737 ,csa_tree_add_7_25_groupi_n_6047);
  nor csa_tree_add_7_25_groupi_g15009(csa_tree_add_7_25_groupi_n_6078 ,csa_tree_add_7_25_groupi_n_5956 ,csa_tree_add_7_25_groupi_n_6030);
  or csa_tree_add_7_25_groupi_g15010(csa_tree_add_7_25_groupi_n_6077 ,csa_tree_add_7_25_groupi_n_5957 ,csa_tree_add_7_25_groupi_n_6029);
  nor csa_tree_add_7_25_groupi_g15011(csa_tree_add_7_25_groupi_n_6076 ,csa_tree_add_7_25_groupi_n_6013 ,csa_tree_add_7_25_groupi_n_5909);
  or csa_tree_add_7_25_groupi_g15012(csa_tree_add_7_25_groupi_n_6075 ,csa_tree_add_7_25_groupi_n_3333 ,csa_tree_add_7_25_groupi_n_6054);
  or csa_tree_add_7_25_groupi_g15013(csa_tree_add_7_25_groupi_n_6074 ,csa_tree_add_7_25_groupi_n_3725 ,csa_tree_add_7_25_groupi_n_6052);
  nor csa_tree_add_7_25_groupi_g15014(csa_tree_add_7_25_groupi_n_6073 ,csa_tree_add_7_25_groupi_n_5949 ,csa_tree_add_7_25_groupi_n_6020);
  or csa_tree_add_7_25_groupi_g15015(csa_tree_add_7_25_groupi_n_6072 ,csa_tree_add_7_25_groupi_n_5950 ,csa_tree_add_7_25_groupi_n_6019);
  or csa_tree_add_7_25_groupi_g15016(csa_tree_add_7_25_groupi_n_6071 ,csa_tree_add_7_25_groupi_n_6018 ,csa_tree_add_7_25_groupi_n_5910);
  nor csa_tree_add_7_25_groupi_g15017(csa_tree_add_7_25_groupi_n_6070 ,csa_tree_add_7_25_groupi_n_6017 ,csa_tree_add_7_25_groupi_n_5911);
  or csa_tree_add_7_25_groupi_g15018(csa_tree_add_7_25_groupi_n_6069 ,csa_tree_add_7_25_groupi_n_6021 ,csa_tree_add_7_25_groupi_n_5898);
  and csa_tree_add_7_25_groupi_g15019(csa_tree_add_7_25_groupi_n_6068 ,csa_tree_add_7_25_groupi_n_6021 ,csa_tree_add_7_25_groupi_n_5898);
  and csa_tree_add_7_25_groupi_g15020(csa_tree_add_7_25_groupi_n_6067 ,csa_tree_add_7_25_groupi_n_6032 ,csa_tree_add_7_25_groupi_n_5854);
  or csa_tree_add_7_25_groupi_g15021(csa_tree_add_7_25_groupi_n_6066 ,csa_tree_add_7_25_groupi_n_3256 ,csa_tree_add_7_25_groupi_n_6050);
  xnor csa_tree_add_7_25_groupi_g15022(csa_tree_add_7_25_groupi_n_6087 ,csa_tree_add_7_25_groupi_n_6000 ,csa_tree_add_7_25_groupi_n_2567);
  nor csa_tree_add_7_25_groupi_g15023(csa_tree_add_7_25_groupi_n_6056 ,csa_tree_add_7_25_groupi_n_2129 ,csa_tree_add_7_25_groupi_n_1810);
  and csa_tree_add_7_25_groupi_g15024(csa_tree_add_7_25_groupi_n_6055 ,csa_tree_add_7_25_groupi_n_5998 ,csa_tree_add_7_25_groupi_n_5980);
  nor csa_tree_add_7_25_groupi_g15025(csa_tree_add_7_25_groupi_n_6054 ,csa_tree_add_7_25_groupi_n_2114 ,csa_tree_add_7_25_groupi_n_1262);
  nor csa_tree_add_7_25_groupi_g15026(csa_tree_add_7_25_groupi_n_6053 ,csa_tree_add_7_25_groupi_n_2093 ,csa_tree_add_7_25_groupi_n_1261);
  nor csa_tree_add_7_25_groupi_g15027(csa_tree_add_7_25_groupi_n_6052 ,csa_tree_add_7_25_groupi_n_2147 ,csa_tree_add_7_25_groupi_n_1810);
  or csa_tree_add_7_25_groupi_g15028(csa_tree_add_7_25_groupi_n_6051 ,csa_tree_add_7_25_groupi_n_2492 ,csa_tree_add_7_25_groupi_n_6000);
  nor csa_tree_add_7_25_groupi_g15029(csa_tree_add_7_25_groupi_n_6050 ,csa_tree_add_7_25_groupi_n_2171 ,csa_tree_add_7_25_groupi_n_1262);
  nor csa_tree_add_7_25_groupi_g15030(csa_tree_add_7_25_groupi_n_6049 ,csa_tree_add_7_25_groupi_n_1937 ,csa_tree_add_7_25_groupi_n_177);
  nor csa_tree_add_7_25_groupi_g15031(csa_tree_add_7_25_groupi_n_6048 ,csa_tree_add_7_25_groupi_n_2022 ,csa_tree_add_7_25_groupi_n_177);
  nor csa_tree_add_7_25_groupi_g15032(csa_tree_add_7_25_groupi_n_6047 ,csa_tree_add_7_25_groupi_n_2042 ,csa_tree_add_7_25_groupi_n_1261);
  nor csa_tree_add_7_25_groupi_g15033(csa_tree_add_7_25_groupi_n_6046 ,csa_tree_add_7_25_groupi_n_2061 ,csa_tree_add_7_25_groupi_n_176);
  nor csa_tree_add_7_25_groupi_g15034(csa_tree_add_7_25_groupi_n_6045 ,csa_tree_add_7_25_groupi_n_3866 ,csa_tree_add_7_25_groupi_n_5966);
  nor csa_tree_add_7_25_groupi_g15035(csa_tree_add_7_25_groupi_n_6044 ,csa_tree_add_7_25_groupi_n_4097 ,csa_tree_add_7_25_groupi_n_5974);
  nor csa_tree_add_7_25_groupi_g15036(csa_tree_add_7_25_groupi_n_6043 ,csa_tree_add_7_25_groupi_n_4063 ,csa_tree_add_7_25_groupi_n_5975);
  nor csa_tree_add_7_25_groupi_g15037(csa_tree_add_7_25_groupi_n_6042 ,csa_tree_add_7_25_groupi_n_3882 ,csa_tree_add_7_25_groupi_n_5965);
  nor csa_tree_add_7_25_groupi_g15038(csa_tree_add_7_25_groupi_n_6041 ,csa_tree_add_7_25_groupi_n_3844 ,csa_tree_add_7_25_groupi_n_5971);
  nor csa_tree_add_7_25_groupi_g15039(csa_tree_add_7_25_groupi_n_6040 ,csa_tree_add_7_25_groupi_n_3868 ,csa_tree_add_7_25_groupi_n_5967);
  nor csa_tree_add_7_25_groupi_g15040(csa_tree_add_7_25_groupi_n_6039 ,csa_tree_add_7_25_groupi_n_3948 ,csa_tree_add_7_25_groupi_n_5972);
  nor csa_tree_add_7_25_groupi_g15041(csa_tree_add_7_25_groupi_n_6038 ,csa_tree_add_7_25_groupi_n_4010 ,csa_tree_add_7_25_groupi_n_5973);
  nor csa_tree_add_7_25_groupi_g15042(csa_tree_add_7_25_groupi_n_6037 ,csa_tree_add_7_25_groupi_n_3496 ,csa_tree_add_7_25_groupi_n_5960);
  or csa_tree_add_7_25_groupi_g15043(csa_tree_add_7_25_groupi_n_6065 ,csa_tree_add_7_25_groupi_n_5744 ,csa_tree_add_7_25_groupi_n_5990);
  or csa_tree_add_7_25_groupi_g15044(csa_tree_add_7_25_groupi_n_6064 ,csa_tree_add_7_25_groupi_n_5761 ,csa_tree_add_7_25_groupi_n_5968);
  or csa_tree_add_7_25_groupi_g15045(csa_tree_add_7_25_groupi_n_6063 ,csa_tree_add_7_25_groupi_n_5752 ,csa_tree_add_7_25_groupi_n_5964);
  or csa_tree_add_7_25_groupi_g15046(csa_tree_add_7_25_groupi_n_6062 ,csa_tree_add_7_25_groupi_n_5778 ,csa_tree_add_7_25_groupi_n_5991);
  or csa_tree_add_7_25_groupi_g15047(csa_tree_add_7_25_groupi_n_6061 ,csa_tree_add_7_25_groupi_n_5774 ,csa_tree_add_7_25_groupi_n_5987);
  or csa_tree_add_7_25_groupi_g15048(csa_tree_add_7_25_groupi_n_6060 ,csa_tree_add_7_25_groupi_n_5771 ,csa_tree_add_7_25_groupi_n_5986);
  or csa_tree_add_7_25_groupi_g15049(csa_tree_add_7_25_groupi_n_6059 ,csa_tree_add_7_25_groupi_n_5768 ,csa_tree_add_7_25_groupi_n_5984);
  or csa_tree_add_7_25_groupi_g15050(csa_tree_add_7_25_groupi_n_6058 ,csa_tree_add_7_25_groupi_n_5766 ,csa_tree_add_7_25_groupi_n_5997);
  or csa_tree_add_7_25_groupi_g15051(csa_tree_add_7_25_groupi_n_6057 ,csa_tree_add_7_25_groupi_n_5779 ,csa_tree_add_7_25_groupi_n_5992);
  not csa_tree_add_7_25_groupi_g15052(csa_tree_add_7_25_groupi_n_6029 ,csa_tree_add_7_25_groupi_n_6030);
  not csa_tree_add_7_25_groupi_g15053(csa_tree_add_7_25_groupi_n_6026 ,csa_tree_add_7_25_groupi_n_6027);
  not csa_tree_add_7_25_groupi_g15054(csa_tree_add_7_25_groupi_n_6019 ,csa_tree_add_7_25_groupi_n_6020);
  not csa_tree_add_7_25_groupi_g15055(csa_tree_add_7_25_groupi_n_6017 ,csa_tree_add_7_25_groupi_n_6018);
  not csa_tree_add_7_25_groupi_g15056(csa_tree_add_7_25_groupi_n_6015 ,csa_tree_add_7_25_groupi_n_6016);
  not csa_tree_add_7_25_groupi_g15057(csa_tree_add_7_25_groupi_n_6013 ,csa_tree_add_7_25_groupi_n_6014);
  xnor csa_tree_add_7_25_groupi_g15058(out2[11] ,csa_tree_add_7_25_groupi_n_5889 ,csa_tree_add_7_25_groupi_n_5892);
  xnor csa_tree_add_7_25_groupi_g15059(csa_tree_add_7_25_groupi_n_6011 ,csa_tree_add_7_25_groupi_n_5914 ,csa_tree_add_7_25_groupi_n_5867);
  xnor csa_tree_add_7_25_groupi_g15060(csa_tree_add_7_25_groupi_n_6010 ,csa_tree_add_7_25_groupi_n_5901 ,csa_tree_add_7_25_groupi_n_5887);
  xnor csa_tree_add_7_25_groupi_g15061(csa_tree_add_7_25_groupi_n_6009 ,csa_tree_add_7_25_groupi_n_5847 ,csa_tree_add_7_25_groupi_n_5917);
  xnor csa_tree_add_7_25_groupi_g15062(csa_tree_add_7_25_groupi_n_6008 ,csa_tree_add_7_25_groupi_n_5905 ,csa_tree_add_7_25_groupi_n_5866);
  xnor csa_tree_add_7_25_groupi_g15063(csa_tree_add_7_25_groupi_n_6007 ,csa_tree_add_7_25_groupi_n_5869 ,csa_tree_add_7_25_groupi_n_5903);
  xnor csa_tree_add_7_25_groupi_g15064(csa_tree_add_7_25_groupi_n_6006 ,csa_tree_add_7_25_groupi_n_5848 ,csa_tree_add_7_25_groupi_n_5899);
  xnor csa_tree_add_7_25_groupi_g15065(csa_tree_add_7_25_groupi_n_6005 ,csa_tree_add_7_25_groupi_n_5844 ,csa_tree_add_7_25_groupi_n_5912);
  xnor csa_tree_add_7_25_groupi_g15066(csa_tree_add_7_25_groupi_n_6004 ,csa_tree_add_7_25_groupi_n_5845 ,csa_tree_add_7_25_groupi_n_5913);
  xnor csa_tree_add_7_25_groupi_g15067(csa_tree_add_7_25_groupi_n_6003 ,csa_tree_add_7_25_groupi_n_5846 ,csa_tree_add_7_25_groupi_n_5915);
  xnor csa_tree_add_7_25_groupi_g15068(csa_tree_add_7_25_groupi_n_6002 ,csa_tree_add_7_25_groupi_n_5890 ,csa_tree_add_7_25_groupi_n_5557);
  xnor csa_tree_add_7_25_groupi_g15069(csa_tree_add_7_25_groupi_n_6001 ,csa_tree_add_7_25_groupi_n_5843 ,csa_tree_add_7_25_groupi_n_5916);
  xnor csa_tree_add_7_25_groupi_g15070(csa_tree_add_7_25_groupi_n_6036 ,csa_tree_add_7_25_groupi_n_5935 ,in3[8]);
  xnor csa_tree_add_7_25_groupi_g15071(csa_tree_add_7_25_groupi_n_6035 ,csa_tree_add_7_25_groupi_n_5932 ,in3[5]);
  xnor csa_tree_add_7_25_groupi_g15072(csa_tree_add_7_25_groupi_n_6034 ,csa_tree_add_7_25_groupi_n_5928 ,in3[11]);
  xnor csa_tree_add_7_25_groupi_g15073(csa_tree_add_7_25_groupi_n_6033 ,csa_tree_add_7_25_groupi_n_5930 ,in3[14]);
  xnor csa_tree_add_7_25_groupi_g15074(csa_tree_add_7_25_groupi_n_6032 ,csa_tree_add_7_25_groupi_n_5931 ,in3[2]);
  xnor csa_tree_add_7_25_groupi_g15075(csa_tree_add_7_25_groupi_n_6031 ,csa_tree_add_7_25_groupi_n_5918 ,csa_tree_add_7_25_groupi_n_5795);
  xnor csa_tree_add_7_25_groupi_g15076(csa_tree_add_7_25_groupi_n_6030 ,csa_tree_add_7_25_groupi_n_5922 ,csa_tree_add_7_25_groupi_n_5793);
  xnor csa_tree_add_7_25_groupi_g15077(csa_tree_add_7_25_groupi_n_6028 ,csa_tree_add_7_25_groupi_n_5923 ,csa_tree_add_7_25_groupi_n_5791);
  xnor csa_tree_add_7_25_groupi_g15078(csa_tree_add_7_25_groupi_n_6027 ,csa_tree_add_7_25_groupi_n_5926 ,csa_tree_add_7_25_groupi_n_5797);
  xnor csa_tree_add_7_25_groupi_g15079(csa_tree_add_7_25_groupi_n_6025 ,csa_tree_add_7_25_groupi_n_5924 ,csa_tree_add_7_25_groupi_n_5792);
  xnor csa_tree_add_7_25_groupi_g15080(csa_tree_add_7_25_groupi_n_6024 ,csa_tree_add_7_25_groupi_n_5920 ,csa_tree_add_7_25_groupi_n_5787);
  xnor csa_tree_add_7_25_groupi_g15081(csa_tree_add_7_25_groupi_n_6023 ,csa_tree_add_7_25_groupi_n_5919 ,csa_tree_add_7_25_groupi_n_5788);
  xnor csa_tree_add_7_25_groupi_g15082(csa_tree_add_7_25_groupi_n_6022 ,csa_tree_add_7_25_groupi_n_5925 ,csa_tree_add_7_25_groupi_n_5789);
  xnor csa_tree_add_7_25_groupi_g15083(csa_tree_add_7_25_groupi_n_6021 ,csa_tree_add_7_25_groupi_n_5934 ,in3[17]);
  xnor csa_tree_add_7_25_groupi_g15084(csa_tree_add_7_25_groupi_n_6020 ,csa_tree_add_7_25_groupi_n_5921 ,csa_tree_add_7_25_groupi_n_5794);
  xnor csa_tree_add_7_25_groupi_g15085(csa_tree_add_7_25_groupi_n_6018 ,csa_tree_add_7_25_groupi_n_5929 ,in3[20]);
  xnor csa_tree_add_7_25_groupi_g15086(csa_tree_add_7_25_groupi_n_6016 ,csa_tree_add_7_25_groupi_n_5936 ,in3[26]);
  xnor csa_tree_add_7_25_groupi_g15087(csa_tree_add_7_25_groupi_n_6014 ,csa_tree_add_7_25_groupi_n_5927 ,in3[23]);
  or csa_tree_add_7_25_groupi_g15088(csa_tree_add_7_25_groupi_n_5999 ,csa_tree_add_7_25_groupi_n_5914 ,csa_tree_add_7_25_groupi_n_5867);
  or csa_tree_add_7_25_groupi_g15089(csa_tree_add_7_25_groupi_n_5998 ,csa_tree_add_7_25_groupi_n_5847 ,csa_tree_add_7_25_groupi_n_5917);
  and csa_tree_add_7_25_groupi_g15090(csa_tree_add_7_25_groupi_n_5997 ,csa_tree_add_7_25_groupi_n_5925 ,csa_tree_add_7_25_groupi_n_5765);
  and csa_tree_add_7_25_groupi_g15091(csa_tree_add_7_25_groupi_n_5996 ,csa_tree_add_7_25_groupi_n_5847 ,csa_tree_add_7_25_groupi_n_5917);
  and csa_tree_add_7_25_groupi_g15092(csa_tree_add_7_25_groupi_n_5995 ,csa_tree_add_7_25_groupi_n_5914 ,csa_tree_add_7_25_groupi_n_5867);
  and csa_tree_add_7_25_groupi_g15093(csa_tree_add_7_25_groupi_n_5994 ,csa_tree_add_7_25_groupi_n_5848 ,csa_tree_add_7_25_groupi_n_5899);
  or csa_tree_add_7_25_groupi_g15094(csa_tree_add_7_25_groupi_n_5993 ,csa_tree_add_7_25_groupi_n_5848 ,csa_tree_add_7_25_groupi_n_5899);
  and csa_tree_add_7_25_groupi_g15095(csa_tree_add_7_25_groupi_n_5992 ,csa_tree_add_7_25_groupi_n_5918 ,csa_tree_add_7_25_groupi_n_5780);
  and csa_tree_add_7_25_groupi_g15096(csa_tree_add_7_25_groupi_n_5991 ,csa_tree_add_7_25_groupi_n_5920 ,csa_tree_add_7_25_groupi_n_5777);
  and csa_tree_add_7_25_groupi_g15097(csa_tree_add_7_25_groupi_n_5990 ,csa_tree_add_7_25_groupi_n_5926 ,csa_tree_add_7_25_groupi_n_5743);
  and csa_tree_add_7_25_groupi_g15098(csa_tree_add_7_25_groupi_n_5989 ,csa_tree_add_7_25_groupi_n_5844 ,csa_tree_add_7_25_groupi_n_5912);
  or csa_tree_add_7_25_groupi_g15099(csa_tree_add_7_25_groupi_n_5988 ,csa_tree_add_7_25_groupi_n_5844 ,csa_tree_add_7_25_groupi_n_5912);
  and csa_tree_add_7_25_groupi_g15100(csa_tree_add_7_25_groupi_n_5987 ,csa_tree_add_7_25_groupi_n_5924 ,csa_tree_add_7_25_groupi_n_5773);
  and csa_tree_add_7_25_groupi_g15101(csa_tree_add_7_25_groupi_n_5986 ,csa_tree_add_7_25_groupi_n_5919 ,csa_tree_add_7_25_groupi_n_5770);
  or csa_tree_add_7_25_groupi_g15102(csa_tree_add_7_25_groupi_n_5985 ,csa_tree_add_7_25_groupi_n_5845 ,csa_tree_add_7_25_groupi_n_5913);
  and csa_tree_add_7_25_groupi_g15103(csa_tree_add_7_25_groupi_n_5984 ,csa_tree_add_7_25_groupi_n_5923 ,csa_tree_add_7_25_groupi_n_5767);
  and csa_tree_add_7_25_groupi_g15104(csa_tree_add_7_25_groupi_n_5983 ,csa_tree_add_7_25_groupi_n_5845 ,csa_tree_add_7_25_groupi_n_5913);
  and csa_tree_add_7_25_groupi_g15105(csa_tree_add_7_25_groupi_n_5982 ,csa_tree_add_7_25_groupi_n_5846 ,csa_tree_add_7_25_groupi_n_5915);
  or csa_tree_add_7_25_groupi_g15106(csa_tree_add_7_25_groupi_n_5981 ,csa_tree_add_7_25_groupi_n_5846 ,csa_tree_add_7_25_groupi_n_5915);
  and csa_tree_add_7_25_groupi_g15107(csa_tree_add_7_25_groupi_n_6000 ,csa_tree_add_7_25_groupi_n_2428 ,csa_tree_add_7_25_groupi_n_5941);
  or csa_tree_add_7_25_groupi_g15108(csa_tree_add_7_25_groupi_n_5978 ,csa_tree_add_7_25_groupi_n_5900 ,csa_tree_add_7_25_groupi_n_5887);
  nor csa_tree_add_7_25_groupi_g15109(csa_tree_add_7_25_groupi_n_5977 ,csa_tree_add_7_25_groupi_n_5868 ,csa_tree_add_7_25_groupi_n_5903);
  or csa_tree_add_7_25_groupi_g15110(csa_tree_add_7_25_groupi_n_5976 ,csa_tree_add_7_25_groupi_n_5869 ,csa_tree_add_7_25_groupi_n_5902);
  or csa_tree_add_7_25_groupi_g15111(csa_tree_add_7_25_groupi_n_5975 ,csa_tree_add_7_25_groupi_n_3319 ,csa_tree_add_7_25_groupi_n_5944);
  or csa_tree_add_7_25_groupi_g15112(csa_tree_add_7_25_groupi_n_5974 ,csa_tree_add_7_25_groupi_n_3315 ,csa_tree_add_7_25_groupi_n_5945);
  or csa_tree_add_7_25_groupi_g15113(csa_tree_add_7_25_groupi_n_5973 ,csa_tree_add_7_25_groupi_n_3313 ,csa_tree_add_7_25_groupi_n_5947);
  or csa_tree_add_7_25_groupi_g15114(csa_tree_add_7_25_groupi_n_5972 ,csa_tree_add_7_25_groupi_n_3698 ,csa_tree_add_7_25_groupi_n_5939);
  or csa_tree_add_7_25_groupi_g15115(csa_tree_add_7_25_groupi_n_5971 ,csa_tree_add_7_25_groupi_n_3699 ,csa_tree_add_7_25_groupi_n_5940);
  nor csa_tree_add_7_25_groupi_g15116(csa_tree_add_7_25_groupi_n_5970 ,csa_tree_add_7_25_groupi_n_5905 ,csa_tree_add_7_25_groupi_n_5865);
  or csa_tree_add_7_25_groupi_g15117(csa_tree_add_7_25_groupi_n_5969 ,csa_tree_add_7_25_groupi_n_5904 ,csa_tree_add_7_25_groupi_n_5866);
  and csa_tree_add_7_25_groupi_g15118(csa_tree_add_7_25_groupi_n_5968 ,csa_tree_add_7_25_groupi_n_5922 ,csa_tree_add_7_25_groupi_n_5760);
  or csa_tree_add_7_25_groupi_g15119(csa_tree_add_7_25_groupi_n_5967 ,csa_tree_add_7_25_groupi_n_3700 ,csa_tree_add_7_25_groupi_n_5942);
  or csa_tree_add_7_25_groupi_g15120(csa_tree_add_7_25_groupi_n_5966 ,csa_tree_add_7_25_groupi_n_3703 ,csa_tree_add_7_25_groupi_n_5943);
  or csa_tree_add_7_25_groupi_g15121(csa_tree_add_7_25_groupi_n_5965 ,csa_tree_add_7_25_groupi_n_3701 ,csa_tree_add_7_25_groupi_n_5946);
  and csa_tree_add_7_25_groupi_g15122(csa_tree_add_7_25_groupi_n_5964 ,csa_tree_add_7_25_groupi_n_5921 ,csa_tree_add_7_25_groupi_n_5751);
  and csa_tree_add_7_25_groupi_g15123(csa_tree_add_7_25_groupi_n_5963 ,csa_tree_add_7_25_groupi_n_5843 ,csa_tree_add_7_25_groupi_n_5916);
  or csa_tree_add_7_25_groupi_g15124(csa_tree_add_7_25_groupi_n_5962 ,csa_tree_add_7_25_groupi_n_5843 ,csa_tree_add_7_25_groupi_n_5916);
  nor csa_tree_add_7_25_groupi_g15125(csa_tree_add_7_25_groupi_n_5961 ,csa_tree_add_7_25_groupi_n_5901 ,csa_tree_add_7_25_groupi_n_5886);
  or csa_tree_add_7_25_groupi_g15126(csa_tree_add_7_25_groupi_n_5960 ,csa_tree_add_7_25_groupi_n_3229 ,csa_tree_add_7_25_groupi_n_5938);
  or csa_tree_add_7_25_groupi_g15127(csa_tree_add_7_25_groupi_n_5980 ,csa_tree_add_7_25_groupi_n_5937 ,csa_tree_add_7_25_groupi_n_5850);
  xnor csa_tree_add_7_25_groupi_g15128(csa_tree_add_7_25_groupi_n_5979 ,csa_tree_add_7_25_groupi_n_5888 ,csa_tree_add_7_25_groupi_n_2568);
  not csa_tree_add_7_25_groupi_g15129(csa_tree_add_7_25_groupi_n_5956 ,csa_tree_add_7_25_groupi_n_5957);
  not csa_tree_add_7_25_groupi_g15130(csa_tree_add_7_25_groupi_n_5954 ,csa_tree_add_7_25_groupi_n_5955);
  not csa_tree_add_7_25_groupi_g15131(csa_tree_add_7_25_groupi_n_5949 ,csa_tree_add_7_25_groupi_n_5950);
  nor csa_tree_add_7_25_groupi_g15132(csa_tree_add_7_25_groupi_n_5947 ,csa_tree_add_7_25_groupi_n_2103 ,csa_tree_add_7_25_groupi_n_1808);
  nor csa_tree_add_7_25_groupi_g15133(csa_tree_add_7_25_groupi_n_5946 ,csa_tree_add_7_25_groupi_n_2157 ,csa_tree_add_7_25_groupi_n_1256);
  nor csa_tree_add_7_25_groupi_g15134(csa_tree_add_7_25_groupi_n_5945 ,csa_tree_add_7_25_groupi_n_2124 ,csa_tree_add_7_25_groupi_n_1255);
  nor csa_tree_add_7_25_groupi_g15135(csa_tree_add_7_25_groupi_n_5944 ,csa_tree_add_7_25_groupi_n_2142 ,csa_tree_add_7_25_groupi_n_154);
  nor csa_tree_add_7_25_groupi_g15136(csa_tree_add_7_25_groupi_n_5943 ,csa_tree_add_7_25_groupi_n_2058 ,csa_tree_add_7_25_groupi_n_1256);
  nor csa_tree_add_7_25_groupi_g15137(csa_tree_add_7_25_groupi_n_5942 ,csa_tree_add_7_25_groupi_n_2049 ,csa_tree_add_7_25_groupi_n_155);
  or csa_tree_add_7_25_groupi_g15138(csa_tree_add_7_25_groupi_n_5941 ,csa_tree_add_7_25_groupi_n_2485 ,csa_tree_add_7_25_groupi_n_5888);
  nor csa_tree_add_7_25_groupi_g15139(csa_tree_add_7_25_groupi_n_5940 ,csa_tree_add_7_25_groupi_n_2031 ,csa_tree_add_7_25_groupi_n_1808);
  nor csa_tree_add_7_25_groupi_g15140(csa_tree_add_7_25_groupi_n_5939 ,csa_tree_add_7_25_groupi_n_554 ,csa_tree_add_7_25_groupi_n_1255);
  nor csa_tree_add_7_25_groupi_g15141(csa_tree_add_7_25_groupi_n_5938 ,csa_tree_add_7_25_groupi_n_2184 ,csa_tree_add_7_25_groupi_n_155);
  and csa_tree_add_7_25_groupi_g15142(csa_tree_add_7_25_groupi_n_5937 ,csa_tree_add_7_25_groupi_n_5889 ,csa_tree_add_7_25_groupi_n_5849);
  nor csa_tree_add_7_25_groupi_g15143(csa_tree_add_7_25_groupi_n_5936 ,csa_tree_add_7_25_groupi_n_3852 ,csa_tree_add_7_25_groupi_n_5859);
  nor csa_tree_add_7_25_groupi_g15144(csa_tree_add_7_25_groupi_n_5935 ,csa_tree_add_7_25_groupi_n_4094 ,csa_tree_add_7_25_groupi_n_5861);
  nor csa_tree_add_7_25_groupi_g15145(csa_tree_add_7_25_groupi_n_5934 ,csa_tree_add_7_25_groupi_n_3894 ,csa_tree_add_7_25_groupi_n_5863);
  or csa_tree_add_7_25_groupi_g15146(csa_tree_add_7_25_groupi_n_5933 ,csa_tree_add_7_25_groupi_n_5444 ,csa_tree_add_7_25_groupi_n_5884);
  nor csa_tree_add_7_25_groupi_g15147(csa_tree_add_7_25_groupi_n_5932 ,csa_tree_add_7_25_groupi_n_4064 ,csa_tree_add_7_25_groupi_n_5862);
  nor csa_tree_add_7_25_groupi_g15148(csa_tree_add_7_25_groupi_n_5931 ,csa_tree_add_7_25_groupi_n_3467 ,csa_tree_add_7_25_groupi_n_5857);
  nor csa_tree_add_7_25_groupi_g15149(csa_tree_add_7_25_groupi_n_5930 ,csa_tree_add_7_25_groupi_n_3883 ,csa_tree_add_7_25_groupi_n_5853);
  nor csa_tree_add_7_25_groupi_g15150(csa_tree_add_7_25_groupi_n_5929 ,csa_tree_add_7_25_groupi_n_3856 ,csa_tree_add_7_25_groupi_n_5855);
  nor csa_tree_add_7_25_groupi_g15151(csa_tree_add_7_25_groupi_n_5928 ,csa_tree_add_7_25_groupi_n_4000 ,csa_tree_add_7_25_groupi_n_5860);
  nor csa_tree_add_7_25_groupi_g15152(csa_tree_add_7_25_groupi_n_5927 ,csa_tree_add_7_25_groupi_n_3840 ,csa_tree_add_7_25_groupi_n_5856);
  or csa_tree_add_7_25_groupi_g15153(csa_tree_add_7_25_groupi_n_5959 ,csa_tree_add_7_25_groupi_n_5660 ,csa_tree_add_7_25_groupi_n_5880);
  or csa_tree_add_7_25_groupi_g15154(csa_tree_add_7_25_groupi_n_5958 ,csa_tree_add_7_25_groupi_n_5631 ,csa_tree_add_7_25_groupi_n_5852);
  or csa_tree_add_7_25_groupi_g15155(csa_tree_add_7_25_groupi_n_5957 ,csa_tree_add_7_25_groupi_n_5642 ,csa_tree_add_7_25_groupi_n_5858);
  or csa_tree_add_7_25_groupi_g15156(csa_tree_add_7_25_groupi_n_5955 ,csa_tree_add_7_25_groupi_n_5645 ,csa_tree_add_7_25_groupi_n_5883);
  or csa_tree_add_7_25_groupi_g15157(csa_tree_add_7_25_groupi_n_5953 ,csa_tree_add_7_25_groupi_n_5669 ,csa_tree_add_7_25_groupi_n_5873);
  or csa_tree_add_7_25_groupi_g15158(csa_tree_add_7_25_groupi_n_5952 ,csa_tree_add_7_25_groupi_n_5651 ,csa_tree_add_7_25_groupi_n_5885);
  or csa_tree_add_7_25_groupi_g15159(csa_tree_add_7_25_groupi_n_5951 ,csa_tree_add_7_25_groupi_n_5655 ,csa_tree_add_7_25_groupi_n_5879);
  or csa_tree_add_7_25_groupi_g15160(csa_tree_add_7_25_groupi_n_5950 ,csa_tree_add_7_25_groupi_n_5668 ,csa_tree_add_7_25_groupi_n_5876);
  or csa_tree_add_7_25_groupi_g15161(csa_tree_add_7_25_groupi_n_5948 ,csa_tree_add_7_25_groupi_n_5663 ,csa_tree_add_7_25_groupi_n_5881);
  not csa_tree_add_7_25_groupi_g15162(csa_tree_add_7_25_groupi_n_5910 ,csa_tree_add_7_25_groupi_n_5911);
  not csa_tree_add_7_25_groupi_g15163(csa_tree_add_7_25_groupi_n_5908 ,csa_tree_add_7_25_groupi_n_5909);
  not csa_tree_add_7_25_groupi_g15164(csa_tree_add_7_25_groupi_n_5906 ,csa_tree_add_7_25_groupi_n_5907);
  not csa_tree_add_7_25_groupi_g15165(csa_tree_add_7_25_groupi_n_5904 ,csa_tree_add_7_25_groupi_n_5905);
  not csa_tree_add_7_25_groupi_g15166(csa_tree_add_7_25_groupi_n_5902 ,csa_tree_add_7_25_groupi_n_5903);
  not csa_tree_add_7_25_groupi_g15167(csa_tree_add_7_25_groupi_n_5900 ,csa_tree_add_7_25_groupi_n_5901);
  xnor csa_tree_add_7_25_groupi_g15168(out2[10] ,csa_tree_add_7_25_groupi_n_5785 ,csa_tree_add_7_25_groupi_n_5796);
  xnor csa_tree_add_7_25_groupi_g15169(csa_tree_add_7_25_groupi_n_5896 ,csa_tree_add_7_25_groupi_n_5735 ,csa_tree_add_7_25_groupi_n_5802);
  xnor csa_tree_add_7_25_groupi_g15170(csa_tree_add_7_25_groupi_n_5895 ,csa_tree_add_7_25_groupi_n_5731 ,csa_tree_add_7_25_groupi_n_5803);
  xnor csa_tree_add_7_25_groupi_g15171(csa_tree_add_7_25_groupi_n_5894 ,csa_tree_add_7_25_groupi_n_5730 ,csa_tree_add_7_25_groupi_n_5805);
  xnor csa_tree_add_7_25_groupi_g15172(csa_tree_add_7_25_groupi_n_5893 ,csa_tree_add_7_25_groupi_n_5804 ,csa_tree_add_7_25_groupi_n_5734);
  xnor csa_tree_add_7_25_groupi_g15173(csa_tree_add_7_25_groupi_n_5892 ,csa_tree_add_7_25_groupi_n_5732 ,csa_tree_add_7_25_groupi_n_5807);
  xnor csa_tree_add_7_25_groupi_g15174(csa_tree_add_7_25_groupi_n_5891 ,csa_tree_add_7_25_groupi_n_5733 ,csa_tree_add_7_25_groupi_n_5806);
  xnor csa_tree_add_7_25_groupi_g15175(csa_tree_add_7_25_groupi_n_5890 ,csa_tree_add_7_25_groupi_n_5820 ,in3[29]);
  xnor csa_tree_add_7_25_groupi_g15176(csa_tree_add_7_25_groupi_n_5926 ,csa_tree_add_7_25_groupi_n_5824 ,in3[26]);
  xnor csa_tree_add_7_25_groupi_g15177(csa_tree_add_7_25_groupi_n_5925 ,csa_tree_add_7_25_groupi_n_5822 ,in3[11]);
  xnor csa_tree_add_7_25_groupi_g15178(csa_tree_add_7_25_groupi_n_5924 ,csa_tree_add_7_25_groupi_n_5819 ,in3[5]);
  xnor csa_tree_add_7_25_groupi_g15179(csa_tree_add_7_25_groupi_n_5923 ,csa_tree_add_7_25_groupi_n_5818 ,in3[8]);
  xnor csa_tree_add_7_25_groupi_g15180(csa_tree_add_7_25_groupi_n_5922 ,csa_tree_add_7_25_groupi_n_5821 ,in3[23]);
  xnor csa_tree_add_7_25_groupi_g15181(csa_tree_add_7_25_groupi_n_5921 ,csa_tree_add_7_25_groupi_n_5823 ,in3[20]);
  xnor csa_tree_add_7_25_groupi_g15182(csa_tree_add_7_25_groupi_n_5920 ,csa_tree_add_7_25_groupi_n_5827 ,in3[17]);
  xnor csa_tree_add_7_25_groupi_g15183(csa_tree_add_7_25_groupi_n_5919 ,csa_tree_add_7_25_groupi_n_5826 ,in3[14]);
  xnor csa_tree_add_7_25_groupi_g15184(csa_tree_add_7_25_groupi_n_5918 ,csa_tree_add_7_25_groupi_n_5825 ,in3[2]);
  xnor csa_tree_add_7_25_groupi_g15185(csa_tree_add_7_25_groupi_n_5917 ,csa_tree_add_7_25_groupi_n_5816 ,csa_tree_add_7_25_groupi_n_5678);
  xnor csa_tree_add_7_25_groupi_g15186(csa_tree_add_7_25_groupi_n_5916 ,csa_tree_add_7_25_groupi_n_5817 ,csa_tree_add_7_25_groupi_n_5674);
  xnor csa_tree_add_7_25_groupi_g15187(csa_tree_add_7_25_groupi_n_5915 ,csa_tree_add_7_25_groupi_n_5815 ,csa_tree_add_7_25_groupi_n_5671);
  xnor csa_tree_add_7_25_groupi_g15188(csa_tree_add_7_25_groupi_n_5914 ,csa_tree_add_7_25_groupi_n_5810 ,csa_tree_add_7_25_groupi_n_5680);
  xnor csa_tree_add_7_25_groupi_g15189(csa_tree_add_7_25_groupi_n_5913 ,csa_tree_add_7_25_groupi_n_5809 ,csa_tree_add_7_25_groupi_n_5675);
  xnor csa_tree_add_7_25_groupi_g15190(csa_tree_add_7_25_groupi_n_5912 ,csa_tree_add_7_25_groupi_n_5814 ,csa_tree_add_7_25_groupi_n_5676);
  xnor csa_tree_add_7_25_groupi_g15191(csa_tree_add_7_25_groupi_n_5911 ,csa_tree_add_7_25_groupi_n_5739 ,csa_tree_add_7_25_groupi_n_5800);
  xnor csa_tree_add_7_25_groupi_g15192(csa_tree_add_7_25_groupi_n_5909 ,csa_tree_add_7_25_groupi_n_5736 ,csa_tree_add_7_25_groupi_n_5799);
  xnor csa_tree_add_7_25_groupi_g15193(csa_tree_add_7_25_groupi_n_5907 ,csa_tree_add_7_25_groupi_n_5738 ,csa_tree_add_7_25_groupi_n_5798);
  xnor csa_tree_add_7_25_groupi_g15194(csa_tree_add_7_25_groupi_n_5905 ,csa_tree_add_7_25_groupi_n_5811 ,csa_tree_add_7_25_groupi_n_5673);
  xnor csa_tree_add_7_25_groupi_g15195(csa_tree_add_7_25_groupi_n_5903 ,csa_tree_add_7_25_groupi_n_5812 ,csa_tree_add_7_25_groupi_n_5672);
  xnor csa_tree_add_7_25_groupi_g15196(csa_tree_add_7_25_groupi_n_5901 ,csa_tree_add_7_25_groupi_n_5808 ,csa_tree_add_7_25_groupi_n_5455);
  xnor csa_tree_add_7_25_groupi_g15197(csa_tree_add_7_25_groupi_n_5899 ,csa_tree_add_7_25_groupi_n_5813 ,csa_tree_add_7_25_groupi_n_5677);
  xnor csa_tree_add_7_25_groupi_g15198(csa_tree_add_7_25_groupi_n_5898 ,csa_tree_add_7_25_groupi_n_5737 ,csa_tree_add_7_25_groupi_n_5790);
  not csa_tree_add_7_25_groupi_g15199(csa_tree_add_7_25_groupi_n_5886 ,csa_tree_add_7_25_groupi_n_5887);
  and csa_tree_add_7_25_groupi_g15200(csa_tree_add_7_25_groupi_n_5885 ,csa_tree_add_7_25_groupi_n_5809 ,csa_tree_add_7_25_groupi_n_5650);
  and csa_tree_add_7_25_groupi_g15201(csa_tree_add_7_25_groupi_n_5884 ,csa_tree_add_7_25_groupi_n_5808 ,csa_tree_add_7_25_groupi_n_5443);
  and csa_tree_add_7_25_groupi_g15202(csa_tree_add_7_25_groupi_n_5883 ,csa_tree_add_7_25_groupi_n_5812 ,csa_tree_add_7_25_groupi_n_5644);
  or csa_tree_add_7_25_groupi_g15203(csa_tree_add_7_25_groupi_n_5882 ,csa_tree_add_7_25_groupi_n_5730 ,csa_tree_add_7_25_groupi_n_5805);
  and csa_tree_add_7_25_groupi_g15204(csa_tree_add_7_25_groupi_n_5881 ,csa_tree_add_7_25_groupi_n_5816 ,csa_tree_add_7_25_groupi_n_5661);
  and csa_tree_add_7_25_groupi_g15205(csa_tree_add_7_25_groupi_n_5880 ,csa_tree_add_7_25_groupi_n_5813 ,csa_tree_add_7_25_groupi_n_5659);
  and csa_tree_add_7_25_groupi_g15206(csa_tree_add_7_25_groupi_n_5879 ,csa_tree_add_7_25_groupi_n_5814 ,csa_tree_add_7_25_groupi_n_5653);
  and csa_tree_add_7_25_groupi_g15207(csa_tree_add_7_25_groupi_n_5878 ,csa_tree_add_7_25_groupi_n_5735 ,csa_tree_add_7_25_groupi_n_5802);
  or csa_tree_add_7_25_groupi_g15208(csa_tree_add_7_25_groupi_n_5877 ,csa_tree_add_7_25_groupi_n_5735 ,csa_tree_add_7_25_groupi_n_5802);
  and csa_tree_add_7_25_groupi_g15209(csa_tree_add_7_25_groupi_n_5876 ,csa_tree_add_7_25_groupi_n_5810 ,csa_tree_add_7_25_groupi_n_5667);
  and csa_tree_add_7_25_groupi_g15210(csa_tree_add_7_25_groupi_n_5875 ,csa_tree_add_7_25_groupi_n_5804 ,csa_tree_add_7_25_groupi_n_5734);
  or csa_tree_add_7_25_groupi_g15211(csa_tree_add_7_25_groupi_n_5874 ,csa_tree_add_7_25_groupi_n_5804 ,csa_tree_add_7_25_groupi_n_5734);
  and csa_tree_add_7_25_groupi_g15212(csa_tree_add_7_25_groupi_n_5873 ,csa_tree_add_7_25_groupi_n_5815 ,csa_tree_add_7_25_groupi_n_5636);
  and csa_tree_add_7_25_groupi_g15213(csa_tree_add_7_25_groupi_n_5872 ,csa_tree_add_7_25_groupi_n_5731 ,csa_tree_add_7_25_groupi_n_5803);
  or csa_tree_add_7_25_groupi_g15214(csa_tree_add_7_25_groupi_n_5871 ,csa_tree_add_7_25_groupi_n_5731 ,csa_tree_add_7_25_groupi_n_5803);
  and csa_tree_add_7_25_groupi_g15215(csa_tree_add_7_25_groupi_n_5870 ,csa_tree_add_7_25_groupi_n_5730 ,csa_tree_add_7_25_groupi_n_5805);
  or csa_tree_add_7_25_groupi_g15216(csa_tree_add_7_25_groupi_n_5889 ,csa_tree_add_7_25_groupi_n_5782 ,csa_tree_add_7_25_groupi_n_5835);
  and csa_tree_add_7_25_groupi_g15217(csa_tree_add_7_25_groupi_n_5888 ,csa_tree_add_7_25_groupi_n_2440 ,csa_tree_add_7_25_groupi_n_5841);
  or csa_tree_add_7_25_groupi_g15218(csa_tree_add_7_25_groupi_n_5887 ,csa_tree_add_7_25_groupi_n_5764 ,csa_tree_add_7_25_groupi_n_5836);
  not csa_tree_add_7_25_groupi_g15219(csa_tree_add_7_25_groupi_n_5868 ,csa_tree_add_7_25_groupi_n_5869);
  not csa_tree_add_7_25_groupi_g15220(csa_tree_add_7_25_groupi_n_5865 ,csa_tree_add_7_25_groupi_n_5866);
  or csa_tree_add_7_25_groupi_g15221(csa_tree_add_7_25_groupi_n_5863 ,csa_tree_add_7_25_groupi_n_3695 ,csa_tree_add_7_25_groupi_n_5832);
  or csa_tree_add_7_25_groupi_g15222(csa_tree_add_7_25_groupi_n_5862 ,csa_tree_add_7_25_groupi_n_3299 ,csa_tree_add_7_25_groupi_n_5837);
  or csa_tree_add_7_25_groupi_g15223(csa_tree_add_7_25_groupi_n_5861 ,csa_tree_add_7_25_groupi_n_3294 ,csa_tree_add_7_25_groupi_n_5838);
  or csa_tree_add_7_25_groupi_g15224(csa_tree_add_7_25_groupi_n_5860 ,csa_tree_add_7_25_groupi_n_3296 ,csa_tree_add_7_25_groupi_n_5840);
  or csa_tree_add_7_25_groupi_g15225(csa_tree_add_7_25_groupi_n_5859 ,csa_tree_add_7_25_groupi_n_3691 ,csa_tree_add_7_25_groupi_n_5829);
  and csa_tree_add_7_25_groupi_g15226(csa_tree_add_7_25_groupi_n_5858 ,csa_tree_add_7_25_groupi_n_5811 ,csa_tree_add_7_25_groupi_n_5641);
  or csa_tree_add_7_25_groupi_g15227(csa_tree_add_7_25_groupi_n_5857 ,csa_tree_add_7_25_groupi_n_3189 ,csa_tree_add_7_25_groupi_n_5830);
  or csa_tree_add_7_25_groupi_g15228(csa_tree_add_7_25_groupi_n_5856 ,csa_tree_add_7_25_groupi_n_3692 ,csa_tree_add_7_25_groupi_n_5828);
  or csa_tree_add_7_25_groupi_g15229(csa_tree_add_7_25_groupi_n_5855 ,csa_tree_add_7_25_groupi_n_3693 ,csa_tree_add_7_25_groupi_n_5831);
  or csa_tree_add_7_25_groupi_g15230(csa_tree_add_7_25_groupi_n_5854 ,csa_tree_add_7_25_groupi_n_5733 ,csa_tree_add_7_25_groupi_n_5806);
  or csa_tree_add_7_25_groupi_g15231(csa_tree_add_7_25_groupi_n_5853 ,csa_tree_add_7_25_groupi_n_3690 ,csa_tree_add_7_25_groupi_n_5839);
  and csa_tree_add_7_25_groupi_g15232(csa_tree_add_7_25_groupi_n_5852 ,csa_tree_add_7_25_groupi_n_5817 ,csa_tree_add_7_25_groupi_n_5630);
  and csa_tree_add_7_25_groupi_g15233(csa_tree_add_7_25_groupi_n_5851 ,csa_tree_add_7_25_groupi_n_5733 ,csa_tree_add_7_25_groupi_n_5806);
  and csa_tree_add_7_25_groupi_g15234(csa_tree_add_7_25_groupi_n_5850 ,csa_tree_add_7_25_groupi_n_5732 ,csa_tree_add_7_25_groupi_n_5807);
  or csa_tree_add_7_25_groupi_g15235(csa_tree_add_7_25_groupi_n_5849 ,csa_tree_add_7_25_groupi_n_5732 ,csa_tree_add_7_25_groupi_n_5807);
  or csa_tree_add_7_25_groupi_g15236(csa_tree_add_7_25_groupi_n_5869 ,csa_tree_add_7_25_groupi_n_5784 ,csa_tree_add_7_25_groupi_n_5842);
  or csa_tree_add_7_25_groupi_g15237(csa_tree_add_7_25_groupi_n_5867 ,csa_tree_add_7_25_groupi_n_5747 ,csa_tree_add_7_25_groupi_n_5833);
  or csa_tree_add_7_25_groupi_g15238(csa_tree_add_7_25_groupi_n_5866 ,csa_tree_add_7_25_groupi_n_5754 ,csa_tree_add_7_25_groupi_n_5834);
  xnor csa_tree_add_7_25_groupi_g15239(csa_tree_add_7_25_groupi_n_5864 ,csa_tree_add_7_25_groupi_n_5786 ,csa_tree_add_7_25_groupi_n_2569);
  and csa_tree_add_7_25_groupi_g15240(csa_tree_add_7_25_groupi_n_5842 ,csa_tree_add_7_25_groupi_n_5736 ,csa_tree_add_7_25_groupi_n_5762);
  or csa_tree_add_7_25_groupi_g15241(csa_tree_add_7_25_groupi_n_5841 ,csa_tree_add_7_25_groupi_n_2497 ,csa_tree_add_7_25_groupi_n_5786);
  nor csa_tree_add_7_25_groupi_g15242(csa_tree_add_7_25_groupi_n_5840 ,csa_tree_add_7_25_groupi_n_2103 ,csa_tree_add_7_25_groupi_n_196);
  nor csa_tree_add_7_25_groupi_g15243(csa_tree_add_7_25_groupi_n_5839 ,csa_tree_add_7_25_groupi_n_2157 ,csa_tree_add_7_25_groupi_n_1286);
  nor csa_tree_add_7_25_groupi_g15244(csa_tree_add_7_25_groupi_n_5838 ,csa_tree_add_7_25_groupi_n_2124 ,csa_tree_add_7_25_groupi_n_1285);
  nor csa_tree_add_7_25_groupi_g15245(csa_tree_add_7_25_groupi_n_5837 ,csa_tree_add_7_25_groupi_n_2142 ,csa_tree_add_7_25_groupi_n_1806);
  and csa_tree_add_7_25_groupi_g15246(csa_tree_add_7_25_groupi_n_5836 ,csa_tree_add_7_25_groupi_n_5738 ,csa_tree_add_7_25_groupi_n_5781);
  and csa_tree_add_7_25_groupi_g15247(csa_tree_add_7_25_groupi_n_5835 ,csa_tree_add_7_25_groupi_n_5783 ,csa_tree_add_7_25_groupi_n_5785);
  and csa_tree_add_7_25_groupi_g15248(csa_tree_add_7_25_groupi_n_5834 ,csa_tree_add_7_25_groupi_n_5739 ,csa_tree_add_7_25_groupi_n_5753);
  and csa_tree_add_7_25_groupi_g15249(csa_tree_add_7_25_groupi_n_5833 ,csa_tree_add_7_25_groupi_n_5746 ,csa_tree_add_7_25_groupi_n_5737);
  nor csa_tree_add_7_25_groupi_g15250(csa_tree_add_7_25_groupi_n_5832 ,csa_tree_add_7_25_groupi_n_2055 ,csa_tree_add_7_25_groupi_n_1286);
  nor csa_tree_add_7_25_groupi_g15251(csa_tree_add_7_25_groupi_n_5831 ,csa_tree_add_7_25_groupi_n_2040 ,csa_tree_add_7_25_groupi_n_196);
  nor csa_tree_add_7_25_groupi_g15252(csa_tree_add_7_25_groupi_n_5830 ,csa_tree_add_7_25_groupi_n_2184 ,csa_tree_add_7_25_groupi_n_1806);
  nor csa_tree_add_7_25_groupi_g15253(csa_tree_add_7_25_groupi_n_5829 ,csa_tree_add_7_25_groupi_n_1795 ,csa_tree_add_7_25_groupi_n_1285);
  nor csa_tree_add_7_25_groupi_g15254(csa_tree_add_7_25_groupi_n_5828 ,csa_tree_add_7_25_groupi_n_2021 ,csa_tree_add_7_25_groupi_n_195);
  nor csa_tree_add_7_25_groupi_g15255(csa_tree_add_7_25_groupi_n_5827 ,csa_tree_add_7_25_groupi_n_3934 ,csa_tree_add_7_25_groupi_n_5748);
  nor csa_tree_add_7_25_groupi_g15256(csa_tree_add_7_25_groupi_n_5826 ,csa_tree_add_7_25_groupi_n_3871 ,csa_tree_add_7_25_groupi_n_5745);
  nor csa_tree_add_7_25_groupi_g15257(csa_tree_add_7_25_groupi_n_5825 ,csa_tree_add_7_25_groupi_n_3387 ,csa_tree_add_7_25_groupi_n_5740);
  nor csa_tree_add_7_25_groupi_g15258(csa_tree_add_7_25_groupi_n_5824 ,csa_tree_add_7_25_groupi_n_3918 ,csa_tree_add_7_25_groupi_n_5750);
  nor csa_tree_add_7_25_groupi_g15259(csa_tree_add_7_25_groupi_n_5823 ,csa_tree_add_7_25_groupi_n_4096 ,csa_tree_add_7_25_groupi_n_5759);
  nor csa_tree_add_7_25_groupi_g15260(csa_tree_add_7_25_groupi_n_5822 ,csa_tree_add_7_25_groupi_n_3998 ,csa_tree_add_7_25_groupi_n_5756);
  nor csa_tree_add_7_25_groupi_g15261(csa_tree_add_7_25_groupi_n_5821 ,csa_tree_add_7_25_groupi_n_3900 ,csa_tree_add_7_25_groupi_n_5749);
  nor csa_tree_add_7_25_groupi_g15262(csa_tree_add_7_25_groupi_n_5820 ,csa_tree_add_7_25_groupi_n_3864 ,csa_tree_add_7_25_groupi_n_5755);
  nor csa_tree_add_7_25_groupi_g15263(csa_tree_add_7_25_groupi_n_5819 ,csa_tree_add_7_25_groupi_n_4060 ,csa_tree_add_7_25_groupi_n_5758);
  nor csa_tree_add_7_25_groupi_g15264(csa_tree_add_7_25_groupi_n_5818 ,csa_tree_add_7_25_groupi_n_4087 ,csa_tree_add_7_25_groupi_n_5757);
  or csa_tree_add_7_25_groupi_g15265(csa_tree_add_7_25_groupi_n_5848 ,csa_tree_add_7_25_groupi_n_5518 ,csa_tree_add_7_25_groupi_n_5741);
  or csa_tree_add_7_25_groupi_g15266(csa_tree_add_7_25_groupi_n_5847 ,csa_tree_add_7_25_groupi_n_5516 ,csa_tree_add_7_25_groupi_n_5742);
  or csa_tree_add_7_25_groupi_g15267(csa_tree_add_7_25_groupi_n_5846 ,csa_tree_add_7_25_groupi_n_5548 ,csa_tree_add_7_25_groupi_n_5769);
  or csa_tree_add_7_25_groupi_g15268(csa_tree_add_7_25_groupi_n_5845 ,csa_tree_add_7_25_groupi_n_5535 ,csa_tree_add_7_25_groupi_n_5772);
  or csa_tree_add_7_25_groupi_g15269(csa_tree_add_7_25_groupi_n_5844 ,csa_tree_add_7_25_groupi_n_5538 ,csa_tree_add_7_25_groupi_n_5775);
  or csa_tree_add_7_25_groupi_g15270(csa_tree_add_7_25_groupi_n_5843 ,csa_tree_add_7_25_groupi_n_5540 ,csa_tree_add_7_25_groupi_n_5776);
  xnor csa_tree_add_7_25_groupi_g15271(out2[9] ,csa_tree_add_7_25_groupi_n_5649 ,csa_tree_add_7_25_groupi_n_5679);
  xnor csa_tree_add_7_25_groupi_g15272(csa_tree_add_7_25_groupi_n_5800 ,csa_tree_add_7_25_groupi_n_5689 ,csa_tree_add_7_25_groupi_n_5571);
  xnor csa_tree_add_7_25_groupi_g15273(csa_tree_add_7_25_groupi_n_5799 ,csa_tree_add_7_25_groupi_n_5694 ,csa_tree_add_7_25_groupi_n_5573);
  xnor csa_tree_add_7_25_groupi_g15274(csa_tree_add_7_25_groupi_n_5798 ,csa_tree_add_7_25_groupi_n_5698 ,csa_tree_add_7_25_groupi_n_5464);
  xnor csa_tree_add_7_25_groupi_g15275(csa_tree_add_7_25_groupi_n_5797 ,csa_tree_add_7_25_groupi_n_5622 ,csa_tree_add_7_25_groupi_n_5687);
  xnor csa_tree_add_7_25_groupi_g15276(csa_tree_add_7_25_groupi_n_5796 ,csa_tree_add_7_25_groupi_n_5625 ,csa_tree_add_7_25_groupi_n_5692);
  xnor csa_tree_add_7_25_groupi_g15277(csa_tree_add_7_25_groupi_n_5795 ,csa_tree_add_7_25_groupi_n_5624 ,csa_tree_add_7_25_groupi_n_5691);
  xnor csa_tree_add_7_25_groupi_g15278(csa_tree_add_7_25_groupi_n_5794 ,csa_tree_add_7_25_groupi_n_5627 ,csa_tree_add_7_25_groupi_n_5685);
  xnor csa_tree_add_7_25_groupi_g15279(csa_tree_add_7_25_groupi_n_5793 ,csa_tree_add_7_25_groupi_n_5618 ,csa_tree_add_7_25_groupi_n_5696);
  xnor csa_tree_add_7_25_groupi_g15280(csa_tree_add_7_25_groupi_n_5792 ,csa_tree_add_7_25_groupi_n_5623 ,csa_tree_add_7_25_groupi_n_5690);
  xnor csa_tree_add_7_25_groupi_g15281(csa_tree_add_7_25_groupi_n_5791 ,csa_tree_add_7_25_groupi_n_5620 ,csa_tree_add_7_25_groupi_n_5699);
  xnor csa_tree_add_7_25_groupi_g15282(csa_tree_add_7_25_groupi_n_5790 ,csa_tree_add_7_25_groupi_n_5700 ,csa_tree_add_7_25_groupi_n_5578);
  xnor csa_tree_add_7_25_groupi_g15283(csa_tree_add_7_25_groupi_n_5789 ,csa_tree_add_7_25_groupi_n_5615 ,csa_tree_add_7_25_groupi_n_5701);
  xnor csa_tree_add_7_25_groupi_g15284(csa_tree_add_7_25_groupi_n_5788 ,csa_tree_add_7_25_groupi_n_5619 ,csa_tree_add_7_25_groupi_n_5702);
  xnor csa_tree_add_7_25_groupi_g15285(csa_tree_add_7_25_groupi_n_5787 ,csa_tree_add_7_25_groupi_n_5616 ,csa_tree_add_7_25_groupi_n_5683);
  xnor csa_tree_add_7_25_groupi_g15286(csa_tree_add_7_25_groupi_n_5817 ,csa_tree_add_7_25_groupi_n_5715 ,in3[17]);
  xnor csa_tree_add_7_25_groupi_g15287(csa_tree_add_7_25_groupi_n_5816 ,csa_tree_add_7_25_groupi_n_5712 ,in3[2]);
  xnor csa_tree_add_7_25_groupi_g15288(csa_tree_add_7_25_groupi_n_5815 ,csa_tree_add_7_25_groupi_n_5710 ,in3[14]);
  xnor csa_tree_add_7_25_groupi_g15289(csa_tree_add_7_25_groupi_n_5814 ,csa_tree_add_7_25_groupi_n_5713 ,in3[8]);
  xnor csa_tree_add_7_25_groupi_g15290(csa_tree_add_7_25_groupi_n_5813 ,csa_tree_add_7_25_groupi_n_5716 ,in3[5]);
  xnor csa_tree_add_7_25_groupi_g15291(csa_tree_add_7_25_groupi_n_5812 ,csa_tree_add_7_25_groupi_n_5717 ,in3[26]);
  xnor csa_tree_add_7_25_groupi_g15292(csa_tree_add_7_25_groupi_n_5811 ,csa_tree_add_7_25_groupi_n_5714 ,in3[23]);
  xnor csa_tree_add_7_25_groupi_g15293(csa_tree_add_7_25_groupi_n_5810 ,csa_tree_add_7_25_groupi_n_5709 ,in3[20]);
  xnor csa_tree_add_7_25_groupi_g15294(csa_tree_add_7_25_groupi_n_5809 ,csa_tree_add_7_25_groupi_n_5718 ,in3[11]);
  xnor csa_tree_add_7_25_groupi_g15295(csa_tree_add_7_25_groupi_n_5808 ,csa_tree_add_7_25_groupi_n_5711 ,in3[29]);
  xnor csa_tree_add_7_25_groupi_g15296(csa_tree_add_7_25_groupi_n_5807 ,csa_tree_add_7_25_groupi_n_5704 ,csa_tree_add_7_25_groupi_n_5561);
  xnor csa_tree_add_7_25_groupi_g15297(csa_tree_add_7_25_groupi_n_5806 ,csa_tree_add_7_25_groupi_n_5708 ,csa_tree_add_7_25_groupi_n_5562);
  xnor csa_tree_add_7_25_groupi_g15298(csa_tree_add_7_25_groupi_n_5805 ,csa_tree_add_7_25_groupi_n_5705 ,csa_tree_add_7_25_groupi_n_5559);
  xnor csa_tree_add_7_25_groupi_g15299(csa_tree_add_7_25_groupi_n_5804 ,csa_tree_add_7_25_groupi_n_5703 ,csa_tree_add_7_25_groupi_n_5560);
  xnor csa_tree_add_7_25_groupi_g15300(csa_tree_add_7_25_groupi_n_5803 ,csa_tree_add_7_25_groupi_n_5706 ,csa_tree_add_7_25_groupi_n_5558);
  xnor csa_tree_add_7_25_groupi_g15301(csa_tree_add_7_25_groupi_n_5802 ,csa_tree_add_7_25_groupi_n_5707 ,csa_tree_add_7_25_groupi_n_5564);
  nor csa_tree_add_7_25_groupi_g15302(csa_tree_add_7_25_groupi_n_5784 ,csa_tree_add_7_25_groupi_n_5693 ,csa_tree_add_7_25_groupi_n_5573);
  or csa_tree_add_7_25_groupi_g15303(csa_tree_add_7_25_groupi_n_5783 ,csa_tree_add_7_25_groupi_n_5625 ,csa_tree_add_7_25_groupi_n_5692);
  and csa_tree_add_7_25_groupi_g15304(csa_tree_add_7_25_groupi_n_5782 ,csa_tree_add_7_25_groupi_n_5625 ,csa_tree_add_7_25_groupi_n_5692);
  or csa_tree_add_7_25_groupi_g15305(csa_tree_add_7_25_groupi_n_5781 ,csa_tree_add_7_25_groupi_n_5698 ,csa_tree_add_7_25_groupi_n_5463);
  or csa_tree_add_7_25_groupi_g15306(csa_tree_add_7_25_groupi_n_5780 ,csa_tree_add_7_25_groupi_n_5624 ,csa_tree_add_7_25_groupi_n_5691);
  and csa_tree_add_7_25_groupi_g15307(csa_tree_add_7_25_groupi_n_5779 ,csa_tree_add_7_25_groupi_n_5624 ,csa_tree_add_7_25_groupi_n_5691);
  and csa_tree_add_7_25_groupi_g15308(csa_tree_add_7_25_groupi_n_5778 ,csa_tree_add_7_25_groupi_n_5616 ,csa_tree_add_7_25_groupi_n_5683);
  or csa_tree_add_7_25_groupi_g15309(csa_tree_add_7_25_groupi_n_5777 ,csa_tree_add_7_25_groupi_n_5616 ,csa_tree_add_7_25_groupi_n_5683);
  and csa_tree_add_7_25_groupi_g15310(csa_tree_add_7_25_groupi_n_5776 ,csa_tree_add_7_25_groupi_n_5703 ,csa_tree_add_7_25_groupi_n_5539);
  and csa_tree_add_7_25_groupi_g15311(csa_tree_add_7_25_groupi_n_5775 ,csa_tree_add_7_25_groupi_n_5707 ,csa_tree_add_7_25_groupi_n_5537);
  and csa_tree_add_7_25_groupi_g15312(csa_tree_add_7_25_groupi_n_5774 ,csa_tree_add_7_25_groupi_n_5623 ,csa_tree_add_7_25_groupi_n_5690);
  or csa_tree_add_7_25_groupi_g15313(csa_tree_add_7_25_groupi_n_5773 ,csa_tree_add_7_25_groupi_n_5623 ,csa_tree_add_7_25_groupi_n_5690);
  and csa_tree_add_7_25_groupi_g15314(csa_tree_add_7_25_groupi_n_5772 ,csa_tree_add_7_25_groupi_n_5706 ,csa_tree_add_7_25_groupi_n_5536);
  and csa_tree_add_7_25_groupi_g15315(csa_tree_add_7_25_groupi_n_5771 ,csa_tree_add_7_25_groupi_n_5619 ,csa_tree_add_7_25_groupi_n_5702);
  or csa_tree_add_7_25_groupi_g15316(csa_tree_add_7_25_groupi_n_5770 ,csa_tree_add_7_25_groupi_n_5619 ,csa_tree_add_7_25_groupi_n_5702);
  and csa_tree_add_7_25_groupi_g15317(csa_tree_add_7_25_groupi_n_5769 ,csa_tree_add_7_25_groupi_n_5705 ,csa_tree_add_7_25_groupi_n_5549);
  and csa_tree_add_7_25_groupi_g15318(csa_tree_add_7_25_groupi_n_5768 ,csa_tree_add_7_25_groupi_n_5620 ,csa_tree_add_7_25_groupi_n_5699);
  or csa_tree_add_7_25_groupi_g15319(csa_tree_add_7_25_groupi_n_5767 ,csa_tree_add_7_25_groupi_n_5620 ,csa_tree_add_7_25_groupi_n_5699);
  and csa_tree_add_7_25_groupi_g15320(csa_tree_add_7_25_groupi_n_5766 ,csa_tree_add_7_25_groupi_n_5615 ,csa_tree_add_7_25_groupi_n_5701);
  or csa_tree_add_7_25_groupi_g15321(csa_tree_add_7_25_groupi_n_5765 ,csa_tree_add_7_25_groupi_n_5615 ,csa_tree_add_7_25_groupi_n_5701);
  nor csa_tree_add_7_25_groupi_g15322(csa_tree_add_7_25_groupi_n_5764 ,csa_tree_add_7_25_groupi_n_5697 ,csa_tree_add_7_25_groupi_n_5464);
  and csa_tree_add_7_25_groupi_g15323(csa_tree_add_7_25_groupi_n_5786 ,csa_tree_add_7_25_groupi_n_2482 ,csa_tree_add_7_25_groupi_n_5728);
  or csa_tree_add_7_25_groupi_g15324(csa_tree_add_7_25_groupi_n_5785 ,csa_tree_add_7_25_groupi_n_5724 ,csa_tree_add_7_25_groupi_n_5664);
  or csa_tree_add_7_25_groupi_g15325(csa_tree_add_7_25_groupi_n_5762 ,csa_tree_add_7_25_groupi_n_5694 ,csa_tree_add_7_25_groupi_n_5572);
  nor csa_tree_add_7_25_groupi_g15326(csa_tree_add_7_25_groupi_n_5761 ,csa_tree_add_7_25_groupi_n_5617 ,csa_tree_add_7_25_groupi_n_5696);
  or csa_tree_add_7_25_groupi_g15327(csa_tree_add_7_25_groupi_n_5760 ,csa_tree_add_7_25_groupi_n_5618 ,csa_tree_add_7_25_groupi_n_5695);
  or csa_tree_add_7_25_groupi_g15328(csa_tree_add_7_25_groupi_n_5759 ,csa_tree_add_7_25_groupi_n_3298 ,csa_tree_add_7_25_groupi_n_5723);
  or csa_tree_add_7_25_groupi_g15329(csa_tree_add_7_25_groupi_n_5758 ,csa_tree_add_7_25_groupi_n_3269 ,csa_tree_add_7_25_groupi_n_5725);
  or csa_tree_add_7_25_groupi_g15330(csa_tree_add_7_25_groupi_n_5757 ,csa_tree_add_7_25_groupi_n_3264 ,csa_tree_add_7_25_groupi_n_5726);
  or csa_tree_add_7_25_groupi_g15331(csa_tree_add_7_25_groupi_n_5756 ,csa_tree_add_7_25_groupi_n_3265 ,csa_tree_add_7_25_groupi_n_5682);
  or csa_tree_add_7_25_groupi_g15332(csa_tree_add_7_25_groupi_n_5755 ,csa_tree_add_7_25_groupi_n_3683 ,csa_tree_add_7_25_groupi_n_5719);
  nor csa_tree_add_7_25_groupi_g15333(csa_tree_add_7_25_groupi_n_5754 ,csa_tree_add_7_25_groupi_n_5688 ,csa_tree_add_7_25_groupi_n_5571);
  or csa_tree_add_7_25_groupi_g15334(csa_tree_add_7_25_groupi_n_5753 ,csa_tree_add_7_25_groupi_n_5689 ,csa_tree_add_7_25_groupi_n_5570);
  nor csa_tree_add_7_25_groupi_g15335(csa_tree_add_7_25_groupi_n_5752 ,csa_tree_add_7_25_groupi_n_5626 ,csa_tree_add_7_25_groupi_n_5685);
  or csa_tree_add_7_25_groupi_g15336(csa_tree_add_7_25_groupi_n_5751 ,csa_tree_add_7_25_groupi_n_5627 ,csa_tree_add_7_25_groupi_n_5684);
  or csa_tree_add_7_25_groupi_g15337(csa_tree_add_7_25_groupi_n_5750 ,csa_tree_add_7_25_groupi_n_3682 ,csa_tree_add_7_25_groupi_n_5721);
  or csa_tree_add_7_25_groupi_g15338(csa_tree_add_7_25_groupi_n_5749 ,csa_tree_add_7_25_groupi_n_3685 ,csa_tree_add_7_25_groupi_n_5722);
  or csa_tree_add_7_25_groupi_g15339(csa_tree_add_7_25_groupi_n_5748 ,csa_tree_add_7_25_groupi_n_3686 ,csa_tree_add_7_25_groupi_n_5729);
  and csa_tree_add_7_25_groupi_g15340(csa_tree_add_7_25_groupi_n_5747 ,csa_tree_add_7_25_groupi_n_5700 ,csa_tree_add_7_25_groupi_n_5578);
  or csa_tree_add_7_25_groupi_g15341(csa_tree_add_7_25_groupi_n_5746 ,csa_tree_add_7_25_groupi_n_5700 ,csa_tree_add_7_25_groupi_n_5578);
  or csa_tree_add_7_25_groupi_g15342(csa_tree_add_7_25_groupi_n_5745 ,csa_tree_add_7_25_groupi_n_3684 ,csa_tree_add_7_25_groupi_n_5727);
  nor csa_tree_add_7_25_groupi_g15343(csa_tree_add_7_25_groupi_n_5744 ,csa_tree_add_7_25_groupi_n_5621 ,csa_tree_add_7_25_groupi_n_5687);
  or csa_tree_add_7_25_groupi_g15344(csa_tree_add_7_25_groupi_n_5743 ,csa_tree_add_7_25_groupi_n_5622 ,csa_tree_add_7_25_groupi_n_5686);
  and csa_tree_add_7_25_groupi_g15345(csa_tree_add_7_25_groupi_n_5742 ,csa_tree_add_7_25_groupi_n_5704 ,csa_tree_add_7_25_groupi_n_5515);
  and csa_tree_add_7_25_groupi_g15346(csa_tree_add_7_25_groupi_n_5741 ,csa_tree_add_7_25_groupi_n_5708 ,csa_tree_add_7_25_groupi_n_5517);
  or csa_tree_add_7_25_groupi_g15347(csa_tree_add_7_25_groupi_n_5740 ,csa_tree_add_7_25_groupi_n_3165 ,csa_tree_add_7_25_groupi_n_5720);
  xnor csa_tree_add_7_25_groupi_g15348(csa_tree_add_7_25_groupi_n_5763 ,csa_tree_add_7_25_groupi_n_5670 ,csa_tree_add_7_25_groupi_n_2570);
  nor csa_tree_add_7_25_groupi_g15349(csa_tree_add_7_25_groupi_n_5729 ,csa_tree_add_7_25_groupi_n_2063 ,csa_tree_add_7_25_groupi_n_172);
  or csa_tree_add_7_25_groupi_g15350(csa_tree_add_7_25_groupi_n_5728 ,csa_tree_add_7_25_groupi_n_2469 ,csa_tree_add_7_25_groupi_n_5670);
  nor csa_tree_add_7_25_groupi_g15351(csa_tree_add_7_25_groupi_n_5727 ,csa_tree_add_7_25_groupi_n_2154 ,csa_tree_add_7_25_groupi_n_192);
  nor csa_tree_add_7_25_groupi_g15352(csa_tree_add_7_25_groupi_n_5726 ,csa_tree_add_7_25_groupi_n_2109 ,csa_tree_add_7_25_groupi_n_1815);
  nor csa_tree_add_7_25_groupi_g15353(csa_tree_add_7_25_groupi_n_5725 ,csa_tree_add_7_25_groupi_n_2193 ,csa_tree_add_7_25_groupi_n_193);
  and csa_tree_add_7_25_groupi_g15354(csa_tree_add_7_25_groupi_n_5724 ,csa_tree_add_7_25_groupi_n_5666 ,csa_tree_add_7_25_groupi_n_5649);
  nor csa_tree_add_7_25_groupi_g15355(csa_tree_add_7_25_groupi_n_5723 ,csa_tree_add_7_25_groupi_n_2039 ,csa_tree_add_7_25_groupi_n_1854);
  nor csa_tree_add_7_25_groupi_g15356(csa_tree_add_7_25_groupi_n_5722 ,csa_tree_add_7_25_groupi_n_2027 ,csa_tree_add_7_25_groupi_n_1816);
  nor csa_tree_add_7_25_groupi_g15357(csa_tree_add_7_25_groupi_n_5721 ,csa_tree_add_7_25_groupi_n_379 ,csa_tree_add_7_25_groupi_n_193);
  nor csa_tree_add_7_25_groupi_g15358(csa_tree_add_7_25_groupi_n_5720 ,csa_tree_add_7_25_groupi_n_2181 ,csa_tree_add_7_25_groupi_n_172);
  nor csa_tree_add_7_25_groupi_g15359(csa_tree_add_7_25_groupi_n_5719 ,csa_tree_add_7_25_groupi_n_1854 ,csa_tree_add_7_25_groupi_n_1318);
  nor csa_tree_add_7_25_groupi_g15360(csa_tree_add_7_25_groupi_n_5718 ,csa_tree_add_7_25_groupi_n_3982 ,csa_tree_add_7_25_groupi_n_5637);
  nor csa_tree_add_7_25_groupi_g15361(csa_tree_add_7_25_groupi_n_5717 ,csa_tree_add_7_25_groupi_n_3829 ,csa_tree_add_7_25_groupi_n_5634);
  nor csa_tree_add_7_25_groupi_g15362(csa_tree_add_7_25_groupi_n_5716 ,csa_tree_add_7_25_groupi_n_4053 ,csa_tree_add_7_25_groupi_n_5640);
  nor csa_tree_add_7_25_groupi_g15363(csa_tree_add_7_25_groupi_n_5715 ,csa_tree_add_7_25_groupi_n_3891 ,csa_tree_add_7_25_groupi_n_5629);
  nor csa_tree_add_7_25_groupi_g15364(csa_tree_add_7_25_groupi_n_5714 ,csa_tree_add_7_25_groupi_n_3919 ,csa_tree_add_7_25_groupi_n_5633);
  nor csa_tree_add_7_25_groupi_g15365(csa_tree_add_7_25_groupi_n_5713 ,csa_tree_add_7_25_groupi_n_4061 ,csa_tree_add_7_25_groupi_n_5639);
  nor csa_tree_add_7_25_groupi_g15366(csa_tree_add_7_25_groupi_n_5712 ,csa_tree_add_7_25_groupi_n_3466 ,csa_tree_add_7_25_groupi_n_5628);
  nor csa_tree_add_7_25_groupi_g15367(csa_tree_add_7_25_groupi_n_5711 ,csa_tree_add_7_25_groupi_n_3841 ,csa_tree_add_7_25_groupi_n_5647);
  nor csa_tree_add_7_25_groupi_g15368(csa_tree_add_7_25_groupi_n_5710 ,csa_tree_add_7_25_groupi_n_4017 ,csa_tree_add_7_25_groupi_n_5638);
  nor csa_tree_add_7_25_groupi_g15369(csa_tree_add_7_25_groupi_n_5709 ,csa_tree_add_7_25_groupi_n_3874 ,csa_tree_add_7_25_groupi_n_5632);
  or csa_tree_add_7_25_groupi_g15370(csa_tree_add_7_25_groupi_n_5739 ,csa_tree_add_7_25_groupi_n_5419 ,csa_tree_add_7_25_groupi_n_5635);
  or csa_tree_add_7_25_groupi_g15371(csa_tree_add_7_25_groupi_n_5738 ,csa_tree_add_7_25_groupi_n_5169 ,csa_tree_add_7_25_groupi_n_5643);
  or csa_tree_add_7_25_groupi_g15372(csa_tree_add_7_25_groupi_n_5737 ,csa_tree_add_7_25_groupi_n_5438 ,csa_tree_add_7_25_groupi_n_5665);
  or csa_tree_add_7_25_groupi_g15373(csa_tree_add_7_25_groupi_n_5736 ,csa_tree_add_7_25_groupi_n_5405 ,csa_tree_add_7_25_groupi_n_5656);
  or csa_tree_add_7_25_groupi_g15374(csa_tree_add_7_25_groupi_n_5735 ,csa_tree_add_7_25_groupi_n_5431 ,csa_tree_add_7_25_groupi_n_5654);
  or csa_tree_add_7_25_groupi_g15375(csa_tree_add_7_25_groupi_n_5734 ,csa_tree_add_7_25_groupi_n_5433 ,csa_tree_add_7_25_groupi_n_5657);
  or csa_tree_add_7_25_groupi_g15376(csa_tree_add_7_25_groupi_n_5733 ,csa_tree_add_7_25_groupi_n_5435 ,csa_tree_add_7_25_groupi_n_5658);
  or csa_tree_add_7_25_groupi_g15377(csa_tree_add_7_25_groupi_n_5732 ,csa_tree_add_7_25_groupi_n_5437 ,csa_tree_add_7_25_groupi_n_5662);
  or csa_tree_add_7_25_groupi_g15378(csa_tree_add_7_25_groupi_n_5731 ,csa_tree_add_7_25_groupi_n_5429 ,csa_tree_add_7_25_groupi_n_5652);
  or csa_tree_add_7_25_groupi_g15379(csa_tree_add_7_25_groupi_n_5730 ,csa_tree_add_7_25_groupi_n_5427 ,csa_tree_add_7_25_groupi_n_5646);
  not csa_tree_add_7_25_groupi_g15380(csa_tree_add_7_25_groupi_n_5697 ,csa_tree_add_7_25_groupi_n_5698);
  not csa_tree_add_7_25_groupi_g15381(csa_tree_add_7_25_groupi_n_5695 ,csa_tree_add_7_25_groupi_n_5696);
  not csa_tree_add_7_25_groupi_g15382(csa_tree_add_7_25_groupi_n_5693 ,csa_tree_add_7_25_groupi_n_5694);
  not csa_tree_add_7_25_groupi_g15383(csa_tree_add_7_25_groupi_n_5688 ,csa_tree_add_7_25_groupi_n_5689);
  not csa_tree_add_7_25_groupi_g15384(csa_tree_add_7_25_groupi_n_5686 ,csa_tree_add_7_25_groupi_n_5687);
  not csa_tree_add_7_25_groupi_g15385(csa_tree_add_7_25_groupi_n_5684 ,csa_tree_add_7_25_groupi_n_5685);
  nor csa_tree_add_7_25_groupi_g15386(csa_tree_add_7_25_groupi_n_5682 ,csa_tree_add_7_25_groupi_n_2163 ,csa_tree_add_7_25_groupi_n_1815);
  xnor csa_tree_add_7_25_groupi_g15387(out2[8] ,csa_tree_add_7_25_groupi_n_5555 ,csa_tree_add_7_25_groupi_n_5563);
  xnor csa_tree_add_7_25_groupi_g15388(csa_tree_add_7_25_groupi_n_5680 ,csa_tree_add_7_25_groupi_n_5534 ,csa_tree_add_7_25_groupi_n_5576);
  xnor csa_tree_add_7_25_groupi_g15389(csa_tree_add_7_25_groupi_n_5679 ,csa_tree_add_7_25_groupi_n_5582 ,csa_tree_add_7_25_groupi_n_5513);
  xnor csa_tree_add_7_25_groupi_g15390(csa_tree_add_7_25_groupi_n_5678 ,csa_tree_add_7_25_groupi_n_5580 ,csa_tree_add_7_25_groupi_n_5511);
  xnor csa_tree_add_7_25_groupi_g15391(csa_tree_add_7_25_groupi_n_5677 ,csa_tree_add_7_25_groupi_n_5577 ,csa_tree_add_7_25_groupi_n_5512);
  xnor csa_tree_add_7_25_groupi_g15392(csa_tree_add_7_25_groupi_n_5676 ,csa_tree_add_7_25_groupi_n_5581 ,csa_tree_add_7_25_groupi_n_5510);
  xnor csa_tree_add_7_25_groupi_g15393(csa_tree_add_7_25_groupi_n_5675 ,csa_tree_add_7_25_groupi_n_5575 ,csa_tree_add_7_25_groupi_n_5509);
  xnor csa_tree_add_7_25_groupi_g15394(csa_tree_add_7_25_groupi_n_5674 ,csa_tree_add_7_25_groupi_n_5579 ,csa_tree_add_7_25_groupi_n_5508);
  xnor csa_tree_add_7_25_groupi_g15395(csa_tree_add_7_25_groupi_n_5673 ,csa_tree_add_7_25_groupi_n_5554 ,csa_tree_add_7_25_groupi_n_5567);
  xnor csa_tree_add_7_25_groupi_g15396(csa_tree_add_7_25_groupi_n_5672 ,csa_tree_add_7_25_groupi_n_5569 ,csa_tree_add_7_25_groupi_n_5552);
  xnor csa_tree_add_7_25_groupi_g15397(csa_tree_add_7_25_groupi_n_5671 ,csa_tree_add_7_25_groupi_n_5574 ,csa_tree_add_7_25_groupi_n_5514);
  xnor csa_tree_add_7_25_groupi_g15398(csa_tree_add_7_25_groupi_n_5708 ,csa_tree_add_7_25_groupi_n_5593 ,in3[5]);
  xnor csa_tree_add_7_25_groupi_g15399(csa_tree_add_7_25_groupi_n_5707 ,csa_tree_add_7_25_groupi_n_5597 ,in3[8]);
  xnor csa_tree_add_7_25_groupi_g15400(csa_tree_add_7_25_groupi_n_5706 ,csa_tree_add_7_25_groupi_n_5601 ,in3[11]);
  xnor csa_tree_add_7_25_groupi_g15401(csa_tree_add_7_25_groupi_n_5705 ,csa_tree_add_7_25_groupi_n_5598 ,in3[14]);
  xnor csa_tree_add_7_25_groupi_g15402(csa_tree_add_7_25_groupi_n_5704 ,csa_tree_add_7_25_groupi_n_5594 ,in3[2]);
  xnor csa_tree_add_7_25_groupi_g15403(csa_tree_add_7_25_groupi_n_5703 ,csa_tree_add_7_25_groupi_n_5595 ,in3[17]);
  xnor csa_tree_add_7_25_groupi_g15404(csa_tree_add_7_25_groupi_n_5702 ,csa_tree_add_7_25_groupi_n_5587 ,csa_tree_add_7_25_groupi_n_5454);
  xnor csa_tree_add_7_25_groupi_g15405(csa_tree_add_7_25_groupi_n_5701 ,csa_tree_add_7_25_groupi_n_5585 ,csa_tree_add_7_25_groupi_n_5453);
  xnor csa_tree_add_7_25_groupi_g15406(csa_tree_add_7_25_groupi_n_5700 ,csa_tree_add_7_25_groupi_n_5600 ,in3[20]);
  xnor csa_tree_add_7_25_groupi_g15407(csa_tree_add_7_25_groupi_n_5699 ,csa_tree_add_7_25_groupi_n_5584 ,csa_tree_add_7_25_groupi_n_5452);
  xnor csa_tree_add_7_25_groupi_g15408(csa_tree_add_7_25_groupi_n_5698 ,csa_tree_add_7_25_groupi_n_5599 ,in3[29]);
  xnor csa_tree_add_7_25_groupi_g15409(csa_tree_add_7_25_groupi_n_5696 ,csa_tree_add_7_25_groupi_n_5592 ,csa_tree_add_7_25_groupi_n_5457);
  xnor csa_tree_add_7_25_groupi_g15410(csa_tree_add_7_25_groupi_n_5694 ,csa_tree_add_7_25_groupi_n_5602 ,in3[26]);
  xnor csa_tree_add_7_25_groupi_g15411(csa_tree_add_7_25_groupi_n_5692 ,csa_tree_add_7_25_groupi_n_5586 ,csa_tree_add_7_25_groupi_n_5449);
  xnor csa_tree_add_7_25_groupi_g15412(csa_tree_add_7_25_groupi_n_5691 ,csa_tree_add_7_25_groupi_n_5589 ,csa_tree_add_7_25_groupi_n_5450);
  xnor csa_tree_add_7_25_groupi_g15413(csa_tree_add_7_25_groupi_n_5690 ,csa_tree_add_7_25_groupi_n_5583 ,csa_tree_add_7_25_groupi_n_5451);
  xnor csa_tree_add_7_25_groupi_g15414(csa_tree_add_7_25_groupi_n_5689 ,csa_tree_add_7_25_groupi_n_5596 ,in3[23]);
  xnor csa_tree_add_7_25_groupi_g15415(csa_tree_add_7_25_groupi_n_5687 ,csa_tree_add_7_25_groupi_n_5590 ,csa_tree_add_7_25_groupi_n_5218);
  xnor csa_tree_add_7_25_groupi_g15416(csa_tree_add_7_25_groupi_n_5685 ,csa_tree_add_7_25_groupi_n_5591 ,csa_tree_add_7_25_groupi_n_5461);
  xnor csa_tree_add_7_25_groupi_g15417(csa_tree_add_7_25_groupi_n_5683 ,csa_tree_add_7_25_groupi_n_5588 ,csa_tree_add_7_25_groupi_n_5458);
  and csa_tree_add_7_25_groupi_g15418(csa_tree_add_7_25_groupi_n_5669 ,csa_tree_add_7_25_groupi_n_5574 ,csa_tree_add_7_25_groupi_n_5514);
  and csa_tree_add_7_25_groupi_g15419(csa_tree_add_7_25_groupi_n_5668 ,csa_tree_add_7_25_groupi_n_5534 ,csa_tree_add_7_25_groupi_n_5576);
  or csa_tree_add_7_25_groupi_g15420(csa_tree_add_7_25_groupi_n_5667 ,csa_tree_add_7_25_groupi_n_5534 ,csa_tree_add_7_25_groupi_n_5576);
  or csa_tree_add_7_25_groupi_g15421(csa_tree_add_7_25_groupi_n_5666 ,csa_tree_add_7_25_groupi_n_5582 ,csa_tree_add_7_25_groupi_n_5513);
  and csa_tree_add_7_25_groupi_g15422(csa_tree_add_7_25_groupi_n_5665 ,csa_tree_add_7_25_groupi_n_5588 ,csa_tree_add_7_25_groupi_n_5445);
  and csa_tree_add_7_25_groupi_g15423(csa_tree_add_7_25_groupi_n_5664 ,csa_tree_add_7_25_groupi_n_5582 ,csa_tree_add_7_25_groupi_n_5513);
  and csa_tree_add_7_25_groupi_g15424(csa_tree_add_7_25_groupi_n_5663 ,csa_tree_add_7_25_groupi_n_5580 ,csa_tree_add_7_25_groupi_n_5511);
  and csa_tree_add_7_25_groupi_g15425(csa_tree_add_7_25_groupi_n_5662 ,csa_tree_add_7_25_groupi_n_5586 ,csa_tree_add_7_25_groupi_n_5436);
  or csa_tree_add_7_25_groupi_g15426(csa_tree_add_7_25_groupi_n_5661 ,csa_tree_add_7_25_groupi_n_5580 ,csa_tree_add_7_25_groupi_n_5511);
  and csa_tree_add_7_25_groupi_g15427(csa_tree_add_7_25_groupi_n_5660 ,csa_tree_add_7_25_groupi_n_5577 ,csa_tree_add_7_25_groupi_n_5512);
  or csa_tree_add_7_25_groupi_g15428(csa_tree_add_7_25_groupi_n_5659 ,csa_tree_add_7_25_groupi_n_5577 ,csa_tree_add_7_25_groupi_n_5512);
  and csa_tree_add_7_25_groupi_g15429(csa_tree_add_7_25_groupi_n_5658 ,csa_tree_add_7_25_groupi_n_5589 ,csa_tree_add_7_25_groupi_n_5434);
  and csa_tree_add_7_25_groupi_g15430(csa_tree_add_7_25_groupi_n_5657 ,csa_tree_add_7_25_groupi_n_5587 ,csa_tree_add_7_25_groupi_n_5432);
  and csa_tree_add_7_25_groupi_g15431(csa_tree_add_7_25_groupi_n_5656 ,csa_tree_add_7_25_groupi_n_5592 ,csa_tree_add_7_25_groupi_n_5404);
  and csa_tree_add_7_25_groupi_g15432(csa_tree_add_7_25_groupi_n_5655 ,csa_tree_add_7_25_groupi_n_5581 ,csa_tree_add_7_25_groupi_n_5510);
  and csa_tree_add_7_25_groupi_g15433(csa_tree_add_7_25_groupi_n_5654 ,csa_tree_add_7_25_groupi_n_5583 ,csa_tree_add_7_25_groupi_n_5430);
  or csa_tree_add_7_25_groupi_g15434(csa_tree_add_7_25_groupi_n_5653 ,csa_tree_add_7_25_groupi_n_5581 ,csa_tree_add_7_25_groupi_n_5510);
  and csa_tree_add_7_25_groupi_g15435(csa_tree_add_7_25_groupi_n_5652 ,csa_tree_add_7_25_groupi_n_5584 ,csa_tree_add_7_25_groupi_n_5428);
  and csa_tree_add_7_25_groupi_g15436(csa_tree_add_7_25_groupi_n_5651 ,csa_tree_add_7_25_groupi_n_5575 ,csa_tree_add_7_25_groupi_n_5509);
  or csa_tree_add_7_25_groupi_g15437(csa_tree_add_7_25_groupi_n_5650 ,csa_tree_add_7_25_groupi_n_5575 ,csa_tree_add_7_25_groupi_n_5509);
  and csa_tree_add_7_25_groupi_g15438(csa_tree_add_7_25_groupi_n_5670 ,csa_tree_add_7_25_groupi_n_2466 ,csa_tree_add_7_25_groupi_n_5609);
  or csa_tree_add_7_25_groupi_g15439(csa_tree_add_7_25_groupi_n_5647 ,csa_tree_add_7_25_groupi_n_3671 ,csa_tree_add_7_25_groupi_n_5603);
  and csa_tree_add_7_25_groupi_g15440(csa_tree_add_7_25_groupi_n_5646 ,csa_tree_add_7_25_groupi_n_5585 ,csa_tree_add_7_25_groupi_n_5426);
  nor csa_tree_add_7_25_groupi_g15441(csa_tree_add_7_25_groupi_n_5645 ,csa_tree_add_7_25_groupi_n_5569 ,csa_tree_add_7_25_groupi_n_5551);
  or csa_tree_add_7_25_groupi_g15442(csa_tree_add_7_25_groupi_n_5644 ,csa_tree_add_7_25_groupi_n_5568 ,csa_tree_add_7_25_groupi_n_5552);
  and csa_tree_add_7_25_groupi_g15443(csa_tree_add_7_25_groupi_n_5643 ,csa_tree_add_7_25_groupi_n_5168 ,csa_tree_add_7_25_groupi_n_5590);
  nor csa_tree_add_7_25_groupi_g15444(csa_tree_add_7_25_groupi_n_5642 ,csa_tree_add_7_25_groupi_n_5553 ,csa_tree_add_7_25_groupi_n_5567);
  or csa_tree_add_7_25_groupi_g15445(csa_tree_add_7_25_groupi_n_5641 ,csa_tree_add_7_25_groupi_n_5554 ,csa_tree_add_7_25_groupi_n_5566);
  or csa_tree_add_7_25_groupi_g15446(csa_tree_add_7_25_groupi_n_5640 ,csa_tree_add_7_25_groupi_n_3251 ,csa_tree_add_7_25_groupi_n_5610);
  or csa_tree_add_7_25_groupi_g15447(csa_tree_add_7_25_groupi_n_5639 ,csa_tree_add_7_25_groupi_n_3248 ,csa_tree_add_7_25_groupi_n_5611);
  or csa_tree_add_7_25_groupi_g15448(csa_tree_add_7_25_groupi_n_5638 ,csa_tree_add_7_25_groupi_n_3247 ,csa_tree_add_7_25_groupi_n_5612);
  or csa_tree_add_7_25_groupi_g15449(csa_tree_add_7_25_groupi_n_5637 ,csa_tree_add_7_25_groupi_n_3249 ,csa_tree_add_7_25_groupi_n_5613);
  or csa_tree_add_7_25_groupi_g15450(csa_tree_add_7_25_groupi_n_5636 ,csa_tree_add_7_25_groupi_n_5574 ,csa_tree_add_7_25_groupi_n_5514);
  and csa_tree_add_7_25_groupi_g15451(csa_tree_add_7_25_groupi_n_5635 ,csa_tree_add_7_25_groupi_n_5591 ,csa_tree_add_7_25_groupi_n_5418);
  or csa_tree_add_7_25_groupi_g15452(csa_tree_add_7_25_groupi_n_5634 ,csa_tree_add_7_25_groupi_n_3672 ,csa_tree_add_7_25_groupi_n_5605);
  or csa_tree_add_7_25_groupi_g15453(csa_tree_add_7_25_groupi_n_5633 ,csa_tree_add_7_25_groupi_n_3680 ,csa_tree_add_7_25_groupi_n_5606);
  or csa_tree_add_7_25_groupi_g15454(csa_tree_add_7_25_groupi_n_5632 ,csa_tree_add_7_25_groupi_n_3670 ,csa_tree_add_7_25_groupi_n_5607);
  and csa_tree_add_7_25_groupi_g15455(csa_tree_add_7_25_groupi_n_5631 ,csa_tree_add_7_25_groupi_n_5579 ,csa_tree_add_7_25_groupi_n_5508);
  or csa_tree_add_7_25_groupi_g15456(csa_tree_add_7_25_groupi_n_5630 ,csa_tree_add_7_25_groupi_n_5579 ,csa_tree_add_7_25_groupi_n_5508);
  or csa_tree_add_7_25_groupi_g15457(csa_tree_add_7_25_groupi_n_5629 ,csa_tree_add_7_25_groupi_n_3668 ,csa_tree_add_7_25_groupi_n_5608);
  or csa_tree_add_7_25_groupi_g15458(csa_tree_add_7_25_groupi_n_5628 ,csa_tree_add_7_25_groupi_n_3093 ,csa_tree_add_7_25_groupi_n_5604);
  or csa_tree_add_7_25_groupi_g15459(csa_tree_add_7_25_groupi_n_5649 ,csa_tree_add_7_25_groupi_n_5614 ,csa_tree_add_7_25_groupi_n_5519);
  xnor csa_tree_add_7_25_groupi_g15460(csa_tree_add_7_25_groupi_n_5648 ,csa_tree_add_7_25_groupi_n_5556 ,csa_tree_add_7_25_groupi_n_2571);
  not csa_tree_add_7_25_groupi_g15461(csa_tree_add_7_25_groupi_n_5626 ,csa_tree_add_7_25_groupi_n_5627);
  not csa_tree_add_7_25_groupi_g15462(csa_tree_add_7_25_groupi_n_5621 ,csa_tree_add_7_25_groupi_n_5622);
  not csa_tree_add_7_25_groupi_g15463(csa_tree_add_7_25_groupi_n_5617 ,csa_tree_add_7_25_groupi_n_5618);
  and csa_tree_add_7_25_groupi_g15464(csa_tree_add_7_25_groupi_n_5614 ,csa_tree_add_7_25_groupi_n_5555 ,csa_tree_add_7_25_groupi_n_5520);
  nor csa_tree_add_7_25_groupi_g15465(csa_tree_add_7_25_groupi_n_5613 ,csa_tree_add_7_25_groupi_n_2099 ,csa_tree_add_7_25_groupi_n_1870);
  nor csa_tree_add_7_25_groupi_g15466(csa_tree_add_7_25_groupi_n_5612 ,csa_tree_add_7_25_groupi_n_2150 ,csa_tree_add_7_25_groupi_n_179);
  nor csa_tree_add_7_25_groupi_g15467(csa_tree_add_7_25_groupi_n_5611 ,csa_tree_add_7_25_groupi_n_2120 ,csa_tree_add_7_25_groupi_n_209);
  nor csa_tree_add_7_25_groupi_g15468(csa_tree_add_7_25_groupi_n_5610 ,csa_tree_add_7_25_groupi_n_2135 ,csa_tree_add_7_25_groupi_n_1812);
  or csa_tree_add_7_25_groupi_g15469(csa_tree_add_7_25_groupi_n_5609 ,csa_tree_add_7_25_groupi_n_2457 ,csa_tree_add_7_25_groupi_n_5556);
  nor csa_tree_add_7_25_groupi_g15470(csa_tree_add_7_25_groupi_n_5608 ,csa_tree_add_7_25_groupi_n_2061 ,csa_tree_add_7_25_groupi_n_179);
  nor csa_tree_add_7_25_groupi_g15471(csa_tree_add_7_25_groupi_n_5607 ,csa_tree_add_7_25_groupi_n_2048 ,csa_tree_add_7_25_groupi_n_208);
  nor csa_tree_add_7_25_groupi_g15472(csa_tree_add_7_25_groupi_n_5606 ,csa_tree_add_7_25_groupi_n_2027 ,csa_tree_add_7_25_groupi_n_1813);
  nor csa_tree_add_7_25_groupi_g15473(csa_tree_add_7_25_groupi_n_5605 ,csa_tree_add_7_25_groupi_n_209 ,csa_tree_add_7_25_groupi_n_1310);
  nor csa_tree_add_7_25_groupi_g15474(csa_tree_add_7_25_groupi_n_5604 ,csa_tree_add_7_25_groupi_n_2177 ,csa_tree_add_7_25_groupi_n_1812);
  nor csa_tree_add_7_25_groupi_g15475(csa_tree_add_7_25_groupi_n_5603 ,csa_tree_add_7_25_groupi_n_1870 ,csa_tree_add_7_25_groupi_n_1322);
  nor csa_tree_add_7_25_groupi_g15476(csa_tree_add_7_25_groupi_n_5602 ,csa_tree_add_7_25_groupi_n_3906 ,csa_tree_add_7_25_groupi_n_5523);
  nor csa_tree_add_7_25_groupi_g15477(csa_tree_add_7_25_groupi_n_5601 ,csa_tree_add_7_25_groupi_n_4098 ,csa_tree_add_7_25_groupi_n_5527);
  nor csa_tree_add_7_25_groupi_g15478(csa_tree_add_7_25_groupi_n_5600 ,csa_tree_add_7_25_groupi_n_3888 ,csa_tree_add_7_25_groupi_n_5522);
  nor csa_tree_add_7_25_groupi_g15479(csa_tree_add_7_25_groupi_n_5599 ,csa_tree_add_7_25_groupi_n_3901 ,csa_tree_add_7_25_groupi_n_5524);
  nor csa_tree_add_7_25_groupi_g15480(csa_tree_add_7_25_groupi_n_5598 ,csa_tree_add_7_25_groupi_n_3981 ,csa_tree_add_7_25_groupi_n_5525);
  nor csa_tree_add_7_25_groupi_g15481(csa_tree_add_7_25_groupi_n_5597 ,csa_tree_add_7_25_groupi_n_4065 ,csa_tree_add_7_25_groupi_n_5526);
  nor csa_tree_add_7_25_groupi_g15482(csa_tree_add_7_25_groupi_n_5596 ,csa_tree_add_7_25_groupi_n_4076 ,csa_tree_add_7_25_groupi_n_5531);
  nor csa_tree_add_7_25_groupi_g15483(csa_tree_add_7_25_groupi_n_5595 ,csa_tree_add_7_25_groupi_n_3853 ,csa_tree_add_7_25_groupi_n_5521);
  nor csa_tree_add_7_25_groupi_g15484(csa_tree_add_7_25_groupi_n_5594 ,csa_tree_add_7_25_groupi_n_3485 ,csa_tree_add_7_25_groupi_n_5528);
  nor csa_tree_add_7_25_groupi_g15485(csa_tree_add_7_25_groupi_n_5593 ,csa_tree_add_7_25_groupi_n_4013 ,csa_tree_add_7_25_groupi_n_5530);
  or csa_tree_add_7_25_groupi_g15486(csa_tree_add_7_25_groupi_n_5627 ,csa_tree_add_7_25_groupi_n_5321 ,csa_tree_add_7_25_groupi_n_5547);
  or csa_tree_add_7_25_groupi_g15487(csa_tree_add_7_25_groupi_n_5625 ,csa_tree_add_7_25_groupi_n_5317 ,csa_tree_add_7_25_groupi_n_5546);
  or csa_tree_add_7_25_groupi_g15488(csa_tree_add_7_25_groupi_n_5624 ,csa_tree_add_7_25_groupi_n_5313 ,csa_tree_add_7_25_groupi_n_5545);
  or csa_tree_add_7_25_groupi_g15489(csa_tree_add_7_25_groupi_n_5623 ,csa_tree_add_7_25_groupi_n_5311 ,csa_tree_add_7_25_groupi_n_5544);
  or csa_tree_add_7_25_groupi_g15490(csa_tree_add_7_25_groupi_n_5622 ,csa_tree_add_7_25_groupi_n_5099 ,csa_tree_add_7_25_groupi_n_5550);
  or csa_tree_add_7_25_groupi_g15491(csa_tree_add_7_25_groupi_n_5620 ,csa_tree_add_7_25_groupi_n_5305 ,csa_tree_add_7_25_groupi_n_5542);
  or csa_tree_add_7_25_groupi_g15492(csa_tree_add_7_25_groupi_n_5619 ,csa_tree_add_7_25_groupi_n_5291 ,csa_tree_add_7_25_groupi_n_5541);
  or csa_tree_add_7_25_groupi_g15493(csa_tree_add_7_25_groupi_n_5618 ,csa_tree_add_7_25_groupi_n_5298 ,csa_tree_add_7_25_groupi_n_5532);
  or csa_tree_add_7_25_groupi_g15494(csa_tree_add_7_25_groupi_n_5616 ,csa_tree_add_7_25_groupi_n_5295 ,csa_tree_add_7_25_groupi_n_5529);
  or csa_tree_add_7_25_groupi_g15495(csa_tree_add_7_25_groupi_n_5615 ,csa_tree_add_7_25_groupi_n_5308 ,csa_tree_add_7_25_groupi_n_5543);
  not csa_tree_add_7_25_groupi_g15496(csa_tree_add_7_25_groupi_n_5572 ,csa_tree_add_7_25_groupi_n_5573);
  not csa_tree_add_7_25_groupi_g15497(csa_tree_add_7_25_groupi_n_5570 ,csa_tree_add_7_25_groupi_n_5571);
  not csa_tree_add_7_25_groupi_g15498(csa_tree_add_7_25_groupi_n_5568 ,csa_tree_add_7_25_groupi_n_5569);
  not csa_tree_add_7_25_groupi_g15499(csa_tree_add_7_25_groupi_n_5566 ,csa_tree_add_7_25_groupi_n_5567);
  xnor csa_tree_add_7_25_groupi_g15500(out2[7] ,csa_tree_add_7_25_groupi_n_5446 ,csa_tree_add_7_25_groupi_n_5448);
  xnor csa_tree_add_7_25_groupi_g15501(csa_tree_add_7_25_groupi_n_5564 ,csa_tree_add_7_25_groupi_n_5471 ,csa_tree_add_7_25_groupi_n_5391);
  xnor csa_tree_add_7_25_groupi_g15502(csa_tree_add_7_25_groupi_n_5563 ,csa_tree_add_7_25_groupi_n_5465 ,csa_tree_add_7_25_groupi_n_5395);
  xnor csa_tree_add_7_25_groupi_g15503(csa_tree_add_7_25_groupi_n_5562 ,csa_tree_add_7_25_groupi_n_5466 ,csa_tree_add_7_25_groupi_n_5393);
  xnor csa_tree_add_7_25_groupi_g15504(csa_tree_add_7_25_groupi_n_5561 ,csa_tree_add_7_25_groupi_n_5467 ,csa_tree_add_7_25_groupi_n_5394);
  xnor csa_tree_add_7_25_groupi_g15505(csa_tree_add_7_25_groupi_n_5560 ,csa_tree_add_7_25_groupi_n_5389 ,csa_tree_add_7_25_groupi_n_5470);
  xnor csa_tree_add_7_25_groupi_g15506(csa_tree_add_7_25_groupi_n_5559 ,csa_tree_add_7_25_groupi_n_5469 ,csa_tree_add_7_25_groupi_n_5390);
  xnor csa_tree_add_7_25_groupi_g15507(csa_tree_add_7_25_groupi_n_5558 ,csa_tree_add_7_25_groupi_n_5468 ,csa_tree_add_7_25_groupi_n_5392);
  xnor csa_tree_add_7_25_groupi_g15508(csa_tree_add_7_25_groupi_n_5557 ,csa_tree_add_7_25_groupi_n_5482 ,csa_tree_add_7_25_groupi_n_1973);
  xnor csa_tree_add_7_25_groupi_g15509(csa_tree_add_7_25_groupi_n_5592 ,csa_tree_add_7_25_groupi_n_5492 ,in3[26]);
  xnor csa_tree_add_7_25_groupi_g15510(csa_tree_add_7_25_groupi_n_5591 ,csa_tree_add_7_25_groupi_n_5488 ,in3[23]);
  xnor csa_tree_add_7_25_groupi_g15511(csa_tree_add_7_25_groupi_n_5590 ,csa_tree_add_7_25_groupi_n_5487 ,in3[29]);
  xnor csa_tree_add_7_25_groupi_g15512(csa_tree_add_7_25_groupi_n_5589 ,csa_tree_add_7_25_groupi_n_5491 ,in3[5]);
  xnor csa_tree_add_7_25_groupi_g15513(csa_tree_add_7_25_groupi_n_5588 ,csa_tree_add_7_25_groupi_n_5489 ,in3[20]);
  xnor csa_tree_add_7_25_groupi_g15514(csa_tree_add_7_25_groupi_n_5587 ,csa_tree_add_7_25_groupi_n_5490 ,in3[17]);
  xnor csa_tree_add_7_25_groupi_g15515(csa_tree_add_7_25_groupi_n_5586 ,csa_tree_add_7_25_groupi_n_5486 ,in3[2]);
  xnor csa_tree_add_7_25_groupi_g15516(csa_tree_add_7_25_groupi_n_5585 ,csa_tree_add_7_25_groupi_n_5485 ,in3[14]);
  xnor csa_tree_add_7_25_groupi_g15517(csa_tree_add_7_25_groupi_n_5584 ,csa_tree_add_7_25_groupi_n_5483 ,in3[11]);
  xnor csa_tree_add_7_25_groupi_g15518(csa_tree_add_7_25_groupi_n_5583 ,csa_tree_add_7_25_groupi_n_5484 ,in3[8]);
  xnor csa_tree_add_7_25_groupi_g15519(csa_tree_add_7_25_groupi_n_5582 ,csa_tree_add_7_25_groupi_n_5480 ,csa_tree_add_7_25_groupi_n_5333);
  xnor csa_tree_add_7_25_groupi_g15520(csa_tree_add_7_25_groupi_n_5581 ,csa_tree_add_7_25_groupi_n_5478 ,csa_tree_add_7_25_groupi_n_5330);
  xnor csa_tree_add_7_25_groupi_g15521(csa_tree_add_7_25_groupi_n_5580 ,csa_tree_add_7_25_groupi_n_5476 ,csa_tree_add_7_25_groupi_n_5332);
  xnor csa_tree_add_7_25_groupi_g15522(csa_tree_add_7_25_groupi_n_5579 ,csa_tree_add_7_25_groupi_n_5475 ,csa_tree_add_7_25_groupi_n_5329);
  xnor csa_tree_add_7_25_groupi_g15523(csa_tree_add_7_25_groupi_n_5578 ,csa_tree_add_7_25_groupi_n_5396 ,csa_tree_add_7_25_groupi_n_5456);
  xnor csa_tree_add_7_25_groupi_g15524(csa_tree_add_7_25_groupi_n_5577 ,csa_tree_add_7_25_groupi_n_5477 ,csa_tree_add_7_25_groupi_n_5331);
  xnor csa_tree_add_7_25_groupi_g15525(csa_tree_add_7_25_groupi_n_5576 ,csa_tree_add_7_25_groupi_n_5473 ,csa_tree_add_7_25_groupi_n_5335);
  xnor csa_tree_add_7_25_groupi_g15526(csa_tree_add_7_25_groupi_n_5575 ,csa_tree_add_7_25_groupi_n_5479 ,csa_tree_add_7_25_groupi_n_5328);
  xnor csa_tree_add_7_25_groupi_g15527(csa_tree_add_7_25_groupi_n_5574 ,csa_tree_add_7_25_groupi_n_5481 ,csa_tree_add_7_25_groupi_n_5327);
  xnor csa_tree_add_7_25_groupi_g15528(csa_tree_add_7_25_groupi_n_5573 ,csa_tree_add_7_25_groupi_n_5397 ,csa_tree_add_7_25_groupi_n_5460);
  xnor csa_tree_add_7_25_groupi_g15529(csa_tree_add_7_25_groupi_n_5571 ,csa_tree_add_7_25_groupi_n_5398 ,csa_tree_add_7_25_groupi_n_5459);
  xnor csa_tree_add_7_25_groupi_g15530(csa_tree_add_7_25_groupi_n_5569 ,csa_tree_add_7_25_groupi_n_5472 ,csa_tree_add_7_25_groupi_n_1);
  xnor csa_tree_add_7_25_groupi_g15531(csa_tree_add_7_25_groupi_n_5567 ,csa_tree_add_7_25_groupi_n_5474 ,csa_tree_add_7_25_groupi_n_5336);
  not csa_tree_add_7_25_groupi_g15532(csa_tree_add_7_25_groupi_n_5553 ,csa_tree_add_7_25_groupi_n_5554);
  not csa_tree_add_7_25_groupi_g15533(csa_tree_add_7_25_groupi_n_5551 ,csa_tree_add_7_25_groupi_n_5552);
  and csa_tree_add_7_25_groupi_g15534(csa_tree_add_7_25_groupi_n_5550 ,csa_tree_add_7_25_groupi_n_5472 ,csa_tree_add_7_25_groupi_n_5104);
  or csa_tree_add_7_25_groupi_g15535(csa_tree_add_7_25_groupi_n_5549 ,csa_tree_add_7_25_groupi_n_5469 ,csa_tree_add_7_25_groupi_n_5390);
  and csa_tree_add_7_25_groupi_g15536(csa_tree_add_7_25_groupi_n_5548 ,csa_tree_add_7_25_groupi_n_5469 ,csa_tree_add_7_25_groupi_n_5390);
  and csa_tree_add_7_25_groupi_g15537(csa_tree_add_7_25_groupi_n_5547 ,csa_tree_add_7_25_groupi_n_5473 ,csa_tree_add_7_25_groupi_n_5319);
  and csa_tree_add_7_25_groupi_g15538(csa_tree_add_7_25_groupi_n_5546 ,csa_tree_add_7_25_groupi_n_5480 ,csa_tree_add_7_25_groupi_n_5316);
  and csa_tree_add_7_25_groupi_g15539(csa_tree_add_7_25_groupi_n_5545 ,csa_tree_add_7_25_groupi_n_5476 ,csa_tree_add_7_25_groupi_n_5312);
  and csa_tree_add_7_25_groupi_g15540(csa_tree_add_7_25_groupi_n_5544 ,csa_tree_add_7_25_groupi_n_5477 ,csa_tree_add_7_25_groupi_n_5310);
  and csa_tree_add_7_25_groupi_g15541(csa_tree_add_7_25_groupi_n_5543 ,csa_tree_add_7_25_groupi_n_5479 ,csa_tree_add_7_25_groupi_n_5307);
  and csa_tree_add_7_25_groupi_g15542(csa_tree_add_7_25_groupi_n_5542 ,csa_tree_add_7_25_groupi_n_5478 ,csa_tree_add_7_25_groupi_n_5284);
  and csa_tree_add_7_25_groupi_g15543(csa_tree_add_7_25_groupi_n_5541 ,csa_tree_add_7_25_groupi_n_5481 ,csa_tree_add_7_25_groupi_n_5301);
  and csa_tree_add_7_25_groupi_g15544(csa_tree_add_7_25_groupi_n_5540 ,csa_tree_add_7_25_groupi_n_5389 ,csa_tree_add_7_25_groupi_n_5470);
  or csa_tree_add_7_25_groupi_g15545(csa_tree_add_7_25_groupi_n_5539 ,csa_tree_add_7_25_groupi_n_5389 ,csa_tree_add_7_25_groupi_n_5470);
  and csa_tree_add_7_25_groupi_g15546(csa_tree_add_7_25_groupi_n_5538 ,csa_tree_add_7_25_groupi_n_5471 ,csa_tree_add_7_25_groupi_n_5391);
  or csa_tree_add_7_25_groupi_g15547(csa_tree_add_7_25_groupi_n_5537 ,csa_tree_add_7_25_groupi_n_5471 ,csa_tree_add_7_25_groupi_n_5391);
  or csa_tree_add_7_25_groupi_g15548(csa_tree_add_7_25_groupi_n_5536 ,csa_tree_add_7_25_groupi_n_5468 ,csa_tree_add_7_25_groupi_n_5392);
  and csa_tree_add_7_25_groupi_g15549(csa_tree_add_7_25_groupi_n_5535 ,csa_tree_add_7_25_groupi_n_5468 ,csa_tree_add_7_25_groupi_n_5392);
  and csa_tree_add_7_25_groupi_g15550(csa_tree_add_7_25_groupi_n_5556 ,csa_tree_add_7_25_groupi_n_2439 ,csa_tree_add_7_25_groupi_n_5506);
  or csa_tree_add_7_25_groupi_g15551(csa_tree_add_7_25_groupi_n_5555 ,csa_tree_add_7_25_groupi_n_5441 ,csa_tree_add_7_25_groupi_n_5500);
  or csa_tree_add_7_25_groupi_g15552(csa_tree_add_7_25_groupi_n_5554 ,csa_tree_add_7_25_groupi_n_5421 ,csa_tree_add_7_25_groupi_n_5504);
  or csa_tree_add_7_25_groupi_g15553(csa_tree_add_7_25_groupi_n_5552 ,csa_tree_add_7_25_groupi_n_5439 ,csa_tree_add_7_25_groupi_n_5505);
  and csa_tree_add_7_25_groupi_g15554(csa_tree_add_7_25_groupi_n_5532 ,csa_tree_add_7_25_groupi_n_5474 ,csa_tree_add_7_25_groupi_n_5297);
  or csa_tree_add_7_25_groupi_g15555(csa_tree_add_7_25_groupi_n_5531 ,csa_tree_add_7_25_groupi_n_3268 ,csa_tree_add_7_25_groupi_n_5499);
  or csa_tree_add_7_25_groupi_g15556(csa_tree_add_7_25_groupi_n_5530 ,csa_tree_add_7_25_groupi_n_3232 ,csa_tree_add_7_25_groupi_n_5496);
  and csa_tree_add_7_25_groupi_g15557(csa_tree_add_7_25_groupi_n_5529 ,csa_tree_add_7_25_groupi_n_5475 ,csa_tree_add_7_25_groupi_n_5294);
  or csa_tree_add_7_25_groupi_g15558(csa_tree_add_7_25_groupi_n_5528 ,csa_tree_add_7_25_groupi_n_3078 ,csa_tree_add_7_25_groupi_n_5501);
  or csa_tree_add_7_25_groupi_g15559(csa_tree_add_7_25_groupi_n_5527 ,csa_tree_add_7_25_groupi_n_3219 ,csa_tree_add_7_25_groupi_n_5495);
  or csa_tree_add_7_25_groupi_g15560(csa_tree_add_7_25_groupi_n_5526 ,csa_tree_add_7_25_groupi_n_3218 ,csa_tree_add_7_25_groupi_n_5494);
  or csa_tree_add_7_25_groupi_g15561(csa_tree_add_7_25_groupi_n_5525 ,csa_tree_add_7_25_groupi_n_3220 ,csa_tree_add_7_25_groupi_n_5493);
  or csa_tree_add_7_25_groupi_g15562(csa_tree_add_7_25_groupi_n_5524 ,csa_tree_add_7_25_groupi_n_3655 ,csa_tree_add_7_25_groupi_n_5502);
  or csa_tree_add_7_25_groupi_g15563(csa_tree_add_7_25_groupi_n_5523 ,csa_tree_add_7_25_groupi_n_3659 ,csa_tree_add_7_25_groupi_n_5507);
  or csa_tree_add_7_25_groupi_g15564(csa_tree_add_7_25_groupi_n_5522 ,csa_tree_add_7_25_groupi_n_3661 ,csa_tree_add_7_25_groupi_n_5498);
  or csa_tree_add_7_25_groupi_g15565(csa_tree_add_7_25_groupi_n_5521 ,csa_tree_add_7_25_groupi_n_3660 ,csa_tree_add_7_25_groupi_n_5497);
  or csa_tree_add_7_25_groupi_g15566(csa_tree_add_7_25_groupi_n_5520 ,csa_tree_add_7_25_groupi_n_5465 ,csa_tree_add_7_25_groupi_n_5395);
  and csa_tree_add_7_25_groupi_g15567(csa_tree_add_7_25_groupi_n_5519 ,csa_tree_add_7_25_groupi_n_5465 ,csa_tree_add_7_25_groupi_n_5395);
  and csa_tree_add_7_25_groupi_g15568(csa_tree_add_7_25_groupi_n_5518 ,csa_tree_add_7_25_groupi_n_5466 ,csa_tree_add_7_25_groupi_n_5393);
  or csa_tree_add_7_25_groupi_g15569(csa_tree_add_7_25_groupi_n_5517 ,csa_tree_add_7_25_groupi_n_5466 ,csa_tree_add_7_25_groupi_n_5393);
  and csa_tree_add_7_25_groupi_g15570(csa_tree_add_7_25_groupi_n_5516 ,csa_tree_add_7_25_groupi_n_5467 ,csa_tree_add_7_25_groupi_n_5394);
  or csa_tree_add_7_25_groupi_g15571(csa_tree_add_7_25_groupi_n_5515 ,csa_tree_add_7_25_groupi_n_5467 ,csa_tree_add_7_25_groupi_n_5394);
  or csa_tree_add_7_25_groupi_g15572(csa_tree_add_7_25_groupi_n_5534 ,csa_tree_add_7_25_groupi_n_5415 ,csa_tree_add_7_25_groupi_n_5503);
  xnor csa_tree_add_7_25_groupi_g15573(csa_tree_add_7_25_groupi_n_5533 ,csa_tree_add_7_25_groupi_n_5447 ,csa_tree_add_7_25_groupi_n_2572);
  nor csa_tree_add_7_25_groupi_g15574(csa_tree_add_7_25_groupi_n_5507 ,csa_tree_add_7_25_groupi_n_1934 ,csa_tree_add_7_25_groupi_n_185);
  or csa_tree_add_7_25_groupi_g15575(csa_tree_add_7_25_groupi_n_5506 ,csa_tree_add_7_25_groupi_n_2474 ,csa_tree_add_7_25_groupi_n_5447);
  and csa_tree_add_7_25_groupi_g15576(csa_tree_add_7_25_groupi_n_5505 ,csa_tree_add_7_25_groupi_n_5397 ,csa_tree_add_7_25_groupi_n_5442);
  and csa_tree_add_7_25_groupi_g15577(csa_tree_add_7_25_groupi_n_5504 ,csa_tree_add_7_25_groupi_n_5398 ,csa_tree_add_7_25_groupi_n_5420);
  and csa_tree_add_7_25_groupi_g15578(csa_tree_add_7_25_groupi_n_5503 ,csa_tree_add_7_25_groupi_n_5396 ,csa_tree_add_7_25_groupi_n_5414);
  nor csa_tree_add_7_25_groupi_g15579(csa_tree_add_7_25_groupi_n_5502 ,csa_tree_add_7_25_groupi_n_1856 ,csa_tree_add_7_25_groupi_n_1319);
  nor csa_tree_add_7_25_groupi_g15580(csa_tree_add_7_25_groupi_n_5501 ,csa_tree_add_7_25_groupi_n_2178 ,csa_tree_add_7_25_groupi_n_1819);
  and csa_tree_add_7_25_groupi_g15581(csa_tree_add_7_25_groupi_n_5500 ,csa_tree_add_7_25_groupi_n_5440 ,csa_tree_add_7_25_groupi_n_5446);
  nor csa_tree_add_7_25_groupi_g15582(csa_tree_add_7_25_groupi_n_5499 ,csa_tree_add_7_25_groupi_n_2022 ,csa_tree_add_7_25_groupi_n_1856);
  nor csa_tree_add_7_25_groupi_g15583(csa_tree_add_7_25_groupi_n_5498 ,csa_tree_add_7_25_groupi_n_2049 ,csa_tree_add_7_25_groupi_n_190);
  nor csa_tree_add_7_25_groupi_g15584(csa_tree_add_7_25_groupi_n_5497 ,csa_tree_add_7_25_groupi_n_2067 ,csa_tree_add_7_25_groupi_n_185);
  nor csa_tree_add_7_25_groupi_g15585(csa_tree_add_7_25_groupi_n_5496 ,csa_tree_add_7_25_groupi_n_2136 ,csa_tree_add_7_25_groupi_n_190);
  nor csa_tree_add_7_25_groupi_g15586(csa_tree_add_7_25_groupi_n_5495 ,csa_tree_add_7_25_groupi_n_2100 ,csa_tree_add_7_25_groupi_n_1818);
  nor csa_tree_add_7_25_groupi_g15587(csa_tree_add_7_25_groupi_n_5494 ,csa_tree_add_7_25_groupi_n_2121 ,csa_tree_add_7_25_groupi_n_189);
  nor csa_tree_add_7_25_groupi_g15588(csa_tree_add_7_25_groupi_n_5493 ,csa_tree_add_7_25_groupi_n_2151 ,csa_tree_add_7_25_groupi_n_1818);
  nor csa_tree_add_7_25_groupi_g15589(csa_tree_add_7_25_groupi_n_5492 ,csa_tree_add_7_25_groupi_n_3854 ,csa_tree_add_7_25_groupi_n_5408);
  nor csa_tree_add_7_25_groupi_g15590(csa_tree_add_7_25_groupi_n_5491 ,csa_tree_add_7_25_groupi_n_4074 ,csa_tree_add_7_25_groupi_n_5413);
  nor csa_tree_add_7_25_groupi_g15591(csa_tree_add_7_25_groupi_n_5490 ,csa_tree_add_7_25_groupi_n_3884 ,csa_tree_add_7_25_groupi_n_5406);
  nor csa_tree_add_7_25_groupi_g15592(csa_tree_add_7_25_groupi_n_5489 ,csa_tree_add_7_25_groupi_n_3846 ,csa_tree_add_7_25_groupi_n_5407);
  nor csa_tree_add_7_25_groupi_g15593(csa_tree_add_7_25_groupi_n_5488 ,csa_tree_add_7_25_groupi_n_4024 ,csa_tree_add_7_25_groupi_n_5417);
  nor csa_tree_add_7_25_groupi_g15594(csa_tree_add_7_25_groupi_n_5487 ,csa_tree_add_7_25_groupi_n_3859 ,csa_tree_add_7_25_groupi_n_5409);
  nor csa_tree_add_7_25_groupi_g15595(csa_tree_add_7_25_groupi_n_5486 ,csa_tree_add_7_25_groupi_n_3481 ,csa_tree_add_7_25_groupi_n_5399);
  nor csa_tree_add_7_25_groupi_g15596(csa_tree_add_7_25_groupi_n_5485 ,csa_tree_add_7_25_groupi_n_4006 ,csa_tree_add_7_25_groupi_n_5422);
  nor csa_tree_add_7_25_groupi_g15597(csa_tree_add_7_25_groupi_n_5484 ,csa_tree_add_7_25_groupi_n_4049 ,csa_tree_add_7_25_groupi_n_5411);
  nor csa_tree_add_7_25_groupi_g15598(csa_tree_add_7_25_groupi_n_5483 ,csa_tree_add_7_25_groupi_n_4062 ,csa_tree_add_7_25_groupi_n_5412);
  nor csa_tree_add_7_25_groupi_g15599(csa_tree_add_7_25_groupi_n_5482 ,csa_tree_add_7_25_groupi_n_3921 ,csa_tree_add_7_25_groupi_n_5403);
  or csa_tree_add_7_25_groupi_g15600(csa_tree_add_7_25_groupi_n_5514 ,csa_tree_add_7_25_groupi_n_5192 ,csa_tree_add_7_25_groupi_n_5410);
  or csa_tree_add_7_25_groupi_g15601(csa_tree_add_7_25_groupi_n_5513 ,csa_tree_add_7_25_groupi_n_5178 ,csa_tree_add_7_25_groupi_n_5402);
  or csa_tree_add_7_25_groupi_g15602(csa_tree_add_7_25_groupi_n_5512 ,csa_tree_add_7_25_groupi_n_5177 ,csa_tree_add_7_25_groupi_n_5401);
  or csa_tree_add_7_25_groupi_g15603(csa_tree_add_7_25_groupi_n_5511 ,csa_tree_add_7_25_groupi_n_5174 ,csa_tree_add_7_25_groupi_n_5400);
  or csa_tree_add_7_25_groupi_g15604(csa_tree_add_7_25_groupi_n_5510 ,csa_tree_add_7_25_groupi_n_5197 ,csa_tree_add_7_25_groupi_n_5425);
  or csa_tree_add_7_25_groupi_g15605(csa_tree_add_7_25_groupi_n_5509 ,csa_tree_add_7_25_groupi_n_5195 ,csa_tree_add_7_25_groupi_n_5424);
  or csa_tree_add_7_25_groupi_g15606(csa_tree_add_7_25_groupi_n_5508 ,csa_tree_add_7_25_groupi_n_5189 ,csa_tree_add_7_25_groupi_n_5416);
  not csa_tree_add_7_25_groupi_g15607(csa_tree_add_7_25_groupi_n_5463 ,csa_tree_add_7_25_groupi_n_5464);
  xnor csa_tree_add_7_25_groupi_g15608(out2[6] ,csa_tree_add_7_25_groupi_n_5304 ,csa_tree_add_7_25_groupi_n_5334);
  xnor csa_tree_add_7_25_groupi_g15609(csa_tree_add_7_25_groupi_n_5461 ,csa_tree_add_7_25_groupi_n_5279 ,csa_tree_add_7_25_groupi_n_5345);
  xnor csa_tree_add_7_25_groupi_g15610(csa_tree_add_7_25_groupi_n_5460 ,csa_tree_add_7_25_groupi_n_5342 ,csa_tree_add_7_25_groupi_n_5120);
  xnor csa_tree_add_7_25_groupi_g15611(csa_tree_add_7_25_groupi_n_5459 ,csa_tree_add_7_25_groupi_n_5356 ,csa_tree_add_7_25_groupi_n_5227);
  xnor csa_tree_add_7_25_groupi_g15612(csa_tree_add_7_25_groupi_n_5458 ,csa_tree_add_7_25_groupi_n_5269 ,csa_tree_add_7_25_groupi_n_5350);
  xnor csa_tree_add_7_25_groupi_g15613(csa_tree_add_7_25_groupi_n_5457 ,csa_tree_add_7_25_groupi_n_5276 ,csa_tree_add_7_25_groupi_n_5347);
  xnor csa_tree_add_7_25_groupi_g15614(csa_tree_add_7_25_groupi_n_5456 ,csa_tree_add_7_25_groupi_n_5343 ,csa_tree_add_7_25_groupi_n_5232);
  xnor csa_tree_add_7_25_groupi_g15615(csa_tree_add_7_25_groupi_n_5455 ,csa_tree_add_7_25_groupi_n_5388 ,csa_tree_add_7_25_groupi_n_5386);
  xnor csa_tree_add_7_25_groupi_g15616(csa_tree_add_7_25_groupi_n_5454 ,csa_tree_add_7_25_groupi_n_5277 ,csa_tree_add_7_25_groupi_n_5349);
  xnor csa_tree_add_7_25_groupi_g15617(csa_tree_add_7_25_groupi_n_5453 ,csa_tree_add_7_25_groupi_n_5274 ,csa_tree_add_7_25_groupi_n_5348);
  xnor csa_tree_add_7_25_groupi_g15618(csa_tree_add_7_25_groupi_n_5452 ,csa_tree_add_7_25_groupi_n_5272 ,csa_tree_add_7_25_groupi_n_5351);
  xnor csa_tree_add_7_25_groupi_g15619(csa_tree_add_7_25_groupi_n_5451 ,csa_tree_add_7_25_groupi_n_5271 ,csa_tree_add_7_25_groupi_n_5352);
  xnor csa_tree_add_7_25_groupi_g15620(csa_tree_add_7_25_groupi_n_5450 ,csa_tree_add_7_25_groupi_n_5270 ,csa_tree_add_7_25_groupi_n_5353);
  xnor csa_tree_add_7_25_groupi_g15621(csa_tree_add_7_25_groupi_n_5449 ,csa_tree_add_7_25_groupi_n_5273 ,csa_tree_add_7_25_groupi_n_5354);
  xnor csa_tree_add_7_25_groupi_g15622(csa_tree_add_7_25_groupi_n_5448 ,csa_tree_add_7_25_groupi_n_5280 ,csa_tree_add_7_25_groupi_n_5357);
  xnor csa_tree_add_7_25_groupi_g15623(csa_tree_add_7_25_groupi_n_5481 ,csa_tree_add_7_25_groupi_n_5371 ,in3[17]);
  xnor csa_tree_add_7_25_groupi_g15624(csa_tree_add_7_25_groupi_n_5480 ,csa_tree_add_7_25_groupi_n_5370 ,in3[2]);
  xnor csa_tree_add_7_25_groupi_g15625(csa_tree_add_7_25_groupi_n_5479 ,csa_tree_add_7_25_groupi_n_5366 ,in3[14]);
  xnor csa_tree_add_7_25_groupi_g15626(csa_tree_add_7_25_groupi_n_5478 ,csa_tree_add_7_25_groupi_n_5372 ,in3[11]);
  xnor csa_tree_add_7_25_groupi_g15627(csa_tree_add_7_25_groupi_n_5477 ,csa_tree_add_7_25_groupi_n_5369 ,in3[8]);
  xnor csa_tree_add_7_25_groupi_g15628(csa_tree_add_7_25_groupi_n_5476 ,csa_tree_add_7_25_groupi_n_5374 ,in3[5]);
  xnor csa_tree_add_7_25_groupi_g15629(csa_tree_add_7_25_groupi_n_5475 ,csa_tree_add_7_25_groupi_n_5368 ,in3[20]);
  xnor csa_tree_add_7_25_groupi_g15630(csa_tree_add_7_25_groupi_n_5474 ,csa_tree_add_7_25_groupi_n_5365 ,in3[26]);
  xnor csa_tree_add_7_25_groupi_g15631(csa_tree_add_7_25_groupi_n_5473 ,csa_tree_add_7_25_groupi_n_5367 ,in3[23]);
  xnor csa_tree_add_7_25_groupi_g15632(csa_tree_add_7_25_groupi_n_5472 ,csa_tree_add_7_25_groupi_n_5373 ,in3[29]);
  xnor csa_tree_add_7_25_groupi_g15633(csa_tree_add_7_25_groupi_n_5471 ,csa_tree_add_7_25_groupi_n_5361 ,csa_tree_add_7_25_groupi_n_5213);
  xnor csa_tree_add_7_25_groupi_g15634(csa_tree_add_7_25_groupi_n_5470 ,csa_tree_add_7_25_groupi_n_5358 ,csa_tree_add_7_25_groupi_n_5219);
  xnor csa_tree_add_7_25_groupi_g15635(csa_tree_add_7_25_groupi_n_5469 ,csa_tree_add_7_25_groupi_n_5364 ,csa_tree_add_7_25_groupi_n_5220);
  xnor csa_tree_add_7_25_groupi_g15636(csa_tree_add_7_25_groupi_n_5468 ,csa_tree_add_7_25_groupi_n_5360 ,csa_tree_add_7_25_groupi_n_5221);
  xnor csa_tree_add_7_25_groupi_g15637(csa_tree_add_7_25_groupi_n_5467 ,csa_tree_add_7_25_groupi_n_5363 ,csa_tree_add_7_25_groupi_n_5217);
  xnor csa_tree_add_7_25_groupi_g15638(csa_tree_add_7_25_groupi_n_5466 ,csa_tree_add_7_25_groupi_n_5362 ,csa_tree_add_7_25_groupi_n_5216);
  xnor csa_tree_add_7_25_groupi_g15639(csa_tree_add_7_25_groupi_n_5465 ,csa_tree_add_7_25_groupi_n_5359 ,csa_tree_add_7_25_groupi_n_5214);
  xnor csa_tree_add_7_25_groupi_g15640(csa_tree_add_7_25_groupi_n_5464 ,csa_tree_add_7_25_groupi_n_5337 ,csa_tree_add_7_25_groupi_n_5156);
  or csa_tree_add_7_25_groupi_g15641(csa_tree_add_7_25_groupi_n_5445 ,csa_tree_add_7_25_groupi_n_5269 ,csa_tree_add_7_25_groupi_n_5350);
  nor csa_tree_add_7_25_groupi_g15642(csa_tree_add_7_25_groupi_n_5444 ,csa_tree_add_7_25_groupi_n_2346 ,csa_tree_add_7_25_groupi_n_5388);
  or csa_tree_add_7_25_groupi_g15643(csa_tree_add_7_25_groupi_n_5443 ,csa_tree_add_7_25_groupi_n_1973 ,csa_tree_add_7_25_groupi_n_5387);
  or csa_tree_add_7_25_groupi_g15644(csa_tree_add_7_25_groupi_n_5442 ,csa_tree_add_7_25_groupi_n_5342 ,csa_tree_add_7_25_groupi_n_5119);
  and csa_tree_add_7_25_groupi_g15645(csa_tree_add_7_25_groupi_n_5441 ,csa_tree_add_7_25_groupi_n_5280 ,csa_tree_add_7_25_groupi_n_5357);
  or csa_tree_add_7_25_groupi_g15646(csa_tree_add_7_25_groupi_n_5440 ,csa_tree_add_7_25_groupi_n_5280 ,csa_tree_add_7_25_groupi_n_5357);
  nor csa_tree_add_7_25_groupi_g15647(csa_tree_add_7_25_groupi_n_5439 ,csa_tree_add_7_25_groupi_n_5341 ,csa_tree_add_7_25_groupi_n_5120);
  and csa_tree_add_7_25_groupi_g15648(csa_tree_add_7_25_groupi_n_5438 ,csa_tree_add_7_25_groupi_n_5269 ,csa_tree_add_7_25_groupi_n_5350);
  and csa_tree_add_7_25_groupi_g15649(csa_tree_add_7_25_groupi_n_5437 ,csa_tree_add_7_25_groupi_n_5273 ,csa_tree_add_7_25_groupi_n_5354);
  or csa_tree_add_7_25_groupi_g15650(csa_tree_add_7_25_groupi_n_5436 ,csa_tree_add_7_25_groupi_n_5273 ,csa_tree_add_7_25_groupi_n_5354);
  and csa_tree_add_7_25_groupi_g15651(csa_tree_add_7_25_groupi_n_5435 ,csa_tree_add_7_25_groupi_n_5270 ,csa_tree_add_7_25_groupi_n_5353);
  or csa_tree_add_7_25_groupi_g15652(csa_tree_add_7_25_groupi_n_5434 ,csa_tree_add_7_25_groupi_n_5270 ,csa_tree_add_7_25_groupi_n_5353);
  and csa_tree_add_7_25_groupi_g15653(csa_tree_add_7_25_groupi_n_5433 ,csa_tree_add_7_25_groupi_n_5277 ,csa_tree_add_7_25_groupi_n_5349);
  or csa_tree_add_7_25_groupi_g15654(csa_tree_add_7_25_groupi_n_5432 ,csa_tree_add_7_25_groupi_n_5277 ,csa_tree_add_7_25_groupi_n_5349);
  and csa_tree_add_7_25_groupi_g15655(csa_tree_add_7_25_groupi_n_5431 ,csa_tree_add_7_25_groupi_n_5271 ,csa_tree_add_7_25_groupi_n_5352);
  or csa_tree_add_7_25_groupi_g15656(csa_tree_add_7_25_groupi_n_5430 ,csa_tree_add_7_25_groupi_n_5271 ,csa_tree_add_7_25_groupi_n_5352);
  and csa_tree_add_7_25_groupi_g15657(csa_tree_add_7_25_groupi_n_5429 ,csa_tree_add_7_25_groupi_n_5272 ,csa_tree_add_7_25_groupi_n_5351);
  or csa_tree_add_7_25_groupi_g15658(csa_tree_add_7_25_groupi_n_5428 ,csa_tree_add_7_25_groupi_n_5272 ,csa_tree_add_7_25_groupi_n_5351);
  and csa_tree_add_7_25_groupi_g15659(csa_tree_add_7_25_groupi_n_5427 ,csa_tree_add_7_25_groupi_n_5274 ,csa_tree_add_7_25_groupi_n_5348);
  or csa_tree_add_7_25_groupi_g15660(csa_tree_add_7_25_groupi_n_5426 ,csa_tree_add_7_25_groupi_n_5274 ,csa_tree_add_7_25_groupi_n_5348);
  and csa_tree_add_7_25_groupi_g15661(csa_tree_add_7_25_groupi_n_5425 ,csa_tree_add_7_25_groupi_n_5361 ,csa_tree_add_7_25_groupi_n_5196);
  and csa_tree_add_7_25_groupi_g15662(csa_tree_add_7_25_groupi_n_5424 ,csa_tree_add_7_25_groupi_n_5360 ,csa_tree_add_7_25_groupi_n_5194);
  and csa_tree_add_7_25_groupi_g15663(csa_tree_add_7_25_groupi_n_5447 ,csa_tree_add_7_25_groupi_n_2477 ,csa_tree_add_7_25_groupi_n_5383);
  or csa_tree_add_7_25_groupi_g15664(csa_tree_add_7_25_groupi_n_5446 ,csa_tree_add_7_25_groupi_n_5324 ,csa_tree_add_7_25_groupi_n_5380);
  or csa_tree_add_7_25_groupi_g15665(csa_tree_add_7_25_groupi_n_5422 ,csa_tree_add_7_25_groupi_n_3217 ,csa_tree_add_7_25_groupi_n_5339);
  nor csa_tree_add_7_25_groupi_g15666(csa_tree_add_7_25_groupi_n_5421 ,csa_tree_add_7_25_groupi_n_5355 ,csa_tree_add_7_25_groupi_n_5227);
  or csa_tree_add_7_25_groupi_g15667(csa_tree_add_7_25_groupi_n_5420 ,csa_tree_add_7_25_groupi_n_5356 ,csa_tree_add_7_25_groupi_n_5226);
  nor csa_tree_add_7_25_groupi_g15668(csa_tree_add_7_25_groupi_n_5419 ,csa_tree_add_7_25_groupi_n_5278 ,csa_tree_add_7_25_groupi_n_5345);
  or csa_tree_add_7_25_groupi_g15669(csa_tree_add_7_25_groupi_n_5418 ,csa_tree_add_7_25_groupi_n_5279 ,csa_tree_add_7_25_groupi_n_5344);
  or csa_tree_add_7_25_groupi_g15670(csa_tree_add_7_25_groupi_n_5417 ,csa_tree_add_7_25_groupi_n_3253 ,csa_tree_add_7_25_groupi_n_5375);
  and csa_tree_add_7_25_groupi_g15671(csa_tree_add_7_25_groupi_n_5416 ,csa_tree_add_7_25_groupi_n_5358 ,csa_tree_add_7_25_groupi_n_5193);
  and csa_tree_add_7_25_groupi_g15672(csa_tree_add_7_25_groupi_n_5415 ,csa_tree_add_7_25_groupi_n_5343 ,csa_tree_add_7_25_groupi_n_5232);
  or csa_tree_add_7_25_groupi_g15673(csa_tree_add_7_25_groupi_n_5414 ,csa_tree_add_7_25_groupi_n_5343 ,csa_tree_add_7_25_groupi_n_5232);
  or csa_tree_add_7_25_groupi_g15674(csa_tree_add_7_25_groupi_n_5413 ,csa_tree_add_7_25_groupi_n_3200 ,csa_tree_add_7_25_groupi_n_5382);
  or csa_tree_add_7_25_groupi_g15675(csa_tree_add_7_25_groupi_n_5412 ,csa_tree_add_7_25_groupi_n_3338 ,csa_tree_add_7_25_groupi_n_5384);
  or csa_tree_add_7_25_groupi_g15676(csa_tree_add_7_25_groupi_n_5411 ,csa_tree_add_7_25_groupi_n_3318 ,csa_tree_add_7_25_groupi_n_5340);
  and csa_tree_add_7_25_groupi_g15677(csa_tree_add_7_25_groupi_n_5410 ,csa_tree_add_7_25_groupi_n_5364 ,csa_tree_add_7_25_groupi_n_5191);
  or csa_tree_add_7_25_groupi_g15678(csa_tree_add_7_25_groupi_n_5409 ,csa_tree_add_7_25_groupi_n_3603 ,csa_tree_add_7_25_groupi_n_5378);
  or csa_tree_add_7_25_groupi_g15679(csa_tree_add_7_25_groupi_n_5408 ,csa_tree_add_7_25_groupi_n_3639 ,csa_tree_add_7_25_groupi_n_5376);
  or csa_tree_add_7_25_groupi_g15680(csa_tree_add_7_25_groupi_n_5407 ,csa_tree_add_7_25_groupi_n_3622 ,csa_tree_add_7_25_groupi_n_5385);
  or csa_tree_add_7_25_groupi_g15681(csa_tree_add_7_25_groupi_n_5406 ,csa_tree_add_7_25_groupi_n_3594 ,csa_tree_add_7_25_groupi_n_5381);
  nor csa_tree_add_7_25_groupi_g15682(csa_tree_add_7_25_groupi_n_5405 ,csa_tree_add_7_25_groupi_n_5275 ,csa_tree_add_7_25_groupi_n_5347);
  or csa_tree_add_7_25_groupi_g15683(csa_tree_add_7_25_groupi_n_5404 ,csa_tree_add_7_25_groupi_n_5276 ,csa_tree_add_7_25_groupi_n_5346);
  or csa_tree_add_7_25_groupi_g15684(csa_tree_add_7_25_groupi_n_5403 ,csa_tree_add_7_25_groupi_n_3055 ,csa_tree_add_7_25_groupi_n_5379);
  and csa_tree_add_7_25_groupi_g15685(csa_tree_add_7_25_groupi_n_5402 ,csa_tree_add_7_25_groupi_n_5359 ,csa_tree_add_7_25_groupi_n_5173);
  and csa_tree_add_7_25_groupi_g15686(csa_tree_add_7_25_groupi_n_5401 ,csa_tree_add_7_25_groupi_n_5362 ,csa_tree_add_7_25_groupi_n_5175);
  and csa_tree_add_7_25_groupi_g15687(csa_tree_add_7_25_groupi_n_5400 ,csa_tree_add_7_25_groupi_n_5363 ,csa_tree_add_7_25_groupi_n_5187);
  or csa_tree_add_7_25_groupi_g15688(csa_tree_add_7_25_groupi_n_5399 ,csa_tree_add_7_25_groupi_n_3074 ,csa_tree_add_7_25_groupi_n_5377);
  xnor csa_tree_add_7_25_groupi_g15689(csa_tree_add_7_25_groupi_n_5423 ,csa_tree_add_7_25_groupi_n_5326 ,csa_tree_add_7_25_groupi_n_2573);
  not csa_tree_add_7_25_groupi_g15690(csa_tree_add_7_25_groupi_n_5387 ,csa_tree_add_7_25_groupi_n_5388);
  nor csa_tree_add_7_25_groupi_g15692(csa_tree_add_7_25_groupi_n_5385 ,csa_tree_add_7_25_groupi_n_261 ,csa_tree_add_7_25_groupi_n_2042);
  nor csa_tree_add_7_25_groupi_g15693(csa_tree_add_7_25_groupi_n_5384 ,csa_tree_add_7_25_groupi_n_2738 ,csa_tree_add_7_25_groupi_n_181);
  or csa_tree_add_7_25_groupi_g15694(csa_tree_add_7_25_groupi_n_5383 ,csa_tree_add_7_25_groupi_n_2486 ,csa_tree_add_7_25_groupi_n_5326);
  nor csa_tree_add_7_25_groupi_g15695(csa_tree_add_7_25_groupi_n_5382 ,csa_tree_add_7_25_groupi_n_2746 ,csa_tree_add_7_25_groupi_n_181);
  nor csa_tree_add_7_25_groupi_g15696(csa_tree_add_7_25_groupi_n_5381 ,csa_tree_add_7_25_groupi_n_2066 ,csa_tree_add_7_25_groupi_n_1836);
  and csa_tree_add_7_25_groupi_g15697(csa_tree_add_7_25_groupi_n_5380 ,csa_tree_add_7_25_groupi_n_5304 ,csa_tree_add_7_25_groupi_n_5323);
  nor csa_tree_add_7_25_groupi_g15698(csa_tree_add_7_25_groupi_n_5379 ,csa_tree_add_7_25_groupi_n_636 ,csa_tree_add_7_25_groupi_n_261);
  nor csa_tree_add_7_25_groupi_g15699(csa_tree_add_7_25_groupi_n_5378 ,csa_tree_add_7_25_groupi_n_483 ,csa_tree_add_7_25_groupi_n_264);
  nor csa_tree_add_7_25_groupi_g15700(csa_tree_add_7_25_groupi_n_5377 ,csa_tree_add_7_25_groupi_n_264 ,csa_tree_add_7_25_groupi_n_2836);
  nor csa_tree_add_7_25_groupi_g15701(csa_tree_add_7_25_groupi_n_5376 ,csa_tree_add_7_25_groupi_n_260 ,csa_tree_add_7_25_groupi_n_1796);
  nor csa_tree_add_7_25_groupi_g15702(csa_tree_add_7_25_groupi_n_5375 ,csa_tree_add_7_25_groupi_n_2030 ,csa_tree_add_7_25_groupi_n_1836);
  nor csa_tree_add_7_25_groupi_g15703(csa_tree_add_7_25_groupi_n_5374 ,csa_tree_add_7_25_groupi_n_4034 ,csa_tree_add_7_25_groupi_n_5292);
  nor csa_tree_add_7_25_groupi_g15704(csa_tree_add_7_25_groupi_n_5373 ,csa_tree_add_7_25_groupi_n_3937 ,csa_tree_add_7_25_groupi_n_5293);
  nor csa_tree_add_7_25_groupi_g15705(csa_tree_add_7_25_groupi_n_5372 ,csa_tree_add_7_25_groupi_n_4088 ,csa_tree_add_7_25_groupi_n_5302);
  nor csa_tree_add_7_25_groupi_g15706(csa_tree_add_7_25_groupi_n_5371 ,csa_tree_add_7_25_groupi_n_3828 ,csa_tree_add_7_25_groupi_n_5285);
  nor csa_tree_add_7_25_groupi_g15707(csa_tree_add_7_25_groupi_n_5370 ,csa_tree_add_7_25_groupi_n_3472 ,csa_tree_add_7_25_groupi_n_5282);
  nor csa_tree_add_7_25_groupi_g15708(csa_tree_add_7_25_groupi_n_5369 ,csa_tree_add_7_25_groupi_n_4045 ,csa_tree_add_7_25_groupi_n_5290);
  nor csa_tree_add_7_25_groupi_g15709(csa_tree_add_7_25_groupi_n_5368 ,csa_tree_add_7_25_groupi_n_3851 ,csa_tree_add_7_25_groupi_n_5286);
  nor csa_tree_add_7_25_groupi_g15710(csa_tree_add_7_25_groupi_n_5367 ,csa_tree_add_7_25_groupi_n_3826 ,csa_tree_add_7_25_groupi_n_5287);
  nor csa_tree_add_7_25_groupi_g15711(csa_tree_add_7_25_groupi_n_5366 ,csa_tree_add_7_25_groupi_n_3983 ,csa_tree_add_7_25_groupi_n_5289);
  nor csa_tree_add_7_25_groupi_g15712(csa_tree_add_7_25_groupi_n_5365 ,csa_tree_add_7_25_groupi_n_3821 ,csa_tree_add_7_25_groupi_n_5288);
  or csa_tree_add_7_25_groupi_g15713(csa_tree_add_7_25_groupi_n_5398 ,csa_tree_add_7_25_groupi_n_5097 ,csa_tree_add_7_25_groupi_n_5296);
  or csa_tree_add_7_25_groupi_g15714(csa_tree_add_7_25_groupi_n_5397 ,csa_tree_add_7_25_groupi_n_4888 ,csa_tree_add_7_25_groupi_n_5299);
  or csa_tree_add_7_25_groupi_g15715(csa_tree_add_7_25_groupi_n_5396 ,csa_tree_add_7_25_groupi_n_5019 ,csa_tree_add_7_25_groupi_n_5318);
  or csa_tree_add_7_25_groupi_g15716(csa_tree_add_7_25_groupi_n_5395 ,csa_tree_add_7_25_groupi_n_5016 ,csa_tree_add_7_25_groupi_n_5315);
  or csa_tree_add_7_25_groupi_g15717(csa_tree_add_7_25_groupi_n_5394 ,csa_tree_add_7_25_groupi_n_5014 ,csa_tree_add_7_25_groupi_n_5325);
  or csa_tree_add_7_25_groupi_g15718(csa_tree_add_7_25_groupi_n_5393 ,csa_tree_add_7_25_groupi_n_5012 ,csa_tree_add_7_25_groupi_n_5309);
  or csa_tree_add_7_25_groupi_g15719(csa_tree_add_7_25_groupi_n_5392 ,csa_tree_add_7_25_groupi_n_5010 ,csa_tree_add_7_25_groupi_n_5306);
  or csa_tree_add_7_25_groupi_g15720(csa_tree_add_7_25_groupi_n_5391 ,csa_tree_add_7_25_groupi_n_4997 ,csa_tree_add_7_25_groupi_n_5320);
  or csa_tree_add_7_25_groupi_g15721(csa_tree_add_7_25_groupi_n_5390 ,csa_tree_add_7_25_groupi_n_5004 ,csa_tree_add_7_25_groupi_n_5300);
  or csa_tree_add_7_25_groupi_g15722(csa_tree_add_7_25_groupi_n_5389 ,csa_tree_add_7_25_groupi_n_5024 ,csa_tree_add_7_25_groupi_n_5314);
  and csa_tree_add_7_25_groupi_g15723(csa_tree_add_7_25_groupi_n_5388 ,csa_tree_add_7_25_groupi_n_5183 ,csa_tree_add_7_25_groupi_n_5322);
  and csa_tree_add_7_25_groupi_g15724(csa_tree_add_7_25_groupi_n_5386 ,csa_tree_add_7_25_groupi_n_3813 ,csa_tree_add_7_25_groupi_n_5283);
  not csa_tree_add_7_25_groupi_g15725(csa_tree_add_7_25_groupi_n_5355 ,csa_tree_add_7_25_groupi_n_5356);
  not csa_tree_add_7_25_groupi_g15726(csa_tree_add_7_25_groupi_n_5346 ,csa_tree_add_7_25_groupi_n_5347);
  not csa_tree_add_7_25_groupi_g15727(csa_tree_add_7_25_groupi_n_5344 ,csa_tree_add_7_25_groupi_n_5345);
  not csa_tree_add_7_25_groupi_g15728(csa_tree_add_7_25_groupi_n_5341 ,csa_tree_add_7_25_groupi_n_5342);
  nor csa_tree_add_7_25_groupi_g15729(csa_tree_add_7_25_groupi_n_5340 ,csa_tree_add_7_25_groupi_n_263 ,csa_tree_add_7_25_groupi_n_2742);
  nor csa_tree_add_7_25_groupi_g15730(csa_tree_add_7_25_groupi_n_5339 ,csa_tree_add_7_25_groupi_n_2750 ,csa_tree_add_7_25_groupi_n_1837);
  xnor csa_tree_add_7_25_groupi_g15731(out2[5] ,csa_tree_add_7_25_groupi_n_5211 ,csa_tree_add_7_25_groupi_n_5215);
  xnor csa_tree_add_7_25_groupi_g15732(csa_tree_add_7_25_groupi_n_5337 ,csa_tree_add_7_25_groupi_n_5281 ,in3[11]);
  xnor csa_tree_add_7_25_groupi_g15733(csa_tree_add_7_25_groupi_n_5336 ,csa_tree_add_7_25_groupi_n_5225 ,csa_tree_add_7_25_groupi_n_5210);
  xnor csa_tree_add_7_25_groupi_g15734(csa_tree_add_7_25_groupi_n_5335 ,csa_tree_add_7_25_groupi_n_5237 ,csa_tree_add_7_25_groupi_n_5159);
  xnor csa_tree_add_7_25_groupi_g15735(csa_tree_add_7_25_groupi_n_5334 ,csa_tree_add_7_25_groupi_n_5160 ,csa_tree_add_7_25_groupi_n_5235);
  xnor csa_tree_add_7_25_groupi_g15736(csa_tree_add_7_25_groupi_n_5333 ,csa_tree_add_7_25_groupi_n_5163 ,csa_tree_add_7_25_groupi_n_5236);
  xnor csa_tree_add_7_25_groupi_g15737(csa_tree_add_7_25_groupi_n_5332 ,csa_tree_add_7_25_groupi_n_5164 ,csa_tree_add_7_25_groupi_n_5234);
  xnor csa_tree_add_7_25_groupi_g15738(csa_tree_add_7_25_groupi_n_5331 ,csa_tree_add_7_25_groupi_n_5165 ,csa_tree_add_7_25_groupi_n_5231);
  xnor csa_tree_add_7_25_groupi_g15739(csa_tree_add_7_25_groupi_n_5330 ,csa_tree_add_7_25_groupi_n_5161 ,csa_tree_add_7_25_groupi_n_5230);
  xnor csa_tree_add_7_25_groupi_g15740(csa_tree_add_7_25_groupi_n_5329 ,csa_tree_add_7_25_groupi_n_5157 ,csa_tree_add_7_25_groupi_n_5233);
  xnor csa_tree_add_7_25_groupi_g15741(csa_tree_add_7_25_groupi_n_5328 ,csa_tree_add_7_25_groupi_n_5162 ,csa_tree_add_7_25_groupi_n_5229);
  xnor csa_tree_add_7_25_groupi_g15742(csa_tree_add_7_25_groupi_n_5327 ,csa_tree_add_7_25_groupi_n_5158 ,csa_tree_add_7_25_groupi_n_5228);
  xnor csa_tree_add_7_25_groupi_g15743(csa_tree_add_7_25_groupi_n_5364 ,csa_tree_add_7_25_groupi_n_5252 ,in3[17]);
  xnor csa_tree_add_7_25_groupi_g15744(csa_tree_add_7_25_groupi_n_5363 ,csa_tree_add_7_25_groupi_n_5251 ,in3[5]);
  xnor csa_tree_add_7_25_groupi_g15745(csa_tree_add_7_25_groupi_n_5362 ,csa_tree_add_7_25_groupi_n_5255 ,in3[8]);
  xnor csa_tree_add_7_25_groupi_g15746(csa_tree_add_7_25_groupi_n_5361 ,csa_tree_add_7_25_groupi_n_5249 ,in3[11]);
  xnor csa_tree_add_7_25_groupi_g15747(csa_tree_add_7_25_groupi_n_5360 ,csa_tree_add_7_25_groupi_n_5248 ,in3[14]);
  xnor csa_tree_add_7_25_groupi_g15748(csa_tree_add_7_25_groupi_n_5359 ,csa_tree_add_7_25_groupi_n_5256 ,in3[2]);
  xnor csa_tree_add_7_25_groupi_g15749(csa_tree_add_7_25_groupi_n_5358 ,csa_tree_add_7_25_groupi_n_5253 ,in3[20]);
  xnor csa_tree_add_7_25_groupi_g15750(csa_tree_add_7_25_groupi_n_5357 ,csa_tree_add_7_25_groupi_n_5243 ,csa_tree_add_7_25_groupi_n_5035);
  xnor csa_tree_add_7_25_groupi_g15751(csa_tree_add_7_25_groupi_n_5356 ,csa_tree_add_7_25_groupi_n_5254 ,in3[26]);
  xnor csa_tree_add_7_25_groupi_g15752(csa_tree_add_7_25_groupi_n_5354 ,csa_tree_add_7_25_groupi_n_5247 ,csa_tree_add_7_25_groupi_n_5033);
  xnor csa_tree_add_7_25_groupi_g15753(csa_tree_add_7_25_groupi_n_5353 ,csa_tree_add_7_25_groupi_n_5246 ,csa_tree_add_7_25_groupi_n_5032);
  xnor csa_tree_add_7_25_groupi_g15754(csa_tree_add_7_25_groupi_n_5352 ,csa_tree_add_7_25_groupi_n_5245 ,csa_tree_add_7_25_groupi_n_5031);
  xnor csa_tree_add_7_25_groupi_g15755(csa_tree_add_7_25_groupi_n_5351 ,csa_tree_add_7_25_groupi_n_5244 ,csa_tree_add_7_25_groupi_n_5030);
  xnor csa_tree_add_7_25_groupi_g15756(csa_tree_add_7_25_groupi_n_5350 ,csa_tree_add_7_25_groupi_n_5240 ,csa_tree_add_7_25_groupi_n_5027);
  xnor csa_tree_add_7_25_groupi_g15757(csa_tree_add_7_25_groupi_n_5349 ,csa_tree_add_7_25_groupi_n_5241 ,csa_tree_add_7_25_groupi_n_5037);
  xnor csa_tree_add_7_25_groupi_g15758(csa_tree_add_7_25_groupi_n_5348 ,csa_tree_add_7_25_groupi_n_5242 ,csa_tree_add_7_25_groupi_n_5029);
  xnor csa_tree_add_7_25_groupi_g15759(csa_tree_add_7_25_groupi_n_5347 ,csa_tree_add_7_25_groupi_n_5238 ,csa_tree_add_7_25_groupi_n_4947);
  xnor csa_tree_add_7_25_groupi_g15760(csa_tree_add_7_25_groupi_n_5345 ,csa_tree_add_7_25_groupi_n_5239 ,csa_tree_add_7_25_groupi_n_5109);
  xnor csa_tree_add_7_25_groupi_g15761(csa_tree_add_7_25_groupi_n_5343 ,csa_tree_add_7_25_groupi_n_5250 ,in3[23]);
  xnor csa_tree_add_7_25_groupi_g15762(csa_tree_add_7_25_groupi_n_5342 ,csa_tree_add_7_25_groupi_n_5257 ,in3[29]);
  and csa_tree_add_7_25_groupi_g15763(csa_tree_add_7_25_groupi_n_5325 ,csa_tree_add_7_25_groupi_n_5247 ,csa_tree_add_7_25_groupi_n_5013);
  and csa_tree_add_7_25_groupi_g15764(csa_tree_add_7_25_groupi_n_5324 ,csa_tree_add_7_25_groupi_n_5160 ,csa_tree_add_7_25_groupi_n_5235);
  or csa_tree_add_7_25_groupi_g15765(csa_tree_add_7_25_groupi_n_5323 ,csa_tree_add_7_25_groupi_n_5160 ,csa_tree_add_7_25_groupi_n_5235);
  or csa_tree_add_7_25_groupi_g15766(csa_tree_add_7_25_groupi_n_5322 ,csa_tree_add_7_25_groupi_n_5182 ,csa_tree_add_7_25_groupi_n_5281);
  and csa_tree_add_7_25_groupi_g15767(csa_tree_add_7_25_groupi_n_5321 ,csa_tree_add_7_25_groupi_n_5237 ,csa_tree_add_7_25_groupi_n_5159);
  and csa_tree_add_7_25_groupi_g15768(csa_tree_add_7_25_groupi_n_5320 ,csa_tree_add_7_25_groupi_n_5245 ,csa_tree_add_7_25_groupi_n_5005);
  or csa_tree_add_7_25_groupi_g15769(csa_tree_add_7_25_groupi_n_5319 ,csa_tree_add_7_25_groupi_n_5237 ,csa_tree_add_7_25_groupi_n_5159);
  and csa_tree_add_7_25_groupi_g15770(csa_tree_add_7_25_groupi_n_5318 ,csa_tree_add_7_25_groupi_n_5240 ,csa_tree_add_7_25_groupi_n_5018);
  and csa_tree_add_7_25_groupi_g15771(csa_tree_add_7_25_groupi_n_5317 ,csa_tree_add_7_25_groupi_n_5163 ,csa_tree_add_7_25_groupi_n_5236);
  or csa_tree_add_7_25_groupi_g15772(csa_tree_add_7_25_groupi_n_5316 ,csa_tree_add_7_25_groupi_n_5163 ,csa_tree_add_7_25_groupi_n_5236);
  and csa_tree_add_7_25_groupi_g15773(csa_tree_add_7_25_groupi_n_5315 ,csa_tree_add_7_25_groupi_n_5243 ,csa_tree_add_7_25_groupi_n_5015);
  and csa_tree_add_7_25_groupi_g15774(csa_tree_add_7_25_groupi_n_5314 ,csa_tree_add_7_25_groupi_n_5241 ,csa_tree_add_7_25_groupi_n_5017);
  and csa_tree_add_7_25_groupi_g15775(csa_tree_add_7_25_groupi_n_5313 ,csa_tree_add_7_25_groupi_n_5164 ,csa_tree_add_7_25_groupi_n_5234);
  or csa_tree_add_7_25_groupi_g15776(csa_tree_add_7_25_groupi_n_5312 ,csa_tree_add_7_25_groupi_n_5164 ,csa_tree_add_7_25_groupi_n_5234);
  and csa_tree_add_7_25_groupi_g15777(csa_tree_add_7_25_groupi_n_5311 ,csa_tree_add_7_25_groupi_n_5165 ,csa_tree_add_7_25_groupi_n_5231);
  or csa_tree_add_7_25_groupi_g15778(csa_tree_add_7_25_groupi_n_5310 ,csa_tree_add_7_25_groupi_n_5165 ,csa_tree_add_7_25_groupi_n_5231);
  and csa_tree_add_7_25_groupi_g15779(csa_tree_add_7_25_groupi_n_5309 ,csa_tree_add_7_25_groupi_n_5246 ,csa_tree_add_7_25_groupi_n_5011);
  and csa_tree_add_7_25_groupi_g15780(csa_tree_add_7_25_groupi_n_5308 ,csa_tree_add_7_25_groupi_n_5162 ,csa_tree_add_7_25_groupi_n_5229);
  or csa_tree_add_7_25_groupi_g15781(csa_tree_add_7_25_groupi_n_5307 ,csa_tree_add_7_25_groupi_n_5162 ,csa_tree_add_7_25_groupi_n_5229);
  and csa_tree_add_7_25_groupi_g15782(csa_tree_add_7_25_groupi_n_5306 ,csa_tree_add_7_25_groupi_n_5244 ,csa_tree_add_7_25_groupi_n_5009);
  and csa_tree_add_7_25_groupi_g15783(csa_tree_add_7_25_groupi_n_5305 ,csa_tree_add_7_25_groupi_n_5161 ,csa_tree_add_7_25_groupi_n_5230);
  and csa_tree_add_7_25_groupi_g15784(csa_tree_add_7_25_groupi_n_5326 ,csa_tree_add_7_25_groupi_n_2424 ,csa_tree_add_7_25_groupi_n_5263);
  or csa_tree_add_7_25_groupi_g15785(csa_tree_add_7_25_groupi_n_5302 ,csa_tree_add_7_25_groupi_n_3166 ,csa_tree_add_7_25_groupi_n_5267);
  or csa_tree_add_7_25_groupi_g15786(csa_tree_add_7_25_groupi_n_5301 ,csa_tree_add_7_25_groupi_n_5158 ,csa_tree_add_7_25_groupi_n_5228);
  and csa_tree_add_7_25_groupi_g15787(csa_tree_add_7_25_groupi_n_5300 ,csa_tree_add_7_25_groupi_n_5242 ,csa_tree_add_7_25_groupi_n_5003);
  and csa_tree_add_7_25_groupi_g15788(csa_tree_add_7_25_groupi_n_5299 ,csa_tree_add_7_25_groupi_n_4887 ,csa_tree_add_7_25_groupi_n_5238);
  nor csa_tree_add_7_25_groupi_g15789(csa_tree_add_7_25_groupi_n_5298 ,csa_tree_add_7_25_groupi_n_5225 ,csa_tree_add_7_25_groupi_n_5209);
  or csa_tree_add_7_25_groupi_g15790(csa_tree_add_7_25_groupi_n_5297 ,csa_tree_add_7_25_groupi_n_5224 ,csa_tree_add_7_25_groupi_n_5210);
  and csa_tree_add_7_25_groupi_g15791(csa_tree_add_7_25_groupi_n_5296 ,csa_tree_add_7_25_groupi_n_5239 ,csa_tree_add_7_25_groupi_n_5098);
  and csa_tree_add_7_25_groupi_g15792(csa_tree_add_7_25_groupi_n_5295 ,csa_tree_add_7_25_groupi_n_5157 ,csa_tree_add_7_25_groupi_n_5233);
  or csa_tree_add_7_25_groupi_g15793(csa_tree_add_7_25_groupi_n_5294 ,csa_tree_add_7_25_groupi_n_5157 ,csa_tree_add_7_25_groupi_n_5233);
  or csa_tree_add_7_25_groupi_g15794(csa_tree_add_7_25_groupi_n_5293 ,csa_tree_add_7_25_groupi_n_3570 ,csa_tree_add_7_25_groupi_n_5264);
  or csa_tree_add_7_25_groupi_g15795(csa_tree_add_7_25_groupi_n_5292 ,csa_tree_add_7_25_groupi_n_3169 ,csa_tree_add_7_25_groupi_n_5258);
  and csa_tree_add_7_25_groupi_g15796(csa_tree_add_7_25_groupi_n_5291 ,csa_tree_add_7_25_groupi_n_5158 ,csa_tree_add_7_25_groupi_n_5228);
  or csa_tree_add_7_25_groupi_g15797(csa_tree_add_7_25_groupi_n_5290 ,csa_tree_add_7_25_groupi_n_3168 ,csa_tree_add_7_25_groupi_n_5222);
  or csa_tree_add_7_25_groupi_g15798(csa_tree_add_7_25_groupi_n_5289 ,csa_tree_add_7_25_groupi_n_3167 ,csa_tree_add_7_25_groupi_n_5223);
  or csa_tree_add_7_25_groupi_g15799(csa_tree_add_7_25_groupi_n_5288 ,csa_tree_add_7_25_groupi_n_3592 ,csa_tree_add_7_25_groupi_n_5262);
  or csa_tree_add_7_25_groupi_g15800(csa_tree_add_7_25_groupi_n_5287 ,csa_tree_add_7_25_groupi_n_3599 ,csa_tree_add_7_25_groupi_n_5261);
  or csa_tree_add_7_25_groupi_g15801(csa_tree_add_7_25_groupi_n_5286 ,csa_tree_add_7_25_groupi_n_3635 ,csa_tree_add_7_25_groupi_n_5260);
  or csa_tree_add_7_25_groupi_g15802(csa_tree_add_7_25_groupi_n_5285 ,csa_tree_add_7_25_groupi_n_3583 ,csa_tree_add_7_25_groupi_n_5259);
  or csa_tree_add_7_25_groupi_g15803(csa_tree_add_7_25_groupi_n_5284 ,csa_tree_add_7_25_groupi_n_5161 ,csa_tree_add_7_25_groupi_n_5230);
  nor csa_tree_add_7_25_groupi_g15804(csa_tree_add_7_25_groupi_n_5283 ,csa_tree_add_7_25_groupi_n_2936 ,csa_tree_add_7_25_groupi_n_5265);
  or csa_tree_add_7_25_groupi_g15805(csa_tree_add_7_25_groupi_n_5282 ,csa_tree_add_7_25_groupi_n_3048 ,csa_tree_add_7_25_groupi_n_5268);
  or csa_tree_add_7_25_groupi_g15806(csa_tree_add_7_25_groupi_n_5304 ,csa_tree_add_7_25_groupi_n_5266 ,csa_tree_add_7_25_groupi_n_5172);
  xnor csa_tree_add_7_25_groupi_g15807(csa_tree_add_7_25_groupi_n_5303 ,csa_tree_add_7_25_groupi_n_5212 ,csa_tree_add_7_25_groupi_n_2574);
  not csa_tree_add_7_25_groupi_g15808(csa_tree_add_7_25_groupi_n_5278 ,csa_tree_add_7_25_groupi_n_5279);
  not csa_tree_add_7_25_groupi_g15809(csa_tree_add_7_25_groupi_n_5275 ,csa_tree_add_7_25_groupi_n_5276);
  nor csa_tree_add_7_25_groupi_g15810(csa_tree_add_7_25_groupi_n_5268 ,csa_tree_add_7_25_groupi_n_339 ,csa_tree_add_7_25_groupi_n_2175);
  nor csa_tree_add_7_25_groupi_g15811(csa_tree_add_7_25_groupi_n_5267 ,csa_tree_add_7_25_groupi_n_2097 ,csa_tree_add_7_25_groupi_n_1845);
  and csa_tree_add_7_25_groupi_g15812(csa_tree_add_7_25_groupi_n_5266 ,csa_tree_add_7_25_groupi_n_5171 ,csa_tree_add_7_25_groupi_n_5211);
  nor csa_tree_add_7_25_groupi_g15813(csa_tree_add_7_25_groupi_n_5265 ,csa_tree_add_7_25_groupi_n_639 ,csa_tree_add_7_25_groupi_n_1845);
  nor csa_tree_add_7_25_groupi_g15814(csa_tree_add_7_25_groupi_n_5264 ,csa_tree_add_7_25_groupi_n_1916 ,csa_tree_add_7_25_groupi_n_132);
  or csa_tree_add_7_25_groupi_g15815(csa_tree_add_7_25_groupi_n_5263 ,csa_tree_add_7_25_groupi_n_2448 ,csa_tree_add_7_25_groupi_n_5212);
  nor csa_tree_add_7_25_groupi_g15816(csa_tree_add_7_25_groupi_n_5262 ,csa_tree_add_7_25_groupi_n_336 ,csa_tree_add_7_25_groupi_n_1795);
  nor csa_tree_add_7_25_groupi_g15817(csa_tree_add_7_25_groupi_n_5261 ,csa_tree_add_7_25_groupi_n_335 ,csa_tree_add_7_25_groupi_n_1106);
  nor csa_tree_add_7_25_groupi_g15818(csa_tree_add_7_25_groupi_n_5260 ,csa_tree_add_7_25_groupi_n_336 ,csa_tree_add_7_25_groupi_n_2034);
  nor csa_tree_add_7_25_groupi_g15819(csa_tree_add_7_25_groupi_n_5259 ,csa_tree_add_7_25_groupi_n_338 ,csa_tree_add_7_25_groupi_n_2782);
  nor csa_tree_add_7_25_groupi_g15820(csa_tree_add_7_25_groupi_n_5258 ,csa_tree_add_7_25_groupi_n_2133 ,csa_tree_add_7_25_groupi_n_1846);
  nor csa_tree_add_7_25_groupi_g15821(csa_tree_add_7_25_groupi_n_5257 ,csa_tree_add_7_25_groupi_n_3941 ,csa_tree_add_7_25_groupi_n_5203);
  nor csa_tree_add_7_25_groupi_g15822(csa_tree_add_7_25_groupi_n_5256 ,csa_tree_add_7_25_groupi_n_3484 ,csa_tree_add_7_25_groupi_n_5170);
  nor csa_tree_add_7_25_groupi_g15823(csa_tree_add_7_25_groupi_n_5255 ,csa_tree_add_7_25_groupi_n_4005 ,csa_tree_add_7_25_groupi_n_5186);
  nor csa_tree_add_7_25_groupi_g15824(csa_tree_add_7_25_groupi_n_5254 ,csa_tree_add_7_25_groupi_n_4054 ,csa_tree_add_7_25_groupi_n_5184);
  nor csa_tree_add_7_25_groupi_g15825(csa_tree_add_7_25_groupi_n_5253 ,csa_tree_add_7_25_groupi_n_3876 ,csa_tree_add_7_25_groupi_n_5180);
  nor csa_tree_add_7_25_groupi_g15826(csa_tree_add_7_25_groupi_n_5252 ,csa_tree_add_7_25_groupi_n_4019 ,csa_tree_add_7_25_groupi_n_5208);
  nor csa_tree_add_7_25_groupi_g15827(csa_tree_add_7_25_groupi_n_5251 ,csa_tree_add_7_25_groupi_n_4091 ,csa_tree_add_7_25_groupi_n_5166);
  nor csa_tree_add_7_25_groupi_g15828(csa_tree_add_7_25_groupi_n_5250 ,csa_tree_add_7_25_groupi_n_3895 ,csa_tree_add_7_25_groupi_n_5181);
  nor csa_tree_add_7_25_groupi_g15829(csa_tree_add_7_25_groupi_n_5249 ,csa_tree_add_7_25_groupi_n_4077 ,csa_tree_add_7_25_groupi_n_5176);
  nor csa_tree_add_7_25_groupi_g15830(csa_tree_add_7_25_groupi_n_5248 ,csa_tree_add_7_25_groupi_n_4084 ,csa_tree_add_7_25_groupi_n_5185);
  and csa_tree_add_7_25_groupi_g15831(csa_tree_add_7_25_groupi_n_5281 ,csa_tree_add_7_25_groupi_n_3893 ,csa_tree_add_7_25_groupi_n_5179);
  or csa_tree_add_7_25_groupi_g15832(csa_tree_add_7_25_groupi_n_5280 ,csa_tree_add_7_25_groupi_n_4913 ,csa_tree_add_7_25_groupi_n_5201);
  or csa_tree_add_7_25_groupi_g15833(csa_tree_add_7_25_groupi_n_5279 ,csa_tree_add_7_25_groupi_n_5022 ,csa_tree_add_7_25_groupi_n_5206);
  or csa_tree_add_7_25_groupi_g15834(csa_tree_add_7_25_groupi_n_5277 ,csa_tree_add_7_25_groupi_n_4926 ,csa_tree_add_7_25_groupi_n_5207);
  or csa_tree_add_7_25_groupi_g15835(csa_tree_add_7_25_groupi_n_5276 ,csa_tree_add_7_25_groupi_n_4815 ,csa_tree_add_7_25_groupi_n_5205);
  or csa_tree_add_7_25_groupi_g15836(csa_tree_add_7_25_groupi_n_5274 ,csa_tree_add_7_25_groupi_n_4921 ,csa_tree_add_7_25_groupi_n_5204);
  or csa_tree_add_7_25_groupi_g15837(csa_tree_add_7_25_groupi_n_5273 ,csa_tree_add_7_25_groupi_n_4917 ,csa_tree_add_7_25_groupi_n_5202);
  or csa_tree_add_7_25_groupi_g15838(csa_tree_add_7_25_groupi_n_5272 ,csa_tree_add_7_25_groupi_n_4916 ,csa_tree_add_7_25_groupi_n_5200);
  or csa_tree_add_7_25_groupi_g15839(csa_tree_add_7_25_groupi_n_5271 ,csa_tree_add_7_25_groupi_n_4922 ,csa_tree_add_7_25_groupi_n_5199);
  or csa_tree_add_7_25_groupi_g15840(csa_tree_add_7_25_groupi_n_5270 ,csa_tree_add_7_25_groupi_n_4924 ,csa_tree_add_7_25_groupi_n_5198);
  or csa_tree_add_7_25_groupi_g15841(csa_tree_add_7_25_groupi_n_5269 ,csa_tree_add_7_25_groupi_n_4902 ,csa_tree_add_7_25_groupi_n_5190);
  not csa_tree_add_7_25_groupi_g15842(csa_tree_add_7_25_groupi_n_5226 ,csa_tree_add_7_25_groupi_n_5227);
  not csa_tree_add_7_25_groupi_g15843(csa_tree_add_7_25_groupi_n_5224 ,csa_tree_add_7_25_groupi_n_5225);
  nor csa_tree_add_7_25_groupi_g15844(csa_tree_add_7_25_groupi_n_5223 ,csa_tree_add_7_25_groupi_n_339 ,csa_tree_add_7_25_groupi_n_2190);
  nor csa_tree_add_7_25_groupi_g15845(csa_tree_add_7_25_groupi_n_5222 ,csa_tree_add_7_25_groupi_n_2118 ,csa_tree_add_7_25_groupi_n_132);
  xnor csa_tree_add_7_25_groupi_g15846(csa_tree_add_7_25_groupi_n_5221 ,csa_tree_add_7_25_groupi_n_4937 ,csa_tree_add_7_25_groupi_n_5125);
  xnor csa_tree_add_7_25_groupi_g15847(csa_tree_add_7_25_groupi_n_5220 ,csa_tree_add_7_25_groupi_n_4933 ,csa_tree_add_7_25_groupi_n_5126);
  xnor csa_tree_add_7_25_groupi_g15848(csa_tree_add_7_25_groupi_n_5219 ,csa_tree_add_7_25_groupi_n_4930 ,csa_tree_add_7_25_groupi_n_5118);
  xnor csa_tree_add_7_25_groupi_g15849(csa_tree_add_7_25_groupi_n_5218 ,csa_tree_add_7_25_groupi_n_1104 ,csa_tree_add_7_25_groupi_n_1108);
  xnor csa_tree_add_7_25_groupi_g15850(csa_tree_add_7_25_groupi_n_5217 ,csa_tree_add_7_25_groupi_n_4932 ,csa_tree_add_7_25_groupi_n_5123);
  xnor csa_tree_add_7_25_groupi_g15851(csa_tree_add_7_25_groupi_n_5216 ,csa_tree_add_7_25_groupi_n_4934 ,csa_tree_add_7_25_groupi_n_5124);
  xnor csa_tree_add_7_25_groupi_g15852(csa_tree_add_7_25_groupi_n_5215 ,csa_tree_add_7_25_groupi_n_4931 ,csa_tree_add_7_25_groupi_n_5121);
  xnor csa_tree_add_7_25_groupi_g15853(csa_tree_add_7_25_groupi_n_5214 ,csa_tree_add_7_25_groupi_n_4938 ,csa_tree_add_7_25_groupi_n_5122);
  xnor csa_tree_add_7_25_groupi_g15854(csa_tree_add_7_25_groupi_n_5213 ,csa_tree_add_7_25_groupi_n_4935 ,csa_tree_add_7_25_groupi_n_5127);
  xnor csa_tree_add_7_25_groupi_g15855(csa_tree_add_7_25_groupi_n_5247 ,csa_tree_add_7_25_groupi_n_5138 ,in3[5]);
  xnor csa_tree_add_7_25_groupi_g15856(csa_tree_add_7_25_groupi_n_5246 ,csa_tree_add_7_25_groupi_n_5141 ,in3[8]);
  xnor csa_tree_add_7_25_groupi_g15857(csa_tree_add_7_25_groupi_n_5245 ,csa_tree_add_7_25_groupi_n_5140 ,in3[11]);
  xnor csa_tree_add_7_25_groupi_g15858(csa_tree_add_7_25_groupi_n_5244 ,csa_tree_add_7_25_groupi_n_5145 ,in3[14]);
  xnor csa_tree_add_7_25_groupi_g15859(csa_tree_add_7_25_groupi_n_5243 ,csa_tree_add_7_25_groupi_n_5147 ,in3[2]);
  xnor csa_tree_add_7_25_groupi_g15860(csa_tree_add_7_25_groupi_n_5242 ,csa_tree_add_7_25_groupi_n_5143 ,in3[17]);
  xnor csa_tree_add_7_25_groupi_g15861(csa_tree_add_7_25_groupi_n_5241 ,csa_tree_add_7_25_groupi_n_5144 ,in3[20]);
  xnor csa_tree_add_7_25_groupi_g15862(csa_tree_add_7_25_groupi_n_5240 ,csa_tree_add_7_25_groupi_n_5146 ,in3[23]);
  xnor csa_tree_add_7_25_groupi_g15863(csa_tree_add_7_25_groupi_n_5239 ,csa_tree_add_7_25_groupi_n_5142 ,in3[26]);
  xnor csa_tree_add_7_25_groupi_g15864(csa_tree_add_7_25_groupi_n_5238 ,csa_tree_add_7_25_groupi_n_5139 ,in3[29]);
  xnor csa_tree_add_7_25_groupi_g15865(csa_tree_add_7_25_groupi_n_5237 ,csa_tree_add_7_25_groupi_n_5133 ,csa_tree_add_7_25_groupi_n_5036);
  xnor csa_tree_add_7_25_groupi_g15866(csa_tree_add_7_25_groupi_n_5236 ,csa_tree_add_7_25_groupi_n_5132 ,csa_tree_add_7_25_groupi_n_4950);
  xnor csa_tree_add_7_25_groupi_g15867(csa_tree_add_7_25_groupi_n_5235 ,csa_tree_add_7_25_groupi_n_5137 ,csa_tree_add_7_25_groupi_n_4949);
  xnor csa_tree_add_7_25_groupi_g15868(csa_tree_add_7_25_groupi_n_5234 ,csa_tree_add_7_25_groupi_n_5129 ,csa_tree_add_7_25_groupi_n_4946);
  xnor csa_tree_add_7_25_groupi_g15869(csa_tree_add_7_25_groupi_n_5233 ,csa_tree_add_7_25_groupi_n_5130 ,csa_tree_add_7_25_groupi_n_4941);
  xnor csa_tree_add_7_25_groupi_g15870(csa_tree_add_7_25_groupi_n_5232 ,csa_tree_add_7_25_groupi_n_4936 ,csa_tree_add_7_25_groupi_n_5111);
  xnor csa_tree_add_7_25_groupi_g15871(csa_tree_add_7_25_groupi_n_5231 ,csa_tree_add_7_25_groupi_n_5131 ,csa_tree_add_7_25_groupi_n_4945);
  xnor csa_tree_add_7_25_groupi_g15872(csa_tree_add_7_25_groupi_n_5230 ,csa_tree_add_7_25_groupi_n_5134 ,csa_tree_add_7_25_groupi_n_4944);
  xnor csa_tree_add_7_25_groupi_g15873(csa_tree_add_7_25_groupi_n_5229 ,csa_tree_add_7_25_groupi_n_5135 ,csa_tree_add_7_25_groupi_n_4943);
  xnor csa_tree_add_7_25_groupi_g15874(csa_tree_add_7_25_groupi_n_5228 ,csa_tree_add_7_25_groupi_n_5128 ,csa_tree_add_7_25_groupi_n_4942);
  xnor csa_tree_add_7_25_groupi_g15875(csa_tree_add_7_25_groupi_n_5227 ,csa_tree_add_7_25_groupi_n_5078 ,csa_tree_add_7_25_groupi_n_5110);
  xnor csa_tree_add_7_25_groupi_g15876(csa_tree_add_7_25_groupi_n_5225 ,csa_tree_add_7_25_groupi_n_5136 ,csa_tree_add_7_25_groupi_n_0);
  not csa_tree_add_7_25_groupi_g15877(csa_tree_add_7_25_groupi_n_5209 ,csa_tree_add_7_25_groupi_n_5210);
  or csa_tree_add_7_25_groupi_g15878(csa_tree_add_7_25_groupi_n_5208 ,csa_tree_add_7_25_groupi_n_3148 ,csa_tree_add_7_25_groupi_n_5117);
  and csa_tree_add_7_25_groupi_g15879(csa_tree_add_7_25_groupi_n_5207 ,csa_tree_add_7_25_groupi_n_5128 ,csa_tree_add_7_25_groupi_n_4925);
  and csa_tree_add_7_25_groupi_g15880(csa_tree_add_7_25_groupi_n_5206 ,csa_tree_add_7_25_groupi_n_5133 ,csa_tree_add_7_25_groupi_n_5021);
  and csa_tree_add_7_25_groupi_g15881(csa_tree_add_7_25_groupi_n_5205 ,csa_tree_add_7_25_groupi_n_5136 ,csa_tree_add_7_25_groupi_n_4814);
  and csa_tree_add_7_25_groupi_g15882(csa_tree_add_7_25_groupi_n_5204 ,csa_tree_add_7_25_groupi_n_5135 ,csa_tree_add_7_25_groupi_n_4920);
  or csa_tree_add_7_25_groupi_g15883(csa_tree_add_7_25_groupi_n_5203 ,csa_tree_add_7_25_groupi_n_3628 ,csa_tree_add_7_25_groupi_n_5152);
  and csa_tree_add_7_25_groupi_g15884(csa_tree_add_7_25_groupi_n_5202 ,csa_tree_add_7_25_groupi_n_5132 ,csa_tree_add_7_25_groupi_n_4914);
  and csa_tree_add_7_25_groupi_g15885(csa_tree_add_7_25_groupi_n_5201 ,csa_tree_add_7_25_groupi_n_5137 ,csa_tree_add_7_25_groupi_n_4915);
  and csa_tree_add_7_25_groupi_g15886(csa_tree_add_7_25_groupi_n_5200 ,csa_tree_add_7_25_groupi_n_5134 ,csa_tree_add_7_25_groupi_n_4918);
  and csa_tree_add_7_25_groupi_g15887(csa_tree_add_7_25_groupi_n_5199 ,csa_tree_add_7_25_groupi_n_5131 ,csa_tree_add_7_25_groupi_n_4923);
  and csa_tree_add_7_25_groupi_g15888(csa_tree_add_7_25_groupi_n_5198 ,csa_tree_add_7_25_groupi_n_5129 ,csa_tree_add_7_25_groupi_n_4927);
  and csa_tree_add_7_25_groupi_g15889(csa_tree_add_7_25_groupi_n_5197 ,csa_tree_add_7_25_groupi_n_4935 ,csa_tree_add_7_25_groupi_n_5127);
  or csa_tree_add_7_25_groupi_g15890(csa_tree_add_7_25_groupi_n_5196 ,csa_tree_add_7_25_groupi_n_4935 ,csa_tree_add_7_25_groupi_n_5127);
  and csa_tree_add_7_25_groupi_g15891(csa_tree_add_7_25_groupi_n_5195 ,csa_tree_add_7_25_groupi_n_4937 ,csa_tree_add_7_25_groupi_n_5125);
  or csa_tree_add_7_25_groupi_g15892(csa_tree_add_7_25_groupi_n_5194 ,csa_tree_add_7_25_groupi_n_4937 ,csa_tree_add_7_25_groupi_n_5125);
  or csa_tree_add_7_25_groupi_g15893(csa_tree_add_7_25_groupi_n_5193 ,csa_tree_add_7_25_groupi_n_4930 ,csa_tree_add_7_25_groupi_n_5118);
  and csa_tree_add_7_25_groupi_g15894(csa_tree_add_7_25_groupi_n_5192 ,csa_tree_add_7_25_groupi_n_4933 ,csa_tree_add_7_25_groupi_n_5126);
  or csa_tree_add_7_25_groupi_g15895(csa_tree_add_7_25_groupi_n_5191 ,csa_tree_add_7_25_groupi_n_4933 ,csa_tree_add_7_25_groupi_n_5126);
  and csa_tree_add_7_25_groupi_g15896(csa_tree_add_7_25_groupi_n_5190 ,csa_tree_add_7_25_groupi_n_5130 ,csa_tree_add_7_25_groupi_n_4886);
  and csa_tree_add_7_25_groupi_g15897(csa_tree_add_7_25_groupi_n_5189 ,csa_tree_add_7_25_groupi_n_4930 ,csa_tree_add_7_25_groupi_n_5118);
  and csa_tree_add_7_25_groupi_g15898(csa_tree_add_7_25_groupi_n_5212 ,csa_tree_add_7_25_groupi_n_2453 ,csa_tree_add_7_25_groupi_n_5149);
  or csa_tree_add_7_25_groupi_g15899(csa_tree_add_7_25_groupi_n_5211 ,csa_tree_add_7_25_groupi_n_5020 ,csa_tree_add_7_25_groupi_n_5148);
  or csa_tree_add_7_25_groupi_g15900(csa_tree_add_7_25_groupi_n_5210 ,csa_tree_add_7_25_groupi_n_5096 ,csa_tree_add_7_25_groupi_n_5150);
  or csa_tree_add_7_25_groupi_g15901(csa_tree_add_7_25_groupi_n_5187 ,csa_tree_add_7_25_groupi_n_4932 ,csa_tree_add_7_25_groupi_n_5123);
  or csa_tree_add_7_25_groupi_g15902(csa_tree_add_7_25_groupi_n_5186 ,csa_tree_add_7_25_groupi_n_3117 ,csa_tree_add_7_25_groupi_n_5114);
  or csa_tree_add_7_25_groupi_g15903(csa_tree_add_7_25_groupi_n_5185 ,csa_tree_add_7_25_groupi_n_3097 ,csa_tree_add_7_25_groupi_n_5113);
  or csa_tree_add_7_25_groupi_g15904(csa_tree_add_7_25_groupi_n_5184 ,csa_tree_add_7_25_groupi_n_2995 ,csa_tree_add_7_25_groupi_n_5154);
  or csa_tree_add_7_25_groupi_g15905(csa_tree_add_7_25_groupi_n_5183 ,in3[11] ,csa_tree_add_7_25_groupi_n_1096);
  and csa_tree_add_7_25_groupi_g15906(csa_tree_add_7_25_groupi_n_5182 ,in3[11] ,csa_tree_add_7_25_groupi_n_1108);
  or csa_tree_add_7_25_groupi_g15907(csa_tree_add_7_25_groupi_n_5181 ,csa_tree_add_7_25_groupi_n_3548 ,csa_tree_add_7_25_groupi_n_5155);
  or csa_tree_add_7_25_groupi_g15908(csa_tree_add_7_25_groupi_n_5180 ,csa_tree_add_7_25_groupi_n_3633 ,csa_tree_add_7_25_groupi_n_5112);
  nor csa_tree_add_7_25_groupi_g15909(csa_tree_add_7_25_groupi_n_5179 ,csa_tree_add_7_25_groupi_n_3030 ,csa_tree_add_7_25_groupi_n_5151);
  and csa_tree_add_7_25_groupi_g15910(csa_tree_add_7_25_groupi_n_5178 ,csa_tree_add_7_25_groupi_n_4938 ,csa_tree_add_7_25_groupi_n_5122);
  and csa_tree_add_7_25_groupi_g15911(csa_tree_add_7_25_groupi_n_5177 ,csa_tree_add_7_25_groupi_n_4934 ,csa_tree_add_7_25_groupi_n_5124);
  or csa_tree_add_7_25_groupi_g15912(csa_tree_add_7_25_groupi_n_5176 ,csa_tree_add_7_25_groupi_n_3113 ,csa_tree_add_7_25_groupi_n_5115);
  or csa_tree_add_7_25_groupi_g15913(csa_tree_add_7_25_groupi_n_5175 ,csa_tree_add_7_25_groupi_n_4934 ,csa_tree_add_7_25_groupi_n_5124);
  and csa_tree_add_7_25_groupi_g15914(csa_tree_add_7_25_groupi_n_5174 ,csa_tree_add_7_25_groupi_n_4932 ,csa_tree_add_7_25_groupi_n_5123);
  or csa_tree_add_7_25_groupi_g15915(csa_tree_add_7_25_groupi_n_5173 ,csa_tree_add_7_25_groupi_n_4938 ,csa_tree_add_7_25_groupi_n_5122);
  and csa_tree_add_7_25_groupi_g15916(csa_tree_add_7_25_groupi_n_5172 ,csa_tree_add_7_25_groupi_n_4931 ,csa_tree_add_7_25_groupi_n_5121);
  or csa_tree_add_7_25_groupi_g15917(csa_tree_add_7_25_groupi_n_5171 ,csa_tree_add_7_25_groupi_n_4931 ,csa_tree_add_7_25_groupi_n_5121);
  or csa_tree_add_7_25_groupi_g15918(csa_tree_add_7_25_groupi_n_5170 ,csa_tree_add_7_25_groupi_n_2974 ,csa_tree_add_7_25_groupi_n_5153);
  nor csa_tree_add_7_25_groupi_g15919(csa_tree_add_7_25_groupi_n_5169 ,csa_tree_add_7_25_groupi_n_5074 ,csa_tree_add_7_25_groupi_n_2345);
  or csa_tree_add_7_25_groupi_g15920(csa_tree_add_7_25_groupi_n_5168 ,csa_tree_add_7_25_groupi_n_5075 ,csa_tree_add_7_25_groupi_n_1096);
  xnor csa_tree_add_7_25_groupi_g15921(out2[4] ,csa_tree_add_7_25_groupi_n_5107 ,csa_tree_add_7_25_groupi_n_5034);
  or csa_tree_add_7_25_groupi_g15922(csa_tree_add_7_25_groupi_n_5166 ,csa_tree_add_7_25_groupi_n_3137 ,csa_tree_add_7_25_groupi_n_5116);
  xnor csa_tree_add_7_25_groupi_g15923(csa_tree_add_7_25_groupi_n_5188 ,csa_tree_add_7_25_groupi_n_5108 ,csa_tree_add_7_25_groupi_n_2578);
  nor csa_tree_add_7_25_groupi_g15925(csa_tree_add_7_25_groupi_n_5155 ,csa_tree_add_7_25_groupi_n_279 ,csa_tree_add_7_25_groupi_n_2018);
  nor csa_tree_add_7_25_groupi_g15926(csa_tree_add_7_25_groupi_n_5154 ,csa_tree_add_7_25_groupi_n_362 ,csa_tree_add_7_25_groupi_n_1830);
  nor csa_tree_add_7_25_groupi_g15927(csa_tree_add_7_25_groupi_n_5153 ,csa_tree_add_7_25_groupi_n_2174 ,csa_tree_add_7_25_groupi_n_1831);
  nor csa_tree_add_7_25_groupi_g15928(csa_tree_add_7_25_groupi_n_5152 ,csa_tree_add_7_25_groupi_n_1879 ,csa_tree_add_7_25_groupi_n_141);
  nor csa_tree_add_7_25_groupi_g15929(csa_tree_add_7_25_groupi_n_5151 ,csa_tree_add_7_25_groupi_n_638 ,csa_tree_add_7_25_groupi_n_280);
  and csa_tree_add_7_25_groupi_g15930(csa_tree_add_7_25_groupi_n_5150 ,csa_tree_add_7_25_groupi_n_5078 ,csa_tree_add_7_25_groupi_n_5095);
  or csa_tree_add_7_25_groupi_g15931(csa_tree_add_7_25_groupi_n_5149 ,csa_tree_add_7_25_groupi_n_2481 ,csa_tree_add_7_25_groupi_n_5108);
  and csa_tree_add_7_25_groupi_g15932(csa_tree_add_7_25_groupi_n_5148 ,csa_tree_add_7_25_groupi_n_5025 ,csa_tree_add_7_25_groupi_n_5107);
  nor csa_tree_add_7_25_groupi_g15933(csa_tree_add_7_25_groupi_n_5147 ,csa_tree_add_7_25_groupi_n_3488 ,csa_tree_add_7_25_groupi_n_5080);
  nor csa_tree_add_7_25_groupi_g15934(csa_tree_add_7_25_groupi_n_5146 ,csa_tree_add_7_25_groupi_n_3809 ,csa_tree_add_7_25_groupi_n_5088);
  nor csa_tree_add_7_25_groupi_g15935(csa_tree_add_7_25_groupi_n_5145 ,csa_tree_add_7_25_groupi_n_3990 ,csa_tree_add_7_25_groupi_n_5089);
  nor csa_tree_add_7_25_groupi_g15936(csa_tree_add_7_25_groupi_n_5144 ,csa_tree_add_7_25_groupi_n_3887 ,csa_tree_add_7_25_groupi_n_5087);
  nor csa_tree_add_7_25_groupi_g15937(csa_tree_add_7_25_groupi_n_5143 ,csa_tree_add_7_25_groupi_n_3822 ,csa_tree_add_7_25_groupi_n_5086);
  nor csa_tree_add_7_25_groupi_g15938(csa_tree_add_7_25_groupi_n_5142 ,csa_tree_add_7_25_groupi_n_4038 ,csa_tree_add_7_25_groupi_n_5100);
  nor csa_tree_add_7_25_groupi_g15939(csa_tree_add_7_25_groupi_n_5141 ,csa_tree_add_7_25_groupi_n_4029 ,csa_tree_add_7_25_groupi_n_5090);
  nor csa_tree_add_7_25_groupi_g15940(csa_tree_add_7_25_groupi_n_5140 ,csa_tree_add_7_25_groupi_n_4068 ,csa_tree_add_7_25_groupi_n_5091);
  nor csa_tree_add_7_25_groupi_g15941(csa_tree_add_7_25_groupi_n_5139 ,csa_tree_add_7_25_groupi_n_3886 ,csa_tree_add_7_25_groupi_n_5102);
  nor csa_tree_add_7_25_groupi_g15942(csa_tree_add_7_25_groupi_n_5138 ,csa_tree_add_7_25_groupi_n_4080 ,csa_tree_add_7_25_groupi_n_5085);
  or csa_tree_add_7_25_groupi_g15943(csa_tree_add_7_25_groupi_n_5165 ,csa_tree_add_7_25_groupi_n_4787 ,csa_tree_add_7_25_groupi_n_5083);
  or csa_tree_add_7_25_groupi_g15944(csa_tree_add_7_25_groupi_n_5164 ,csa_tree_add_7_25_groupi_n_4782 ,csa_tree_add_7_25_groupi_n_5082);
  or csa_tree_add_7_25_groupi_g15945(csa_tree_add_7_25_groupi_n_5163 ,csa_tree_add_7_25_groupi_n_4778 ,csa_tree_add_7_25_groupi_n_5081);
  or csa_tree_add_7_25_groupi_g15946(csa_tree_add_7_25_groupi_n_5162 ,csa_tree_add_7_25_groupi_n_4811 ,csa_tree_add_7_25_groupi_n_5101);
  or csa_tree_add_7_25_groupi_g15947(csa_tree_add_7_25_groupi_n_5161 ,csa_tree_add_7_25_groupi_n_4808 ,csa_tree_add_7_25_groupi_n_5106);
  or csa_tree_add_7_25_groupi_g15948(csa_tree_add_7_25_groupi_n_5160 ,csa_tree_add_7_25_groupi_n_4777 ,csa_tree_add_7_25_groupi_n_5092);
  or csa_tree_add_7_25_groupi_g15949(csa_tree_add_7_25_groupi_n_5159 ,csa_tree_add_7_25_groupi_n_4982 ,csa_tree_add_7_25_groupi_n_5094);
  or csa_tree_add_7_25_groupi_g15950(csa_tree_add_7_25_groupi_n_5158 ,csa_tree_add_7_25_groupi_n_4813 ,csa_tree_add_7_25_groupi_n_5103);
  or csa_tree_add_7_25_groupi_g15951(csa_tree_add_7_25_groupi_n_5157 ,csa_tree_add_7_25_groupi_n_4802 ,csa_tree_add_7_25_groupi_n_5105);
  and csa_tree_add_7_25_groupi_g15952(csa_tree_add_7_25_groupi_n_5156 ,csa_tree_add_7_25_groupi_n_3899 ,csa_tree_add_7_25_groupi_n_5084);
  not csa_tree_add_7_25_groupi_g15953(csa_tree_add_7_25_groupi_n_5119 ,csa_tree_add_7_25_groupi_n_5120);
  nor csa_tree_add_7_25_groupi_g15954(csa_tree_add_7_25_groupi_n_5117 ,csa_tree_add_7_25_groupi_n_302 ,csa_tree_add_7_25_groupi_n_2073);
  nor csa_tree_add_7_25_groupi_g15955(csa_tree_add_7_25_groupi_n_5116 ,csa_tree_add_7_25_groupi_n_303 ,csa_tree_add_7_25_groupi_n_2132);
  nor csa_tree_add_7_25_groupi_g15956(csa_tree_add_7_25_groupi_n_5115 ,csa_tree_add_7_25_groupi_n_303 ,csa_tree_add_7_25_groupi_n_2096);
  nor csa_tree_add_7_25_groupi_g15957(csa_tree_add_7_25_groupi_n_5114 ,csa_tree_add_7_25_groupi_n_2117 ,csa_tree_add_7_25_groupi_n_1830);
  nor csa_tree_add_7_25_groupi_g15958(csa_tree_add_7_25_groupi_n_5113 ,csa_tree_add_7_25_groupi_n_280 ,csa_tree_add_7_25_groupi_n_2189);
  nor csa_tree_add_7_25_groupi_g15959(csa_tree_add_7_25_groupi_n_5112 ,csa_tree_add_7_25_groupi_n_2034 ,csa_tree_add_7_25_groupi_n_141);
  xnor csa_tree_add_7_25_groupi_g15960(csa_tree_add_7_25_groupi_n_5111 ,csa_tree_add_7_25_groupi_n_5047 ,csa_tree_add_7_25_groupi_n_4851);
  xnor csa_tree_add_7_25_groupi_g15961(csa_tree_add_7_25_groupi_n_5110 ,csa_tree_add_7_25_groupi_n_5043 ,csa_tree_add_7_25_groupi_n_4845);
  xnor csa_tree_add_7_25_groupi_g15962(csa_tree_add_7_25_groupi_n_5109 ,csa_tree_add_7_25_groupi_n_4988 ,csa_tree_add_7_25_groupi_n_5041);
  xnor csa_tree_add_7_25_groupi_g15964(csa_tree_add_7_25_groupi_n_5137 ,csa_tree_add_7_25_groupi_n_5058 ,in3[2]);
  xnor csa_tree_add_7_25_groupi_g15965(csa_tree_add_7_25_groupi_n_5136 ,csa_tree_add_7_25_groupi_n_5056 ,in3[29]);
  xnor csa_tree_add_7_25_groupi_g15966(csa_tree_add_7_25_groupi_n_5135 ,csa_tree_add_7_25_groupi_n_5053 ,in3[17]);
  xnor csa_tree_add_7_25_groupi_g15967(csa_tree_add_7_25_groupi_n_5134 ,csa_tree_add_7_25_groupi_n_5059 ,in3[14]);
  xnor csa_tree_add_7_25_groupi_g15968(csa_tree_add_7_25_groupi_n_5133 ,csa_tree_add_7_25_groupi_n_5055 ,in3[26]);
  xnor csa_tree_add_7_25_groupi_g15969(csa_tree_add_7_25_groupi_n_5132 ,csa_tree_add_7_25_groupi_n_5060 ,in3[5]);
  xnor csa_tree_add_7_25_groupi_g15970(csa_tree_add_7_25_groupi_n_5131 ,csa_tree_add_7_25_groupi_n_5061 ,in3[11]);
  xnor csa_tree_add_7_25_groupi_g15971(csa_tree_add_7_25_groupi_n_5130 ,csa_tree_add_7_25_groupi_n_5054 ,in3[23]);
  xnor csa_tree_add_7_25_groupi_g15972(csa_tree_add_7_25_groupi_n_5129 ,csa_tree_add_7_25_groupi_n_5062 ,in3[8]);
  xnor csa_tree_add_7_25_groupi_g15973(csa_tree_add_7_25_groupi_n_5128 ,csa_tree_add_7_25_groupi_n_5057 ,in3[20]);
  xnor csa_tree_add_7_25_groupi_g15974(csa_tree_add_7_25_groupi_n_5127 ,csa_tree_add_7_25_groupi_n_5052 ,csa_tree_add_7_25_groupi_n_4837);
  xnor csa_tree_add_7_25_groupi_g15975(csa_tree_add_7_25_groupi_n_5126 ,csa_tree_add_7_25_groupi_n_5044 ,csa_tree_add_7_25_groupi_n_4835);
  xnor csa_tree_add_7_25_groupi_g15976(csa_tree_add_7_25_groupi_n_5125 ,csa_tree_add_7_25_groupi_n_5046 ,csa_tree_add_7_25_groupi_n_4836);
  xnor csa_tree_add_7_25_groupi_g15977(csa_tree_add_7_25_groupi_n_5124 ,csa_tree_add_7_25_groupi_n_5049 ,csa_tree_add_7_25_groupi_n_4832);
  xnor csa_tree_add_7_25_groupi_g15978(csa_tree_add_7_25_groupi_n_5123 ,csa_tree_add_7_25_groupi_n_5050 ,csa_tree_add_7_25_groupi_n_4833);
  xnor csa_tree_add_7_25_groupi_g15979(csa_tree_add_7_25_groupi_n_5122 ,csa_tree_add_7_25_groupi_n_5051 ,csa_tree_add_7_25_groupi_n_4829);
  xnor csa_tree_add_7_25_groupi_g15980(csa_tree_add_7_25_groupi_n_5121 ,csa_tree_add_7_25_groupi_n_5048 ,csa_tree_add_7_25_groupi_n_4830);
  xnor csa_tree_add_7_25_groupi_g15981(csa_tree_add_7_25_groupi_n_5120 ,csa_tree_add_7_25_groupi_n_5028 ,csa_tree_add_7_25_groupi_n_4883);
  xnor csa_tree_add_7_25_groupi_g15982(csa_tree_add_7_25_groupi_n_5118 ,csa_tree_add_7_25_groupi_n_5045 ,csa_tree_add_7_25_groupi_n_4834);
  and csa_tree_add_7_25_groupi_g15983(csa_tree_add_7_25_groupi_n_5106 ,csa_tree_add_7_25_groupi_n_5052 ,csa_tree_add_7_25_groupi_n_4809);
  and csa_tree_add_7_25_groupi_g15984(csa_tree_add_7_25_groupi_n_5105 ,csa_tree_add_7_25_groupi_n_5045 ,csa_tree_add_7_25_groupi_n_4816);
  or csa_tree_add_7_25_groupi_g15985(csa_tree_add_7_25_groupi_n_5104 ,csa_tree_add_7_25_groupi_n_1104 ,csa_tree_add_7_25_groupi_n_5076);
  and csa_tree_add_7_25_groupi_g15986(csa_tree_add_7_25_groupi_n_5103 ,csa_tree_add_7_25_groupi_n_5044 ,csa_tree_add_7_25_groupi_n_4812);
  or csa_tree_add_7_25_groupi_g15987(csa_tree_add_7_25_groupi_n_5102 ,csa_tree_add_7_25_groupi_n_3629 ,csa_tree_add_7_25_groupi_n_5067);
  and csa_tree_add_7_25_groupi_g15988(csa_tree_add_7_25_groupi_n_5101 ,csa_tree_add_7_25_groupi_n_5046 ,csa_tree_add_7_25_groupi_n_4810);
  or csa_tree_add_7_25_groupi_g15989(csa_tree_add_7_25_groupi_n_5100 ,csa_tree_add_7_25_groupi_n_3245 ,csa_tree_add_7_25_groupi_n_5065);
  nor csa_tree_add_7_25_groupi_g15990(csa_tree_add_7_25_groupi_n_5099 ,csa_tree_add_7_25_groupi_n_5075 ,csa_tree_add_7_25_groupi_n_5077);
  or csa_tree_add_7_25_groupi_g15991(csa_tree_add_7_25_groupi_n_5098 ,csa_tree_add_7_25_groupi_n_4988 ,csa_tree_add_7_25_groupi_n_5040);
  nor csa_tree_add_7_25_groupi_g15992(csa_tree_add_7_25_groupi_n_5097 ,csa_tree_add_7_25_groupi_n_4987 ,csa_tree_add_7_25_groupi_n_5041);
  nor csa_tree_add_7_25_groupi_g15993(csa_tree_add_7_25_groupi_n_5096 ,csa_tree_add_7_25_groupi_n_5042 ,csa_tree_add_7_25_groupi_n_4845);
  or csa_tree_add_7_25_groupi_g15994(csa_tree_add_7_25_groupi_n_5095 ,csa_tree_add_7_25_groupi_n_5043 ,csa_tree_add_7_25_groupi_n_4844);
  and csa_tree_add_7_25_groupi_g15995(csa_tree_add_7_25_groupi_n_5094 ,csa_tree_add_7_25_groupi_n_5047 ,csa_tree_add_7_25_groupi_n_4981);
  and csa_tree_add_7_25_groupi_g15996(csa_tree_add_7_25_groupi_n_5108 ,csa_tree_add_7_25_groupi_n_2443 ,csa_tree_add_7_25_groupi_n_5070);
  or csa_tree_add_7_25_groupi_g15997(csa_tree_add_7_25_groupi_n_5107 ,csa_tree_add_7_25_groupi_n_4928 ,csa_tree_add_7_25_groupi_n_5071);
  and csa_tree_add_7_25_groupi_g15998(csa_tree_add_7_25_groupi_n_5092 ,csa_tree_add_7_25_groupi_n_5048 ,csa_tree_add_7_25_groupi_n_4780);
  or csa_tree_add_7_25_groupi_g15999(csa_tree_add_7_25_groupi_n_5091 ,csa_tree_add_7_25_groupi_n_3118 ,csa_tree_add_7_25_groupi_n_5039);
  or csa_tree_add_7_25_groupi_g16000(csa_tree_add_7_25_groupi_n_5090 ,csa_tree_add_7_25_groupi_n_3116 ,csa_tree_add_7_25_groupi_n_5068);
  or csa_tree_add_7_25_groupi_g16001(csa_tree_add_7_25_groupi_n_5089 ,csa_tree_add_7_25_groupi_n_3114 ,csa_tree_add_7_25_groupi_n_5038);
  or csa_tree_add_7_25_groupi_g16002(csa_tree_add_7_25_groupi_n_5088 ,csa_tree_add_7_25_groupi_n_3647 ,csa_tree_add_7_25_groupi_n_5064);
  or csa_tree_add_7_25_groupi_g16003(csa_tree_add_7_25_groupi_n_5087 ,csa_tree_add_7_25_groupi_n_3569 ,csa_tree_add_7_25_groupi_n_5063);
  or csa_tree_add_7_25_groupi_g16004(csa_tree_add_7_25_groupi_n_5086 ,csa_tree_add_7_25_groupi_n_3632 ,csa_tree_add_7_25_groupi_n_5069);
  or csa_tree_add_7_25_groupi_g16005(csa_tree_add_7_25_groupi_n_5085 ,csa_tree_add_7_25_groupi_n_3138 ,csa_tree_add_7_25_groupi_n_5072);
  nor csa_tree_add_7_25_groupi_g16006(csa_tree_add_7_25_groupi_n_5084 ,csa_tree_add_7_25_groupi_n_2978 ,csa_tree_add_7_25_groupi_n_5073);
  and csa_tree_add_7_25_groupi_g16007(csa_tree_add_7_25_groupi_n_5083 ,csa_tree_add_7_25_groupi_n_5049 ,csa_tree_add_7_25_groupi_n_4786);
  and csa_tree_add_7_25_groupi_g16008(csa_tree_add_7_25_groupi_n_5082 ,csa_tree_add_7_25_groupi_n_5050 ,csa_tree_add_7_25_groupi_n_4781);
  and csa_tree_add_7_25_groupi_g16009(csa_tree_add_7_25_groupi_n_5081 ,csa_tree_add_7_25_groupi_n_5051 ,csa_tree_add_7_25_groupi_n_4779);
  or csa_tree_add_7_25_groupi_g16010(csa_tree_add_7_25_groupi_n_5080 ,csa_tree_add_7_25_groupi_n_2985 ,csa_tree_add_7_25_groupi_n_5066);
  xnor csa_tree_add_7_25_groupi_g16011(out2[3] ,csa_tree_add_7_25_groupi_n_5008 ,csa_tree_add_7_25_groupi_n_4948);
  xnor csa_tree_add_7_25_groupi_g16012(csa_tree_add_7_25_groupi_n_5093 ,csa_tree_add_7_25_groupi_n_5026 ,csa_tree_add_7_25_groupi_n_2583);
  not csa_tree_add_7_25_groupi_g16013(csa_tree_add_7_25_groupi_n_5076 ,csa_tree_add_7_25_groupi_n_5077);
  not csa_tree_add_7_25_groupi_g16014(csa_tree_add_7_25_groupi_n_5075 ,csa_tree_add_7_25_groupi_n_5074);
  nor csa_tree_add_7_25_groupi_g16015(csa_tree_add_7_25_groupi_n_5073 ,csa_tree_add_7_25_groupi_n_549 ,csa_tree_add_7_25_groupi_n_283);
  nor csa_tree_add_7_25_groupi_g16016(csa_tree_add_7_25_groupi_n_5072 ,csa_tree_add_7_25_groupi_n_2130 ,csa_tree_add_7_25_groupi_n_1827);
  and csa_tree_add_7_25_groupi_g16017(csa_tree_add_7_25_groupi_n_5071 ,csa_tree_add_7_25_groupi_n_4919 ,csa_tree_add_7_25_groupi_n_5008);
  or csa_tree_add_7_25_groupi_g16018(csa_tree_add_7_25_groupi_n_5070 ,csa_tree_add_7_25_groupi_n_2422 ,csa_tree_add_7_25_groupi_n_5026);
  nor csa_tree_add_7_25_groupi_g16019(csa_tree_add_7_25_groupi_n_5069 ,csa_tree_add_7_25_groupi_n_2070 ,csa_tree_add_7_25_groupi_n_1828);
  nor csa_tree_add_7_25_groupi_g16020(csa_tree_add_7_25_groupi_n_5068 ,csa_tree_add_7_25_groupi_n_2115 ,csa_tree_add_7_25_groupi_n_187);
  nor csa_tree_add_7_25_groupi_g16021(csa_tree_add_7_25_groupi_n_5067 ,csa_tree_add_7_25_groupi_n_315 ,csa_tree_add_7_25_groupi_n_1322);
  nor csa_tree_add_7_25_groupi_g16022(csa_tree_add_7_25_groupi_n_5066 ,csa_tree_add_7_25_groupi_n_282 ,csa_tree_add_7_25_groupi_n_2172);
  nor csa_tree_add_7_25_groupi_g16023(csa_tree_add_7_25_groupi_n_5065 ,csa_tree_add_7_25_groupi_n_315 ,csa_tree_add_7_25_groupi_n_1309);
  nor csa_tree_add_7_25_groupi_g16024(csa_tree_add_7_25_groupi_n_5064 ,csa_tree_add_7_25_groupi_n_314 ,csa_tree_add_7_25_groupi_n_2019);
  nor csa_tree_add_7_25_groupi_g16025(csa_tree_add_7_25_groupi_n_5063 ,csa_tree_add_7_25_groupi_n_2039 ,csa_tree_add_7_25_groupi_n_1827);
  nor csa_tree_add_7_25_groupi_g16026(csa_tree_add_7_25_groupi_n_5062 ,csa_tree_add_7_25_groupi_n_4083 ,csa_tree_add_7_25_groupi_n_4996);
  nor csa_tree_add_7_25_groupi_g16027(csa_tree_add_7_25_groupi_n_5061 ,csa_tree_add_7_25_groupi_n_4022 ,csa_tree_add_7_25_groupi_n_5006);
  nor csa_tree_add_7_25_groupi_g16028(csa_tree_add_7_25_groupi_n_5060 ,csa_tree_add_7_25_groupi_n_4073 ,csa_tree_add_7_25_groupi_n_4999);
  nor csa_tree_add_7_25_groupi_g16029(csa_tree_add_7_25_groupi_n_5059 ,csa_tree_add_7_25_groupi_n_3989 ,csa_tree_add_7_25_groupi_n_4998);
  nor csa_tree_add_7_25_groupi_g16030(csa_tree_add_7_25_groupi_n_5058 ,csa_tree_add_7_25_groupi_n_3492 ,csa_tree_add_7_25_groupi_n_4990);
  nor csa_tree_add_7_25_groupi_g16031(csa_tree_add_7_25_groupi_n_5057 ,csa_tree_add_7_25_groupi_n_3808 ,csa_tree_add_7_25_groupi_n_4993);
  nor csa_tree_add_7_25_groupi_g16032(csa_tree_add_7_25_groupi_n_5056 ,csa_tree_add_7_25_groupi_n_3928 ,csa_tree_add_7_25_groupi_n_5001);
  nor csa_tree_add_7_25_groupi_g16033(csa_tree_add_7_25_groupi_n_5055 ,csa_tree_add_7_25_groupi_n_3925 ,csa_tree_add_7_25_groupi_n_4995);
  nor csa_tree_add_7_25_groupi_g16034(csa_tree_add_7_25_groupi_n_5054 ,csa_tree_add_7_25_groupi_n_3946 ,csa_tree_add_7_25_groupi_n_4994);
  nor csa_tree_add_7_25_groupi_g16035(csa_tree_add_7_25_groupi_n_5053 ,csa_tree_add_7_25_groupi_n_4085 ,csa_tree_add_7_25_groupi_n_5000);
  or csa_tree_add_7_25_groupi_g16036(csa_tree_add_7_25_groupi_n_5078 ,csa_tree_add_7_25_groupi_n_4557 ,csa_tree_add_7_25_groupi_n_5002);
  and csa_tree_add_7_25_groupi_g16037(csa_tree_add_7_25_groupi_n_5077 ,csa_tree_add_7_25_groupi_n_4894 ,csa_tree_add_7_25_groupi_n_5023);
  and csa_tree_add_7_25_groupi_g16038(csa_tree_add_7_25_groupi_n_5074 ,csa_tree_add_7_25_groupi_n_3923 ,csa_tree_add_7_25_groupi_n_4991);
  not csa_tree_add_7_25_groupi_g16039(csa_tree_add_7_25_groupi_n_5042 ,csa_tree_add_7_25_groupi_n_5043);
  not csa_tree_add_7_25_groupi_g16040(csa_tree_add_7_25_groupi_n_5040 ,csa_tree_add_7_25_groupi_n_5041);
  nor csa_tree_add_7_25_groupi_g16041(csa_tree_add_7_25_groupi_n_5039 ,csa_tree_add_7_25_groupi_n_283 ,csa_tree_add_7_25_groupi_n_2094);
  nor csa_tree_add_7_25_groupi_g16042(csa_tree_add_7_25_groupi_n_5038 ,csa_tree_add_7_25_groupi_n_2148 ,csa_tree_add_7_25_groupi_n_187);
  xnor csa_tree_add_7_25_groupi_g16043(csa_tree_add_7_25_groupi_n_5037 ,csa_tree_add_7_25_groupi_n_4954 ,csa_tree_add_7_25_groupi_n_4907);
  xnor csa_tree_add_7_25_groupi_g16044(csa_tree_add_7_25_groupi_n_5036 ,csa_tree_add_7_25_groupi_n_4884 ,csa_tree_add_7_25_groupi_n_4957);
  xnor csa_tree_add_7_25_groupi_g16045(csa_tree_add_7_25_groupi_n_5035 ,csa_tree_add_7_25_groupi_n_4962 ,csa_tree_add_7_25_groupi_n_4912);
  xnor csa_tree_add_7_25_groupi_g16046(csa_tree_add_7_25_groupi_n_5034 ,csa_tree_add_7_25_groupi_n_4960 ,csa_tree_add_7_25_groupi_n_4905);
  xnor csa_tree_add_7_25_groupi_g16047(csa_tree_add_7_25_groupi_n_5033 ,csa_tree_add_7_25_groupi_n_4963 ,csa_tree_add_7_25_groupi_n_4904);
  xnor csa_tree_add_7_25_groupi_g16048(csa_tree_add_7_25_groupi_n_5032 ,csa_tree_add_7_25_groupi_n_4961 ,csa_tree_add_7_25_groupi_n_4911);
  xnor csa_tree_add_7_25_groupi_g16049(csa_tree_add_7_25_groupi_n_5031 ,csa_tree_add_7_25_groupi_n_4959 ,csa_tree_add_7_25_groupi_n_4910);
  xnor csa_tree_add_7_25_groupi_g16050(csa_tree_add_7_25_groupi_n_5030 ,csa_tree_add_7_25_groupi_n_4958 ,csa_tree_add_7_25_groupi_n_4909);
  xnor csa_tree_add_7_25_groupi_g16051(csa_tree_add_7_25_groupi_n_5029 ,csa_tree_add_7_25_groupi_n_4956 ,csa_tree_add_7_25_groupi_n_4908);
  xnor csa_tree_add_7_25_groupi_g16052(csa_tree_add_7_25_groupi_n_5028 ,csa_tree_add_7_25_groupi_n_4989 ,in3[8]);
  xnor csa_tree_add_7_25_groupi_g16053(csa_tree_add_7_25_groupi_n_5027 ,csa_tree_add_7_25_groupi_n_4955 ,csa_tree_add_7_25_groupi_n_4906);
  xnor csa_tree_add_7_25_groupi_g16054(csa_tree_add_7_25_groupi_n_5052 ,csa_tree_add_7_25_groupi_n_4972 ,in3[14]);
  xnor csa_tree_add_7_25_groupi_g16055(csa_tree_add_7_25_groupi_n_5051 ,csa_tree_add_7_25_groupi_n_4970 ,in3[5]);
  xnor csa_tree_add_7_25_groupi_g16056(csa_tree_add_7_25_groupi_n_5050 ,csa_tree_add_7_25_groupi_n_4971 ,in3[8]);
  xnor csa_tree_add_7_25_groupi_g16057(csa_tree_add_7_25_groupi_n_5049 ,csa_tree_add_7_25_groupi_n_4973 ,in3[11]);
  xnor csa_tree_add_7_25_groupi_g16058(csa_tree_add_7_25_groupi_n_5048 ,csa_tree_add_7_25_groupi_n_4974 ,in3[2]);
  xnor csa_tree_add_7_25_groupi_g16059(csa_tree_add_7_25_groupi_n_5047 ,csa_tree_add_7_25_groupi_n_4967 ,in3[26]);
  xnor csa_tree_add_7_25_groupi_g16060(csa_tree_add_7_25_groupi_n_5046 ,csa_tree_add_7_25_groupi_n_4965 ,in3[17]);
  xnor csa_tree_add_7_25_groupi_g16061(csa_tree_add_7_25_groupi_n_5045 ,csa_tree_add_7_25_groupi_n_4968 ,in3[23]);
  xnor csa_tree_add_7_25_groupi_g16062(csa_tree_add_7_25_groupi_n_5044 ,csa_tree_add_7_25_groupi_n_4969 ,in3[20]);
  xnor csa_tree_add_7_25_groupi_g16063(csa_tree_add_7_25_groupi_n_5043 ,csa_tree_add_7_25_groupi_n_4966 ,in3[29]);
  xnor csa_tree_add_7_25_groupi_g16064(csa_tree_add_7_25_groupi_n_5041 ,csa_tree_add_7_25_groupi_n_4964 ,csa_tree_add_7_25_groupi_n_4616);
  or csa_tree_add_7_25_groupi_g16065(csa_tree_add_7_25_groupi_n_5025 ,csa_tree_add_7_25_groupi_n_4960 ,csa_tree_add_7_25_groupi_n_4905);
  and csa_tree_add_7_25_groupi_g16066(csa_tree_add_7_25_groupi_n_5024 ,csa_tree_add_7_25_groupi_n_4954 ,csa_tree_add_7_25_groupi_n_4907);
  or csa_tree_add_7_25_groupi_g16067(csa_tree_add_7_25_groupi_n_5023 ,csa_tree_add_7_25_groupi_n_4893 ,csa_tree_add_7_25_groupi_n_4989);
  and csa_tree_add_7_25_groupi_g16068(csa_tree_add_7_25_groupi_n_5022 ,csa_tree_add_7_25_groupi_n_4884 ,csa_tree_add_7_25_groupi_n_4957);
  or csa_tree_add_7_25_groupi_g16069(csa_tree_add_7_25_groupi_n_5021 ,csa_tree_add_7_25_groupi_n_4884 ,csa_tree_add_7_25_groupi_n_4957);
  and csa_tree_add_7_25_groupi_g16070(csa_tree_add_7_25_groupi_n_5020 ,csa_tree_add_7_25_groupi_n_4960 ,csa_tree_add_7_25_groupi_n_4905);
  and csa_tree_add_7_25_groupi_g16071(csa_tree_add_7_25_groupi_n_5019 ,csa_tree_add_7_25_groupi_n_4955 ,csa_tree_add_7_25_groupi_n_4906);
  or csa_tree_add_7_25_groupi_g16072(csa_tree_add_7_25_groupi_n_5018 ,csa_tree_add_7_25_groupi_n_4955 ,csa_tree_add_7_25_groupi_n_4906);
  or csa_tree_add_7_25_groupi_g16073(csa_tree_add_7_25_groupi_n_5017 ,csa_tree_add_7_25_groupi_n_4954 ,csa_tree_add_7_25_groupi_n_4907);
  and csa_tree_add_7_25_groupi_g16074(csa_tree_add_7_25_groupi_n_5016 ,csa_tree_add_7_25_groupi_n_4962 ,csa_tree_add_7_25_groupi_n_4912);
  or csa_tree_add_7_25_groupi_g16075(csa_tree_add_7_25_groupi_n_5015 ,csa_tree_add_7_25_groupi_n_4962 ,csa_tree_add_7_25_groupi_n_4912);
  and csa_tree_add_7_25_groupi_g16076(csa_tree_add_7_25_groupi_n_5014 ,csa_tree_add_7_25_groupi_n_4963 ,csa_tree_add_7_25_groupi_n_4904);
  or csa_tree_add_7_25_groupi_g16077(csa_tree_add_7_25_groupi_n_5013 ,csa_tree_add_7_25_groupi_n_4963 ,csa_tree_add_7_25_groupi_n_4904);
  and csa_tree_add_7_25_groupi_g16078(csa_tree_add_7_25_groupi_n_5012 ,csa_tree_add_7_25_groupi_n_4961 ,csa_tree_add_7_25_groupi_n_4911);
  or csa_tree_add_7_25_groupi_g16079(csa_tree_add_7_25_groupi_n_5011 ,csa_tree_add_7_25_groupi_n_4961 ,csa_tree_add_7_25_groupi_n_4911);
  and csa_tree_add_7_25_groupi_g16080(csa_tree_add_7_25_groupi_n_5010 ,csa_tree_add_7_25_groupi_n_4958 ,csa_tree_add_7_25_groupi_n_4909);
  or csa_tree_add_7_25_groupi_g16081(csa_tree_add_7_25_groupi_n_5009 ,csa_tree_add_7_25_groupi_n_4958 ,csa_tree_add_7_25_groupi_n_4909);
  and csa_tree_add_7_25_groupi_g16082(csa_tree_add_7_25_groupi_n_5026 ,csa_tree_add_7_25_groupi_n_2465 ,csa_tree_add_7_25_groupi_n_4985);
  or csa_tree_add_7_25_groupi_g16083(csa_tree_add_7_25_groupi_n_5006 ,csa_tree_add_7_25_groupi_n_3099 ,csa_tree_add_7_25_groupi_n_4952);
  or csa_tree_add_7_25_groupi_g16084(csa_tree_add_7_25_groupi_n_5005 ,csa_tree_add_7_25_groupi_n_4959 ,csa_tree_add_7_25_groupi_n_4910);
  and csa_tree_add_7_25_groupi_g16085(csa_tree_add_7_25_groupi_n_5004 ,csa_tree_add_7_25_groupi_n_4956 ,csa_tree_add_7_25_groupi_n_4908);
  or csa_tree_add_7_25_groupi_g16086(csa_tree_add_7_25_groupi_n_5003 ,csa_tree_add_7_25_groupi_n_4956 ,csa_tree_add_7_25_groupi_n_4908);
  and csa_tree_add_7_25_groupi_g16087(csa_tree_add_7_25_groupi_n_5002 ,csa_tree_add_7_25_groupi_n_4556 ,csa_tree_add_7_25_groupi_n_4964);
  or csa_tree_add_7_25_groupi_g16088(csa_tree_add_7_25_groupi_n_5001 ,csa_tree_add_7_25_groupi_n_3638 ,csa_tree_add_7_25_groupi_n_4979);
  or csa_tree_add_7_25_groupi_g16089(csa_tree_add_7_25_groupi_n_5000 ,csa_tree_add_7_25_groupi_n_3147 ,csa_tree_add_7_25_groupi_n_4984);
  or csa_tree_add_7_25_groupi_g16090(csa_tree_add_7_25_groupi_n_4999 ,csa_tree_add_7_25_groupi_n_3141 ,csa_tree_add_7_25_groupi_n_4980);
  or csa_tree_add_7_25_groupi_g16091(csa_tree_add_7_25_groupi_n_4998 ,csa_tree_add_7_25_groupi_n_3127 ,csa_tree_add_7_25_groupi_n_4953);
  and csa_tree_add_7_25_groupi_g16092(csa_tree_add_7_25_groupi_n_4997 ,csa_tree_add_7_25_groupi_n_4959 ,csa_tree_add_7_25_groupi_n_4910);
  or csa_tree_add_7_25_groupi_g16093(csa_tree_add_7_25_groupi_n_4996 ,csa_tree_add_7_25_groupi_n_3111 ,csa_tree_add_7_25_groupi_n_4951);
  or csa_tree_add_7_25_groupi_g16094(csa_tree_add_7_25_groupi_n_4995 ,csa_tree_add_7_25_groupi_n_3602 ,csa_tree_add_7_25_groupi_n_4977);
  or csa_tree_add_7_25_groupi_g16095(csa_tree_add_7_25_groupi_n_4994 ,csa_tree_add_7_25_groupi_n_3575 ,csa_tree_add_7_25_groupi_n_4976);
  or csa_tree_add_7_25_groupi_g16096(csa_tree_add_7_25_groupi_n_4993 ,csa_tree_add_7_25_groupi_n_3555 ,csa_tree_add_7_25_groupi_n_4975);
  xnor csa_tree_add_7_25_groupi_g16097(out2[2] ,csa_tree_add_7_25_groupi_n_4940 ,csa_tree_add_7_25_groupi_n_4831);
  nor csa_tree_add_7_25_groupi_g16098(csa_tree_add_7_25_groupi_n_4991 ,csa_tree_add_7_25_groupi_n_2950 ,csa_tree_add_7_25_groupi_n_4986);
  or csa_tree_add_7_25_groupi_g16099(csa_tree_add_7_25_groupi_n_4990 ,csa_tree_add_7_25_groupi_n_3035 ,csa_tree_add_7_25_groupi_n_4978);
  or csa_tree_add_7_25_groupi_g16100(csa_tree_add_7_25_groupi_n_5008 ,csa_tree_add_7_25_groupi_n_4784 ,csa_tree_add_7_25_groupi_n_4983);
  xnor csa_tree_add_7_25_groupi_g16101(csa_tree_add_7_25_groupi_n_5007 ,csa_tree_add_7_25_groupi_n_4939 ,csa_tree_add_7_25_groupi_n_2575);
  not csa_tree_add_7_25_groupi_g16102(csa_tree_add_7_25_groupi_n_4987 ,csa_tree_add_7_25_groupi_n_4988);
  nor csa_tree_add_7_25_groupi_g16103(csa_tree_add_7_25_groupi_n_4986 ,csa_tree_add_7_25_groupi_n_548 ,csa_tree_add_7_25_groupi_n_252);
  or csa_tree_add_7_25_groupi_g16104(csa_tree_add_7_25_groupi_n_4985 ,csa_tree_add_7_25_groupi_n_2421 ,csa_tree_add_7_25_groupi_n_4939);
  nor csa_tree_add_7_25_groupi_g16105(csa_tree_add_7_25_groupi_n_4984 ,csa_tree_add_7_25_groupi_n_2069 ,csa_tree_add_7_25_groupi_n_1825);
  and csa_tree_add_7_25_groupi_g16106(csa_tree_add_7_25_groupi_n_4983 ,csa_tree_add_7_25_groupi_n_4785 ,csa_tree_add_7_25_groupi_n_4940);
  and csa_tree_add_7_25_groupi_g16107(csa_tree_add_7_25_groupi_n_4982 ,csa_tree_add_7_25_groupi_n_4851 ,csa_tree_add_7_25_groupi_n_4936);
  or csa_tree_add_7_25_groupi_g16108(csa_tree_add_7_25_groupi_n_4981 ,csa_tree_add_7_25_groupi_n_4851 ,csa_tree_add_7_25_groupi_n_4936);
  nor csa_tree_add_7_25_groupi_g16109(csa_tree_add_7_25_groupi_n_4980 ,csa_tree_add_7_25_groupi_n_2165 ,csa_tree_add_7_25_groupi_n_1824);
  nor csa_tree_add_7_25_groupi_g16110(csa_tree_add_7_25_groupi_n_4979 ,csa_tree_add_7_25_groupi_n_1878 ,csa_tree_add_7_25_groupi_n_148);
  nor csa_tree_add_7_25_groupi_g16111(csa_tree_add_7_25_groupi_n_4978 ,csa_tree_add_7_25_groupi_n_254 ,csa_tree_add_7_25_groupi_n_2168);
  nor csa_tree_add_7_25_groupi_g16112(csa_tree_add_7_25_groupi_n_4977 ,csa_tree_add_7_25_groupi_n_740 ,csa_tree_add_7_25_groupi_n_255);
  nor csa_tree_add_7_25_groupi_g16113(csa_tree_add_7_25_groupi_n_4976 ,csa_tree_add_7_25_groupi_n_252 ,csa_tree_add_7_25_groupi_n_2197);
  nor csa_tree_add_7_25_groupi_g16114(csa_tree_add_7_25_groupi_n_4975 ,csa_tree_add_7_25_groupi_n_251 ,csa_tree_add_7_25_groupi_n_2052);
  nor csa_tree_add_7_25_groupi_g16115(csa_tree_add_7_25_groupi_n_4974 ,csa_tree_add_7_25_groupi_n_3487 ,csa_tree_add_7_25_groupi_n_4889);
  nor csa_tree_add_7_25_groupi_g16116(csa_tree_add_7_25_groupi_n_4973 ,csa_tree_add_7_25_groupi_n_4014 ,csa_tree_add_7_25_groupi_n_4897);
  nor csa_tree_add_7_25_groupi_g16117(csa_tree_add_7_25_groupi_n_4972 ,csa_tree_add_7_25_groupi_n_4089 ,csa_tree_add_7_25_groupi_n_4898);
  nor csa_tree_add_7_25_groupi_g16118(csa_tree_add_7_25_groupi_n_4971 ,csa_tree_add_7_25_groupi_n_4048 ,csa_tree_add_7_25_groupi_n_4896);
  nor csa_tree_add_7_25_groupi_g16119(csa_tree_add_7_25_groupi_n_4970 ,csa_tree_add_7_25_groupi_n_3997 ,csa_tree_add_7_25_groupi_n_4899);
  nor csa_tree_add_7_25_groupi_g16120(csa_tree_add_7_25_groupi_n_4969 ,csa_tree_add_7_25_groupi_n_3857 ,csa_tree_add_7_25_groupi_n_4891);
  nor csa_tree_add_7_25_groupi_g16121(csa_tree_add_7_25_groupi_n_4968 ,csa_tree_add_7_25_groupi_n_3855 ,csa_tree_add_7_25_groupi_n_4892);
  nor csa_tree_add_7_25_groupi_g16122(csa_tree_add_7_25_groupi_n_4967 ,csa_tree_add_7_25_groupi_n_3834 ,csa_tree_add_7_25_groupi_n_4895);
  nor csa_tree_add_7_25_groupi_g16123(csa_tree_add_7_25_groupi_n_4966 ,csa_tree_add_7_25_groupi_n_3827 ,csa_tree_add_7_25_groupi_n_4901);
  nor csa_tree_add_7_25_groupi_g16124(csa_tree_add_7_25_groupi_n_4965 ,csa_tree_add_7_25_groupi_n_4058 ,csa_tree_add_7_25_groupi_n_4900);
  and csa_tree_add_7_25_groupi_g16125(csa_tree_add_7_25_groupi_n_4989 ,csa_tree_add_7_25_groupi_n_3904 ,csa_tree_add_7_25_groupi_n_4890);
  or csa_tree_add_7_25_groupi_g16126(csa_tree_add_7_25_groupi_n_4988 ,csa_tree_add_7_25_groupi_n_4479 ,csa_tree_add_7_25_groupi_n_4929);
  nor csa_tree_add_7_25_groupi_g16127(csa_tree_add_7_25_groupi_n_4953 ,csa_tree_add_7_25_groupi_n_2144 ,csa_tree_add_7_25_groupi_n_148);
  nor csa_tree_add_7_25_groupi_g16128(csa_tree_add_7_25_groupi_n_4952 ,csa_tree_add_7_25_groupi_n_255 ,csa_tree_add_7_25_groupi_n_2090);
  nor csa_tree_add_7_25_groupi_g16129(csa_tree_add_7_25_groupi_n_4951 ,csa_tree_add_7_25_groupi_n_2111 ,csa_tree_add_7_25_groupi_n_1824);
  xnor csa_tree_add_7_25_groupi_g16130(csa_tree_add_7_25_groupi_n_4950 ,csa_tree_add_7_25_groupi_n_4854 ,csa_tree_add_7_25_groupi_n_4793);
  xnor csa_tree_add_7_25_groupi_g16131(csa_tree_add_7_25_groupi_n_4949 ,csa_tree_add_7_25_groupi_n_4850 ,csa_tree_add_7_25_groupi_n_4800);
  xnor csa_tree_add_7_25_groupi_g16132(csa_tree_add_7_25_groupi_n_4948 ,csa_tree_add_7_25_groupi_n_4853 ,csa_tree_add_7_25_groupi_n_4801);
  xnor csa_tree_add_7_25_groupi_g16133(csa_tree_add_7_25_groupi_n_4947 ,csa_tree_add_7_25_groupi_n_1102 ,csa_tree_add_7_25_groupi_n_1107);
  xnor csa_tree_add_7_25_groupi_g16134(csa_tree_add_7_25_groupi_n_4946 ,csa_tree_add_7_25_groupi_n_4855 ,csa_tree_add_7_25_groupi_n_4799);
  xnor csa_tree_add_7_25_groupi_g16135(csa_tree_add_7_25_groupi_n_4945 ,csa_tree_add_7_25_groupi_n_4852 ,csa_tree_add_7_25_groupi_n_4798);
  xnor csa_tree_add_7_25_groupi_g16136(csa_tree_add_7_25_groupi_n_4944 ,csa_tree_add_7_25_groupi_n_4849 ,csa_tree_add_7_25_groupi_n_4797);
  xnor csa_tree_add_7_25_groupi_g16137(csa_tree_add_7_25_groupi_n_4943 ,csa_tree_add_7_25_groupi_n_4848 ,csa_tree_add_7_25_groupi_n_4796);
  xnor csa_tree_add_7_25_groupi_g16138(csa_tree_add_7_25_groupi_n_4942 ,csa_tree_add_7_25_groupi_n_4847 ,csa_tree_add_7_25_groupi_n_4795);
  xnor csa_tree_add_7_25_groupi_g16139(csa_tree_add_7_25_groupi_n_4941 ,csa_tree_add_7_25_groupi_n_4846 ,csa_tree_add_7_25_groupi_n_4794);
  xnor csa_tree_add_7_25_groupi_g16140(csa_tree_add_7_25_groupi_n_4964 ,csa_tree_add_7_25_groupi_n_4864 ,in3[29]);
  xnor csa_tree_add_7_25_groupi_g16141(csa_tree_add_7_25_groupi_n_4963 ,csa_tree_add_7_25_groupi_n_4861 ,in3[8]);
  xnor csa_tree_add_7_25_groupi_g16142(csa_tree_add_7_25_groupi_n_4962 ,csa_tree_add_7_25_groupi_n_4858 ,in3[5]);
  xnor csa_tree_add_7_25_groupi_g16143(csa_tree_add_7_25_groupi_n_4961 ,csa_tree_add_7_25_groupi_n_4863 ,in3[11]);
  xnor csa_tree_add_7_25_groupi_g16144(csa_tree_add_7_25_groupi_n_4960 ,csa_tree_add_7_25_groupi_n_4859 ,in3[2]);
  xnor csa_tree_add_7_25_groupi_g16145(csa_tree_add_7_25_groupi_n_4959 ,csa_tree_add_7_25_groupi_n_4866 ,in3[14]);
  xnor csa_tree_add_7_25_groupi_g16146(csa_tree_add_7_25_groupi_n_4958 ,csa_tree_add_7_25_groupi_n_4860 ,in3[17]);
  xnor csa_tree_add_7_25_groupi_g16147(csa_tree_add_7_25_groupi_n_4957 ,csa_tree_add_7_25_groupi_n_4856 ,csa_tree_add_7_25_groupi_n_4505);
  xnor csa_tree_add_7_25_groupi_g16148(csa_tree_add_7_25_groupi_n_4956 ,csa_tree_add_7_25_groupi_n_4862 ,in3[20]);
  xnor csa_tree_add_7_25_groupi_g16149(csa_tree_add_7_25_groupi_n_4955 ,csa_tree_add_7_25_groupi_n_4865 ,in3[26]);
  xnor csa_tree_add_7_25_groupi_g16150(csa_tree_add_7_25_groupi_n_4954 ,csa_tree_add_7_25_groupi_n_4857 ,in3[23]);
  and csa_tree_add_7_25_groupi_g16151(csa_tree_add_7_25_groupi_n_4929 ,csa_tree_add_7_25_groupi_n_4476 ,csa_tree_add_7_25_groupi_n_4856);
  and csa_tree_add_7_25_groupi_g16152(csa_tree_add_7_25_groupi_n_4928 ,csa_tree_add_7_25_groupi_n_4853 ,csa_tree_add_7_25_groupi_n_4801);
  or csa_tree_add_7_25_groupi_g16153(csa_tree_add_7_25_groupi_n_4927 ,csa_tree_add_7_25_groupi_n_4855 ,csa_tree_add_7_25_groupi_n_4799);
  and csa_tree_add_7_25_groupi_g16154(csa_tree_add_7_25_groupi_n_4926 ,csa_tree_add_7_25_groupi_n_4847 ,csa_tree_add_7_25_groupi_n_4795);
  or csa_tree_add_7_25_groupi_g16155(csa_tree_add_7_25_groupi_n_4925 ,csa_tree_add_7_25_groupi_n_4847 ,csa_tree_add_7_25_groupi_n_4795);
  and csa_tree_add_7_25_groupi_g16156(csa_tree_add_7_25_groupi_n_4924 ,csa_tree_add_7_25_groupi_n_4855 ,csa_tree_add_7_25_groupi_n_4799);
  or csa_tree_add_7_25_groupi_g16157(csa_tree_add_7_25_groupi_n_4923 ,csa_tree_add_7_25_groupi_n_4852 ,csa_tree_add_7_25_groupi_n_4798);
  and csa_tree_add_7_25_groupi_g16158(csa_tree_add_7_25_groupi_n_4922 ,csa_tree_add_7_25_groupi_n_4852 ,csa_tree_add_7_25_groupi_n_4798);
  and csa_tree_add_7_25_groupi_g16159(csa_tree_add_7_25_groupi_n_4921 ,csa_tree_add_7_25_groupi_n_4848 ,csa_tree_add_7_25_groupi_n_4796);
  or csa_tree_add_7_25_groupi_g16160(csa_tree_add_7_25_groupi_n_4920 ,csa_tree_add_7_25_groupi_n_4848 ,csa_tree_add_7_25_groupi_n_4796);
  or csa_tree_add_7_25_groupi_g16161(csa_tree_add_7_25_groupi_n_4919 ,csa_tree_add_7_25_groupi_n_4853 ,csa_tree_add_7_25_groupi_n_4801);
  or csa_tree_add_7_25_groupi_g16162(csa_tree_add_7_25_groupi_n_4918 ,csa_tree_add_7_25_groupi_n_4849 ,csa_tree_add_7_25_groupi_n_4797);
  and csa_tree_add_7_25_groupi_g16163(csa_tree_add_7_25_groupi_n_4917 ,csa_tree_add_7_25_groupi_n_4854 ,csa_tree_add_7_25_groupi_n_4793);
  and csa_tree_add_7_25_groupi_g16164(csa_tree_add_7_25_groupi_n_4916 ,csa_tree_add_7_25_groupi_n_4849 ,csa_tree_add_7_25_groupi_n_4797);
  or csa_tree_add_7_25_groupi_g16165(csa_tree_add_7_25_groupi_n_4915 ,csa_tree_add_7_25_groupi_n_4850 ,csa_tree_add_7_25_groupi_n_4800);
  or csa_tree_add_7_25_groupi_g16166(csa_tree_add_7_25_groupi_n_4914 ,csa_tree_add_7_25_groupi_n_4854 ,csa_tree_add_7_25_groupi_n_4793);
  and csa_tree_add_7_25_groupi_g16167(csa_tree_add_7_25_groupi_n_4913 ,csa_tree_add_7_25_groupi_n_4850 ,csa_tree_add_7_25_groupi_n_4800);
  or csa_tree_add_7_25_groupi_g16168(csa_tree_add_7_25_groupi_n_4940 ,csa_tree_add_7_25_groupi_n_4700 ,csa_tree_add_7_25_groupi_n_4874);
  and csa_tree_add_7_25_groupi_g16169(csa_tree_add_7_25_groupi_n_4939 ,csa_tree_add_7_25_groupi_n_2420 ,csa_tree_add_7_25_groupi_n_4880);
  or csa_tree_add_7_25_groupi_g16170(csa_tree_add_7_25_groupi_n_4938 ,csa_tree_add_7_25_groupi_n_4695 ,csa_tree_add_7_25_groupi_n_4867);
  or csa_tree_add_7_25_groupi_g16171(csa_tree_add_7_25_groupi_n_4937 ,csa_tree_add_7_25_groupi_n_4712 ,csa_tree_add_7_25_groupi_n_4868);
  or csa_tree_add_7_25_groupi_g16172(csa_tree_add_7_25_groupi_n_4936 ,csa_tree_add_7_25_groupi_n_4703 ,csa_tree_add_7_25_groupi_n_4872);
  or csa_tree_add_7_25_groupi_g16173(csa_tree_add_7_25_groupi_n_4935 ,csa_tree_add_7_25_groupi_n_4692 ,csa_tree_add_7_25_groupi_n_4870);
  or csa_tree_add_7_25_groupi_g16174(csa_tree_add_7_25_groupi_n_4934 ,csa_tree_add_7_25_groupi_n_4699 ,csa_tree_add_7_25_groupi_n_4871);
  or csa_tree_add_7_25_groupi_g16175(csa_tree_add_7_25_groupi_n_4933 ,csa_tree_add_7_25_groupi_n_4704 ,csa_tree_add_7_25_groupi_n_4881);
  or csa_tree_add_7_25_groupi_g16176(csa_tree_add_7_25_groupi_n_4932 ,csa_tree_add_7_25_groupi_n_4707 ,csa_tree_add_7_25_groupi_n_4873);
  or csa_tree_add_7_25_groupi_g16177(csa_tree_add_7_25_groupi_n_4931 ,csa_tree_add_7_25_groupi_n_4696 ,csa_tree_add_7_25_groupi_n_4869);
  or csa_tree_add_7_25_groupi_g16178(csa_tree_add_7_25_groupi_n_4930 ,csa_tree_add_7_25_groupi_n_4708 ,csa_tree_add_7_25_groupi_n_4879);
  and csa_tree_add_7_25_groupi_g16179(csa_tree_add_7_25_groupi_n_4902 ,csa_tree_add_7_25_groupi_n_4846 ,csa_tree_add_7_25_groupi_n_4794);
  or csa_tree_add_7_25_groupi_g16180(csa_tree_add_7_25_groupi_n_4901 ,csa_tree_add_7_25_groupi_n_3610 ,csa_tree_add_7_25_groupi_n_4876);
  or csa_tree_add_7_25_groupi_g16181(csa_tree_add_7_25_groupi_n_4900 ,csa_tree_add_7_25_groupi_n_3151 ,csa_tree_add_7_25_groupi_n_4843);
  or csa_tree_add_7_25_groupi_g16182(csa_tree_add_7_25_groupi_n_4899 ,csa_tree_add_7_25_groupi_n_3143 ,csa_tree_add_7_25_groupi_n_4842);
  or csa_tree_add_7_25_groupi_g16183(csa_tree_add_7_25_groupi_n_4898 ,csa_tree_add_7_25_groupi_n_3112 ,csa_tree_add_7_25_groupi_n_4841);
  or csa_tree_add_7_25_groupi_g16184(csa_tree_add_7_25_groupi_n_4897 ,csa_tree_add_7_25_groupi_n_3110 ,csa_tree_add_7_25_groupi_n_4840);
  or csa_tree_add_7_25_groupi_g16185(csa_tree_add_7_25_groupi_n_4896 ,csa_tree_add_7_25_groupi_n_3128 ,csa_tree_add_7_25_groupi_n_4839);
  or csa_tree_add_7_25_groupi_g16186(csa_tree_add_7_25_groupi_n_4895 ,csa_tree_add_7_25_groupi_n_3596 ,csa_tree_add_7_25_groupi_n_4878);
  or csa_tree_add_7_25_groupi_g16187(csa_tree_add_7_25_groupi_n_4894 ,in3[8] ,csa_tree_add_7_25_groupi_n_1098);
  and csa_tree_add_7_25_groupi_g16188(csa_tree_add_7_25_groupi_n_4893 ,in3[8] ,csa_tree_add_7_25_groupi_n_1107);
  or csa_tree_add_7_25_groupi_g16189(csa_tree_add_7_25_groupi_n_4892 ,csa_tree_add_7_25_groupi_n_3611 ,csa_tree_add_7_25_groupi_n_4882);
  or csa_tree_add_7_25_groupi_g16190(csa_tree_add_7_25_groupi_n_4891 ,csa_tree_add_7_25_groupi_n_3571 ,csa_tree_add_7_25_groupi_n_4838);
  nor csa_tree_add_7_25_groupi_g16191(csa_tree_add_7_25_groupi_n_4890 ,csa_tree_add_7_25_groupi_n_2983 ,csa_tree_add_7_25_groupi_n_4875);
  or csa_tree_add_7_25_groupi_g16192(csa_tree_add_7_25_groupi_n_4889 ,csa_tree_add_7_25_groupi_n_3033 ,csa_tree_add_7_25_groupi_n_4877);
  nor csa_tree_add_7_25_groupi_g16193(csa_tree_add_7_25_groupi_n_4888 ,csa_tree_add_7_25_groupi_n_4771 ,csa_tree_add_7_25_groupi_n_2344);
  or csa_tree_add_7_25_groupi_g16194(csa_tree_add_7_25_groupi_n_4887 ,csa_tree_add_7_25_groupi_n_4772 ,csa_tree_add_7_25_groupi_n_1098);
  or csa_tree_add_7_25_groupi_g16195(csa_tree_add_7_25_groupi_n_4886 ,csa_tree_add_7_25_groupi_n_4846 ,csa_tree_add_7_25_groupi_n_4794);
  xnor csa_tree_add_7_25_groupi_g16196(out2[1] ,csa_tree_add_7_25_groupi_n_4826 ,csa_tree_add_7_25_groupi_n_4725);
  xnor csa_tree_add_7_25_groupi_g16197(csa_tree_add_7_25_groupi_n_4912 ,csa_tree_add_7_25_groupi_n_4828 ,csa_tree_add_7_25_groupi_n_4726);
  xnor csa_tree_add_7_25_groupi_g16198(csa_tree_add_7_25_groupi_n_4911 ,csa_tree_add_7_25_groupi_n_4825 ,csa_tree_add_7_25_groupi_n_4723);
  xnor csa_tree_add_7_25_groupi_g16199(csa_tree_add_7_25_groupi_n_4910 ,csa_tree_add_7_25_groupi_n_4821 ,csa_tree_add_7_25_groupi_n_4722);
  xnor csa_tree_add_7_25_groupi_g16200(csa_tree_add_7_25_groupi_n_4909 ,csa_tree_add_7_25_groupi_n_4819 ,csa_tree_add_7_25_groupi_n_4721);
  xnor csa_tree_add_7_25_groupi_g16201(csa_tree_add_7_25_groupi_n_4908 ,csa_tree_add_7_25_groupi_n_4822 ,csa_tree_add_7_25_groupi_n_4720);
  xnor csa_tree_add_7_25_groupi_g16202(csa_tree_add_7_25_groupi_n_4907 ,csa_tree_add_7_25_groupi_n_4824 ,csa_tree_add_7_25_groupi_n_4719);
  xnor csa_tree_add_7_25_groupi_g16203(csa_tree_add_7_25_groupi_n_4906 ,csa_tree_add_7_25_groupi_n_4823 ,csa_tree_add_7_25_groupi_n_4728);
  xnor csa_tree_add_7_25_groupi_g16204(csa_tree_add_7_25_groupi_n_4905 ,csa_tree_add_7_25_groupi_n_4827 ,csa_tree_add_7_25_groupi_n_4727);
  xnor csa_tree_add_7_25_groupi_g16205(csa_tree_add_7_25_groupi_n_4904 ,csa_tree_add_7_25_groupi_n_4818 ,csa_tree_add_7_25_groupi_n_4724);
  xnor csa_tree_add_7_25_groupi_g16206(csa_tree_add_7_25_groupi_n_4903 ,csa_tree_add_7_25_groupi_n_4820 ,csa_tree_add_7_25_groupi_n_2585);
  nor csa_tree_add_7_25_groupi_g16208(csa_tree_add_7_25_groupi_n_4882 ,csa_tree_add_7_25_groupi_n_306 ,csa_tree_add_7_25_groupi_n_2024);
  and csa_tree_add_7_25_groupi_g16209(csa_tree_add_7_25_groupi_n_4881 ,csa_tree_add_7_25_groupi_n_4709 ,csa_tree_add_7_25_groupi_n_4822);
  or csa_tree_add_7_25_groupi_g16210(csa_tree_add_7_25_groupi_n_4880 ,csa_tree_add_7_25_groupi_n_2490 ,csa_tree_add_7_25_groupi_n_4820);
  and csa_tree_add_7_25_groupi_g16211(csa_tree_add_7_25_groupi_n_4879 ,csa_tree_add_7_25_groupi_n_4711 ,csa_tree_add_7_25_groupi_n_4824);
  nor csa_tree_add_7_25_groupi_g16212(csa_tree_add_7_25_groupi_n_4878 ,csa_tree_add_7_25_groupi_n_1861 ,csa_tree_add_7_25_groupi_n_1309);
  nor csa_tree_add_7_25_groupi_g16213(csa_tree_add_7_25_groupi_n_4877 ,csa_tree_add_7_25_groupi_n_2183 ,csa_tree_add_7_25_groupi_n_1861);
  nor csa_tree_add_7_25_groupi_g16214(csa_tree_add_7_25_groupi_n_4876 ,csa_tree_add_7_25_groupi_n_1878 ,csa_tree_add_7_25_groupi_n_145);
  nor csa_tree_add_7_25_groupi_g16215(csa_tree_add_7_25_groupi_n_4875 ,csa_tree_add_7_25_groupi_n_639 ,csa_tree_add_7_25_groupi_n_289);
  and csa_tree_add_7_25_groupi_g16216(csa_tree_add_7_25_groupi_n_4874 ,csa_tree_add_7_25_groupi_n_4705 ,csa_tree_add_7_25_groupi_n_4826);
  and csa_tree_add_7_25_groupi_g16217(csa_tree_add_7_25_groupi_n_4873 ,csa_tree_add_7_25_groupi_n_4710 ,csa_tree_add_7_25_groupi_n_4818);
  and csa_tree_add_7_25_groupi_g16218(csa_tree_add_7_25_groupi_n_4872 ,csa_tree_add_7_25_groupi_n_4702 ,csa_tree_add_7_25_groupi_n_4823);
  and csa_tree_add_7_25_groupi_g16219(csa_tree_add_7_25_groupi_n_4871 ,csa_tree_add_7_25_groupi_n_4701 ,csa_tree_add_7_25_groupi_n_4825);
  and csa_tree_add_7_25_groupi_g16220(csa_tree_add_7_25_groupi_n_4870 ,csa_tree_add_7_25_groupi_n_4697 ,csa_tree_add_7_25_groupi_n_4821);
  and csa_tree_add_7_25_groupi_g16221(csa_tree_add_7_25_groupi_n_4869 ,csa_tree_add_7_25_groupi_n_4694 ,csa_tree_add_7_25_groupi_n_4827);
  and csa_tree_add_7_25_groupi_g16222(csa_tree_add_7_25_groupi_n_4868 ,csa_tree_add_7_25_groupi_n_4698 ,csa_tree_add_7_25_groupi_n_4819);
  and csa_tree_add_7_25_groupi_g16223(csa_tree_add_7_25_groupi_n_4867 ,csa_tree_add_7_25_groupi_n_4693 ,csa_tree_add_7_25_groupi_n_4828);
  nor csa_tree_add_7_25_groupi_g16224(csa_tree_add_7_25_groupi_n_4866 ,csa_tree_add_7_25_groupi_n_4067 ,csa_tree_add_7_25_groupi_n_4803);
  nor csa_tree_add_7_25_groupi_g16225(csa_tree_add_7_25_groupi_n_4865 ,csa_tree_add_7_25_groupi_n_3944 ,csa_tree_add_7_25_groupi_n_4790);
  nor csa_tree_add_7_25_groupi_g16226(csa_tree_add_7_25_groupi_n_4864 ,csa_tree_add_7_25_groupi_n_3996 ,csa_tree_add_7_25_groupi_n_4806);
  nor csa_tree_add_7_25_groupi_g16227(csa_tree_add_7_25_groupi_n_4863 ,csa_tree_add_7_25_groupi_n_4051 ,csa_tree_add_7_25_groupi_n_4817);
  nor csa_tree_add_7_25_groupi_g16228(csa_tree_add_7_25_groupi_n_4862 ,csa_tree_add_7_25_groupi_n_3949 ,csa_tree_add_7_25_groupi_n_4788);
  nor csa_tree_add_7_25_groupi_g16229(csa_tree_add_7_25_groupi_n_4861 ,csa_tree_add_7_25_groupi_n_4046 ,csa_tree_add_7_25_groupi_n_4791);
  nor csa_tree_add_7_25_groupi_g16230(csa_tree_add_7_25_groupi_n_4860 ,csa_tree_add_7_25_groupi_n_4070 ,csa_tree_add_7_25_groupi_n_4805);
  nor csa_tree_add_7_25_groupi_g16231(csa_tree_add_7_25_groupi_n_4859 ,csa_tree_add_7_25_groupi_n_3471 ,csa_tree_add_7_25_groupi_n_4776);
  nor csa_tree_add_7_25_groupi_g16232(csa_tree_add_7_25_groupi_n_4858 ,csa_tree_add_7_25_groupi_n_4030 ,csa_tree_add_7_25_groupi_n_4804);
  nor csa_tree_add_7_25_groupi_g16233(csa_tree_add_7_25_groupi_n_4857 ,csa_tree_add_7_25_groupi_n_3898 ,csa_tree_add_7_25_groupi_n_4789);
  or csa_tree_add_7_25_groupi_g16234(csa_tree_add_7_25_groupi_n_4884 ,csa_tree_add_7_25_groupi_n_4444 ,csa_tree_add_7_25_groupi_n_4807);
  and csa_tree_add_7_25_groupi_g16235(csa_tree_add_7_25_groupi_n_4883 ,csa_tree_add_7_25_groupi_n_3869 ,csa_tree_add_7_25_groupi_n_4783);
  not csa_tree_add_7_25_groupi_g16236(csa_tree_add_7_25_groupi_n_4844 ,csa_tree_add_7_25_groupi_n_4845);
  nor csa_tree_add_7_25_groupi_g16237(csa_tree_add_7_25_groupi_n_4843 ,csa_tree_add_7_25_groupi_n_305 ,csa_tree_add_7_25_groupi_n_2057);
  nor csa_tree_add_7_25_groupi_g16238(csa_tree_add_7_25_groupi_n_4842 ,csa_tree_add_7_25_groupi_n_288 ,csa_tree_add_7_25_groupi_n_2141);
  nor csa_tree_add_7_25_groupi_g16239(csa_tree_add_7_25_groupi_n_4841 ,csa_tree_add_7_25_groupi_n_306 ,csa_tree_add_7_25_groupi_n_2156);
  nor csa_tree_add_7_25_groupi_g16240(csa_tree_add_7_25_groupi_n_4840 ,csa_tree_add_7_25_groupi_n_2102 ,csa_tree_add_7_25_groupi_n_145);
  nor csa_tree_add_7_25_groupi_g16241(csa_tree_add_7_25_groupi_n_4839 ,csa_tree_add_7_25_groupi_n_289 ,csa_tree_add_7_25_groupi_n_2123);
  nor csa_tree_add_7_25_groupi_g16242(csa_tree_add_7_25_groupi_n_4838 ,csa_tree_add_7_25_groupi_n_2052 ,csa_tree_add_7_25_groupi_n_1862);
  xnor csa_tree_add_7_25_groupi_g16243(csa_tree_add_7_25_groupi_n_4837 ,csa_tree_add_7_25_groupi_n_4740 ,csa_tree_add_7_25_groupi_n_4683);
  xnor csa_tree_add_7_25_groupi_g16244(csa_tree_add_7_25_groupi_n_4836 ,csa_tree_add_7_25_groupi_n_4739 ,csa_tree_add_7_25_groupi_n_4677);
  xnor csa_tree_add_7_25_groupi_g16245(csa_tree_add_7_25_groupi_n_4835 ,csa_tree_add_7_25_groupi_n_4738 ,csa_tree_add_7_25_groupi_n_4684);
  xnor csa_tree_add_7_25_groupi_g16246(csa_tree_add_7_25_groupi_n_4834 ,csa_tree_add_7_25_groupi_n_4737 ,csa_tree_add_7_25_groupi_n_4685);
  xnor csa_tree_add_7_25_groupi_g16248(csa_tree_add_7_25_groupi_n_4833 ,csa_tree_add_7_25_groupi_n_4736 ,csa_tree_add_7_25_groupi_n_4681);
  xnor csa_tree_add_7_25_groupi_g16249(csa_tree_add_7_25_groupi_n_4832 ,csa_tree_add_7_25_groupi_n_4741 ,csa_tree_add_7_25_groupi_n_4682);
  xnor csa_tree_add_7_25_groupi_g16250(csa_tree_add_7_25_groupi_n_4831 ,csa_tree_add_7_25_groupi_n_4742 ,csa_tree_add_7_25_groupi_n_4679);
  xnor csa_tree_add_7_25_groupi_g16251(csa_tree_add_7_25_groupi_n_4830 ,csa_tree_add_7_25_groupi_n_4744 ,csa_tree_add_7_25_groupi_n_4678);
  xnor csa_tree_add_7_25_groupi_g16252(csa_tree_add_7_25_groupi_n_4829 ,csa_tree_add_7_25_groupi_n_4743 ,csa_tree_add_7_25_groupi_n_4680);
  xnor csa_tree_add_7_25_groupi_g16253(csa_tree_add_7_25_groupi_n_4856 ,csa_tree_add_7_25_groupi_n_4751 ,in3[29]);
  xnor csa_tree_add_7_25_groupi_g16254(csa_tree_add_7_25_groupi_n_4855 ,csa_tree_add_7_25_groupi_n_4753 ,in3[11]);
  xnor csa_tree_add_7_25_groupi_g16255(csa_tree_add_7_25_groupi_n_4854 ,csa_tree_add_7_25_groupi_n_4746 ,in3[8]);
  xnor csa_tree_add_7_25_groupi_g16256(csa_tree_add_7_25_groupi_n_4853 ,csa_tree_add_7_25_groupi_n_4748 ,in3[2]);
  xnor csa_tree_add_7_25_groupi_g16257(csa_tree_add_7_25_groupi_n_4852 ,csa_tree_add_7_25_groupi_n_4755 ,in3[14]);
  xnor csa_tree_add_7_25_groupi_g16258(csa_tree_add_7_25_groupi_n_4851 ,csa_tree_add_7_25_groupi_n_4745 ,csa_tree_add_7_25_groupi_n_4504);
  xnor csa_tree_add_7_25_groupi_g16259(csa_tree_add_7_25_groupi_n_4850 ,csa_tree_add_7_25_groupi_n_4749 ,in3[5]);
  xnor csa_tree_add_7_25_groupi_g16260(csa_tree_add_7_25_groupi_n_4849 ,csa_tree_add_7_25_groupi_n_4747 ,in3[17]);
  xnor csa_tree_add_7_25_groupi_g16261(csa_tree_add_7_25_groupi_n_4848 ,csa_tree_add_7_25_groupi_n_4754 ,in3[20]);
  xnor csa_tree_add_7_25_groupi_g16262(csa_tree_add_7_25_groupi_n_4847 ,csa_tree_add_7_25_groupi_n_4750 ,in3[23]);
  xnor csa_tree_add_7_25_groupi_g16263(csa_tree_add_7_25_groupi_n_4846 ,csa_tree_add_7_25_groupi_n_4752 ,in3[26]);
  xnor csa_tree_add_7_25_groupi_g16264(csa_tree_add_7_25_groupi_n_4845 ,csa_tree_add_7_25_groupi_n_4718 ,csa_tree_add_7_25_groupi_n_4554);
  or csa_tree_add_7_25_groupi_g16265(csa_tree_add_7_25_groupi_n_4817 ,csa_tree_add_7_25_groupi_n_3105 ,csa_tree_add_7_25_groupi_n_4731);
  or csa_tree_add_7_25_groupi_g16266(csa_tree_add_7_25_groupi_n_4816 ,csa_tree_add_7_25_groupi_n_4737 ,csa_tree_add_7_25_groupi_n_4685);
  nor csa_tree_add_7_25_groupi_g16267(csa_tree_add_7_25_groupi_n_4815 ,csa_tree_add_7_25_groupi_n_4772 ,csa_tree_add_7_25_groupi_n_4774);
  or csa_tree_add_7_25_groupi_g16268(csa_tree_add_7_25_groupi_n_4814 ,csa_tree_add_7_25_groupi_n_1102 ,csa_tree_add_7_25_groupi_n_4773);
  and csa_tree_add_7_25_groupi_g16269(csa_tree_add_7_25_groupi_n_4813 ,csa_tree_add_7_25_groupi_n_4738 ,csa_tree_add_7_25_groupi_n_4684);
  or csa_tree_add_7_25_groupi_g16270(csa_tree_add_7_25_groupi_n_4812 ,csa_tree_add_7_25_groupi_n_4738 ,csa_tree_add_7_25_groupi_n_4684);
  and csa_tree_add_7_25_groupi_g16271(csa_tree_add_7_25_groupi_n_4811 ,csa_tree_add_7_25_groupi_n_4739 ,csa_tree_add_7_25_groupi_n_4677);
  or csa_tree_add_7_25_groupi_g16272(csa_tree_add_7_25_groupi_n_4810 ,csa_tree_add_7_25_groupi_n_4739 ,csa_tree_add_7_25_groupi_n_4677);
  or csa_tree_add_7_25_groupi_g16273(csa_tree_add_7_25_groupi_n_4809 ,csa_tree_add_7_25_groupi_n_4740 ,csa_tree_add_7_25_groupi_n_4683);
  and csa_tree_add_7_25_groupi_g16274(csa_tree_add_7_25_groupi_n_4808 ,csa_tree_add_7_25_groupi_n_4740 ,csa_tree_add_7_25_groupi_n_4683);
  and csa_tree_add_7_25_groupi_g16275(csa_tree_add_7_25_groupi_n_4807 ,csa_tree_add_7_25_groupi_n_4745 ,csa_tree_add_7_25_groupi_n_4445);
  or csa_tree_add_7_25_groupi_g16276(csa_tree_add_7_25_groupi_n_4806 ,csa_tree_add_7_25_groupi_n_3024 ,csa_tree_add_7_25_groupi_n_4756);
  or csa_tree_add_7_25_groupi_g16277(csa_tree_add_7_25_groupi_n_4805 ,csa_tree_add_7_25_groupi_n_3146 ,csa_tree_add_7_25_groupi_n_4734);
  or csa_tree_add_7_25_groupi_g16278(csa_tree_add_7_25_groupi_n_4804 ,csa_tree_add_7_25_groupi_n_3134 ,csa_tree_add_7_25_groupi_n_4733);
  or csa_tree_add_7_25_groupi_g16279(csa_tree_add_7_25_groupi_n_4803 ,csa_tree_add_7_25_groupi_n_3107 ,csa_tree_add_7_25_groupi_n_4732);
  and csa_tree_add_7_25_groupi_g16280(csa_tree_add_7_25_groupi_n_4802 ,csa_tree_add_7_25_groupi_n_4737 ,csa_tree_add_7_25_groupi_n_4685);
  or csa_tree_add_7_25_groupi_g16281(csa_tree_add_7_25_groupi_n_4828 ,csa_tree_add_7_25_groupi_n_4588 ,csa_tree_add_7_25_groupi_n_4759);
  or csa_tree_add_7_25_groupi_g16282(csa_tree_add_7_25_groupi_n_4827 ,csa_tree_add_7_25_groupi_n_4555 ,csa_tree_add_7_25_groupi_n_4760);
  or csa_tree_add_7_25_groupi_g16283(csa_tree_add_7_25_groupi_n_4826 ,csa_tree_add_7_25_groupi_n_4592 ,csa_tree_add_7_25_groupi_n_4764);
  or csa_tree_add_7_25_groupi_g16284(csa_tree_add_7_25_groupi_n_4825 ,csa_tree_add_7_25_groupi_n_4598 ,csa_tree_add_7_25_groupi_n_4765);
  or csa_tree_add_7_25_groupi_g16285(csa_tree_add_7_25_groupi_n_4824 ,csa_tree_add_7_25_groupi_n_4599 ,csa_tree_add_7_25_groupi_n_4770);
  or csa_tree_add_7_25_groupi_g16286(csa_tree_add_7_25_groupi_n_4823 ,csa_tree_add_7_25_groupi_n_4572 ,csa_tree_add_7_25_groupi_n_4758);
  or csa_tree_add_7_25_groupi_g16287(csa_tree_add_7_25_groupi_n_4822 ,csa_tree_add_7_25_groupi_n_4600 ,csa_tree_add_7_25_groupi_n_4766);
  or csa_tree_add_7_25_groupi_g16288(csa_tree_add_7_25_groupi_n_4821 ,csa_tree_add_7_25_groupi_n_4583 ,csa_tree_add_7_25_groupi_n_4769);
  and csa_tree_add_7_25_groupi_g16289(csa_tree_add_7_25_groupi_n_4820 ,csa_tree_add_7_25_groupi_n_2463 ,csa_tree_add_7_25_groupi_n_4768);
  or csa_tree_add_7_25_groupi_g16290(csa_tree_add_7_25_groupi_n_4819 ,csa_tree_add_7_25_groupi_n_4589 ,csa_tree_add_7_25_groupi_n_4762);
  or csa_tree_add_7_25_groupi_g16291(csa_tree_add_7_25_groupi_n_4818 ,csa_tree_add_7_25_groupi_n_4587 ,csa_tree_add_7_25_groupi_n_4761);
  or csa_tree_add_7_25_groupi_g16292(csa_tree_add_7_25_groupi_n_4791 ,csa_tree_add_7_25_groupi_n_3100 ,csa_tree_add_7_25_groupi_n_4730);
  or csa_tree_add_7_25_groupi_g16293(csa_tree_add_7_25_groupi_n_4790 ,csa_tree_add_7_25_groupi_n_3586 ,csa_tree_add_7_25_groupi_n_4763);
  or csa_tree_add_7_25_groupi_g16294(csa_tree_add_7_25_groupi_n_4789 ,csa_tree_add_7_25_groupi_n_3588 ,csa_tree_add_7_25_groupi_n_4735);
  or csa_tree_add_7_25_groupi_g16295(csa_tree_add_7_25_groupi_n_4788 ,csa_tree_add_7_25_groupi_n_3562 ,csa_tree_add_7_25_groupi_n_4729);
  and csa_tree_add_7_25_groupi_g16296(csa_tree_add_7_25_groupi_n_4787 ,csa_tree_add_7_25_groupi_n_4741 ,csa_tree_add_7_25_groupi_n_4682);
  or csa_tree_add_7_25_groupi_g16297(csa_tree_add_7_25_groupi_n_4786 ,csa_tree_add_7_25_groupi_n_4741 ,csa_tree_add_7_25_groupi_n_4682);
  or csa_tree_add_7_25_groupi_g16298(csa_tree_add_7_25_groupi_n_4785 ,csa_tree_add_7_25_groupi_n_4742 ,csa_tree_add_7_25_groupi_n_4679);
  and csa_tree_add_7_25_groupi_g16299(csa_tree_add_7_25_groupi_n_4784 ,csa_tree_add_7_25_groupi_n_4742 ,csa_tree_add_7_25_groupi_n_4679);
  nor csa_tree_add_7_25_groupi_g16300(csa_tree_add_7_25_groupi_n_4783 ,csa_tree_add_7_25_groupi_n_2947 ,csa_tree_add_7_25_groupi_n_4757);
  and csa_tree_add_7_25_groupi_g16301(csa_tree_add_7_25_groupi_n_4782 ,csa_tree_add_7_25_groupi_n_4736 ,csa_tree_add_7_25_groupi_n_4681);
  or csa_tree_add_7_25_groupi_g16302(csa_tree_add_7_25_groupi_n_4781 ,csa_tree_add_7_25_groupi_n_4736 ,csa_tree_add_7_25_groupi_n_4681);
  or csa_tree_add_7_25_groupi_g16303(csa_tree_add_7_25_groupi_n_4780 ,csa_tree_add_7_25_groupi_n_4744 ,csa_tree_add_7_25_groupi_n_4678);
  or csa_tree_add_7_25_groupi_g16304(csa_tree_add_7_25_groupi_n_4779 ,csa_tree_add_7_25_groupi_n_4743 ,csa_tree_add_7_25_groupi_n_4680);
  and csa_tree_add_7_25_groupi_g16305(csa_tree_add_7_25_groupi_n_4778 ,csa_tree_add_7_25_groupi_n_4743 ,csa_tree_add_7_25_groupi_n_4680);
  and csa_tree_add_7_25_groupi_g16306(csa_tree_add_7_25_groupi_n_4777 ,csa_tree_add_7_25_groupi_n_4744 ,csa_tree_add_7_25_groupi_n_4678);
  or csa_tree_add_7_25_groupi_g16307(csa_tree_add_7_25_groupi_n_4776 ,csa_tree_add_7_25_groupi_n_3036 ,csa_tree_add_7_25_groupi_n_4767);
  xnor csa_tree_add_7_25_groupi_g16308(out2[0] ,csa_tree_add_7_25_groupi_n_4691 ,csa_tree_add_7_25_groupi_n_4614);
  xnor csa_tree_add_7_25_groupi_g16309(csa_tree_add_7_25_groupi_n_4801 ,csa_tree_add_7_25_groupi_n_4689 ,csa_tree_add_7_25_groupi_n_4613);
  xnor csa_tree_add_7_25_groupi_g16310(csa_tree_add_7_25_groupi_n_4800 ,csa_tree_add_7_25_groupi_n_4690 ,csa_tree_add_7_25_groupi_n_4612);
  xnor csa_tree_add_7_25_groupi_g16311(csa_tree_add_7_25_groupi_n_4799 ,csa_tree_add_7_25_groupi_n_4687 ,csa_tree_add_7_25_groupi_n_4615);
  xnor csa_tree_add_7_25_groupi_g16312(csa_tree_add_7_25_groupi_n_4798 ,csa_tree_add_7_25_groupi_n_4688 ,csa_tree_add_7_25_groupi_n_4621);
  xnor csa_tree_add_7_25_groupi_g16313(csa_tree_add_7_25_groupi_n_4797 ,csa_tree_add_7_25_groupi_n_4715 ,csa_tree_add_7_25_groupi_n_4617);
  xnor csa_tree_add_7_25_groupi_g16314(csa_tree_add_7_25_groupi_n_4796 ,csa_tree_add_7_25_groupi_n_4713 ,csa_tree_add_7_25_groupi_n_4618);
  xnor csa_tree_add_7_25_groupi_g16315(csa_tree_add_7_25_groupi_n_4795 ,csa_tree_add_7_25_groupi_n_4714 ,csa_tree_add_7_25_groupi_n_4619);
  xnor csa_tree_add_7_25_groupi_g16316(csa_tree_add_7_25_groupi_n_4794 ,csa_tree_add_7_25_groupi_n_4717 ,csa_tree_add_7_25_groupi_n_4620);
  xnor csa_tree_add_7_25_groupi_g16317(csa_tree_add_7_25_groupi_n_4793 ,csa_tree_add_7_25_groupi_n_4686 ,csa_tree_add_7_25_groupi_n_4611);
  xnor csa_tree_add_7_25_groupi_g16318(csa_tree_add_7_25_groupi_n_4792 ,csa_tree_add_7_25_groupi_n_4716 ,csa_tree_add_7_25_groupi_n_2582);
  not csa_tree_add_7_25_groupi_g16319(csa_tree_add_7_25_groupi_n_4773 ,csa_tree_add_7_25_groupi_n_4774);
  not csa_tree_add_7_25_groupi_g16320(csa_tree_add_7_25_groupi_n_4772 ,csa_tree_add_7_25_groupi_n_4771);
  and csa_tree_add_7_25_groupi_g16321(csa_tree_add_7_25_groupi_n_4770 ,csa_tree_add_7_25_groupi_n_4594 ,csa_tree_add_7_25_groupi_n_4714);
  and csa_tree_add_7_25_groupi_g16322(csa_tree_add_7_25_groupi_n_4769 ,csa_tree_add_7_25_groupi_n_4591 ,csa_tree_add_7_25_groupi_n_4688);
  or csa_tree_add_7_25_groupi_g16323(csa_tree_add_7_25_groupi_n_4768 ,csa_tree_add_7_25_groupi_n_2438 ,csa_tree_add_7_25_groupi_n_4716);
  nor csa_tree_add_7_25_groupi_g16324(csa_tree_add_7_25_groupi_n_4767 ,csa_tree_add_7_25_groupi_n_309 ,csa_tree_add_7_25_groupi_n_2187);
  and csa_tree_add_7_25_groupi_g16325(csa_tree_add_7_25_groupi_n_4766 ,csa_tree_add_7_25_groupi_n_4596 ,csa_tree_add_7_25_groupi_n_4713);
  and csa_tree_add_7_25_groupi_g16326(csa_tree_add_7_25_groupi_n_4765 ,csa_tree_add_7_25_groupi_n_4597 ,csa_tree_add_7_25_groupi_n_4687);
  and csa_tree_add_7_25_groupi_g16327(csa_tree_add_7_25_groupi_n_4764 ,csa_tree_add_7_25_groupi_n_4593 ,csa_tree_add_7_25_groupi_n_4691);
  nor csa_tree_add_7_25_groupi_g16328(csa_tree_add_7_25_groupi_n_4763 ,csa_tree_add_7_25_groupi_n_555 ,csa_tree_add_7_25_groupi_n_1858);
  and csa_tree_add_7_25_groupi_g16329(csa_tree_add_7_25_groupi_n_4762 ,csa_tree_add_7_25_groupi_n_4595 ,csa_tree_add_7_25_groupi_n_4715);
  and csa_tree_add_7_25_groupi_g16330(csa_tree_add_7_25_groupi_n_4761 ,csa_tree_add_7_25_groupi_n_4586 ,csa_tree_add_7_25_groupi_n_4686);
  and csa_tree_add_7_25_groupi_g16331(csa_tree_add_7_25_groupi_n_4760 ,csa_tree_add_7_25_groupi_n_4584 ,csa_tree_add_7_25_groupi_n_4689);
  and csa_tree_add_7_25_groupi_g16332(csa_tree_add_7_25_groupi_n_4759 ,csa_tree_add_7_25_groupi_n_4585 ,csa_tree_add_7_25_groupi_n_4690);
  and csa_tree_add_7_25_groupi_g16333(csa_tree_add_7_25_groupi_n_4758 ,csa_tree_add_7_25_groupi_n_4571 ,csa_tree_add_7_25_groupi_n_4717);
  nor csa_tree_add_7_25_groupi_g16334(csa_tree_add_7_25_groupi_n_4757 ,csa_tree_add_7_25_groupi_n_638 ,csa_tree_add_7_25_groupi_n_150);
  nor csa_tree_add_7_25_groupi_g16335(csa_tree_add_7_25_groupi_n_4756 ,csa_tree_add_7_25_groupi_n_1859 ,csa_tree_add_7_25_groupi_n_1319);
  nor csa_tree_add_7_25_groupi_g16336(csa_tree_add_7_25_groupi_n_4755 ,csa_tree_add_7_25_groupi_n_4078 ,csa_tree_add_7_25_groupi_n_4672);
  nor csa_tree_add_7_25_groupi_g16337(csa_tree_add_7_25_groupi_n_4754 ,csa_tree_add_7_25_groupi_n_3835 ,csa_tree_add_7_25_groupi_n_4667);
  nor csa_tree_add_7_25_groupi_g16338(csa_tree_add_7_25_groupi_n_4753 ,csa_tree_add_7_25_groupi_n_4028 ,csa_tree_add_7_25_groupi_n_4671);
  nor csa_tree_add_7_25_groupi_g16339(csa_tree_add_7_25_groupi_n_4752 ,csa_tree_add_7_25_groupi_n_3833 ,csa_tree_add_7_25_groupi_n_4669);
  nor csa_tree_add_7_25_groupi_g16340(csa_tree_add_7_25_groupi_n_4751 ,csa_tree_add_7_25_groupi_n_3947 ,csa_tree_add_7_25_groupi_n_4675);
  nor csa_tree_add_7_25_groupi_g16341(csa_tree_add_7_25_groupi_n_4750 ,csa_tree_add_7_25_groupi_n_3848 ,csa_tree_add_7_25_groupi_n_4668);
  nor csa_tree_add_7_25_groupi_g16342(csa_tree_add_7_25_groupi_n_4749 ,csa_tree_add_7_25_groupi_n_4042 ,csa_tree_add_7_25_groupi_n_4673);
  nor csa_tree_add_7_25_groupi_g16343(csa_tree_add_7_25_groupi_n_4748 ,csa_tree_add_7_25_groupi_n_3477 ,csa_tree_add_7_25_groupi_n_4666);
  nor csa_tree_add_7_25_groupi_g16344(csa_tree_add_7_25_groupi_n_4747 ,csa_tree_add_7_25_groupi_n_4095 ,csa_tree_add_7_25_groupi_n_4674);
  nor csa_tree_add_7_25_groupi_g16345(csa_tree_add_7_25_groupi_n_4746 ,csa_tree_add_7_25_groupi_n_4041 ,csa_tree_add_7_25_groupi_n_4670);
  and csa_tree_add_7_25_groupi_g16346(csa_tree_add_7_25_groupi_n_4774 ,csa_tree_add_7_25_groupi_n_4561 ,csa_tree_add_7_25_groupi_n_4706);
  and csa_tree_add_7_25_groupi_g16347(csa_tree_add_7_25_groupi_n_4771 ,csa_tree_add_7_25_groupi_n_3837 ,csa_tree_add_7_25_groupi_n_4665);
  nor csa_tree_add_7_25_groupi_g16348(csa_tree_add_7_25_groupi_n_4735 ,csa_tree_add_7_25_groupi_n_309 ,csa_tree_add_7_25_groupi_n_2025);
  nor csa_tree_add_7_25_groupi_g16349(csa_tree_add_7_25_groupi_n_4734 ,csa_tree_add_7_25_groupi_n_333 ,csa_tree_add_7_25_groupi_n_2054);
  nor csa_tree_add_7_25_groupi_g16350(csa_tree_add_7_25_groupi_n_4733 ,csa_tree_add_7_25_groupi_n_332 ,csa_tree_add_7_25_groupi_n_2139);
  nor csa_tree_add_7_25_groupi_g16351(csa_tree_add_7_25_groupi_n_4732 ,csa_tree_add_7_25_groupi_n_308 ,csa_tree_add_7_25_groupi_n_2160);
  nor csa_tree_add_7_25_groupi_g16352(csa_tree_add_7_25_groupi_n_4731 ,csa_tree_add_7_25_groupi_n_2106 ,csa_tree_add_7_25_groupi_n_150);
  nor csa_tree_add_7_25_groupi_g16353(csa_tree_add_7_25_groupi_n_4730 ,csa_tree_add_7_25_groupi_n_333 ,csa_tree_add_7_25_groupi_n_2127);
  nor csa_tree_add_7_25_groupi_g16354(csa_tree_add_7_25_groupi_n_4729 ,csa_tree_add_7_25_groupi_n_2045 ,csa_tree_add_7_25_groupi_n_1859);
  xnor csa_tree_add_7_25_groupi_g16355(csa_tree_add_7_25_groupi_n_4728 ,csa_tree_add_7_25_groupi_n_4636 ,csa_tree_add_7_25_groupi_n_4406);
  xnor csa_tree_add_7_25_groupi_g16356(csa_tree_add_7_25_groupi_n_4727 ,csa_tree_add_7_25_groupi_n_4630 ,csa_tree_add_7_25_groupi_n_4575);
  xnor csa_tree_add_7_25_groupi_g16357(csa_tree_add_7_25_groupi_n_4726 ,csa_tree_add_7_25_groupi_n_4631 ,csa_tree_add_7_25_groupi_n_4582);
  xnor csa_tree_add_7_25_groupi_g16358(csa_tree_add_7_25_groupi_n_4725 ,csa_tree_add_7_25_groupi_n_4633 ,csa_tree_add_7_25_groupi_n_4574);
  xnor csa_tree_add_7_25_groupi_g16359(csa_tree_add_7_25_groupi_n_4724 ,csa_tree_add_7_25_groupi_n_4632 ,csa_tree_add_7_25_groupi_n_4581);
  xnor csa_tree_add_7_25_groupi_g16360(csa_tree_add_7_25_groupi_n_4723 ,csa_tree_add_7_25_groupi_n_4634 ,csa_tree_add_7_25_groupi_n_4580);
  xnor csa_tree_add_7_25_groupi_g16361(csa_tree_add_7_25_groupi_n_4722 ,csa_tree_add_7_25_groupi_n_4635 ,csa_tree_add_7_25_groupi_n_4579);
  xnor csa_tree_add_7_25_groupi_g16362(csa_tree_add_7_25_groupi_n_4721 ,csa_tree_add_7_25_groupi_n_4637 ,csa_tree_add_7_25_groupi_n_4578);
  xnor csa_tree_add_7_25_groupi_g16363(csa_tree_add_7_25_groupi_n_4720 ,csa_tree_add_7_25_groupi_n_4629 ,csa_tree_add_7_25_groupi_n_4577);
  xnor csa_tree_add_7_25_groupi_g16364(csa_tree_add_7_25_groupi_n_4719 ,csa_tree_add_7_25_groupi_n_4628 ,csa_tree_add_7_25_groupi_n_4576);
  xnor csa_tree_add_7_25_groupi_g16365(csa_tree_add_7_25_groupi_n_4718 ,csa_tree_add_7_25_groupi_n_4664 ,in3[5]);
  xnor csa_tree_add_7_25_groupi_g16366(csa_tree_add_7_25_groupi_n_4745 ,csa_tree_add_7_25_groupi_n_4647 ,in3[29]);
  xnor csa_tree_add_7_25_groupi_g16367(csa_tree_add_7_25_groupi_n_4744 ,csa_tree_add_7_25_groupi_n_4639 ,in3[5]);
  xnor csa_tree_add_7_25_groupi_g16368(csa_tree_add_7_25_groupi_n_4743 ,csa_tree_add_7_25_groupi_n_4642 ,in3[8]);
  xnor csa_tree_add_7_25_groupi_g16369(csa_tree_add_7_25_groupi_n_4742 ,csa_tree_add_7_25_groupi_n_4646 ,in3[2]);
  xnor csa_tree_add_7_25_groupi_g16370(csa_tree_add_7_25_groupi_n_4741 ,csa_tree_add_7_25_groupi_n_4641 ,in3[14]);
  xnor csa_tree_add_7_25_groupi_g16371(csa_tree_add_7_25_groupi_n_4740 ,csa_tree_add_7_25_groupi_n_4640 ,in3[17]);
  xnor csa_tree_add_7_25_groupi_g16372(csa_tree_add_7_25_groupi_n_4739 ,csa_tree_add_7_25_groupi_n_4643 ,in3[20]);
  xnor csa_tree_add_7_25_groupi_g16373(csa_tree_add_7_25_groupi_n_4738 ,csa_tree_add_7_25_groupi_n_4644 ,in3[23]);
  xnor csa_tree_add_7_25_groupi_g16374(csa_tree_add_7_25_groupi_n_4737 ,csa_tree_add_7_25_groupi_n_4645 ,in3[26]);
  xnor csa_tree_add_7_25_groupi_g16375(csa_tree_add_7_25_groupi_n_4736 ,csa_tree_add_7_25_groupi_n_4638 ,in3[11]);
  and csa_tree_add_7_25_groupi_g16376(csa_tree_add_7_25_groupi_n_4712 ,csa_tree_add_7_25_groupi_n_4637 ,csa_tree_add_7_25_groupi_n_4578);
  or csa_tree_add_7_25_groupi_g16377(csa_tree_add_7_25_groupi_n_4711 ,csa_tree_add_7_25_groupi_n_4628 ,csa_tree_add_7_25_groupi_n_4576);
  or csa_tree_add_7_25_groupi_g16378(csa_tree_add_7_25_groupi_n_4710 ,csa_tree_add_7_25_groupi_n_4632 ,csa_tree_add_7_25_groupi_n_4581);
  or csa_tree_add_7_25_groupi_g16379(csa_tree_add_7_25_groupi_n_4709 ,csa_tree_add_7_25_groupi_n_4629 ,csa_tree_add_7_25_groupi_n_4577);
  and csa_tree_add_7_25_groupi_g16380(csa_tree_add_7_25_groupi_n_4708 ,csa_tree_add_7_25_groupi_n_4628 ,csa_tree_add_7_25_groupi_n_4576);
  and csa_tree_add_7_25_groupi_g16381(csa_tree_add_7_25_groupi_n_4707 ,csa_tree_add_7_25_groupi_n_4632 ,csa_tree_add_7_25_groupi_n_4581);
  or csa_tree_add_7_25_groupi_g16382(csa_tree_add_7_25_groupi_n_4706 ,csa_tree_add_7_25_groupi_n_4562 ,csa_tree_add_7_25_groupi_n_4664);
  or csa_tree_add_7_25_groupi_g16383(csa_tree_add_7_25_groupi_n_4705 ,csa_tree_add_7_25_groupi_n_4633 ,csa_tree_add_7_25_groupi_n_4574);
  and csa_tree_add_7_25_groupi_g16384(csa_tree_add_7_25_groupi_n_4704 ,csa_tree_add_7_25_groupi_n_4629 ,csa_tree_add_7_25_groupi_n_4577);
  and csa_tree_add_7_25_groupi_g16385(csa_tree_add_7_25_groupi_n_4703 ,csa_tree_add_7_25_groupi_n_4636 ,csa_tree_add_7_25_groupi_n_4406);
  or csa_tree_add_7_25_groupi_g16386(csa_tree_add_7_25_groupi_n_4702 ,csa_tree_add_7_25_groupi_n_4636 ,csa_tree_add_7_25_groupi_n_4406);
  or csa_tree_add_7_25_groupi_g16387(csa_tree_add_7_25_groupi_n_4701 ,csa_tree_add_7_25_groupi_n_4634 ,csa_tree_add_7_25_groupi_n_4580);
  and csa_tree_add_7_25_groupi_g16388(csa_tree_add_7_25_groupi_n_4700 ,csa_tree_add_7_25_groupi_n_4633 ,csa_tree_add_7_25_groupi_n_4574);
  and csa_tree_add_7_25_groupi_g16389(csa_tree_add_7_25_groupi_n_4699 ,csa_tree_add_7_25_groupi_n_4634 ,csa_tree_add_7_25_groupi_n_4580);
  or csa_tree_add_7_25_groupi_g16390(csa_tree_add_7_25_groupi_n_4698 ,csa_tree_add_7_25_groupi_n_4637 ,csa_tree_add_7_25_groupi_n_4578);
  or csa_tree_add_7_25_groupi_g16391(csa_tree_add_7_25_groupi_n_4697 ,csa_tree_add_7_25_groupi_n_4635 ,csa_tree_add_7_25_groupi_n_4579);
  and csa_tree_add_7_25_groupi_g16392(csa_tree_add_7_25_groupi_n_4696 ,csa_tree_add_7_25_groupi_n_4630 ,csa_tree_add_7_25_groupi_n_4575);
  and csa_tree_add_7_25_groupi_g16393(csa_tree_add_7_25_groupi_n_4695 ,csa_tree_add_7_25_groupi_n_4631 ,csa_tree_add_7_25_groupi_n_4582);
  or csa_tree_add_7_25_groupi_g16394(csa_tree_add_7_25_groupi_n_4694 ,csa_tree_add_7_25_groupi_n_4630 ,csa_tree_add_7_25_groupi_n_4575);
  or csa_tree_add_7_25_groupi_g16395(csa_tree_add_7_25_groupi_n_4693 ,csa_tree_add_7_25_groupi_n_4631 ,csa_tree_add_7_25_groupi_n_4582);
  and csa_tree_add_7_25_groupi_g16396(csa_tree_add_7_25_groupi_n_4692 ,csa_tree_add_7_25_groupi_n_4635 ,csa_tree_add_7_25_groupi_n_4579);
  or csa_tree_add_7_25_groupi_g16397(csa_tree_add_7_25_groupi_n_4717 ,csa_tree_add_7_25_groupi_n_4475 ,csa_tree_add_7_25_groupi_n_4659);
  and csa_tree_add_7_25_groupi_g16398(csa_tree_add_7_25_groupi_n_4716 ,csa_tree_add_7_25_groupi_n_2435 ,csa_tree_add_7_25_groupi_n_4660);
  or csa_tree_add_7_25_groupi_g16399(csa_tree_add_7_25_groupi_n_4715 ,csa_tree_add_7_25_groupi_n_4473 ,csa_tree_add_7_25_groupi_n_4658);
  or csa_tree_add_7_25_groupi_g16400(csa_tree_add_7_25_groupi_n_4714 ,csa_tree_add_7_25_groupi_n_4481 ,csa_tree_add_7_25_groupi_n_4662);
  or csa_tree_add_7_25_groupi_g16401(csa_tree_add_7_25_groupi_n_4713 ,csa_tree_add_7_25_groupi_n_4477 ,csa_tree_add_7_25_groupi_n_4661);
  or csa_tree_add_7_25_groupi_g16402(csa_tree_add_7_25_groupi_n_4675 ,csa_tree_add_7_25_groupi_n_3581 ,csa_tree_add_7_25_groupi_n_4650);
  or csa_tree_add_7_25_groupi_g16403(csa_tree_add_7_25_groupi_n_4674 ,csa_tree_add_7_25_groupi_n_3154 ,csa_tree_add_7_25_groupi_n_4626);
  or csa_tree_add_7_25_groupi_g16404(csa_tree_add_7_25_groupi_n_4673 ,csa_tree_add_7_25_groupi_n_3144 ,csa_tree_add_7_25_groupi_n_4625);
  or csa_tree_add_7_25_groupi_g16405(csa_tree_add_7_25_groupi_n_4672 ,csa_tree_add_7_25_groupi_n_3120 ,csa_tree_add_7_25_groupi_n_4623);
  or csa_tree_add_7_25_groupi_g16406(csa_tree_add_7_25_groupi_n_4671 ,csa_tree_add_7_25_groupi_n_3126 ,csa_tree_add_7_25_groupi_n_4624);
  or csa_tree_add_7_25_groupi_g16407(csa_tree_add_7_25_groupi_n_4670 ,csa_tree_add_7_25_groupi_n_3115 ,csa_tree_add_7_25_groupi_n_4622);
  or csa_tree_add_7_25_groupi_g16408(csa_tree_add_7_25_groupi_n_4669 ,csa_tree_add_7_25_groupi_n_3636 ,csa_tree_add_7_25_groupi_n_4663);
  or csa_tree_add_7_25_groupi_g16409(csa_tree_add_7_25_groupi_n_4668 ,csa_tree_add_7_25_groupi_n_3564 ,csa_tree_add_7_25_groupi_n_4648);
  or csa_tree_add_7_25_groupi_g16410(csa_tree_add_7_25_groupi_n_4667 ,csa_tree_add_7_25_groupi_n_3565 ,csa_tree_add_7_25_groupi_n_4627);
  or csa_tree_add_7_25_groupi_g16411(csa_tree_add_7_25_groupi_n_4666 ,csa_tree_add_7_25_groupi_n_2919 ,csa_tree_add_7_25_groupi_n_4649);
  nor csa_tree_add_7_25_groupi_g16412(csa_tree_add_7_25_groupi_n_4665 ,csa_tree_add_7_25_groupi_n_2990 ,csa_tree_add_7_25_groupi_n_4651);
  or csa_tree_add_7_25_groupi_g16413(csa_tree_add_7_25_groupi_n_4691 ,csa_tree_add_7_25_groupi_n_4544 ,csa_tree_add_7_25_groupi_n_4657);
  or csa_tree_add_7_25_groupi_g16414(csa_tree_add_7_25_groupi_n_4690 ,csa_tree_add_7_25_groupi_n_4447 ,csa_tree_add_7_25_groupi_n_4655);
  or csa_tree_add_7_25_groupi_g16415(csa_tree_add_7_25_groupi_n_4689 ,csa_tree_add_7_25_groupi_n_4448 ,csa_tree_add_7_25_groupi_n_4653);
  or csa_tree_add_7_25_groupi_g16416(csa_tree_add_7_25_groupi_n_4688 ,csa_tree_add_7_25_groupi_n_4456 ,csa_tree_add_7_25_groupi_n_4652);
  or csa_tree_add_7_25_groupi_g16417(csa_tree_add_7_25_groupi_n_4687 ,csa_tree_add_7_25_groupi_n_4454 ,csa_tree_add_7_25_groupi_n_4656);
  or csa_tree_add_7_25_groupi_g16418(csa_tree_add_7_25_groupi_n_4686 ,csa_tree_add_7_25_groupi_n_4451 ,csa_tree_add_7_25_groupi_n_4654);
  xnor csa_tree_add_7_25_groupi_g16419(csa_tree_add_7_25_groupi_n_4685 ,csa_tree_add_7_25_groupi_n_4602 ,csa_tree_add_7_25_groupi_n_4509);
  xnor csa_tree_add_7_25_groupi_g16420(csa_tree_add_7_25_groupi_n_4684 ,csa_tree_add_7_25_groupi_n_4608 ,csa_tree_add_7_25_groupi_n_4506);
  xnor csa_tree_add_7_25_groupi_g16421(csa_tree_add_7_25_groupi_n_4683 ,csa_tree_add_7_25_groupi_n_4609 ,csa_tree_add_7_25_groupi_n_4508);
  xnor csa_tree_add_7_25_groupi_g16422(csa_tree_add_7_25_groupi_n_4682 ,csa_tree_add_7_25_groupi_n_4607 ,csa_tree_add_7_25_groupi_n_4502);
  xnor csa_tree_add_7_25_groupi_g16423(csa_tree_add_7_25_groupi_n_4681 ,csa_tree_add_7_25_groupi_n_4601 ,csa_tree_add_7_25_groupi_n_4503);
  xnor csa_tree_add_7_25_groupi_g16424(csa_tree_add_7_25_groupi_n_4680 ,csa_tree_add_7_25_groupi_n_4605 ,csa_tree_add_7_25_groupi_n_4499);
  xnor csa_tree_add_7_25_groupi_g16425(csa_tree_add_7_25_groupi_n_4679 ,csa_tree_add_7_25_groupi_n_4604 ,csa_tree_add_7_25_groupi_n_4501);
  xnor csa_tree_add_7_25_groupi_g16426(csa_tree_add_7_25_groupi_n_4678 ,csa_tree_add_7_25_groupi_n_4603 ,csa_tree_add_7_25_groupi_n_4500);
  xnor csa_tree_add_7_25_groupi_g16427(csa_tree_add_7_25_groupi_n_4677 ,csa_tree_add_7_25_groupi_n_4606 ,csa_tree_add_7_25_groupi_n_4507);
  xnor csa_tree_add_7_25_groupi_g16428(csa_tree_add_7_25_groupi_n_4676 ,csa_tree_add_7_25_groupi_n_4610 ,csa_tree_add_7_25_groupi_n_2576);
  nor csa_tree_add_7_25_groupi_g16429(csa_tree_add_7_25_groupi_n_4663 ,csa_tree_add_7_25_groupi_n_741 ,csa_tree_add_7_25_groupi_n_271);
  and csa_tree_add_7_25_groupi_g16430(csa_tree_add_7_25_groupi_n_4662 ,csa_tree_add_7_25_groupi_n_4488 ,csa_tree_add_7_25_groupi_n_4608);
  and csa_tree_add_7_25_groupi_g16431(csa_tree_add_7_25_groupi_n_4661 ,csa_tree_add_7_25_groupi_n_4472 ,csa_tree_add_7_25_groupi_n_4606);
  or csa_tree_add_7_25_groupi_g16432(csa_tree_add_7_25_groupi_n_4660 ,csa_tree_add_7_25_groupi_n_2451 ,csa_tree_add_7_25_groupi_n_4610);
  and csa_tree_add_7_25_groupi_g16433(csa_tree_add_7_25_groupi_n_4659 ,csa_tree_add_7_25_groupi_n_4474 ,csa_tree_add_7_25_groupi_n_4602);
  and csa_tree_add_7_25_groupi_g16434(csa_tree_add_7_25_groupi_n_4658 ,csa_tree_add_7_25_groupi_n_4484 ,csa_tree_add_7_25_groupi_n_4609);
  nor csa_tree_add_7_25_groupi_g16435(csa_tree_add_7_25_groupi_n_4657 ,csa_tree_add_7_25_groupi_n_4545 ,csa_tree_add_7_25_groupi_n_4590);
  and csa_tree_add_7_25_groupi_g16436(csa_tree_add_7_25_groupi_n_4656 ,csa_tree_add_7_25_groupi_n_4453 ,csa_tree_add_7_25_groupi_n_4601);
  and csa_tree_add_7_25_groupi_g16437(csa_tree_add_7_25_groupi_n_4655 ,csa_tree_add_7_25_groupi_n_4450 ,csa_tree_add_7_25_groupi_n_4603);
  and csa_tree_add_7_25_groupi_g16438(csa_tree_add_7_25_groupi_n_4654 ,csa_tree_add_7_25_groupi_n_4452 ,csa_tree_add_7_25_groupi_n_4605);
  and csa_tree_add_7_25_groupi_g16439(csa_tree_add_7_25_groupi_n_4653 ,csa_tree_add_7_25_groupi_n_4449 ,csa_tree_add_7_25_groupi_n_4604);
  and csa_tree_add_7_25_groupi_g16440(csa_tree_add_7_25_groupi_n_4652 ,csa_tree_add_7_25_groupi_n_4455 ,csa_tree_add_7_25_groupi_n_4607);
  nor csa_tree_add_7_25_groupi_g16441(csa_tree_add_7_25_groupi_n_4651 ,csa_tree_add_7_25_groupi_n_551 ,csa_tree_add_7_25_groupi_n_1821);
  nor csa_tree_add_7_25_groupi_g16442(csa_tree_add_7_25_groupi_n_4650 ,csa_tree_add_7_25_groupi_n_1917 ,csa_tree_add_7_25_groupi_n_174);
  nor csa_tree_add_7_25_groupi_g16443(csa_tree_add_7_25_groupi_n_4649 ,csa_tree_add_7_25_groupi_n_2169 ,csa_tree_add_7_25_groupi_n_1822);
  nor csa_tree_add_7_25_groupi_g16444(csa_tree_add_7_25_groupi_n_4648 ,csa_tree_add_7_25_groupi_n_320 ,csa_tree_add_7_25_groupi_n_2028);
  nor csa_tree_add_7_25_groupi_g16445(csa_tree_add_7_25_groupi_n_4647 ,csa_tree_add_7_25_groupi_n_3830 ,csa_tree_add_7_25_groupi_n_4569);
  nor csa_tree_add_7_25_groupi_g16446(csa_tree_add_7_25_groupi_n_4646 ,csa_tree_add_7_25_groupi_n_3476 ,csa_tree_add_7_25_groupi_n_4558);
  nor csa_tree_add_7_25_groupi_g16447(csa_tree_add_7_25_groupi_n_4645 ,csa_tree_add_7_25_groupi_n_3938 ,csa_tree_add_7_25_groupi_n_4563);
  nor csa_tree_add_7_25_groupi_g16448(csa_tree_add_7_25_groupi_n_4644 ,csa_tree_add_7_25_groupi_n_3931 ,csa_tree_add_7_25_groupi_n_4560);
  nor csa_tree_add_7_25_groupi_g16449(csa_tree_add_7_25_groupi_n_4643 ,csa_tree_add_7_25_groupi_n_4090 ,csa_tree_add_7_25_groupi_n_4570);
  nor csa_tree_add_7_25_groupi_g16450(csa_tree_add_7_25_groupi_n_4642 ,csa_tree_add_7_25_groupi_n_4043 ,csa_tree_add_7_25_groupi_n_4566);
  nor csa_tree_add_7_25_groupi_g16451(csa_tree_add_7_25_groupi_n_4641 ,csa_tree_add_7_25_groupi_n_4044 ,csa_tree_add_7_25_groupi_n_4565);
  nor csa_tree_add_7_25_groupi_g16452(csa_tree_add_7_25_groupi_n_4640 ,csa_tree_add_7_25_groupi_n_4079 ,csa_tree_add_7_25_groupi_n_4568);
  nor csa_tree_add_7_25_groupi_g16453(csa_tree_add_7_25_groupi_n_4639 ,csa_tree_add_7_25_groupi_n_3992 ,csa_tree_add_7_25_groupi_n_4567);
  nor csa_tree_add_7_25_groupi_g16454(csa_tree_add_7_25_groupi_n_4638 ,csa_tree_add_7_25_groupi_n_4047 ,csa_tree_add_7_25_groupi_n_4564);
  and csa_tree_add_7_25_groupi_g16455(csa_tree_add_7_25_groupi_n_4664 ,csa_tree_add_7_25_groupi_n_3933 ,csa_tree_add_7_25_groupi_n_4559);
  nor csa_tree_add_7_25_groupi_g16456(csa_tree_add_7_25_groupi_n_4627 ,csa_tree_add_7_25_groupi_n_271 ,csa_tree_add_7_25_groupi_n_2043);
  nor csa_tree_add_7_25_groupi_g16457(csa_tree_add_7_25_groupi_n_4626 ,csa_tree_add_7_25_groupi_n_321 ,csa_tree_add_7_25_groupi_n_2058);
  nor csa_tree_add_7_25_groupi_g16458(csa_tree_add_7_25_groupi_n_4625 ,csa_tree_add_7_25_groupi_n_270 ,csa_tree_add_7_25_groupi_n_2166);
  nor csa_tree_add_7_25_groupi_g16459(csa_tree_add_7_25_groupi_n_4624 ,csa_tree_add_7_25_groupi_n_2091 ,csa_tree_add_7_25_groupi_n_1821);
  nor csa_tree_add_7_25_groupi_g16460(csa_tree_add_7_25_groupi_n_4623 ,csa_tree_add_7_25_groupi_n_321 ,csa_tree_add_7_25_groupi_n_2145);
  nor csa_tree_add_7_25_groupi_g16461(csa_tree_add_7_25_groupi_n_4622 ,csa_tree_add_7_25_groupi_n_2112 ,csa_tree_add_7_25_groupi_n_174);
  xnor csa_tree_add_7_25_groupi_g16462(csa_tree_add_7_25_groupi_n_4621 ,csa_tree_add_7_25_groupi_n_4521 ,csa_tree_add_7_25_groupi_n_4466);
  xnor csa_tree_add_7_25_groupi_g16463(csa_tree_add_7_25_groupi_n_4620 ,csa_tree_add_7_25_groupi_n_4517 ,csa_tree_add_7_25_groupi_n_4352);
  xnor csa_tree_add_7_25_groupi_g16464(csa_tree_add_7_25_groupi_n_4619 ,csa_tree_add_7_25_groupi_n_4518 ,csa_tree_add_7_25_groupi_n_4463);
  xnor csa_tree_add_7_25_groupi_g16465(csa_tree_add_7_25_groupi_n_4618 ,csa_tree_add_7_25_groupi_n_4519 ,csa_tree_add_7_25_groupi_n_4464);
  xnor csa_tree_add_7_25_groupi_g16466(csa_tree_add_7_25_groupi_n_4617 ,csa_tree_add_7_25_groupi_n_4520 ,csa_tree_add_7_25_groupi_n_4465);
  xnor csa_tree_add_7_25_groupi_g16467(csa_tree_add_7_25_groupi_n_4616 ,csa_tree_add_7_25_groupi_n_1094 ,csa_tree_add_7_25_groupi_n_1109);
  xnor csa_tree_add_7_25_groupi_g16468(csa_tree_add_7_25_groupi_n_4615 ,csa_tree_add_7_25_groupi_n_4522 ,csa_tree_add_7_25_groupi_n_4467);
  xnor csa_tree_add_7_25_groupi_g16469(csa_tree_add_7_25_groupi_n_4614 ,csa_tree_add_7_25_groupi_n_4523 ,csa_tree_add_7_25_groupi_n_4468);
  xnor csa_tree_add_7_25_groupi_g16470(csa_tree_add_7_25_groupi_n_4613 ,csa_tree_add_7_25_groupi_n_4526 ,csa_tree_add_7_25_groupi_n_4461);
  xnor csa_tree_add_7_25_groupi_g16471(csa_tree_add_7_25_groupi_n_4612 ,csa_tree_add_7_25_groupi_n_4525 ,csa_tree_add_7_25_groupi_n_4469);
  xnor csa_tree_add_7_25_groupi_g16472(csa_tree_add_7_25_groupi_n_4611 ,csa_tree_add_7_25_groupi_n_4524 ,csa_tree_add_7_25_groupi_n_4462);
  xnor csa_tree_add_7_25_groupi_g16473(csa_tree_add_7_25_groupi_n_4637 ,csa_tree_add_7_25_groupi_n_4531 ,in3[20]);
  xnor csa_tree_add_7_25_groupi_g16474(csa_tree_add_7_25_groupi_n_4636 ,csa_tree_add_7_25_groupi_n_4533 ,in3[29]);
  xnor csa_tree_add_7_25_groupi_g16475(csa_tree_add_7_25_groupi_n_4635 ,csa_tree_add_7_25_groupi_n_4530 ,in3[17]);
  xnor csa_tree_add_7_25_groupi_g16476(csa_tree_add_7_25_groupi_n_4634 ,csa_tree_add_7_25_groupi_n_4528 ,in3[14]);
  xnor csa_tree_add_7_25_groupi_g16477(csa_tree_add_7_25_groupi_n_4633 ,csa_tree_add_7_25_groupi_n_4535 ,in3[2]);
  xnor csa_tree_add_7_25_groupi_g16478(csa_tree_add_7_25_groupi_n_4632 ,csa_tree_add_7_25_groupi_n_4534 ,in3[11]);
  xnor csa_tree_add_7_25_groupi_g16479(csa_tree_add_7_25_groupi_n_4631 ,csa_tree_add_7_25_groupi_n_4536 ,in3[8]);
  xnor csa_tree_add_7_25_groupi_g16480(csa_tree_add_7_25_groupi_n_4630 ,csa_tree_add_7_25_groupi_n_4527 ,in3[5]);
  xnor csa_tree_add_7_25_groupi_g16481(csa_tree_add_7_25_groupi_n_4629 ,csa_tree_add_7_25_groupi_n_4532 ,in3[23]);
  xnor csa_tree_add_7_25_groupi_g16482(csa_tree_add_7_25_groupi_n_4628 ,csa_tree_add_7_25_groupi_n_4529 ,in3[26]);
  and csa_tree_add_7_25_groupi_g16483(csa_tree_add_7_25_groupi_n_4600 ,csa_tree_add_7_25_groupi_n_4519 ,csa_tree_add_7_25_groupi_n_4464);
  and csa_tree_add_7_25_groupi_g16484(csa_tree_add_7_25_groupi_n_4599 ,csa_tree_add_7_25_groupi_n_4518 ,csa_tree_add_7_25_groupi_n_4463);
  and csa_tree_add_7_25_groupi_g16485(csa_tree_add_7_25_groupi_n_4598 ,csa_tree_add_7_25_groupi_n_4522 ,csa_tree_add_7_25_groupi_n_4467);
  or csa_tree_add_7_25_groupi_g16486(csa_tree_add_7_25_groupi_n_4597 ,csa_tree_add_7_25_groupi_n_4522 ,csa_tree_add_7_25_groupi_n_4467);
  or csa_tree_add_7_25_groupi_g16487(csa_tree_add_7_25_groupi_n_4596 ,csa_tree_add_7_25_groupi_n_4519 ,csa_tree_add_7_25_groupi_n_4464);
  or csa_tree_add_7_25_groupi_g16488(csa_tree_add_7_25_groupi_n_4595 ,csa_tree_add_7_25_groupi_n_4520 ,csa_tree_add_7_25_groupi_n_4465);
  or csa_tree_add_7_25_groupi_g16489(csa_tree_add_7_25_groupi_n_4594 ,csa_tree_add_7_25_groupi_n_4518 ,csa_tree_add_7_25_groupi_n_4463);
  or csa_tree_add_7_25_groupi_g16490(csa_tree_add_7_25_groupi_n_4593 ,csa_tree_add_7_25_groupi_n_4523 ,csa_tree_add_7_25_groupi_n_4468);
  and csa_tree_add_7_25_groupi_g16491(csa_tree_add_7_25_groupi_n_4592 ,csa_tree_add_7_25_groupi_n_4523 ,csa_tree_add_7_25_groupi_n_4468);
  or csa_tree_add_7_25_groupi_g16492(csa_tree_add_7_25_groupi_n_4591 ,csa_tree_add_7_25_groupi_n_4521 ,csa_tree_add_7_25_groupi_n_4466);
  nor csa_tree_add_7_25_groupi_g16493(csa_tree_add_7_25_groupi_n_4590 ,csa_tree_add_7_25_groupi_n_4365 ,csa_tree_add_7_25_groupi_n_4539);
  and csa_tree_add_7_25_groupi_g16494(csa_tree_add_7_25_groupi_n_4589 ,csa_tree_add_7_25_groupi_n_4520 ,csa_tree_add_7_25_groupi_n_4465);
  and csa_tree_add_7_25_groupi_g16495(csa_tree_add_7_25_groupi_n_4588 ,csa_tree_add_7_25_groupi_n_4525 ,csa_tree_add_7_25_groupi_n_4469);
  and csa_tree_add_7_25_groupi_g16496(csa_tree_add_7_25_groupi_n_4587 ,csa_tree_add_7_25_groupi_n_4524 ,csa_tree_add_7_25_groupi_n_4462);
  or csa_tree_add_7_25_groupi_g16497(csa_tree_add_7_25_groupi_n_4586 ,csa_tree_add_7_25_groupi_n_4524 ,csa_tree_add_7_25_groupi_n_4462);
  or csa_tree_add_7_25_groupi_g16498(csa_tree_add_7_25_groupi_n_4585 ,csa_tree_add_7_25_groupi_n_4525 ,csa_tree_add_7_25_groupi_n_4469);
  or csa_tree_add_7_25_groupi_g16499(csa_tree_add_7_25_groupi_n_4584 ,csa_tree_add_7_25_groupi_n_4526 ,csa_tree_add_7_25_groupi_n_4461);
  and csa_tree_add_7_25_groupi_g16500(csa_tree_add_7_25_groupi_n_4583 ,csa_tree_add_7_25_groupi_n_4521 ,csa_tree_add_7_25_groupi_n_4466);
  and csa_tree_add_7_25_groupi_g16501(csa_tree_add_7_25_groupi_n_4610 ,csa_tree_add_7_25_groupi_n_2487 ,csa_tree_add_7_25_groupi_n_4547);
  or csa_tree_add_7_25_groupi_g16502(csa_tree_add_7_25_groupi_n_4609 ,csa_tree_add_7_25_groupi_n_4364 ,csa_tree_add_7_25_groupi_n_4537);
  or csa_tree_add_7_25_groupi_g16503(csa_tree_add_7_25_groupi_n_4608 ,csa_tree_add_7_25_groupi_n_4366 ,csa_tree_add_7_25_groupi_n_4546);
  or csa_tree_add_7_25_groupi_g16504(csa_tree_add_7_25_groupi_n_4607 ,csa_tree_add_7_25_groupi_n_4357 ,csa_tree_add_7_25_groupi_n_4551);
  or csa_tree_add_7_25_groupi_g16505(csa_tree_add_7_25_groupi_n_4606 ,csa_tree_add_7_25_groupi_n_4358 ,csa_tree_add_7_25_groupi_n_4543);
  or csa_tree_add_7_25_groupi_g16506(csa_tree_add_7_25_groupi_n_4605 ,csa_tree_add_7_25_groupi_n_4346 ,csa_tree_add_7_25_groupi_n_4540);
  or csa_tree_add_7_25_groupi_g16507(csa_tree_add_7_25_groupi_n_4604 ,csa_tree_add_7_25_groupi_n_4336 ,csa_tree_add_7_25_groupi_n_4542);
  or csa_tree_add_7_25_groupi_g16508(csa_tree_add_7_25_groupi_n_4603 ,csa_tree_add_7_25_groupi_n_4345 ,csa_tree_add_7_25_groupi_n_4541);
  or csa_tree_add_7_25_groupi_g16509(csa_tree_add_7_25_groupi_n_4602 ,csa_tree_add_7_25_groupi_n_4353 ,csa_tree_add_7_25_groupi_n_4538);
  or csa_tree_add_7_25_groupi_g16510(csa_tree_add_7_25_groupi_n_4601 ,csa_tree_add_7_25_groupi_n_4363 ,csa_tree_add_7_25_groupi_n_4549);
  and csa_tree_add_7_25_groupi_g16511(csa_tree_add_7_25_groupi_n_4572 ,csa_tree_add_7_25_groupi_n_4517 ,csa_tree_add_7_25_groupi_n_4352);
  or csa_tree_add_7_25_groupi_g16512(csa_tree_add_7_25_groupi_n_4571 ,csa_tree_add_7_25_groupi_n_4517 ,csa_tree_add_7_25_groupi_n_4352);
  or csa_tree_add_7_25_groupi_g16513(csa_tree_add_7_25_groupi_n_4570 ,csa_tree_add_7_25_groupi_n_3174 ,csa_tree_add_7_25_groupi_n_4510);
  or csa_tree_add_7_25_groupi_g16514(csa_tree_add_7_25_groupi_n_4569 ,csa_tree_add_7_25_groupi_n_3653 ,csa_tree_add_7_25_groupi_n_4550);
  or csa_tree_add_7_25_groupi_g16515(csa_tree_add_7_25_groupi_n_4568 ,csa_tree_add_7_25_groupi_n_3153 ,csa_tree_add_7_25_groupi_n_4515);
  or csa_tree_add_7_25_groupi_g16516(csa_tree_add_7_25_groupi_n_4567 ,csa_tree_add_7_25_groupi_n_3133 ,csa_tree_add_7_25_groupi_n_4514);
  or csa_tree_add_7_25_groupi_g16517(csa_tree_add_7_25_groupi_n_4566 ,csa_tree_add_7_25_groupi_n_3123 ,csa_tree_add_7_25_groupi_n_4511);
  or csa_tree_add_7_25_groupi_g16518(csa_tree_add_7_25_groupi_n_4565 ,csa_tree_add_7_25_groupi_n_3125 ,csa_tree_add_7_25_groupi_n_4513);
  or csa_tree_add_7_25_groupi_g16519(csa_tree_add_7_25_groupi_n_4564 ,csa_tree_add_7_25_groupi_n_3131 ,csa_tree_add_7_25_groupi_n_4512);
  or csa_tree_add_7_25_groupi_g16520(csa_tree_add_7_25_groupi_n_4563 ,csa_tree_add_7_25_groupi_n_3572 ,csa_tree_add_7_25_groupi_n_4553);
  and csa_tree_add_7_25_groupi_g16521(csa_tree_add_7_25_groupi_n_4562 ,in3[5] ,csa_tree_add_7_25_groupi_n_1100);
  or csa_tree_add_7_25_groupi_g16522(csa_tree_add_7_25_groupi_n_4561 ,in3[5] ,csa_tree_add_7_25_groupi_n_1109);
  or csa_tree_add_7_25_groupi_g16523(csa_tree_add_7_25_groupi_n_4560 ,csa_tree_add_7_25_groupi_n_3646 ,csa_tree_add_7_25_groupi_n_4516);
  nor csa_tree_add_7_25_groupi_g16524(csa_tree_add_7_25_groupi_n_4559 ,csa_tree_add_7_25_groupi_n_2968 ,csa_tree_add_7_25_groupi_n_4548);
  or csa_tree_add_7_25_groupi_g16525(csa_tree_add_7_25_groupi_n_4558 ,csa_tree_add_7_25_groupi_n_2941 ,csa_tree_add_7_25_groupi_n_4552);
  nor csa_tree_add_7_25_groupi_g16526(csa_tree_add_7_25_groupi_n_4557 ,csa_tree_add_7_25_groupi_n_4442 ,csa_tree_add_7_25_groupi_n_2343);
  or csa_tree_add_7_25_groupi_g16527(csa_tree_add_7_25_groupi_n_4556 ,csa_tree_add_7_25_groupi_n_2342 ,csa_tree_add_7_25_groupi_n_1100);
  and csa_tree_add_7_25_groupi_g16528(csa_tree_add_7_25_groupi_n_4555 ,csa_tree_add_7_25_groupi_n_4526 ,csa_tree_add_7_25_groupi_n_4461);
  xnor csa_tree_add_7_25_groupi_g16529(csa_tree_add_7_25_groupi_n_4582 ,csa_tree_add_7_25_groupi_n_4496 ,csa_tree_add_7_25_groupi_n_4384);
  xnor csa_tree_add_7_25_groupi_g16530(csa_tree_add_7_25_groupi_n_4581 ,csa_tree_add_7_25_groupi_n_4492 ,csa_tree_add_7_25_groupi_n_4385);
  xnor csa_tree_add_7_25_groupi_g16531(csa_tree_add_7_25_groupi_n_4580 ,csa_tree_add_7_25_groupi_n_4489 ,csa_tree_add_7_25_groupi_n_4386);
  xnor csa_tree_add_7_25_groupi_g16532(csa_tree_add_7_25_groupi_n_4579 ,csa_tree_add_7_25_groupi_n_4498 ,csa_tree_add_7_25_groupi_n_4387);
  xnor csa_tree_add_7_25_groupi_g16533(csa_tree_add_7_25_groupi_n_4578 ,csa_tree_add_7_25_groupi_n_4490 ,csa_tree_add_7_25_groupi_n_4388);
  xnor csa_tree_add_7_25_groupi_g16534(csa_tree_add_7_25_groupi_n_4577 ,csa_tree_add_7_25_groupi_n_4493 ,csa_tree_add_7_25_groupi_n_4389);
  xnor csa_tree_add_7_25_groupi_g16535(csa_tree_add_7_25_groupi_n_4576 ,csa_tree_add_7_25_groupi_n_4497 ,csa_tree_add_7_25_groupi_n_4381);
  xnor csa_tree_add_7_25_groupi_g16536(csa_tree_add_7_25_groupi_n_4575 ,csa_tree_add_7_25_groupi_n_4494 ,csa_tree_add_7_25_groupi_n_4383);
  xnor csa_tree_add_7_25_groupi_g16537(csa_tree_add_7_25_groupi_n_4574 ,csa_tree_add_7_25_groupi_n_4495 ,csa_tree_add_7_25_groupi_n_4382);
  xnor csa_tree_add_7_25_groupi_g16538(csa_tree_add_7_25_groupi_n_4573 ,csa_tree_add_7_25_groupi_n_4491 ,csa_tree_add_7_25_groupi_n_2587);
  nor csa_tree_add_7_25_groupi_g16540(csa_tree_add_7_25_groupi_n_4553 ,csa_tree_add_7_25_groupi_n_741 ,csa_tree_add_7_25_groupi_n_258);
  nor csa_tree_add_7_25_groupi_g16541(csa_tree_add_7_25_groupi_n_4552 ,csa_tree_add_7_25_groupi_n_2085 ,csa_tree_add_7_25_groupi_n_157);
  and csa_tree_add_7_25_groupi_g16542(csa_tree_add_7_25_groupi_n_4551 ,csa_tree_add_7_25_groupi_n_4367 ,csa_tree_add_7_25_groupi_n_4489);
  nor csa_tree_add_7_25_groupi_g16543(csa_tree_add_7_25_groupi_n_4550 ,csa_tree_add_7_25_groupi_n_266 ,csa_tree_add_7_25_groupi_n_1842);
  and csa_tree_add_7_25_groupi_g16544(csa_tree_add_7_25_groupi_n_4549 ,csa_tree_add_7_25_groupi_n_4359 ,csa_tree_add_7_25_groupi_n_4492);
  nor csa_tree_add_7_25_groupi_g16545(csa_tree_add_7_25_groupi_n_4548 ,csa_tree_add_7_25_groupi_n_552 ,csa_tree_add_7_25_groupi_n_157);
  or csa_tree_add_7_25_groupi_g16546(csa_tree_add_7_25_groupi_n_4547 ,csa_tree_add_7_25_groupi_n_2444 ,csa_tree_add_7_25_groupi_n_4491);
  and csa_tree_add_7_25_groupi_g16547(csa_tree_add_7_25_groupi_n_4546 ,csa_tree_add_7_25_groupi_n_4362 ,csa_tree_add_7_25_groupi_n_4493);
  nor csa_tree_add_7_25_groupi_g16548(csa_tree_add_7_25_groupi_n_4545 ,csa_tree_add_7_25_groupi_n_4411 ,csa_tree_add_7_25_groupi_n_4471);
  nor csa_tree_add_7_25_groupi_g16549(csa_tree_add_7_25_groupi_n_4544 ,csa_tree_add_7_25_groupi_n_4412 ,csa_tree_add_7_25_groupi_n_4470);
  and csa_tree_add_7_25_groupi_g16550(csa_tree_add_7_25_groupi_n_4543 ,csa_tree_add_7_25_groupi_n_4360 ,csa_tree_add_7_25_groupi_n_4490);
  and csa_tree_add_7_25_groupi_g16551(csa_tree_add_7_25_groupi_n_4542 ,csa_tree_add_7_25_groupi_n_4348 ,csa_tree_add_7_25_groupi_n_4495);
  and csa_tree_add_7_25_groupi_g16552(csa_tree_add_7_25_groupi_n_4541 ,csa_tree_add_7_25_groupi_n_4349 ,csa_tree_add_7_25_groupi_n_4494);
  and csa_tree_add_7_25_groupi_g16553(csa_tree_add_7_25_groupi_n_4540 ,csa_tree_add_7_25_groupi_n_4347 ,csa_tree_add_7_25_groupi_n_4496);
  nor csa_tree_add_7_25_groupi_g16554(csa_tree_add_7_25_groupi_n_4539 ,csa_tree_add_7_25_groupi_n_4354 ,csa_tree_add_7_25_groupi_n_4478);
  and csa_tree_add_7_25_groupi_g16555(csa_tree_add_7_25_groupi_n_4538 ,csa_tree_add_7_25_groupi_n_4355 ,csa_tree_add_7_25_groupi_n_4497);
  and csa_tree_add_7_25_groupi_g16556(csa_tree_add_7_25_groupi_n_4537 ,csa_tree_add_7_25_groupi_n_4361 ,csa_tree_add_7_25_groupi_n_4498);
  nor csa_tree_add_7_25_groupi_g16557(csa_tree_add_7_25_groupi_n_4536 ,csa_tree_add_7_25_groupi_n_4037 ,csa_tree_add_7_25_groupi_n_4458);
  nor csa_tree_add_7_25_groupi_g16558(csa_tree_add_7_25_groupi_n_4535 ,csa_tree_add_7_25_groupi_n_3463 ,csa_tree_add_7_25_groupi_n_4446);
  nor csa_tree_add_7_25_groupi_g16559(csa_tree_add_7_25_groupi_n_4534 ,csa_tree_add_7_25_groupi_n_4023 ,csa_tree_add_7_25_groupi_n_4443);
  nor csa_tree_add_7_25_groupi_g16560(csa_tree_add_7_25_groupi_n_4533 ,csa_tree_add_7_25_groupi_n_3885 ,csa_tree_add_7_25_groupi_n_4485);
  nor csa_tree_add_7_25_groupi_g16561(csa_tree_add_7_25_groupi_n_4532 ,csa_tree_add_7_25_groupi_n_4007 ,csa_tree_add_7_25_groupi_n_4482);
  nor csa_tree_add_7_25_groupi_g16562(csa_tree_add_7_25_groupi_n_4531 ,csa_tree_add_7_25_groupi_n_3988 ,csa_tree_add_7_25_groupi_n_4483);
  nor csa_tree_add_7_25_groupi_g16563(csa_tree_add_7_25_groupi_n_4530 ,csa_tree_add_7_25_groupi_n_4018 ,csa_tree_add_7_25_groupi_n_4486);
  nor csa_tree_add_7_25_groupi_g16564(csa_tree_add_7_25_groupi_n_4529 ,csa_tree_add_7_25_groupi_n_3811 ,csa_tree_add_7_25_groupi_n_4457);
  nor csa_tree_add_7_25_groupi_g16565(csa_tree_add_7_25_groupi_n_4528 ,csa_tree_add_7_25_groupi_n_4057 ,csa_tree_add_7_25_groupi_n_4459);
  nor csa_tree_add_7_25_groupi_g16566(csa_tree_add_7_25_groupi_n_4527 ,csa_tree_add_7_25_groupi_n_3995 ,csa_tree_add_7_25_groupi_n_4487);
  and csa_tree_add_7_25_groupi_g16567(csa_tree_add_7_25_groupi_n_4554 ,csa_tree_add_7_25_groupi_n_3831 ,csa_tree_add_7_25_groupi_n_4480);
  nor csa_tree_add_7_25_groupi_g16568(csa_tree_add_7_25_groupi_n_4516 ,csa_tree_add_7_25_groupi_n_330 ,csa_tree_add_7_25_groupi_n_2021);
  nor csa_tree_add_7_25_groupi_g16569(csa_tree_add_7_25_groupi_n_4515 ,csa_tree_add_7_25_groupi_n_257 ,csa_tree_add_7_25_groupi_n_2069);
  nor csa_tree_add_7_25_groupi_g16570(csa_tree_add_7_25_groupi_n_4514 ,csa_tree_add_7_25_groupi_n_258 ,csa_tree_add_7_25_groupi_n_2088);
  nor csa_tree_add_7_25_groupi_g16571(csa_tree_add_7_25_groupi_n_4513 ,csa_tree_add_7_25_groupi_n_330 ,csa_tree_add_7_25_groupi_n_2082);
  nor csa_tree_add_7_25_groupi_g16572(csa_tree_add_7_25_groupi_n_4512 ,csa_tree_add_7_25_groupi_n_2076 ,csa_tree_add_7_25_groupi_n_1842);
  nor csa_tree_add_7_25_groupi_g16573(csa_tree_add_7_25_groupi_n_4511 ,csa_tree_add_7_25_groupi_n_329 ,csa_tree_add_7_25_groupi_n_2079);
  nor csa_tree_add_7_25_groupi_g16574(csa_tree_add_7_25_groupi_n_4510 ,csa_tree_add_7_25_groupi_n_2046 ,csa_tree_add_7_25_groupi_n_1843);
  xnor csa_tree_add_7_25_groupi_g16575(csa_tree_add_7_25_groupi_n_4509 ,csa_tree_add_7_25_groupi_n_4276 ,csa_tree_add_7_25_groupi_n_4401);
  xnor csa_tree_add_7_25_groupi_g16576(csa_tree_add_7_25_groupi_n_4508 ,csa_tree_add_7_25_groupi_n_4398 ,csa_tree_add_7_25_groupi_n_4409);
  xnor csa_tree_add_7_25_groupi_g16577(csa_tree_add_7_25_groupi_n_4507 ,csa_tree_add_7_25_groupi_n_4399 ,csa_tree_add_7_25_groupi_n_4408);
  xnor csa_tree_add_7_25_groupi_g16578(csa_tree_add_7_25_groupi_n_4506 ,csa_tree_add_7_25_groupi_n_4400 ,csa_tree_add_7_25_groupi_n_4407);
  xnor csa_tree_add_7_25_groupi_g16579(csa_tree_add_7_25_groupi_n_4505 ,csa_tree_add_7_25_groupi_n_1090 ,csa_tree_add_7_25_groupi_n_4369);
  xnor csa_tree_add_7_25_groupi_g16580(csa_tree_add_7_25_groupi_n_4504 ,csa_tree_add_7_25_groupi_n_4370 ,csa_tree_add_7_25_groupi_n_4392);
  xnor csa_tree_add_7_25_groupi_g16581(csa_tree_add_7_25_groupi_n_4503 ,csa_tree_add_7_25_groupi_n_4395 ,csa_tree_add_7_25_groupi_n_4405);
  xnor csa_tree_add_7_25_groupi_g16582(csa_tree_add_7_25_groupi_n_4502 ,csa_tree_add_7_25_groupi_n_4397 ,csa_tree_add_7_25_groupi_n_4396);
  xnor csa_tree_add_7_25_groupi_g16583(csa_tree_add_7_25_groupi_n_4501 ,csa_tree_add_7_25_groupi_n_4394 ,csa_tree_add_7_25_groupi_n_4402);
  xnor csa_tree_add_7_25_groupi_g16584(csa_tree_add_7_25_groupi_n_4500 ,csa_tree_add_7_25_groupi_n_4393 ,csa_tree_add_7_25_groupi_n_4403);
  xnor csa_tree_add_7_25_groupi_g16585(csa_tree_add_7_25_groupi_n_4499 ,csa_tree_add_7_25_groupi_n_4410 ,csa_tree_add_7_25_groupi_n_4404);
  xnor csa_tree_add_7_25_groupi_g16586(csa_tree_add_7_25_groupi_n_4526 ,csa_tree_add_7_25_groupi_n_4418 ,in3[5]);
  xnor csa_tree_add_7_25_groupi_g16587(csa_tree_add_7_25_groupi_n_4525 ,csa_tree_add_7_25_groupi_n_4415 ,in3[8]);
  xnor csa_tree_add_7_25_groupi_g16588(csa_tree_add_7_25_groupi_n_4524 ,csa_tree_add_7_25_groupi_n_4420 ,in3[11]);
  xnor csa_tree_add_7_25_groupi_g16589(csa_tree_add_7_25_groupi_n_4523 ,csa_tree_add_7_25_groupi_n_4419 ,in3[2]);
  xnor csa_tree_add_7_25_groupi_g16590(csa_tree_add_7_25_groupi_n_4522 ,csa_tree_add_7_25_groupi_n_4413 ,in3[14]);
  xnor csa_tree_add_7_25_groupi_g16591(csa_tree_add_7_25_groupi_n_4521 ,csa_tree_add_7_25_groupi_n_4421 ,in3[17]);
  xnor csa_tree_add_7_25_groupi_g16592(csa_tree_add_7_25_groupi_n_4520 ,csa_tree_add_7_25_groupi_n_4417 ,in3[20]);
  xnor csa_tree_add_7_25_groupi_g16593(csa_tree_add_7_25_groupi_n_4519 ,csa_tree_add_7_25_groupi_n_4422 ,in3[23]);
  xnor csa_tree_add_7_25_groupi_g16594(csa_tree_add_7_25_groupi_n_4518 ,csa_tree_add_7_25_groupi_n_4414 ,in3[26]);
  xnor csa_tree_add_7_25_groupi_g16595(csa_tree_add_7_25_groupi_n_4517 ,csa_tree_add_7_25_groupi_n_4416 ,in3[29]);
  or csa_tree_add_7_25_groupi_g16596(csa_tree_add_7_25_groupi_n_4488 ,csa_tree_add_7_25_groupi_n_4400 ,csa_tree_add_7_25_groupi_n_4407);
  or csa_tree_add_7_25_groupi_g16597(csa_tree_add_7_25_groupi_n_4487 ,csa_tree_add_7_25_groupi_n_3135 ,csa_tree_add_7_25_groupi_n_4436);
  or csa_tree_add_7_25_groupi_g16598(csa_tree_add_7_25_groupi_n_4486 ,csa_tree_add_7_25_groupi_n_3152 ,csa_tree_add_7_25_groupi_n_4434);
  or csa_tree_add_7_25_groupi_g16599(csa_tree_add_7_25_groupi_n_4485 ,csa_tree_add_7_25_groupi_n_3607 ,csa_tree_add_7_25_groupi_n_4427);
  or csa_tree_add_7_25_groupi_g16600(csa_tree_add_7_25_groupi_n_4484 ,csa_tree_add_7_25_groupi_n_4398 ,csa_tree_add_7_25_groupi_n_4409);
  or csa_tree_add_7_25_groupi_g16601(csa_tree_add_7_25_groupi_n_4483 ,csa_tree_add_7_25_groupi_n_3177 ,csa_tree_add_7_25_groupi_n_4433);
  or csa_tree_add_7_25_groupi_g16602(csa_tree_add_7_25_groupi_n_4482 ,csa_tree_add_7_25_groupi_n_3215 ,csa_tree_add_7_25_groupi_n_2);
  and csa_tree_add_7_25_groupi_g16603(csa_tree_add_7_25_groupi_n_4481 ,csa_tree_add_7_25_groupi_n_4400 ,csa_tree_add_7_25_groupi_n_4407);
  nor csa_tree_add_7_25_groupi_g16604(csa_tree_add_7_25_groupi_n_4480 ,csa_tree_add_7_25_groupi_n_3371 ,csa_tree_add_7_25_groupi_n_4425);
  and csa_tree_add_7_25_groupi_g16605(csa_tree_add_7_25_groupi_n_4479 ,csa_tree_add_7_25_groupi_n_1972 ,csa_tree_add_7_25_groupi_n_1094);
  nor csa_tree_add_7_25_groupi_g16606(csa_tree_add_7_25_groupi_n_4478 ,csa_tree_add_7_25_groupi_n_4314 ,csa_tree_add_7_25_groupi_n_4430);
  and csa_tree_add_7_25_groupi_g16607(csa_tree_add_7_25_groupi_n_4477 ,csa_tree_add_7_25_groupi_n_4399 ,csa_tree_add_7_25_groupi_n_4408);
  or csa_tree_add_7_25_groupi_g16608(csa_tree_add_7_25_groupi_n_4476 ,csa_tree_add_7_25_groupi_n_4369 ,csa_tree_add_7_25_groupi_n_1090);
  and csa_tree_add_7_25_groupi_g16609(csa_tree_add_7_25_groupi_n_4475 ,csa_tree_add_7_25_groupi_n_4276 ,csa_tree_add_7_25_groupi_n_4401);
  or csa_tree_add_7_25_groupi_g16610(csa_tree_add_7_25_groupi_n_4474 ,csa_tree_add_7_25_groupi_n_4276 ,csa_tree_add_7_25_groupi_n_4401);
  and csa_tree_add_7_25_groupi_g16611(csa_tree_add_7_25_groupi_n_4473 ,csa_tree_add_7_25_groupi_n_4398 ,csa_tree_add_7_25_groupi_n_4409);
  or csa_tree_add_7_25_groupi_g16612(csa_tree_add_7_25_groupi_n_4472 ,csa_tree_add_7_25_groupi_n_4399 ,csa_tree_add_7_25_groupi_n_4408);
  or csa_tree_add_7_25_groupi_g16613(csa_tree_add_7_25_groupi_n_4498 ,csa_tree_add_7_25_groupi_n_4274 ,csa_tree_add_7_25_groupi_n_4423);
  or csa_tree_add_7_25_groupi_g16614(csa_tree_add_7_25_groupi_n_4497 ,csa_tree_add_7_25_groupi_n_4302 ,csa_tree_add_7_25_groupi_n_4424);
  or csa_tree_add_7_25_groupi_g16615(csa_tree_add_7_25_groupi_n_4496 ,csa_tree_add_7_25_groupi_n_4300 ,csa_tree_add_7_25_groupi_n_4440);
  or csa_tree_add_7_25_groupi_g16616(csa_tree_add_7_25_groupi_n_4495 ,csa_tree_add_7_25_groupi_n_4316 ,csa_tree_add_7_25_groupi_n_4431);
  or csa_tree_add_7_25_groupi_g16617(csa_tree_add_7_25_groupi_n_4494 ,csa_tree_add_7_25_groupi_n_4272 ,csa_tree_add_7_25_groupi_n_4432);
  or csa_tree_add_7_25_groupi_g16618(csa_tree_add_7_25_groupi_n_4493 ,csa_tree_add_7_25_groupi_n_4315 ,csa_tree_add_7_25_groupi_n_4438);
  or csa_tree_add_7_25_groupi_g16619(csa_tree_add_7_25_groupi_n_4492 ,csa_tree_add_7_25_groupi_n_4304 ,csa_tree_add_7_25_groupi_n_4441);
  and csa_tree_add_7_25_groupi_g16620(csa_tree_add_7_25_groupi_n_4491 ,csa_tree_add_7_25_groupi_n_2460 ,csa_tree_add_7_25_groupi_n_4435);
  or csa_tree_add_7_25_groupi_g16621(csa_tree_add_7_25_groupi_n_4490 ,csa_tree_add_7_25_groupi_n_4275 ,csa_tree_add_7_25_groupi_n_4426);
  or csa_tree_add_7_25_groupi_g16622(csa_tree_add_7_25_groupi_n_4489 ,csa_tree_add_7_25_groupi_n_4313 ,csa_tree_add_7_25_groupi_n_4439);
  not csa_tree_add_7_25_groupi_g16623(csa_tree_add_7_25_groupi_n_4471 ,csa_tree_add_7_25_groupi_n_4470);
  or csa_tree_add_7_25_groupi_g16624(csa_tree_add_7_25_groupi_n_4459 ,csa_tree_add_7_25_groupi_n_3122 ,csa_tree_add_7_25_groupi_n_4390);
  or csa_tree_add_7_25_groupi_g16625(csa_tree_add_7_25_groupi_n_4458 ,csa_tree_add_7_25_groupi_n_3104 ,csa_tree_add_7_25_groupi_n_4437);
  or csa_tree_add_7_25_groupi_g16626(csa_tree_add_7_25_groupi_n_4457 ,csa_tree_add_7_25_groupi_n_3584 ,csa_tree_add_7_25_groupi_n_4429);
  and csa_tree_add_7_25_groupi_g16627(csa_tree_add_7_25_groupi_n_4456 ,csa_tree_add_7_25_groupi_n_4397 ,csa_tree_add_7_25_groupi_n_4396);
  or csa_tree_add_7_25_groupi_g16628(csa_tree_add_7_25_groupi_n_4455 ,csa_tree_add_7_25_groupi_n_4397 ,csa_tree_add_7_25_groupi_n_4396);
  and csa_tree_add_7_25_groupi_g16629(csa_tree_add_7_25_groupi_n_4454 ,csa_tree_add_7_25_groupi_n_4395 ,csa_tree_add_7_25_groupi_n_4405);
  or csa_tree_add_7_25_groupi_g16630(csa_tree_add_7_25_groupi_n_4453 ,csa_tree_add_7_25_groupi_n_4395 ,csa_tree_add_7_25_groupi_n_4405);
  or csa_tree_add_7_25_groupi_g16631(csa_tree_add_7_25_groupi_n_4452 ,csa_tree_add_7_25_groupi_n_4410 ,csa_tree_add_7_25_groupi_n_4404);
  and csa_tree_add_7_25_groupi_g16632(csa_tree_add_7_25_groupi_n_4451 ,csa_tree_add_7_25_groupi_n_4410 ,csa_tree_add_7_25_groupi_n_4404);
  or csa_tree_add_7_25_groupi_g16633(csa_tree_add_7_25_groupi_n_4450 ,csa_tree_add_7_25_groupi_n_4393 ,csa_tree_add_7_25_groupi_n_4403);
  or csa_tree_add_7_25_groupi_g16634(csa_tree_add_7_25_groupi_n_4449 ,csa_tree_add_7_25_groupi_n_4394 ,csa_tree_add_7_25_groupi_n_4402);
  and csa_tree_add_7_25_groupi_g16635(csa_tree_add_7_25_groupi_n_4448 ,csa_tree_add_7_25_groupi_n_4394 ,csa_tree_add_7_25_groupi_n_4402);
  and csa_tree_add_7_25_groupi_g16636(csa_tree_add_7_25_groupi_n_4447 ,csa_tree_add_7_25_groupi_n_4393 ,csa_tree_add_7_25_groupi_n_4403);
  or csa_tree_add_7_25_groupi_g16637(csa_tree_add_7_25_groupi_n_4446 ,csa_tree_add_7_25_groupi_n_2980 ,csa_tree_add_7_25_groupi_n_4428);
  or csa_tree_add_7_25_groupi_g16638(csa_tree_add_7_25_groupi_n_4445 ,csa_tree_add_7_25_groupi_n_4392 ,csa_tree_add_7_25_groupi_n_4370);
  and csa_tree_add_7_25_groupi_g16639(csa_tree_add_7_25_groupi_n_4444 ,csa_tree_add_7_25_groupi_n_4392 ,csa_tree_add_7_25_groupi_n_4370);
  or csa_tree_add_7_25_groupi_g16640(csa_tree_add_7_25_groupi_n_4443 ,csa_tree_add_7_25_groupi_n_3103 ,csa_tree_add_7_25_groupi_n_4391);
  xnor csa_tree_add_7_25_groupi_g16641(csa_tree_add_7_25_groupi_n_4470 ,csa_tree_add_7_25_groupi_n_4160 ,csa_tree_add_7_25_groupi_n_4332);
  xnor csa_tree_add_7_25_groupi_g16642(csa_tree_add_7_25_groupi_n_4469 ,csa_tree_add_7_25_groupi_n_4375 ,csa_tree_add_7_25_groupi_n_4330);
  xnor csa_tree_add_7_25_groupi_g16643(csa_tree_add_7_25_groupi_n_4468 ,csa_tree_add_7_25_groupi_n_4379 ,csa_tree_add_7_25_groupi_n_4331);
  xnor csa_tree_add_7_25_groupi_g16644(csa_tree_add_7_25_groupi_n_4467 ,csa_tree_add_7_25_groupi_n_4378 ,csa_tree_add_7_25_groupi_n_4333);
  xnor csa_tree_add_7_25_groupi_g16645(csa_tree_add_7_25_groupi_n_4466 ,csa_tree_add_7_25_groupi_n_4372 ,csa_tree_add_7_25_groupi_n_4326);
  xnor csa_tree_add_7_25_groupi_g16646(csa_tree_add_7_25_groupi_n_4465 ,csa_tree_add_7_25_groupi_n_4374 ,csa_tree_add_7_25_groupi_n_4325);
  xnor csa_tree_add_7_25_groupi_g16647(csa_tree_add_7_25_groupi_n_4464 ,csa_tree_add_7_25_groupi_n_4380 ,csa_tree_add_7_25_groupi_n_4324);
  xnor csa_tree_add_7_25_groupi_g16648(csa_tree_add_7_25_groupi_n_4463 ,csa_tree_add_7_25_groupi_n_4377 ,csa_tree_add_7_25_groupi_n_4327);
  xnor csa_tree_add_7_25_groupi_g16649(csa_tree_add_7_25_groupi_n_4462 ,csa_tree_add_7_25_groupi_n_4373 ,csa_tree_add_7_25_groupi_n_4328);
  xnor csa_tree_add_7_25_groupi_g16650(csa_tree_add_7_25_groupi_n_4461 ,csa_tree_add_7_25_groupi_n_4376 ,csa_tree_add_7_25_groupi_n_4329);
  xnor csa_tree_add_7_25_groupi_g16651(csa_tree_add_7_25_groupi_n_4460 ,csa_tree_add_7_25_groupi_n_4371 ,csa_tree_add_7_25_groupi_n_2580);
  and csa_tree_add_7_25_groupi_g16653(csa_tree_add_7_25_groupi_n_4441 ,csa_tree_add_7_25_groupi_n_4308 ,csa_tree_add_7_25_groupi_n_4373);
  and csa_tree_add_7_25_groupi_g16654(csa_tree_add_7_25_groupi_n_4440 ,csa_tree_add_7_25_groupi_n_4319 ,csa_tree_add_7_25_groupi_n_4375);
  and csa_tree_add_7_25_groupi_g16655(csa_tree_add_7_25_groupi_n_4439 ,csa_tree_add_7_25_groupi_n_4312 ,csa_tree_add_7_25_groupi_n_4378);
  and csa_tree_add_7_25_groupi_g16656(csa_tree_add_7_25_groupi_n_4438 ,csa_tree_add_7_25_groupi_n_4303 ,csa_tree_add_7_25_groupi_n_4380);
  nor csa_tree_add_7_25_groupi_g16657(csa_tree_add_7_25_groupi_n_4437 ,csa_tree_add_7_25_groupi_n_295 ,csa_tree_add_7_25_groupi_n_2114);
  nor csa_tree_add_7_25_groupi_g16658(csa_tree_add_7_25_groupi_n_4436 ,csa_tree_add_7_25_groupi_n_2129 ,csa_tree_add_7_25_groupi_n_1839);
  or csa_tree_add_7_25_groupi_g16659(csa_tree_add_7_25_groupi_n_4435 ,csa_tree_add_7_25_groupi_n_2491 ,csa_tree_add_7_25_groupi_n_4371);
  nor csa_tree_add_7_25_groupi_g16660(csa_tree_add_7_25_groupi_n_4434 ,csa_tree_add_7_25_groupi_n_2072 ,csa_tree_add_7_25_groupi_n_204);
  nor csa_tree_add_7_25_groupi_g16661(csa_tree_add_7_25_groupi_n_4433 ,csa_tree_add_7_25_groupi_n_2040 ,csa_tree_add_7_25_groupi_n_1839);
  and csa_tree_add_7_25_groupi_g16662(csa_tree_add_7_25_groupi_n_4432 ,csa_tree_add_7_25_groupi_n_4318 ,csa_tree_add_7_25_groupi_n_4376);
  and csa_tree_add_7_25_groupi_g16663(csa_tree_add_7_25_groupi_n_4431 ,csa_tree_add_7_25_groupi_n_4310 ,csa_tree_add_7_25_groupi_n_4379);
  nor csa_tree_add_7_25_groupi_g16664(csa_tree_add_7_25_groupi_n_4430 ,csa_tree_add_7_25_groupi_n_4260 ,csa_tree_add_7_25_groupi_n_4368);
  nor csa_tree_add_7_25_groupi_g16666(csa_tree_add_7_25_groupi_n_4429 ,csa_tree_add_7_25_groupi_n_555 ,csa_tree_add_7_25_groupi_n_268);
  nor csa_tree_add_7_25_groupi_g16667(csa_tree_add_7_25_groupi_n_4428 ,csa_tree_add_7_25_groupi_n_268 ,csa_tree_add_7_25_groupi_n_2171);
  nor csa_tree_add_7_25_groupi_g16668(csa_tree_add_7_25_groupi_n_4427 ,csa_tree_add_7_25_groupi_n_483 ,csa_tree_add_7_25_groupi_n_295);
  and csa_tree_add_7_25_groupi_g16669(csa_tree_add_7_25_groupi_n_4426 ,csa_tree_add_7_25_groupi_n_4298 ,csa_tree_add_7_25_groupi_n_4374);
  nor csa_tree_add_7_25_groupi_g16670(csa_tree_add_7_25_groupi_n_4425 ,csa_tree_add_7_25_groupi_n_552 ,csa_tree_add_7_25_groupi_n_204);
  and csa_tree_add_7_25_groupi_g16671(csa_tree_add_7_25_groupi_n_4424 ,csa_tree_add_7_25_groupi_n_4307 ,csa_tree_add_7_25_groupi_n_4377);
  and csa_tree_add_7_25_groupi_g16672(csa_tree_add_7_25_groupi_n_4423 ,csa_tree_add_7_25_groupi_n_4306 ,csa_tree_add_7_25_groupi_n_4372);
  nor csa_tree_add_7_25_groupi_g16673(csa_tree_add_7_25_groupi_n_4422 ,csa_tree_add_7_25_groupi_n_3867 ,csa_tree_add_7_25_groupi_n_4350);
  nor csa_tree_add_7_25_groupi_g16674(csa_tree_add_7_25_groupi_n_4421 ,csa_tree_add_7_25_groupi_n_4082 ,csa_tree_add_7_25_groupi_n_4342);
  nor csa_tree_add_7_25_groupi_g16675(csa_tree_add_7_25_groupi_n_4420 ,csa_tree_add_7_25_groupi_n_4052 ,csa_tree_add_7_25_groupi_n_4339);
  nor csa_tree_add_7_25_groupi_g16676(csa_tree_add_7_25_groupi_n_4419 ,csa_tree_add_7_25_groupi_n_3464 ,csa_tree_add_7_25_groupi_n_4334);
  nor csa_tree_add_7_25_groupi_g16677(csa_tree_add_7_25_groupi_n_4418 ,csa_tree_add_7_25_groupi_n_4066 ,csa_tree_add_7_25_groupi_n_4341);
  nor csa_tree_add_7_25_groupi_g16678(csa_tree_add_7_25_groupi_n_4417 ,csa_tree_add_7_25_groupi_n_3987 ,csa_tree_add_7_25_groupi_n_4344);
  nor csa_tree_add_7_25_groupi_g16679(csa_tree_add_7_25_groupi_n_4416 ,csa_tree_add_7_25_groupi_n_3845 ,csa_tree_add_7_25_groupi_n_4343);
  nor csa_tree_add_7_25_groupi_g16680(csa_tree_add_7_25_groupi_n_4415 ,csa_tree_add_7_25_groupi_n_4026 ,csa_tree_add_7_25_groupi_n_4338);
  nor csa_tree_add_7_25_groupi_g16681(csa_tree_add_7_25_groupi_n_4414 ,csa_tree_add_7_25_groupi_n_3910 ,csa_tree_add_7_25_groupi_n_4337);
  nor csa_tree_add_7_25_groupi_g16682(csa_tree_add_7_25_groupi_n_4413 ,csa_tree_add_7_25_groupi_n_4059 ,csa_tree_add_7_25_groupi_n_4340);
  and csa_tree_add_7_25_groupi_g16683(csa_tree_add_7_25_groupi_n_4442 ,csa_tree_add_7_25_groupi_n_3929 ,csa_tree_add_7_25_groupi_n_4335);
  not csa_tree_add_7_25_groupi_g16684(csa_tree_add_7_25_groupi_n_4412 ,csa_tree_add_7_25_groupi_n_4411);
  nor csa_tree_add_7_25_groupi_g16685(csa_tree_add_7_25_groupi_n_4391 ,csa_tree_add_7_25_groupi_n_294 ,csa_tree_add_7_25_groupi_n_2093);
  nor csa_tree_add_7_25_groupi_g16686(csa_tree_add_7_25_groupi_n_4390 ,csa_tree_add_7_25_groupi_n_2147 ,csa_tree_add_7_25_groupi_n_1840);
  xnor csa_tree_add_7_25_groupi_g16687(csa_tree_add_7_25_groupi_n_4411 ,csa_tree_add_7_25_groupi_n_4288 ,in3[2]);
  xnor csa_tree_add_7_25_groupi_g16688(csa_tree_add_7_25_groupi_n_4389 ,csa_tree_add_7_25_groupi_n_4199 ,csa_tree_add_7_25_groupi_n_4278);
  xnor csa_tree_add_7_25_groupi_g16689(csa_tree_add_7_25_groupi_n_4388 ,csa_tree_add_7_25_groupi_n_4200 ,csa_tree_add_7_25_groupi_n_4279);
  xnor csa_tree_add_7_25_groupi_g16690(csa_tree_add_7_25_groupi_n_4387 ,csa_tree_add_7_25_groupi_n_4201 ,csa_tree_add_7_25_groupi_n_4280);
  xnor csa_tree_add_7_25_groupi_g16691(csa_tree_add_7_25_groupi_n_4386 ,csa_tree_add_7_25_groupi_n_4202 ,csa_tree_add_7_25_groupi_n_4281);
  xnor csa_tree_add_7_25_groupi_g16692(csa_tree_add_7_25_groupi_n_4385 ,csa_tree_add_7_25_groupi_n_4203 ,csa_tree_add_7_25_groupi_n_4282);
  xnor csa_tree_add_7_25_groupi_g16693(csa_tree_add_7_25_groupi_n_4384 ,csa_tree_add_7_25_groupi_n_4206 ,csa_tree_add_7_25_groupi_n_4283);
  xnor csa_tree_add_7_25_groupi_g16694(csa_tree_add_7_25_groupi_n_4383 ,csa_tree_add_7_25_groupi_n_4207 ,csa_tree_add_7_25_groupi_n_4284);
  xnor csa_tree_add_7_25_groupi_g16695(csa_tree_add_7_25_groupi_n_4382 ,csa_tree_add_7_25_groupi_n_4205 ,csa_tree_add_7_25_groupi_n_4285);
  xnor csa_tree_add_7_25_groupi_g16696(csa_tree_add_7_25_groupi_n_4381 ,csa_tree_add_7_25_groupi_n_4111 ,csa_tree_add_7_25_groupi_n_4277);
  xnor csa_tree_add_7_25_groupi_g16697(csa_tree_add_7_25_groupi_n_4410 ,csa_tree_add_7_25_groupi_n_4292 ,in3[11]);
  xnor csa_tree_add_7_25_groupi_g16698(csa_tree_add_7_25_groupi_n_4409 ,csa_tree_add_7_25_groupi_n_4247 ,csa_tree_add_7_25_groupi_n_4255);
  xnor csa_tree_add_7_25_groupi_g16699(csa_tree_add_7_25_groupi_n_4408 ,csa_tree_add_7_25_groupi_n_4240 ,csa_tree_add_7_25_groupi_n_4256);
  xnor csa_tree_add_7_25_groupi_g16700(csa_tree_add_7_25_groupi_n_4407 ,csa_tree_add_7_25_groupi_n_4243 ,csa_tree_add_7_25_groupi_n_4258);
  xnor csa_tree_add_7_25_groupi_g16701(csa_tree_add_7_25_groupi_n_4406 ,csa_tree_add_7_25_groupi_n_4185 ,csa_tree_add_7_25_groupi_n_4321);
  xnor csa_tree_add_7_25_groupi_g16702(csa_tree_add_7_25_groupi_n_4405 ,csa_tree_add_7_25_groupi_n_4244 ,csa_tree_add_7_25_groupi_n_4253);
  xnor csa_tree_add_7_25_groupi_g16703(csa_tree_add_7_25_groupi_n_4404 ,csa_tree_add_7_25_groupi_n_4216 ,csa_tree_add_7_25_groupi_n_4250);
  xnor csa_tree_add_7_25_groupi_g16704(csa_tree_add_7_25_groupi_n_4403 ,csa_tree_add_7_25_groupi_n_4246 ,csa_tree_add_7_25_groupi_n_4252);
  xnor csa_tree_add_7_25_groupi_g16705(csa_tree_add_7_25_groupi_n_4402 ,csa_tree_add_7_25_groupi_n_4248 ,csa_tree_add_7_25_groupi_n_4251);
  xnor csa_tree_add_7_25_groupi_g16706(csa_tree_add_7_25_groupi_n_4401 ,csa_tree_add_7_25_groupi_n_4293 ,in3[29]);
  xnor csa_tree_add_7_25_groupi_g16707(csa_tree_add_7_25_groupi_n_4400 ,csa_tree_add_7_25_groupi_n_4289 ,in3[26]);
  xnor csa_tree_add_7_25_groupi_g16708(csa_tree_add_7_25_groupi_n_4399 ,csa_tree_add_7_25_groupi_n_4291 ,in3[23]);
  xnor csa_tree_add_7_25_groupi_g16709(csa_tree_add_7_25_groupi_n_4398 ,csa_tree_add_7_25_groupi_n_4259 ,in3[20]);
  xnor csa_tree_add_7_25_groupi_g16710(csa_tree_add_7_25_groupi_n_4397 ,csa_tree_add_7_25_groupi_n_4290 ,in3[17]);
  xnor csa_tree_add_7_25_groupi_g16711(csa_tree_add_7_25_groupi_n_4396 ,csa_tree_add_7_25_groupi_n_4241 ,csa_tree_add_7_25_groupi_n_4254);
  xnor csa_tree_add_7_25_groupi_g16712(csa_tree_add_7_25_groupi_n_4395 ,csa_tree_add_7_25_groupi_n_4287 ,in3[14]);
  xnor csa_tree_add_7_25_groupi_g16713(csa_tree_add_7_25_groupi_n_4394 ,csa_tree_add_7_25_groupi_n_4257 ,in3[5]);
  xnor csa_tree_add_7_25_groupi_g16714(csa_tree_add_7_25_groupi_n_4393 ,csa_tree_add_7_25_groupi_n_4294 ,in3[8]);
  or csa_tree_add_7_25_groupi_g16715(csa_tree_add_7_25_groupi_n_4392 ,csa_tree_add_7_25_groupi_n_4356 ,csa_tree_add_7_25_groupi_n_2341);
  nor csa_tree_add_7_25_groupi_g16717(csa_tree_add_7_25_groupi_n_4368 ,csa_tree_add_7_25_groupi_n_4226 ,csa_tree_add_7_25_groupi_n_4295);
  or csa_tree_add_7_25_groupi_g16718(csa_tree_add_7_25_groupi_n_4367 ,csa_tree_add_7_25_groupi_n_4202 ,csa_tree_add_7_25_groupi_n_4281);
  and csa_tree_add_7_25_groupi_g16719(csa_tree_add_7_25_groupi_n_4366 ,csa_tree_add_7_25_groupi_n_4199 ,csa_tree_add_7_25_groupi_n_4278);
  and csa_tree_add_7_25_groupi_g16720(csa_tree_add_7_25_groupi_n_4365 ,csa_tree_add_7_25_groupi_n_4286 ,csa_tree_add_7_25_groupi_n_4218);
  and csa_tree_add_7_25_groupi_g16721(csa_tree_add_7_25_groupi_n_4364 ,csa_tree_add_7_25_groupi_n_4201 ,csa_tree_add_7_25_groupi_n_4280);
  and csa_tree_add_7_25_groupi_g16722(csa_tree_add_7_25_groupi_n_4363 ,csa_tree_add_7_25_groupi_n_4203 ,csa_tree_add_7_25_groupi_n_4282);
  or csa_tree_add_7_25_groupi_g16723(csa_tree_add_7_25_groupi_n_4362 ,csa_tree_add_7_25_groupi_n_4199 ,csa_tree_add_7_25_groupi_n_4278);
  or csa_tree_add_7_25_groupi_g16724(csa_tree_add_7_25_groupi_n_4361 ,csa_tree_add_7_25_groupi_n_4201 ,csa_tree_add_7_25_groupi_n_4280);
  or csa_tree_add_7_25_groupi_g16725(csa_tree_add_7_25_groupi_n_4360 ,csa_tree_add_7_25_groupi_n_4200 ,csa_tree_add_7_25_groupi_n_4279);
  or csa_tree_add_7_25_groupi_g16726(csa_tree_add_7_25_groupi_n_4359 ,csa_tree_add_7_25_groupi_n_4203 ,csa_tree_add_7_25_groupi_n_4282);
  and csa_tree_add_7_25_groupi_g16727(csa_tree_add_7_25_groupi_n_4358 ,csa_tree_add_7_25_groupi_n_4200 ,csa_tree_add_7_25_groupi_n_4279);
  and csa_tree_add_7_25_groupi_g16728(csa_tree_add_7_25_groupi_n_4357 ,csa_tree_add_7_25_groupi_n_4202 ,csa_tree_add_7_25_groupi_n_4281);
  nor csa_tree_add_7_25_groupi_g16729(csa_tree_add_7_25_groupi_n_4356 ,in3[2] ,csa_tree_add_7_25_groupi_n_4322);
  or csa_tree_add_7_25_groupi_g16730(csa_tree_add_7_25_groupi_n_4355 ,csa_tree_add_7_25_groupi_n_4111 ,csa_tree_add_7_25_groupi_n_4277);
  nor csa_tree_add_7_25_groupi_g16731(csa_tree_add_7_25_groupi_n_4354 ,csa_tree_add_7_25_groupi_n_4286 ,csa_tree_add_7_25_groupi_n_4218);
  and csa_tree_add_7_25_groupi_g16732(csa_tree_add_7_25_groupi_n_4353 ,csa_tree_add_7_25_groupi_n_4111 ,csa_tree_add_7_25_groupi_n_4277);
  or csa_tree_add_7_25_groupi_g16733(csa_tree_add_7_25_groupi_n_4380 ,csa_tree_add_7_25_groupi_n_4220 ,csa_tree_add_7_25_groupi_n_4320);
  or csa_tree_add_7_25_groupi_g16734(csa_tree_add_7_25_groupi_n_4379 ,csa_tree_add_7_25_groupi_n_4239 ,csa_tree_add_7_25_groupi_n_4296);
  or csa_tree_add_7_25_groupi_g16735(csa_tree_add_7_25_groupi_n_4378 ,csa_tree_add_7_25_groupi_n_4231 ,csa_tree_add_7_25_groupi_n_4311);
  or csa_tree_add_7_25_groupi_g16736(csa_tree_add_7_25_groupi_n_4377 ,csa_tree_add_7_25_groupi_n_4224 ,csa_tree_add_7_25_groupi_n_4309);
  or csa_tree_add_7_25_groupi_g16737(csa_tree_add_7_25_groupi_n_4376 ,csa_tree_add_7_25_groupi_n_4234 ,csa_tree_add_7_25_groupi_n_4297);
  or csa_tree_add_7_25_groupi_g16738(csa_tree_add_7_25_groupi_n_4375 ,csa_tree_add_7_25_groupi_n_4236 ,csa_tree_add_7_25_groupi_n_4299);
  or csa_tree_add_7_25_groupi_g16739(csa_tree_add_7_25_groupi_n_4374 ,csa_tree_add_7_25_groupi_n_4221 ,csa_tree_add_7_25_groupi_n_4301);
  or csa_tree_add_7_25_groupi_g16740(csa_tree_add_7_25_groupi_n_4373 ,csa_tree_add_7_25_groupi_n_4232 ,csa_tree_add_7_25_groupi_n_4317);
  or csa_tree_add_7_25_groupi_g16741(csa_tree_add_7_25_groupi_n_4372 ,csa_tree_add_7_25_groupi_n_4230 ,csa_tree_add_7_25_groupi_n_4273);
  and csa_tree_add_7_25_groupi_g16742(csa_tree_add_7_25_groupi_n_4371 ,csa_tree_add_7_25_groupi_n_2495 ,csa_tree_add_7_25_groupi_n_4305);
  and csa_tree_add_7_25_groupi_g16743(csa_tree_add_7_25_groupi_n_4370 ,csa_tree_add_7_25_groupi_n_4186 ,csa_tree_add_7_25_groupi_n_4321);
  or csa_tree_add_7_25_groupi_g16744(csa_tree_add_7_25_groupi_n_4369 ,csa_tree_add_7_25_groupi_n_1092 ,csa_tree_add_7_25_groupi_n_4323);
  or csa_tree_add_7_25_groupi_g16745(csa_tree_add_7_25_groupi_n_4350 ,csa_tree_add_7_25_groupi_n_3630 ,csa_tree_add_7_25_groupi_n_4267);
  or csa_tree_add_7_25_groupi_g16746(csa_tree_add_7_25_groupi_n_4349 ,csa_tree_add_7_25_groupi_n_4207 ,csa_tree_add_7_25_groupi_n_4284);
  or csa_tree_add_7_25_groupi_g16747(csa_tree_add_7_25_groupi_n_4348 ,csa_tree_add_7_25_groupi_n_4205 ,csa_tree_add_7_25_groupi_n_4285);
  or csa_tree_add_7_25_groupi_g16748(csa_tree_add_7_25_groupi_n_4347 ,csa_tree_add_7_25_groupi_n_4206 ,csa_tree_add_7_25_groupi_n_4283);
  and csa_tree_add_7_25_groupi_g16749(csa_tree_add_7_25_groupi_n_4346 ,csa_tree_add_7_25_groupi_n_4206 ,csa_tree_add_7_25_groupi_n_4283);
  and csa_tree_add_7_25_groupi_g16750(csa_tree_add_7_25_groupi_n_4345 ,csa_tree_add_7_25_groupi_n_4207 ,csa_tree_add_7_25_groupi_n_4284);
  or csa_tree_add_7_25_groupi_g16751(csa_tree_add_7_25_groupi_n_4344 ,csa_tree_add_7_25_groupi_n_3179 ,csa_tree_add_7_25_groupi_n_4266);
  or csa_tree_add_7_25_groupi_g16752(csa_tree_add_7_25_groupi_n_4343 ,csa_tree_add_7_25_groupi_n_3643 ,csa_tree_add_7_25_groupi_n_4270);
  or csa_tree_add_7_25_groupi_g16753(csa_tree_add_7_25_groupi_n_4342 ,csa_tree_add_7_25_groupi_n_3156 ,csa_tree_add_7_25_groupi_n_4265);
  or csa_tree_add_7_25_groupi_g16754(csa_tree_add_7_25_groupi_n_4341 ,csa_tree_add_7_25_groupi_n_3139 ,csa_tree_add_7_25_groupi_n_4264);
  or csa_tree_add_7_25_groupi_g16755(csa_tree_add_7_25_groupi_n_4340 ,csa_tree_add_7_25_groupi_n_3108 ,csa_tree_add_7_25_groupi_n_4262);
  or csa_tree_add_7_25_groupi_g16756(csa_tree_add_7_25_groupi_n_4339 ,csa_tree_add_7_25_groupi_n_3124 ,csa_tree_add_7_25_groupi_n_4263);
  or csa_tree_add_7_25_groupi_g16757(csa_tree_add_7_25_groupi_n_4338 ,csa_tree_add_7_25_groupi_n_3101 ,csa_tree_add_7_25_groupi_n_4261);
  or csa_tree_add_7_25_groupi_g16758(csa_tree_add_7_25_groupi_n_4337 ,csa_tree_add_7_25_groupi_n_3560 ,csa_tree_add_7_25_groupi_n_4268);
  and csa_tree_add_7_25_groupi_g16759(csa_tree_add_7_25_groupi_n_4336 ,csa_tree_add_7_25_groupi_n_4205 ,csa_tree_add_7_25_groupi_n_4285);
  nor csa_tree_add_7_25_groupi_g16760(csa_tree_add_7_25_groupi_n_4335 ,csa_tree_add_7_25_groupi_n_3025 ,csa_tree_add_7_25_groupi_n_4271);
  or csa_tree_add_7_25_groupi_g16761(csa_tree_add_7_25_groupi_n_4334 ,csa_tree_add_7_25_groupi_n_2969 ,csa_tree_add_7_25_groupi_n_4269);
  xnor csa_tree_add_7_25_groupi_g16762(csa_tree_add_7_25_groupi_n_4333 ,csa_tree_add_7_25_groupi_n_4213 ,in2[17]);
  xnor csa_tree_add_7_25_groupi_g16763(csa_tree_add_7_25_groupi_n_4332 ,csa_tree_add_7_25_groupi_n_4249 ,in2[4]);
  xnor csa_tree_add_7_25_groupi_g16764(csa_tree_add_7_25_groupi_n_4331 ,csa_tree_add_7_25_groupi_n_4208 ,in2[5]);
  xnor csa_tree_add_7_25_groupi_g16765(csa_tree_add_7_25_groupi_n_4330 ,csa_tree_add_7_25_groupi_n_4210 ,in2[11]);
  xnor csa_tree_add_7_25_groupi_g16766(csa_tree_add_7_25_groupi_n_4329 ,csa_tree_add_7_25_groupi_n_4209 ,in2[8]);
  xnor csa_tree_add_7_25_groupi_g16767(csa_tree_add_7_25_groupi_n_4328 ,csa_tree_add_7_25_groupi_n_4211 ,in2[14]);
  xnor csa_tree_add_7_25_groupi_g16768(csa_tree_add_7_25_groupi_n_4327 ,csa_tree_add_7_25_groupi_n_4212 ,in2[29]);
  xnor csa_tree_add_7_25_groupi_g16769(csa_tree_add_7_25_groupi_n_4326 ,csa_tree_add_7_25_groupi_n_4214 ,in2[20]);
  xnor csa_tree_add_7_25_groupi_g16770(csa_tree_add_7_25_groupi_n_4325 ,csa_tree_add_7_25_groupi_n_4215 ,in2[23]);
  xnor csa_tree_add_7_25_groupi_g16771(csa_tree_add_7_25_groupi_n_4324 ,csa_tree_add_7_25_groupi_n_4204 ,in2[26]);
  xnor csa_tree_add_7_25_groupi_g16772(csa_tree_add_7_25_groupi_n_4352 ,csa_tree_add_7_25_groupi_n_4245 ,csa_tree_add_7_25_groupi_n_4138);
  xnor csa_tree_add_7_25_groupi_g16773(csa_tree_add_7_25_groupi_n_4351 ,csa_tree_add_7_25_groupi_n_4242 ,csa_tree_add_7_25_groupi_n_2584);
  not csa_tree_add_7_25_groupi_g16774(csa_tree_add_7_25_groupi_n_4323 ,csa_tree_add_7_25_groupi_n_4322);
  and csa_tree_add_7_25_groupi_g16775(csa_tree_add_7_25_groupi_n_4320 ,csa_tree_add_7_25_groupi_n_4240 ,csa_tree_add_7_25_groupi_n_4222);
  or csa_tree_add_7_25_groupi_g16776(csa_tree_add_7_25_groupi_n_4319 ,in2[11] ,csa_tree_add_7_25_groupi_n_4210);
  or csa_tree_add_7_25_groupi_g16777(csa_tree_add_7_25_groupi_n_4318 ,in2[8] ,csa_tree_add_7_25_groupi_n_4209);
  and csa_tree_add_7_25_groupi_g16778(csa_tree_add_7_25_groupi_n_4317 ,csa_tree_add_7_25_groupi_n_4216 ,csa_tree_add_7_25_groupi_n_4237);
  and csa_tree_add_7_25_groupi_g16779(csa_tree_add_7_25_groupi_n_4316 ,in2[5] ,csa_tree_add_7_25_groupi_n_4208);
  and csa_tree_add_7_25_groupi_g16780(csa_tree_add_7_25_groupi_n_4315 ,in2[26] ,csa_tree_add_7_25_groupi_n_4204);
  and csa_tree_add_7_25_groupi_g16781(csa_tree_add_7_25_groupi_n_4314 ,in2[2] ,csa_tree_add_7_25_groupi_n_4217);
  and csa_tree_add_7_25_groupi_g16782(csa_tree_add_7_25_groupi_n_4313 ,in2[17] ,csa_tree_add_7_25_groupi_n_4213);
  or csa_tree_add_7_25_groupi_g16783(csa_tree_add_7_25_groupi_n_4312 ,in2[17] ,csa_tree_add_7_25_groupi_n_4213);
  and csa_tree_add_7_25_groupi_g16784(csa_tree_add_7_25_groupi_n_4311 ,csa_tree_add_7_25_groupi_n_4244 ,csa_tree_add_7_25_groupi_n_4229);
  or csa_tree_add_7_25_groupi_g16785(csa_tree_add_7_25_groupi_n_4310 ,in2[5] ,csa_tree_add_7_25_groupi_n_4208);
  and csa_tree_add_7_25_groupi_g16786(csa_tree_add_7_25_groupi_n_4309 ,csa_tree_add_7_25_groupi_n_4243 ,csa_tree_add_7_25_groupi_n_4225);
  or csa_tree_add_7_25_groupi_g16787(csa_tree_add_7_25_groupi_n_4308 ,in2[14] ,csa_tree_add_7_25_groupi_n_4211);
  or csa_tree_add_7_25_groupi_g16788(csa_tree_add_7_25_groupi_n_4307 ,in2[29] ,csa_tree_add_7_25_groupi_n_4212);
  or csa_tree_add_7_25_groupi_g16789(csa_tree_add_7_25_groupi_n_4306 ,in2[20] ,csa_tree_add_7_25_groupi_n_4214);
  or csa_tree_add_7_25_groupi_g16790(csa_tree_add_7_25_groupi_n_4305 ,csa_tree_add_7_25_groupi_n_2417 ,csa_tree_add_7_25_groupi_n_4242);
  and csa_tree_add_7_25_groupi_g16791(csa_tree_add_7_25_groupi_n_4304 ,in2[14] ,csa_tree_add_7_25_groupi_n_4211);
  or csa_tree_add_7_25_groupi_g16792(csa_tree_add_7_25_groupi_n_4303 ,in2[26] ,csa_tree_add_7_25_groupi_n_4204);
  and csa_tree_add_7_25_groupi_g16793(csa_tree_add_7_25_groupi_n_4302 ,in2[29] ,csa_tree_add_7_25_groupi_n_4212);
  and csa_tree_add_7_25_groupi_g16794(csa_tree_add_7_25_groupi_n_4301 ,csa_tree_add_7_25_groupi_n_4247 ,csa_tree_add_7_25_groupi_n_4223);
  and csa_tree_add_7_25_groupi_g16795(csa_tree_add_7_25_groupi_n_4300 ,in2[11] ,csa_tree_add_7_25_groupi_n_4210);
  and csa_tree_add_7_25_groupi_g16796(csa_tree_add_7_25_groupi_n_4299 ,csa_tree_add_7_25_groupi_n_4246 ,csa_tree_add_7_25_groupi_n_4235);
  or csa_tree_add_7_25_groupi_g16797(csa_tree_add_7_25_groupi_n_4298 ,in2[23] ,csa_tree_add_7_25_groupi_n_4215);
  and csa_tree_add_7_25_groupi_g16798(csa_tree_add_7_25_groupi_n_4297 ,csa_tree_add_7_25_groupi_n_4248 ,csa_tree_add_7_25_groupi_n_4233);
  and csa_tree_add_7_25_groupi_g16799(csa_tree_add_7_25_groupi_n_4296 ,csa_tree_add_7_25_groupi_n_4249 ,csa_tree_add_7_25_groupi_n_4238);
  nor csa_tree_add_7_25_groupi_g16800(csa_tree_add_7_25_groupi_n_4295 ,csa_tree_add_7_25_groupi_n_4219 ,csa_tree_add_7_25_groupi_n_4227);
  nor csa_tree_add_7_25_groupi_g16801(csa_tree_add_7_25_groupi_n_4294 ,csa_tree_add_7_25_groupi_n_4093 ,csa_tree_add_7_25_groupi_n_4193);
  nor csa_tree_add_7_25_groupi_g16802(csa_tree_add_7_25_groupi_n_4293 ,csa_tree_add_7_25_groupi_n_3843 ,csa_tree_add_7_25_groupi_n_4192);
  nor csa_tree_add_7_25_groupi_g16803(csa_tree_add_7_25_groupi_n_4292 ,csa_tree_add_7_25_groupi_n_4056 ,csa_tree_add_7_25_groupi_n_4197);
  nor csa_tree_add_7_25_groupi_g16804(csa_tree_add_7_25_groupi_n_4291 ,csa_tree_add_7_25_groupi_n_3870 ,csa_tree_add_7_25_groupi_n_4190);
  and csa_tree_add_7_25_groupi_g16805(csa_tree_add_7_25_groupi_n_4322 ,csa_tree_add_7_25_groupi_n_3917 ,csa_tree_add_7_25_groupi_n_4189);
  nor csa_tree_add_7_25_groupi_g16806(csa_tree_add_7_25_groupi_n_4290 ,csa_tree_add_7_25_groupi_n_4081 ,csa_tree_add_7_25_groupi_n_4196);
  nor csa_tree_add_7_25_groupi_g16807(csa_tree_add_7_25_groupi_n_4289 ,csa_tree_add_7_25_groupi_n_3810 ,csa_tree_add_7_25_groupi_n_4191);
  nor csa_tree_add_7_25_groupi_g16808(csa_tree_add_7_25_groupi_n_4288 ,csa_tree_add_7_25_groupi_n_3490 ,csa_tree_add_7_25_groupi_n_4188);
  nor csa_tree_add_7_25_groupi_g16809(csa_tree_add_7_25_groupi_n_4287 ,csa_tree_add_7_25_groupi_n_4036 ,csa_tree_add_7_25_groupi_n_4194);
  and csa_tree_add_7_25_groupi_g16810(csa_tree_add_7_25_groupi_n_4321 ,csa_tree_add_7_25_groupi_n_4139 ,csa_tree_add_7_25_groupi_n_4245);
  and csa_tree_add_7_25_groupi_g16811(csa_tree_add_7_25_groupi_n_4275 ,in2[23] ,csa_tree_add_7_25_groupi_n_4215);
  and csa_tree_add_7_25_groupi_g16812(csa_tree_add_7_25_groupi_n_4274 ,in2[20] ,csa_tree_add_7_25_groupi_n_4214);
  and csa_tree_add_7_25_groupi_g16813(csa_tree_add_7_25_groupi_n_4273 ,csa_tree_add_7_25_groupi_n_4241 ,csa_tree_add_7_25_groupi_n_4228);
  and csa_tree_add_7_25_groupi_g16814(csa_tree_add_7_25_groupi_n_4272 ,in2[8] ,csa_tree_add_7_25_groupi_n_4209);
  nor csa_tree_add_7_25_groupi_g16815(csa_tree_add_7_25_groupi_n_4271 ,csa_tree_add_7_25_groupi_n_549 ,csa_tree_add_7_25_groupi_n_274);
  nor csa_tree_add_7_25_groupi_g16816(csa_tree_add_7_25_groupi_n_4270 ,csa_tree_add_7_25_groupi_n_206 ,csa_tree_add_7_25_groupi_n_1318);
  nor csa_tree_add_7_25_groupi_g16817(csa_tree_add_7_25_groupi_n_4269 ,csa_tree_add_7_25_groupi_n_2169 ,csa_tree_add_7_25_groupi_n_1873);
  nor csa_tree_add_7_25_groupi_g16818(csa_tree_add_7_25_groupi_n_4268 ,csa_tree_add_7_25_groupi_n_1873 ,csa_tree_add_7_25_groupi_n_1796);
  nor csa_tree_add_7_25_groupi_g16819(csa_tree_add_7_25_groupi_n_4267 ,csa_tree_add_7_25_groupi_n_327 ,csa_tree_add_7_25_groupi_n_2025);
  nor csa_tree_add_7_25_groupi_g16820(csa_tree_add_7_25_groupi_n_4266 ,csa_tree_add_7_25_groupi_n_327 ,csa_tree_add_7_25_groupi_n_2051);
  nor csa_tree_add_7_25_groupi_g16821(csa_tree_add_7_25_groupi_n_4265 ,csa_tree_add_7_25_groupi_n_274 ,csa_tree_add_7_25_groupi_n_2054);
  nor csa_tree_add_7_25_groupi_g16822(csa_tree_add_7_25_groupi_n_4264 ,csa_tree_add_7_25_groupi_n_326 ,csa_tree_add_7_25_groupi_n_2166);
  nor csa_tree_add_7_25_groupi_g16823(csa_tree_add_7_25_groupi_n_4263 ,csa_tree_add_7_25_groupi_n_2091 ,csa_tree_add_7_25_groupi_n_206);
  nor csa_tree_add_7_25_groupi_g16824(csa_tree_add_7_25_groupi_n_4262 ,csa_tree_add_7_25_groupi_n_273 ,csa_tree_add_7_25_groupi_n_2145);
  nor csa_tree_add_7_25_groupi_g16825(csa_tree_add_7_25_groupi_n_4261 ,csa_tree_add_7_25_groupi_n_2112 ,csa_tree_add_7_25_groupi_n_1872);
  nor csa_tree_add_7_25_groupi_g16826(csa_tree_add_7_25_groupi_n_4260 ,in2[2] ,csa_tree_add_7_25_groupi_n_4217);
  nor csa_tree_add_7_25_groupi_g16827(csa_tree_add_7_25_groupi_n_4259 ,csa_tree_add_7_25_groupi_n_3986 ,csa_tree_add_7_25_groupi_n_4187);
  xnor csa_tree_add_7_25_groupi_g16828(csa_tree_add_7_25_groupi_n_4258 ,csa_tree_add_7_25_groupi_n_4153 ,in2[28]);
  nor csa_tree_add_7_25_groupi_g16829(csa_tree_add_7_25_groupi_n_4257 ,csa_tree_add_7_25_groupi_n_4069 ,csa_tree_add_7_25_groupi_n_4195);
  xnor csa_tree_add_7_25_groupi_g16830(csa_tree_add_7_25_groupi_n_4256 ,csa_tree_add_7_25_groupi_n_4162 ,in2[25]);
  xnor csa_tree_add_7_25_groupi_g16831(csa_tree_add_7_25_groupi_n_4255 ,csa_tree_add_7_25_groupi_n_4161 ,in2[22]);
  xnor csa_tree_add_7_25_groupi_g16832(csa_tree_add_7_25_groupi_n_4254 ,csa_tree_add_7_25_groupi_n_4157 ,in2[19]);
  xnor csa_tree_add_7_25_groupi_g16833(csa_tree_add_7_25_groupi_n_4253 ,csa_tree_add_7_25_groupi_n_4158 ,in2[16]);
  xnor csa_tree_add_7_25_groupi_g16834(csa_tree_add_7_25_groupi_n_4252 ,csa_tree_add_7_25_groupi_n_4156 ,in2[10]);
  xnor csa_tree_add_7_25_groupi_g16835(csa_tree_add_7_25_groupi_n_4251 ,csa_tree_add_7_25_groupi_n_4155 ,in2[7]);
  xnor csa_tree_add_7_25_groupi_g16836(csa_tree_add_7_25_groupi_n_4286 ,csa_tree_add_7_25_groupi_n_4167 ,in3[2]);
  xnor csa_tree_add_7_25_groupi_g16837(csa_tree_add_7_25_groupi_n_4250 ,csa_tree_add_7_25_groupi_n_4154 ,in2[13]);
  xnor csa_tree_add_7_25_groupi_g16838(csa_tree_add_7_25_groupi_n_4285 ,csa_tree_add_7_25_groupi_n_4170 ,in3[5]);
  xnor csa_tree_add_7_25_groupi_g16839(csa_tree_add_7_25_groupi_n_4284 ,csa_tree_add_7_25_groupi_n_4168 ,in3[8]);
  xnor csa_tree_add_7_25_groupi_g16840(csa_tree_add_7_25_groupi_n_4283 ,csa_tree_add_7_25_groupi_n_4140 ,in3[11]);
  xnor csa_tree_add_7_25_groupi_g16841(csa_tree_add_7_25_groupi_n_4282 ,csa_tree_add_7_25_groupi_n_4165 ,in3[14]);
  xnor csa_tree_add_7_25_groupi_g16842(csa_tree_add_7_25_groupi_n_4281 ,csa_tree_add_7_25_groupi_n_4164 ,in3[17]);
  xnor csa_tree_add_7_25_groupi_g16843(csa_tree_add_7_25_groupi_n_4280 ,csa_tree_add_7_25_groupi_n_4169 ,in3[20]);
  xnor csa_tree_add_7_25_groupi_g16844(csa_tree_add_7_25_groupi_n_4279 ,csa_tree_add_7_25_groupi_n_4171 ,in3[23]);
  xnor csa_tree_add_7_25_groupi_g16845(csa_tree_add_7_25_groupi_n_4278 ,csa_tree_add_7_25_groupi_n_4172 ,in3[26]);
  xnor csa_tree_add_7_25_groupi_g16846(csa_tree_add_7_25_groupi_n_4277 ,csa_tree_add_7_25_groupi_n_4166 ,in3[29]);
  xnor csa_tree_add_7_25_groupi_g16847(csa_tree_add_7_25_groupi_n_4276 ,csa_tree_add_7_25_groupi_n_4100 ,csa_tree_add_7_25_groupi_n_4141);
  nor csa_tree_add_7_25_groupi_g16848(csa_tree_add_7_25_groupi_n_4239 ,csa_tree_add_7_25_groupi_n_2413 ,csa_tree_add_7_25_groupi_n_4160);
  or csa_tree_add_7_25_groupi_g16849(csa_tree_add_7_25_groupi_n_4238 ,in2[4] ,csa_tree_add_7_25_groupi_n_4159);
  or csa_tree_add_7_25_groupi_g16850(csa_tree_add_7_25_groupi_n_4237 ,in2[13] ,csa_tree_add_7_25_groupi_n_4154);
  and csa_tree_add_7_25_groupi_g16851(csa_tree_add_7_25_groupi_n_4236 ,in2[10] ,csa_tree_add_7_25_groupi_n_4156);
  or csa_tree_add_7_25_groupi_g16852(csa_tree_add_7_25_groupi_n_4235 ,in2[10] ,csa_tree_add_7_25_groupi_n_4156);
  and csa_tree_add_7_25_groupi_g16853(csa_tree_add_7_25_groupi_n_4234 ,in2[7] ,csa_tree_add_7_25_groupi_n_4155);
  or csa_tree_add_7_25_groupi_g16854(csa_tree_add_7_25_groupi_n_4233 ,in2[7] ,csa_tree_add_7_25_groupi_n_4155);
  and csa_tree_add_7_25_groupi_g16855(csa_tree_add_7_25_groupi_n_4232 ,in2[13] ,csa_tree_add_7_25_groupi_n_4154);
  and csa_tree_add_7_25_groupi_g16856(csa_tree_add_7_25_groupi_n_4231 ,in2[16] ,csa_tree_add_7_25_groupi_n_4158);
  and csa_tree_add_7_25_groupi_g16857(csa_tree_add_7_25_groupi_n_4230 ,in2[19] ,csa_tree_add_7_25_groupi_n_4157);
  or csa_tree_add_7_25_groupi_g16858(csa_tree_add_7_25_groupi_n_4229 ,in2[16] ,csa_tree_add_7_25_groupi_n_4158);
  or csa_tree_add_7_25_groupi_g16859(csa_tree_add_7_25_groupi_n_4228 ,in2[19] ,csa_tree_add_7_25_groupi_n_4157);
  nor csa_tree_add_7_25_groupi_g16860(csa_tree_add_7_25_groupi_n_4227 ,in2[1] ,csa_tree_add_7_25_groupi_n_4163);
  and csa_tree_add_7_25_groupi_g16861(csa_tree_add_7_25_groupi_n_4226 ,in2[1] ,csa_tree_add_7_25_groupi_n_4163);
  or csa_tree_add_7_25_groupi_g16862(csa_tree_add_7_25_groupi_n_4225 ,in2[28] ,csa_tree_add_7_25_groupi_n_4153);
  and csa_tree_add_7_25_groupi_g16863(csa_tree_add_7_25_groupi_n_4224 ,in2[28] ,csa_tree_add_7_25_groupi_n_4153);
  or csa_tree_add_7_25_groupi_g16864(csa_tree_add_7_25_groupi_n_4223 ,in2[22] ,csa_tree_add_7_25_groupi_n_4161);
  or csa_tree_add_7_25_groupi_g16865(csa_tree_add_7_25_groupi_n_4222 ,in2[25] ,csa_tree_add_7_25_groupi_n_4162);
  and csa_tree_add_7_25_groupi_g16866(csa_tree_add_7_25_groupi_n_4221 ,in2[22] ,csa_tree_add_7_25_groupi_n_4161);
  and csa_tree_add_7_25_groupi_g16867(csa_tree_add_7_25_groupi_n_4220 ,in2[25] ,csa_tree_add_7_25_groupi_n_4162);
  nor csa_tree_add_7_25_groupi_g16868(csa_tree_add_7_25_groupi_n_4219 ,csa_tree_add_7_25_groupi_n_2496 ,csa_tree_add_7_25_groupi_n_4174);
  or csa_tree_add_7_25_groupi_g16869(csa_tree_add_7_25_groupi_n_4249 ,csa_tree_add_7_25_groupi_n_2442 ,csa_tree_add_7_25_groupi_n_4184);
  or csa_tree_add_7_25_groupi_g16870(csa_tree_add_7_25_groupi_n_4248 ,csa_tree_add_7_25_groupi_n_2454 ,csa_tree_add_7_25_groupi_n_4176);
  or csa_tree_add_7_25_groupi_g16871(csa_tree_add_7_25_groupi_n_4247 ,csa_tree_add_7_25_groupi_n_2488 ,csa_tree_add_7_25_groupi_n_4179);
  or csa_tree_add_7_25_groupi_g16872(csa_tree_add_7_25_groupi_n_4246 ,csa_tree_add_7_25_groupi_n_2446 ,csa_tree_add_7_25_groupi_n_4178);
  or csa_tree_add_7_25_groupi_g16873(csa_tree_add_7_25_groupi_n_4245 ,csa_tree_add_7_25_groupi_n_4135 ,csa_tree_add_7_25_groupi_n_4175);
  or csa_tree_add_7_25_groupi_g16874(csa_tree_add_7_25_groupi_n_4244 ,csa_tree_add_7_25_groupi_n_2425 ,csa_tree_add_7_25_groupi_n_4183);
  or csa_tree_add_7_25_groupi_g16875(csa_tree_add_7_25_groupi_n_4243 ,csa_tree_add_7_25_groupi_n_2431 ,csa_tree_add_7_25_groupi_n_4180);
  and csa_tree_add_7_25_groupi_g16876(csa_tree_add_7_25_groupi_n_4242 ,csa_tree_add_7_25_groupi_n_2430 ,csa_tree_add_7_25_groupi_n_4173);
  or csa_tree_add_7_25_groupi_g16877(csa_tree_add_7_25_groupi_n_4241 ,csa_tree_add_7_25_groupi_n_2471 ,csa_tree_add_7_25_groupi_n_4182);
  or csa_tree_add_7_25_groupi_g16878(csa_tree_add_7_25_groupi_n_4240 ,csa_tree_add_7_25_groupi_n_2437 ,csa_tree_add_7_25_groupi_n_4181);
  or csa_tree_add_7_25_groupi_g16879(csa_tree_add_7_25_groupi_n_4197 ,csa_tree_add_7_25_groupi_n_3109 ,csa_tree_add_7_25_groupi_n_4144);
  or csa_tree_add_7_25_groupi_g16880(csa_tree_add_7_25_groupi_n_4196 ,csa_tree_add_7_25_groupi_n_3155 ,csa_tree_add_7_25_groupi_n_4152);
  or csa_tree_add_7_25_groupi_g16881(csa_tree_add_7_25_groupi_n_4195 ,csa_tree_add_7_25_groupi_n_3136 ,csa_tree_add_7_25_groupi_n_4146);
  or csa_tree_add_7_25_groupi_g16882(csa_tree_add_7_25_groupi_n_4194 ,csa_tree_add_7_25_groupi_n_3132 ,csa_tree_add_7_25_groupi_n_4145);
  or csa_tree_add_7_25_groupi_g16883(csa_tree_add_7_25_groupi_n_4193 ,csa_tree_add_7_25_groupi_n_3102 ,csa_tree_add_7_25_groupi_n_4143);
  or csa_tree_add_7_25_groupi_g16884(csa_tree_add_7_25_groupi_n_4192 ,csa_tree_add_7_25_groupi_n_3645 ,csa_tree_add_7_25_groupi_n_4147);
  or csa_tree_add_7_25_groupi_g16885(csa_tree_add_7_25_groupi_n_4191 ,csa_tree_add_7_25_groupi_n_3642 ,csa_tree_add_7_25_groupi_n_4150);
  or csa_tree_add_7_25_groupi_g16886(csa_tree_add_7_25_groupi_n_4190 ,csa_tree_add_7_25_groupi_n_3577 ,csa_tree_add_7_25_groupi_n_4149);
  nor csa_tree_add_7_25_groupi_g16887(csa_tree_add_7_25_groupi_n_4189 ,csa_tree_add_7_25_groupi_n_3038 ,csa_tree_add_7_25_groupi_n_4142);
  or csa_tree_add_7_25_groupi_g16888(csa_tree_add_7_25_groupi_n_4188 ,csa_tree_add_7_25_groupi_n_3009 ,csa_tree_add_7_25_groupi_n_4151);
  or csa_tree_add_7_25_groupi_g16889(csa_tree_add_7_25_groupi_n_4187 ,csa_tree_add_7_25_groupi_n_3180 ,csa_tree_add_7_25_groupi_n_4148);
  xnor csa_tree_add_7_25_groupi_g16890(csa_tree_add_7_25_groupi_n_4218 ,csa_tree_add_7_25_groupi_n_4116 ,csa_tree_add_7_25_groupi_n_2594);
  xnor csa_tree_add_7_25_groupi_g16891(csa_tree_add_7_25_groupi_n_4217 ,csa_tree_add_7_25_groupi_n_4130 ,in3[2]);
  or csa_tree_add_7_25_groupi_g16892(csa_tree_add_7_25_groupi_n_4216 ,csa_tree_add_7_25_groupi_n_2455 ,csa_tree_add_7_25_groupi_n_4177);
  xnor csa_tree_add_7_25_groupi_g16893(csa_tree_add_7_25_groupi_n_4215 ,csa_tree_add_7_25_groupi_n_4129 ,in3[23]);
  xnor csa_tree_add_7_25_groupi_g16894(csa_tree_add_7_25_groupi_n_4214 ,csa_tree_add_7_25_groupi_n_4126 ,in3[20]);
  xnor csa_tree_add_7_25_groupi_g16895(csa_tree_add_7_25_groupi_n_4213 ,csa_tree_add_7_25_groupi_n_4121 ,in3[17]);
  xnor csa_tree_add_7_25_groupi_g16896(csa_tree_add_7_25_groupi_n_4212 ,csa_tree_add_7_25_groupi_n_4128 ,in3[29]);
  xnor csa_tree_add_7_25_groupi_g16897(csa_tree_add_7_25_groupi_n_4211 ,csa_tree_add_7_25_groupi_n_4123 ,in3[14]);
  xnor csa_tree_add_7_25_groupi_g16898(csa_tree_add_7_25_groupi_n_4210 ,csa_tree_add_7_25_groupi_n_4125 ,in3[11]);
  xnor csa_tree_add_7_25_groupi_g16899(csa_tree_add_7_25_groupi_n_4209 ,csa_tree_add_7_25_groupi_n_4127 ,in3[8]);
  xnor csa_tree_add_7_25_groupi_g16900(csa_tree_add_7_25_groupi_n_4208 ,csa_tree_add_7_25_groupi_n_4122 ,in3[5]);
  xnor csa_tree_add_7_25_groupi_g16901(csa_tree_add_7_25_groupi_n_4207 ,csa_tree_add_7_25_groupi_n_4117 ,csa_tree_add_7_25_groupi_n_2596);
  xnor csa_tree_add_7_25_groupi_g16902(csa_tree_add_7_25_groupi_n_4206 ,csa_tree_add_7_25_groupi_n_4120 ,csa_tree_add_7_25_groupi_n_2593);
  xnor csa_tree_add_7_25_groupi_g16903(csa_tree_add_7_25_groupi_n_4205 ,csa_tree_add_7_25_groupi_n_4118 ,csa_tree_add_7_25_groupi_n_2595);
  xnor csa_tree_add_7_25_groupi_g16904(csa_tree_add_7_25_groupi_n_4204 ,csa_tree_add_7_25_groupi_n_4124 ,in3[26]);
  xnor csa_tree_add_7_25_groupi_g16905(csa_tree_add_7_25_groupi_n_4203 ,csa_tree_add_7_25_groupi_n_4115 ,csa_tree_add_7_25_groupi_n_2592);
  xnor csa_tree_add_7_25_groupi_g16906(csa_tree_add_7_25_groupi_n_4202 ,csa_tree_add_7_25_groupi_n_4114 ,csa_tree_add_7_25_groupi_n_2591);
  xnor csa_tree_add_7_25_groupi_g16907(csa_tree_add_7_25_groupi_n_4201 ,csa_tree_add_7_25_groupi_n_4113 ,csa_tree_add_7_25_groupi_n_2590);
  xnor csa_tree_add_7_25_groupi_g16908(csa_tree_add_7_25_groupi_n_4200 ,csa_tree_add_7_25_groupi_n_4112 ,csa_tree_add_7_25_groupi_n_2589);
  xnor csa_tree_add_7_25_groupi_g16909(csa_tree_add_7_25_groupi_n_4199 ,csa_tree_add_7_25_groupi_n_4119 ,csa_tree_add_7_25_groupi_n_2588);
  xnor csa_tree_add_7_25_groupi_g16910(csa_tree_add_7_25_groupi_n_4198 ,csa_tree_add_7_25_groupi_n_4137 ,csa_tree_add_7_25_groupi_n_2577);
  not csa_tree_add_7_25_groupi_g16911(csa_tree_add_7_25_groupi_n_4186 ,csa_tree_add_7_25_groupi_n_4185);
  and csa_tree_add_7_25_groupi_g16912(csa_tree_add_7_25_groupi_n_4184 ,csa_tree_add_7_25_groupi_n_2462 ,csa_tree_add_7_25_groupi_n_4116);
  and csa_tree_add_7_25_groupi_g16913(csa_tree_add_7_25_groupi_n_4183 ,csa_tree_add_7_25_groupi_n_2427 ,csa_tree_add_7_25_groupi_n_4115);
  and csa_tree_add_7_25_groupi_g16914(csa_tree_add_7_25_groupi_n_4182 ,csa_tree_add_7_25_groupi_n_2459 ,csa_tree_add_7_25_groupi_n_4114);
  and csa_tree_add_7_25_groupi_g16915(csa_tree_add_7_25_groupi_n_4181 ,csa_tree_add_7_25_groupi_n_2418 ,csa_tree_add_7_25_groupi_n_4112);
  and csa_tree_add_7_25_groupi_g16916(csa_tree_add_7_25_groupi_n_4180 ,csa_tree_add_7_25_groupi_n_2450 ,csa_tree_add_7_25_groupi_n_4119);
  and csa_tree_add_7_25_groupi_g16917(csa_tree_add_7_25_groupi_n_4179 ,csa_tree_add_7_25_groupi_n_2484 ,csa_tree_add_7_25_groupi_n_4113);
  and csa_tree_add_7_25_groupi_g16918(csa_tree_add_7_25_groupi_n_4178 ,csa_tree_add_7_25_groupi_n_2472 ,csa_tree_add_7_25_groupi_n_4117);
  and csa_tree_add_7_25_groupi_g16919(csa_tree_add_7_25_groupi_n_4177 ,csa_tree_add_7_25_groupi_n_2419 ,csa_tree_add_7_25_groupi_n_4120);
  and csa_tree_add_7_25_groupi_g16920(csa_tree_add_7_25_groupi_n_4176 ,csa_tree_add_7_25_groupi_n_2458 ,csa_tree_add_7_25_groupi_n_4118);
  nor csa_tree_add_7_25_groupi_g16921(csa_tree_add_7_25_groupi_n_4175 ,csa_tree_add_7_25_groupi_n_4101 ,csa_tree_add_7_25_groupi_n_4131);
  nor csa_tree_add_7_25_groupi_g16922(csa_tree_add_7_25_groupi_n_4174 ,csa_tree_add_7_25_groupi_n_2479 ,csa_tree_add_7_25_groupi_n_4103);
  or csa_tree_add_7_25_groupi_g16923(csa_tree_add_7_25_groupi_n_4173 ,csa_tree_add_7_25_groupi_n_2494 ,csa_tree_add_7_25_groupi_n_4137);
  nor csa_tree_add_7_25_groupi_g16924(csa_tree_add_7_25_groupi_n_4172 ,csa_tree_add_7_25_groupi_n_3932 ,csa_tree_add_7_25_groupi_n_4134);
  nor csa_tree_add_7_25_groupi_g16925(csa_tree_add_7_25_groupi_n_4171 ,csa_tree_add_7_25_groupi_n_3812 ,csa_tree_add_7_25_groupi_n_4105);
  nor csa_tree_add_7_25_groupi_g16926(csa_tree_add_7_25_groupi_n_4170 ,csa_tree_add_7_25_groupi_n_4004 ,csa_tree_add_7_25_groupi_n_4102);
  nor csa_tree_add_7_25_groupi_g16927(csa_tree_add_7_25_groupi_n_4169 ,csa_tree_add_7_25_groupi_n_3984 ,csa_tree_add_7_25_groupi_n_4133);
  nor csa_tree_add_7_25_groupi_g16928(csa_tree_add_7_25_groupi_n_4168 ,csa_tree_add_7_25_groupi_n_4072 ,csa_tree_add_7_25_groupi_n_4107);
  nor csa_tree_add_7_25_groupi_g16929(csa_tree_add_7_25_groupi_n_4167 ,csa_tree_add_7_25_groupi_n_3480 ,csa_tree_add_7_25_groupi_n_4104);
  nor csa_tree_add_7_25_groupi_g16930(csa_tree_add_7_25_groupi_n_4166 ,csa_tree_add_7_25_groupi_n_3839 ,csa_tree_add_7_25_groupi_n_4132);
  nor csa_tree_add_7_25_groupi_g16931(csa_tree_add_7_25_groupi_n_4165 ,csa_tree_add_7_25_groupi_n_4055 ,csa_tree_add_7_25_groupi_n_4106);
  nor csa_tree_add_7_25_groupi_g16932(csa_tree_add_7_25_groupi_n_4164 ,csa_tree_add_7_25_groupi_n_4075 ,csa_tree_add_7_25_groupi_n_4136);
  and csa_tree_add_7_25_groupi_g16933(csa_tree_add_7_25_groupi_n_4185 ,csa_tree_add_7_25_groupi_n_3927 ,csa_tree_add_7_25_groupi_n_4109);
  not csa_tree_add_7_25_groupi_g16934(csa_tree_add_7_25_groupi_n_4159 ,csa_tree_add_7_25_groupi_n_4160);
  nor csa_tree_add_7_25_groupi_g16935(csa_tree_add_7_25_groupi_n_4152 ,csa_tree_add_7_25_groupi_n_324 ,csa_tree_add_7_25_groupi_n_2060);
  nor csa_tree_add_7_25_groupi_g16936(csa_tree_add_7_25_groupi_n_4151 ,csa_tree_add_7_25_groupi_n_2186 ,csa_tree_add_7_25_groupi_n_1833);
  nor csa_tree_add_7_25_groupi_g16937(csa_tree_add_7_25_groupi_n_4150 ,csa_tree_add_7_25_groupi_n_379 ,csa_tree_add_7_25_groupi_n_1833);
  nor csa_tree_add_7_25_groupi_g16938(csa_tree_add_7_25_groupi_n_4149 ,csa_tree_add_7_25_groupi_n_2028 ,csa_tree_add_7_25_groupi_n_159);
  nor csa_tree_add_7_25_groupi_g16939(csa_tree_add_7_25_groupi_n_4148 ,csa_tree_add_7_25_groupi_n_248 ,csa_tree_add_7_25_groupi_n_2046);
  nor csa_tree_add_7_25_groupi_g16940(csa_tree_add_7_25_groupi_n_4147 ,csa_tree_add_7_25_groupi_n_241 ,csa_tree_add_7_25_groupi_n_249);
  nor csa_tree_add_7_25_groupi_g16941(csa_tree_add_7_25_groupi_n_4146 ,csa_tree_add_7_25_groupi_n_249 ,csa_tree_add_7_25_groupi_n_2138);
  nor csa_tree_add_7_25_groupi_g16942(csa_tree_add_7_25_groupi_n_4145 ,csa_tree_add_7_25_groupi_n_324 ,csa_tree_add_7_25_groupi_n_2159);
  nor csa_tree_add_7_25_groupi_g16943(csa_tree_add_7_25_groupi_n_4144 ,csa_tree_add_7_25_groupi_n_2105 ,csa_tree_add_7_25_groupi_n_1834);
  nor csa_tree_add_7_25_groupi_g16944(csa_tree_add_7_25_groupi_n_4143 ,csa_tree_add_7_25_groupi_n_323 ,csa_tree_add_7_25_groupi_n_2126);
  nor csa_tree_add_7_25_groupi_g16945(csa_tree_add_7_25_groupi_n_4142 ,csa_tree_add_7_25_groupi_n_636 ,csa_tree_add_7_25_groupi_n_159);
  xnor csa_tree_add_7_25_groupi_g16946(csa_tree_add_7_25_groupi_n_4141 ,csa_tree_add_7_25_groupi_n_4101 ,in2[31]);
  xnor csa_tree_add_7_25_groupi_g16947(csa_tree_add_7_25_groupi_n_4163 ,csa_tree_add_7_25_groupi_n_1092 ,csa_tree_add_7_25_groupi_n_3951);
  nor csa_tree_add_7_25_groupi_g16948(csa_tree_add_7_25_groupi_n_4140 ,csa_tree_add_7_25_groupi_n_3980 ,csa_tree_add_7_25_groupi_n_4108);
  xnor csa_tree_add_7_25_groupi_g16949(csa_tree_add_7_25_groupi_n_4162 ,csa_tree_add_7_25_groupi_n_4027 ,in3[26]);
  xnor csa_tree_add_7_25_groupi_g16950(csa_tree_add_7_25_groupi_n_4161 ,csa_tree_add_7_25_groupi_n_3959 ,in3[23]);
  xnor csa_tree_add_7_25_groupi_g16951(csa_tree_add_7_25_groupi_n_4160 ,csa_tree_add_7_25_groupi_n_3955 ,in3[5]);
  xnor csa_tree_add_7_25_groupi_g16952(csa_tree_add_7_25_groupi_n_4158 ,csa_tree_add_7_25_groupi_n_3954 ,in3[17]);
  xnor csa_tree_add_7_25_groupi_g16953(csa_tree_add_7_25_groupi_n_4157 ,csa_tree_add_7_25_groupi_n_3953 ,in3[20]);
  xnor csa_tree_add_7_25_groupi_g16954(csa_tree_add_7_25_groupi_n_4156 ,csa_tree_add_7_25_groupi_n_3956 ,in3[11]);
  xnor csa_tree_add_7_25_groupi_g16955(csa_tree_add_7_25_groupi_n_4155 ,csa_tree_add_7_25_groupi_n_3957 ,in3[8]);
  xnor csa_tree_add_7_25_groupi_g16956(csa_tree_add_7_25_groupi_n_4154 ,csa_tree_add_7_25_groupi_n_3958 ,in3[14]);
  xnor csa_tree_add_7_25_groupi_g16957(csa_tree_add_7_25_groupi_n_4153 ,csa_tree_add_7_25_groupi_n_3952 ,in3[29]);
  not csa_tree_add_7_25_groupi_g16958(csa_tree_add_7_25_groupi_n_4139 ,csa_tree_add_7_25_groupi_n_4138);
  or csa_tree_add_7_25_groupi_g16959(csa_tree_add_7_25_groupi_n_4136 ,csa_tree_add_7_25_groupi_n_3150 ,csa_tree_add_7_25_groupi_n_3977);
  nor csa_tree_add_7_25_groupi_g16960(csa_tree_add_7_25_groupi_n_4135 ,csa_tree_add_7_25_groupi_n_2412 ,csa_tree_add_7_25_groupi_n_4100);
  or csa_tree_add_7_25_groupi_g16961(csa_tree_add_7_25_groupi_n_4134 ,csa_tree_add_7_25_groupi_n_3679 ,csa_tree_add_7_25_groupi_n_3974);
  or csa_tree_add_7_25_groupi_g16962(csa_tree_add_7_25_groupi_n_4133 ,csa_tree_add_7_25_groupi_n_3176 ,csa_tree_add_7_25_groupi_n_3976);
  or csa_tree_add_7_25_groupi_g16963(csa_tree_add_7_25_groupi_n_4132 ,csa_tree_add_7_25_groupi_n_3673 ,csa_tree_add_7_25_groupi_n_3960);
  and csa_tree_add_7_25_groupi_g16964(csa_tree_add_7_25_groupi_n_4131 ,csa_tree_add_7_25_groupi_n_2412 ,csa_tree_add_7_25_groupi_n_4100);
  nor csa_tree_add_7_25_groupi_g16965(csa_tree_add_7_25_groupi_n_4130 ,csa_tree_add_7_25_groupi_n_3483 ,csa_tree_add_7_25_groupi_n_3962);
  nor csa_tree_add_7_25_groupi_g16966(csa_tree_add_7_25_groupi_n_4129 ,csa_tree_add_7_25_groupi_n_3838 ,csa_tree_add_7_25_groupi_n_3968);
  nor csa_tree_add_7_25_groupi_g16967(csa_tree_add_7_25_groupi_n_4128 ,csa_tree_add_7_25_groupi_n_3836 ,csa_tree_add_7_25_groupi_n_3970);
  nor csa_tree_add_7_25_groupi_g16968(csa_tree_add_7_25_groupi_n_4127 ,csa_tree_add_7_25_groupi_n_3849 ,csa_tree_add_7_25_groupi_n_3971);
  nor csa_tree_add_7_25_groupi_g16969(csa_tree_add_7_25_groupi_n_4126 ,csa_tree_add_7_25_groupi_n_3896 ,csa_tree_add_7_25_groupi_n_3966);
  nor csa_tree_add_7_25_groupi_g16970(csa_tree_add_7_25_groupi_n_4125 ,csa_tree_add_7_25_groupi_n_3920 ,csa_tree_add_7_25_groupi_n_3973);
  nor csa_tree_add_7_25_groupi_g16971(csa_tree_add_7_25_groupi_n_4124 ,csa_tree_add_7_25_groupi_n_3902 ,csa_tree_add_7_25_groupi_n_3967);
  nor csa_tree_add_7_25_groupi_g16972(csa_tree_add_7_25_groupi_n_4123 ,csa_tree_add_7_25_groupi_n_3943 ,csa_tree_add_7_25_groupi_n_3969);
  nor csa_tree_add_7_25_groupi_g16973(csa_tree_add_7_25_groupi_n_4122 ,csa_tree_add_7_25_groupi_n_4031 ,csa_tree_add_7_25_groupi_n_3964);
  nor csa_tree_add_7_25_groupi_g16974(csa_tree_add_7_25_groupi_n_4121 ,csa_tree_add_7_25_groupi_n_3890 ,csa_tree_add_7_25_groupi_n_3972);
  and csa_tree_add_7_25_groupi_g16975(csa_tree_add_7_25_groupi_n_4138 ,csa_tree_add_7_25_groupi_n_3935 ,csa_tree_add_7_25_groupi_n_3965);
  and csa_tree_add_7_25_groupi_g16976(csa_tree_add_7_25_groupi_n_4137 ,csa_tree_add_7_25_groupi_n_2416 ,csa_tree_add_7_25_groupi_n_4001);
  nor csa_tree_add_7_25_groupi_g16977(csa_tree_add_7_25_groupi_n_4109 ,csa_tree_add_7_25_groupi_n_3043 ,csa_tree_add_7_25_groupi_n_3961);
  or csa_tree_add_7_25_groupi_g16978(csa_tree_add_7_25_groupi_n_4108 ,csa_tree_add_7_25_groupi_n_3130 ,csa_tree_add_7_25_groupi_n_4020);
  or csa_tree_add_7_25_groupi_g16979(csa_tree_add_7_25_groupi_n_4107 ,csa_tree_add_7_25_groupi_n_3119 ,csa_tree_add_7_25_groupi_n_3979);
  or csa_tree_add_7_25_groupi_g16980(csa_tree_add_7_25_groupi_n_4106 ,csa_tree_add_7_25_groupi_n_3106 ,csa_tree_add_7_25_groupi_n_3985);
  or csa_tree_add_7_25_groupi_g16981(csa_tree_add_7_25_groupi_n_4105 ,csa_tree_add_7_25_groupi_n_3669 ,csa_tree_add_7_25_groupi_n_3975);
  or csa_tree_add_7_25_groupi_g16982(csa_tree_add_7_25_groupi_n_4104 ,csa_tree_add_7_25_groupi_n_3041 ,csa_tree_add_7_25_groupi_n_3963);
  xnor csa_tree_add_7_25_groupi_g16983(csa_tree_add_7_25_groupi_n_4103 ,csa_tree_add_7_25_groupi_n_1226 ,csa_tree_add_7_25_groupi_n_3744);
  or csa_tree_add_7_25_groupi_g16984(csa_tree_add_7_25_groupi_n_4102 ,csa_tree_add_7_25_groupi_n_3140 ,csa_tree_add_7_25_groupi_n_3978);
  xnor csa_tree_add_7_25_groupi_g16985(csa_tree_add_7_25_groupi_n_4120 ,csa_tree_add_7_25_groupi_n_3539 ,in3[14]);
  xnor csa_tree_add_7_25_groupi_g16986(csa_tree_add_7_25_groupi_n_4119 ,csa_tree_add_7_25_groupi_n_3542 ,in3[29]);
  xnor csa_tree_add_7_25_groupi_g16987(csa_tree_add_7_25_groupi_n_4118 ,csa_tree_add_7_25_groupi_n_3540 ,in3[8]);
  xnor csa_tree_add_7_25_groupi_g16988(csa_tree_add_7_25_groupi_n_4117 ,csa_tree_add_7_25_groupi_n_3543 ,in3[11]);
  xnor csa_tree_add_7_25_groupi_g16989(csa_tree_add_7_25_groupi_n_4116 ,csa_tree_add_7_25_groupi_n_3537 ,in3[5]);
  xnor csa_tree_add_7_25_groupi_g16990(csa_tree_add_7_25_groupi_n_4115 ,csa_tree_add_7_25_groupi_n_3544 ,in3[17]);
  xnor csa_tree_add_7_25_groupi_g16991(csa_tree_add_7_25_groupi_n_4114 ,csa_tree_add_7_25_groupi_n_3538 ,in3[20]);
  xnor csa_tree_add_7_25_groupi_g16992(csa_tree_add_7_25_groupi_n_4113 ,csa_tree_add_7_25_groupi_n_3541 ,in3[23]);
  xnor csa_tree_add_7_25_groupi_g16993(csa_tree_add_7_25_groupi_n_4112 ,csa_tree_add_7_25_groupi_n_3536 ,in3[26]);
  xnor csa_tree_add_7_25_groupi_g16994(csa_tree_add_7_25_groupi_n_4111 ,csa_tree_add_7_25_groupi_n_3743 ,in2[30]);
  xnor csa_tree_add_7_25_groupi_g16995(csa_tree_add_7_25_groupi_n_4110 ,csa_tree_add_7_25_groupi_n_3950 ,csa_tree_add_7_25_groupi_n_2581);
  or csa_tree_add_7_25_groupi_g16996(csa_tree_add_7_25_groupi_n_4099 ,csa_tree_add_7_25_groupi_n_3260 ,csa_tree_add_7_25_groupi_n_3799);
  or csa_tree_add_7_25_groupi_g16997(csa_tree_add_7_25_groupi_n_4098 ,csa_tree_add_7_25_groupi_n_3057 ,csa_tree_add_7_25_groupi_n_3662);
  or csa_tree_add_7_25_groupi_g16998(csa_tree_add_7_25_groupi_n_4097 ,csa_tree_add_7_25_groupi_n_3194 ,csa_tree_add_7_25_groupi_n_3704);
  or csa_tree_add_7_25_groupi_g16999(csa_tree_add_7_25_groupi_n_4096 ,csa_tree_add_7_25_groupi_n_3095 ,csa_tree_add_7_25_groupi_n_3689);
  or csa_tree_add_7_25_groupi_g17000(csa_tree_add_7_25_groupi_n_4095 ,csa_tree_add_7_25_groupi_n_2927 ,csa_tree_add_7_25_groupi_n_3651);
  or csa_tree_add_7_25_groupi_g17001(csa_tree_add_7_25_groupi_n_4094 ,csa_tree_add_7_25_groupi_n_3160 ,csa_tree_add_7_25_groupi_n_3697);
  or csa_tree_add_7_25_groupi_g17002(csa_tree_add_7_25_groupi_n_4093 ,csa_tree_add_7_25_groupi_n_2934 ,csa_tree_add_7_25_groupi_n_3648);
  or csa_tree_add_7_25_groupi_g17003(csa_tree_add_7_25_groupi_n_4092 ,csa_tree_add_7_25_groupi_n_3276 ,csa_tree_add_7_25_groupi_n_3754);
  or csa_tree_add_7_25_groupi_g17004(csa_tree_add_7_25_groupi_n_4091 ,csa_tree_add_7_25_groupi_n_3015 ,csa_tree_add_7_25_groupi_n_3568);
  or csa_tree_add_7_25_groupi_g17005(csa_tree_add_7_25_groupi_n_4090 ,csa_tree_add_7_25_groupi_n_2996 ,csa_tree_add_7_25_groupi_n_3613);
  or csa_tree_add_7_25_groupi_g17006(csa_tree_add_7_25_groupi_n_4089 ,csa_tree_add_7_25_groupi_n_2930 ,csa_tree_add_7_25_groupi_n_3634);
  or csa_tree_add_7_25_groupi_g17007(csa_tree_add_7_25_groupi_n_4088 ,csa_tree_add_7_25_groupi_n_2955 ,csa_tree_add_7_25_groupi_n_3595);
  or csa_tree_add_7_25_groupi_g17008(csa_tree_add_7_25_groupi_n_4087 ,csa_tree_add_7_25_groupi_n_3094 ,csa_tree_add_7_25_groupi_n_3688);
  or csa_tree_add_7_25_groupi_g17009(csa_tree_add_7_25_groupi_n_4086 ,csa_tree_add_7_25_groupi_n_3258 ,csa_tree_add_7_25_groupi_n_3746);
  or csa_tree_add_7_25_groupi_g17010(csa_tree_add_7_25_groupi_n_4085 ,csa_tree_add_7_25_groupi_n_3001 ,csa_tree_add_7_25_groupi_n_3614);
  or csa_tree_add_7_25_groupi_g17011(csa_tree_add_7_25_groupi_n_4084 ,csa_tree_add_7_25_groupi_n_2913 ,csa_tree_add_7_25_groupi_n_3644);
  or csa_tree_add_7_25_groupi_g17012(csa_tree_add_7_25_groupi_n_4083 ,csa_tree_add_7_25_groupi_n_2952 ,csa_tree_add_7_25_groupi_n_3606);
  or csa_tree_add_7_25_groupi_g17013(csa_tree_add_7_25_groupi_n_4082 ,csa_tree_add_7_25_groupi_n_2920 ,csa_tree_add_7_25_groupi_n_3609);
  or csa_tree_add_7_25_groupi_g17014(csa_tree_add_7_25_groupi_n_4081 ,csa_tree_add_7_25_groupi_n_3013 ,csa_tree_add_7_25_groupi_n_3624);
  or csa_tree_add_7_25_groupi_g17015(csa_tree_add_7_25_groupi_n_4080 ,csa_tree_add_7_25_groupi_n_2979 ,csa_tree_add_7_25_groupi_n_3553);
  or csa_tree_add_7_25_groupi_g17016(csa_tree_add_7_25_groupi_n_4079 ,csa_tree_add_7_25_groupi_n_3029 ,csa_tree_add_7_25_groupi_n_3600);
  or csa_tree_add_7_25_groupi_g17017(csa_tree_add_7_25_groupi_n_4078 ,csa_tree_add_7_25_groupi_n_3006 ,csa_tree_add_7_25_groupi_n_3554);
  or csa_tree_add_7_25_groupi_g17018(csa_tree_add_7_25_groupi_n_4077 ,csa_tree_add_7_25_groupi_n_2922 ,csa_tree_add_7_25_groupi_n_3626);
  or csa_tree_add_7_25_groupi_g17019(csa_tree_add_7_25_groupi_n_4076 ,csa_tree_add_7_25_groupi_n_3072 ,csa_tree_add_7_25_groupi_n_3654);
  or csa_tree_add_7_25_groupi_g17020(csa_tree_add_7_25_groupi_n_4075 ,csa_tree_add_7_25_groupi_n_2944 ,csa_tree_add_7_25_groupi_n_3678);
  or csa_tree_add_7_25_groupi_g17021(csa_tree_add_7_25_groupi_n_4074 ,csa_tree_add_7_25_groupi_n_3052 ,csa_tree_add_7_25_groupi_n_3587);
  or csa_tree_add_7_25_groupi_g17022(csa_tree_add_7_25_groupi_n_4073 ,csa_tree_add_7_25_groupi_n_3027 ,csa_tree_add_7_25_groupi_n_3619);
  or csa_tree_add_7_25_groupi_g17023(csa_tree_add_7_25_groupi_n_4072 ,csa_tree_add_7_25_groupi_n_2915 ,csa_tree_add_7_25_groupi_n_3677);
  or csa_tree_add_7_25_groupi_g17024(csa_tree_add_7_25_groupi_n_4071 ,csa_tree_add_7_25_groupi_n_3380 ,csa_tree_add_7_25_groupi_n_3779);
  or csa_tree_add_7_25_groupi_g17025(csa_tree_add_7_25_groupi_n_4070 ,csa_tree_add_7_25_groupi_n_3016 ,csa_tree_add_7_25_groupi_n_3547);
  or csa_tree_add_7_25_groupi_g17026(csa_tree_add_7_25_groupi_n_4069 ,csa_tree_add_7_25_groupi_n_3007 ,csa_tree_add_7_25_groupi_n_3579);
  or csa_tree_add_7_25_groupi_g17027(csa_tree_add_7_25_groupi_n_4068 ,csa_tree_add_7_25_groupi_n_2973 ,csa_tree_add_7_25_groupi_n_3741);
  or csa_tree_add_7_25_groupi_g17028(csa_tree_add_7_25_groupi_n_4067 ,csa_tree_add_7_25_groupi_n_2958 ,csa_tree_add_7_25_groupi_n_3615);
  or csa_tree_add_7_25_groupi_g17029(csa_tree_add_7_25_groupi_n_4066 ,csa_tree_add_7_25_groupi_n_3037 ,csa_tree_add_7_25_groupi_n_3567);
  or csa_tree_add_7_25_groupi_g17030(csa_tree_add_7_25_groupi_n_4065 ,csa_tree_add_7_25_groupi_n_3076 ,csa_tree_add_7_25_groupi_n_3656);
  or csa_tree_add_7_25_groupi_g17031(csa_tree_add_7_25_groupi_n_4064 ,csa_tree_add_7_25_groupi_n_3164 ,csa_tree_add_7_25_groupi_n_3696);
  or csa_tree_add_7_25_groupi_g17032(csa_tree_add_7_25_groupi_n_4063 ,csa_tree_add_7_25_groupi_n_3196 ,csa_tree_add_7_25_groupi_n_3705);
  or csa_tree_add_7_25_groupi_g17033(csa_tree_add_7_25_groupi_n_4062 ,csa_tree_add_7_25_groupi_n_3049 ,csa_tree_add_7_25_groupi_n_3649);
  or csa_tree_add_7_25_groupi_g17034(csa_tree_add_7_25_groupi_n_4061 ,csa_tree_add_7_25_groupi_n_3084 ,csa_tree_add_7_25_groupi_n_3665);
  or csa_tree_add_7_25_groupi_g17035(csa_tree_add_7_25_groupi_n_4060 ,csa_tree_add_7_25_groupi_n_3092 ,csa_tree_add_7_25_groupi_n_3687);
  or csa_tree_add_7_25_groupi_g17036(csa_tree_add_7_25_groupi_n_4059 ,csa_tree_add_7_25_groupi_n_3032 ,csa_tree_add_7_25_groupi_n_3552);
  or csa_tree_add_7_25_groupi_g17037(csa_tree_add_7_25_groupi_n_4058 ,csa_tree_add_7_25_groupi_n_3040 ,csa_tree_add_7_25_groupi_n_3616);
  or csa_tree_add_7_25_groupi_g17038(csa_tree_add_7_25_groupi_n_4057 ,csa_tree_add_7_25_groupi_n_2918 ,csa_tree_add_7_25_groupi_n_3549);
  or csa_tree_add_7_25_groupi_g17039(csa_tree_add_7_25_groupi_n_4056 ,csa_tree_add_7_25_groupi_n_2956 ,csa_tree_add_7_25_groupi_n_3601);
  or csa_tree_add_7_25_groupi_g17040(csa_tree_add_7_25_groupi_n_4055 ,csa_tree_add_7_25_groupi_n_2970 ,csa_tree_add_7_25_groupi_n_3675);
  or csa_tree_add_7_25_groupi_g17041(csa_tree_add_7_25_groupi_n_4054 ,csa_tree_add_7_25_groupi_n_3238 ,csa_tree_add_7_25_groupi_n_3559);
  or csa_tree_add_7_25_groupi_g17042(csa_tree_add_7_25_groupi_n_4053 ,csa_tree_add_7_25_groupi_n_3082 ,csa_tree_add_7_25_groupi_n_3674);
  or csa_tree_add_7_25_groupi_g17043(csa_tree_add_7_25_groupi_n_4052 ,csa_tree_add_7_25_groupi_n_2962 ,csa_tree_add_7_25_groupi_n_3621);
  or csa_tree_add_7_25_groupi_g17044(csa_tree_add_7_25_groupi_n_4051 ,csa_tree_add_7_25_groupi_n_3011 ,csa_tree_add_7_25_groupi_n_3625);
  or csa_tree_add_7_25_groupi_g17045(csa_tree_add_7_25_groupi_n_4050 ,csa_tree_add_7_25_groupi_n_3221 ,csa_tree_add_7_25_groupi_n_3738);
  or csa_tree_add_7_25_groupi_g17046(csa_tree_add_7_25_groupi_n_4049 ,csa_tree_add_7_25_groupi_n_3050 ,csa_tree_add_7_25_groupi_n_3640);
  or csa_tree_add_7_25_groupi_g17047(csa_tree_add_7_25_groupi_n_4048 ,csa_tree_add_7_25_groupi_n_2971 ,csa_tree_add_7_25_groupi_n_3617);
  or csa_tree_add_7_25_groupi_g17048(csa_tree_add_7_25_groupi_n_4047 ,csa_tree_add_7_25_groupi_n_3031 ,csa_tree_add_7_25_groupi_n_3593);
  or csa_tree_add_7_25_groupi_g17049(csa_tree_add_7_25_groupi_n_4046 ,csa_tree_add_7_25_groupi_n_3028 ,csa_tree_add_7_25_groupi_n_3591);
  or csa_tree_add_7_25_groupi_g17050(csa_tree_add_7_25_groupi_n_4045 ,csa_tree_add_7_25_groupi_n_2975 ,csa_tree_add_7_25_groupi_n_3620);
  or csa_tree_add_7_25_groupi_g17051(csa_tree_add_7_25_groupi_n_4044 ,csa_tree_add_7_25_groupi_n_2964 ,csa_tree_add_7_25_groupi_n_3623);
  or csa_tree_add_7_25_groupi_g17052(csa_tree_add_7_25_groupi_n_4043 ,csa_tree_add_7_25_groupi_n_3008 ,csa_tree_add_7_25_groupi_n_3589);
  or csa_tree_add_7_25_groupi_g17053(csa_tree_add_7_25_groupi_n_4042 ,csa_tree_add_7_25_groupi_n_2946 ,csa_tree_add_7_25_groupi_n_3597);
  or csa_tree_add_7_25_groupi_g17054(csa_tree_add_7_25_groupi_n_4041 ,csa_tree_add_7_25_groupi_n_2942 ,csa_tree_add_7_25_groupi_n_3608);
  or csa_tree_add_7_25_groupi_g17055(csa_tree_add_7_25_groupi_n_4040 ,csa_tree_add_7_25_groupi_n_3226 ,csa_tree_add_7_25_groupi_n_3739);
  or csa_tree_add_7_25_groupi_g17056(csa_tree_add_7_25_groupi_n_4039 ,csa_tree_add_7_25_groupi_n_3227 ,csa_tree_add_7_25_groupi_n_3707);
  or csa_tree_add_7_25_groupi_g17057(csa_tree_add_7_25_groupi_n_4038 ,csa_tree_add_7_25_groupi_n_2954 ,csa_tree_add_7_25_groupi_n_3605);
  or csa_tree_add_7_25_groupi_g17058(csa_tree_add_7_25_groupi_n_4037 ,csa_tree_add_7_25_groupi_n_2953 ,csa_tree_add_7_25_groupi_n_3566);
  or csa_tree_add_7_25_groupi_g17059(csa_tree_add_7_25_groupi_n_4036 ,csa_tree_add_7_25_groupi_n_3012 ,csa_tree_add_7_25_groupi_n_3578);
  or csa_tree_add_7_25_groupi_g17060(csa_tree_add_7_25_groupi_n_4035 ,csa_tree_add_7_25_groupi_n_3408 ,csa_tree_add_7_25_groupi_n_3766);
  or csa_tree_add_7_25_groupi_g17061(csa_tree_add_7_25_groupi_n_4034 ,csa_tree_add_7_25_groupi_n_3198 ,csa_tree_add_7_25_groupi_n_3561);
  or csa_tree_add_7_25_groupi_g17062(csa_tree_add_7_25_groupi_n_4033 ,csa_tree_add_7_25_groupi_n_3458 ,csa_tree_add_7_25_groupi_n_3803);
  or csa_tree_add_7_25_groupi_g17063(csa_tree_add_7_25_groupi_n_4032 ,csa_tree_add_7_25_groupi_n_3462 ,csa_tree_add_7_25_groupi_n_3802);
  or csa_tree_add_7_25_groupi_g17064(csa_tree_add_7_25_groupi_n_4031 ,csa_tree_add_7_25_groupi_n_3142 ,csa_tree_add_7_25_groupi_n_3731);
  or csa_tree_add_7_25_groupi_g17065(csa_tree_add_7_25_groupi_n_4030 ,csa_tree_add_7_25_groupi_n_2932 ,csa_tree_add_7_25_groupi_n_3598);
  or csa_tree_add_7_25_groupi_g17066(csa_tree_add_7_25_groupi_n_4029 ,csa_tree_add_7_25_groupi_n_3014 ,csa_tree_add_7_25_groupi_n_3576);
  or csa_tree_add_7_25_groupi_g17067(csa_tree_add_7_25_groupi_n_4028 ,csa_tree_add_7_25_groupi_n_2966 ,csa_tree_add_7_25_groupi_n_3618);
  nor csa_tree_add_7_25_groupi_g17068(csa_tree_add_7_25_groupi_n_4027 ,csa_tree_add_7_25_groupi_n_2899 ,csa_tree_add_7_25_groupi_n_3915);
  or csa_tree_add_7_25_groupi_g17069(csa_tree_add_7_25_groupi_n_4101 ,csa_tree_add_7_25_groupi_n_2380 ,csa_tree_add_7_25_groupi_n_3743);
  and csa_tree_add_7_25_groupi_g17070(csa_tree_add_7_25_groupi_n_4100 ,csa_tree_add_7_25_groupi_n_2912 ,csa_tree_add_7_25_groupi_n_3879);
  or csa_tree_add_7_25_groupi_g17071(csa_tree_add_7_25_groupi_n_4026 ,csa_tree_add_7_25_groupi_n_2928 ,csa_tree_add_7_25_groupi_n_3557);
  or csa_tree_add_7_25_groupi_g17072(csa_tree_add_7_25_groupi_n_4025 ,csa_tree_add_7_25_groupi_n_3469 ,csa_tree_add_7_25_groupi_n_3797);
  or csa_tree_add_7_25_groupi_g17073(csa_tree_add_7_25_groupi_n_4024 ,csa_tree_add_7_25_groupi_n_3045 ,csa_tree_add_7_25_groupi_n_3652);
  or csa_tree_add_7_25_groupi_g17074(csa_tree_add_7_25_groupi_n_4023 ,csa_tree_add_7_25_groupi_n_3010 ,csa_tree_add_7_25_groupi_n_3627);
  or csa_tree_add_7_25_groupi_g17075(csa_tree_add_7_25_groupi_n_4022 ,csa_tree_add_7_25_groupi_n_2984 ,csa_tree_add_7_25_groupi_n_3641);
  or csa_tree_add_7_25_groupi_g17076(csa_tree_add_7_25_groupi_n_4021 ,csa_tree_add_7_25_groupi_n_3309 ,csa_tree_add_7_25_groupi_n_3761);
  nor csa_tree_add_7_25_groupi_g17077(csa_tree_add_7_25_groupi_n_4020 ,csa_tree_add_7_25_groupi_n_292 ,csa_tree_add_7_25_groupi_n_2076);
  or csa_tree_add_7_25_groupi_g17078(csa_tree_add_7_25_groupi_n_4019 ,csa_tree_add_7_25_groupi_n_2972 ,csa_tree_add_7_25_groupi_n_3573);
  or csa_tree_add_7_25_groupi_g17079(csa_tree_add_7_25_groupi_n_4018 ,csa_tree_add_7_25_groupi_n_3019 ,csa_tree_add_7_25_groupi_n_3590);
  or csa_tree_add_7_25_groupi_g17080(csa_tree_add_7_25_groupi_n_4017 ,csa_tree_add_7_25_groupi_n_3079 ,csa_tree_add_7_25_groupi_n_3667);
  or csa_tree_add_7_25_groupi_g17081(csa_tree_add_7_25_groupi_n_4016 ,csa_tree_add_7_25_groupi_n_3452 ,csa_tree_add_7_25_groupi_n_3788);
  or csa_tree_add_7_25_groupi_g17082(csa_tree_add_7_25_groupi_n_4015 ,csa_tree_add_7_25_groupi_n_3222 ,csa_tree_add_7_25_groupi_n_3715);
  or csa_tree_add_7_25_groupi_g17083(csa_tree_add_7_25_groupi_n_4014 ,csa_tree_add_7_25_groupi_n_2997 ,csa_tree_add_7_25_groupi_n_3631);
  or csa_tree_add_7_25_groupi_g17084(csa_tree_add_7_25_groupi_n_4013 ,csa_tree_add_7_25_groupi_n_3065 ,csa_tree_add_7_25_groupi_n_3658);
  or csa_tree_add_7_25_groupi_g17085(csa_tree_add_7_25_groupi_n_4012 ,csa_tree_add_7_25_groupi_n_3331 ,csa_tree_add_7_25_groupi_n_3763);
  or csa_tree_add_7_25_groupi_g17086(csa_tree_add_7_25_groupi_n_4011 ,csa_tree_add_7_25_groupi_n_3416 ,csa_tree_add_7_25_groupi_n_3787);
  or csa_tree_add_7_25_groupi_g17087(csa_tree_add_7_25_groupi_n_4010 ,csa_tree_add_7_25_groupi_n_3193 ,csa_tree_add_7_25_groupi_n_3702);
  or csa_tree_add_7_25_groupi_g17088(csa_tree_add_7_25_groupi_n_4009 ,csa_tree_add_7_25_groupi_n_3303 ,csa_tree_add_7_25_groupi_n_3756);
  or csa_tree_add_7_25_groupi_g17089(csa_tree_add_7_25_groupi_n_4008 ,csa_tree_add_7_25_groupi_n_3403 ,csa_tree_add_7_25_groupi_n_3782);
  or csa_tree_add_7_25_groupi_g17090(csa_tree_add_7_25_groupi_n_4007 ,csa_tree_add_7_25_groupi_n_2960 ,csa_tree_add_7_25_groupi_n_3580);
  or csa_tree_add_7_25_groupi_g17091(csa_tree_add_7_25_groupi_n_4006 ,csa_tree_add_7_25_groupi_n_3047 ,csa_tree_add_7_25_groupi_n_3563);
  or csa_tree_add_7_25_groupi_g17092(csa_tree_add_7_25_groupi_n_4005 ,csa_tree_add_7_25_groupi_n_3022 ,csa_tree_add_7_25_groupi_n_3582);
  or csa_tree_add_7_25_groupi_g17093(csa_tree_add_7_25_groupi_n_4004 ,csa_tree_add_7_25_groupi_n_2982 ,csa_tree_add_7_25_groupi_n_3666);
  or csa_tree_add_7_25_groupi_g17094(csa_tree_add_7_25_groupi_n_4003 ,csa_tree_add_7_25_groupi_n_3280 ,csa_tree_add_7_25_groupi_n_3749);
  or csa_tree_add_7_25_groupi_g17095(csa_tree_add_7_25_groupi_n_4002 ,csa_tree_add_7_25_groupi_n_3383 ,csa_tree_add_7_25_groupi_n_3776);
  or csa_tree_add_7_25_groupi_g17096(csa_tree_add_7_25_groupi_n_4001 ,csa_tree_add_7_25_groupi_n_2470 ,csa_tree_add_7_25_groupi_n_3950);
  or csa_tree_add_7_25_groupi_g17097(csa_tree_add_7_25_groupi_n_4000 ,csa_tree_add_7_25_groupi_n_3163 ,csa_tree_add_7_25_groupi_n_3694);
  or csa_tree_add_7_25_groupi_g17098(csa_tree_add_7_25_groupi_n_3999 ,csa_tree_add_7_25_groupi_n_3459 ,csa_tree_add_7_25_groupi_n_3801);
  or csa_tree_add_7_25_groupi_g17099(csa_tree_add_7_25_groupi_n_3998 ,csa_tree_add_7_25_groupi_n_3088 ,csa_tree_add_7_25_groupi_n_3681);
  or csa_tree_add_7_25_groupi_g17100(csa_tree_add_7_25_groupi_n_3997 ,csa_tree_add_7_25_groupi_n_3004 ,csa_tree_add_7_25_groupi_n_3604);
  or csa_tree_add_7_25_groupi_g17101(csa_tree_add_7_25_groupi_n_3996 ,csa_tree_add_7_25_groupi_n_3291 ,csa_tree_add_7_25_groupi_n_3556);
  or csa_tree_add_7_25_groupi_g17102(csa_tree_add_7_25_groupi_n_3995 ,csa_tree_add_7_25_groupi_n_3023 ,csa_tree_add_7_25_groupi_n_3585);
  or csa_tree_add_7_25_groupi_g17103(csa_tree_add_7_25_groupi_n_3994 ,csa_tree_add_7_25_groupi_n_3352 ,csa_tree_add_7_25_groupi_n_3773);
  or csa_tree_add_7_25_groupi_g17104(csa_tree_add_7_25_groupi_n_3993 ,csa_tree_add_7_25_groupi_n_3461 ,csa_tree_add_7_25_groupi_n_3800);
  or csa_tree_add_7_25_groupi_g17105(csa_tree_add_7_25_groupi_n_3992 ,csa_tree_add_7_25_groupi_n_2933 ,csa_tree_add_7_25_groupi_n_3612);
  or csa_tree_add_7_25_groupi_g17106(csa_tree_add_7_25_groupi_n_3991 ,csa_tree_add_7_25_groupi_n_3327 ,csa_tree_add_7_25_groupi_n_3764);
  or csa_tree_add_7_25_groupi_g17107(csa_tree_add_7_25_groupi_n_3990 ,csa_tree_add_7_25_groupi_n_2917 ,csa_tree_add_7_25_groupi_n_3546);
  or csa_tree_add_7_25_groupi_g17108(csa_tree_add_7_25_groupi_n_3989 ,csa_tree_add_7_25_groupi_n_2939 ,csa_tree_add_7_25_groupi_n_3650);
  or csa_tree_add_7_25_groupi_g17109(csa_tree_add_7_25_groupi_n_3988 ,csa_tree_add_7_25_groupi_n_2948 ,csa_tree_add_7_25_groupi_n_3551);
  or csa_tree_add_7_25_groupi_g17110(csa_tree_add_7_25_groupi_n_3987 ,csa_tree_add_7_25_groupi_n_2965 ,csa_tree_add_7_25_groupi_n_3550);
  or csa_tree_add_7_25_groupi_g17111(csa_tree_add_7_25_groupi_n_3986 ,csa_tree_add_7_25_groupi_n_2929 ,csa_tree_add_7_25_groupi_n_3574);
  nor csa_tree_add_7_25_groupi_g17112(csa_tree_add_7_25_groupi_n_3985 ,csa_tree_add_7_25_groupi_n_2082 ,csa_tree_add_7_25_groupi_n_143);
  or csa_tree_add_7_25_groupi_g17113(csa_tree_add_7_25_groupi_n_3984 ,csa_tree_add_7_25_groupi_n_3002 ,csa_tree_add_7_25_groupi_n_3664);
  or csa_tree_add_7_25_groupi_g17114(csa_tree_add_7_25_groupi_n_3983 ,csa_tree_add_7_25_groupi_n_2989 ,csa_tree_add_7_25_groupi_n_3558);
  or csa_tree_add_7_25_groupi_g17115(csa_tree_add_7_25_groupi_n_3982 ,csa_tree_add_7_25_groupi_n_3081 ,csa_tree_add_7_25_groupi_n_3663);
  or csa_tree_add_7_25_groupi_g17116(csa_tree_add_7_25_groupi_n_3981 ,csa_tree_add_7_25_groupi_n_3056 ,csa_tree_add_7_25_groupi_n_3657);
  or csa_tree_add_7_25_groupi_g17117(csa_tree_add_7_25_groupi_n_3980 ,csa_tree_add_7_25_groupi_n_2986 ,csa_tree_add_7_25_groupi_n_3676);
  nor csa_tree_add_7_25_groupi_g17118(csa_tree_add_7_25_groupi_n_3979 ,csa_tree_add_7_25_groupi_n_2079 ,csa_tree_add_7_25_groupi_n_1868);
  nor csa_tree_add_7_25_groupi_g17119(csa_tree_add_7_25_groupi_n_3978 ,csa_tree_add_7_25_groupi_n_2088 ,csa_tree_add_7_25_groupi_n_1867);
  nor csa_tree_add_7_25_groupi_g17120(csa_tree_add_7_25_groupi_n_3977 ,csa_tree_add_7_25_groupi_n_318 ,csa_tree_add_7_25_groupi_n_2064);
  nor csa_tree_add_7_25_groupi_g17121(csa_tree_add_7_25_groupi_n_3976 ,csa_tree_add_7_25_groupi_n_318 ,csa_tree_add_7_25_groupi_n_2037);
  nor csa_tree_add_7_25_groupi_g17122(csa_tree_add_7_25_groupi_n_3975 ,csa_tree_add_7_25_groupi_n_317 ,csa_tree_add_7_25_groupi_n_2018);
  nor csa_tree_add_7_25_groupi_g17123(csa_tree_add_7_25_groupi_n_3974 ,csa_tree_add_7_25_groupi_n_291 ,csa_tree_add_7_25_groupi_n_1310);
  or csa_tree_add_7_25_groupi_g17124(csa_tree_add_7_25_groupi_n_3973 ,csa_tree_add_7_25_groupi_n_3720 ,csa_tree_add_7_25_groupi_n_3714);
  or csa_tree_add_7_25_groupi_g17125(csa_tree_add_7_25_groupi_n_3972 ,csa_tree_add_7_25_groupi_n_3721 ,csa_tree_add_7_25_groupi_n_3733);
  or csa_tree_add_7_25_groupi_g17126(csa_tree_add_7_25_groupi_n_3971 ,csa_tree_add_7_25_groupi_n_3724 ,csa_tree_add_7_25_groupi_n_3732);
  or csa_tree_add_7_25_groupi_g17127(csa_tree_add_7_25_groupi_n_3970 ,csa_tree_add_7_25_groupi_n_3711 ,csa_tree_add_7_25_groupi_n_3712);
  or csa_tree_add_7_25_groupi_g17128(csa_tree_add_7_25_groupi_n_3969 ,csa_tree_add_7_25_groupi_n_3723 ,csa_tree_add_7_25_groupi_n_3717);
  or csa_tree_add_7_25_groupi_g17129(csa_tree_add_7_25_groupi_n_3968 ,csa_tree_add_7_25_groupi_n_3708 ,csa_tree_add_7_25_groupi_n_3730);
  or csa_tree_add_7_25_groupi_g17130(csa_tree_add_7_25_groupi_n_3967 ,csa_tree_add_7_25_groupi_n_3728 ,csa_tree_add_7_25_groupi_n_3718);
  or csa_tree_add_7_25_groupi_g17131(csa_tree_add_7_25_groupi_n_3966 ,csa_tree_add_7_25_groupi_n_3734 ,csa_tree_add_7_25_groupi_n_3727);
  nor csa_tree_add_7_25_groupi_g17132(csa_tree_add_7_25_groupi_n_3965 ,csa_tree_add_7_25_groupi_n_3060 ,csa_tree_add_7_25_groupi_n_3545);
  or csa_tree_add_7_25_groupi_g17133(csa_tree_add_7_25_groupi_n_3964 ,csa_tree_add_7_25_groupi_n_3070 ,csa_tree_add_7_25_groupi_n_3736);
  nor csa_tree_add_7_25_groupi_g17134(csa_tree_add_7_25_groupi_n_3963 ,csa_tree_add_7_25_groupi_n_2085 ,csa_tree_add_7_25_groupi_n_143);
  or csa_tree_add_7_25_groupi_g17135(csa_tree_add_7_25_groupi_n_3962 ,csa_tree_add_7_25_groupi_n_2963 ,csa_tree_add_7_25_groupi_n_3709);
  nor csa_tree_add_7_25_groupi_g17136(csa_tree_add_7_25_groupi_n_3961 ,csa_tree_add_7_25_groupi_n_635 ,csa_tree_add_7_25_groupi_n_292);
  nor csa_tree_add_7_25_groupi_g17137(csa_tree_add_7_25_groupi_n_3960 ,csa_tree_add_7_25_groupi_n_1868 ,csa_tree_add_7_25_groupi_n_1321);
  nor csa_tree_add_7_25_groupi_g17138(csa_tree_add_7_25_groupi_n_3959 ,csa_tree_add_7_25_groupi_n_2901 ,csa_tree_add_7_25_groupi_n_3860);
  nor csa_tree_add_7_25_groupi_g17139(csa_tree_add_7_25_groupi_n_3958 ,csa_tree_add_7_25_groupi_n_3271 ,csa_tree_add_7_25_groupi_n_3729);
  nor csa_tree_add_7_25_groupi_g17140(csa_tree_add_7_25_groupi_n_3957 ,csa_tree_add_7_25_groupi_n_3357 ,csa_tree_add_7_25_groupi_n_3713);
  nor csa_tree_add_7_25_groupi_g17141(csa_tree_add_7_25_groupi_n_3956 ,csa_tree_add_7_25_groupi_n_3358 ,csa_tree_add_7_25_groupi_n_3710);
  or csa_tree_add_7_25_groupi_g17142(csa_tree_add_7_25_groupi_n_3955 ,csa_tree_add_7_25_groupi_n_3201 ,csa_tree_add_7_25_groupi_n_3719);
  nor csa_tree_add_7_25_groupi_g17143(csa_tree_add_7_25_groupi_n_3954 ,csa_tree_add_7_25_groupi_n_3204 ,csa_tree_add_7_25_groupi_n_3726);
  nor csa_tree_add_7_25_groupi_g17144(csa_tree_add_7_25_groupi_n_3953 ,csa_tree_add_7_25_groupi_n_3230 ,csa_tree_add_7_25_groupi_n_3706);
  nor csa_tree_add_7_25_groupi_g17145(csa_tree_add_7_25_groupi_n_3952 ,csa_tree_add_7_25_groupi_n_2904 ,csa_tree_add_7_25_groupi_n_3862);
  or csa_tree_add_7_25_groupi_g17146(csa_tree_add_7_25_groupi_n_3951 ,csa_tree_add_7_25_groupi_n_3064 ,csa_tree_add_7_25_groupi_n_3722);
  or csa_tree_add_7_25_groupi_g17147(csa_tree_add_7_25_groupi_n_3949 ,csa_tree_add_7_25_groupi_n_3005 ,csa_tree_add_7_25_groupi_n_3173);
  or csa_tree_add_7_25_groupi_g17148(csa_tree_add_7_25_groupi_n_3948 ,csa_tree_add_7_25_groupi_n_3044 ,csa_tree_add_7_25_groupi_n_3359);
  or csa_tree_add_7_25_groupi_g17149(csa_tree_add_7_25_groupi_n_3947 ,csa_tree_add_7_25_groupi_n_3017 ,csa_tree_add_7_25_groupi_n_3287);
  or csa_tree_add_7_25_groupi_g17150(csa_tree_add_7_25_groupi_n_3946 ,csa_tree_add_7_25_groupi_n_2977 ,csa_tree_add_7_25_groupi_n_3209);
  or csa_tree_add_7_25_groupi_g17151(csa_tree_add_7_25_groupi_n_3945 ,csa_tree_add_7_25_groupi_n_3329 ,csa_tree_add_7_25_groupi_n_3409);
  or csa_tree_add_7_25_groupi_g17152(csa_tree_add_7_25_groupi_n_3944 ,csa_tree_add_7_25_groupi_n_3020 ,csa_tree_add_7_25_groupi_n_3241);
  or csa_tree_add_7_25_groupi_g17153(csa_tree_add_7_25_groupi_n_3943 ,csa_tree_add_7_25_groupi_n_3071 ,csa_tree_add_7_25_groupi_n_3121);
  or csa_tree_add_7_25_groupi_g17154(csa_tree_add_7_25_groupi_n_3942 ,csa_tree_add_7_25_groupi_n_3350 ,csa_tree_add_7_25_groupi_n_3425);
  or csa_tree_add_7_25_groupi_g17155(csa_tree_add_7_25_groupi_n_3941 ,csa_tree_add_7_25_groupi_n_2943 ,csa_tree_add_7_25_groupi_n_3293);
  or csa_tree_add_7_25_groupi_g17156(csa_tree_add_7_25_groupi_n_3940 ,csa_tree_add_7_25_groupi_n_3426 ,csa_tree_add_7_25_groupi_n_3454);
  or csa_tree_add_7_25_groupi_g17157(csa_tree_add_7_25_groupi_n_3939 ,csa_tree_add_7_25_groupi_n_3225 ,csa_tree_add_7_25_groupi_n_3356);
  or csa_tree_add_7_25_groupi_g17158(csa_tree_add_7_25_groupi_n_3938 ,csa_tree_add_7_25_groupi_n_2940 ,csa_tree_add_7_25_groupi_n_3239);
  or csa_tree_add_7_25_groupi_g17159(csa_tree_add_7_25_groupi_n_3937 ,csa_tree_add_7_25_groupi_n_2921 ,csa_tree_add_7_25_groupi_n_3302);
  or csa_tree_add_7_25_groupi_g17160(csa_tree_add_7_25_groupi_n_3936 ,csa_tree_add_7_25_groupi_n_3308 ,csa_tree_add_7_25_groupi_n_3394);
  and csa_tree_add_7_25_groupi_g17161(csa_tree_add_7_25_groupi_n_3935 ,csa_tree_add_7_25_groupi_n_2831 ,csa_tree_add_7_25_groupi_n_3366);
  or csa_tree_add_7_25_groupi_g17162(csa_tree_add_7_25_groupi_n_3934 ,csa_tree_add_7_25_groupi_n_3096 ,csa_tree_add_7_25_groupi_n_3270);
  and csa_tree_add_7_25_groupi_g17163(csa_tree_add_7_25_groupi_n_3933 ,csa_tree_add_7_25_groupi_n_2723 ,csa_tree_add_7_25_groupi_n_3372);
  or csa_tree_add_7_25_groupi_g17164(csa_tree_add_7_25_groupi_n_3932 ,csa_tree_add_7_25_groupi_n_2923 ,csa_tree_add_7_25_groupi_n_3235);
  or csa_tree_add_7_25_groupi_g17165(csa_tree_add_7_25_groupi_n_3931 ,csa_tree_add_7_25_groupi_n_2924 ,csa_tree_add_7_25_groupi_n_3213);
  or csa_tree_add_7_25_groupi_g17166(csa_tree_add_7_25_groupi_n_3930 ,csa_tree_add_7_25_groupi_n_3378 ,csa_tree_add_7_25_groupi_n_3437);
  and csa_tree_add_7_25_groupi_g17167(csa_tree_add_7_25_groupi_n_3929 ,csa_tree_add_7_25_groupi_n_2726 ,csa_tree_add_7_25_groupi_n_3367);
  or csa_tree_add_7_25_groupi_g17168(csa_tree_add_7_25_groupi_n_3928 ,csa_tree_add_7_25_groupi_n_2951 ,csa_tree_add_7_25_groupi_n_3286);
  and csa_tree_add_7_25_groupi_g17169(csa_tree_add_7_25_groupi_n_3927 ,csa_tree_add_7_25_groupi_n_2735 ,csa_tree_add_7_25_groupi_n_3364);
  or csa_tree_add_7_25_groupi_g17170(csa_tree_add_7_25_groupi_n_3926 ,csa_tree_add_7_25_groupi_n_3228 ,csa_tree_add_7_25_groupi_n_3390);
  or csa_tree_add_7_25_groupi_g17171(csa_tree_add_7_25_groupi_n_3925 ,csa_tree_add_7_25_groupi_n_3003 ,csa_tree_add_7_25_groupi_n_3236);
  or csa_tree_add_7_25_groupi_g17172(csa_tree_add_7_25_groupi_n_3924 ,csa_tree_add_7_25_groupi_n_3351 ,csa_tree_add_7_25_groupi_n_3422);
  and csa_tree_add_7_25_groupi_g17173(csa_tree_add_7_25_groupi_n_3923 ,csa_tree_add_7_25_groupi_n_2720 ,csa_tree_add_7_25_groupi_n_3362);
  or csa_tree_add_7_25_groupi_g17174(csa_tree_add_7_25_groupi_n_3922 ,csa_tree_add_7_25_groupi_n_3400 ,csa_tree_add_7_25_groupi_n_3440);
  or csa_tree_add_7_25_groupi_g17175(csa_tree_add_7_25_groupi_n_3921 ,csa_tree_add_7_25_groupi_n_2737 ,csa_tree_add_7_25_groupi_n_3397);
  or csa_tree_add_7_25_groupi_g17176(csa_tree_add_7_25_groupi_n_3920 ,csa_tree_add_7_25_groupi_n_3063 ,csa_tree_add_7_25_groupi_n_3098);
  or csa_tree_add_7_25_groupi_g17177(csa_tree_add_7_25_groupi_n_3919 ,csa_tree_add_7_25_groupi_n_3085 ,csa_tree_add_7_25_groupi_n_3297);
  or csa_tree_add_7_25_groupi_g17178(csa_tree_add_7_25_groupi_n_3918 ,csa_tree_add_7_25_groupi_n_3087 ,csa_tree_add_7_25_groupi_n_3335);
  and csa_tree_add_7_25_groupi_g17179(csa_tree_add_7_25_groupi_n_3917 ,csa_tree_add_7_25_groupi_n_2729 ,csa_tree_add_7_25_groupi_n_3361);
  or csa_tree_add_7_25_groupi_g17180(csa_tree_add_7_25_groupi_n_3916 ,csa_tree_add_7_25_groupi_n_3443 ,csa_tree_add_7_25_groupi_n_3495);
  or csa_tree_add_7_25_groupi_g17181(csa_tree_add_7_25_groupi_n_3915 ,csa_tree_add_7_25_groupi_n_3188 ,csa_tree_add_7_25_groupi_n_3273);
  or csa_tree_add_7_25_groupi_g17182(csa_tree_add_7_25_groupi_n_3914 ,csa_tree_add_7_25_groupi_n_3353 ,csa_tree_add_7_25_groupi_n_3424);
  or csa_tree_add_7_25_groupi_g17183(csa_tree_add_7_25_groupi_n_3913 ,csa_tree_add_7_25_groupi_n_3257 ,csa_tree_add_7_25_groupi_n_3343);
  or csa_tree_add_7_25_groupi_g17184(csa_tree_add_7_25_groupi_n_3912 ,csa_tree_add_7_25_groupi_n_3305 ,csa_tree_add_7_25_groupi_n_3398);
  or csa_tree_add_7_25_groupi_g17185(csa_tree_add_7_25_groupi_n_3911 ,csa_tree_add_7_25_groupi_n_3347 ,csa_tree_add_7_25_groupi_n_3420);
  or csa_tree_add_7_25_groupi_g17186(csa_tree_add_7_25_groupi_n_3910 ,csa_tree_add_7_25_groupi_n_3021 ,csa_tree_add_7_25_groupi_n_3244);
  or csa_tree_add_7_25_groupi_g17187(csa_tree_add_7_25_groupi_n_3909 ,csa_tree_add_7_25_groupi_n_3307 ,csa_tree_add_7_25_groupi_n_3412);
  or csa_tree_add_7_25_groupi_g17188(csa_tree_add_7_25_groupi_n_3908 ,csa_tree_add_7_25_groupi_n_3278 ,csa_tree_add_7_25_groupi_n_3375);
  or csa_tree_add_7_25_groupi_g17189(csa_tree_add_7_25_groupi_n_3907 ,csa_tree_add_7_25_groupi_n_3261 ,csa_tree_add_7_25_groupi_n_3354);
  or csa_tree_add_7_25_groupi_g17190(csa_tree_add_7_25_groupi_n_3906 ,csa_tree_add_7_25_groupi_n_3073 ,csa_tree_add_7_25_groupi_n_3301);
  or csa_tree_add_7_25_groupi_g17191(csa_tree_add_7_25_groupi_n_3905 ,csa_tree_add_7_25_groupi_n_3430 ,csa_tree_add_7_25_groupi_n_3453);
  and csa_tree_add_7_25_groupi_g17192(csa_tree_add_7_25_groupi_n_3904 ,csa_tree_add_7_25_groupi_n_2719 ,csa_tree_add_7_25_groupi_n_3369);
  or csa_tree_add_7_25_groupi_g17193(csa_tree_add_7_25_groupi_n_3903 ,csa_tree_add_7_25_groupi_n_3306 ,csa_tree_add_7_25_groupi_n_3406);
  or csa_tree_add_7_25_groupi_g17194(csa_tree_add_7_25_groupi_n_3902 ,csa_tree_add_7_25_groupi_n_3066 ,csa_tree_add_7_25_groupi_n_3243);
  or csa_tree_add_7_25_groupi_g17195(csa_tree_add_7_25_groupi_n_3901 ,csa_tree_add_7_25_groupi_n_3068 ,csa_tree_add_7_25_groupi_n_3324);
  or csa_tree_add_7_25_groupi_g17196(csa_tree_add_7_25_groupi_n_3900 ,csa_tree_add_7_25_groupi_n_3089 ,csa_tree_add_7_25_groupi_n_3311);
  and csa_tree_add_7_25_groupi_g17197(csa_tree_add_7_25_groupi_n_3899 ,csa_tree_add_7_25_groupi_n_2728 ,csa_tree_add_7_25_groupi_n_3370);
  or csa_tree_add_7_25_groupi_g17198(csa_tree_add_7_25_groupi_n_3898 ,csa_tree_add_7_25_groupi_n_2991 ,csa_tree_add_7_25_groupi_n_3207);
  or csa_tree_add_7_25_groupi_g17199(csa_tree_add_7_25_groupi_n_3897 ,csa_tree_add_7_25_groupi_n_3419 ,csa_tree_add_7_25_groupi_n_3449);
  or csa_tree_add_7_25_groupi_g17200(csa_tree_add_7_25_groupi_n_3896 ,csa_tree_add_7_25_groupi_n_3075 ,csa_tree_add_7_25_groupi_n_3178);
  or csa_tree_add_7_25_groupi_g17201(csa_tree_add_7_25_groupi_n_3895 ,csa_tree_add_7_25_groupi_n_2992 ,csa_tree_add_7_25_groupi_n_3212);
  or csa_tree_add_7_25_groupi_g17202(csa_tree_add_7_25_groupi_n_3894 ,csa_tree_add_7_25_groupi_n_3159 ,csa_tree_add_7_25_groupi_n_3300);
  and csa_tree_add_7_25_groupi_g17203(csa_tree_add_7_25_groupi_n_3893 ,csa_tree_add_7_25_groupi_n_2722 ,csa_tree_add_7_25_groupi_n_3363);
  or csa_tree_add_7_25_groupi_g17204(csa_tree_add_7_25_groupi_n_3892 ,csa_tree_add_7_25_groupi_n_3279 ,csa_tree_add_7_25_groupi_n_3391);
  or csa_tree_add_7_25_groupi_g17205(csa_tree_add_7_25_groupi_n_3891 ,csa_tree_add_7_25_groupi_n_3077 ,csa_tree_add_7_25_groupi_n_3254);
  or csa_tree_add_7_25_groupi_g17206(csa_tree_add_7_25_groupi_n_3890 ,csa_tree_add_7_25_groupi_n_3061 ,csa_tree_add_7_25_groupi_n_3145);
  or csa_tree_add_7_25_groupi_g17207(csa_tree_add_7_25_groupi_n_3889 ,csa_tree_add_7_25_groupi_n_3428 ,csa_tree_add_7_25_groupi_n_3457);
  or csa_tree_add_7_25_groupi_g17208(csa_tree_add_7_25_groupi_n_3888 ,csa_tree_add_7_25_groupi_n_3069 ,csa_tree_add_7_25_groupi_n_3250);
  or csa_tree_add_7_25_groupi_g17209(csa_tree_add_7_25_groupi_n_3887 ,csa_tree_add_7_25_groupi_n_2967 ,csa_tree_add_7_25_groupi_n_3170);
  or csa_tree_add_7_25_groupi_g17210(csa_tree_add_7_25_groupi_n_3886 ,csa_tree_add_7_25_groupi_n_2961 ,csa_tree_add_7_25_groupi_n_3290);
  or csa_tree_add_7_25_groupi_g17211(csa_tree_add_7_25_groupi_n_3885 ,csa_tree_add_7_25_groupi_n_2998 ,csa_tree_add_7_25_groupi_n_3289);
  or csa_tree_add_7_25_groupi_g17212(csa_tree_add_7_25_groupi_n_3884 ,csa_tree_add_7_25_groupi_n_3046 ,csa_tree_add_7_25_groupi_n_3203);
  or csa_tree_add_7_25_groupi_g17213(csa_tree_add_7_25_groupi_n_3883 ,csa_tree_add_7_25_groupi_n_3161 ,csa_tree_add_7_25_groupi_n_3295);
  or csa_tree_add_7_25_groupi_g17214(csa_tree_add_7_25_groupi_n_3882 ,csa_tree_add_7_25_groupi_n_3192 ,csa_tree_add_7_25_groupi_n_3314);
  or csa_tree_add_7_25_groupi_g17215(csa_tree_add_7_25_groupi_n_3881 ,csa_tree_add_7_25_groupi_n_3274 ,csa_tree_add_7_25_groupi_n_3377);
  or csa_tree_add_7_25_groupi_g17216(csa_tree_add_7_25_groupi_n_3880 ,csa_tree_add_7_25_groupi_n_3304 ,csa_tree_add_7_25_groupi_n_3393);
  and csa_tree_add_7_25_groupi_g17217(csa_tree_add_7_25_groupi_n_3879 ,csa_tree_add_7_25_groupi_n_3396 ,csa_tree_add_7_25_groupi_n_3386);
  or csa_tree_add_7_25_groupi_g17218(csa_tree_add_7_25_groupi_n_3878 ,csa_tree_add_7_25_groupi_n_3414 ,csa_tree_add_7_25_groupi_n_3448);
  or csa_tree_add_7_25_groupi_g17219(csa_tree_add_7_25_groupi_n_3877 ,csa_tree_add_7_25_groupi_n_3431 ,csa_tree_add_7_25_groupi_n_3456);
  or csa_tree_add_7_25_groupi_g17220(csa_tree_add_7_25_groupi_n_3876 ,csa_tree_add_7_25_groupi_n_2945 ,csa_tree_add_7_25_groupi_n_3172);
  or csa_tree_add_7_25_groupi_g17221(csa_tree_add_7_25_groupi_n_3875 ,csa_tree_add_7_25_groupi_n_3223 ,csa_tree_add_7_25_groupi_n_3341);
  or csa_tree_add_7_25_groupi_g17222(csa_tree_add_7_25_groupi_n_3874 ,csa_tree_add_7_25_groupi_n_3080 ,csa_tree_add_7_25_groupi_n_3267);
  or csa_tree_add_7_25_groupi_g17223(csa_tree_add_7_25_groupi_n_3873 ,csa_tree_add_7_25_groupi_n_3349 ,csa_tree_add_7_25_groupi_n_3421);
  or csa_tree_add_7_25_groupi_g17224(csa_tree_add_7_25_groupi_n_3872 ,csa_tree_add_7_25_groupi_n_3445 ,csa_tree_add_7_25_groupi_n_3470);
  or csa_tree_add_7_25_groupi_g17225(csa_tree_add_7_25_groupi_n_3871 ,csa_tree_add_7_25_groupi_n_3090 ,csa_tree_add_7_25_groupi_n_3266);
  or csa_tree_add_7_25_groupi_g17226(csa_tree_add_7_25_groupi_n_3870 ,csa_tree_add_7_25_groupi_n_2926 ,csa_tree_add_7_25_groupi_n_3205);
  and csa_tree_add_7_25_groupi_g17227(csa_tree_add_7_25_groupi_n_3869 ,csa_tree_add_7_25_groupi_n_2724 ,csa_tree_add_7_25_groupi_n_3368);
  or csa_tree_add_7_25_groupi_g17228(csa_tree_add_7_25_groupi_n_3868 ,csa_tree_add_7_25_groupi_n_3185 ,csa_tree_add_7_25_groupi_n_3323);
  or csa_tree_add_7_25_groupi_g17229(csa_tree_add_7_25_groupi_n_3867 ,csa_tree_add_7_25_groupi_n_2935 ,csa_tree_add_7_25_groupi_n_3216);
  or csa_tree_add_7_25_groupi_g17230(csa_tree_add_7_25_groupi_n_3866 ,csa_tree_add_7_25_groupi_n_3197 ,csa_tree_add_7_25_groupi_n_3321);
  or csa_tree_add_7_25_groupi_g17231(csa_tree_add_7_25_groupi_n_3865 ,csa_tree_add_7_25_groupi_n_3379 ,csa_tree_add_7_25_groupi_n_3436);
  or csa_tree_add_7_25_groupi_g17232(csa_tree_add_7_25_groupi_n_3864 ,csa_tree_add_7_25_groupi_n_3091 ,csa_tree_add_7_25_groupi_n_3355);
  or csa_tree_add_7_25_groupi_g17233(csa_tree_add_7_25_groupi_n_3863 ,csa_tree_add_7_25_groupi_n_3277 ,csa_tree_add_7_25_groupi_n_3374);
  or csa_tree_add_7_25_groupi_g17234(csa_tree_add_7_25_groupi_n_3862 ,csa_tree_add_7_25_groupi_n_3186 ,csa_tree_add_7_25_groupi_n_3317);
  or csa_tree_add_7_25_groupi_g17235(csa_tree_add_7_25_groupi_n_3861 ,csa_tree_add_7_25_groupi_n_3441 ,csa_tree_add_7_25_groupi_n_3482);
  or csa_tree_add_7_25_groupi_g17236(csa_tree_add_7_25_groupi_n_3860 ,csa_tree_add_7_25_groupi_n_3498 ,csa_tree_add_7_25_groupi_n_3252);
  or csa_tree_add_7_25_groupi_g17237(csa_tree_add_7_25_groupi_n_3859 ,csa_tree_add_7_25_groupi_n_3053 ,csa_tree_add_7_25_groupi_n_3316);
  or csa_tree_add_7_25_groupi_g17238(csa_tree_add_7_25_groupi_n_3858 ,csa_tree_add_7_25_groupi_n_3275 ,csa_tree_add_7_25_groupi_n_3399);
  or csa_tree_add_7_25_groupi_g17239(csa_tree_add_7_25_groupi_n_3857 ,csa_tree_add_7_25_groupi_n_2916 ,csa_tree_add_7_25_groupi_n_3175);
  or csa_tree_add_7_25_groupi_g17240(csa_tree_add_7_25_groupi_n_3856 ,csa_tree_add_7_25_groupi_n_3162 ,csa_tree_add_7_25_groupi_n_3312);
  or csa_tree_add_7_25_groupi_g17241(csa_tree_add_7_25_groupi_n_3855 ,csa_tree_add_7_25_groupi_n_2938 ,csa_tree_add_7_25_groupi_n_3211);
  or csa_tree_add_7_25_groupi_g17242(csa_tree_add_7_25_groupi_n_3854 ,csa_tree_add_7_25_groupi_n_3054 ,csa_tree_add_7_25_groupi_n_3272);
  or csa_tree_add_7_25_groupi_g17243(csa_tree_add_7_25_groupi_n_3853 ,csa_tree_add_7_25_groupi_n_3059 ,csa_tree_add_7_25_groupi_n_3234);
  or csa_tree_add_7_25_groupi_g17244(csa_tree_add_7_25_groupi_n_3852 ,csa_tree_add_7_25_groupi_n_3158 ,csa_tree_add_7_25_groupi_n_3342);
  or csa_tree_add_7_25_groupi_g17245(csa_tree_add_7_25_groupi_n_3851 ,csa_tree_add_7_25_groupi_n_2994 ,csa_tree_add_7_25_groupi_n_3202);
  or csa_tree_add_7_25_groupi_g17246(csa_tree_add_7_25_groupi_n_3850 ,csa_tree_add_7_25_groupi_n_3402 ,csa_tree_add_7_25_groupi_n_3447);
  or csa_tree_add_7_25_groupi_g17247(csa_tree_add_7_25_groupi_n_3849 ,csa_tree_add_7_25_groupi_n_3067 ,csa_tree_add_7_25_groupi_n_3129);
  or csa_tree_add_7_25_groupi_g17248(csa_tree_add_7_25_groupi_n_3848 ,csa_tree_add_7_25_groupi_n_2949 ,csa_tree_add_7_25_groupi_n_3208);
  nor csa_tree_add_7_25_groupi_g17249(csa_tree_add_7_25_groupi_n_3847 ,csa_tree_add_7_25_groupi_n_764 ,csa_tree_add_7_25_groupi_n_1418);
  or csa_tree_add_7_25_groupi_g17250(csa_tree_add_7_25_groupi_n_3846 ,csa_tree_add_7_25_groupi_n_3051 ,csa_tree_add_7_25_groupi_n_3231);
  or csa_tree_add_7_25_groupi_g17251(csa_tree_add_7_25_groupi_n_3845 ,csa_tree_add_7_25_groupi_n_3026 ,csa_tree_add_7_25_groupi_n_3288);
  or csa_tree_add_7_25_groupi_g17252(csa_tree_add_7_25_groupi_n_3844 ,csa_tree_add_7_25_groupi_n_3190 ,csa_tree_add_7_25_groupi_n_3340);
  or csa_tree_add_7_25_groupi_g17253(csa_tree_add_7_25_groupi_n_3843 ,csa_tree_add_7_25_groupi_n_2914 ,csa_tree_add_7_25_groupi_n_3284);
  or csa_tree_add_7_25_groupi_g17254(csa_tree_add_7_25_groupi_n_3842 ,csa_tree_add_7_25_groupi_n_3259 ,csa_tree_add_7_25_groupi_n_3360);
  or csa_tree_add_7_25_groupi_g17255(csa_tree_add_7_25_groupi_n_3841 ,csa_tree_add_7_25_groupi_n_3083 ,csa_tree_add_7_25_groupi_n_3339);
  or csa_tree_add_7_25_groupi_g17256(csa_tree_add_7_25_groupi_n_3840 ,csa_tree_add_7_25_groupi_n_3157 ,csa_tree_add_7_25_groupi_n_3322);
  or csa_tree_add_7_25_groupi_g17257(csa_tree_add_7_25_groupi_n_3839 ,csa_tree_add_7_25_groupi_n_3000 ,csa_tree_add_7_25_groupi_n_3283);
  or csa_tree_add_7_25_groupi_g17258(csa_tree_add_7_25_groupi_n_3838 ,csa_tree_add_7_25_groupi_n_3058 ,csa_tree_add_7_25_groupi_n_3210);
  and csa_tree_add_7_25_groupi_g17259(csa_tree_add_7_25_groupi_n_3837 ,csa_tree_add_7_25_groupi_n_2718 ,csa_tree_add_7_25_groupi_n_3365);
  or csa_tree_add_7_25_groupi_g17260(csa_tree_add_7_25_groupi_n_3836 ,csa_tree_add_7_25_groupi_n_3062 ,csa_tree_add_7_25_groupi_n_3292);
  or csa_tree_add_7_25_groupi_g17261(csa_tree_add_7_25_groupi_n_3835 ,csa_tree_add_7_25_groupi_n_3042 ,csa_tree_add_7_25_groupi_n_3181);
  or csa_tree_add_7_25_groupi_g17262(csa_tree_add_7_25_groupi_n_3834 ,csa_tree_add_7_25_groupi_n_2988 ,csa_tree_add_7_25_groupi_n_3246);
  or csa_tree_add_7_25_groupi_g17263(csa_tree_add_7_25_groupi_n_3833 ,csa_tree_add_7_25_groupi_n_2957 ,csa_tree_add_7_25_groupi_n_3240);
  or csa_tree_add_7_25_groupi_g17264(csa_tree_add_7_25_groupi_n_3832 ,csa_tree_add_7_25_groupi_n_3427 ,csa_tree_add_7_25_groupi_n_3455);
  and csa_tree_add_7_25_groupi_g17265(csa_tree_add_7_25_groupi_n_3831 ,csa_tree_add_7_25_groupi_n_2725 ,csa_tree_add_7_25_groupi_n_2925);
  or csa_tree_add_7_25_groupi_g17266(csa_tree_add_7_25_groupi_n_3830 ,csa_tree_add_7_25_groupi_n_2987 ,csa_tree_add_7_25_groupi_n_3285);
  or csa_tree_add_7_25_groupi_g17267(csa_tree_add_7_25_groupi_n_3829 ,csa_tree_add_7_25_groupi_n_3086 ,csa_tree_add_7_25_groupi_n_3320);
  or csa_tree_add_7_25_groupi_g17268(csa_tree_add_7_25_groupi_n_3828 ,csa_tree_add_7_25_groupi_n_2931 ,csa_tree_add_7_25_groupi_n_3182);
  or csa_tree_add_7_25_groupi_g17269(csa_tree_add_7_25_groupi_n_3827 ,csa_tree_add_7_25_groupi_n_3018 ,csa_tree_add_7_25_groupi_n_3282);
  or csa_tree_add_7_25_groupi_g17270(csa_tree_add_7_25_groupi_n_3826 ,csa_tree_add_7_25_groupi_n_2981 ,csa_tree_add_7_25_groupi_n_3233);
  or csa_tree_add_7_25_groupi_g17271(csa_tree_add_7_25_groupi_n_3825 ,csa_tree_add_7_25_groupi_n_3328 ,csa_tree_add_7_25_groupi_n_3411);
  or csa_tree_add_7_25_groupi_g17272(csa_tree_add_7_25_groupi_n_3824 ,csa_tree_add_7_25_groupi_n_3382 ,csa_tree_add_7_25_groupi_n_3434);
  or csa_tree_add_7_25_groupi_g17273(csa_tree_add_7_25_groupi_n_3823 ,csa_tree_add_7_25_groupi_n_3224 ,csa_tree_add_7_25_groupi_n_3334);
  or csa_tree_add_7_25_groupi_g17274(csa_tree_add_7_25_groupi_n_3822 ,csa_tree_add_7_25_groupi_n_2959 ,csa_tree_add_7_25_groupi_n_3149);
  or csa_tree_add_7_25_groupi_g17275(csa_tree_add_7_25_groupi_n_3821 ,csa_tree_add_7_25_groupi_n_2999 ,csa_tree_add_7_25_groupi_n_3263);
  or csa_tree_add_7_25_groupi_g17276(csa_tree_add_7_25_groupi_n_3820 ,csa_tree_add_7_25_groupi_n_3255 ,csa_tree_add_7_25_groupi_n_3388);
  or csa_tree_add_7_25_groupi_g17277(csa_tree_add_7_25_groupi_n_3819 ,csa_tree_add_7_25_groupi_n_3384 ,csa_tree_add_7_25_groupi_n_3433);
  or csa_tree_add_7_25_groupi_g17278(csa_tree_add_7_25_groupi_n_3818 ,csa_tree_add_7_25_groupi_n_3418 ,csa_tree_add_7_25_groupi_n_3450);
  or csa_tree_add_7_25_groupi_g17279(csa_tree_add_7_25_groupi_n_3817 ,csa_tree_add_7_25_groupi_n_3262 ,csa_tree_add_7_25_groupi_n_3345);
  or csa_tree_add_7_25_groupi_g17280(csa_tree_add_7_25_groupi_n_3816 ,csa_tree_add_7_25_groupi_n_3401 ,csa_tree_add_7_25_groupi_n_3438);
  or csa_tree_add_7_25_groupi_g17281(csa_tree_add_7_25_groupi_n_3815 ,csa_tree_add_7_25_groupi_n_3404 ,csa_tree_add_7_25_groupi_n_3439);
  or csa_tree_add_7_25_groupi_g17282(csa_tree_add_7_25_groupi_n_3814 ,csa_tree_add_7_25_groupi_n_3326 ,csa_tree_add_7_25_groupi_n_3413);
  and csa_tree_add_7_25_groupi_g17283(csa_tree_add_7_25_groupi_n_3813 ,csa_tree_add_7_25_groupi_n_2727 ,csa_tree_add_7_25_groupi_n_3389);
  or csa_tree_add_7_25_groupi_g17284(csa_tree_add_7_25_groupi_n_3812 ,csa_tree_add_7_25_groupi_n_2976 ,csa_tree_add_7_25_groupi_n_3206);
  or csa_tree_add_7_25_groupi_g17285(csa_tree_add_7_25_groupi_n_3811 ,csa_tree_add_7_25_groupi_n_2937 ,csa_tree_add_7_25_groupi_n_3237);
  or csa_tree_add_7_25_groupi_g17286(csa_tree_add_7_25_groupi_n_3810 ,csa_tree_add_7_25_groupi_n_3034 ,csa_tree_add_7_25_groupi_n_3242);
  or csa_tree_add_7_25_groupi_g17287(csa_tree_add_7_25_groupi_n_3809 ,csa_tree_add_7_25_groupi_n_3039 ,csa_tree_add_7_25_groupi_n_3214);
  or csa_tree_add_7_25_groupi_g17288(csa_tree_add_7_25_groupi_n_3808 ,csa_tree_add_7_25_groupi_n_2993 ,csa_tree_add_7_25_groupi_n_3171);
  nor csa_tree_add_7_25_groupi_g17289(csa_tree_add_7_25_groupi_n_3807 ,csa_tree_add_7_25_groupi_n_641 ,csa_tree_add_7_25_groupi_n_1538);
  nor csa_tree_add_7_25_groupi_g17290(csa_tree_add_7_25_groupi_n_3806 ,csa_tree_add_7_25_groupi_n_951 ,csa_tree_add_7_25_groupi_n_1466);
  nor csa_tree_add_7_25_groupi_g17291(csa_tree_add_7_25_groupi_n_3805 ,csa_tree_add_7_25_groupi_n_644 ,csa_tree_add_7_25_groupi_n_1715);
  nor csa_tree_add_7_25_groupi_g17292(csa_tree_add_7_25_groupi_n_3804 ,csa_tree_add_7_25_groupi_n_624 ,csa_tree_add_7_25_groupi_n_1388);
  nor csa_tree_add_7_25_groupi_g17293(csa_tree_add_7_25_groupi_n_3803 ,csa_tree_add_7_25_groupi_n_626 ,csa_tree_add_7_25_groupi_n_1496);
  nor csa_tree_add_7_25_groupi_g17294(csa_tree_add_7_25_groupi_n_3802 ,csa_tree_add_7_25_groupi_n_626 ,csa_tree_add_7_25_groupi_n_1565);
  nor csa_tree_add_7_25_groupi_g17295(csa_tree_add_7_25_groupi_n_3801 ,csa_tree_add_7_25_groupi_n_994 ,csa_tree_add_7_25_groupi_n_1421);
  nor csa_tree_add_7_25_groupi_g17296(csa_tree_add_7_25_groupi_n_3800 ,csa_tree_add_7_25_groupi_n_999 ,csa_tree_add_7_25_groupi_n_1514);
  nor csa_tree_add_7_25_groupi_g17297(csa_tree_add_7_25_groupi_n_3799 ,csa_tree_add_7_25_groupi_n_767 ,csa_tree_add_7_25_groupi_n_1544);
  nor csa_tree_add_7_25_groupi_g17298(csa_tree_add_7_25_groupi_n_3798 ,csa_tree_add_7_25_groupi_n_64 ,csa_tree_add_7_25_groupi_n_1480);
  nor csa_tree_add_7_25_groupi_g17299(csa_tree_add_7_25_groupi_n_3797 ,csa_tree_add_7_25_groupi_n_1003 ,csa_tree_add_7_25_groupi_n_1385);
  nor csa_tree_add_7_25_groupi_g17300(csa_tree_add_7_25_groupi_n_3796 ,csa_tree_add_7_25_groupi_n_114 ,csa_tree_add_7_25_groupi_n_1679);
  nor csa_tree_add_7_25_groupi_g17301(csa_tree_add_7_25_groupi_n_3795 ,csa_tree_add_7_25_groupi_n_996 ,csa_tree_add_7_25_groupi_n_1516);
  nor csa_tree_add_7_25_groupi_g17302(csa_tree_add_7_25_groupi_n_3794 ,csa_tree_add_7_25_groupi_n_463 ,csa_tree_add_7_25_groupi_n_1504);
  nor csa_tree_add_7_25_groupi_g17303(csa_tree_add_7_25_groupi_n_3793 ,csa_tree_add_7_25_groupi_n_481 ,csa_tree_add_7_25_groupi_n_1540);
  nor csa_tree_add_7_25_groupi_g17304(csa_tree_add_7_25_groupi_n_3792 ,csa_tree_add_7_25_groupi_n_1881 ,csa_tree_add_7_25_groupi_n_1409);
  nor csa_tree_add_7_25_groupi_g17305(csa_tree_add_7_25_groupi_n_3791 ,csa_tree_add_7_25_groupi_n_1883 ,csa_tree_add_7_25_groupi_n_1483);
  nor csa_tree_add_7_25_groupi_g17306(csa_tree_add_7_25_groupi_n_3790 ,csa_tree_add_7_25_groupi_n_1887 ,csa_tree_add_7_25_groupi_n_1471);
  nor csa_tree_add_7_25_groupi_g17307(csa_tree_add_7_25_groupi_n_3789 ,csa_tree_add_7_25_groupi_n_477 ,csa_tree_add_7_25_groupi_n_1528);
  nor csa_tree_add_7_25_groupi_g17308(csa_tree_add_7_25_groupi_n_3788 ,csa_tree_add_7_25_groupi_n_468 ,csa_tree_add_7_25_groupi_n_1408);
  nor csa_tree_add_7_25_groupi_g17309(csa_tree_add_7_25_groupi_n_3787 ,csa_tree_add_7_25_groupi_n_466 ,csa_tree_add_7_25_groupi_n_1453);
  nor csa_tree_add_7_25_groupi_g17310(csa_tree_add_7_25_groupi_n_3786 ,csa_tree_add_7_25_groupi_n_478 ,csa_tree_add_7_25_groupi_n_1546);
  nor csa_tree_add_7_25_groupi_g17311(csa_tree_add_7_25_groupi_n_3785 ,csa_tree_add_7_25_groupi_n_469 ,csa_tree_add_7_25_groupi_n_1468);
  nor csa_tree_add_7_25_groupi_g17312(csa_tree_add_7_25_groupi_n_3784 ,csa_tree_add_7_25_groupi_n_442 ,csa_tree_add_7_25_groupi_n_1493);
  nor csa_tree_add_7_25_groupi_g17313(csa_tree_add_7_25_groupi_n_3783 ,csa_tree_add_7_25_groupi_n_486 ,csa_tree_add_7_25_groupi_n_1382);
  nor csa_tree_add_7_25_groupi_g17314(csa_tree_add_7_25_groupi_n_3782 ,csa_tree_add_7_25_groupi_n_442 ,csa_tree_add_7_25_groupi_n_1459);
  nor csa_tree_add_7_25_groupi_g17315(csa_tree_add_7_25_groupi_n_3781 ,csa_tree_add_7_25_groupi_n_445 ,csa_tree_add_7_25_groupi_n_1477);
  nor csa_tree_add_7_25_groupi_g17316(csa_tree_add_7_25_groupi_n_3780 ,csa_tree_add_7_25_groupi_n_486 ,csa_tree_add_7_25_groupi_n_2009);
  nor csa_tree_add_7_25_groupi_g17317(csa_tree_add_7_25_groupi_n_3779 ,csa_tree_add_7_25_groupi_n_454 ,csa_tree_add_7_25_groupi_n_1504);
  nor csa_tree_add_7_25_groupi_g17318(csa_tree_add_7_25_groupi_n_3778 ,csa_tree_add_7_25_groupi_n_451 ,csa_tree_add_7_25_groupi_n_2010);
  nor csa_tree_add_7_25_groupi_g17319(csa_tree_add_7_25_groupi_n_3777 ,csa_tree_add_7_25_groupi_n_460 ,csa_tree_add_7_25_groupi_n_1540);
  nor csa_tree_add_7_25_groupi_g17320(csa_tree_add_7_25_groupi_n_3776 ,csa_tree_add_7_25_groupi_n_298 ,csa_tree_add_7_25_groupi_n_1457);
  nor csa_tree_add_7_25_groupi_g17321(csa_tree_add_7_25_groupi_n_3775 ,csa_tree_add_7_25_groupi_n_457 ,csa_tree_add_7_25_groupi_n_1567);
  nor csa_tree_add_7_25_groupi_g17322(csa_tree_add_7_25_groupi_n_3774 ,csa_tree_add_7_25_groupi_n_454 ,csa_tree_add_7_25_groupi_n_1475);
  nor csa_tree_add_7_25_groupi_g17323(csa_tree_add_7_25_groupi_n_3773 ,csa_tree_add_7_25_groupi_n_439 ,csa_tree_add_7_25_groupi_n_1453);
  nor csa_tree_add_7_25_groupi_g17324(csa_tree_add_7_25_groupi_n_3772 ,csa_tree_add_7_25_groupi_n_409 ,csa_tree_add_7_25_groupi_n_1409);
  nor csa_tree_add_7_25_groupi_g17325(csa_tree_add_7_25_groupi_n_3771 ,csa_tree_add_7_25_groupi_n_348 ,csa_tree_add_7_25_groupi_n_1468);
  nor csa_tree_add_7_25_groupi_g17326(csa_tree_add_7_25_groupi_n_3770 ,csa_tree_add_7_25_groupi_n_424 ,csa_tree_add_7_25_groupi_n_1556);
  nor csa_tree_add_7_25_groupi_g17327(csa_tree_add_7_25_groupi_n_3769 ,csa_tree_add_7_25_groupi_n_391 ,csa_tree_add_7_25_groupi_n_1382);
  nor csa_tree_add_7_25_groupi_g17328(csa_tree_add_7_25_groupi_n_3768 ,csa_tree_add_7_25_groupi_n_397 ,csa_tree_add_7_25_groupi_n_1493);
  nor csa_tree_add_7_25_groupi_g17329(csa_tree_add_7_25_groupi_n_3767 ,csa_tree_add_7_25_groupi_n_370 ,csa_tree_add_7_25_groupi_n_1528);
  nor csa_tree_add_7_25_groupi_g17330(csa_tree_add_7_25_groupi_n_3766 ,csa_tree_add_7_25_groupi_n_368 ,csa_tree_add_7_25_groupi_n_1475);
  nor csa_tree_add_7_25_groupi_g17331(csa_tree_add_7_25_groupi_n_3765 ,csa_tree_add_7_25_groupi_n_382 ,csa_tree_add_7_25_groupi_n_1787);
  nor csa_tree_add_7_25_groupi_g17332(csa_tree_add_7_25_groupi_n_3764 ,csa_tree_add_7_25_groupi_n_377 ,csa_tree_add_7_25_groupi_n_1457);
  nor csa_tree_add_7_25_groupi_g17333(csa_tree_add_7_25_groupi_n_3763 ,csa_tree_add_7_25_groupi_n_371 ,csa_tree_add_7_25_groupi_n_1546);
  nor csa_tree_add_7_25_groupi_g17334(csa_tree_add_7_25_groupi_n_3762 ,csa_tree_add_7_25_groupi_n_540 ,csa_tree_add_7_25_groupi_n_1559);
  nor csa_tree_add_7_25_groupi_g17335(csa_tree_add_7_25_groupi_n_3761 ,csa_tree_add_7_25_groupi_n_557 ,csa_tree_add_7_25_groupi_n_1459);
  nor csa_tree_add_7_25_groupi_g17336(csa_tree_add_7_25_groupi_n_3760 ,csa_tree_add_7_25_groupi_n_385 ,csa_tree_add_7_25_groupi_n_1733);
  nor csa_tree_add_7_25_groupi_g17337(csa_tree_add_7_25_groupi_n_3759 ,csa_tree_add_7_25_groupi_n_430 ,csa_tree_add_7_25_groupi_n_1567);
  nor csa_tree_add_7_25_groupi_g17338(csa_tree_add_7_25_groupi_n_3758 ,csa_tree_add_7_25_groupi_n_412 ,csa_tree_add_7_25_groupi_n_1477);
  nor csa_tree_add_7_25_groupi_g17339(csa_tree_add_7_25_groupi_n_3757 ,csa_tree_add_7_25_groupi_n_558 ,csa_tree_add_7_25_groupi_n_1516);
  nor csa_tree_add_7_25_groupi_g17340(csa_tree_add_7_25_groupi_n_3756 ,csa_tree_add_7_25_groupi_n_561 ,csa_tree_add_7_25_groupi_n_1480);
  nor csa_tree_add_7_25_groupi_g17341(csa_tree_add_7_25_groupi_n_3755 ,csa_tree_add_7_25_groupi_n_415 ,csa_tree_add_7_25_groupi_n_2006);
  nor csa_tree_add_7_25_groupi_g17342(csa_tree_add_7_25_groupi_n_3754 ,csa_tree_add_7_25_groupi_n_418 ,csa_tree_add_7_25_groupi_n_1483);
  nor csa_tree_add_7_25_groupi_g17343(csa_tree_add_7_25_groupi_n_3753 ,csa_tree_add_7_25_groupi_n_762 ,csa_tree_add_7_25_groupi_n_1471);
  nor csa_tree_add_7_25_groupi_g17344(csa_tree_add_7_25_groupi_n_3752 ,csa_tree_add_7_25_groupi_n_564 ,csa_tree_add_7_25_groupi_n_1529);
  nor csa_tree_add_7_25_groupi_g17345(csa_tree_add_7_25_groupi_n_3751 ,csa_tree_add_7_25_groupi_n_567 ,csa_tree_add_7_25_groupi_n_1571);
  nor csa_tree_add_7_25_groupi_g17346(csa_tree_add_7_25_groupi_n_3750 ,csa_tree_add_7_25_groupi_n_400 ,csa_tree_add_7_25_groupi_n_1342);
  nor csa_tree_add_7_25_groupi_g17347(csa_tree_add_7_25_groupi_n_3749 ,csa_tree_add_7_25_groupi_n_354 ,csa_tree_add_7_25_groupi_n_1547);
  nor csa_tree_add_7_25_groupi_g17348(csa_tree_add_7_25_groupi_n_3748 ,csa_tree_add_7_25_groupi_n_344 ,csa_tree_add_7_25_groupi_n_1726);
  nor csa_tree_add_7_25_groupi_g17349(csa_tree_add_7_25_groupi_n_3747 ,csa_tree_add_7_25_groupi_n_765 ,csa_tree_add_7_25_groupi_n_1783);
  nor csa_tree_add_7_25_groupi_g17350(csa_tree_add_7_25_groupi_n_3746 ,csa_tree_add_7_25_groupi_n_768 ,csa_tree_add_7_25_groupi_n_1460);
  nor csa_tree_add_7_25_groupi_g17351(csa_tree_add_7_25_groupi_n_3745 ,csa_tree_add_7_25_groupi_n_570 ,csa_tree_add_7_25_groupi_n_1744);
  or csa_tree_add_7_25_groupi_g17352(csa_tree_add_7_25_groupi_n_3744 ,csa_tree_add_7_25_groupi_n_30 ,csa_tree_add_7_25_groupi_n_2909);
  and csa_tree_add_7_25_groupi_g17353(csa_tree_add_7_25_groupi_n_3950 ,csa_tree_add_7_25_groupi_n_2456 ,csa_tree_add_7_25_groupi_n_3478);
  nor csa_tree_add_7_25_groupi_g17354(csa_tree_add_7_25_groupi_n_3741 ,csa_tree_add_7_25_groupi_n_671 ,csa_tree_add_7_25_groupi_n_1535);
  nor csa_tree_add_7_25_groupi_g17355(csa_tree_add_7_25_groupi_n_3740 ,csa_tree_add_7_25_groupi_n_573 ,csa_tree_add_7_25_groupi_n_1995);
  nor csa_tree_add_7_25_groupi_g17356(csa_tree_add_7_25_groupi_n_3739 ,csa_tree_add_7_25_groupi_n_471 ,csa_tree_add_7_25_groupi_n_2007);
  nor csa_tree_add_7_25_groupi_g17357(csa_tree_add_7_25_groupi_n_3738 ,csa_tree_add_7_25_groupi_n_773 ,csa_tree_add_7_25_groupi_n_1598);
  nor csa_tree_add_7_25_groupi_g17358(csa_tree_add_7_25_groupi_n_3737 ,csa_tree_add_7_25_groupi_n_771 ,csa_tree_add_7_25_groupi_n_1555);
  nor csa_tree_add_7_25_groupi_g17359(csa_tree_add_7_25_groupi_n_3736 ,csa_tree_add_7_25_groupi_n_285 ,csa_tree_add_7_25_groupi_n_2130);
  nor csa_tree_add_7_25_groupi_g17360(csa_tree_add_7_25_groupi_n_3735 ,csa_tree_add_7_25_groupi_n_774 ,csa_tree_add_7_25_groupi_n_1904);
  nor csa_tree_add_7_25_groupi_g17361(csa_tree_add_7_25_groupi_n_3734 ,csa_tree_add_7_25_groupi_n_582 ,csa_tree_add_7_25_groupi_n_1995);
  nor csa_tree_add_7_25_groupi_g17362(csa_tree_add_7_25_groupi_n_3733 ,csa_tree_add_7_25_groupi_n_2055 ,csa_tree_add_7_25_groupi_n_1865);
  nor csa_tree_add_7_25_groupi_g17363(csa_tree_add_7_25_groupi_n_3732 ,csa_tree_add_7_25_groupi_n_2115 ,csa_tree_add_7_25_groupi_n_1864);
  nor csa_tree_add_7_25_groupi_g17364(csa_tree_add_7_25_groupi_n_3731 ,csa_tree_add_7_25_groupi_n_585 ,csa_tree_add_7_25_groupi_n_1484);
  nor csa_tree_add_7_25_groupi_g17365(csa_tree_add_7_25_groupi_n_3730 ,csa_tree_add_7_25_groupi_n_2024 ,csa_tree_add_7_25_groupi_n_166);
  or csa_tree_add_7_25_groupi_g17366(csa_tree_add_7_25_groupi_n_3729 ,csa_tree_add_7_25_groupi_n_3195 ,csa_tree_add_7_25_groupi_n_2902);
  nor csa_tree_add_7_25_groupi_g17367(csa_tree_add_7_25_groupi_n_3728 ,csa_tree_add_7_25_groupi_n_936 ,csa_tree_add_7_25_groupi_n_1905);
  nor csa_tree_add_7_25_groupi_g17368(csa_tree_add_7_25_groupi_n_3727 ,csa_tree_add_7_25_groupi_n_312 ,csa_tree_add_7_25_groupi_n_2051);
  or csa_tree_add_7_25_groupi_g17369(csa_tree_add_7_25_groupi_n_3726 ,csa_tree_add_7_25_groupi_n_3187 ,csa_tree_add_7_25_groupi_n_2905);
  nor csa_tree_add_7_25_groupi_g17370(csa_tree_add_7_25_groupi_n_3725 ,csa_tree_add_7_25_groupi_n_780 ,csa_tree_add_7_25_groupi_n_1478);
  nor csa_tree_add_7_25_groupi_g17371(csa_tree_add_7_25_groupi_n_3724 ,csa_tree_add_7_25_groupi_n_939 ,csa_tree_add_7_25_groupi_n_1637);
  nor csa_tree_add_7_25_groupi_g17372(csa_tree_add_7_25_groupi_n_3723 ,csa_tree_add_7_25_groupi_n_543 ,csa_tree_add_7_25_groupi_n_1379);
  or csa_tree_add_7_25_groupi_g17373(csa_tree_add_7_25_groupi_n_3722 ,csa_tree_add_7_25_groupi_n_2646 ,csa_tree_add_7_25_groupi_n_2910);
  nor csa_tree_add_7_25_groupi_g17374(csa_tree_add_7_25_groupi_n_3721 ,csa_tree_add_7_25_groupi_n_546 ,csa_tree_add_7_25_groupi_n_1786);
  nor csa_tree_add_7_25_groupi_g17375(csa_tree_add_7_25_groupi_n_3720 ,csa_tree_add_7_25_groupi_n_576 ,csa_tree_add_7_25_groupi_n_1517);
  or csa_tree_add_7_25_groupi_g17376(csa_tree_add_7_25_groupi_n_3719 ,csa_tree_add_7_25_groupi_n_3385 ,csa_tree_add_7_25_groupi_n_2897);
  nor csa_tree_add_7_25_groupi_g17377(csa_tree_add_7_25_groupi_n_3718 ,csa_tree_add_7_25_groupi_n_362 ,csa_tree_add_7_25_groupi_n_286);
  nor csa_tree_add_7_25_groupi_g17378(csa_tree_add_7_25_groupi_n_3717 ,csa_tree_add_7_25_groupi_n_311 ,csa_tree_add_7_25_groupi_n_2148);
  nor csa_tree_add_7_25_groupi_g17379(csa_tree_add_7_25_groupi_n_3716 ,csa_tree_add_7_25_groupi_n_588 ,csa_tree_add_7_25_groupi_n_1733);
  nor csa_tree_add_7_25_groupi_g17380(csa_tree_add_7_25_groupi_n_3715 ,csa_tree_add_7_25_groupi_n_472 ,csa_tree_add_7_25_groupi_n_1513);
  nor csa_tree_add_7_25_groupi_g17381(csa_tree_add_7_25_groupi_n_3714 ,csa_tree_add_7_25_groupi_n_312 ,csa_tree_add_7_25_groupi_n_2094);
  or csa_tree_add_7_25_groupi_g17382(csa_tree_add_7_25_groupi_n_3713 ,csa_tree_add_7_25_groupi_n_3184 ,csa_tree_add_7_25_groupi_n_2898);
  nor csa_tree_add_7_25_groupi_g17383(csa_tree_add_7_25_groupi_n_3712 ,csa_tree_add_7_25_groupi_n_1865 ,csa_tree_add_7_25_groupi_n_1321);
  nor csa_tree_add_7_25_groupi_g17384(csa_tree_add_7_25_groupi_n_3711 ,csa_tree_add_7_25_groupi_n_579 ,csa_tree_add_7_25_groupi_n_42);
  or csa_tree_add_7_25_groupi_g17385(csa_tree_add_7_25_groupi_n_3710 ,csa_tree_add_7_25_groupi_n_3191 ,csa_tree_add_7_25_groupi_n_2900);
  nor csa_tree_add_7_25_groupi_g17386(csa_tree_add_7_25_groupi_n_3709 ,csa_tree_add_7_25_groupi_n_286 ,csa_tree_add_7_25_groupi_n_2172);
  nor csa_tree_add_7_25_groupi_g17387(csa_tree_add_7_25_groupi_n_3708 ,csa_tree_add_7_25_groupi_n_581 ,csa_tree_add_7_25_groupi_n_1744);
  nor csa_tree_add_7_25_groupi_g17388(csa_tree_add_7_25_groupi_n_3707 ,csa_tree_add_7_25_groupi_n_388 ,csa_tree_add_7_25_groupi_n_1481);
  or csa_tree_add_7_25_groupi_g17389(csa_tree_add_7_25_groupi_n_3706 ,csa_tree_add_7_25_groupi_n_3183 ,csa_tree_add_7_25_groupi_n_2903);
  nor csa_tree_add_7_25_groupi_g17390(csa_tree_add_7_25_groupi_n_3705 ,csa_tree_add_7_25_groupi_n_834 ,csa_tree_add_7_25_groupi_n_1678);
  nor csa_tree_add_7_25_groupi_g17391(csa_tree_add_7_25_groupi_n_3704 ,csa_tree_add_7_25_groupi_n_840 ,csa_tree_add_7_25_groupi_n_1543);
  nor csa_tree_add_7_25_groupi_g17392(csa_tree_add_7_25_groupi_n_3703 ,csa_tree_add_7_25_groupi_n_786 ,csa_tree_add_7_25_groupi_n_1408);
  nor csa_tree_add_7_25_groupi_g17393(csa_tree_add_7_25_groupi_n_3702 ,csa_tree_add_7_25_groupi_n_789 ,csa_tree_add_7_25_groupi_n_1534);
  nor csa_tree_add_7_25_groupi_g17394(csa_tree_add_7_25_groupi_n_3701 ,csa_tree_add_7_25_groupi_n_833 ,csa_tree_add_7_25_groupi_n_1472);
  nor csa_tree_add_7_25_groupi_g17395(csa_tree_add_7_25_groupi_n_3700 ,csa_tree_add_7_25_groupi_n_839 ,csa_tree_add_7_25_groupi_n_1994);
  nor csa_tree_add_7_25_groupi_g17396(csa_tree_add_7_25_groupi_n_3699 ,csa_tree_add_7_25_groupi_n_427 ,csa_tree_add_7_25_groupi_n_1774);
  nor csa_tree_add_7_25_groupi_g17397(csa_tree_add_7_25_groupi_n_3698 ,csa_tree_add_7_25_groupi_n_433 ,csa_tree_add_7_25_groupi_n_1295);
  nor csa_tree_add_7_25_groupi_g17398(csa_tree_add_7_25_groupi_n_3697 ,csa_tree_add_7_25_groupi_n_795 ,csa_tree_add_7_25_groupi_n_1636);
  nor csa_tree_add_7_25_groupi_g17399(csa_tree_add_7_25_groupi_n_3696 ,csa_tree_add_7_25_groupi_n_647 ,csa_tree_add_7_25_groupi_n_1597);
  nor csa_tree_add_7_25_groupi_g17400(csa_tree_add_7_25_groupi_n_3695 ,csa_tree_add_7_25_groupi_n_611 ,csa_tree_add_7_25_groupi_n_1784);
  nor csa_tree_add_7_25_groupi_g17401(csa_tree_add_7_25_groupi_n_3694 ,csa_tree_add_7_25_groupi_n_845 ,csa_tree_add_7_25_groupi_n_1513);
  nor csa_tree_add_7_25_groupi_g17402(csa_tree_add_7_25_groupi_n_3693 ,csa_tree_add_7_25_groupi_n_650 ,csa_tree_add_7_25_groupi_n_1994);
  nor csa_tree_add_7_25_groupi_g17403(csa_tree_add_7_25_groupi_n_3692 ,csa_tree_add_7_25_groupi_n_436 ,csa_tree_add_7_25_groupi_n_1727);
  nor csa_tree_add_7_25_groupi_g17404(csa_tree_add_7_25_groupi_n_3691 ,csa_tree_add_7_25_groupi_n_594 ,csa_tree_add_7_25_groupi_n_1907);
  nor csa_tree_add_7_25_groupi_g17405(csa_tree_add_7_25_groupi_n_3690 ,csa_tree_add_7_25_groupi_n_606 ,csa_tree_add_7_25_groupi_n_1384);
  nor csa_tree_add_7_25_groupi_g17406(csa_tree_add_7_25_groupi_n_3689 ,csa_tree_add_7_25_groupi_n_669 ,csa_tree_add_7_25_groupi_n_1568);
  nor csa_tree_add_7_25_groupi_g17407(csa_tree_add_7_25_groupi_n_3688 ,csa_tree_add_7_25_groupi_n_660 ,csa_tree_add_7_25_groupi_n_1543);
  nor csa_tree_add_7_25_groupi_g17408(csa_tree_add_7_25_groupi_n_3687 ,csa_tree_add_7_25_groupi_n_656 ,csa_tree_add_7_25_groupi_n_1678);
  nor csa_tree_add_7_25_groupi_g17409(csa_tree_add_7_25_groupi_n_3686 ,csa_tree_add_7_25_groupi_n_665 ,csa_tree_add_7_25_groupi_n_1343);
  nor csa_tree_add_7_25_groupi_g17410(csa_tree_add_7_25_groupi_n_3685 ,csa_tree_add_7_25_groupi_n_851 ,csa_tree_add_7_25_groupi_n_1732);
  nor csa_tree_add_7_25_groupi_g17411(csa_tree_add_7_25_groupi_n_3684 ,csa_tree_add_7_25_groupi_n_827 ,csa_tree_add_7_25_groupi_n_1378);
  nor csa_tree_add_7_25_groupi_g17412(csa_tree_add_7_25_groupi_n_3683 ,csa_tree_add_7_25_groupi_n_659 ,csa_tree_add_7_25_groupi_n_533);
  nor csa_tree_add_7_25_groupi_g17413(csa_tree_add_7_25_groupi_n_3682 ,csa_tree_add_7_25_groupi_n_668 ,csa_tree_add_7_25_groupi_n_134);
  nor csa_tree_add_7_25_groupi_g17414(csa_tree_add_7_25_groupi_n_3681 ,csa_tree_add_7_25_groupi_n_609 ,csa_tree_add_7_25_groupi_n_1417);
  nor csa_tree_add_7_25_groupi_g17415(csa_tree_add_7_25_groupi_n_3680 ,csa_tree_add_7_25_groupi_n_618 ,csa_tree_add_7_25_groupi_n_1156);
  nor csa_tree_add_7_25_groupi_g17416(csa_tree_add_7_25_groupi_n_3679 ,csa_tree_add_7_25_groupi_n_776 ,csa_tree_add_7_25_groupi_n_198);
  nor csa_tree_add_7_25_groupi_g17417(csa_tree_add_7_25_groupi_n_3678 ,csa_tree_add_7_25_groupi_n_791 ,csa_tree_add_7_25_groupi_n_1163);
  nor csa_tree_add_7_25_groupi_g17418(csa_tree_add_7_25_groupi_n_3677 ,csa_tree_add_7_25_groupi_n_44 ,csa_tree_add_7_25_groupi_n_1714);
  nor csa_tree_add_7_25_groupi_g17419(csa_tree_add_7_25_groupi_n_3676 ,csa_tree_add_7_25_groupi_n_777 ,csa_tree_add_7_25_groupi_n_1537);
  nor csa_tree_add_7_25_groupi_g17420(csa_tree_add_7_25_groupi_n_3675 ,csa_tree_add_7_25_groupi_n_929 ,csa_tree_add_7_25_groupi_n_1384);
  nor csa_tree_add_7_25_groupi_g17421(csa_tree_add_7_25_groupi_n_3674 ,csa_tree_add_7_25_groupi_n_696 ,csa_tree_add_7_25_groupi_n_1465);
  nor csa_tree_add_7_25_groupi_g17422(csa_tree_add_7_25_groupi_n_3673 ,csa_tree_add_7_25_groupi_n_1044 ,csa_tree_add_7_25_groupi_n_534);
  nor csa_tree_add_7_25_groupi_g17423(csa_tree_add_7_25_groupi_n_3672 ,csa_tree_add_7_25_groupi_n_683 ,csa_tree_add_7_25_groupi_n_1300);
  nor csa_tree_add_7_25_groupi_g17424(csa_tree_add_7_25_groupi_n_3671 ,csa_tree_add_7_25_groupi_n_692 ,csa_tree_add_7_25_groupi_n_533);
  nor csa_tree_add_7_25_groupi_g17425(csa_tree_add_7_25_groupi_n_3670 ,csa_tree_add_7_25_groupi_n_863 ,csa_tree_add_7_25_groupi_n_1154);
  nor csa_tree_add_7_25_groupi_g17426(csa_tree_add_7_25_groupi_n_3669 ,csa_tree_add_7_25_groupi_n_1047 ,csa_tree_add_7_25_groupi_n_1772);
  nor csa_tree_add_7_25_groupi_g17427(csa_tree_add_7_25_groupi_n_3668 ,csa_tree_add_7_25_groupi_n_966 ,csa_tree_add_7_25_groupi_n_2195);
  nor csa_tree_add_7_25_groupi_g17428(csa_tree_add_7_25_groupi_n_3667 ,csa_tree_add_7_25_groupi_n_686 ,csa_tree_add_7_25_groupi_n_1387);
  nor csa_tree_add_7_25_groupi_g17429(csa_tree_add_7_25_groupi_n_3666 ,csa_tree_add_7_25_groupi_n_963 ,csa_tree_add_7_25_groupi_n_1420);
  nor csa_tree_add_7_25_groupi_g17430(csa_tree_add_7_25_groupi_n_3665 ,csa_tree_add_7_25_groupi_n_695 ,csa_tree_add_7_25_groupi_n_1564);
  nor csa_tree_add_7_25_groupi_g17431(csa_tree_add_7_25_groupi_n_3664 ,csa_tree_add_7_25_groupi_n_932 ,csa_tree_add_7_25_groupi_n_1558);
  nor csa_tree_add_7_25_groupi_g17432(csa_tree_add_7_25_groupi_n_3663 ,csa_tree_add_7_25_groupi_n_617 ,csa_tree_add_7_25_groupi_n_1535);
  nor csa_tree_add_7_25_groupi_g17433(csa_tree_add_7_25_groupi_n_3662 ,csa_tree_add_7_25_groupi_n_701 ,csa_tree_add_7_25_groupi_n_1505);
  nor csa_tree_add_7_25_groupi_g17434(csa_tree_add_7_25_groupi_n_3661 ,csa_tree_add_7_25_groupi_n_878 ,csa_tree_add_7_25_groupi_n_1151);
  nor csa_tree_add_7_25_groupi_g17435(csa_tree_add_7_25_groupi_n_3660 ,csa_tree_add_7_25_groupi_n_1035 ,csa_tree_add_7_25_groupi_n_2195);
  nor csa_tree_add_7_25_groupi_g17436(csa_tree_add_7_25_groupi_n_3659 ,csa_tree_add_7_25_groupi_n_975 ,csa_tree_add_7_25_groupi_n_1300);
  nor csa_tree_add_7_25_groupi_g17437(csa_tree_add_7_25_groupi_n_3658 ,csa_tree_add_7_25_groupi_n_620 ,csa_tree_add_7_25_groupi_n_1598);
  nor csa_tree_add_7_25_groupi_g17438(csa_tree_add_7_25_groupi_n_3657 ,csa_tree_add_7_25_groupi_n_704 ,csa_tree_add_7_25_groupi_n_1495);
  nor csa_tree_add_7_25_groupi_g17439(csa_tree_add_7_25_groupi_n_3656 ,csa_tree_add_7_25_groupi_n_756 ,csa_tree_add_7_25_groupi_n_1637);
  nor csa_tree_add_7_25_groupi_g17440(csa_tree_add_7_25_groupi_n_3655 ,csa_tree_add_7_25_groupi_n_867 ,csa_tree_add_7_25_groupi_n_941);
  nor csa_tree_add_7_25_groupi_g17441(csa_tree_add_7_25_groupi_n_3654 ,csa_tree_add_7_25_groupi_n_879 ,csa_tree_add_7_25_groupi_n_1157);
  nor csa_tree_add_7_25_groupi_g17442(csa_tree_add_7_25_groupi_n_3653 ,csa_tree_add_7_25_groupi_n_714 ,csa_tree_add_7_25_groupi_n_536);
  nor csa_tree_add_7_25_groupi_g17443(csa_tree_add_7_25_groupi_n_3652 ,csa_tree_add_7_25_groupi_n_824 ,csa_tree_add_7_25_groupi_n_1771);
  nor csa_tree_add_7_25_groupi_g17444(csa_tree_add_7_25_groupi_n_3651 ,csa_tree_add_7_25_groupi_n_698 ,csa_tree_add_7_25_groupi_n_1162);
  nor csa_tree_add_7_25_groupi_g17445(csa_tree_add_7_25_groupi_n_3650 ,csa_tree_add_7_25_groupi_n_752 ,csa_tree_add_7_25_groupi_n_1379);
  nor csa_tree_add_7_25_groupi_g17446(csa_tree_add_7_25_groupi_n_3649 ,csa_tree_add_7_25_groupi_n_818 ,csa_tree_add_7_25_groupi_n_1537);
  nor csa_tree_add_7_25_groupi_g17447(csa_tree_add_7_25_groupi_n_3648 ,csa_tree_add_7_25_groupi_n_689 ,csa_tree_add_7_25_groupi_n_1541);
  nor csa_tree_add_7_25_groupi_g17448(csa_tree_add_7_25_groupi_n_3647 ,csa_tree_add_7_25_groupi_n_860 ,csa_tree_add_7_25_groupi_n_1775);
  nor csa_tree_add_7_25_groupi_g17449(csa_tree_add_7_25_groupi_n_3646 ,csa_tree_add_7_25_groupi_n_782 ,csa_tree_add_7_25_groupi_n_1727);
  nor csa_tree_add_7_25_groupi_g17450(csa_tree_add_7_25_groupi_n_3645 ,csa_tree_add_7_25_groupi_n_725 ,csa_tree_add_7_25_groupi_n_537);
  nor csa_tree_add_7_25_groupi_g17451(csa_tree_add_7_25_groupi_n_3644 ,csa_tree_add_7_25_groupi_n_836 ,csa_tree_add_7_25_groupi_n_1469);
  nor csa_tree_add_7_25_groupi_g17452(csa_tree_add_7_25_groupi_n_3643 ,csa_tree_add_7_25_groupi_n_848 ,csa_tree_add_7_25_groupi_n_42);
  nor csa_tree_add_7_25_groupi_g17453(csa_tree_add_7_25_groupi_n_3642 ,csa_tree_add_7_25_groupi_n_54 ,csa_tree_add_7_25_groupi_n_1295);
  nor csa_tree_add_7_25_groupi_g17454(csa_tree_add_7_25_groupi_n_3641 ,csa_tree_add_7_25_groupi_n_758 ,csa_tree_add_7_25_groupi_n_1381);
  nor csa_tree_add_7_25_groupi_g17455(csa_tree_add_7_25_groupi_n_3640 ,csa_tree_add_7_25_groupi_n_825 ,csa_tree_add_7_25_groupi_n_1564);
  nor csa_tree_add_7_25_groupi_g17456(csa_tree_add_7_25_groupi_n_3639 ,csa_tree_add_7_25_groupi_n_728 ,csa_tree_add_7_25_groupi_n_1294);
  nor csa_tree_add_7_25_groupi_g17457(csa_tree_add_7_25_groupi_n_3638 ,csa_tree_add_7_25_groupi_n_82 ,csa_tree_add_7_25_groupi_n_536);
  nor csa_tree_add_7_25_groupi_g17458(csa_tree_add_7_25_groupi_n_3637 ,csa_tree_add_7_25_groupi_n_403 ,csa_tree_add_7_25_groupi_n_1495);
  nor csa_tree_add_7_25_groupi_g17459(csa_tree_add_7_25_groupi_n_3636 ,csa_tree_add_7_25_groupi_n_716 ,csa_tree_add_7_25_groupi_n_1294);
  nor csa_tree_add_7_25_groupi_g17460(csa_tree_add_7_25_groupi_n_3635 ,csa_tree_add_7_25_groupi_n_800 ,csa_tree_add_7_25_groupi_n_1154);
  nor csa_tree_add_7_25_groupi_g17461(csa_tree_add_7_25_groupi_n_3634 ,csa_tree_add_7_25_groupi_n_908 ,csa_tree_add_7_25_groupi_n_1474);
  nor csa_tree_add_7_25_groupi_g17462(csa_tree_add_7_25_groupi_n_3633 ,csa_tree_add_7_25_groupi_n_890 ,csa_tree_add_7_25_groupi_n_1150);
  nor csa_tree_add_7_25_groupi_g17463(csa_tree_add_7_25_groupi_n_3632 ,csa_tree_add_7_25_groupi_n_92 ,csa_tree_add_7_25_groupi_n_2006);
  nor csa_tree_add_7_25_groupi_g17464(csa_tree_add_7_25_groupi_n_3631 ,csa_tree_add_7_25_groupi_n_806 ,csa_tree_add_7_25_groupi_n_1517);
  nor csa_tree_add_7_25_groupi_g17465(csa_tree_add_7_25_groupi_n_3630 ,csa_tree_add_7_25_groupi_n_875 ,csa_tree_add_7_25_groupi_n_1775);
  nor csa_tree_add_7_25_groupi_g17466(csa_tree_add_7_25_groupi_n_3629 ,csa_tree_add_7_25_groupi_n_672 ,csa_tree_add_7_25_groupi_n_527);
  nor csa_tree_add_7_25_groupi_g17467(csa_tree_add_7_25_groupi_n_3628 ,csa_tree_add_7_25_groupi_n_72 ,csa_tree_add_7_25_groupi_n_528);
  nor csa_tree_add_7_25_groupi_g17468(csa_tree_add_7_25_groupi_n_3627 ,csa_tree_add_7_25_groupi_n_707 ,csa_tree_add_7_25_groupi_n_1381);
  nor csa_tree_add_7_25_groupi_g17469(csa_tree_add_7_25_groupi_n_3626 ,csa_tree_add_7_25_groupi_n_837 ,csa_tree_add_7_25_groupi_n_1529);
  nor csa_tree_add_7_25_groupi_g17470(csa_tree_add_7_25_groupi_n_3625 ,csa_tree_add_7_25_groupi_n_749 ,csa_tree_add_7_25_groupi_n_1514);
  nor csa_tree_add_7_25_groupi_g17471(csa_tree_add_7_25_groupi_n_3624 ,csa_tree_add_7_25_groupi_n_690 ,csa_tree_add_7_25_groupi_n_1786);
  nor csa_tree_add_7_25_groupi_g17472(csa_tree_add_7_25_groupi_n_3623 ,csa_tree_add_7_25_groupi_n_46 ,csa_tree_add_7_25_groupi_n_1472);
  nor csa_tree_add_7_25_groupi_g17473(csa_tree_add_7_25_groupi_n_3622 ,csa_tree_add_7_25_groupi_n_1026 ,csa_tree_add_7_25_groupi_n_1568);
  nor csa_tree_add_7_25_groupi_g17474(csa_tree_add_7_25_groupi_n_3621 ,csa_tree_add_7_25_groupi_n_86 ,csa_tree_add_7_25_groupi_n_1534);
  nor csa_tree_add_7_25_groupi_g17475(csa_tree_add_7_25_groupi_n_3620 ,csa_tree_add_7_25_groupi_n_812 ,csa_tree_add_7_25_groupi_n_1492);
  nor csa_tree_add_7_25_groupi_g17476(csa_tree_add_7_25_groupi_n_3619 ,csa_tree_add_7_25_groupi_n_753 ,csa_tree_add_7_25_groupi_n_1454);
  nor csa_tree_add_7_25_groupi_g17477(csa_tree_add_7_25_groupi_n_3618 ,csa_tree_add_7_25_groupi_n_99 ,csa_tree_add_7_25_groupi_n_1505);
  nor csa_tree_add_7_25_groupi_g17478(csa_tree_add_7_25_groupi_n_3617 ,csa_tree_add_7_25_groupi_n_84 ,csa_tree_add_7_25_groupi_n_1481);
  nor csa_tree_add_7_25_groupi_g17479(csa_tree_add_7_25_groupi_n_3616 ,csa_tree_add_7_25_groupi_n_909 ,csa_tree_add_7_25_groupi_n_2007);
  nor csa_tree_add_7_25_groupi_g17480(csa_tree_add_7_25_groupi_n_3615 ,csa_tree_add_7_25_groupi_n_797 ,csa_tree_add_7_25_groupi_n_1474);
  nor csa_tree_add_7_25_groupi_g17481(csa_tree_add_7_25_groupi_n_3614 ,csa_tree_add_7_25_groupi_n_911 ,csa_tree_add_7_25_groupi_n_2009);
  nor csa_tree_add_7_25_groupi_g17482(csa_tree_add_7_25_groupi_n_3613 ,csa_tree_add_7_25_groupi_n_917 ,csa_tree_add_7_25_groupi_n_1558);
  nor csa_tree_add_7_25_groupi_g17483(csa_tree_add_7_25_groupi_n_3612 ,csa_tree_add_7_25_groupi_n_713 ,csa_tree_add_7_25_groupi_n_1420);
  nor csa_tree_add_7_25_groupi_g17484(csa_tree_add_7_25_groupi_n_3611 ,csa_tree_add_7_25_groupi_n_869 ,csa_tree_add_7_25_groupi_n_1745);
  nor csa_tree_add_7_25_groupi_g17485(csa_tree_add_7_25_groupi_n_3610 ,csa_tree_add_7_25_groupi_n_1080 ,csa_tree_add_7_25_groupi_n_534);
  nor csa_tree_add_7_25_groupi_g17486(csa_tree_add_7_25_groupi_n_3609 ,csa_tree_add_7_25_groupi_n_849 ,csa_tree_add_7_25_groupi_n_1163);
  nor csa_tree_add_7_25_groupi_g17487(csa_tree_add_7_25_groupi_n_3608 ,csa_tree_add_7_25_groupi_n_857 ,csa_tree_add_7_25_groupi_n_1492);
  nor csa_tree_add_7_25_groupi_g17488(csa_tree_add_7_25_groupi_n_3607 ,csa_tree_add_7_25_groupi_n_746 ,csa_tree_add_7_25_groupi_n_527);
  nor csa_tree_add_7_25_groupi_g17489(csa_tree_add_7_25_groupi_n_3606 ,csa_tree_add_7_25_groupi_n_1029 ,csa_tree_add_7_25_groupi_n_1547);
  nor csa_tree_add_7_25_groupi_g17490(csa_tree_add_7_25_groupi_n_3605 ,csa_tree_add_7_25_groupi_n_719 ,csa_tree_add_7_25_groupi_n_168);
  nor csa_tree_add_7_25_groupi_g17491(csa_tree_add_7_25_groupi_n_3604 ,csa_tree_add_7_25_groupi_n_1062 ,csa_tree_add_7_25_groupi_n_1456);
  nor csa_tree_add_7_25_groupi_g17492(csa_tree_add_7_25_groupi_n_3603 ,csa_tree_add_7_25_groupi_n_1068 ,csa_tree_add_7_25_groupi_n_528);
  nor csa_tree_add_7_25_groupi_g17493(csa_tree_add_7_25_groupi_n_3602 ,csa_tree_add_7_25_groupi_n_1032 ,csa_tree_add_7_25_groupi_n_198);
  nor csa_tree_add_7_25_groupi_g17494(csa_tree_add_7_25_groupi_n_3601 ,csa_tree_add_7_25_groupi_n_902 ,csa_tree_add_7_25_groupi_n_1417);
  nor csa_tree_add_7_25_groupi_g17495(csa_tree_add_7_25_groupi_n_3600 ,csa_tree_add_7_25_groupi_n_710 ,csa_tree_add_7_25_groupi_n_1784);
  nor csa_tree_add_7_25_groupi_g17496(csa_tree_add_7_25_groupi_n_3599 ,csa_tree_add_7_25_groupi_n_78 ,csa_tree_add_7_25_groupi_n_1771);
  nor csa_tree_add_7_25_groupi_g17497(csa_tree_add_7_25_groupi_n_3598 ,csa_tree_add_7_25_groupi_n_50 ,csa_tree_add_7_25_groupi_n_1484);
  nor csa_tree_add_7_25_groupi_g17498(csa_tree_add_7_25_groupi_n_3597 ,csa_tree_add_7_25_groupi_n_1005 ,csa_tree_add_7_25_groupi_n_1456);
  nor csa_tree_add_7_25_groupi_g17499(csa_tree_add_7_25_groupi_n_3596 ,csa_tree_add_7_25_groupi_n_972 ,csa_tree_add_7_25_groupi_n_168);
  nor csa_tree_add_7_25_groupi_g17500(csa_tree_add_7_25_groupi_n_3595 ,csa_tree_add_7_25_groupi_n_801 ,csa_tree_add_7_25_groupi_n_1538);
  nor csa_tree_add_7_25_groupi_g17501(csa_tree_add_7_25_groupi_n_3594 ,csa_tree_add_7_25_groupi_n_1086 ,csa_tree_add_7_25_groupi_n_1783);
  nor csa_tree_add_7_25_groupi_g17502(csa_tree_add_7_25_groupi_n_3593 ,csa_tree_add_7_25_groupi_n_1050 ,csa_tree_add_7_25_groupi_n_1418);
  nor csa_tree_add_7_25_groupi_g17503(csa_tree_add_7_25_groupi_n_3592 ,csa_tree_add_7_25_groupi_n_920 ,csa_tree_add_7_25_groupi_n_202);
  nor csa_tree_add_7_25_groupi_g17504(csa_tree_add_7_25_groupi_n_3591 ,csa_tree_add_7_25_groupi_n_750 ,csa_tree_add_7_25_groupi_n_1544);
  nor csa_tree_add_7_25_groupi_g17505(csa_tree_add_7_25_groupi_n_3590 ,csa_tree_add_7_25_groupi_n_74 ,csa_tree_add_7_25_groupi_n_2010);
  nor csa_tree_add_7_25_groupi_g17506(csa_tree_add_7_25_groupi_n_3589 ,csa_tree_add_7_25_groupi_n_981 ,csa_tree_add_7_25_groupi_n_1636);
  nor csa_tree_add_7_25_groupi_g17507(csa_tree_add_7_25_groupi_n_3588 ,csa_tree_add_7_25_groupi_n_884 ,csa_tree_add_7_25_groupi_n_1157);
  nor csa_tree_add_7_25_groupi_g17508(csa_tree_add_7_25_groupi_n_3587 ,csa_tree_add_7_25_groupi_n_731 ,csa_tree_add_7_25_groupi_n_1460);
  nor csa_tree_add_7_25_groupi_g17509(csa_tree_add_7_25_groupi_n_3586 ,csa_tree_add_7_25_groupi_n_1038 ,csa_tree_add_7_25_groupi_n_134);
  nor csa_tree_add_7_25_groupi_g17510(csa_tree_add_7_25_groupi_n_3585 ,csa_tree_add_7_25_groupi_n_708 ,csa_tree_add_7_25_groupi_n_1679);
  nor csa_tree_add_7_25_groupi_g17511(csa_tree_add_7_25_groupi_n_3584 ,csa_tree_add_7_25_groupi_n_893 ,csa_tree_add_7_25_groupi_n_1301);
  nor csa_tree_add_7_25_groupi_g17512(csa_tree_add_7_25_groupi_n_3583 ,csa_tree_add_7_25_groupi_n_1056 ,csa_tree_add_7_25_groupi_n_1787);
  nor csa_tree_add_7_25_groupi_g17513(csa_tree_add_7_25_groupi_n_3582 ,csa_tree_add_7_25_groupi_n_737 ,csa_tree_add_7_25_groupi_n_1541);
  nor csa_tree_add_7_25_groupi_g17514(csa_tree_add_7_25_groupi_n_3581 ,csa_tree_add_7_25_groupi_n_1014 ,csa_tree_add_7_25_groupi_n_941);
  nor csa_tree_add_7_25_groupi_g17515(csa_tree_add_7_25_groupi_n_3580 ,csa_tree_add_7_25_groupi_n_1011 ,csa_tree_add_7_25_groupi_n_1726);
  nor csa_tree_add_7_25_groupi_g17516(csa_tree_add_7_25_groupi_n_3579 ,csa_tree_add_7_25_groupi_n_1008 ,csa_tree_add_7_25_groupi_n_1597);
  nor csa_tree_add_7_25_groupi_g17517(csa_tree_add_7_25_groupi_n_3578 ,csa_tree_add_7_25_groupi_n_1020 ,csa_tree_add_7_25_groupi_n_1478);
  nor csa_tree_add_7_25_groupi_g17518(csa_tree_add_7_25_groupi_n_3577 ,csa_tree_add_7_25_groupi_n_954 ,csa_tree_add_7_25_groupi_n_1732);
  nor csa_tree_add_7_25_groupi_g17519(csa_tree_add_7_25_groupi_n_3576 ,csa_tree_add_7_25_groupi_n_1017 ,csa_tree_add_7_25_groupi_n_1714);
  nor csa_tree_add_7_25_groupi_g17520(csa_tree_add_7_25_groupi_n_3575 ,csa_tree_add_7_25_groupi_n_957 ,csa_tree_add_7_25_groupi_n_1772);
  nor csa_tree_add_7_25_groupi_g17521(csa_tree_add_7_25_groupi_n_3574 ,csa_tree_add_7_25_groupi_n_905 ,csa_tree_add_7_25_groupi_n_1570);
  nor csa_tree_add_7_25_groupi_g17522(csa_tree_add_7_25_groupi_n_3573 ,csa_tree_add_7_25_groupi_n_1074 ,csa_tree_add_7_25_groupi_n_1343);
  nor csa_tree_add_7_25_groupi_g17523(csa_tree_add_7_25_groupi_n_3572 ,csa_tree_add_7_25_groupi_n_984 ,csa_tree_add_7_25_groupi_n_1301);
  nor csa_tree_add_7_25_groupi_g17524(csa_tree_add_7_25_groupi_n_3571 ,csa_tree_add_7_25_groupi_n_872 ,csa_tree_add_7_25_groupi_n_1555);
  nor csa_tree_add_7_25_groupi_g17525(csa_tree_add_7_25_groupi_n_3570 ,csa_tree_add_7_25_groupi_n_1059 ,csa_tree_add_7_25_groupi_n_537);
  nor csa_tree_add_7_25_groupi_g17526(csa_tree_add_7_25_groupi_n_3569 ,csa_tree_add_7_25_groupi_n_1065 ,csa_tree_add_7_25_groupi_n_1151);
  nor csa_tree_add_7_25_groupi_g17527(csa_tree_add_7_25_groupi_n_3568 ,csa_tree_add_7_25_groupi_n_1083 ,csa_tree_add_7_25_groupi_n_1454);
  nor csa_tree_add_7_25_groupi_g17528(csa_tree_add_7_25_groupi_n_3567 ,csa_tree_add_7_25_groupi_n_674 ,csa_tree_add_7_25_groupi_n_1465);
  nor csa_tree_add_7_25_groupi_g17529(csa_tree_add_7_25_groupi_n_3566 ,csa_tree_add_7_25_groupi_n_1023 ,csa_tree_add_7_25_groupi_n_1565);
  nor csa_tree_add_7_25_groupi_g17530(csa_tree_add_7_25_groupi_n_3565 ,csa_tree_add_7_25_groupi_n_1041 ,csa_tree_add_7_25_groupi_n_1571);
  nor csa_tree_add_7_25_groupi_g17531(csa_tree_add_7_25_groupi_n_3564 ,csa_tree_add_7_25_groupi_n_614 ,csa_tree_add_7_25_groupi_n_1745);
  nor csa_tree_add_7_25_groupi_g17532(csa_tree_add_7_25_groupi_n_3563 ,csa_tree_add_7_25_groupi_n_735 ,csa_tree_add_7_25_groupi_n_1385);
  nor csa_tree_add_7_25_groupi_g17533(csa_tree_add_7_25_groupi_n_3562 ,csa_tree_add_7_25_groupi_n_1053 ,csa_tree_add_7_25_groupi_n_1556);
  nor csa_tree_add_7_25_groupi_g17534(csa_tree_add_7_25_groupi_n_3561 ,csa_tree_add_7_25_groupi_n_960 ,csa_tree_add_7_25_groupi_n_1421);
  nor csa_tree_add_7_25_groupi_g17535(csa_tree_add_7_25_groupi_n_3560 ,csa_tree_add_7_25_groupi_n_1071 ,csa_tree_add_7_25_groupi_n_202);
  nor csa_tree_add_7_25_groupi_g17536(csa_tree_add_7_25_groupi_n_3559 ,csa_tree_add_7_25_groupi_n_987 ,csa_tree_add_7_25_groupi_n_1908);
  nor csa_tree_add_7_25_groupi_g17537(csa_tree_add_7_25_groupi_n_3558 ,csa_tree_add_7_25_groupi_n_923 ,csa_tree_add_7_25_groupi_n_1378);
  nor csa_tree_add_7_25_groupi_g17538(csa_tree_add_7_25_groupi_n_3557 ,csa_tree_add_7_25_groupi_n_1077 ,csa_tree_add_7_25_groupi_n_1715);
  nor csa_tree_add_7_25_groupi_g17539(csa_tree_add_7_25_groupi_n_3556 ,csa_tree_add_7_25_groupi_n_948 ,csa_tree_add_7_25_groupi_n_942);
  nor csa_tree_add_7_25_groupi_g17540(csa_tree_add_7_25_groupi_n_3555 ,csa_tree_add_7_25_groupi_n_914 ,csa_tree_add_7_25_groupi_n_1153);
  nor csa_tree_add_7_25_groupi_g17541(csa_tree_add_7_25_groupi_n_3554 ,csa_tree_add_7_25_groupi_n_654 ,csa_tree_add_7_25_groupi_n_1469);
  nor csa_tree_add_7_25_groupi_g17542(csa_tree_add_7_25_groupi_n_3553 ,csa_tree_add_7_25_groupi_n_978 ,csa_tree_add_7_25_groupi_n_1466);
  nor csa_tree_add_7_25_groupi_g17543(csa_tree_add_7_25_groupi_n_3552 ,csa_tree_add_7_25_groupi_n_969 ,csa_tree_add_7_25_groupi_n_1387);
  nor csa_tree_add_7_25_groupi_g17544(csa_tree_add_7_25_groupi_n_3551 ,csa_tree_add_7_25_groupi_n_945 ,csa_tree_add_7_25_groupi_n_1570);
  nor csa_tree_add_7_25_groupi_g17545(csa_tree_add_7_25_groupi_n_3550 ,csa_tree_add_7_25_groupi_n_677 ,csa_tree_add_7_25_groupi_n_1559);
  nor csa_tree_add_7_25_groupi_g17546(csa_tree_add_7_25_groupi_n_3549 ,csa_tree_add_7_25_groupi_n_896 ,csa_tree_add_7_25_groupi_n_1496);
  nor csa_tree_add_7_25_groupi_g17547(csa_tree_add_7_25_groupi_n_3548 ,csa_tree_add_7_25_groupi_n_743 ,csa_tree_add_7_25_groupi_n_1774);
  nor csa_tree_add_7_25_groupi_g17548(csa_tree_add_7_25_groupi_n_3547 ,csa_tree_add_7_25_groupi_n_887 ,csa_tree_add_7_25_groupi_n_1342);
  nor csa_tree_add_7_25_groupi_g17549(csa_tree_add_7_25_groupi_n_3546 ,csa_tree_add_7_25_groupi_n_722 ,csa_tree_add_7_25_groupi_n_1388);
  nor csa_tree_add_7_25_groupi_g17550(csa_tree_add_7_25_groupi_n_3545 ,csa_tree_add_7_25_groupi_n_635 ,csa_tree_add_7_25_groupi_n_166);
  or csa_tree_add_7_25_groupi_g17551(csa_tree_add_7_25_groupi_n_3544 ,csa_tree_add_7_25_groupi_n_581 ,csa_tree_add_7_25_groupi_n_2895);
  or csa_tree_add_7_25_groupi_g17552(csa_tree_add_7_25_groupi_n_3543 ,csa_tree_add_7_25_groupi_n_584 ,csa_tree_add_7_25_groupi_n_2892);
  or csa_tree_add_7_25_groupi_g17553(csa_tree_add_7_25_groupi_n_3542 ,csa_tree_add_7_25_groupi_n_28 ,csa_tree_add_7_25_groupi_n_2911);
  or csa_tree_add_7_25_groupi_g17554(csa_tree_add_7_25_groupi_n_3541 ,csa_tree_add_7_25_groupi_n_30 ,csa_tree_add_7_25_groupi_n_2906);
  or csa_tree_add_7_25_groupi_g17555(csa_tree_add_7_25_groupi_n_3540 ,csa_tree_add_7_25_groupi_n_28 ,csa_tree_add_7_25_groupi_n_2891);
  or csa_tree_add_7_25_groupi_g17556(csa_tree_add_7_25_groupi_n_3539 ,csa_tree_add_7_25_groupi_n_542 ,csa_tree_add_7_25_groupi_n_2893);
  or csa_tree_add_7_25_groupi_g17557(csa_tree_add_7_25_groupi_n_3538 ,csa_tree_add_7_25_groupi_n_545 ,csa_tree_add_7_25_groupi_n_2896);
  or csa_tree_add_7_25_groupi_g17558(csa_tree_add_7_25_groupi_n_3537 ,csa_tree_add_7_25_groupi_n_575 ,csa_tree_add_7_25_groupi_n_2894);
  or csa_tree_add_7_25_groupi_g17559(csa_tree_add_7_25_groupi_n_3536 ,csa_tree_add_7_25_groupi_n_578 ,csa_tree_add_7_25_groupi_n_2908);
  or csa_tree_add_7_25_groupi_g17560(csa_tree_add_7_25_groupi_n_3743 ,csa_tree_add_7_25_groupi_n_543 ,csa_tree_add_7_25_groupi_n_2907);
  xnor csa_tree_add_7_25_groupi_g17561(csa_tree_add_7_25_groupi_n_3742 ,csa_tree_add_7_25_groupi_n_2890 ,csa_tree_add_7_25_groupi_n_2579);
  not csa_tree_add_7_25_groupi_g17562(csa_tree_add_7_25_groupi_n_3534 ,csa_tree_add_7_25_groupi_n_3532);
  not csa_tree_add_7_25_groupi_g17563(csa_tree_add_7_25_groupi_n_3533 ,csa_tree_add_7_25_groupi_n_3532);
  not csa_tree_add_7_25_groupi_g17564(csa_tree_add_7_25_groupi_n_3531 ,csa_tree_add_7_25_groupi_n_3528);
  not csa_tree_add_7_25_groupi_g17565(csa_tree_add_7_25_groupi_n_3530 ,csa_tree_add_7_25_groupi_n_3528);
  not csa_tree_add_7_25_groupi_g17566(csa_tree_add_7_25_groupi_n_3529 ,csa_tree_add_7_25_groupi_n_3528);
  not csa_tree_add_7_25_groupi_g17568(csa_tree_add_7_25_groupi_n_3527 ,csa_tree_add_7_25_groupi_n_1990);
  not csa_tree_add_7_25_groupi_g17569(csa_tree_add_7_25_groupi_n_3525 ,csa_tree_add_7_25_groupi_n_1990);
  not csa_tree_add_7_25_groupi_g17570(csa_tree_add_7_25_groupi_n_3524 ,csa_tree_add_7_25_groupi_n_3526);
  not csa_tree_add_7_25_groupi_g17571(csa_tree_add_7_25_groupi_n_3523 ,csa_tree_add_7_25_groupi_n_1117);
  not csa_tree_add_7_25_groupi_g17573(csa_tree_add_7_25_groupi_n_3522 ,csa_tree_add_7_25_groupi_n_3521);
  not csa_tree_add_7_25_groupi_g17574(csa_tree_add_7_25_groupi_n_3520 ,csa_tree_add_7_25_groupi_n_1117);
  not csa_tree_add_7_25_groupi_g17575(csa_tree_add_7_25_groupi_n_3519 ,csa_tree_add_7_25_groupi_n_3521);
  not csa_tree_add_7_25_groupi_g17576(csa_tree_add_7_25_groupi_n_3518 ,csa_tree_add_7_25_groupi_n_3516);
  not csa_tree_add_7_25_groupi_g17577(csa_tree_add_7_25_groupi_n_3517 ,csa_tree_add_7_25_groupi_n_1987);
  not csa_tree_add_7_25_groupi_g17578(csa_tree_add_7_25_groupi_n_3515 ,csa_tree_add_7_25_groupi_n_1987);
  not csa_tree_add_7_25_groupi_g17579(csa_tree_add_7_25_groupi_n_3514 ,csa_tree_add_7_25_groupi_n_3516);
  not csa_tree_add_7_25_groupi_g17580(csa_tree_add_7_25_groupi_n_3513 ,csa_tree_add_7_25_groupi_n_3511);
  not csa_tree_add_7_25_groupi_g17581(csa_tree_add_7_25_groupi_n_3512 ,csa_tree_add_7_25_groupi_n_1981);
  not csa_tree_add_7_25_groupi_g17582(csa_tree_add_7_25_groupi_n_3510 ,csa_tree_add_7_25_groupi_n_1981);
  not csa_tree_add_7_25_groupi_g17583(csa_tree_add_7_25_groupi_n_3509 ,csa_tree_add_7_25_groupi_n_3511);
  not csa_tree_add_7_25_groupi_g17584(csa_tree_add_7_25_groupi_n_3508 ,csa_tree_add_7_25_groupi_n_3506);
  not csa_tree_add_7_25_groupi_g17585(csa_tree_add_7_25_groupi_n_3507 ,csa_tree_add_7_25_groupi_n_1977);
  not csa_tree_add_7_25_groupi_g17586(csa_tree_add_7_25_groupi_n_3505 ,csa_tree_add_7_25_groupi_n_1977);
  not csa_tree_add_7_25_groupi_g17587(csa_tree_add_7_25_groupi_n_3504 ,csa_tree_add_7_25_groupi_n_3506);
  not csa_tree_add_7_25_groupi_g17588(csa_tree_add_7_25_groupi_n_3503 ,csa_tree_add_7_25_groupi_n_3501);
  not csa_tree_add_7_25_groupi_g17589(csa_tree_add_7_25_groupi_n_3502 ,csa_tree_add_7_25_groupi_n_1975);
  not csa_tree_add_7_25_groupi_g17590(csa_tree_add_7_25_groupi_n_3500 ,csa_tree_add_7_25_groupi_n_1975);
  not csa_tree_add_7_25_groupi_g17591(csa_tree_add_7_25_groupi_n_3499 ,csa_tree_add_7_25_groupi_n_3501);
  nor csa_tree_add_7_25_groupi_g17592(csa_tree_add_7_25_groupi_n_3498 ,csa_tree_add_7_25_groupi_n_584 ,csa_tree_add_7_25_groupi_n_1757);
  or csa_tree_add_7_25_groupi_g17593(csa_tree_add_7_25_groupi_n_3497 ,csa_tree_add_7_25_groupi_n_2644 ,csa_tree_add_7_25_groupi_n_2819);
  or csa_tree_add_7_25_groupi_g17594(csa_tree_add_7_25_groupi_n_3496 ,csa_tree_add_7_25_groupi_n_2650 ,csa_tree_add_7_25_groupi_n_2721);
  nor csa_tree_add_7_25_groupi_g17595(csa_tree_add_7_25_groupi_n_3495 ,csa_tree_add_7_25_groupi_n_642 ,csa_tree_add_7_25_groupi_n_1406);
  or csa_tree_add_7_25_groupi_g17596(csa_tree_add_7_25_groupi_n_3494 ,csa_tree_add_7_25_groupi_n_2634 ,csa_tree_add_7_25_groupi_n_2824);
  or csa_tree_add_7_25_groupi_g17597(csa_tree_add_7_25_groupi_n_3493 ,csa_tree_add_7_25_groupi_n_2628 ,csa_tree_add_7_25_groupi_n_2817);
  or csa_tree_add_7_25_groupi_g17598(csa_tree_add_7_25_groupi_n_3492 ,csa_tree_add_7_25_groupi_n_2609 ,csa_tree_add_7_25_groupi_n_2712);
  or csa_tree_add_7_25_groupi_g17599(csa_tree_add_7_25_groupi_n_3491 ,csa_tree_add_7_25_groupi_n_2636 ,csa_tree_add_7_25_groupi_n_2827);
  or csa_tree_add_7_25_groupi_g17600(csa_tree_add_7_25_groupi_n_3490 ,csa_tree_add_7_25_groupi_n_2608 ,csa_tree_add_7_25_groupi_n_2713);
  or csa_tree_add_7_25_groupi_g17601(csa_tree_add_7_25_groupi_n_3489 ,csa_tree_add_7_25_groupi_n_2642 ,csa_tree_add_7_25_groupi_n_2832);
  or csa_tree_add_7_25_groupi_g17602(csa_tree_add_7_25_groupi_n_3488 ,csa_tree_add_7_25_groupi_n_2602 ,csa_tree_add_7_25_groupi_n_2710);
  or csa_tree_add_7_25_groupi_g17603(csa_tree_add_7_25_groupi_n_3487 ,csa_tree_add_7_25_groupi_n_2610 ,csa_tree_add_7_25_groupi_n_2715);
  or csa_tree_add_7_25_groupi_g17604(csa_tree_add_7_25_groupi_n_3486 ,csa_tree_add_7_25_groupi_n_2632 ,csa_tree_add_7_25_groupi_n_2815);
  or csa_tree_add_7_25_groupi_g17605(csa_tree_add_7_25_groupi_n_3485 ,csa_tree_add_7_25_groupi_n_2678 ,csa_tree_add_7_25_groupi_n_2717);
  or csa_tree_add_7_25_groupi_g17606(csa_tree_add_7_25_groupi_n_3484 ,csa_tree_add_7_25_groupi_n_2601 ,csa_tree_add_7_25_groupi_n_2708);
  or csa_tree_add_7_25_groupi_g17607(csa_tree_add_7_25_groupi_n_3483 ,csa_tree_add_7_25_groupi_n_2613 ,csa_tree_add_7_25_groupi_n_2734);
  nor csa_tree_add_7_25_groupi_g17608(csa_tree_add_7_25_groupi_n_3482 ,csa_tree_add_7_25_groupi_n_950 ,csa_tree_add_7_25_groupi_n_1373);
  or csa_tree_add_7_25_groupi_g17609(csa_tree_add_7_25_groupi_n_3481 ,csa_tree_add_7_25_groupi_n_2598 ,csa_tree_add_7_25_groupi_n_2733);
  or csa_tree_add_7_25_groupi_g17610(csa_tree_add_7_25_groupi_n_3480 ,csa_tree_add_7_25_groupi_n_2605 ,csa_tree_add_7_25_groupi_n_2731);
  or csa_tree_add_7_25_groupi_g17611(csa_tree_add_7_25_groupi_n_3479 ,csa_tree_add_7_25_groupi_n_2630 ,csa_tree_add_7_25_groupi_n_2808);
  or csa_tree_add_7_25_groupi_g17612(csa_tree_add_7_25_groupi_n_3478 ,csa_tree_add_7_25_groupi_n_2434 ,csa_tree_add_7_25_groupi_n_2890);
  or csa_tree_add_7_25_groupi_g17613(csa_tree_add_7_25_groupi_n_3477 ,csa_tree_add_7_25_groupi_n_2606 ,csa_tree_add_7_25_groupi_n_2711);
  or csa_tree_add_7_25_groupi_g17614(csa_tree_add_7_25_groupi_n_3476 ,csa_tree_add_7_25_groupi_n_2603 ,csa_tree_add_7_25_groupi_n_2707);
  or csa_tree_add_7_25_groupi_g17615(csa_tree_add_7_25_groupi_n_3475 ,csa_tree_add_7_25_groupi_n_2633 ,csa_tree_add_7_25_groupi_n_2804);
  or csa_tree_add_7_25_groupi_g17616(csa_tree_add_7_25_groupi_n_3474 ,csa_tree_add_7_25_groupi_n_2641 ,csa_tree_add_7_25_groupi_n_2830);
  or csa_tree_add_7_25_groupi_g17617(csa_tree_add_7_25_groupi_n_3473 ,csa_tree_add_7_25_groupi_n_2627 ,csa_tree_add_7_25_groupi_n_2820);
  or csa_tree_add_7_25_groupi_g17618(csa_tree_add_7_25_groupi_n_3472 ,csa_tree_add_7_25_groupi_n_2604 ,csa_tree_add_7_25_groupi_n_2714);
  or csa_tree_add_7_25_groupi_g17619(csa_tree_add_7_25_groupi_n_3471 ,csa_tree_add_7_25_groupi_n_2612 ,csa_tree_add_7_25_groupi_n_2716);
  nor csa_tree_add_7_25_groupi_g17620(csa_tree_add_7_25_groupi_n_3470 ,csa_tree_add_7_25_groupi_n_645 ,csa_tree_add_7_25_groupi_n_1403);
  nor csa_tree_add_7_25_groupi_g17621(csa_tree_add_7_25_groupi_n_3469 ,csa_tree_add_7_25_groupi_n_645 ,csa_tree_add_7_25_groupi_n_1412);
  or csa_tree_add_7_25_groupi_g17622(csa_tree_add_7_25_groupi_n_3468 ,csa_tree_add_7_25_groupi_n_2629 ,csa_tree_add_7_25_groupi_n_2813);
  or csa_tree_add_7_25_groupi_g17623(csa_tree_add_7_25_groupi_n_3467 ,csa_tree_add_7_25_groupi_n_2651 ,csa_tree_add_7_25_groupi_n_2736);
  or csa_tree_add_7_25_groupi_g17624(csa_tree_add_7_25_groupi_n_3466 ,csa_tree_add_7_25_groupi_n_2659 ,csa_tree_add_7_25_groupi_n_2730);
  or csa_tree_add_7_25_groupi_g17625(csa_tree_add_7_25_groupi_n_3465 ,csa_tree_add_7_25_groupi_n_2631 ,csa_tree_add_7_25_groupi_n_2807);
  or csa_tree_add_7_25_groupi_g17626(csa_tree_add_7_25_groupi_n_3464 ,csa_tree_add_7_25_groupi_n_2607 ,csa_tree_add_7_25_groupi_n_2706);
  or csa_tree_add_7_25_groupi_g17627(csa_tree_add_7_25_groupi_n_3463 ,csa_tree_add_7_25_groupi_n_2611 ,csa_tree_add_7_25_groupi_n_2709);
  nor csa_tree_add_7_25_groupi_g17628(csa_tree_add_7_25_groupi_n_3462 ,csa_tree_add_7_25_groupi_n_641 ,csa_tree_add_7_25_groupi_n_1367);
  nor csa_tree_add_7_25_groupi_g17629(csa_tree_add_7_25_groupi_n_3461 ,csa_tree_add_7_25_groupi_n_951 ,csa_tree_add_7_25_groupi_n_1700);
  nor csa_tree_add_7_25_groupi_g17630(csa_tree_add_7_25_groupi_n_3460 ,csa_tree_add_7_25_groupi_n_644 ,csa_tree_add_7_25_groupi_n_1463);
  nor csa_tree_add_7_25_groupi_g17631(csa_tree_add_7_25_groupi_n_3459 ,csa_tree_add_7_25_groupi_n_623 ,csa_tree_add_7_25_groupi_n_1442);
  nor csa_tree_add_7_25_groupi_g17632(csa_tree_add_7_25_groupi_n_3458 ,csa_tree_add_7_25_groupi_n_642 ,csa_tree_add_7_25_groupi_n_1487);
  nor csa_tree_add_7_25_groupi_g17633(csa_tree_add_7_25_groupi_n_3457 ,csa_tree_add_7_25_groupi_n_627 ,csa_tree_add_7_25_groupi_n_1352);
  nor csa_tree_add_7_25_groupi_g17634(csa_tree_add_7_25_groupi_n_3456 ,csa_tree_add_7_25_groupi_n_630 ,csa_tree_add_7_25_groupi_n_1245);
  nor csa_tree_add_7_25_groupi_g17635(csa_tree_add_7_25_groupi_n_3455 ,csa_tree_add_7_25_groupi_n_101 ,csa_tree_add_7_25_groupi_n_1236);
  nor csa_tree_add_7_25_groupi_g17636(csa_tree_add_7_25_groupi_n_3454 ,csa_tree_add_7_25_groupi_n_1000 ,csa_tree_add_7_25_groupi_n_1230);
  nor csa_tree_add_7_25_groupi_g17637(csa_tree_add_7_25_groupi_n_3453 ,csa_tree_add_7_25_groupi_n_629 ,csa_tree_add_7_25_groupi_n_1242);
  nor csa_tree_add_7_25_groupi_g17638(csa_tree_add_7_25_groupi_n_3452 ,csa_tree_add_7_25_groupi_n_632 ,csa_tree_add_7_25_groupi_n_1148);
  nor csa_tree_add_7_25_groupi_g17639(csa_tree_add_7_25_groupi_n_3451 ,csa_tree_add_7_25_groupi_n_1002 ,csa_tree_add_7_25_groupi_n_1639);
  nor csa_tree_add_7_25_groupi_g17640(csa_tree_add_7_25_groupi_n_3450 ,csa_tree_add_7_25_groupi_n_1089 ,csa_tree_add_7_25_groupi_n_1621);
  nor csa_tree_add_7_25_groupi_g17641(csa_tree_add_7_25_groupi_n_3449 ,csa_tree_add_7_25_groupi_n_104 ,csa_tree_add_7_25_groupi_n_1603);
  nor csa_tree_add_7_25_groupi_g17642(csa_tree_add_7_25_groupi_n_3448 ,csa_tree_add_7_25_groupi_n_633 ,csa_tree_add_7_25_groupi_n_1612);
  nor csa_tree_add_7_25_groupi_g17643(csa_tree_add_7_25_groupi_n_3447 ,csa_tree_add_7_25_groupi_n_1889 ,csa_tree_add_7_25_groupi_n_1325);
  nor csa_tree_add_7_25_groupi_g17644(csa_tree_add_7_25_groupi_n_3446 ,csa_tree_add_7_25_groupi_n_215 ,csa_tree_add_7_25_groupi_n_1639);
  nor csa_tree_add_7_25_groupi_g17645(csa_tree_add_7_25_groupi_n_3445 ,csa_tree_add_7_25_groupi_n_629 ,csa_tree_add_7_25_groupi_n_1502);
  nor csa_tree_add_7_25_groupi_g17646(csa_tree_add_7_25_groupi_n_3444 ,csa_tree_add_7_25_groupi_n_994 ,csa_tree_add_7_25_groupi_n_1490);
  nor csa_tree_add_7_25_groupi_g17647(csa_tree_add_7_25_groupi_n_3443 ,csa_tree_add_7_25_groupi_n_999 ,csa_tree_add_7_25_groupi_n_1526);
  nor csa_tree_add_7_25_groupi_g17648(csa_tree_add_7_25_groupi_n_3442 ,csa_tree_add_7_25_groupi_n_627 ,csa_tree_add_7_25_groupi_n_1233);
  nor csa_tree_add_7_25_groupi_g17649(csa_tree_add_7_25_groupi_n_3441 ,csa_tree_add_7_25_groupi_n_630 ,csa_tree_add_7_25_groupi_n_1439);
  nor csa_tree_add_7_25_groupi_g17650(csa_tree_add_7_25_groupi_n_3440 ,csa_tree_add_7_25_groupi_n_239 ,csa_tree_add_7_25_groupi_n_1621);
  nor csa_tree_add_7_25_groupi_g17651(csa_tree_add_7_25_groupi_n_3439 ,csa_tree_add_7_25_groupi_n_462 ,csa_tree_add_7_25_groupi_n_1612);
  nor csa_tree_add_7_25_groupi_g17652(csa_tree_add_7_25_groupi_n_3438 ,csa_tree_add_7_25_groupi_n_463 ,csa_tree_add_7_25_groupi_n_1603);
  nor csa_tree_add_7_25_groupi_g17653(csa_tree_add_7_25_groupi_n_3437 ,csa_tree_add_7_25_groupi_n_220 ,csa_tree_add_7_25_groupi_n_1330);
  nor csa_tree_add_7_25_groupi_g17654(csa_tree_add_7_25_groupi_n_3436 ,csa_tree_add_7_25_groupi_n_1891 ,csa_tree_add_7_25_groupi_n_1239);
  nor csa_tree_add_7_25_groupi_g17655(csa_tree_add_7_25_groupi_n_3435 ,csa_tree_add_7_25_groupi_n_1893 ,csa_tree_add_7_25_groupi_n_1645);
  nor csa_tree_add_7_25_groupi_g17656(csa_tree_add_7_25_groupi_n_3434 ,csa_tree_add_7_25_groupi_n_1895 ,csa_tree_add_7_25_groupi_n_1594);
  nor csa_tree_add_7_25_groupi_g17657(csa_tree_add_7_25_groupi_n_3433 ,csa_tree_add_7_25_groupi_n_232 ,csa_tree_add_7_25_groupi_n_1627);
  nor csa_tree_add_7_25_groupi_g17658(csa_tree_add_7_25_groupi_n_3432 ,csa_tree_add_7_25_groupi_n_466 ,csa_tree_add_7_25_groupi_n_1360);
  nor csa_tree_add_7_25_groupi_g17659(csa_tree_add_7_25_groupi_n_3431 ,csa_tree_add_7_25_groupi_n_115 ,csa_tree_add_7_25_groupi_n_1334);
  nor csa_tree_add_7_25_groupi_g17660(csa_tree_add_7_25_groupi_n_3430 ,csa_tree_add_7_25_groupi_n_115 ,csa_tree_add_7_25_groupi_n_1550);
  nor csa_tree_add_7_25_groupi_g17661(csa_tree_add_7_25_groupi_n_3429 ,csa_tree_add_7_25_groupi_n_996 ,csa_tree_add_7_25_groupi_n_1666);
  nor csa_tree_add_7_25_groupi_g17662(csa_tree_add_7_25_groupi_n_3428 ,csa_tree_add_7_25_groupi_n_632 ,csa_tree_add_7_25_groupi_n_1781);
  nor csa_tree_add_7_25_groupi_g17663(csa_tree_add_7_25_groupi_n_3427 ,csa_tree_add_7_25_groupi_n_1002 ,csa_tree_add_7_25_groupi_n_1676);
  nor csa_tree_add_7_25_groupi_g17664(csa_tree_add_7_25_groupi_n_3426 ,csa_tree_add_7_25_groupi_n_1089 ,csa_tree_add_7_25_groupi_n_1376);
  nor csa_tree_add_7_25_groupi_g17665(csa_tree_add_7_25_groupi_n_3425 ,csa_tree_add_7_25_groupi_n_448 ,csa_tree_add_7_25_groupi_n_1997);
  nor csa_tree_add_7_25_groupi_g17666(csa_tree_add_7_25_groupi_n_3424 ,csa_tree_add_7_25_groupi_n_1897 ,csa_tree_add_7_25_groupi_n_1325);
  nor csa_tree_add_7_25_groupi_g17667(csa_tree_add_7_25_groupi_n_3423 ,csa_tree_add_7_25_groupi_n_1899 ,csa_tree_add_7_25_groupi_n_1648);
  nor csa_tree_add_7_25_groupi_g17668(csa_tree_add_7_25_groupi_n_3422 ,csa_tree_add_7_25_groupi_n_229 ,csa_tree_add_7_25_groupi_n_1633);
  nor csa_tree_add_7_25_groupi_g17669(csa_tree_add_7_25_groupi_n_3421 ,csa_tree_add_7_25_groupi_n_235 ,csa_tree_add_7_25_groupi_n_1615);
  nor csa_tree_add_7_25_groupi_g17670(csa_tree_add_7_25_groupi_n_3420 ,csa_tree_add_7_25_groupi_n_448 ,csa_tree_add_7_25_groupi_n_1606);
  nor csa_tree_add_7_25_groupi_g17671(csa_tree_add_7_25_groupi_n_3419 ,csa_tree_add_7_25_groupi_n_1881 ,csa_tree_add_7_25_groupi_n_1507);
  nor csa_tree_add_7_25_groupi_g17672(csa_tree_add_7_25_groupi_n_3418 ,csa_tree_add_7_25_groupi_n_1883 ,csa_tree_add_7_25_groupi_n_1444);
  nor csa_tree_add_7_25_groupi_g17673(csa_tree_add_7_25_groupi_n_3417 ,csa_tree_add_7_25_groupi_n_1887 ,csa_tree_add_7_25_groupi_n_1166);
  nor csa_tree_add_7_25_groupi_g17674(csa_tree_add_7_25_groupi_n_3416 ,csa_tree_add_7_25_groupi_n_1889 ,csa_tree_add_7_25_groupi_n_1519);
  nor csa_tree_add_7_25_groupi_g17675(csa_tree_add_7_25_groupi_n_3415 ,csa_tree_add_7_25_groupi_n_214 ,csa_tree_add_7_25_groupi_n_1666);
  nor csa_tree_add_7_25_groupi_g17676(csa_tree_add_7_25_groupi_n_3414 ,csa_tree_add_7_25_groupi_n_238 ,csa_tree_add_7_25_groupi_n_1531);
  nor csa_tree_add_7_25_groupi_g17677(csa_tree_add_7_25_groupi_n_3413 ,csa_tree_add_7_25_groupi_n_451 ,csa_tree_add_7_25_groupi_n_1337);
  nor csa_tree_add_7_25_groupi_g17678(csa_tree_add_7_25_groupi_n_3412 ,csa_tree_add_7_25_groupi_n_243 ,csa_tree_add_7_25_groupi_n_1720);
  nor csa_tree_add_7_25_groupi_g17679(csa_tree_add_7_25_groupi_n_3411 ,csa_tree_add_7_25_groupi_n_1885 ,csa_tree_add_7_25_groupi_n_1663);
  nor csa_tree_add_7_25_groupi_g17680(csa_tree_add_7_25_groupi_n_3410 ,csa_tree_add_7_25_groupi_n_223 ,csa_tree_add_7_25_groupi_n_1364);
  nor csa_tree_add_7_25_groupi_g17681(csa_tree_add_7_25_groupi_n_3409 ,csa_tree_add_7_25_groupi_n_226 ,csa_tree_add_7_25_groupi_n_1601);
  nor csa_tree_add_7_25_groupi_g17682(csa_tree_add_7_25_groupi_n_3408 ,csa_tree_add_7_25_groupi_n_459 ,csa_tree_add_7_25_groupi_n_1631);
  nor csa_tree_add_7_25_groupi_g17683(csa_tree_add_7_25_groupi_n_3407 ,csa_tree_add_7_25_groupi_n_298 ,csa_tree_add_7_25_groupi_n_1391);
  nor csa_tree_add_7_25_groupi_g17684(csa_tree_add_7_25_groupi_n_3406 ,csa_tree_add_7_25_groupi_n_217 ,csa_tree_add_7_25_groupi_n_1793);
  nor csa_tree_add_7_25_groupi_g17685(csa_tree_add_7_25_groupi_n_3405 ,csa_tree_add_7_25_groupi_n_478 ,csa_tree_add_7_25_groupi_n_1672);
  nor csa_tree_add_7_25_groupi_g17686(csa_tree_add_7_25_groupi_n_3404 ,csa_tree_add_7_25_groupi_n_469 ,csa_tree_add_7_25_groupi_n_1369);
  nor csa_tree_add_7_25_groupi_g17687(csa_tree_add_7_25_groupi_n_3403 ,csa_tree_add_7_25_groupi_n_221 ,csa_tree_add_7_25_groupi_n_1522);
  nor csa_tree_add_7_25_groupi_g17688(csa_tree_add_7_25_groupi_n_3402 ,csa_tree_add_7_25_groupi_n_1891 ,csa_tree_add_7_25_groupi_n_2003);
  nor csa_tree_add_7_25_groupi_g17689(csa_tree_add_7_25_groupi_n_3401 ,csa_tree_add_7_25_groupi_n_1893 ,csa_tree_add_7_25_groupi_n_1510);
  nor csa_tree_add_7_25_groupi_g17690(csa_tree_add_7_25_groupi_n_3400 ,csa_tree_add_7_25_groupi_n_1895 ,csa_tree_add_7_25_groupi_n_1498);
  nor csa_tree_add_7_25_groupi_g17691(csa_tree_add_7_25_groupi_n_3399 ,csa_tree_add_7_25_groupi_n_365 ,csa_tree_add_7_25_groupi_n_1721);
  nor csa_tree_add_7_25_groupi_g17692(csa_tree_add_7_25_groupi_n_3398 ,csa_tree_add_7_25_groupi_n_408 ,csa_tree_add_7_25_groupi_n_1661);
  nor csa_tree_add_7_25_groupi_g17693(csa_tree_add_7_25_groupi_n_3397 ,csa_tree_add_7_25_groupi_n_831 ,csa_tree_add_7_25_groupi_n_504);
  or csa_tree_add_7_25_groupi_g17694(csa_tree_add_7_25_groupi_n_3396 ,csa_tree_add_7_25_groupi_n_44 ,csa_tree_add_7_25_groupi_n_495);
  nor csa_tree_add_7_25_groupi_g17695(csa_tree_add_7_25_groupi_n_3395 ,csa_tree_add_7_25_groupi_n_438 ,csa_tree_add_7_25_groupi_n_1643);
  nor csa_tree_add_7_25_groupi_g17696(csa_tree_add_7_25_groupi_n_3394 ,csa_tree_add_7_25_groupi_n_397 ,csa_tree_add_7_25_groupi_n_1625);
  nor csa_tree_add_7_25_groupi_g17697(csa_tree_add_7_25_groupi_n_3393 ,csa_tree_add_7_25_groupi_n_423 ,csa_tree_add_7_25_groupi_n_1397);
  nor csa_tree_add_7_25_groupi_g17698(csa_tree_add_7_25_groupi_n_3392 ,csa_tree_add_7_25_groupi_n_390 ,csa_tree_add_7_25_groupi_n_1400);
  nor csa_tree_add_7_25_groupi_g17699(csa_tree_add_7_25_groupi_n_3391 ,csa_tree_add_7_25_groupi_n_368 ,csa_tree_add_7_25_groupi_n_1337);
  nor csa_tree_add_7_25_groupi_g17700(csa_tree_add_7_25_groupi_n_3390 ,csa_tree_add_7_25_groupi_n_341 ,csa_tree_add_7_25_groupi_n_1931);
  or csa_tree_add_7_25_groupi_g17701(csa_tree_add_7_25_groupi_n_3389 ,csa_tree_add_7_25_groupi_n_88 ,csa_tree_add_7_25_groupi_n_497);
  nor csa_tree_add_7_25_groupi_g17702(csa_tree_add_7_25_groupi_n_3388 ,csa_tree_add_7_25_groupi_n_421 ,csa_tree_add_7_25_groupi_n_1760);
  or csa_tree_add_7_25_groupi_g17703(csa_tree_add_7_25_groupi_n_3387 ,csa_tree_add_7_25_groupi_n_2655 ,csa_tree_add_7_25_groupi_n_2732);
  or csa_tree_add_7_25_groupi_g17704(csa_tree_add_7_25_groupi_n_3386 ,csa_tree_add_7_25_groupi_n_935 ,csa_tree_add_7_25_groupi_n_512);
  nor csa_tree_add_7_25_groupi_g17705(csa_tree_add_7_25_groupi_n_3385 ,csa_tree_add_7_25_groupi_n_935 ,csa_tree_add_7_25_groupi_n_1423);
  nor csa_tree_add_7_25_groupi_g17706(csa_tree_add_7_25_groupi_n_3384 ,csa_tree_add_7_25_groupi_n_445 ,csa_tree_add_7_25_groupi_n_1450);
  nor csa_tree_add_7_25_groupi_g17707(csa_tree_add_7_25_groupi_n_3383 ,csa_tree_add_7_25_groupi_n_485 ,csa_tree_add_7_25_groupi_n_1340);
  nor csa_tree_add_7_25_groupi_g17708(csa_tree_add_7_25_groupi_n_3382 ,csa_tree_add_7_25_groupi_n_447 ,csa_tree_add_7_25_groupi_n_1414);
  nor csa_tree_add_7_25_groupi_g17709(csa_tree_add_7_25_groupi_n_3381 ,csa_tree_add_7_25_groupi_n_1897 ,csa_tree_add_7_25_groupi_n_1681);
  nor csa_tree_add_7_25_groupi_g17710(csa_tree_add_7_25_groupi_n_3380 ,csa_tree_add_7_25_groupi_n_1899 ,csa_tree_add_7_25_groupi_n_1435);
  nor csa_tree_add_7_25_groupi_g17711(csa_tree_add_7_25_groupi_n_3379 ,csa_tree_add_7_25_groupi_n_230 ,csa_tree_add_7_25_groupi_n_1777);
  nor csa_tree_add_7_25_groupi_g17712(csa_tree_add_7_25_groupi_n_3378 ,csa_tree_add_7_25_groupi_n_236 ,csa_tree_add_7_25_groupi_n_1735);
  nor csa_tree_add_7_25_groupi_g17713(csa_tree_add_7_25_groupi_n_3377 ,csa_tree_add_7_25_groupi_n_374 ,csa_tree_add_7_25_groupi_n_1657);
  nor csa_tree_add_7_25_groupi_g17714(csa_tree_add_7_25_groupi_n_3376 ,csa_tree_add_7_25_groupi_n_357 ,csa_tree_add_7_25_groupi_n_1364);
  nor csa_tree_add_7_25_groupi_g17715(csa_tree_add_7_25_groupi_n_3375 ,csa_tree_add_7_25_groupi_n_381 ,csa_tree_add_7_25_groupi_n_1601);
  nor csa_tree_add_7_25_groupi_g17716(csa_tree_add_7_25_groupi_n_3374 ,csa_tree_add_7_25_groupi_n_376 ,csa_tree_add_7_25_groupi_n_1631);
  nor csa_tree_add_7_25_groupi_g17717(csa_tree_add_7_25_groupi_n_3373 ,csa_tree_add_7_25_groupi_n_374 ,csa_tree_add_7_25_groupi_n_1391);
  or csa_tree_add_7_25_groupi_g17718(csa_tree_add_7_25_groupi_n_3372 ,csa_tree_add_7_25_groupi_n_50 ,csa_tree_add_7_25_groupi_n_497);
  nor csa_tree_add_7_25_groupi_g17719(csa_tree_add_7_25_groupi_n_3371 ,csa_tree_add_7_25_groupi_n_699 ,csa_tree_add_7_25_groupi_n_501);
  or csa_tree_add_7_25_groupi_g17720(csa_tree_add_7_25_groupi_n_3370 ,csa_tree_add_7_25_groupi_n_78 ,csa_tree_add_7_25_groupi_n_498);
  or csa_tree_add_7_25_groupi_g17721(csa_tree_add_7_25_groupi_n_3369 ,csa_tree_add_7_25_groupi_n_92 ,csa_tree_add_7_25_groupi_n_500);
  or csa_tree_add_7_25_groupi_g17722(csa_tree_add_7_25_groupi_n_3368 ,csa_tree_add_7_25_groupi_n_82 ,csa_tree_add_7_25_groupi_n_494);
  or csa_tree_add_7_25_groupi_g17723(csa_tree_add_7_25_groupi_n_3367 ,csa_tree_add_7_25_groupi_n_26 ,csa_tree_add_7_25_groupi_n_494);
  or csa_tree_add_7_25_groupi_g17724(csa_tree_add_7_25_groupi_n_3366 ,csa_tree_add_7_25_groupi_n_54 ,csa_tree_add_7_25_groupi_n_498);
  or csa_tree_add_7_25_groupi_g17725(csa_tree_add_7_25_groupi_n_3365 ,csa_tree_add_7_25_groupi_n_84 ,csa_tree_add_7_25_groupi_n_495);
  or csa_tree_add_7_25_groupi_g17726(csa_tree_add_7_25_groupi_n_3364 ,csa_tree_add_7_25_groupi_n_86 ,csa_tree_add_7_25_groupi_n_504);
  or csa_tree_add_7_25_groupi_g17727(csa_tree_add_7_25_groupi_n_3363 ,csa_tree_add_7_25_groupi_n_112 ,csa_tree_add_7_25_groupi_n_503);
  or csa_tree_add_7_25_groupi_g17728(csa_tree_add_7_25_groupi_n_3362 ,csa_tree_add_7_25_groupi_n_72 ,csa_tree_add_7_25_groupi_n_503);
  or csa_tree_add_7_25_groupi_g17729(csa_tree_add_7_25_groupi_n_3361 ,csa_tree_add_7_25_groupi_n_74 ,csa_tree_add_7_25_groupi_n_500);
  nor csa_tree_add_7_25_groupi_g17730(csa_tree_add_7_25_groupi_n_3360 ,csa_tree_add_7_25_groupi_n_384 ,csa_tree_add_7_25_groupi_n_1789);
  nor csa_tree_add_7_25_groupi_g17731(csa_tree_add_7_25_groupi_n_3359 ,csa_tree_add_7_25_groupi_n_406 ,csa_tree_add_7_25_groupi_n_524);
  nor csa_tree_add_7_25_groupi_g17732(csa_tree_add_7_25_groupi_n_3358 ,csa_tree_add_7_25_groupi_n_792 ,csa_tree_add_7_25_groupi_n_1606);
  nor csa_tree_add_7_25_groupi_g17733(csa_tree_add_7_25_groupi_n_3357 ,csa_tree_add_7_25_groupi_n_822 ,csa_tree_add_7_25_groupi_n_1615);
  nor csa_tree_add_7_25_groupi_g17734(csa_tree_add_7_25_groupi_n_3356 ,csa_tree_add_7_25_groupi_n_762 ,csa_tree_add_7_25_groupi_n_1747);
  nor csa_tree_add_7_25_groupi_g17735(csa_tree_add_7_25_groupi_n_3355 ,csa_tree_add_7_25_groupi_n_600 ,csa_tree_add_7_25_groupi_n_1306);
  nor csa_tree_add_7_25_groupi_g17736(csa_tree_add_7_25_groupi_n_3354 ,csa_tree_add_7_25_groupi_n_350 ,csa_tree_add_7_25_groupi_n_1663);
  nor csa_tree_add_7_25_groupi_g17737(csa_tree_add_7_25_groupi_n_3353 ,csa_tree_add_7_25_groupi_n_456 ,csa_tree_add_7_25_groupi_n_1777);
  nor csa_tree_add_7_25_groupi_g17738(csa_tree_add_7_25_groupi_n_3352 ,csa_tree_add_7_25_groupi_n_453 ,csa_tree_add_7_25_groupi_n_1522);
  nor csa_tree_add_7_25_groupi_g17739(csa_tree_add_7_25_groupi_n_3351 ,csa_tree_add_7_25_groupi_n_450 ,csa_tree_add_7_25_groupi_n_1448);
  nor csa_tree_add_7_25_groupi_g17740(csa_tree_add_7_25_groupi_n_3350 ,csa_tree_add_7_25_groupi_n_246 ,csa_tree_add_7_25_groupi_n_297);
  nor csa_tree_add_7_25_groupi_g17741(csa_tree_add_7_25_groupi_n_3349 ,csa_tree_add_7_25_groupi_n_224 ,csa_tree_add_7_25_groupi_n_1562);
  nor csa_tree_add_7_25_groupi_g17742(csa_tree_add_7_25_groupi_n_3348 ,csa_tree_add_7_25_groupi_n_227 ,csa_tree_add_7_25_groupi_n_1394);
  nor csa_tree_add_7_25_groupi_g17743(csa_tree_add_7_25_groupi_n_3347 ,csa_tree_add_7_25_groupi_n_460 ,csa_tree_add_7_25_groupi_n_1433);
  nor csa_tree_add_7_25_groupi_g17744(csa_tree_add_7_25_groupi_n_3346 ,csa_tree_add_7_25_groupi_n_429 ,csa_tree_add_7_25_groupi_n_1648);
  nor csa_tree_add_7_25_groupi_g17745(csa_tree_add_7_25_groupi_n_3345 ,csa_tree_add_7_25_groupi_n_411 ,csa_tree_add_7_25_groupi_n_1360);
  nor csa_tree_add_7_25_groupi_g17746(csa_tree_add_7_25_groupi_n_3344 ,csa_tree_add_7_25_groupi_n_351 ,csa_tree_add_7_25_groupi_n_1594);
  nor csa_tree_add_7_25_groupi_g17747(csa_tree_add_7_25_groupi_n_3343 ,csa_tree_add_7_25_groupi_n_560 ,csa_tree_add_7_25_groupi_n_1633);
  nor csa_tree_add_7_25_groupi_g17748(csa_tree_add_7_25_groupi_n_3342 ,csa_tree_add_7_25_groupi_n_475 ,csa_tree_add_7_25_groupi_n_1303);
  nor csa_tree_add_7_25_groupi_g17749(csa_tree_add_7_25_groupi_n_3341 ,csa_tree_add_7_25_groupi_n_417 ,csa_tree_add_7_25_groupi_n_1330);
  nor csa_tree_add_7_25_groupi_g17750(csa_tree_add_7_25_groupi_n_3340 ,csa_tree_add_7_25_groupi_n_393 ,csa_tree_add_7_25_groupi_n_124);
  nor csa_tree_add_7_25_groupi_g17751(csa_tree_add_7_25_groupi_n_3339 ,csa_tree_add_7_25_groupi_n_648 ,csa_tree_add_7_25_groupi_n_129);
  nor csa_tree_add_7_25_groupi_g17752(csa_tree_add_7_25_groupi_n_3338 ,csa_tree_add_7_25_groupi_n_684 ,csa_tree_add_7_25_groupi_n_1607);
  nor csa_tree_add_7_25_groupi_g17753(csa_tree_add_7_25_groupi_n_3337 ,csa_tree_add_7_25_groupi_n_563 ,csa_tree_add_7_25_groupi_n_1661);
  nor csa_tree_add_7_25_groupi_g17754(csa_tree_add_7_25_groupi_n_3336 ,csa_tree_add_7_25_groupi_n_566 ,csa_tree_add_7_25_groupi_n_1645);
  nor csa_tree_add_7_25_groupi_g17755(csa_tree_add_7_25_groupi_n_3335 ,csa_tree_add_7_25_groupi_n_603 ,csa_tree_add_7_25_groupi_n_524);
  nor csa_tree_add_7_25_groupi_g17756(csa_tree_add_7_25_groupi_n_3334 ,csa_tree_add_7_25_groupi_n_761 ,csa_tree_add_7_25_groupi_n_1627);
  nor csa_tree_add_7_25_groupi_g17757(csa_tree_add_7_25_groupi_n_3333 ,csa_tree_add_7_25_groupi_n_353 ,csa_tree_add_7_25_groupi_n_1616);
  nor csa_tree_add_7_25_groupi_g17758(csa_tree_add_7_25_groupi_n_3332 ,csa_tree_add_7_25_groupi_n_345 ,csa_tree_add_7_25_groupi_n_1610);
  nor csa_tree_add_7_25_groupi_g17759(csa_tree_add_7_25_groupi_n_3331 ,csa_tree_add_7_25_groupi_n_396 ,csa_tree_add_7_25_groupi_n_1369);
  nor csa_tree_add_7_25_groupi_g17760(csa_tree_add_7_25_groupi_n_3330 ,csa_tree_add_7_25_groupi_n_244 ,csa_tree_add_7_25_groupi_n_1670);
  nor csa_tree_add_7_25_groupi_g17761(csa_tree_add_7_25_groupi_n_3329 ,csa_tree_add_7_25_groupi_n_218 ,csa_tree_add_7_25_groupi_n_1510);
  nor csa_tree_add_7_25_groupi_g17762(csa_tree_add_7_25_groupi_n_3328 ,csa_tree_add_7_25_groupi_n_409 ,csa_tree_add_7_25_groupi_n_1346);
  nor csa_tree_add_7_25_groupi_g17763(csa_tree_add_7_25_groupi_n_3327 ,csa_tree_add_7_25_groupi_n_439 ,csa_tree_add_7_25_groupi_n_1340);
  nor csa_tree_add_7_25_groupi_g17764(csa_tree_add_7_25_groupi_n_3326 ,csa_tree_add_7_25_groupi_n_348 ,csa_tree_add_7_25_groupi_n_1729);
  nor csa_tree_add_7_25_groupi_g17765(csa_tree_add_7_25_groupi_n_3325 ,csa_tree_add_7_25_groupi_n_424 ,csa_tree_add_7_25_groupi_n_1498);
  nor csa_tree_add_7_25_groupi_g17766(csa_tree_add_7_25_groupi_n_3324 ,csa_tree_add_7_25_groupi_n_597 ,csa_tree_add_7_25_groupi_n_1306);
  nor csa_tree_add_7_25_groupi_g17767(csa_tree_add_7_25_groupi_n_3323 ,csa_tree_add_7_25_groupi_n_359 ,csa_tree_add_7_25_groupi_n_1793);
  nor csa_tree_add_7_25_groupi_g17768(csa_tree_add_7_25_groupi_n_3322 ,csa_tree_add_7_25_groupi_n_591 ,csa_tree_add_7_25_groupi_n_1760);
  nor csa_tree_add_7_25_groupi_g17769(csa_tree_add_7_25_groupi_n_3321 ,csa_tree_add_7_25_groupi_n_765 ,csa_tree_add_7_25_groupi_n_1657);
  nor csa_tree_add_7_25_groupi_g17770(csa_tree_add_7_25_groupi_n_3320 ,csa_tree_add_7_25_groupi_n_795 ,csa_tree_add_7_25_groupi_n_1313);
  nor csa_tree_add_7_25_groupi_g17771(csa_tree_add_7_25_groupi_n_3319 ,csa_tree_add_7_25_groupi_n_768 ,csa_tree_add_7_25_groupi_n_1649);
  nor csa_tree_add_7_25_groupi_g17772(csa_tree_add_7_25_groupi_n_3318 ,csa_tree_add_7_25_groupi_n_693 ,csa_tree_add_7_25_groupi_n_1619);
  nor csa_tree_add_7_25_groupi_g17773(csa_tree_add_7_25_groupi_n_3317 ,csa_tree_add_7_25_groupi_n_930 ,csa_tree_add_7_25_groupi_n_1901);
  nor csa_tree_add_7_25_groupi_g17774(csa_tree_add_7_25_groupi_n_3316 ,csa_tree_add_7_25_groupi_n_864 ,csa_tree_add_7_25_groupi_n_1902);
  nor csa_tree_add_7_25_groupi_g17775(csa_tree_add_7_25_groupi_n_3315 ,csa_tree_add_7_25_groupi_n_569 ,csa_tree_add_7_25_groupi_n_1595);
  nor csa_tree_add_7_25_groupi_g17776(csa_tree_add_7_25_groupi_n_3314 ,csa_tree_add_7_25_groupi_n_572 ,csa_tree_add_7_25_groupi_n_1634);
  nor csa_tree_add_7_25_groupi_g17777(csa_tree_add_7_25_groupi_n_3313 ,csa_tree_add_7_25_groupi_n_402 ,csa_tree_add_7_25_groupi_n_1361);
  nor csa_tree_add_7_25_groupi_g17778(csa_tree_add_7_25_groupi_n_3312 ,csa_tree_add_7_25_groupi_n_771 ,csa_tree_add_7_25_groupi_n_2016);
  nor csa_tree_add_7_25_groupi_g17779(csa_tree_add_7_25_groupi_n_3311 ,csa_tree_add_7_25_groupi_n_786 ,csa_tree_add_7_25_groupi_n_1750);
  nor csa_tree_add_7_25_groupi_g17780(csa_tree_add_7_25_groupi_n_3310 ,csa_tree_add_7_25_groupi_n_539 ,csa_tree_add_7_25_groupi_n_1394);
  nor csa_tree_add_7_25_groupi_g17781(csa_tree_add_7_25_groupi_n_3309 ,csa_tree_add_7_25_groupi_n_364 ,csa_tree_add_7_25_groupi_n_1423);
  nor csa_tree_add_7_25_groupi_g17782(csa_tree_add_7_25_groupi_n_3308 ,csa_tree_add_7_25_groupi_n_367 ,csa_tree_add_7_25_groupi_n_1448);
  nor csa_tree_add_7_25_groupi_g17783(csa_tree_add_7_25_groupi_n_3307 ,csa_tree_add_7_25_groupi_n_373 ,csa_tree_add_7_25_groupi_n_1756);
  nor csa_tree_add_7_25_groupi_g17784(csa_tree_add_7_25_groupi_n_3306 ,csa_tree_add_7_25_groupi_n_356 ,csa_tree_add_7_25_groupi_n_136);
  nor csa_tree_add_7_25_groupi_g17785(csa_tree_add_7_25_groupi_n_3305 ,csa_tree_add_7_25_groupi_n_382 ,csa_tree_add_7_25_groupi_n_1781);
  nor csa_tree_add_7_25_groupi_g17786(csa_tree_add_7_25_groupi_n_3304 ,csa_tree_add_7_25_groupi_n_377 ,csa_tree_add_7_25_groupi_n_1433);
  nor csa_tree_add_7_25_groupi_g17787(csa_tree_add_7_25_groupi_n_3303 ,csa_tree_add_7_25_groupi_n_371 ,csa_tree_add_7_25_groupi_n_1562);
  nor csa_tree_add_7_25_groupi_g17788(csa_tree_add_7_25_groupi_n_3302 ,csa_tree_add_7_25_groupi_n_702 ,csa_tree_add_7_25_groupi_n_1848);
  nor csa_tree_add_7_25_groupi_g17789(csa_tree_add_7_25_groupi_n_3301 ,csa_tree_add_7_25_groupi_n_657 ,csa_tree_add_7_25_groupi_n_1922);
  nor csa_tree_add_7_25_groupi_g17790(csa_tree_add_7_25_groupi_n_3300 ,csa_tree_add_7_25_groupi_n_774 ,csa_tree_add_7_25_groupi_n_1655);
  nor csa_tree_add_7_25_groupi_g17791(csa_tree_add_7_25_groupi_n_3299 ,csa_tree_add_7_25_groupi_n_780 ,csa_tree_add_7_25_groupi_n_1652);
  nor csa_tree_add_7_25_groupi_g17792(csa_tree_add_7_25_groupi_n_3298 ,csa_tree_add_7_25_groupi_n_789 ,csa_tree_add_7_25_groupi_n_2015);
  nor csa_tree_add_7_25_groupi_g17793(csa_tree_add_7_25_groupi_n_3297 ,csa_tree_add_7_25_groupi_n_612 ,csa_tree_add_7_25_groupi_n_1751);
  nor csa_tree_add_7_25_groupi_g17794(csa_tree_add_7_25_groupi_n_3296 ,csa_tree_add_7_25_groupi_n_587 ,csa_tree_add_7_25_groupi_n_1604);
  nor csa_tree_add_7_25_groupi_g17795(csa_tree_add_7_25_groupi_n_3295 ,csa_tree_add_7_25_groupi_n_779 ,csa_tree_add_7_25_groupi_n_1358);
  nor csa_tree_add_7_25_groupi_g17796(csa_tree_add_7_25_groupi_n_3294 ,csa_tree_add_7_25_groupi_n_387 ,csa_tree_add_7_25_groupi_n_1613);
  nor csa_tree_add_7_25_groupi_g17797(csa_tree_add_7_25_groupi_n_3293 ,csa_tree_add_7_25_groupi_n_819 ,csa_tree_add_7_25_groupi_n_1316);
  nor csa_tree_add_7_25_groupi_g17798(csa_tree_add_7_25_groupi_n_3292 ,csa_tree_add_7_25_groupi_n_726 ,csa_tree_add_7_25_groupi_n_129);
  nor csa_tree_add_7_25_groupi_g17799(csa_tree_add_7_25_groupi_n_3291 ,csa_tree_add_7_25_groupi_n_759 ,csa_tree_add_7_25_groupi_n_1849);
  nor csa_tree_add_7_25_groupi_g17800(csa_tree_add_7_25_groupi_n_3290 ,csa_tree_add_7_25_groupi_n_813 ,csa_tree_add_7_25_groupi_n_1307);
  nor csa_tree_add_7_25_groupi_g17801(csa_tree_add_7_25_groupi_n_3289 ,csa_tree_add_7_25_groupi_n_717 ,csa_tree_add_7_25_groupi_n_183);
  nor csa_tree_add_7_25_groupi_g17802(csa_tree_add_7_25_groupi_n_3288 ,csa_tree_add_7_25_groupi_n_783 ,csa_tree_add_7_25_groupi_n_1848);
  nor csa_tree_add_7_25_groupi_g17803(csa_tree_add_7_25_groupi_n_3287 ,csa_tree_add_7_25_groupi_n_807 ,csa_tree_add_7_25_groupi_n_183);
  nor csa_tree_add_7_25_groupi_g17804(csa_tree_add_7_25_groupi_n_3286 ,csa_tree_add_7_25_groupi_n_891 ,csa_tree_add_7_25_groupi_n_1307);
  nor csa_tree_add_7_25_groupi_g17805(csa_tree_add_7_25_groupi_n_3285 ,csa_tree_add_7_25_groupi_n_798 ,csa_tree_add_7_25_groupi_n_122);
  nor csa_tree_add_7_25_groupi_g17806(csa_tree_add_7_25_groupi_n_3284 ,csa_tree_add_7_25_groupi_n_747 ,csa_tree_add_7_25_groupi_n_1315);
  nor csa_tree_add_7_25_groupi_g17807(csa_tree_add_7_25_groupi_n_3283 ,csa_tree_add_7_25_groupi_n_876 ,csa_tree_add_7_25_groupi_n_1316);
  nor csa_tree_add_7_25_groupi_g17808(csa_tree_add_7_25_groupi_n_3282 ,csa_tree_add_7_25_groupi_n_861 ,csa_tree_add_7_25_groupi_n_1315);
  nor csa_tree_add_7_25_groupi_g17809(csa_tree_add_7_25_groupi_n_3281 ,csa_tree_add_7_25_groupi_n_414 ,csa_tree_add_7_25_groupi_n_1681);
  nor csa_tree_add_7_25_groupi_g17810(csa_tree_add_7_25_groupi_n_3280 ,csa_tree_add_7_25_groupi_n_420 ,csa_tree_add_7_25_groupi_n_1414);
  nor csa_tree_add_7_25_groupi_g17811(csa_tree_add_7_25_groupi_n_3279 ,csa_tree_add_7_25_groupi_n_385 ,csa_tree_add_7_25_groupi_n_1718);
  nor csa_tree_add_7_25_groupi_g17812(csa_tree_add_7_25_groupi_n_3278 ,csa_tree_add_7_25_groupi_n_351 ,csa_tree_add_7_25_groupi_n_1435);
  nor csa_tree_add_7_25_groupi_g17813(csa_tree_add_7_25_groupi_n_3277 ,csa_tree_add_7_25_groupi_n_430 ,csa_tree_add_7_25_groupi_n_1450);
  nor csa_tree_add_7_25_groupi_g17814(csa_tree_add_7_25_groupi_n_3276 ,csa_tree_add_7_25_groupi_n_412 ,csa_tree_add_7_25_groupi_n_1519);
  nor csa_tree_add_7_25_groupi_g17815(csa_tree_add_7_25_groupi_n_3275 ,csa_tree_add_7_25_groupi_n_558 ,csa_tree_add_7_25_groupi_n_1769);
  nor csa_tree_add_7_25_groupi_g17816(csa_tree_add_7_25_groupi_n_3274 ,csa_tree_add_7_25_groupi_n_561 ,csa_tree_add_7_25_groupi_n_1711);
  nor csa_tree_add_7_25_groupi_g17817(csa_tree_add_7_25_groupi_n_3273 ,csa_tree_add_7_25_groupi_n_1045 ,csa_tree_add_7_25_groupi_n_1304);
  nor csa_tree_add_7_25_groupi_g17818(csa_tree_add_7_25_groupi_n_3272 ,csa_tree_add_7_25_groupi_n_965 ,csa_tree_add_7_25_groupi_n_1303);
  nor csa_tree_add_7_25_groupi_g17819(csa_tree_add_7_25_groupi_n_3271 ,csa_tree_add_7_25_groupi_n_1048 ,csa_tree_add_7_25_groupi_n_1628);
  nor csa_tree_add_7_25_groupi_g17820(csa_tree_add_7_25_groupi_n_3270 ,csa_tree_add_7_25_groupi_n_834 ,csa_tree_add_7_25_groupi_n_1324);
  nor csa_tree_add_7_25_groupi_g17821(csa_tree_add_7_25_groupi_n_3269 ,csa_tree_add_7_25_groupi_n_840 ,csa_tree_add_7_25_groupi_n_1646);
  nor csa_tree_add_7_25_groupi_g17822(csa_tree_add_7_25_groupi_n_3268 ,csa_tree_add_7_25_groupi_n_666 ,csa_tree_add_7_25_groupi_n_1748);
  nor csa_tree_add_7_25_groupi_g17823(csa_tree_add_7_25_groupi_n_3267 ,csa_tree_add_7_25_groupi_n_846 ,csa_tree_add_7_25_groupi_n_1790);
  nor csa_tree_add_7_25_groupi_g17824(csa_tree_add_7_25_groupi_n_3266 ,csa_tree_add_7_25_groupi_n_426 ,csa_tree_add_7_25_groupi_n_1622);
  nor csa_tree_add_7_25_groupi_g17825(csa_tree_add_7_25_groupi_n_3265 ,csa_tree_add_7_25_groupi_n_432 ,csa_tree_add_7_25_groupi_n_1609);
  nor csa_tree_add_7_25_groupi_g17826(csa_tree_add_7_25_groupi_n_3264 ,csa_tree_add_7_25_groupi_n_599 ,csa_tree_add_7_25_groupi_n_1618);
  nor csa_tree_add_7_25_groupi_g17827(csa_tree_add_7_25_groupi_n_3263 ,csa_tree_add_7_25_groupi_n_1036 ,csa_tree_add_7_25_groupi_n_152);
  nor csa_tree_add_7_25_groupi_g17828(csa_tree_add_7_25_groupi_n_3262 ,csa_tree_add_7_25_groupi_n_342 ,csa_tree_add_7_25_groupi_n_1507);
  nor csa_tree_add_7_25_groupi_g17829(csa_tree_add_7_25_groupi_n_3261 ,csa_tree_add_7_25_groupi_n_761 ,csa_tree_add_7_25_groupi_n_1711);
  nor csa_tree_add_7_25_groupi_g17830(csa_tree_add_7_25_groupi_n_3260 ,csa_tree_add_7_25_groupi_n_418 ,csa_tree_add_7_25_groupi_n_1531);
  nor csa_tree_add_7_25_groupi_g17831(csa_tree_add_7_25_groupi_n_3259 ,csa_tree_add_7_25_groupi_n_564 ,csa_tree_add_7_25_groupi_n_1735);
  nor csa_tree_add_7_25_groupi_g17832(csa_tree_add_7_25_groupi_n_3258 ,csa_tree_add_7_25_groupi_n_567 ,csa_tree_add_7_25_groupi_n_1424);
  nor csa_tree_add_7_25_groupi_g17833(csa_tree_add_7_25_groupi_n_3257 ,csa_tree_add_7_25_groupi_n_400 ,csa_tree_add_7_25_groupi_n_1444);
  nor csa_tree_add_7_25_groupi_g17834(csa_tree_add_7_25_groupi_n_3256 ,csa_tree_add_7_25_groupi_n_354 ,csa_tree_add_7_25_groupi_n_1672);
  nor csa_tree_add_7_25_groupi_g17835(csa_tree_add_7_25_groupi_n_3255 ,csa_tree_add_7_25_groupi_n_345 ,csa_tree_add_7_25_groupi_n_1765);
  nor csa_tree_add_7_25_groupi_g17836(csa_tree_add_7_25_groupi_n_3254 ,csa_tree_add_7_25_groupi_n_651 ,csa_tree_add_7_25_groupi_n_1660);
  nor csa_tree_add_7_25_groupi_g17837(csa_tree_add_7_25_groupi_n_3253 ,csa_tree_add_7_25_groupi_n_687 ,csa_tree_add_7_25_groupi_n_1721);
  nor csa_tree_add_7_25_groupi_g17838(csa_tree_add_7_25_groupi_n_3252 ,csa_tree_add_7_25_groupi_n_962 ,csa_tree_add_7_25_groupi_n_1799);
  nor csa_tree_add_7_25_groupi_g17839(csa_tree_add_7_25_groupi_n_3251 ,csa_tree_add_7_25_groupi_n_435 ,csa_tree_add_7_25_groupi_n_1640);
  nor csa_tree_add_7_25_groupi_g17840(csa_tree_add_7_25_groupi_n_3250 ,csa_tree_add_7_25_groupi_n_852 ,csa_tree_add_7_25_groupi_n_1792);
  nor csa_tree_add_7_25_groupi_g17841(csa_tree_add_7_25_groupi_n_3249 ,csa_tree_add_7_25_groupi_n_651 ,csa_tree_add_7_25_groupi_n_1600);
  nor csa_tree_add_7_25_groupi_g17842(csa_tree_add_7_25_groupi_n_3248 ,csa_tree_add_7_25_groupi_n_605 ,csa_tree_add_7_25_groupi_n_1390);
  nor csa_tree_add_7_25_groupi_g17843(csa_tree_add_7_25_groupi_n_3247 ,csa_tree_add_7_25_groupi_n_647 ,csa_tree_add_7_25_groupi_n_1357);
  nor csa_tree_add_7_25_groupi_g17844(csa_tree_add_7_25_groupi_n_3246 ,csa_tree_add_7_25_groupi_n_882 ,csa_tree_add_7_25_groupi_n_1313);
  nor csa_tree_add_7_25_groupi_g17845(csa_tree_add_7_25_groupi_n_3245 ,csa_tree_add_7_25_groupi_n_816 ,csa_tree_add_7_25_groupi_n_200);
  nor csa_tree_add_7_25_groupi_g17846(csa_tree_add_7_25_groupi_n_3244 ,csa_tree_add_7_25_groupi_n_900 ,csa_tree_add_7_25_groupi_n_1312);
  nor csa_tree_add_7_25_groupi_g17847(csa_tree_add_7_25_groupi_n_3243 ,csa_tree_add_7_25_groupi_n_804 ,csa_tree_add_7_25_groupi_n_507);
  nor csa_tree_add_7_25_groupi_g17848(csa_tree_add_7_25_groupi_n_3242 ,csa_tree_add_7_25_groupi_n_663 ,csa_tree_add_7_25_groupi_n_525);
  nor csa_tree_add_7_25_groupi_g17849(csa_tree_add_7_25_groupi_n_3241 ,csa_tree_add_7_25_groupi_n_810 ,csa_tree_add_7_25_groupi_n_525);
  nor csa_tree_add_7_25_groupi_g17850(csa_tree_add_7_25_groupi_n_3240 ,csa_tree_add_7_25_groupi_n_855 ,csa_tree_add_7_25_groupi_n_507);
  nor csa_tree_add_7_25_groupi_g17851(csa_tree_add_7_25_groupi_n_3239 ,csa_tree_add_7_25_groupi_n_681 ,csa_tree_add_7_25_groupi_n_1304);
  nor csa_tree_add_7_25_groupi_g17852(csa_tree_add_7_25_groupi_n_3238 ,csa_tree_add_7_25_groupi_n_729 ,csa_tree_add_7_25_groupi_n_200);
  nor csa_tree_add_7_25_groupi_g17853(csa_tree_add_7_25_groupi_n_3237 ,csa_tree_add_7_25_groupi_n_858 ,csa_tree_add_7_25_groupi_n_1312);
  nor csa_tree_add_7_25_groupi_g17854(csa_tree_add_7_25_groupi_n_3236 ,csa_tree_add_7_25_groupi_n_927 ,csa_tree_add_7_25_groupi_n_152);
  nor csa_tree_add_7_25_groupi_g17855(csa_tree_add_7_25_groupi_n_3235 ,csa_tree_add_7_25_groupi_n_843 ,csa_tree_add_7_25_groupi_n_506);
  nor csa_tree_add_7_25_groupi_g17856(csa_tree_add_7_25_groupi_n_3234 ,csa_tree_add_7_25_groupi_n_827 ,csa_tree_add_7_25_groupi_n_1324);
  nor csa_tree_add_7_25_groupi_g17857(csa_tree_add_7_25_groupi_n_3233 ,csa_tree_add_7_25_groupi_n_974 ,csa_tree_add_7_25_groupi_n_1747);
  nor csa_tree_add_7_25_groupi_g17858(csa_tree_add_7_25_groupi_n_3232 ,csa_tree_add_7_25_groupi_n_660 ,csa_tree_add_7_25_groupi_n_1651);
  nor csa_tree_add_7_25_groupi_g17859(csa_tree_add_7_25_groupi_n_3231 ,csa_tree_add_7_25_groupi_n_696 ,csa_tree_add_7_25_groupi_n_1331);
  nor csa_tree_add_7_25_groupi_g17860(csa_tree_add_7_25_groupi_n_3230 ,csa_tree_add_7_25_groupi_n_933 ,csa_tree_add_7_25_groupi_n_1998);
  nor csa_tree_add_7_25_groupi_g17861(csa_tree_add_7_25_groupi_n_3229 ,csa_tree_add_7_25_groupi_n_405 ,csa_tree_add_7_25_groupi_n_1682);
  nor csa_tree_add_7_25_groupi_g17862(csa_tree_add_7_25_groupi_n_3228 ,csa_tree_add_7_25_groupi_n_394 ,csa_tree_add_7_25_groupi_n_522);
  nor csa_tree_add_7_25_groupi_g17863(csa_tree_add_7_25_groupi_n_3227 ,csa_tree_add_7_25_groupi_n_360 ,csa_tree_add_7_25_groupi_n_1415);
  nor csa_tree_add_7_25_groupi_g17864(csa_tree_add_7_25_groupi_n_3226 ,csa_tree_add_7_25_groupi_n_764 ,csa_tree_add_7_25_groupi_n_1346);
  nor csa_tree_add_7_25_groupi_g17865(csa_tree_add_7_25_groupi_n_3225 ,csa_tree_add_7_25_groupi_n_767 ,csa_tree_add_7_25_groupi_n_1741);
  nor csa_tree_add_7_25_groupi_g17866(csa_tree_add_7_25_groupi_n_3224 ,csa_tree_add_7_25_groupi_n_570 ,csa_tree_add_7_25_groupi_n_1451);
  nor csa_tree_add_7_25_groupi_g17867(csa_tree_add_7_25_groupi_n_3223 ,csa_tree_add_7_25_groupi_n_573 ,csa_tree_add_7_25_groupi_n_1718);
  nor csa_tree_add_7_25_groupi_g17868(csa_tree_add_7_25_groupi_n_3222 ,csa_tree_add_7_25_groupi_n_403 ,csa_tree_add_7_25_groupi_n_1436);
  nor csa_tree_add_7_25_groupi_g17869(csa_tree_add_7_25_groupi_n_3221 ,csa_tree_add_7_25_groupi_n_406 ,csa_tree_add_7_25_groupi_n_1328);
  nor csa_tree_add_7_25_groupi_g17870(csa_tree_add_7_25_groupi_n_3220 ,csa_tree_add_7_25_groupi_n_669 ,csa_tree_add_7_25_groupi_n_1630);
  nor csa_tree_add_7_25_groupi_g17871(csa_tree_add_7_25_groupi_n_3219 ,csa_tree_add_7_25_groupi_n_608 ,csa_tree_add_7_25_groupi_n_1402);
  nor csa_tree_add_7_25_groupi_g17872(csa_tree_add_7_25_groupi_n_3218 ,csa_tree_add_7_25_groupi_n_596 ,csa_tree_add_7_25_groupi_n_1405);
  nor csa_tree_add_7_25_groupi_g17873(csa_tree_add_7_25_groupi_n_3217 ,csa_tree_add_7_25_groupi_n_864 ,csa_tree_add_7_25_groupi_n_1411);
  nor csa_tree_add_7_25_groupi_g17874(csa_tree_add_7_25_groupi_n_3216 ,csa_tree_add_7_25_groupi_n_918 ,csa_tree_add_7_25_groupi_n_1759);
  nor csa_tree_add_7_25_groupi_g17875(csa_tree_add_7_25_groupi_n_3215 ,csa_tree_add_7_25_groupi_n_1006 ,csa_tree_add_7_25_groupi_n_1720);
  nor csa_tree_add_7_25_groupi_g17876(csa_tree_add_7_25_groupi_n_3214 ,csa_tree_add_7_25_groupi_n_921 ,csa_tree_add_7_25_groupi_n_1753);
  nor csa_tree_add_7_25_groupi_g17877(csa_tree_add_7_25_groupi_n_3213 ,csa_tree_add_7_25_groupi_n_885 ,csa_tree_add_7_25_groupi_n_1750);
  nor csa_tree_add_7_25_groupi_g17878(csa_tree_add_7_25_groupi_n_3212 ,csa_tree_add_7_25_groupi_n_1027 ,csa_tree_add_7_25_groupi_n_1754);
  nor csa_tree_add_7_25_groupi_g17879(csa_tree_add_7_25_groupi_n_3211 ,csa_tree_add_7_25_groupi_n_720 ,csa_tree_add_7_25_groupi_n_1759);
  nor csa_tree_add_7_25_groupi_g17880(csa_tree_add_7_25_groupi_n_3210 ,csa_tree_add_7_25_groupi_n_903 ,csa_tree_add_7_25_groupi_n_1798);
  nor csa_tree_add_7_25_groupi_g17881(csa_tree_add_7_25_groupi_n_3209 ,csa_tree_add_7_25_groupi_n_738 ,csa_tree_add_7_25_groupi_n_1751);
  nor csa_tree_add_7_25_groupi_g17882(csa_tree_add_7_25_groupi_n_3208 ,csa_tree_add_7_25_groupi_n_870 ,csa_tree_add_7_25_groupi_n_1753);
  nor csa_tree_add_7_25_groupi_g17883(csa_tree_add_7_25_groupi_n_3207 ,csa_tree_add_7_25_groupi_n_912 ,csa_tree_add_7_25_groupi_n_1748);
  nor csa_tree_add_7_25_groupi_g17884(csa_tree_add_7_25_groupi_n_3206 ,csa_tree_add_7_25_groupi_n_675 ,csa_tree_add_7_25_groupi_n_1754);
  nor csa_tree_add_7_25_groupi_g17885(csa_tree_add_7_25_groupi_n_3205 ,csa_tree_add_7_25_groupi_n_894 ,csa_tree_add_7_25_groupi_n_1798);
  nor csa_tree_add_7_25_groupi_g17886(csa_tree_add_7_25_groupi_n_3204 ,csa_tree_add_7_25_groupi_n_776 ,csa_tree_add_7_25_groupi_n_1664);
  nor csa_tree_add_7_25_groupi_g17887(csa_tree_add_7_25_groupi_n_3203 ,csa_tree_add_7_25_groupi_n_830 ,csa_tree_add_7_25_groupi_n_1238);
  nor csa_tree_add_7_25_groupi_g17888(csa_tree_add_7_25_groupi_n_3202 ,csa_tree_add_7_25_groupi_n_621 ,csa_tree_add_7_25_groupi_n_1998);
  nor csa_tree_add_7_25_groupi_g17889(csa_tree_add_7_25_groupi_n_3201 ,csa_tree_add_7_25_groupi_n_791 ,csa_tree_add_7_25_groupi_n_1363);
  nor csa_tree_add_7_25_groupi_g17890(csa_tree_add_7_25_groupi_n_3200 ,csa_tree_add_7_25_groupi_n_683 ,csa_tree_add_7_25_groupi_n_1372);
  and csa_tree_add_7_25_groupi_g17891(csa_tree_add_7_25_groupi_n_3535 ,csa_tree_add_7_25_groupi_n_2822 ,csa_tree_add_7_25_groupi_n_2805);
  or csa_tree_add_7_25_groupi_g17892(csa_tree_add_7_25_groupi_n_3532 ,csa_tree_add_7_25_groupi_n_2810 ,csa_tree_add_7_25_groupi_n_2814);
  or csa_tree_add_7_25_groupi_g17893(csa_tree_add_7_25_groupi_n_3528 ,csa_tree_add_7_25_groupi_n_2834 ,csa_tree_add_7_25_groupi_n_2816);
  or csa_tree_add_7_25_groupi_g17894(csa_tree_add_7_25_groupi_n_3526 ,csa_tree_add_7_25_groupi_n_2823 ,csa_tree_add_7_25_groupi_n_2833);
  or csa_tree_add_7_25_groupi_g17895(csa_tree_add_7_25_groupi_n_3521 ,csa_tree_add_7_25_groupi_n_2812 ,csa_tree_add_7_25_groupi_n_2826);
  or csa_tree_add_7_25_groupi_g17896(csa_tree_add_7_25_groupi_n_3516 ,csa_tree_add_7_25_groupi_n_2825 ,csa_tree_add_7_25_groupi_n_2829);
  or csa_tree_add_7_25_groupi_g17897(csa_tree_add_7_25_groupi_n_3511 ,csa_tree_add_7_25_groupi_n_2806 ,csa_tree_add_7_25_groupi_n_2818);
  or csa_tree_add_7_25_groupi_g17898(csa_tree_add_7_25_groupi_n_3506 ,csa_tree_add_7_25_groupi_n_2821 ,csa_tree_add_7_25_groupi_n_2835);
  or csa_tree_add_7_25_groupi_g17899(csa_tree_add_7_25_groupi_n_3501 ,csa_tree_add_7_25_groupi_n_2828 ,csa_tree_add_7_25_groupi_n_2809);
  nor csa_tree_add_7_25_groupi_g17900(csa_tree_add_7_25_groupi_n_3198 ,csa_tree_add_7_25_groupi_n_1069 ,csa_tree_add_7_25_groupi_n_1520);
  nor csa_tree_add_7_25_groupi_g17901(csa_tree_add_7_25_groupi_n_3197 ,csa_tree_add_7_25_groupi_n_474 ,csa_tree_add_7_25_groupi_n_2003);
  nor csa_tree_add_7_25_groupi_g17902(csa_tree_add_7_25_groupi_n_3196 ,csa_tree_add_7_25_groupi_n_590 ,csa_tree_add_7_25_groupi_n_1333);
  nor csa_tree_add_7_25_groupi_g17903(csa_tree_add_7_25_groupi_n_3195 ,csa_tree_add_7_25_groupi_n_938 ,csa_tree_add_7_25_groupi_n_1349);
  nor csa_tree_add_7_25_groupi_g17904(csa_tree_add_7_25_groupi_n_3194 ,csa_tree_add_7_25_groupi_n_770 ,csa_tree_add_7_25_groupi_n_1355);
  nor csa_tree_add_7_25_groupi_g17905(csa_tree_add_7_25_groupi_n_3193 ,csa_tree_add_7_25_groupi_n_773 ,csa_tree_add_7_25_groupi_n_1427);
  nor csa_tree_add_7_25_groupi_g17906(csa_tree_add_7_25_groupi_n_3192 ,csa_tree_add_7_25_groupi_n_779 ,csa_tree_add_7_25_groupi_n_1445);
  nor csa_tree_add_7_25_groupi_g17907(csa_tree_add_7_25_groupi_n_3191 ,csa_tree_add_7_25_groupi_n_542 ,csa_tree_add_7_25_groupi_n_1508);
  nor csa_tree_add_7_25_groupi_g17908(csa_tree_add_7_25_groupi_n_3190 ,csa_tree_add_7_25_groupi_n_588 ,csa_tree_add_7_25_groupi_n_1763);
  nor csa_tree_add_7_25_groupi_g17909(csa_tree_add_7_25_groupi_n_3189 ,csa_tree_add_7_25_groupi_n_472 ,csa_tree_add_7_25_groupi_n_1685);
  nor csa_tree_add_7_25_groupi_g17910(csa_tree_add_7_25_groupi_n_3188 ,csa_tree_add_7_25_groupi_n_545 ,csa_tree_add_7_25_groupi_n_1298);
  nor csa_tree_add_7_25_groupi_g17911(csa_tree_add_7_25_groupi_n_3187 ,csa_tree_add_7_25_groupi_n_575 ,csa_tree_add_7_25_groupi_n_1345);
  nor csa_tree_add_7_25_groupi_g17912(csa_tree_add_7_25_groupi_n_3186 ,csa_tree_add_7_25_groupi_n_578 ,csa_tree_add_7_25_groupi_n_516);
  nor csa_tree_add_7_25_groupi_g17913(csa_tree_add_7_25_groupi_n_3185 ,csa_tree_add_7_25_groupi_n_388 ,csa_tree_add_7_25_groupi_n_1739);
  nor csa_tree_add_7_25_groupi_g17914(csa_tree_add_7_25_groupi_n_3184 ,csa_tree_add_7_25_groupi_n_582 ,csa_tree_add_7_25_groupi_n_1532);
  nor csa_tree_add_7_25_groupi_g17915(csa_tree_add_7_25_groupi_n_3183 ,csa_tree_add_7_25_groupi_n_585 ,csa_tree_add_7_25_groupi_n_1739);
  nor csa_tree_add_7_25_groupi_g17916(csa_tree_add_7_25_groupi_n_3182 ,csa_tree_add_7_25_groupi_n_705 ,csa_tree_add_7_25_groupi_n_1351);
  nor csa_tree_add_7_25_groupi_g17917(csa_tree_add_7_25_groupi_n_3181 ,csa_tree_add_7_25_groupi_n_1081 ,csa_tree_add_7_25_groupi_n_2015);
  nor csa_tree_add_7_25_groupi_g17918(csa_tree_add_7_25_groupi_n_3180 ,csa_tree_add_7_25_groupi_n_1012 ,csa_tree_add_7_25_groupi_n_2013);
  nor csa_tree_add_7_25_groupi_g17919(csa_tree_add_7_25_groupi_n_3179 ,csa_tree_add_7_25_groupi_n_711 ,csa_tree_add_7_25_groupi_n_2013);
  nor csa_tree_add_7_25_groupi_g17920(csa_tree_add_7_25_groupi_n_3178 ,csa_tree_add_7_25_groupi_n_1009 ,csa_tree_add_7_25_groupi_n_1792);
  nor csa_tree_add_7_25_groupi_g17921(csa_tree_add_7_25_groupi_n_3177 ,csa_tree_add_7_25_groupi_n_1015 ,csa_tree_add_7_25_groupi_n_1336);
  nor csa_tree_add_7_25_groupi_g17922(csa_tree_add_7_25_groupi_n_3176 ,csa_tree_add_7_25_groupi_n_1072 ,csa_tree_add_7_25_groupi_n_1790);
  nor csa_tree_add_7_25_groupi_g17923(csa_tree_add_7_25_groupi_n_3175 ,csa_tree_add_7_25_groupi_n_1018 ,csa_tree_add_7_25_groupi_n_2016);
  nor csa_tree_add_7_25_groupi_g17924(csa_tree_add_7_25_groupi_n_3174 ,csa_tree_add_7_25_groupi_n_1039 ,csa_tree_add_7_25_groupi_n_2012);
  nor csa_tree_add_7_25_groupi_g17925(csa_tree_add_7_25_groupi_n_3173 ,csa_tree_add_7_25_groupi_n_1030 ,csa_tree_add_7_25_groupi_n_1789);
  nor csa_tree_add_7_25_groupi_g17926(csa_tree_add_7_25_groupi_n_3172 ,csa_tree_add_7_25_groupi_n_1087 ,csa_tree_add_7_25_groupi_n_1331);
  nor csa_tree_add_7_25_groupi_g17927(csa_tree_add_7_25_groupi_n_3171 ,csa_tree_add_7_25_groupi_n_1075 ,csa_tree_add_7_25_groupi_n_2012);
  nor csa_tree_add_7_25_groupi_g17928(csa_tree_add_7_25_groupi_n_3170 ,csa_tree_add_7_25_groupi_n_1057 ,csa_tree_add_7_25_groupi_n_1336);
  nor csa_tree_add_7_25_groupi_g17929(csa_tree_add_7_25_groupi_n_3169 ,csa_tree_add_7_25_groupi_n_755 ,csa_tree_add_7_25_groupi_n_1244);
  nor csa_tree_add_7_25_groupi_g17930(csa_tree_add_7_25_groupi_n_3168 ,csa_tree_add_7_25_groupi_n_866 ,csa_tree_add_7_25_groupi_n_1229);
  nor csa_tree_add_7_25_groupi_g17931(csa_tree_add_7_25_groupi_n_3167 ,csa_tree_add_7_25_groupi_n_878 ,csa_tree_add_7_25_groupi_n_1235);
  nor csa_tree_add_7_25_groupi_g17932(csa_tree_add_7_25_groupi_n_3166 ,csa_tree_add_7_25_groupi_n_701 ,csa_tree_add_7_25_groupi_n_1241);
  nor csa_tree_add_7_25_groupi_g17933(csa_tree_add_7_25_groupi_n_3165 ,csa_tree_add_7_25_groupi_n_602 ,csa_tree_add_7_25_groupi_n_1673);
  nor csa_tree_add_7_25_groupi_g17934(csa_tree_add_7_25_groupi_n_3164 ,csa_tree_add_7_25_groupi_n_785 ,csa_tree_add_7_25_groupi_n_1327);
  nor csa_tree_add_7_25_groupi_g17935(csa_tree_add_7_25_groupi_n_3163 ,csa_tree_add_7_25_groupi_n_788 ,csa_tree_add_7_25_groupi_n_1549);
  nor csa_tree_add_7_25_groupi_g17936(csa_tree_add_7_25_groupi_n_3162 ,csa_tree_add_7_25_groupi_n_833 ,csa_tree_add_7_25_groupi_n_1730);
  nor csa_tree_add_7_25_groupi_g17937(csa_tree_add_7_25_groupi_n_3161 ,csa_tree_add_7_25_groupi_n_839 ,csa_tree_add_7_25_groupi_n_1675);
  nor csa_tree_add_7_25_groupi_g17938(csa_tree_add_7_25_groupi_n_3160 ,csa_tree_add_7_25_groupi_n_427 ,csa_tree_add_7_25_groupi_n_1375);
  nor csa_tree_add_7_25_groupi_g17939(csa_tree_add_7_25_groupi_n_3159 ,csa_tree_add_7_25_groupi_n_433 ,csa_tree_add_7_25_groupi_n_1345);
  nor csa_tree_add_7_25_groupi_g17940(csa_tree_add_7_25_groupi_n_3158 ,csa_tree_add_7_25_groupi_n_600 ,csa_tree_add_7_25_groupi_n_1911);
  nor csa_tree_add_7_25_groupi_g17941(csa_tree_add_7_25_groupi_n_3157 ,csa_tree_add_7_25_groupi_n_603 ,csa_tree_add_7_25_groupi_n_1756);
  nor csa_tree_add_7_25_groupi_g17942(csa_tree_add_7_25_groupi_n_3156 ,csa_tree_add_7_25_groupi_n_1051 ,csa_tree_add_7_25_groupi_n_1239);
  nor csa_tree_add_7_25_groupi_g17943(csa_tree_add_7_25_groupi_n_3155 ,csa_tree_add_7_25_groupi_n_1024 ,csa_tree_add_7_25_groupi_n_1147);
  nor csa_tree_add_7_25_groupi_g17944(csa_tree_add_7_25_groupi_n_3154 ,csa_tree_add_7_25_groupi_n_1063 ,csa_tree_add_7_25_groupi_n_1660);
  nor csa_tree_add_7_25_groupi_g17945(csa_tree_add_7_25_groupi_n_3153 ,csa_tree_add_7_25_groupi_n_1054 ,csa_tree_add_7_25_groupi_n_1352);
  nor csa_tree_add_7_25_groupi_g17946(csa_tree_add_7_25_groupi_n_3152 ,csa_tree_add_7_25_groupi_n_1042 ,csa_tree_add_7_25_groupi_n_1658);
  nor csa_tree_add_7_25_groupi_g17947(csa_tree_add_7_25_groupi_n_3151 ,csa_tree_add_7_25_groupi_n_1066 ,csa_tree_add_7_25_groupi_n_1148);
  nor csa_tree_add_7_25_groupi_g17948(csa_tree_add_7_25_groupi_n_3150 ,csa_tree_add_7_25_groupi_n_1078 ,csa_tree_add_7_25_groupi_n_1654);
  nor csa_tree_add_7_25_groupi_g17949(csa_tree_add_7_25_groupi_n_3149 ,csa_tree_add_7_25_groupi_n_1060 ,csa_tree_add_7_25_groupi_n_1351);
  nor csa_tree_add_7_25_groupi_g17950(csa_tree_add_7_25_groupi_n_3148 ,csa_tree_add_7_25_groupi_n_732 ,csa_tree_add_7_25_groupi_n_1658);
  nor csa_tree_add_7_25_groupi_g17951(csa_tree_add_7_25_groupi_n_3147 ,csa_tree_add_7_25_groupi_n_1084 ,csa_tree_add_7_25_groupi_n_1664);
  nor csa_tree_add_7_25_groupi_g17952(csa_tree_add_7_25_groupi_n_3146 ,csa_tree_add_7_25_groupi_n_1033 ,csa_tree_add_7_25_groupi_n_1654);
  nor csa_tree_add_7_25_groupi_g17953(csa_tree_add_7_25_groupi_n_3145 ,csa_tree_add_7_25_groupi_n_1021 ,csa_tree_add_7_25_groupi_n_1655);
  nor csa_tree_add_7_25_groupi_g17954(csa_tree_add_7_25_groupi_n_3144 ,csa_tree_add_7_25_groupi_n_971 ,csa_tree_add_7_25_groupi_n_1652);
  nor csa_tree_add_7_25_groupi_g17955(csa_tree_add_7_25_groupi_n_3143 ,csa_tree_add_7_25_groupi_n_977 ,csa_tree_add_7_25_groupi_n_1640);
  nor csa_tree_add_7_25_groupi_g17956(csa_tree_add_7_25_groupi_n_3142 ,csa_tree_add_7_25_groupi_n_953 ,csa_tree_add_7_25_groupi_n_1373);
  nor csa_tree_add_7_25_groupi_g17957(csa_tree_add_7_25_groupi_n_3141 ,csa_tree_add_7_25_groupi_n_986 ,csa_tree_add_7_25_groupi_n_1363);
  nor csa_tree_add_7_25_groupi_g17958(csa_tree_add_7_25_groupi_n_3140 ,csa_tree_add_7_25_groupi_n_968 ,csa_tree_add_7_25_groupi_n_1646);
  nor csa_tree_add_7_25_groupi_g17959(csa_tree_add_7_25_groupi_n_3139 ,csa_tree_add_7_25_groupi_n_980 ,csa_tree_add_7_25_groupi_n_1642);
  nor csa_tree_add_7_25_groupi_g17960(csa_tree_add_7_25_groupi_n_3138 ,csa_tree_add_7_25_groupi_n_959 ,csa_tree_add_7_25_groupi_n_1649);
  nor csa_tree_add_7_25_groupi_g17961(csa_tree_add_7_25_groupi_n_3137 ,csa_tree_add_7_25_groupi_n_734 ,csa_tree_add_7_25_groupi_n_1643);
  nor csa_tree_add_7_25_groupi_g17962(csa_tree_add_7_25_groupi_n_3136 ,csa_tree_add_7_25_groupi_n_944 ,csa_tree_add_7_25_groupi_n_1651);
  nor csa_tree_add_7_25_groupi_g17963(csa_tree_add_7_25_groupi_n_3135 ,csa_tree_add_7_25_groupi_n_615 ,csa_tree_add_7_25_groupi_n_1642);
  nor csa_tree_add_7_25_groupi_g17964(csa_tree_add_7_25_groupi_n_3134 ,csa_tree_add_7_25_groupi_n_956 ,csa_tree_add_7_25_groupi_n_1372);
  nor csa_tree_add_7_25_groupi_g17965(csa_tree_add_7_25_groupi_n_3133 ,csa_tree_add_7_25_groupi_n_947 ,csa_tree_add_7_25_groupi_n_1245);
  nor csa_tree_add_7_25_groupi_g17966(csa_tree_add_7_25_groupi_n_3132 ,csa_tree_add_7_25_groupi_n_897 ,csa_tree_add_7_25_groupi_n_1358);
  nor csa_tree_add_7_25_groupi_g17967(csa_tree_add_7_25_groupi_n_3131 ,csa_tree_add_7_25_groupi_n_887 ,csa_tree_add_7_25_groupi_n_1610);
  nor csa_tree_add_7_25_groupi_g17968(csa_tree_add_7_25_groupi_n_3130 ,csa_tree_add_7_25_groupi_n_678 ,csa_tree_add_7_25_groupi_n_1604);
  nor csa_tree_add_7_25_groupi_g17969(csa_tree_add_7_25_groupi_n_3129 ,csa_tree_add_7_25_groupi_n_906 ,csa_tree_add_7_25_groupi_n_1619);
  nor csa_tree_add_7_25_groupi_g17970(csa_tree_add_7_25_groupi_n_3128 ,csa_tree_add_7_25_groupi_n_723 ,csa_tree_add_7_25_groupi_n_1613);
  nor csa_tree_add_7_25_groupi_g17971(csa_tree_add_7_25_groupi_n_3127 ,csa_tree_add_7_25_groupi_n_744 ,csa_tree_add_7_25_groupi_n_1622);
  nor csa_tree_add_7_25_groupi_g17972(csa_tree_add_7_25_groupi_n_3126 ,csa_tree_add_7_25_groupi_n_872 ,csa_tree_add_7_25_groupi_n_1403);
  nor csa_tree_add_7_25_groupi_g17973(csa_tree_add_7_25_groupi_n_3125 ,csa_tree_add_7_25_groupi_n_749 ,csa_tree_add_7_25_groupi_n_1412);
  nor csa_tree_add_7_25_groupi_g17974(csa_tree_add_7_25_groupi_n_3124 ,csa_tree_add_7_25_groupi_n_983 ,csa_tree_add_7_25_groupi_n_1600);
  nor csa_tree_add_7_25_groupi_g17975(csa_tree_add_7_25_groupi_n_3123 ,csa_tree_add_7_25_groupi_n_797 ,csa_tree_add_7_25_groupi_n_1406);
  nor csa_tree_add_7_25_groupi_g17976(csa_tree_add_7_25_groupi_n_3122 ,csa_tree_add_7_25_groupi_n_653 ,csa_tree_add_7_25_groupi_n_1630);
  nor csa_tree_add_7_25_groupi_g17977(csa_tree_add_7_25_groupi_n_3121 ,csa_tree_add_7_25_groupi_n_689 ,csa_tree_add_7_25_groupi_n_1628);
  nor csa_tree_add_7_25_groupi_g17978(csa_tree_add_7_25_groupi_n_3120 ,csa_tree_add_7_25_groupi_n_908 ,csa_tree_add_7_25_groupi_n_1624);
  nor csa_tree_add_7_25_groupi_g17979(csa_tree_add_7_25_groupi_n_3119 ,csa_tree_add_7_25_groupi_n_848 ,csa_tree_add_7_25_groupi_n_1390);
  nor csa_tree_add_7_25_groupi_g17980(csa_tree_add_7_25_groupi_n_3118 ,csa_tree_add_7_25_groupi_n_924 ,csa_tree_add_7_25_groupi_n_1361);
  nor csa_tree_add_7_25_groupi_g17981(csa_tree_add_7_25_groupi_n_3117 ,csa_tree_add_7_25_groupi_n_824 ,csa_tree_add_7_25_groupi_n_1595);
  nor csa_tree_add_7_25_groupi_g17982(csa_tree_add_7_25_groupi_n_3116 ,csa_tree_add_7_25_groupi_n_800 ,csa_tree_add_7_25_groupi_n_1399);
  nor csa_tree_add_7_25_groupi_g17983(csa_tree_add_7_25_groupi_n_3115 ,csa_tree_add_7_25_groupi_n_806 ,csa_tree_add_7_25_groupi_n_1616);
  nor csa_tree_add_7_25_groupi_g17984(csa_tree_add_7_25_groupi_n_3114 ,csa_tree_add_7_25_groupi_n_812 ,csa_tree_add_7_25_groupi_n_1634);
  nor csa_tree_add_7_25_groupi_g17985(csa_tree_add_7_25_groupi_n_3113 ,csa_tree_add_7_25_groupi_n_818 ,csa_tree_add_7_25_groupi_n_1396);
  nor csa_tree_add_7_25_groupi_g17986(csa_tree_add_7_25_groupi_n_3112 ,csa_tree_add_7_25_groupi_n_671 ,csa_tree_add_7_25_groupi_n_1625);
  nor csa_tree_add_7_25_groupi_g17987(csa_tree_add_7_25_groupi_n_3111 ,csa_tree_add_7_25_groupi_n_836 ,csa_tree_add_7_25_groupi_n_1400);
  nor csa_tree_add_7_25_groupi_g17988(csa_tree_add_7_25_groupi_n_3110 ,csa_tree_add_7_25_groupi_n_860 ,csa_tree_add_7_25_groupi_n_1607);
  nor csa_tree_add_7_25_groupi_g17989(csa_tree_add_7_25_groupi_n_3109 ,csa_tree_add_7_25_groupi_n_707 ,csa_tree_add_7_25_groupi_n_1397);
  nor csa_tree_add_7_25_groupi_g17990(csa_tree_add_7_25_groupi_n_3108 ,csa_tree_add_7_25_groupi_n_714 ,csa_tree_add_7_25_groupi_n_1357);
  nor csa_tree_add_7_25_groupi_g17991(csa_tree_add_7_25_groupi_n_3107 ,csa_tree_add_7_25_groupi_n_915 ,csa_tree_add_7_25_groupi_n_1624);
  nor csa_tree_add_7_25_groupi_g17992(csa_tree_add_7_25_groupi_n_3106 ,csa_tree_add_7_25_groupi_n_875 ,csa_tree_add_7_25_groupi_n_1411);
  nor csa_tree_add_7_25_groupi_g17993(csa_tree_add_7_25_groupi_n_3105 ,csa_tree_add_7_25_groupi_n_752 ,csa_tree_add_7_25_groupi_n_1609);
  nor csa_tree_add_7_25_groupi_g17994(csa_tree_add_7_25_groupi_n_3104 ,csa_tree_add_7_25_groupi_n_698 ,csa_tree_add_7_25_groupi_n_1618);
  nor csa_tree_add_7_25_groupi_g17995(csa_tree_add_7_25_groupi_n_3103 ,csa_tree_add_7_25_groupi_n_716 ,csa_tree_add_7_25_groupi_n_1396);
  nor csa_tree_add_7_25_groupi_g17996(csa_tree_add_7_25_groupi_n_3102 ,csa_tree_add_7_25_groupi_n_746 ,csa_tree_add_7_25_groupi_n_1399);
  nor csa_tree_add_7_25_groupi_g17997(csa_tree_add_7_25_groupi_n_3101 ,csa_tree_add_7_25_groupi_n_782 ,csa_tree_add_7_25_groupi_n_1405);
  nor csa_tree_add_7_25_groupi_g17998(csa_tree_add_7_25_groupi_n_3100 ,csa_tree_add_7_25_groupi_n_758 ,csa_tree_add_7_25_groupi_n_1230);
  nor csa_tree_add_7_25_groupi_g17999(csa_tree_add_7_25_groupi_n_3099 ,csa_tree_add_7_25_groupi_n_890 ,csa_tree_add_7_25_groupi_n_1402);
  nor csa_tree_add_7_25_groupi_g18000(csa_tree_add_7_25_groupi_n_3098 ,csa_tree_add_7_25_groupi_n_725 ,csa_tree_add_7_25_groupi_n_1242);
  nor csa_tree_add_7_25_groupi_g18001(csa_tree_add_7_25_groupi_n_3097 ,csa_tree_add_7_25_groupi_n_728 ,csa_tree_add_7_25_groupi_n_1236);
  nor csa_tree_add_7_25_groupi_g18002(csa_tree_add_7_25_groupi_n_3096 ,csa_tree_add_7_25_groupi_n_794 ,csa_tree_add_7_25_groupi_n_1712);
  nor csa_tree_add_7_25_groupi_g18003(csa_tree_add_7_25_groupi_n_3095 ,csa_tree_add_7_25_groupi_n_611 ,csa_tree_add_7_25_groupi_n_1717);
  nor csa_tree_add_7_25_groupi_g18004(csa_tree_add_7_25_groupi_n_3094 ,csa_tree_add_7_25_groupi_n_845 ,csa_tree_add_7_25_groupi_n_1354);
  nor csa_tree_add_7_25_groupi_g18005(csa_tree_add_7_25_groupi_n_3093 ,csa_tree_add_7_25_groupi_n_650 ,csa_tree_add_7_25_groupi_n_1667);
  nor csa_tree_add_7_25_groupi_g18006(csa_tree_add_7_25_groupi_n_3092 ,csa_tree_add_7_25_groupi_n_436 ,csa_tree_add_7_25_groupi_n_1333);
  nor csa_tree_add_7_25_groupi_g18007(csa_tree_add_7_25_groupi_n_3091 ,csa_tree_add_7_25_groupi_n_97 ,csa_tree_add_7_25_groupi_n_612);
  nor csa_tree_add_7_25_groupi_g18008(csa_tree_add_7_25_groupi_n_3090 ,csa_tree_add_7_25_groupi_n_606 ,csa_tree_add_7_25_groupi_n_1348);
  nor csa_tree_add_7_25_groupi_g18009(csa_tree_add_7_25_groupi_n_3089 ,csa_tree_add_7_25_groupi_n_648 ,csa_tree_add_7_25_groupi_n_1766);
  nor csa_tree_add_7_25_groupi_g18010(csa_tree_add_7_25_groupi_n_3088 ,csa_tree_add_7_25_groupi_n_794 ,csa_tree_add_7_25_groupi_n_1426);
  nor csa_tree_add_7_25_groupi_g18011(csa_tree_add_7_25_groupi_n_3087 ,csa_tree_add_7_25_groupi_n_594 ,csa_tree_add_7_25_groupi_n_170);
  nor csa_tree_add_7_25_groupi_g18012(csa_tree_add_7_25_groupi_n_3086 ,csa_tree_add_7_25_groupi_n_656 ,csa_tree_add_7_25_groupi_n_1298);
  nor csa_tree_add_7_25_groupi_g18013(csa_tree_add_7_25_groupi_n_3085 ,csa_tree_add_7_25_groupi_n_665 ,csa_tree_add_7_25_groupi_n_1768);
  nor csa_tree_add_7_25_groupi_g18014(csa_tree_add_7_25_groupi_n_3084 ,csa_tree_add_7_25_groupi_n_851 ,csa_tree_add_7_25_groupi_n_1375);
  nor csa_tree_add_7_25_groupi_g18015(csa_tree_add_7_25_groupi_n_3083 ,csa_tree_add_7_25_groupi_n_828 ,csa_tree_add_7_25_groupi_n_531);
  nor csa_tree_add_7_25_groupi_g18016(csa_tree_add_7_25_groupi_n_3082 ,csa_tree_add_7_25_groupi_n_659 ,csa_tree_add_7_25_groupi_n_1441);
  nor csa_tree_add_7_25_groupi_g18017(csa_tree_add_7_25_groupi_n_3081 ,csa_tree_add_7_25_groupi_n_668 ,csa_tree_add_7_25_groupi_n_1549);
  nor csa_tree_add_7_25_groupi_g18018(csa_tree_add_7_25_groupi_n_3080 ,csa_tree_add_7_25_groupi_n_609 ,csa_tree_add_7_25_groupi_n_1736);
  nor csa_tree_add_7_25_groupi_g18019(csa_tree_add_7_25_groupi_n_3079 ,csa_tree_add_7_25_groupi_n_828 ,csa_tree_add_7_25_groupi_n_1675);
  nor csa_tree_add_7_25_groupi_g18020(csa_tree_add_7_25_groupi_n_3078 ,csa_tree_add_7_25_groupi_n_657 ,csa_tree_add_7_25_groupi_n_1684);
  nor csa_tree_add_7_25_groupi_g18021(csa_tree_add_7_25_groupi_n_3077 ,csa_tree_add_7_25_groupi_n_666 ,csa_tree_add_7_25_groupi_n_1780);
  nor csa_tree_add_7_25_groupi_g18022(csa_tree_add_7_25_groupi_n_3076 ,csa_tree_add_7_25_groupi_n_692 ,csa_tree_add_7_25_groupi_n_1366);
  nor csa_tree_add_7_25_groupi_g18023(csa_tree_add_7_25_groupi_n_3075 ,csa_tree_add_7_25_groupi_n_821 ,csa_tree_add_7_25_groupi_n_246);
  nor csa_tree_add_7_25_groupi_g18024(csa_tree_add_7_25_groupi_n_3074 ,csa_tree_add_7_25_groupi_n_863 ,csa_tree_add_7_25_groupi_n_1393);
  nor csa_tree_add_7_25_groupi_g18025(csa_tree_add_7_25_groupi_n_3073 ,csa_tree_add_7_25_groupi_n_966 ,csa_tree_add_7_25_groupi_n_1292);
  nor csa_tree_add_7_25_groupi_g18026(csa_tree_add_7_25_groupi_n_3072 ,csa_tree_add_7_25_groupi_n_686 ,csa_tree_add_7_25_groupi_n_1769);
  nor csa_tree_add_7_25_groupi_g18027(csa_tree_add_7_25_groupi_n_3071 ,csa_tree_add_7_25_groupi_n_929 ,csa_tree_add_7_25_groupi_n_1486);
  nor csa_tree_add_7_25_groupi_g18028(csa_tree_add_7_25_groupi_n_3070 ,csa_tree_add_7_25_groupi_n_1044 ,csa_tree_add_7_25_groupi_n_1438);
  nor csa_tree_add_7_25_groupi_g18029(csa_tree_add_7_25_groupi_n_3069 ,csa_tree_add_7_25_groupi_n_695 ,csa_tree_add_7_25_groupi_n_162);
  nor csa_tree_add_7_25_groupi_g18030(csa_tree_add_7_25_groupi_n_3068 ,csa_tree_add_7_25_groupi_n_95 ,csa_tree_add_7_25_groupi_n_618);
  nor csa_tree_add_7_25_groupi_g18031(csa_tree_add_7_25_groupi_n_3067 ,csa_tree_add_7_25_groupi_n_1047 ,csa_tree_add_7_25_groupi_n_1525);
  nor csa_tree_add_7_25_groupi_g18032(csa_tree_add_7_25_groupi_n_3066 ,csa_tree_add_7_25_groupi_n_963 ,csa_tree_add_7_25_groupi_n_1297);
  nor csa_tree_add_7_25_groupi_g18033(csa_tree_add_7_25_groupi_n_3065 ,csa_tree_add_7_25_groupi_n_830 ,csa_tree_add_7_25_groupi_n_1328);
  nor csa_tree_add_7_25_groupi_g18034(csa_tree_add_7_25_groupi_n_3064 ,csa_tree_add_7_25_groupi_n_932 ,csa_tree_add_7_25_groupi_n_1462);
  nor csa_tree_add_7_25_groupi_g18035(csa_tree_add_7_25_groupi_n_3063 ,csa_tree_add_7_25_groupi_n_777 ,csa_tree_add_7_25_groupi_n_1699);
  nor csa_tree_add_7_25_groupi_g18036(csa_tree_add_7_25_groupi_n_3062 ,csa_tree_add_7_25_groupi_n_792 ,csa_tree_add_7_25_groupi_n_992);
  nor csa_tree_add_7_25_groupi_g18037(csa_tree_add_7_25_groupi_n_3061 ,csa_tree_add_7_25_groupi_n_821 ,csa_tree_add_7_25_groupi_n_2001);
  nor csa_tree_add_7_25_groupi_g18038(csa_tree_add_7_25_groupi_n_3060 ,csa_tree_add_7_25_groupi_n_930 ,csa_tree_add_7_25_groupi_n_513);
  nor csa_tree_add_7_25_groupi_g18039(csa_tree_add_7_25_groupi_n_3059 ,csa_tree_add_7_25_groupi_n_684 ,csa_tree_add_7_25_groupi_n_2000);
  nor csa_tree_add_7_25_groupi_g18040(csa_tree_add_7_25_groupi_n_3058 ,csa_tree_add_7_25_groupi_n_106 ,csa_tree_add_7_25_groupi_n_1757);
  nor csa_tree_add_7_25_groupi_g18041(csa_tree_add_7_25_groupi_n_3057 ,csa_tree_add_7_25_groupi_n_693 ,csa_tree_add_7_25_groupi_n_1501);
  nor csa_tree_add_7_25_groupi_g18042(csa_tree_add_7_25_groupi_n_3056 ,csa_tree_add_7_25_groupi_n_617 ,csa_tree_add_7_25_groupi_n_1489);
  nor csa_tree_add_7_25_groupi_g18043(csa_tree_add_7_25_groupi_n_3055 ,csa_tree_add_7_25_groupi_n_1035 ,csa_tree_add_7_25_groupi_n_518);
  nor csa_tree_add_7_25_groupi_g18044(csa_tree_add_7_25_groupi_n_3054 ,csa_tree_add_7_25_groupi_n_975 ,csa_tree_add_7_25_groupi_n_521);
  nor csa_tree_add_7_25_groupi_g18045(csa_tree_add_7_25_groupi_n_3053 ,csa_tree_add_7_25_groupi_n_991 ,csa_tree_add_7_25_groupi_n_621);
  nor csa_tree_add_7_25_groupi_g18046(csa_tree_add_7_25_groupi_n_3052 ,csa_tree_add_7_25_groupi_n_704 ,csa_tree_add_7_25_groupi_n_1523);
  nor csa_tree_add_7_25_groupi_g18047(csa_tree_add_7_25_groupi_n_3051 ,csa_tree_add_7_25_groupi_n_756 ,csa_tree_add_7_25_groupi_n_1913);
  nor csa_tree_add_7_25_groupi_g18048(csa_tree_add_7_25_groupi_n_3050 ,csa_tree_add_7_25_groupi_n_866 ,csa_tree_add_7_25_groupi_n_1355);
  nor csa_tree_add_7_25_groupi_g18049(csa_tree_add_7_25_groupi_n_3049 ,csa_tree_add_7_25_groupi_n_620 ,csa_tree_add_7_25_groupi_n_1427);
  nor csa_tree_add_7_25_groupi_g18050(csa_tree_add_7_25_groupi_n_3048 ,csa_tree_add_7_25_groupi_n_702 ,csa_tree_add_7_25_groupi_n_1232);
  nor csa_tree_add_7_25_groupi_g18051(csa_tree_add_7_25_groupi_n_3047 ,csa_tree_add_7_25_groupi_n_88 ,csa_tree_add_7_25_groupi_n_1349);
  nor csa_tree_add_7_25_groupi_g18052(csa_tree_add_7_25_groupi_n_3046 ,csa_tree_add_7_25_groupi_n_867 ,csa_tree_add_7_25_groupi_n_1166);
  nor csa_tree_add_7_25_groupi_g18053(csa_tree_add_7_25_groupi_n_3045 ,csa_tree_add_7_25_groupi_n_879 ,csa_tree_add_7_25_groupi_n_1763);
  nor csa_tree_add_7_25_groupi_g18054(csa_tree_add_7_25_groupi_n_3044 ,csa_tree_add_7_25_groupi_n_475 ,csa_tree_add_7_25_groupi_n_1297);
  nor csa_tree_add_7_25_groupi_g18055(csa_tree_add_7_25_groupi_n_3043 ,csa_tree_add_7_25_groupi_n_803 ,csa_tree_add_7_25_groupi_n_1925);
  nor csa_tree_add_7_25_groupi_g18056(csa_tree_add_7_25_groupi_n_3042 ,csa_tree_add_7_25_groupi_n_680 ,csa_tree_add_7_25_groupi_n_1851);
  nor csa_tree_add_7_25_groupi_g18057(csa_tree_add_7_25_groupi_n_3041 ,csa_tree_add_7_25_groupi_n_842 ,csa_tree_add_7_25_groupi_n_1685);
  nor csa_tree_add_7_25_groupi_g18058(csa_tree_add_7_25_groupi_n_3040 ,csa_tree_add_7_25_groupi_n_809 ,csa_tree_add_7_25_groupi_n_2000);
  nor csa_tree_add_7_25_groupi_g18059(csa_tree_add_7_25_groupi_n_3039 ,csa_tree_add_7_25_groupi_n_926 ,csa_tree_add_7_25_groupi_n_1724);
  nor csa_tree_add_7_25_groupi_g18060(csa_tree_add_7_25_groupi_n_3038 ,csa_tree_add_7_25_groupi_n_674 ,csa_tree_add_7_25_groupi_n_510);
  nor csa_tree_add_7_25_groupi_g18061(csa_tree_add_7_25_groupi_n_3037 ,csa_tree_add_7_25_groupi_n_662 ,csa_tree_add_7_25_groupi_n_1438);
  nor csa_tree_add_7_25_groupi_g18062(csa_tree_add_7_25_groupi_n_3036 ,csa_tree_add_7_25_groupi_n_911 ,csa_tree_add_7_25_groupi_n_1667);
  nor csa_tree_add_7_25_groupi_g18063(csa_tree_add_7_25_groupi_n_3035 ,csa_tree_add_7_25_groupi_n_737 ,csa_tree_add_7_25_groupi_n_1463);
  nor csa_tree_add_7_25_groupi_g18064(csa_tree_add_7_25_groupi_n_3034 ,csa_tree_add_7_25_groupi_n_1071 ,csa_tree_add_7_25_groupi_n_139);
  nor csa_tree_add_7_25_groupi_g18065(csa_tree_add_7_25_groupi_n_3033 ,csa_tree_add_7_25_groupi_n_881 ,csa_tree_add_7_25_groupi_n_1393);
  nor csa_tree_add_7_25_groupi_g18066(csa_tree_add_7_25_groupi_n_3032 ,csa_tree_add_7_25_groupi_n_893 ,csa_tree_add_7_25_groupi_n_1499);
  nor csa_tree_add_7_25_groupi_g18067(csa_tree_add_7_25_groupi_n_3031 ,csa_tree_add_7_25_groupi_n_857 ,csa_tree_add_7_25_groupi_n_1511);
  nor csa_tree_add_7_25_groupi_g18068(csa_tree_add_7_25_groupi_n_3030 ,csa_tree_add_7_25_groupi_n_815 ,csa_tree_add_7_25_groupi_n_518);
  nor csa_tree_add_7_25_groupi_g18069(csa_tree_add_7_25_groupi_n_3029 ,csa_tree_add_7_25_groupi_n_1005 ,csa_tree_add_7_25_groupi_n_1159);
  nor csa_tree_add_7_25_groupi_g18070(csa_tree_add_7_25_groupi_n_3028 ,csa_tree_add_7_25_groupi_n_854 ,csa_tree_add_7_25_groupi_n_1370);
  nor csa_tree_add_7_25_groupi_g18071(csa_tree_add_7_25_groupi_n_3027 ,csa_tree_add_7_25_groupi_n_719 ,csa_tree_add_7_25_groupi_n_1339);
  nor csa_tree_add_7_25_groupi_g18072(csa_tree_add_7_25_groupi_n_3026 ,csa_tree_add_7_25_groupi_n_1011 ,csa_tree_add_7_25_groupi_n_515);
  nor csa_tree_add_7_25_groupi_g18073(csa_tree_add_7_25_groupi_n_3025 ,csa_tree_add_7_25_groupi_n_1023 ,csa_tree_add_7_25_groupi_n_519);
  nor csa_tree_add_7_25_groupi_g18074(csa_tree_add_7_25_groupi_n_3024 ,csa_tree_add_7_25_groupi_n_873 ,csa_tree_add_7_25_groupi_n_530);
  nor csa_tree_add_7_25_groupi_g18075(csa_tree_add_7_25_groupi_n_3023 ,csa_tree_add_7_25_groupi_n_899 ,csa_tree_add_7_25_groupi_n_1520);
  nor csa_tree_add_7_25_groupi_g18076(csa_tree_add_7_25_groupi_n_3022 ,csa_tree_add_7_25_groupi_n_920 ,csa_tree_add_7_25_groupi_n_1525);
  nor csa_tree_add_7_25_groupi_g18077(csa_tree_add_7_25_groupi_n_3021 ,csa_tree_add_7_25_groupi_n_945 ,csa_tree_add_7_25_groupi_n_170);
  nor csa_tree_add_7_25_groupi_g18078(csa_tree_add_7_25_groupi_n_3020 ,csa_tree_add_7_25_groupi_n_1080 ,csa_tree_add_7_25_groupi_n_1291);
  nor csa_tree_add_7_25_groupi_g18079(csa_tree_add_7_25_groupi_n_3019 ,csa_tree_add_7_25_groupi_n_917 ,csa_tree_add_7_25_groupi_n_2004);
  nor csa_tree_add_7_25_groupi_g18080(csa_tree_add_7_25_groupi_n_3018 ,csa_tree_add_7_25_groupi_n_1029 ,csa_tree_add_7_25_groupi_n_530);
  nor csa_tree_add_7_25_groupi_g18081(csa_tree_add_7_25_groupi_n_3017 ,csa_tree_add_7_25_groupi_n_888 ,csa_tree_add_7_25_groupi_n_516);
  nor csa_tree_add_7_25_groupi_g18082(csa_tree_add_7_25_groupi_n_3016 ,csa_tree_add_7_25_groupi_n_1062 ,csa_tree_add_7_25_groupi_n_1778);
  nor csa_tree_add_7_25_groupi_g18083(csa_tree_add_7_25_groupi_n_3015 ,csa_tree_add_7_25_groupi_n_1056 ,csa_tree_add_7_25_groupi_n_1339);
  nor csa_tree_add_7_25_groupi_g18084(csa_tree_add_7_25_groupi_n_3014 ,csa_tree_add_7_25_groupi_n_1074 ,csa_tree_add_7_25_groupi_n_1561);
  nor csa_tree_add_7_25_groupi_g18085(csa_tree_add_7_25_groupi_n_3013 ,csa_tree_add_7_25_groupi_n_1077 ,csa_tree_add_7_25_groupi_n_1780);
  nor csa_tree_add_7_25_groupi_g18086(csa_tree_add_7_25_groupi_n_3012 ,csa_tree_add_7_25_groupi_n_969 ,csa_tree_add_7_25_groupi_n_1489);
  nor csa_tree_add_7_25_groupi_g18087(csa_tree_add_7_25_groupi_n_3011 ,csa_tree_add_7_25_groupi_n_972 ,csa_tree_add_7_25_groupi_n_1501);
  nor csa_tree_add_7_25_groupi_g18088(csa_tree_add_7_25_groupi_n_3010 ,csa_tree_add_7_25_groupi_n_710 ,csa_tree_add_7_25_groupi_n_1432);
  nor csa_tree_add_7_25_groupi_g18089(csa_tree_add_7_25_groupi_n_3009 ,csa_tree_add_7_25_groupi_n_896 ,csa_tree_add_7_25_groupi_n_1673);
  nor csa_tree_add_7_25_groupi_g18090(csa_tree_add_7_25_groupi_n_3008 ,csa_tree_add_7_25_groupi_n_1014 ,csa_tree_add_7_25_groupi_n_1532);
  nor csa_tree_add_7_25_groupi_g18091(csa_tree_add_7_25_groupi_n_3007 ,csa_tree_add_7_25_groupi_n_677 ,csa_tree_add_7_25_groupi_n_1424);
  nor csa_tree_add_7_25_groupi_g18092(csa_tree_add_7_25_groupi_n_3006 ,csa_tree_add_7_25_groupi_n_1038 ,csa_tree_add_7_25_groupi_n_1447);
  nor csa_tree_add_7_25_groupi_g18093(csa_tree_add_7_25_groupi_n_3005 ,csa_tree_add_7_25_groupi_n_869 ,csa_tree_add_7_25_groupi_n_1738);
  nor csa_tree_add_7_25_groupi_g18094(csa_tree_add_7_25_groupi_n_3004 ,csa_tree_add_7_25_groupi_n_1032 ,csa_tree_add_7_25_groupi_n_1334);
  nor csa_tree_add_7_25_groupi_g18095(csa_tree_add_7_25_groupi_n_3003 ,csa_tree_add_7_25_groupi_n_1017 ,csa_tree_add_7_25_groupi_n_522);
  nor csa_tree_add_7_25_groupi_g18096(csa_tree_add_7_25_groupi_n_3002 ,csa_tree_add_7_25_groupi_n_902 ,csa_tree_add_7_25_groupi_n_1729);
  nor csa_tree_add_7_25_groupi_g18097(csa_tree_add_7_25_groupi_n_3001 ,csa_tree_add_7_25_groupi_n_1065 ,csa_tree_add_7_25_groupi_n_1160);
  nor csa_tree_add_7_25_groupi_g18098(csa_tree_add_7_25_groupi_n_3000 ,csa_tree_add_7_25_groupi_n_1008 ,csa_tree_add_7_25_groupi_n_95);
  nor csa_tree_add_7_25_groupi_g18099(csa_tree_add_7_25_groupi_n_2999 ,csa_tree_add_7_25_groupi_n_1026 ,csa_tree_add_7_25_groupi_n_164);
  nor csa_tree_add_7_25_groupi_g18100(csa_tree_add_7_25_groupi_n_2998 ,csa_tree_add_7_25_groupi_n_1050 ,csa_tree_add_7_25_groupi_n_531);
  nor csa_tree_add_7_25_groupi_g18101(csa_tree_add_7_25_groupi_n_2997 ,csa_tree_add_7_25_groupi_n_957 ,csa_tree_add_7_25_groupi_n_1508);
  nor csa_tree_add_7_25_groupi_g18102(csa_tree_add_7_25_groupi_n_2996 ,csa_tree_add_7_25_groupi_n_1041 ,csa_tree_add_7_25_groupi_n_1736);
  nor csa_tree_add_7_25_groupi_g18103(csa_tree_add_7_25_groupi_n_2995 ,csa_tree_add_7_25_groupi_n_1059 ,csa_tree_add_7_25_groupi_n_164);
  nor csa_tree_add_7_25_groupi_g18104(csa_tree_add_7_25_groupi_n_2994 ,csa_tree_add_7_25_groupi_n_1068 ,csa_tree_add_7_25_groupi_n_1852);
  nor csa_tree_add_7_25_groupi_g18105(csa_tree_add_7_25_groupi_n_2993 ,csa_tree_add_7_25_groupi_n_978 ,csa_tree_add_7_25_groupi_n_136);
  nor csa_tree_add_7_25_groupi_g18106(csa_tree_add_7_25_groupi_n_2992 ,csa_tree_add_7_25_groupi_n_960 ,csa_tree_add_7_25_groupi_n_1741);
  nor csa_tree_add_7_25_groupi_g18107(csa_tree_add_7_25_groupi_n_2991 ,csa_tree_add_7_25_groupi_n_909 ,csa_tree_add_7_25_groupi_n_1762);
  nor csa_tree_add_7_25_groupi_g18108(csa_tree_add_7_25_groupi_n_2990 ,csa_tree_add_7_25_groupi_n_1053 ,csa_tree_add_7_25_groupi_n_512);
  nor csa_tree_add_7_25_groupi_g18109(csa_tree_add_7_25_groupi_n_2989 ,csa_tree_add_7_25_groupi_n_1086 ,csa_tree_add_7_25_groupi_n_1445);
  nor csa_tree_add_7_25_groupi_g18110(csa_tree_add_7_25_groupi_n_2988 ,csa_tree_add_7_25_groupi_n_914 ,csa_tree_add_7_25_groupi_n_521);
  nor csa_tree_add_7_25_groupi_g18111(csa_tree_add_7_25_groupi_n_2987 ,csa_tree_add_7_25_groupi_n_989 ,csa_tree_add_7_25_groupi_n_615);
  nor csa_tree_add_7_25_groupi_g18112(csa_tree_add_7_25_groupi_n_2986 ,csa_tree_add_7_25_groupi_n_1020 ,csa_tree_add_7_25_groupi_n_1432);
  nor csa_tree_add_7_25_groupi_g18113(csa_tree_add_7_25_groupi_n_2985 ,csa_tree_add_7_25_groupi_n_923 ,csa_tree_add_7_25_groupi_n_1669);
  nor csa_tree_add_7_25_groupi_g18114(csa_tree_add_7_25_groupi_n_2984 ,csa_tree_add_7_25_groupi_n_722 ,csa_tree_add_7_25_groupi_n_1436);
  nor csa_tree_add_7_25_groupi_g18115(csa_tree_add_7_25_groupi_n_2983 ,csa_tree_add_7_25_groupi_n_753 ,csa_tree_add_7_25_groupi_n_126);
  nor csa_tree_add_7_25_groupi_g18116(csa_tree_add_7_25_groupi_n_2982 ,csa_tree_add_7_25_groupi_n_954 ,csa_tree_add_7_25_groupi_n_1327);
  nor csa_tree_add_7_25_groupi_g18117(csa_tree_add_7_25_groupi_n_2981 ,csa_tree_add_7_25_groupi_n_731 ,csa_tree_add_7_25_groupi_n_1723);
  nor csa_tree_add_7_25_groupi_g18118(csa_tree_add_7_25_groupi_n_2980 ,csa_tree_add_7_25_groupi_n_654 ,csa_tree_add_7_25_groupi_n_1682);
  nor csa_tree_add_7_25_groupi_g18119(csa_tree_add_7_25_groupi_n_2979 ,csa_tree_add_7_25_groupi_n_1083 ,csa_tree_add_7_25_groupi_n_1523);
  nor csa_tree_add_7_25_groupi_g18120(csa_tree_add_7_25_groupi_n_2978 ,csa_tree_add_7_25_groupi_n_987 ,csa_tree_add_7_25_groupi_n_513);
  nor csa_tree_add_7_25_groupi_g18121(csa_tree_add_7_25_groupi_n_2977 ,csa_tree_add_7_25_groupi_n_672 ,csa_tree_add_7_25_groupi_n_1762);
  nor csa_tree_add_7_25_groupi_g18122(csa_tree_add_7_25_groupi_n_2976 ,csa_tree_add_7_25_groupi_n_905 ,csa_tree_add_7_25_groupi_n_1766);
  nor csa_tree_add_7_25_groupi_g18123(csa_tree_add_7_25_groupi_n_2975 ,csa_tree_add_7_25_groupi_n_735 ,csa_tree_add_7_25_groupi_n_1561);
  nor csa_tree_add_7_25_groupi_g18124(csa_tree_add_7_25_groupi_n_2974 ,csa_tree_add_7_25_groupi_n_825 ,csa_tree_add_7_25_groupi_n_1670);
  nor csa_tree_add_7_25_groupi_g18125(csa_tree_add_7_25_groupi_n_2973 ,csa_tree_add_7_25_groupi_n_743 ,csa_tree_add_7_25_groupi_n_1550);
  nor csa_tree_add_7_25_groupi_g18126(csa_tree_add_7_25_groupi_n_2972 ,csa_tree_add_7_25_groupi_n_801 ,csa_tree_add_7_25_groupi_n_2001);
  nor csa_tree_add_7_25_groupi_g18127(csa_tree_add_7_25_groupi_n_2971 ,csa_tree_add_7_25_groupi_n_759 ,csa_tree_add_7_25_groupi_n_1415);
  nor csa_tree_add_7_25_groupi_g18128(csa_tree_add_7_25_groupi_n_2970 ,csa_tree_add_7_25_groupi_n_690 ,csa_tree_add_7_25_groupi_n_1447);
  nor csa_tree_add_7_25_groupi_g18129(csa_tree_add_7_25_groupi_n_2969 ,csa_tree_add_7_25_groupi_n_981 ,csa_tree_add_7_25_groupi_n_1684);
  nor csa_tree_add_7_25_groupi_g18130(csa_tree_add_7_25_groupi_n_2968 ,csa_tree_add_7_25_groupi_n_699 ,csa_tree_add_7_25_groupi_n_510);
  nor csa_tree_add_7_25_groupi_g18131(csa_tree_add_7_25_groupi_n_2967 ,csa_tree_add_7_25_groupi_n_837 ,csa_tree_add_7_25_groupi_n_162);
  nor csa_tree_add_7_25_groupi_g18132(csa_tree_add_7_25_groupi_n_2966 ,csa_tree_add_7_25_groupi_n_948 ,csa_tree_add_7_25_groupi_n_1426);
  nor csa_tree_add_7_25_groupi_g18133(csa_tree_add_7_25_groupi_n_2965 ,csa_tree_add_7_25_groupi_n_708 ,csa_tree_add_7_25_groupi_n_1730);
  nor csa_tree_add_7_25_groupi_g18134(csa_tree_add_7_25_groupi_n_2964 ,csa_tree_add_7_25_groupi_n_717 ,csa_tree_add_7_25_groupi_n_1451);
  nor csa_tree_add_7_25_groupi_g18135(csa_tree_add_7_25_groupi_n_2963 ,csa_tree_add_7_25_groupi_n_726 ,csa_tree_add_7_25_groupi_n_1669);
  nor csa_tree_add_7_25_groupi_g18136(csa_tree_add_7_25_groupi_n_2962 ,csa_tree_add_7_25_groupi_n_747 ,csa_tree_add_7_25_groupi_n_1511);
  nor csa_tree_add_7_25_groupi_g18137(csa_tree_add_7_25_groupi_n_2961 ,csa_tree_add_7_25_groupi_n_891 ,csa_tree_add_7_25_groupi_n_989);
  nor csa_tree_add_7_25_groupi_g18138(csa_tree_add_7_25_groupi_n_2960 ,csa_tree_add_7_25_groupi_n_984 ,csa_tree_add_7_25_groupi_n_1742);
  nor csa_tree_add_7_25_groupi_g18139(csa_tree_add_7_25_groupi_n_2959 ,csa_tree_add_7_25_groupi_n_926 ,csa_tree_add_7_25_groupi_n_1712);
  nor csa_tree_add_7_25_groupi_g18140(csa_tree_add_7_25_groupi_n_2958 ,csa_tree_add_7_25_groupi_n_807 ,csa_tree_add_7_25_groupi_n_1676);
  nor csa_tree_add_7_25_groupi_g18141(csa_tree_add_7_25_groupi_n_2957 ,csa_tree_add_7_25_groupi_n_884 ,csa_tree_add_7_25_groupi_n_1910);
  nor csa_tree_add_7_25_groupi_g18142(csa_tree_add_7_25_groupi_n_2956 ,csa_tree_add_7_25_groupi_n_849 ,csa_tree_add_7_25_groupi_n_1699);
  nor csa_tree_add_7_25_groupi_g18143(csa_tree_add_7_25_groupi_n_2955 ,csa_tree_add_7_25_groupi_n_819 ,csa_tree_add_7_25_groupi_n_1502);
  nor csa_tree_add_7_25_groupi_g18144(csa_tree_add_7_25_groupi_n_2954 ,csa_tree_add_7_25_groupi_n_738 ,csa_tree_add_7_25_groupi_n_1928);
  nor csa_tree_add_7_25_groupi_g18145(csa_tree_add_7_25_groupi_n_2953 ,csa_tree_add_7_25_groupi_n_713 ,csa_tree_add_7_25_groupi_n_1376);
  nor csa_tree_add_7_25_groupi_g18146(csa_tree_add_7_25_groupi_n_2952 ,csa_tree_add_7_25_groupi_n_861 ,csa_tree_add_7_25_groupi_n_1354);
  nor csa_tree_add_7_25_groupi_g18147(csa_tree_add_7_25_groupi_n_2951 ,csa_tree_add_7_25_groupi_n_881 ,csa_tree_add_7_25_groupi_n_991);
  nor csa_tree_add_7_25_groupi_g18148(csa_tree_add_7_25_groupi_n_2950 ,csa_tree_add_7_25_groupi_n_720 ,csa_tree_add_7_25_groupi_n_519);
  nor csa_tree_add_7_25_groupi_g18149(csa_tree_add_7_25_groupi_n_2949 ,csa_tree_add_7_25_groupi_n_750 ,csa_tree_add_7_25_groupi_n_1765);
  nor csa_tree_add_7_25_groupi_g18150(csa_tree_add_7_25_groupi_n_2948 ,csa_tree_add_7_25_groupi_n_783 ,csa_tree_add_7_25_groupi_n_1738);
  nor csa_tree_add_7_25_groupi_g18151(csa_tree_add_7_25_groupi_n_2947 ,csa_tree_add_7_25_groupi_n_854 ,csa_tree_add_7_25_groupi_n_126);
  nor csa_tree_add_7_25_groupi_g18152(csa_tree_add_7_25_groupi_n_2946 ,csa_tree_add_7_25_groupi_n_798 ,csa_tree_add_7_25_groupi_n_1441);
  nor csa_tree_add_7_25_groupi_g18153(csa_tree_add_7_25_groupi_n_2945 ,csa_tree_add_7_25_groupi_n_813 ,csa_tree_add_7_25_groupi_n_1851);
  nor csa_tree_add_7_25_groupi_g18154(csa_tree_add_7_25_groupi_n_2944 ,csa_tree_add_7_25_groupi_n_803 ,csa_tree_add_7_25_groupi_n_2004);
  nor csa_tree_add_7_25_groupi_g18155(csa_tree_add_7_25_groupi_n_2943 ,csa_tree_add_7_25_groupi_n_815 ,csa_tree_add_7_25_groupi_n_97);
  nor csa_tree_add_7_25_groupi_g18156(csa_tree_add_7_25_groupi_n_2942 ,csa_tree_add_7_25_groupi_n_680 ,csa_tree_add_7_25_groupi_n_1370);
  nor csa_tree_add_7_25_groupi_g18157(csa_tree_add_7_25_groupi_n_2941 ,csa_tree_add_7_25_groupi_n_888 ,csa_tree_add_7_25_groupi_n_1462);
  nor csa_tree_add_7_25_groupi_g18158(csa_tree_add_7_25_groupi_n_2940 ,csa_tree_add_7_25_groupi_n_614 ,csa_tree_add_7_25_groupi_n_1291);
  nor csa_tree_add_7_25_groupi_g18159(csa_tree_add_7_25_groupi_n_2939 ,csa_tree_add_7_25_groupi_n_52 ,csa_tree_add_7_25_groupi_n_1348);
  nor csa_tree_add_7_25_groupi_g18160(csa_tree_add_7_25_groupi_n_2938 ,csa_tree_add_7_25_groupi_n_809 ,csa_tree_add_7_25_groupi_n_1742);
  nor csa_tree_add_7_25_groupi_g18161(csa_tree_add_7_25_groupi_n_2937 ,csa_tree_add_7_25_groupi_n_899 ,csa_tree_add_7_25_groupi_n_139);
  nor csa_tree_add_7_25_groupi_g18162(csa_tree_add_7_25_groupi_n_2936 ,csa_tree_add_7_25_groupi_n_729 ,csa_tree_add_7_25_groupi_n_509);
  nor csa_tree_add_7_25_groupi_g18163(csa_tree_add_7_25_groupi_n_2935 ,csa_tree_add_7_25_groupi_n_662 ,csa_tree_add_7_25_groupi_n_1768);
  nor csa_tree_add_7_25_groupi_g18164(csa_tree_add_7_25_groupi_n_2934 ,csa_tree_add_7_25_groupi_n_876 ,csa_tree_add_7_25_groupi_n_1366);
  nor csa_tree_add_7_25_groupi_g18165(csa_tree_add_7_25_groupi_n_2933 ,csa_tree_add_7_25_groupi_n_62 ,csa_tree_add_7_25_groupi_n_1439);
  nor csa_tree_add_7_25_groupi_g18166(csa_tree_add_7_25_groupi_n_2932 ,csa_tree_add_7_25_groupi_n_873 ,csa_tree_add_7_25_groupi_n_1442);
  nor csa_tree_add_7_25_groupi_g18167(csa_tree_add_7_25_groupi_n_2931 ,csa_tree_add_7_25_groupi_n_76 ,csa_tree_add_7_25_groupi_n_1165);
  nor csa_tree_add_7_25_groupi_g18168(csa_tree_add_7_25_groupi_n_2930 ,csa_tree_add_7_25_groupi_n_912 ,csa_tree_add_7_25_groupi_n_1499);
  nor csa_tree_add_7_25_groupi_g18169(csa_tree_add_7_25_groupi_n_2929 ,csa_tree_add_7_25_groupi_n_842 ,csa_tree_add_7_25_groupi_n_1717);
  nor csa_tree_add_7_25_groupi_g18170(csa_tree_add_7_25_groupi_n_2928 ,csa_tree_add_7_25_groupi_n_894 ,csa_tree_add_7_25_groupi_n_1526);
  nor csa_tree_add_7_25_groupi_g18171(csa_tree_add_7_25_groupi_n_2927 ,csa_tree_add_7_25_groupi_n_90 ,csa_tree_add_7_25_groupi_n_1778);
  nor csa_tree_add_7_25_groupi_g18172(csa_tree_add_7_25_groupi_n_2926 ,csa_tree_add_7_25_groupi_n_675 ,csa_tree_add_7_25_groupi_n_1724);
  or csa_tree_add_7_25_groupi_g18173(csa_tree_add_7_25_groupi_n_2925 ,csa_tree_add_7_25_groupi_n_32 ,csa_tree_add_7_25_groupi_n_509);
  nor csa_tree_add_7_25_groupi_g18174(csa_tree_add_7_25_groupi_n_2924 ,csa_tree_add_7_25_groupi_n_56 ,csa_tree_add_7_25_groupi_n_1723);
  nor csa_tree_add_7_25_groupi_g18175(csa_tree_add_7_25_groupi_n_2923 ,csa_tree_add_7_25_groupi_n_903 ,csa_tree_add_7_25_groupi_n_1292);
  nor csa_tree_add_7_25_groupi_g18176(csa_tree_add_7_25_groupi_n_2922 ,csa_tree_add_7_25_groupi_n_921 ,csa_tree_add_7_25_groupi_n_1700);
  nor csa_tree_add_7_25_groupi_g18177(csa_tree_add_7_25_groupi_n_2921 ,csa_tree_add_7_25_groupi_n_108 ,csa_tree_add_7_25_groupi_n_515);
  nor csa_tree_add_7_25_groupi_g18178(csa_tree_add_7_25_groupi_n_2920 ,csa_tree_add_7_25_groupi_n_58 ,csa_tree_add_7_25_groupi_n_1160);
  nor csa_tree_add_7_25_groupi_g18179(csa_tree_add_7_25_groupi_n_2919 ,csa_tree_add_7_25_groupi_n_110 ,csa_tree_add_7_25_groupi_n_1233);
  nor csa_tree_add_7_25_groupi_g18180(csa_tree_add_7_25_groupi_n_2918 ,csa_tree_add_7_25_groupi_n_711 ,csa_tree_add_7_25_groupi_n_1486);
  nor csa_tree_add_7_25_groupi_g18181(csa_tree_add_7_25_groupi_n_2917 ,csa_tree_add_7_25_groupi_n_70 ,csa_tree_add_7_25_groupi_n_1490);
  nor csa_tree_add_7_25_groupi_g18182(csa_tree_add_7_25_groupi_n_2916 ,csa_tree_add_7_25_groupi_n_80 ,csa_tree_add_7_25_groupi_n_1914);
  nor csa_tree_add_7_25_groupi_g18183(csa_tree_add_7_25_groupi_n_2915 ,csa_tree_add_7_25_groupi_n_60 ,csa_tree_add_7_25_groupi_n_1367);
  nor csa_tree_add_7_25_groupi_g18184(csa_tree_add_7_25_groupi_n_2914 ,csa_tree_add_7_25_groupi_n_48 ,csa_tree_add_7_25_groupi_n_94);
  nor csa_tree_add_7_25_groupi_g18185(csa_tree_add_7_25_groupi_n_2913 ,csa_tree_add_7_25_groupi_n_68 ,csa_tree_add_7_25_groupi_n_1487);
  or csa_tree_add_7_25_groupi_g18186(csa_tree_add_7_25_groupi_n_2912 ,csa_tree_add_7_25_groupi_n_212 ,csa_tree_add_7_25_groupi_n_548);
  and csa_tree_add_7_25_groupi_g18187(csa_tree_add_7_25_groupi_n_2911 ,csa_tree_add_7_25_groupi_n_241 ,csa_tree_add_7_25_groupi_n_122);
  nor csa_tree_add_7_25_groupi_g18188(csa_tree_add_7_25_groupi_n_2910 ,csa_tree_add_7_25_groupi_n_212 ,csa_tree_add_7_25_groupi_n_2084);
  and csa_tree_add_7_25_groupi_g18189(csa_tree_add_7_25_groupi_n_2909 ,csa_tree_add_7_25_groupi_n_2084 ,csa_tree_add_7_25_groupi_n_1232);
  and csa_tree_add_7_25_groupi_g18190(csa_tree_add_7_25_groupi_n_2908 ,csa_tree_add_7_25_groupi_n_554 ,csa_tree_add_7_25_groupi_n_506);
  and csa_tree_add_7_25_groupi_g18191(csa_tree_add_7_25_groupi_n_2907 ,csa_tree_add_7_25_groupi_n_551 ,csa_tree_add_7_25_groupi_n_501);
  and csa_tree_add_7_25_groupi_g18192(csa_tree_add_7_25_groupi_n_2906 ,csa_tree_add_7_25_groupi_n_1106 ,csa_tree_add_7_25_groupi_n_124);
  nor csa_tree_add_7_25_groupi_g18193(csa_tree_add_7_25_groupi_n_2905 ,csa_tree_add_7_25_groupi_n_1876 ,csa_tree_add_7_25_groupi_n_1992);
  nor csa_tree_add_7_25_groupi_g18194(csa_tree_add_7_25_groupi_n_2904 ,csa_tree_add_7_25_groupi_n_300 ,csa_tree_add_7_25_groupi_n_266);
  nor csa_tree_add_7_25_groupi_g18195(csa_tree_add_7_25_groupi_n_2903 ,csa_tree_add_7_25_groupi_n_1875 ,csa_tree_add_7_25_groupi_n_2033);
  nor csa_tree_add_7_25_groupi_g18196(csa_tree_add_7_25_groupi_n_2902 ,csa_tree_add_7_25_groupi_n_277 ,csa_tree_add_7_25_groupi_n_2081);
  nor csa_tree_add_7_25_groupi_g18197(csa_tree_add_7_25_groupi_n_2901 ,csa_tree_add_7_25_groupi_n_1875 ,csa_tree_add_7_25_groupi_n_2197);
  nor csa_tree_add_7_25_groupi_g18198(csa_tree_add_7_25_groupi_n_2900 ,csa_tree_add_7_25_groupi_n_276 ,csa_tree_add_7_25_groupi_n_2075);
  nor csa_tree_add_7_25_groupi_g18199(csa_tree_add_7_25_groupi_n_2899 ,csa_tree_add_7_25_groupi_n_740 ,csa_tree_add_7_25_groupi_n_277);
  nor csa_tree_add_7_25_groupi_g18200(csa_tree_add_7_25_groupi_n_2898 ,csa_tree_add_7_25_groupi_n_300 ,csa_tree_add_7_25_groupi_n_2078);
  nor csa_tree_add_7_25_groupi_g18201(csa_tree_add_7_25_groupi_n_2897 ,csa_tree_add_7_25_groupi_n_211 ,csa_tree_add_7_25_groupi_n_2087);
  and csa_tree_add_7_25_groupi_g18202(csa_tree_add_7_25_groupi_n_2896 ,csa_tree_add_7_25_groupi_n_2033 ,csa_tree_add_7_25_groupi_n_1997);
  and csa_tree_add_7_25_groupi_g18203(csa_tree_add_7_25_groupi_n_2895 ,csa_tree_add_7_25_groupi_n_1992 ,csa_tree_add_7_25_groupi_n_1238);
  and csa_tree_add_7_25_groupi_g18204(csa_tree_add_7_25_groupi_n_2894 ,csa_tree_add_7_25_groupi_n_2087 ,csa_tree_add_7_25_groupi_n_1244);
  and csa_tree_add_7_25_groupi_g18205(csa_tree_add_7_25_groupi_n_2893 ,csa_tree_add_7_25_groupi_n_2081 ,csa_tree_add_7_25_groupi_n_1235);
  and csa_tree_add_7_25_groupi_g18206(csa_tree_add_7_25_groupi_n_2892 ,csa_tree_add_7_25_groupi_n_2075 ,csa_tree_add_7_25_groupi_n_1241);
  and csa_tree_add_7_25_groupi_g18207(csa_tree_add_7_25_groupi_n_2891 ,csa_tree_add_7_25_groupi_n_2078 ,csa_tree_add_7_25_groupi_n_1229);
  xnor csa_tree_add_7_25_groupi_g18208(csa_tree_add_7_25_groupi_n_3199 ,csa_tree_add_7_25_groupi_n_2475 ,csa_tree_add_7_25_groupi_n_2586);
  not csa_tree_add_7_25_groupi_g18209(csa_tree_add_7_25_groupi_n_2886 ,csa_tree_add_7_25_groupi_n_2884);
  not csa_tree_add_7_25_groupi_g18210(csa_tree_add_7_25_groupi_n_2885 ,csa_tree_add_7_25_groupi_n_2884);
  not csa_tree_add_7_25_groupi_g18211(csa_tree_add_7_25_groupi_n_2883 ,csa_tree_add_7_25_groupi_n_2881);
  not csa_tree_add_7_25_groupi_g18212(csa_tree_add_7_25_groupi_n_2882 ,csa_tree_add_7_25_groupi_n_2881);
  not csa_tree_add_7_25_groupi_g18213(csa_tree_add_7_25_groupi_n_2880 ,csa_tree_add_7_25_groupi_n_2878);
  not csa_tree_add_7_25_groupi_g18214(csa_tree_add_7_25_groupi_n_2879 ,csa_tree_add_7_25_groupi_n_2878);
  not csa_tree_add_7_25_groupi_g18215(csa_tree_add_7_25_groupi_n_2877 ,csa_tree_add_7_25_groupi_n_2874);
  not csa_tree_add_7_25_groupi_g18216(csa_tree_add_7_25_groupi_n_2876 ,csa_tree_add_7_25_groupi_n_2874);
  not csa_tree_add_7_25_groupi_g18217(csa_tree_add_7_25_groupi_n_2875 ,csa_tree_add_7_25_groupi_n_2874);
  not csa_tree_add_7_25_groupi_g18218(csa_tree_add_7_25_groupi_n_2873 ,csa_tree_add_7_25_groupi_n_2870);
  not csa_tree_add_7_25_groupi_g18219(csa_tree_add_7_25_groupi_n_2872 ,csa_tree_add_7_25_groupi_n_2870);
  not csa_tree_add_7_25_groupi_g18220(csa_tree_add_7_25_groupi_n_2871 ,csa_tree_add_7_25_groupi_n_2870);
  not csa_tree_add_7_25_groupi_g18221(csa_tree_add_7_25_groupi_n_2869 ,csa_tree_add_7_25_groupi_n_1116);
  not csa_tree_add_7_25_groupi_g18223(csa_tree_add_7_25_groupi_n_2868 ,csa_tree_add_7_25_groupi_n_2867);
  not csa_tree_add_7_25_groupi_g18224(csa_tree_add_7_25_groupi_n_2866 ,csa_tree_add_7_25_groupi_n_1116);
  not csa_tree_add_7_25_groupi_g18225(csa_tree_add_7_25_groupi_n_2865 ,csa_tree_add_7_25_groupi_n_2867);
  not csa_tree_add_7_25_groupi_g18226(csa_tree_add_7_25_groupi_n_2864 ,csa_tree_add_7_25_groupi_n_2862);
  not csa_tree_add_7_25_groupi_g18227(csa_tree_add_7_25_groupi_n_2863 ,csa_tree_add_7_25_groupi_n_1989);
  not csa_tree_add_7_25_groupi_g18228(csa_tree_add_7_25_groupi_n_2861 ,csa_tree_add_7_25_groupi_n_1989);
  not csa_tree_add_7_25_groupi_g18229(csa_tree_add_7_25_groupi_n_2860 ,csa_tree_add_7_25_groupi_n_2862);
  not csa_tree_add_7_25_groupi_g18230(csa_tree_add_7_25_groupi_n_2859 ,csa_tree_add_7_25_groupi_n_2857);
  not csa_tree_add_7_25_groupi_g18231(csa_tree_add_7_25_groupi_n_2858 ,csa_tree_add_7_25_groupi_n_1985);
  not csa_tree_add_7_25_groupi_g18232(csa_tree_add_7_25_groupi_n_2856 ,csa_tree_add_7_25_groupi_n_1985);
  not csa_tree_add_7_25_groupi_g18233(csa_tree_add_7_25_groupi_n_2855 ,csa_tree_add_7_25_groupi_n_2857);
  not csa_tree_add_7_25_groupi_g18234(csa_tree_add_7_25_groupi_n_2854 ,csa_tree_add_7_25_groupi_n_2852);
  not csa_tree_add_7_25_groupi_g18235(csa_tree_add_7_25_groupi_n_2853 ,csa_tree_add_7_25_groupi_n_1983);
  not csa_tree_add_7_25_groupi_g18236(csa_tree_add_7_25_groupi_n_2851 ,csa_tree_add_7_25_groupi_n_1983);
  not csa_tree_add_7_25_groupi_g18237(csa_tree_add_7_25_groupi_n_2850 ,csa_tree_add_7_25_groupi_n_2852);
  not csa_tree_add_7_25_groupi_g18238(csa_tree_add_7_25_groupi_n_2849 ,csa_tree_add_7_25_groupi_n_2847);
  not csa_tree_add_7_25_groupi_g18239(csa_tree_add_7_25_groupi_n_2848 ,csa_tree_add_7_25_groupi_n_1979);
  not csa_tree_add_7_25_groupi_g18240(csa_tree_add_7_25_groupi_n_2846 ,csa_tree_add_7_25_groupi_n_1979);
  not csa_tree_add_7_25_groupi_g18241(csa_tree_add_7_25_groupi_n_2845 ,csa_tree_add_7_25_groupi_n_2847);
  not csa_tree_add_7_25_groupi_g18242(csa_tree_add_7_25_groupi_n_2844 ,csa_tree_add_7_25_groupi_n_2842);
  not csa_tree_add_7_25_groupi_g18243(csa_tree_add_7_25_groupi_n_2843 ,csa_tree_add_7_25_groupi_n_1967);
  not csa_tree_add_7_25_groupi_g18244(csa_tree_add_7_25_groupi_n_2841 ,csa_tree_add_7_25_groupi_n_1967);
  not csa_tree_add_7_25_groupi_g18245(csa_tree_add_7_25_groupi_n_2840 ,csa_tree_add_7_25_groupi_n_2842);
  not csa_tree_add_7_25_groupi_g18246(csa_tree_add_7_25_groupi_n_2839 ,csa_tree_add_7_25_groupi_n_160);
  not csa_tree_add_7_25_groupi_g18247(csa_tree_add_7_25_groupi_n_2838 ,csa_tree_add_7_25_groupi_n_1248);
  not csa_tree_add_7_25_groupi_g18251(csa_tree_add_7_25_groupi_n_2337 ,csa_tree_add_7_25_groupi_n_1248);
  not csa_tree_add_7_25_groupi_g18252(csa_tree_add_7_25_groupi_n_2336 ,csa_tree_add_7_25_groupi_n_2837);
  not csa_tree_add_7_25_groupi_g18253(csa_tree_add_7_25_groupi_n_2836 ,csa_tree_add_7_25_groupi_n_160);
  nor csa_tree_add_7_25_groupi_g18255(csa_tree_add_7_25_groupi_n_2835 ,in3[11] ,csa_tree_add_7_25_groupi_n_2675);
  nor csa_tree_add_7_25_groupi_g18256(csa_tree_add_7_25_groupi_n_2834 ,csa_tree_add_7_25_groupi_n_2352 ,csa_tree_add_7_25_groupi_n_2680);
  nor csa_tree_add_7_25_groupi_g18257(csa_tree_add_7_25_groupi_n_2833 ,in3[17] ,csa_tree_add_7_25_groupi_n_2667);
  nor csa_tree_add_7_25_groupi_g18258(csa_tree_add_7_25_groupi_n_2832 ,csa_tree_add_7_25_groupi_n_394 ,csa_tree_add_7_25_groupi_n_1553);
  or csa_tree_add_7_25_groupi_g18259(csa_tree_add_7_25_groupi_n_2831 ,csa_tree_add_7_25_groupi_n_938 ,csa_tree_add_7_25_groupi_n_117);
  nor csa_tree_add_7_25_groupi_g18260(csa_tree_add_7_25_groupi_n_2830 ,csa_tree_add_7_25_groupi_n_342 ,csa_tree_add_7_25_groupi_n_1688);
  nor csa_tree_add_7_25_groupi_g18261(csa_tree_add_7_25_groupi_n_2829 ,in3[5] ,csa_tree_add_7_25_groupi_n_2663);
  nor csa_tree_add_7_25_groupi_g18262(csa_tree_add_7_25_groupi_n_2828 ,csa_tree_add_7_25_groupi_n_1227 ,csa_tree_add_7_25_groupi_n_2674);
  nor csa_tree_add_7_25_groupi_g18263(csa_tree_add_7_25_groupi_n_2827 ,csa_tree_add_7_25_groupi_n_415 ,csa_tree_add_7_25_groupi_n_1694);
  nor csa_tree_add_7_25_groupi_g18264(csa_tree_add_7_25_groupi_n_2826 ,in3[14] ,csa_tree_add_7_25_groupi_n_2670);
  nor csa_tree_add_7_25_groupi_g18265(csa_tree_add_7_25_groupi_n_2825 ,csa_tree_add_7_25_groupi_n_2381 ,csa_tree_add_7_25_groupi_n_2673);
  nor csa_tree_add_7_25_groupi_g18266(csa_tree_add_7_25_groupi_n_2824 ,csa_tree_add_7_25_groupi_n_357 ,csa_tree_add_7_25_groupi_n_1696);
  nor csa_tree_add_7_25_groupi_g18267(csa_tree_add_7_25_groupi_n_2823 ,csa_tree_add_7_25_groupi_n_2351 ,csa_tree_add_7_25_groupi_n_2677);
  or csa_tree_add_7_25_groupi_g18268(csa_tree_add_7_25_groupi_n_2822 ,csa_tree_add_7_25_groupi_n_2384 ,csa_tree_add_7_25_groupi_n_2676);
  nor csa_tree_add_7_25_groupi_g18269(csa_tree_add_7_25_groupi_n_2821 ,csa_tree_add_7_25_groupi_n_2349 ,csa_tree_add_7_25_groupi_n_2669);
  nor csa_tree_add_7_25_groupi_g18270(csa_tree_add_7_25_groupi_n_2820 ,csa_tree_add_7_25_groupi_n_391 ,csa_tree_add_7_25_groupi_n_1690);
  nor csa_tree_add_7_25_groupi_g18271(csa_tree_add_7_25_groupi_n_2819 ,csa_tree_add_7_25_groupi_n_591 ,csa_tree_add_7_25_groupi_n_1705);
  nor csa_tree_add_7_25_groupi_g18272(csa_tree_add_7_25_groupi_n_2818 ,in3[8] ,csa_tree_add_7_25_groupi_n_2666);
  nor csa_tree_add_7_25_groupi_g18273(csa_tree_add_7_25_groupi_n_2817 ,csa_tree_add_7_25_groupi_n_1885 ,csa_tree_add_7_25_groupi_n_1703);
  nor csa_tree_add_7_25_groupi_g18274(csa_tree_add_7_25_groupi_n_2816 ,in3[20] ,csa_tree_add_7_25_groupi_n_2668);
  nor csa_tree_add_7_25_groupi_g18275(csa_tree_add_7_25_groupi_n_2815 ,csa_tree_add_7_25_groupi_n_997 ,csa_tree_add_7_25_groupi_n_1690);
  nor csa_tree_add_7_25_groupi_g18276(csa_tree_add_7_25_groupi_n_2814 ,in3[23] ,csa_tree_add_7_25_groupi_n_2672);
  nor csa_tree_add_7_25_groupi_g18277(csa_tree_add_7_25_groupi_n_2813 ,csa_tree_add_7_25_groupi_n_441 ,csa_tree_add_7_25_groupi_n_1703);
  nor csa_tree_add_7_25_groupi_g18278(csa_tree_add_7_25_groupi_n_2812 ,csa_tree_add_7_25_groupi_n_2350 ,csa_tree_add_7_25_groupi_n_2681);
  nor csa_tree_add_7_25_groupi_g18279(csa_tree_add_7_25_groupi_n_2811 ,csa_tree_add_7_25_groupi_n_624 ,csa_tree_add_7_25_groupi_n_1705);
  nor csa_tree_add_7_25_groupi_g18280(csa_tree_add_7_25_groupi_n_2810 ,csa_tree_add_7_25_groupi_n_2353 ,csa_tree_add_7_25_groupi_n_2664);
  and csa_tree_add_7_25_groupi_g18281(csa_tree_add_7_25_groupi_n_2809 ,csa_tree_add_7_25_groupi_n_1226 ,csa_tree_add_7_25_groupi_n_2665);
  nor csa_tree_add_7_25_groupi_g18282(csa_tree_add_7_25_groupi_n_2808 ,csa_tree_add_7_25_groupi_n_233 ,csa_tree_add_7_25_groupi_n_1696);
  nor csa_tree_add_7_25_groupi_g18283(csa_tree_add_7_25_groupi_n_2807 ,csa_tree_add_7_25_groupi_n_480 ,csa_tree_add_7_25_groupi_n_1706);
  nor csa_tree_add_7_25_groupi_g18284(csa_tree_add_7_25_groupi_n_2806 ,csa_tree_add_7_25_groupi_n_2382 ,csa_tree_add_7_25_groupi_n_2671);
  or csa_tree_add_7_25_groupi_g18285(csa_tree_add_7_25_groupi_n_2805 ,in3[26] ,csa_tree_add_7_25_groupi_n_2679);
  nor csa_tree_add_7_25_groupi_g18286(csa_tree_add_7_25_groupi_n_2804 ,csa_tree_add_7_25_groupi_n_102 ,csa_tree_add_7_25_groupi_n_1709);
  and csa_tree_add_7_25_groupi_g18287(csa_tree_add_7_25_groupi_n_2890 ,csa_tree_add_7_25_groupi_n_2423 ,csa_tree_add_7_25_groupi_n_2660);
  or csa_tree_add_7_25_groupi_g18288(csa_tree_add_7_25_groupi_n_2889 ,in3[31] ,csa_tree_add_7_25_groupi_n_2615);
  or csa_tree_add_7_25_groupi_g18289(csa_tree_add_7_25_groupi_n_2888 ,csa_tree_add_7_25_groupi_n_2373 ,csa_tree_add_7_25_groupi_n_2615);
  and csa_tree_add_7_25_groupi_g18290(csa_tree_add_7_25_groupi_n_2887 ,csa_tree_add_7_25_groupi_n_2657 ,csa_tree_add_7_25_groupi_n_2639);
  and csa_tree_add_7_25_groupi_g18291(csa_tree_add_7_25_groupi_n_2884 ,csa_tree_add_7_25_groupi_n_2698 ,csa_tree_add_7_25_groupi_n_2616);
  and csa_tree_add_7_25_groupi_g18292(csa_tree_add_7_25_groupi_n_2881 ,csa_tree_add_7_25_groupi_n_2616 ,csa_tree_add_7_25_groupi_n_2699);
  or csa_tree_add_7_25_groupi_g18293(csa_tree_add_7_25_groupi_n_2878 ,csa_tree_add_7_25_groupi_n_2638 ,csa_tree_add_7_25_groupi_n_2658);
  or csa_tree_add_7_25_groupi_g18294(csa_tree_add_7_25_groupi_n_2874 ,csa_tree_add_7_25_groupi_n_2648 ,csa_tree_add_7_25_groupi_n_2647);
  or csa_tree_add_7_25_groupi_g18295(csa_tree_add_7_25_groupi_n_2870 ,csa_tree_add_7_25_groupi_n_2662 ,csa_tree_add_7_25_groupi_n_2640);
  or csa_tree_add_7_25_groupi_g18296(csa_tree_add_7_25_groupi_n_2867 ,csa_tree_add_7_25_groupi_n_2661 ,csa_tree_add_7_25_groupi_n_2645);
  or csa_tree_add_7_25_groupi_g18297(csa_tree_add_7_25_groupi_n_2862 ,csa_tree_add_7_25_groupi_n_2654 ,csa_tree_add_7_25_groupi_n_2649);
  or csa_tree_add_7_25_groupi_g18298(csa_tree_add_7_25_groupi_n_2857 ,csa_tree_add_7_25_groupi_n_2637 ,csa_tree_add_7_25_groupi_n_2635);
  or csa_tree_add_7_25_groupi_g18299(csa_tree_add_7_25_groupi_n_2852 ,csa_tree_add_7_25_groupi_n_2656 ,csa_tree_add_7_25_groupi_n_2643);
  or csa_tree_add_7_25_groupi_g18300(csa_tree_add_7_25_groupi_n_2847 ,csa_tree_add_7_25_groupi_n_2653 ,csa_tree_add_7_25_groupi_n_2652);
  and csa_tree_add_7_25_groupi_g18301(csa_tree_add_7_25_groupi_n_2842 ,in3[0] ,csa_tree_add_7_25_groupi_n_2626);
  and csa_tree_add_7_25_groupi_g18302(csa_tree_add_7_25_groupi_n_2837 ,in3[0] ,csa_tree_add_7_25_groupi_n_2625);
  not csa_tree_add_7_25_groupi_g18303(csa_tree_add_7_25_groupi_n_2802 ,csa_tree_add_7_25_groupi_n_2800);
  not csa_tree_add_7_25_groupi_g18304(csa_tree_add_7_25_groupi_n_2801 ,csa_tree_add_7_25_groupi_n_2800);
  not csa_tree_add_7_25_groupi_g18305(csa_tree_add_7_25_groupi_n_2799 ,csa_tree_add_7_25_groupi_n_2797);
  not csa_tree_add_7_25_groupi_g18306(csa_tree_add_7_25_groupi_n_2798 ,csa_tree_add_7_25_groupi_n_2797);
  not csa_tree_add_7_25_groupi_g18307(csa_tree_add_7_25_groupi_n_2796 ,csa_tree_add_7_25_groupi_n_2793);
  not csa_tree_add_7_25_groupi_g18308(csa_tree_add_7_25_groupi_n_2795 ,csa_tree_add_7_25_groupi_n_2793);
  not csa_tree_add_7_25_groupi_g18309(csa_tree_add_7_25_groupi_n_2794 ,csa_tree_add_7_25_groupi_n_2793);
  not csa_tree_add_7_25_groupi_g18311(csa_tree_add_7_25_groupi_n_2792 ,csa_tree_add_7_25_groupi_n_1111);
  not csa_tree_add_7_25_groupi_g18312(csa_tree_add_7_25_groupi_n_2790 ,csa_tree_add_7_25_groupi_n_1111);
  not csa_tree_add_7_25_groupi_g18313(csa_tree_add_7_25_groupi_n_2334 ,csa_tree_add_7_25_groupi_n_2791);
  not csa_tree_add_7_25_groupi_g18316(csa_tree_add_7_25_groupi_n_2789 ,csa_tree_add_7_25_groupi_n_1110);
  not csa_tree_add_7_25_groupi_g18318(csa_tree_add_7_25_groupi_n_2788 ,csa_tree_add_7_25_groupi_n_2787);
  not csa_tree_add_7_25_groupi_g18319(csa_tree_add_7_25_groupi_n_2786 ,csa_tree_add_7_25_groupi_n_1110);
  not csa_tree_add_7_25_groupi_g18320(csa_tree_add_7_25_groupi_n_2785 ,csa_tree_add_7_25_groupi_n_2787);
  not csa_tree_add_7_25_groupi_g18322(csa_tree_add_7_25_groupi_n_2330 ,csa_tree_add_7_25_groupi_n_2784);
  not csa_tree_add_7_25_groupi_g18324(csa_tree_add_7_25_groupi_n_2783 ,csa_tree_add_7_25_groupi_n_2784);
  not csa_tree_add_7_25_groupi_g18325(csa_tree_add_7_25_groupi_n_2329 ,csa_tree_add_7_25_groupi_n_1112);
  not csa_tree_add_7_25_groupi_g18328(csa_tree_add_7_25_groupi_n_2782 ,csa_tree_add_7_25_groupi_n_1251);
  not csa_tree_add_7_25_groupi_g18329(csa_tree_add_7_25_groupi_n_2781 ,csa_tree_add_7_25_groupi_n_1249);
  not csa_tree_add_7_25_groupi_g18332(csa_tree_add_7_25_groupi_n_2327 ,csa_tree_add_7_25_groupi_n_1249);
  not csa_tree_add_7_25_groupi_g18333(csa_tree_add_7_25_groupi_n_2326 ,csa_tree_add_7_25_groupi_n_2780);
  not csa_tree_add_7_25_groupi_g18334(csa_tree_add_7_25_groupi_n_2779 ,csa_tree_add_7_25_groupi_n_1251);
  not csa_tree_add_7_25_groupi_g18336(csa_tree_add_7_25_groupi_n_2778 ,csa_tree_add_7_25_groupi_n_2776);
  not csa_tree_add_7_25_groupi_g18337(csa_tree_add_7_25_groupi_n_2777 ,csa_tree_add_7_25_groupi_n_1965);
  not csa_tree_add_7_25_groupi_g18338(csa_tree_add_7_25_groupi_n_2775 ,csa_tree_add_7_25_groupi_n_1965);
  not csa_tree_add_7_25_groupi_g18339(csa_tree_add_7_25_groupi_n_2774 ,csa_tree_add_7_25_groupi_n_2776);
  not csa_tree_add_7_25_groupi_g18340(csa_tree_add_7_25_groupi_n_2773 ,csa_tree_add_7_25_groupi_n_2771);
  not csa_tree_add_7_25_groupi_g18341(csa_tree_add_7_25_groupi_n_2772 ,csa_tree_add_7_25_groupi_n_1963);
  not csa_tree_add_7_25_groupi_g18342(csa_tree_add_7_25_groupi_n_2770 ,csa_tree_add_7_25_groupi_n_1963);
  not csa_tree_add_7_25_groupi_g18343(csa_tree_add_7_25_groupi_n_2769 ,csa_tree_add_7_25_groupi_n_2771);
  not csa_tree_add_7_25_groupi_g18344(csa_tree_add_7_25_groupi_n_2768 ,csa_tree_add_7_25_groupi_n_2766);
  not csa_tree_add_7_25_groupi_g18345(csa_tree_add_7_25_groupi_n_2767 ,csa_tree_add_7_25_groupi_n_1961);
  not csa_tree_add_7_25_groupi_g18346(csa_tree_add_7_25_groupi_n_2765 ,csa_tree_add_7_25_groupi_n_1961);
  not csa_tree_add_7_25_groupi_g18347(csa_tree_add_7_25_groupi_n_2764 ,csa_tree_add_7_25_groupi_n_2766);
  not csa_tree_add_7_25_groupi_g18348(csa_tree_add_7_25_groupi_n_2763 ,csa_tree_add_7_25_groupi_n_2761);
  not csa_tree_add_7_25_groupi_g18349(csa_tree_add_7_25_groupi_n_2762 ,csa_tree_add_7_25_groupi_n_1959);
  not csa_tree_add_7_25_groupi_g18350(csa_tree_add_7_25_groupi_n_2760 ,csa_tree_add_7_25_groupi_n_1959);
  not csa_tree_add_7_25_groupi_g18351(csa_tree_add_7_25_groupi_n_2759 ,csa_tree_add_7_25_groupi_n_2761);
  not csa_tree_add_7_25_groupi_g18352(csa_tree_add_7_25_groupi_n_2758 ,csa_tree_add_7_25_groupi_n_2756);
  not csa_tree_add_7_25_groupi_g18353(csa_tree_add_7_25_groupi_n_2757 ,csa_tree_add_7_25_groupi_n_1957);
  not csa_tree_add_7_25_groupi_g18354(csa_tree_add_7_25_groupi_n_2755 ,csa_tree_add_7_25_groupi_n_1957);
  not csa_tree_add_7_25_groupi_g18355(csa_tree_add_7_25_groupi_n_2754 ,csa_tree_add_7_25_groupi_n_2756);
  not csa_tree_add_7_25_groupi_g18356(csa_tree_add_7_25_groupi_n_2753 ,csa_tree_add_7_25_groupi_n_127);
  not csa_tree_add_7_25_groupi_g18357(csa_tree_add_7_25_groupi_n_2752 ,csa_tree_add_7_25_groupi_n_1246);
  not csa_tree_add_7_25_groupi_g18361(csa_tree_add_7_25_groupi_n_2325 ,csa_tree_add_7_25_groupi_n_1246);
  not csa_tree_add_7_25_groupi_g18362(csa_tree_add_7_25_groupi_n_2324 ,csa_tree_add_7_25_groupi_n_2751);
  not csa_tree_add_7_25_groupi_g18363(csa_tree_add_7_25_groupi_n_2750 ,csa_tree_add_7_25_groupi_n_127);
  not csa_tree_add_7_25_groupi_g18365(csa_tree_add_7_25_groupi_n_2749 ,csa_tree_add_7_25_groupi_n_130);
  not csa_tree_add_7_25_groupi_g18366(csa_tree_add_7_25_groupi_n_2748 ,csa_tree_add_7_25_groupi_n_1253);
  not csa_tree_add_7_25_groupi_g18370(csa_tree_add_7_25_groupi_n_2322 ,csa_tree_add_7_25_groupi_n_1253);
  not csa_tree_add_7_25_groupi_g18371(csa_tree_add_7_25_groupi_n_2321 ,csa_tree_add_7_25_groupi_n_2747);
  not csa_tree_add_7_25_groupi_g18372(csa_tree_add_7_25_groupi_n_2746 ,csa_tree_add_7_25_groupi_n_130);
  not csa_tree_add_7_25_groupi_g18374(csa_tree_add_7_25_groupi_n_2745 ,csa_tree_add_7_25_groupi_n_146);
  not csa_tree_add_7_25_groupi_g18375(csa_tree_add_7_25_groupi_n_2744 ,csa_tree_add_7_25_groupi_n_1252);
  not csa_tree_add_7_25_groupi_g18379(csa_tree_add_7_25_groupi_n_2319 ,csa_tree_add_7_25_groupi_n_1252);
  not csa_tree_add_7_25_groupi_g18380(csa_tree_add_7_25_groupi_n_2318 ,csa_tree_add_7_25_groupi_n_2743);
  not csa_tree_add_7_25_groupi_g18381(csa_tree_add_7_25_groupi_n_2742 ,csa_tree_add_7_25_groupi_n_146);
  not csa_tree_add_7_25_groupi_g18383(csa_tree_add_7_25_groupi_n_2741 ,csa_tree_add_7_25_groupi_n_137);
  not csa_tree_add_7_25_groupi_g18384(csa_tree_add_7_25_groupi_n_2740 ,csa_tree_add_7_25_groupi_n_1247);
  not csa_tree_add_7_25_groupi_g18388(csa_tree_add_7_25_groupi_n_2316 ,csa_tree_add_7_25_groupi_n_1247);
  not csa_tree_add_7_25_groupi_g18389(csa_tree_add_7_25_groupi_n_2315 ,csa_tree_add_7_25_groupi_n_2739);
  not csa_tree_add_7_25_groupi_g18390(csa_tree_add_7_25_groupi_n_2738 ,csa_tree_add_7_25_groupi_n_137);
  nor csa_tree_add_7_25_groupi_g18392(csa_tree_add_7_25_groupi_n_2737 ,csa_tree_add_7_25_groupi_n_112 ,csa_tree_add_7_25_groupi_n_120);
  nor csa_tree_add_7_25_groupi_g18393(csa_tree_add_7_25_groupi_n_2736 ,csa_tree_add_7_25_groupi_n_846 ,csa_tree_add_7_25_groupi_n_1697);
  or csa_tree_add_7_25_groupi_g18394(csa_tree_add_7_25_groupi_n_2735 ,csa_tree_add_7_25_groupi_n_22 ,csa_tree_add_7_25_groupi_n_491);
  nor csa_tree_add_7_25_groupi_g18395(csa_tree_add_7_25_groupi_n_2734 ,csa_tree_add_7_25_groupi_n_576 ,csa_tree_add_7_25_groupi_n_1693);
  nor csa_tree_add_7_25_groupi_g18396(csa_tree_add_7_25_groupi_n_2733 ,csa_tree_add_7_25_groupi_n_732 ,csa_tree_add_7_25_groupi_n_1708);
  nor csa_tree_add_7_25_groupi_g18397(csa_tree_add_7_25_groupi_n_2732 ,csa_tree_add_7_25_groupi_n_852 ,csa_tree_add_7_25_groupi_n_1693);
  nor csa_tree_add_7_25_groupi_g18398(csa_tree_add_7_25_groupi_n_2731 ,csa_tree_add_7_25_groupi_n_822 ,csa_tree_add_7_25_groupi_n_1552);
  nor csa_tree_add_7_25_groupi_g18399(csa_tree_add_7_25_groupi_n_2730 ,csa_tree_add_7_25_groupi_n_831 ,csa_tree_add_7_25_groupi_n_1687);
  or csa_tree_add_7_25_groupi_g18400(csa_tree_add_7_25_groupi_n_2729 ,csa_tree_add_7_25_groupi_n_36 ,csa_tree_add_7_25_groupi_n_117);
  or csa_tree_add_7_25_groupi_g18401(csa_tree_add_7_25_groupi_n_2728 ,csa_tree_add_7_25_groupi_n_34 ,csa_tree_add_7_25_groupi_n_489);
  or csa_tree_add_7_25_groupi_g18402(csa_tree_add_7_25_groupi_n_2727 ,csa_tree_add_7_25_groupi_n_8 ,csa_tree_add_7_25_groupi_n_119);
  or csa_tree_add_7_25_groupi_g18403(csa_tree_add_7_25_groupi_n_2726 ,csa_tree_add_7_25_groupi_n_10 ,csa_tree_add_7_25_groupi_n_488);
  or csa_tree_add_7_25_groupi_g18404(csa_tree_add_7_25_groupi_n_2725 ,csa_tree_add_7_25_groupi_n_16 ,csa_tree_add_7_25_groupi_n_488);
  or csa_tree_add_7_25_groupi_g18405(csa_tree_add_7_25_groupi_n_2724 ,csa_tree_add_7_25_groupi_n_12 ,csa_tree_add_7_25_groupi_n_489);
  or csa_tree_add_7_25_groupi_g18406(csa_tree_add_7_25_groupi_n_2723 ,csa_tree_add_7_25_groupi_n_26 ,csa_tree_add_7_25_groupi_n_491);
  or csa_tree_add_7_25_groupi_g18407(csa_tree_add_7_25_groupi_n_2722 ,csa_tree_add_7_25_groupi_n_14 ,csa_tree_add_7_25_groupi_n_492);
  nor csa_tree_add_7_25_groupi_g18408(csa_tree_add_7_25_groupi_n_2721 ,csa_tree_add_7_25_groupi_n_785 ,csa_tree_add_7_25_groupi_n_1709);
  or csa_tree_add_7_25_groupi_g18409(csa_tree_add_7_25_groupi_n_2720 ,csa_tree_add_7_25_groupi_n_40 ,csa_tree_add_7_25_groupi_n_492);
  or csa_tree_add_7_25_groupi_g18410(csa_tree_add_7_25_groupi_n_2719 ,csa_tree_add_7_25_groupi_n_18 ,csa_tree_add_7_25_groupi_n_119);
  or csa_tree_add_7_25_groupi_g18411(csa_tree_add_7_25_groupi_n_2718 ,csa_tree_add_7_25_groupi_n_99 ,csa_tree_add_7_25_groupi_n_1919);
  nor csa_tree_add_7_25_groupi_g18412(csa_tree_add_7_25_groupi_n_2717 ,csa_tree_add_7_25_groupi_n_705 ,csa_tree_add_7_25_groupi_n_1691);
  nor csa_tree_add_7_25_groupi_g18413(csa_tree_add_7_25_groupi_n_2716 ,csa_tree_add_7_25_groupi_n_681 ,csa_tree_add_7_25_groupi_n_1687);
  nor csa_tree_add_7_25_groupi_g18414(csa_tree_add_7_25_groupi_n_2715 ,csa_tree_add_7_25_groupi_n_855 ,csa_tree_add_7_25_groupi_n_1702);
  nor csa_tree_add_7_25_groupi_g18415(csa_tree_add_7_25_groupi_n_2714 ,csa_tree_add_7_25_groupi_n_816 ,csa_tree_add_7_25_groupi_n_1697);
  nor csa_tree_add_7_25_groupi_g18416(csa_tree_add_7_25_groupi_n_2713 ,csa_tree_add_7_25_groupi_n_804 ,csa_tree_add_7_25_groupi_n_1702);
  nor csa_tree_add_7_25_groupi_g18417(csa_tree_add_7_25_groupi_n_2712 ,csa_tree_add_7_25_groupi_n_810 ,csa_tree_add_7_25_groupi_n_1706);
  nor csa_tree_add_7_25_groupi_g18418(csa_tree_add_7_25_groupi_n_2711 ,csa_tree_add_7_25_groupi_n_858 ,csa_tree_add_7_25_groupi_n_1694);
  nor csa_tree_add_7_25_groupi_g18419(csa_tree_add_7_25_groupi_n_2710 ,csa_tree_add_7_25_groupi_n_882 ,csa_tree_add_7_25_groupi_n_1708);
  nor csa_tree_add_7_25_groupi_g18420(csa_tree_add_7_25_groupi_n_2709 ,csa_tree_add_7_25_groupi_n_663 ,csa_tree_add_7_25_groupi_n_1691);
  nor csa_tree_add_7_25_groupi_g18421(csa_tree_add_7_25_groupi_n_2708 ,csa_tree_add_7_25_groupi_n_927 ,csa_tree_add_7_25_groupi_n_1552);
  nor csa_tree_add_7_25_groupi_g18422(csa_tree_add_7_25_groupi_n_2707 ,csa_tree_add_7_25_groupi_n_900 ,csa_tree_add_7_25_groupi_n_1688);
  nor csa_tree_add_7_25_groupi_g18423(csa_tree_add_7_25_groupi_n_2706 ,csa_tree_add_7_25_groupi_n_843 ,csa_tree_add_7_25_groupi_n_1553);
  and csa_tree_add_7_25_groupi_g18424(csa_tree_add_7_25_groupi_n_2803 ,csa_tree_add_7_25_groupi_n_2600 ,csa_tree_add_7_25_groupi_n_2599);
  and csa_tree_add_7_25_groupi_g18425(csa_tree_add_7_25_groupi_n_2800 ,csa_tree_add_7_25_groupi_n_2694 ,csa_tree_add_7_25_groupi_n_2617);
  and csa_tree_add_7_25_groupi_g18426(csa_tree_add_7_25_groupi_n_2797 ,csa_tree_add_7_25_groupi_n_2617 ,csa_tree_add_7_25_groupi_n_2695);
  and csa_tree_add_7_25_groupi_g18427(csa_tree_add_7_25_groupi_n_2793 ,csa_tree_add_7_25_groupi_n_2618 ,csa_tree_add_7_25_groupi_n_2689);
  and csa_tree_add_7_25_groupi_g18428(csa_tree_add_7_25_groupi_n_2791 ,csa_tree_add_7_25_groupi_n_2688 ,csa_tree_add_7_25_groupi_n_2618);
  and csa_tree_add_7_25_groupi_g18429(csa_tree_add_7_25_groupi_n_2787 ,csa_tree_add_7_25_groupi_n_2619 ,csa_tree_add_7_25_groupi_n_2693);
  and csa_tree_add_7_25_groupi_g18430(csa_tree_add_7_25_groupi_n_2784 ,csa_tree_add_7_25_groupi_n_2692 ,csa_tree_add_7_25_groupi_n_2619);
  and csa_tree_add_7_25_groupi_g18431(csa_tree_add_7_25_groupi_n_2780 ,csa_tree_add_7_25_groupi_n_2696 ,csa_tree_add_7_25_groupi_n_2620);
  and csa_tree_add_7_25_groupi_g18432(csa_tree_add_7_25_groupi_n_2776 ,csa_tree_add_7_25_groupi_n_2620 ,csa_tree_add_7_25_groupi_n_2697);
  and csa_tree_add_7_25_groupi_g18433(csa_tree_add_7_25_groupi_n_2771 ,csa_tree_add_7_25_groupi_n_2621 ,csa_tree_add_7_25_groupi_n_2701);
  and csa_tree_add_7_25_groupi_g18434(csa_tree_add_7_25_groupi_n_2766 ,csa_tree_add_7_25_groupi_n_2623 ,csa_tree_add_7_25_groupi_n_2703);
  and csa_tree_add_7_25_groupi_g18435(csa_tree_add_7_25_groupi_n_2761 ,csa_tree_add_7_25_groupi_n_2624 ,csa_tree_add_7_25_groupi_n_2705);
  and csa_tree_add_7_25_groupi_g18436(csa_tree_add_7_25_groupi_n_2756 ,csa_tree_add_7_25_groupi_n_2622 ,csa_tree_add_7_25_groupi_n_2691);
  and csa_tree_add_7_25_groupi_g18437(csa_tree_add_7_25_groupi_n_2751 ,csa_tree_add_7_25_groupi_n_2702 ,csa_tree_add_7_25_groupi_n_2623);
  and csa_tree_add_7_25_groupi_g18438(csa_tree_add_7_25_groupi_n_2747 ,csa_tree_add_7_25_groupi_n_2700 ,csa_tree_add_7_25_groupi_n_2621);
  and csa_tree_add_7_25_groupi_g18439(csa_tree_add_7_25_groupi_n_2743 ,csa_tree_add_7_25_groupi_n_2704 ,csa_tree_add_7_25_groupi_n_2624);
  and csa_tree_add_7_25_groupi_g18440(csa_tree_add_7_25_groupi_n_2739 ,csa_tree_add_7_25_groupi_n_2690 ,csa_tree_add_7_25_groupi_n_2622);
  not csa_tree_add_7_25_groupi_g18441(csa_tree_add_7_25_groupi_n_2705 ,csa_tree_add_7_25_groupi_n_2704);
  not csa_tree_add_7_25_groupi_g18442(csa_tree_add_7_25_groupi_n_2703 ,csa_tree_add_7_25_groupi_n_2702);
  not csa_tree_add_7_25_groupi_g18443(csa_tree_add_7_25_groupi_n_2701 ,csa_tree_add_7_25_groupi_n_2700);
  not csa_tree_add_7_25_groupi_g18444(csa_tree_add_7_25_groupi_n_2699 ,csa_tree_add_7_25_groupi_n_2698);
  not csa_tree_add_7_25_groupi_g18445(csa_tree_add_7_25_groupi_n_2697 ,csa_tree_add_7_25_groupi_n_2696);
  not csa_tree_add_7_25_groupi_g18446(csa_tree_add_7_25_groupi_n_2695 ,csa_tree_add_7_25_groupi_n_2694);
  not csa_tree_add_7_25_groupi_g18447(csa_tree_add_7_25_groupi_n_2693 ,csa_tree_add_7_25_groupi_n_2692);
  not csa_tree_add_7_25_groupi_g18448(csa_tree_add_7_25_groupi_n_2691 ,csa_tree_add_7_25_groupi_n_2690);
  not csa_tree_add_7_25_groupi_g18449(csa_tree_add_7_25_groupi_n_2689 ,csa_tree_add_7_25_groupi_n_2688);
  not csa_tree_add_7_25_groupi_g18450(csa_tree_add_7_25_groupi_n_2686 ,csa_tree_add_7_25_groupi_n_2684);
  not csa_tree_add_7_25_groupi_g18451(csa_tree_add_7_25_groupi_n_2685 ,csa_tree_add_7_25_groupi_n_1971);
  not csa_tree_add_7_25_groupi_g18452(csa_tree_add_7_25_groupi_n_2683 ,csa_tree_add_7_25_groupi_n_1971);
  not csa_tree_add_7_25_groupi_g18453(csa_tree_add_7_25_groupi_n_2682 ,csa_tree_add_7_25_groupi_n_2684);
  or csa_tree_add_7_25_groupi_g18454(csa_tree_add_7_25_groupi_n_2681 ,csa_tree_add_7_25_groupi_n_2368 ,csa_tree_add_7_25_groupi_n_2543);
  or csa_tree_add_7_25_groupi_g18455(csa_tree_add_7_25_groupi_n_2680 ,csa_tree_add_7_25_groupi_n_2372 ,csa_tree_add_7_25_groupi_n_2549);
  or csa_tree_add_7_25_groupi_g18456(csa_tree_add_7_25_groupi_n_2679 ,in3[27] ,csa_tree_add_7_25_groupi_n_2558);
  nor csa_tree_add_7_25_groupi_g18457(csa_tree_add_7_25_groupi_n_2678 ,csa_tree_add_7_25_groupi_n_687 ,csa_tree_add_7_25_groupi_n_1430);
  or csa_tree_add_7_25_groupi_g18458(csa_tree_add_7_25_groupi_n_2677 ,csa_tree_add_7_25_groupi_n_2369 ,csa_tree_add_7_25_groupi_n_2547);
  or csa_tree_add_7_25_groupi_g18459(csa_tree_add_7_25_groupi_n_2676 ,csa_tree_add_7_25_groupi_n_2370 ,csa_tree_add_7_25_groupi_n_2523);
  or csa_tree_add_7_25_groupi_g18460(csa_tree_add_7_25_groupi_n_2675 ,in3[12] ,csa_tree_add_7_25_groupi_n_2540);
  or csa_tree_add_7_25_groupi_g18461(csa_tree_add_7_25_groupi_n_2674 ,csa_tree_add_7_25_groupi_n_2406 ,csa_tree_add_7_25_groupi_n_2535);
  or csa_tree_add_7_25_groupi_g18462(csa_tree_add_7_25_groupi_n_2673 ,csa_tree_add_7_25_groupi_n_2407 ,csa_tree_add_7_25_groupi_n_2525);
  or csa_tree_add_7_25_groupi_g18463(csa_tree_add_7_25_groupi_n_2672 ,in3[24] ,csa_tree_add_7_25_groupi_n_2554);
  or csa_tree_add_7_25_groupi_g18464(csa_tree_add_7_25_groupi_n_2671 ,csa_tree_add_7_25_groupi_n_2371 ,csa_tree_add_7_25_groupi_n_2529);
  or csa_tree_add_7_25_groupi_g18465(csa_tree_add_7_25_groupi_n_2670 ,in3[15] ,csa_tree_add_7_25_groupi_n_2542);
  or csa_tree_add_7_25_groupi_g18466(csa_tree_add_7_25_groupi_n_2669 ,csa_tree_add_7_25_groupi_n_2404 ,csa_tree_add_7_25_groupi_n_2537);
  or csa_tree_add_7_25_groupi_g18467(csa_tree_add_7_25_groupi_n_2668 ,in3[21] ,csa_tree_add_7_25_groupi_n_2552);
  or csa_tree_add_7_25_groupi_g18468(csa_tree_add_7_25_groupi_n_2667 ,in3[18] ,csa_tree_add_7_25_groupi_n_2546);
  or csa_tree_add_7_25_groupi_g18469(csa_tree_add_7_25_groupi_n_2666 ,in3[9] ,csa_tree_add_7_25_groupi_n_2532);
  nor csa_tree_add_7_25_groupi_g18470(csa_tree_add_7_25_groupi_n_2665 ,in3[3] ,csa_tree_add_7_25_groupi_n_2534);
  or csa_tree_add_7_25_groupi_g18471(csa_tree_add_7_25_groupi_n_2664 ,csa_tree_add_7_25_groupi_n_2405 ,csa_tree_add_7_25_groupi_n_2555);
  or csa_tree_add_7_25_groupi_g18472(csa_tree_add_7_25_groupi_n_2663 ,in3[6] ,csa_tree_add_7_25_groupi_n_2528);
  and csa_tree_add_7_25_groupi_g18473(csa_tree_add_7_25_groupi_n_2662 ,in3[17] ,csa_tree_add_7_25_groupi_n_2504);
  and csa_tree_add_7_25_groupi_g18474(csa_tree_add_7_25_groupi_n_2661 ,in3[14] ,csa_tree_add_7_25_groupi_n_2514);
  nor csa_tree_add_7_25_groupi_g18476(csa_tree_add_7_25_groupi_n_2659 ,csa_tree_add_7_25_groupi_n_597 ,csa_tree_add_7_25_groupi_n_1574);
  nor csa_tree_add_7_25_groupi_g18477(csa_tree_add_7_25_groupi_n_2658 ,in3[23] ,csa_tree_add_7_25_groupi_n_2517);
  or csa_tree_add_7_25_groupi_g18478(csa_tree_add_7_25_groupi_n_2657 ,csa_tree_add_7_25_groupi_n_2384 ,csa_tree_add_7_25_groupi_n_2507);
  and csa_tree_add_7_25_groupi_g18479(csa_tree_add_7_25_groupi_n_2656 ,in3[2] ,csa_tree_add_7_25_groupi_n_2515);
  nor csa_tree_add_7_25_groupi_g18480(csa_tree_add_7_25_groupi_n_2655 ,csa_tree_add_7_25_groupi_n_593 ,csa_tree_add_7_25_groupi_n_1580);
  and csa_tree_add_7_25_groupi_g18481(csa_tree_add_7_25_groupi_n_2654 ,in3[11] ,csa_tree_add_7_25_groupi_n_2513);
  and csa_tree_add_7_25_groupi_g18482(csa_tree_add_7_25_groupi_n_2653 ,in3[5] ,csa_tree_add_7_25_groupi_n_2500);
  nor csa_tree_add_7_25_groupi_g18483(csa_tree_add_7_25_groupi_n_2652 ,in3[5] ,csa_tree_add_7_25_groupi_n_2509);
  nor csa_tree_add_7_25_groupi_g18484(csa_tree_add_7_25_groupi_n_2651 ,csa_tree_add_7_25_groupi_n_788 ,csa_tree_add_7_25_groupi_n_1582);
  nor csa_tree_add_7_25_groupi_g18485(csa_tree_add_7_25_groupi_n_2650 ,csa_tree_add_7_25_groupi_n_770 ,csa_tree_add_7_25_groupi_n_1576);
  nor csa_tree_add_7_25_groupi_g18486(csa_tree_add_7_25_groupi_n_2649 ,in3[11] ,csa_tree_add_7_25_groupi_n_2508);
  and csa_tree_add_7_25_groupi_g18487(csa_tree_add_7_25_groupi_n_2648 ,in3[20] ,csa_tree_add_7_25_groupi_n_2506);
  nor csa_tree_add_7_25_groupi_g18488(csa_tree_add_7_25_groupi_n_2647 ,in3[20] ,csa_tree_add_7_25_groupi_n_2512);
  nor csa_tree_add_7_25_groupi_g18489(csa_tree_add_7_25_groupi_n_2646 ,csa_tree_add_7_25_groupi_n_579 ,csa_tree_add_7_25_groupi_n_1588);
  nor csa_tree_add_7_25_groupi_g18490(csa_tree_add_7_25_groupi_n_2645 ,in3[14] ,csa_tree_add_7_25_groupi_n_2505);
  nor csa_tree_add_7_25_groupi_g18491(csa_tree_add_7_25_groupi_n_2644 ,csa_tree_add_7_25_groupi_n_360 ,csa_tree_add_7_25_groupi_n_1586);
  nor csa_tree_add_7_25_groupi_g18492(csa_tree_add_7_25_groupi_n_2643 ,in3[2] ,csa_tree_add_7_25_groupi_n_2503);
  nor csa_tree_add_7_25_groupi_g18493(csa_tree_add_7_25_groupi_n_2642 ,csa_tree_add_7_25_groupi_n_399 ,csa_tree_add_7_25_groupi_n_1576);
  nor csa_tree_add_7_25_groupi_g18494(csa_tree_add_7_25_groupi_n_2641 ,csa_tree_add_7_25_groupi_n_421 ,csa_tree_add_7_25_groupi_n_1586);
  nor csa_tree_add_7_25_groupi_g18495(csa_tree_add_7_25_groupi_n_2640 ,in3[17] ,csa_tree_add_7_25_groupi_n_2511);
  or csa_tree_add_7_25_groupi_g18496(csa_tree_add_7_25_groupi_n_2639 ,in3[26] ,csa_tree_add_7_25_groupi_n_2516);
  and csa_tree_add_7_25_groupi_g18497(csa_tree_add_7_25_groupi_n_2638 ,in3[23] ,csa_tree_add_7_25_groupi_n_2501);
  and csa_tree_add_7_25_groupi_g18498(csa_tree_add_7_25_groupi_n_2637 ,in3[8] ,csa_tree_add_7_25_groupi_n_2510);
  nor csa_tree_add_7_25_groupi_g18499(csa_tree_add_7_25_groupi_n_2636 ,csa_tree_add_7_25_groupi_n_365 ,csa_tree_add_7_25_groupi_n_1588);
  nor csa_tree_add_7_25_groupi_g18500(csa_tree_add_7_25_groupi_n_2635 ,in3[8] ,csa_tree_add_7_25_groupi_n_2502);
  nor csa_tree_add_7_25_groupi_g18501(csa_tree_add_7_25_groupi_n_2634 ,csa_tree_add_7_25_groupi_n_347 ,csa_tree_add_7_25_groupi_n_1582);
  nor csa_tree_add_7_25_groupi_g18502(csa_tree_add_7_25_groupi_n_2633 ,csa_tree_add_7_25_groupi_n_623 ,csa_tree_add_7_25_groupi_n_1589);
  nor csa_tree_add_7_25_groupi_g18503(csa_tree_add_7_25_groupi_n_2632 ,csa_tree_add_7_25_groupi_n_66 ,csa_tree_add_7_25_groupi_n_1592);
  nor csa_tree_add_7_25_groupi_g18504(csa_tree_add_7_25_groupi_n_2631 ,csa_tree_add_7_25_groupi_n_633 ,csa_tree_add_7_25_groupi_n_1583);
  nor csa_tree_add_7_25_groupi_g18505(csa_tree_add_7_25_groupi_n_2630 ,csa_tree_add_7_25_groupi_n_481 ,csa_tree_add_7_25_groupi_n_1579);
  nor csa_tree_add_7_25_groupi_g18506(csa_tree_add_7_25_groupi_n_2629 ,csa_tree_add_7_25_groupi_n_465 ,csa_tree_add_7_25_groupi_n_1591);
  nor csa_tree_add_7_25_groupi_g18507(csa_tree_add_7_25_groupi_n_2628 ,csa_tree_add_7_25_groupi_n_444 ,csa_tree_add_7_25_groupi_n_1579);
  nor csa_tree_add_7_25_groupi_g18508(csa_tree_add_7_25_groupi_n_2627 ,csa_tree_add_7_25_groupi_n_457 ,csa_tree_add_7_25_groupi_n_1429);
  or csa_tree_add_7_25_groupi_g18509(csa_tree_add_7_25_groupi_n_2704 ,csa_tree_add_7_25_groupi_n_2526 ,csa_tree_add_7_25_groupi_n_2527);
  or csa_tree_add_7_25_groupi_g18510(csa_tree_add_7_25_groupi_n_2702 ,csa_tree_add_7_25_groupi_n_2538 ,csa_tree_add_7_25_groupi_n_2539);
  or csa_tree_add_7_25_groupi_g18511(csa_tree_add_7_25_groupi_n_2700 ,csa_tree_add_7_25_groupi_n_2536 ,csa_tree_add_7_25_groupi_n_2533);
  or csa_tree_add_7_25_groupi_g18512(csa_tree_add_7_25_groupi_n_2698 ,csa_tree_add_7_25_groupi_n_2524 ,csa_tree_add_7_25_groupi_n_2557);
  or csa_tree_add_7_25_groupi_g18513(csa_tree_add_7_25_groupi_n_2696 ,csa_tree_add_7_25_groupi_n_2544 ,csa_tree_add_7_25_groupi_n_2541);
  or csa_tree_add_7_25_groupi_g18514(csa_tree_add_7_25_groupi_n_2694 ,csa_tree_add_7_25_groupi_n_2556 ,csa_tree_add_7_25_groupi_n_2553);
  or csa_tree_add_7_25_groupi_g18515(csa_tree_add_7_25_groupi_n_2692 ,csa_tree_add_7_25_groupi_n_2548 ,csa_tree_add_7_25_groupi_n_2545);
  or csa_tree_add_7_25_groupi_g18516(csa_tree_add_7_25_groupi_n_2690 ,csa_tree_add_7_25_groupi_n_2530 ,csa_tree_add_7_25_groupi_n_2531);
  or csa_tree_add_7_25_groupi_g18517(csa_tree_add_7_25_groupi_n_2688 ,csa_tree_add_7_25_groupi_n_2550 ,csa_tree_add_7_25_groupi_n_2551);
  or csa_tree_add_7_25_groupi_g18518(csa_tree_add_7_25_groupi_n_2687 ,csa_tree_add_7_25_groupi_n_2385 ,csa_tree_add_7_25_groupi_n_2480);
  and csa_tree_add_7_25_groupi_g18519(csa_tree_add_7_25_groupi_n_2684 ,csa_tree_add_7_25_groupi_n_2409 ,csa_tree_add_7_25_groupi_n_2476);
  not csa_tree_add_7_25_groupi_g18520(csa_tree_add_7_25_groupi_n_2626 ,csa_tree_add_7_25_groupi_n_2625);
  nor csa_tree_add_7_25_groupi_g18521(csa_tree_add_7_25_groupi_n_2613 ,csa_tree_add_7_25_groupi_n_933 ,csa_tree_add_7_25_groupi_n_1573);
  nor csa_tree_add_7_25_groupi_g18522(csa_tree_add_7_25_groupi_n_2612 ,csa_tree_add_7_25_groupi_n_870 ,csa_tree_add_7_25_groupi_n_1592);
  nor csa_tree_add_7_25_groupi_g18523(csa_tree_add_7_25_groupi_n_2611 ,csa_tree_add_7_25_groupi_n_918 ,csa_tree_add_7_25_groupi_n_1577);
  nor csa_tree_add_7_25_groupi_g18524(csa_tree_add_7_25_groupi_n_2610 ,csa_tree_add_7_25_groupi_n_915 ,csa_tree_add_7_25_groupi_n_1573);
  nor csa_tree_add_7_25_groupi_g18525(csa_tree_add_7_25_groupi_n_2609 ,csa_tree_add_7_25_groupi_n_723 ,csa_tree_add_7_25_groupi_n_1585);
  nor csa_tree_add_7_25_groupi_g18526(csa_tree_add_7_25_groupi_n_2608 ,csa_tree_add_7_25_groupi_n_678 ,csa_tree_add_7_25_groupi_n_1583);
  nor csa_tree_add_7_25_groupi_g18527(csa_tree_add_7_25_groupi_n_2607 ,csa_tree_add_7_25_groupi_n_897 ,csa_tree_add_7_25_groupi_n_1585);
  nor csa_tree_add_7_25_groupi_g18528(csa_tree_add_7_25_groupi_n_2606 ,csa_tree_add_7_25_groupi_n_885 ,csa_tree_add_7_25_groupi_n_1589);
  nor csa_tree_add_7_25_groupi_g18529(csa_tree_add_7_25_groupi_n_2605 ,csa_tree_add_7_25_groupi_n_906 ,csa_tree_add_7_25_groupi_n_1580);
  nor csa_tree_add_7_25_groupi_g18530(csa_tree_add_7_25_groupi_n_2604 ,csa_tree_add_7_25_groupi_n_734 ,csa_tree_add_7_25_groupi_n_1591);
  nor csa_tree_add_7_25_groupi_g18531(csa_tree_add_7_25_groupi_n_2603 ,csa_tree_add_7_25_groupi_n_653 ,csa_tree_add_7_25_groupi_n_1577);
  nor csa_tree_add_7_25_groupi_g18532(csa_tree_add_7_25_groupi_n_2602 ,csa_tree_add_7_25_groupi_n_744 ,csa_tree_add_7_25_groupi_n_1429);
  nor csa_tree_add_7_25_groupi_g18533(csa_tree_add_7_25_groupi_n_2601 ,csa_tree_add_7_25_groupi_n_924 ,csa_tree_add_7_25_groupi_n_1574);
  or csa_tree_add_7_25_groupi_g18534(csa_tree_add_7_25_groupi_n_2600 ,csa_tree_add_7_25_groupi_n_2385 ,csa_tree_add_7_25_groupi_n_2498);
  or csa_tree_add_7_25_groupi_g18535(csa_tree_add_7_25_groupi_n_2599 ,in3[29] ,csa_tree_add_7_25_groupi_n_2499);
  nor csa_tree_add_7_25_groupi_g18536(csa_tree_add_7_25_groupi_n_2598 ,csa_tree_add_7_25_groupi_n_755 ,csa_tree_add_7_25_groupi_n_1430);
  xnor csa_tree_add_7_25_groupi_g18537(csa_tree_add_7_25_groupi_n_2597 ,in1[31] ,in1[30]);
  xnor csa_tree_add_7_25_groupi_g18538(csa_tree_add_7_25_groupi_n_2625 ,csa_tree_add_7_25_groupi_n_1227 ,in3[1]);
  xnor csa_tree_add_7_25_groupi_g18539(csa_tree_add_7_25_groupi_n_2596 ,in3[11] ,in2[9]);
  xnor csa_tree_add_7_25_groupi_g18540(csa_tree_add_7_25_groupi_n_2624 ,csa_tree_add_7_25_groupi_n_2407 ,in3[5]);
  xnor csa_tree_add_7_25_groupi_g18541(csa_tree_add_7_25_groupi_n_2595 ,in3[8] ,in2[6]);
  xnor csa_tree_add_7_25_groupi_g18542(csa_tree_add_7_25_groupi_n_2623 ,csa_tree_add_7_25_groupi_n_2404 ,in3[11]);
  xnor csa_tree_add_7_25_groupi_g18543(csa_tree_add_7_25_groupi_n_2622 ,csa_tree_add_7_25_groupi_n_2371 ,in3[8]);
  xnor csa_tree_add_7_25_groupi_g18544(csa_tree_add_7_25_groupi_n_2594 ,in3[5] ,in2[3]);
  xnor csa_tree_add_7_25_groupi_g18545(csa_tree_add_7_25_groupi_n_2621 ,csa_tree_add_7_25_groupi_n_2406 ,in3[2]);
  xnor csa_tree_add_7_25_groupi_g18546(csa_tree_add_7_25_groupi_n_2620 ,csa_tree_add_7_25_groupi_n_2368 ,in3[14]);
  xnor csa_tree_add_7_25_groupi_g18547(csa_tree_add_7_25_groupi_n_2593 ,in3[14] ,in2[12]);
  xnor csa_tree_add_7_25_groupi_g18548(csa_tree_add_7_25_groupi_n_2592 ,in3[17] ,in2[15]);
  xnor csa_tree_add_7_25_groupi_g18549(csa_tree_add_7_25_groupi_n_2619 ,csa_tree_add_7_25_groupi_n_2369 ,in3[17]);
  xnor csa_tree_add_7_25_groupi_g18550(csa_tree_add_7_25_groupi_n_2591 ,in3[20] ,in2[18]);
  xnor csa_tree_add_7_25_groupi_g18551(csa_tree_add_7_25_groupi_n_2618 ,csa_tree_add_7_25_groupi_n_2372 ,in3[20]);
  xnor csa_tree_add_7_25_groupi_g18552(csa_tree_add_7_25_groupi_n_2590 ,in3[23] ,in2[21]);
  xnor csa_tree_add_7_25_groupi_g18553(csa_tree_add_7_25_groupi_n_2617 ,csa_tree_add_7_25_groupi_n_2405 ,in3[23]);
  xnor csa_tree_add_7_25_groupi_g18554(csa_tree_add_7_25_groupi_n_2616 ,csa_tree_add_7_25_groupi_n_2370 ,in3[26]);
  xnor csa_tree_add_7_25_groupi_g18555(csa_tree_add_7_25_groupi_n_2589 ,in3[26] ,in2[24]);
  xnor csa_tree_add_7_25_groupi_g18556(csa_tree_add_7_25_groupi_n_2588 ,in3[29] ,in2[27]);
  xnor csa_tree_add_7_25_groupi_g18557(csa_tree_add_7_25_groupi_n_2615 ,in3[30] ,in3[29]);
  xnor csa_tree_add_7_25_groupi_g18558(csa_tree_add_7_25_groupi_n_2587 ,in1[8] ,in1[7]);
  xnor csa_tree_add_7_25_groupi_g18559(csa_tree_add_7_25_groupi_n_2586 ,in1[2] ,in1[1]);
  xnor csa_tree_add_7_25_groupi_g18560(csa_tree_add_7_25_groupi_n_2585 ,in1[11] ,in1[10]);
  xnor csa_tree_add_7_25_groupi_g18561(csa_tree_add_7_25_groupi_n_2584 ,in1[6] ,in1[5]);
  xnor csa_tree_add_7_25_groupi_g18562(csa_tree_add_7_25_groupi_n_2583 ,in1[13] ,in1[12]);
  xnor csa_tree_add_7_25_groupi_g18563(csa_tree_add_7_25_groupi_n_2582 ,in1[10] ,in1[9]);
  xnor csa_tree_add_7_25_groupi_g18564(csa_tree_add_7_25_groupi_n_2581 ,in1[4] ,in1[3]);
  xnor csa_tree_add_7_25_groupi_g18565(csa_tree_add_7_25_groupi_n_2580 ,in1[7] ,in1[6]);
  xnor csa_tree_add_7_25_groupi_g18566(csa_tree_add_7_25_groupi_n_2579 ,in1[3] ,in1[2]);
  xnor csa_tree_add_7_25_groupi_g18567(csa_tree_add_7_25_groupi_n_2578 ,in1[14] ,in1[13]);
  xnor csa_tree_add_7_25_groupi_g18568(csa_tree_add_7_25_groupi_n_2577 ,in1[5] ,in1[4]);
  xnor csa_tree_add_7_25_groupi_g18569(csa_tree_add_7_25_groupi_n_2576 ,in1[9] ,in1[8]);
  xnor csa_tree_add_7_25_groupi_g18570(csa_tree_add_7_25_groupi_n_2575 ,in1[12] ,in1[11]);
  xnor csa_tree_add_7_25_groupi_g18571(csa_tree_add_7_25_groupi_n_2574 ,in1[15] ,in1[14]);
  xnor csa_tree_add_7_25_groupi_g18572(csa_tree_add_7_25_groupi_n_2573 ,in1[16] ,in1[15]);
  xnor csa_tree_add_7_25_groupi_g18573(csa_tree_add_7_25_groupi_n_2572 ,in1[17] ,in1[16]);
  xnor csa_tree_add_7_25_groupi_g18574(csa_tree_add_7_25_groupi_n_2571 ,in1[18] ,in1[17]);
  xnor csa_tree_add_7_25_groupi_g18575(csa_tree_add_7_25_groupi_n_2570 ,in1[19] ,in1[18]);
  xnor csa_tree_add_7_25_groupi_g18576(csa_tree_add_7_25_groupi_n_2569 ,in1[20] ,in1[19]);
  xnor csa_tree_add_7_25_groupi_g18577(csa_tree_add_7_25_groupi_n_2568 ,in1[21] ,in1[20]);
  xnor csa_tree_add_7_25_groupi_g18578(csa_tree_add_7_25_groupi_n_2567 ,in1[22] ,in1[21]);
  xnor csa_tree_add_7_25_groupi_g18579(csa_tree_add_7_25_groupi_n_2566 ,in1[23] ,in1[22]);
  xnor csa_tree_add_7_25_groupi_g18580(csa_tree_add_7_25_groupi_n_2565 ,in1[24] ,in1[23]);
  xnor csa_tree_add_7_25_groupi_g18581(csa_tree_add_7_25_groupi_n_2564 ,in1[25] ,in1[24]);
  xnor csa_tree_add_7_25_groupi_g18582(csa_tree_add_7_25_groupi_n_2563 ,in1[26] ,in1[25]);
  xnor csa_tree_add_7_25_groupi_g18583(csa_tree_add_7_25_groupi_n_2562 ,in1[27] ,in1[26]);
  xnor csa_tree_add_7_25_groupi_g18584(csa_tree_add_7_25_groupi_n_2561 ,in1[28] ,in1[27]);
  xnor csa_tree_add_7_25_groupi_g18585(csa_tree_add_7_25_groupi_n_2560 ,in1[29] ,in1[28]);
  xnor csa_tree_add_7_25_groupi_g18586(csa_tree_add_7_25_groupi_n_2559 ,in1[30] ,in1[29]);
  xnor csa_tree_add_7_25_groupi_g18587(csa_tree_add_7_25_groupi_n_2614 ,in1[1] ,in1[0]);
  not csa_tree_add_7_25_groupi_g18588(csa_tree_add_7_25_groupi_n_2558 ,csa_tree_add_7_25_groupi_n_2557);
  not csa_tree_add_7_25_groupi_g18589(csa_tree_add_7_25_groupi_n_2556 ,csa_tree_add_7_25_groupi_n_2555);
  not csa_tree_add_7_25_groupi_g18590(csa_tree_add_7_25_groupi_n_2554 ,csa_tree_add_7_25_groupi_n_2553);
  not csa_tree_add_7_25_groupi_g18591(csa_tree_add_7_25_groupi_n_2552 ,csa_tree_add_7_25_groupi_n_2551);
  not csa_tree_add_7_25_groupi_g18592(csa_tree_add_7_25_groupi_n_2550 ,csa_tree_add_7_25_groupi_n_2549);
  not csa_tree_add_7_25_groupi_g18593(csa_tree_add_7_25_groupi_n_2548 ,csa_tree_add_7_25_groupi_n_2547);
  not csa_tree_add_7_25_groupi_g18594(csa_tree_add_7_25_groupi_n_2546 ,csa_tree_add_7_25_groupi_n_2545);
  not csa_tree_add_7_25_groupi_g18595(csa_tree_add_7_25_groupi_n_2544 ,csa_tree_add_7_25_groupi_n_2543);
  not csa_tree_add_7_25_groupi_g18596(csa_tree_add_7_25_groupi_n_2542 ,csa_tree_add_7_25_groupi_n_2541);
  not csa_tree_add_7_25_groupi_g18597(csa_tree_add_7_25_groupi_n_2540 ,csa_tree_add_7_25_groupi_n_2539);
  not csa_tree_add_7_25_groupi_g18598(csa_tree_add_7_25_groupi_n_2538 ,csa_tree_add_7_25_groupi_n_2537);
  not csa_tree_add_7_25_groupi_g18599(csa_tree_add_7_25_groupi_n_2536 ,csa_tree_add_7_25_groupi_n_2535);
  not csa_tree_add_7_25_groupi_g18600(csa_tree_add_7_25_groupi_n_2534 ,csa_tree_add_7_25_groupi_n_2533);
  not csa_tree_add_7_25_groupi_g18601(csa_tree_add_7_25_groupi_n_2532 ,csa_tree_add_7_25_groupi_n_2531);
  not csa_tree_add_7_25_groupi_g18602(csa_tree_add_7_25_groupi_n_2530 ,csa_tree_add_7_25_groupi_n_2529);
  not csa_tree_add_7_25_groupi_g18603(csa_tree_add_7_25_groupi_n_2528 ,csa_tree_add_7_25_groupi_n_2527);
  not csa_tree_add_7_25_groupi_g18604(csa_tree_add_7_25_groupi_n_2526 ,csa_tree_add_7_25_groupi_n_2525);
  not csa_tree_add_7_25_groupi_g18605(csa_tree_add_7_25_groupi_n_2524 ,csa_tree_add_7_25_groupi_n_2523);
  not csa_tree_add_7_25_groupi_g18606(csa_tree_add_7_25_groupi_n_2522 ,csa_tree_add_7_25_groupi_n_2520);
  not csa_tree_add_7_25_groupi_g18607(csa_tree_add_7_25_groupi_n_2521 ,csa_tree_add_7_25_groupi_n_1969);
  not csa_tree_add_7_25_groupi_g18608(csa_tree_add_7_25_groupi_n_2519 ,csa_tree_add_7_25_groupi_n_1969);
  not csa_tree_add_7_25_groupi_g18609(csa_tree_add_7_25_groupi_n_2518 ,csa_tree_add_7_25_groupi_n_2520);
  or csa_tree_add_7_25_groupi_g18610(csa_tree_add_7_25_groupi_n_2517 ,csa_tree_add_7_25_groupi_n_2375 ,in3[24]);
  or csa_tree_add_7_25_groupi_g18611(csa_tree_add_7_25_groupi_n_2516 ,csa_tree_add_7_25_groupi_n_2378 ,in3[27]);
  nor csa_tree_add_7_25_groupi_g18612(csa_tree_add_7_25_groupi_n_2515 ,csa_tree_add_7_25_groupi_n_2406 ,in3[4]);
  nor csa_tree_add_7_25_groupi_g18613(csa_tree_add_7_25_groupi_n_2514 ,csa_tree_add_7_25_groupi_n_2368 ,in3[16]);
  nor csa_tree_add_7_25_groupi_g18614(csa_tree_add_7_25_groupi_n_2513 ,csa_tree_add_7_25_groupi_n_2404 ,in3[13]);
  or csa_tree_add_7_25_groupi_g18615(csa_tree_add_7_25_groupi_n_2512 ,csa_tree_add_7_25_groupi_n_2411 ,in3[21]);
  or csa_tree_add_7_25_groupi_g18616(csa_tree_add_7_25_groupi_n_2511 ,csa_tree_add_7_25_groupi_n_2377 ,in3[18]);
  nor csa_tree_add_7_25_groupi_g18617(csa_tree_add_7_25_groupi_n_2510 ,csa_tree_add_7_25_groupi_n_2371 ,in3[10]);
  or csa_tree_add_7_25_groupi_g18618(csa_tree_add_7_25_groupi_n_2509 ,csa_tree_add_7_25_groupi_n_2374 ,in3[6]);
  or csa_tree_add_7_25_groupi_g18619(csa_tree_add_7_25_groupi_n_2508 ,csa_tree_add_7_25_groupi_n_2414 ,in3[12]);
  or csa_tree_add_7_25_groupi_g18620(csa_tree_add_7_25_groupi_n_2507 ,csa_tree_add_7_25_groupi_n_2370 ,in3[28]);
  nor csa_tree_add_7_25_groupi_g18621(csa_tree_add_7_25_groupi_n_2506 ,csa_tree_add_7_25_groupi_n_2372 ,in3[22]);
  or csa_tree_add_7_25_groupi_g18622(csa_tree_add_7_25_groupi_n_2505 ,csa_tree_add_7_25_groupi_n_2410 ,in3[15]);
  nor csa_tree_add_7_25_groupi_g18623(csa_tree_add_7_25_groupi_n_2504 ,csa_tree_add_7_25_groupi_n_2369 ,in3[19]);
  or csa_tree_add_7_25_groupi_g18624(csa_tree_add_7_25_groupi_n_2503 ,csa_tree_add_7_25_groupi_n_2379 ,in3[3]);
  or csa_tree_add_7_25_groupi_g18625(csa_tree_add_7_25_groupi_n_2502 ,csa_tree_add_7_25_groupi_n_2376 ,in3[9]);
  nor csa_tree_add_7_25_groupi_g18626(csa_tree_add_7_25_groupi_n_2501 ,csa_tree_add_7_25_groupi_n_2405 ,in3[25]);
  nor csa_tree_add_7_25_groupi_g18627(csa_tree_add_7_25_groupi_n_2500 ,csa_tree_add_7_25_groupi_n_2407 ,in3[7]);
  or csa_tree_add_7_25_groupi_g18628(csa_tree_add_7_25_groupi_n_2499 ,csa_tree_add_7_25_groupi_n_2373 ,in3[30]);
  or csa_tree_add_7_25_groupi_g18629(csa_tree_add_7_25_groupi_n_2498 ,csa_tree_add_7_25_groupi_n_2408 ,in3[31]);
  nor csa_tree_add_7_25_groupi_g18630(csa_tree_add_7_25_groupi_n_2497 ,in1[20] ,in1[19]);
  and csa_tree_add_7_25_groupi_g18631(csa_tree_add_7_25_groupi_n_2496 ,in3[2] ,in2[0]);
  or csa_tree_add_7_25_groupi_g18632(csa_tree_add_7_25_groupi_n_2495 ,csa_tree_add_7_25_groupi_n_62 ,csa_tree_add_7_25_groupi_n_46);
  nor csa_tree_add_7_25_groupi_g18633(csa_tree_add_7_25_groupi_n_2494 ,in1[5] ,in1[4]);
  nor csa_tree_add_7_25_groupi_g18635(csa_tree_add_7_25_groupi_n_2492 ,in1[22] ,in1[21]);
  nor csa_tree_add_7_25_groupi_g18636(csa_tree_add_7_25_groupi_n_2491 ,in1[7] ,in1[6]);
  nor csa_tree_add_7_25_groupi_g18637(csa_tree_add_7_25_groupi_n_2490 ,in1[11] ,in1[10]);
  nor csa_tree_add_7_25_groupi_g18638(csa_tree_add_7_25_groupi_n_2489 ,in1[30] ,in1[29]);
  and csa_tree_add_7_25_groupi_g18639(csa_tree_add_7_25_groupi_n_2488 ,in3[23] ,in2[21]);
  or csa_tree_add_7_25_groupi_g18640(csa_tree_add_7_25_groupi_n_2487 ,csa_tree_add_7_25_groupi_n_110 ,csa_tree_add_7_25_groupi_n_90);
  nor csa_tree_add_7_25_groupi_g18641(csa_tree_add_7_25_groupi_n_2486 ,in1[16] ,in1[15]);
  nor csa_tree_add_7_25_groupi_g18642(csa_tree_add_7_25_groupi_n_2485 ,in1[21] ,in1[20]);
  or csa_tree_add_7_25_groupi_g18643(csa_tree_add_7_25_groupi_n_2484 ,in3[23] ,in2[21]);
  nor csa_tree_add_7_25_groupi_g18644(csa_tree_add_7_25_groupi_n_2483 ,in1[28] ,in1[27]);
  or csa_tree_add_7_25_groupi_g18645(csa_tree_add_7_25_groupi_n_2482 ,csa_tree_add_7_25_groupi_n_590 ,csa_tree_add_7_25_groupi_n_599);
  nor csa_tree_add_7_25_groupi_g18646(csa_tree_add_7_25_groupi_n_2481 ,in1[14] ,in1[13]);
  or csa_tree_add_7_25_groupi_g18647(csa_tree_add_7_25_groupi_n_2480 ,csa_tree_add_7_25_groupi_n_2373 ,csa_tree_add_7_25_groupi_n_2408);
  nor csa_tree_add_7_25_groupi_g18648(csa_tree_add_7_25_groupi_n_2479 ,in3[2] ,in2[0]);
  or csa_tree_add_7_25_groupi_g18649(csa_tree_add_7_25_groupi_n_2478 ,csa_tree_add_7_25_groupi_n_224 ,csa_tree_add_7_25_groupi_n_244);
  or csa_tree_add_7_25_groupi_g18650(csa_tree_add_7_25_groupi_n_2477 ,csa_tree_add_7_25_groupi_n_608 ,csa_tree_add_7_25_groupi_n_20);
  and csa_tree_add_7_25_groupi_g18651(csa_tree_add_7_25_groupi_n_2557 ,in3[29] ,csa_tree_add_7_25_groupi_n_2378);
  or csa_tree_add_7_25_groupi_g18652(csa_tree_add_7_25_groupi_n_2555 ,csa_tree_add_7_25_groupi_n_2375 ,in3[26]);
  and csa_tree_add_7_25_groupi_g18653(csa_tree_add_7_25_groupi_n_2553 ,in3[26] ,csa_tree_add_7_25_groupi_n_2375);
  and csa_tree_add_7_25_groupi_g18654(csa_tree_add_7_25_groupi_n_2551 ,in3[23] ,csa_tree_add_7_25_groupi_n_2411);
  or csa_tree_add_7_25_groupi_g18655(csa_tree_add_7_25_groupi_n_2549 ,csa_tree_add_7_25_groupi_n_2411 ,in3[23]);
  or csa_tree_add_7_25_groupi_g18656(csa_tree_add_7_25_groupi_n_2547 ,csa_tree_add_7_25_groupi_n_2377 ,in3[20]);
  and csa_tree_add_7_25_groupi_g18657(csa_tree_add_7_25_groupi_n_2545 ,in3[20] ,csa_tree_add_7_25_groupi_n_2377);
  or csa_tree_add_7_25_groupi_g18658(csa_tree_add_7_25_groupi_n_2543 ,csa_tree_add_7_25_groupi_n_2410 ,in3[17]);
  and csa_tree_add_7_25_groupi_g18659(csa_tree_add_7_25_groupi_n_2541 ,in3[17] ,csa_tree_add_7_25_groupi_n_2410);
  and csa_tree_add_7_25_groupi_g18660(csa_tree_add_7_25_groupi_n_2539 ,in3[14] ,csa_tree_add_7_25_groupi_n_2414);
  nor csa_tree_add_7_25_groupi_g18661(csa_tree_add_7_25_groupi_n_2476 ,csa_tree_add_7_25_groupi_n_2383 ,in3[1]);
  or csa_tree_add_7_25_groupi_g18662(csa_tree_add_7_25_groupi_n_2537 ,csa_tree_add_7_25_groupi_n_2414 ,in3[14]);
  or csa_tree_add_7_25_groupi_g18663(csa_tree_add_7_25_groupi_n_2535 ,csa_tree_add_7_25_groupi_n_2379 ,in3[5]);
  and csa_tree_add_7_25_groupi_g18664(csa_tree_add_7_25_groupi_n_2533 ,in3[5] ,csa_tree_add_7_25_groupi_n_2379);
  and csa_tree_add_7_25_groupi_g18665(csa_tree_add_7_25_groupi_n_2531 ,in3[11] ,csa_tree_add_7_25_groupi_n_2376);
  or csa_tree_add_7_25_groupi_g18666(csa_tree_add_7_25_groupi_n_2529 ,csa_tree_add_7_25_groupi_n_2376 ,in3[11]);
  and csa_tree_add_7_25_groupi_g18667(csa_tree_add_7_25_groupi_n_2527 ,in3[8] ,csa_tree_add_7_25_groupi_n_2374);
  or csa_tree_add_7_25_groupi_g18668(csa_tree_add_7_25_groupi_n_2525 ,csa_tree_add_7_25_groupi_n_2374 ,in3[8]);
  or csa_tree_add_7_25_groupi_g18669(csa_tree_add_7_25_groupi_n_2523 ,csa_tree_add_7_25_groupi_n_2378 ,in3[29]);
  and csa_tree_add_7_25_groupi_g18670(csa_tree_add_7_25_groupi_n_2520 ,in3[1] ,csa_tree_add_7_25_groupi_n_2409);
  nor csa_tree_add_7_25_groupi_g18671(csa_tree_add_7_25_groupi_n_2474 ,in1[17] ,in1[16]);
  nor csa_tree_add_7_25_groupi_g18672(csa_tree_add_7_25_groupi_n_2473 ,in1[24] ,in1[23]);
  or csa_tree_add_7_25_groupi_g18673(csa_tree_add_7_25_groupi_n_2472 ,in3[11] ,in2[9]);
  and csa_tree_add_7_25_groupi_g18674(csa_tree_add_7_25_groupi_n_2471 ,in3[20] ,in2[18]);
  nor csa_tree_add_7_25_groupi_g18675(csa_tree_add_7_25_groupi_n_2470 ,in1[4] ,in1[3]);
  nor csa_tree_add_7_25_groupi_g18676(csa_tree_add_7_25_groupi_n_2469 ,in1[19] ,in1[18]);
  or csa_tree_add_7_25_groupi_g18677(csa_tree_add_7_25_groupi_n_2468 ,csa_tree_add_7_25_groupi_n_38 ,csa_tree_add_7_25_groupi_n_102);
  or csa_tree_add_7_25_groupi_g18678(csa_tree_add_7_25_groupi_n_2467 ,csa_tree_add_7_25_groupi_n_215 ,csa_tree_add_7_25_groupi_n_233);
  or csa_tree_add_7_25_groupi_g18679(csa_tree_add_7_25_groupi_n_2466 ,csa_tree_add_7_25_groupi_n_602 ,csa_tree_add_7_25_groupi_n_605);
  or csa_tree_add_7_25_groupi_g18680(csa_tree_add_7_25_groupi_n_2465 ,csa_tree_add_7_25_groupi_n_68 ,csa_tree_add_7_25_groupi_n_70);
  nor csa_tree_add_7_25_groupi_g18681(csa_tree_add_7_25_groupi_n_2464 ,in1[31] ,in1[30]);
  or csa_tree_add_7_25_groupi_g18682(csa_tree_add_7_25_groupi_n_2463 ,csa_tree_add_7_25_groupi_n_52 ,csa_tree_add_7_25_groupi_n_80);
  or csa_tree_add_7_25_groupi_g18683(csa_tree_add_7_25_groupi_n_2462 ,in3[5] ,in2[3]);
  or csa_tree_add_7_25_groupi_g18684(csa_tree_add_7_25_groupi_n_2461 ,csa_tree_add_7_25_groupi_n_64 ,csa_tree_add_7_25_groupi_n_239);
  or csa_tree_add_7_25_groupi_g18685(csa_tree_add_7_25_groupi_n_2460 ,csa_tree_add_7_25_groupi_n_12 ,csa_tree_add_7_25_groupi_n_56);
  or csa_tree_add_7_25_groupi_g18686(csa_tree_add_7_25_groupi_n_2459 ,in3[20] ,in2[18]);
  or csa_tree_add_7_25_groupi_g18687(csa_tree_add_7_25_groupi_n_2458 ,in3[8] ,in2[6]);
  nor csa_tree_add_7_25_groupi_g18688(csa_tree_add_7_25_groupi_n_2457 ,in1[18] ,in1[17]);
  or csa_tree_add_7_25_groupi_g18689(csa_tree_add_7_25_groupi_n_2456 ,csa_tree_add_7_25_groupi_n_48 ,csa_tree_add_7_25_groupi_n_60);
  and csa_tree_add_7_25_groupi_g18690(csa_tree_add_7_25_groupi_n_2455 ,in3[14] ,in2[12]);
  and csa_tree_add_7_25_groupi_g18691(csa_tree_add_7_25_groupi_n_2454 ,in3[8] ,in2[6]);
  or csa_tree_add_7_25_groupi_g18692(csa_tree_add_7_25_groupi_n_2453 ,csa_tree_add_7_25_groupi_n_24 ,csa_tree_add_7_25_groupi_n_76);
  nor csa_tree_add_7_25_groupi_g18693(csa_tree_add_7_25_groupi_n_2452 ,in1[25] ,in1[24]);
  nor csa_tree_add_7_25_groupi_g18694(csa_tree_add_7_25_groupi_n_2451 ,in1[9] ,in1[8]);
  or csa_tree_add_7_25_groupi_g18695(csa_tree_add_7_25_groupi_n_2450 ,in3[29] ,in2[27]);
  or csa_tree_add_7_25_groupi_g18696(csa_tree_add_7_25_groupi_n_2449 ,csa_tree_add_7_25_groupi_n_230 ,csa_tree_add_7_25_groupi_n_227);
  nor csa_tree_add_7_25_groupi_g18697(csa_tree_add_7_25_groupi_n_2448 ,in1[15] ,in1[14]);
  nor csa_tree_add_7_25_groupi_g18698(csa_tree_add_7_25_groupi_n_2447 ,in1[27] ,in1[26]);
  and csa_tree_add_7_25_groupi_g18699(csa_tree_add_7_25_groupi_n_2446 ,in3[11] ,in2[9]);
  nor csa_tree_add_7_25_groupi_g18700(csa_tree_add_7_25_groupi_n_2445 ,in1[23] ,in1[22]);
  nor csa_tree_add_7_25_groupi_g18701(csa_tree_add_7_25_groupi_n_2444 ,in1[8] ,in1[7]);
  or csa_tree_add_7_25_groupi_g18702(csa_tree_add_7_25_groupi_n_2443 ,csa_tree_add_7_25_groupi_n_108 ,csa_tree_add_7_25_groupi_n_8);
  and csa_tree_add_7_25_groupi_g18703(csa_tree_add_7_25_groupi_n_2442 ,in3[5] ,in2[3]);
  nor csa_tree_add_7_25_groupi_g18704(csa_tree_add_7_25_groupi_n_2441 ,in1[29] ,in1[28]);
  or csa_tree_add_7_25_groupi_g18705(csa_tree_add_7_25_groupi_n_2440 ,csa_tree_add_7_25_groupi_n_569 ,csa_tree_add_7_25_groupi_n_587);
  or csa_tree_add_7_25_groupi_g18706(csa_tree_add_7_25_groupi_n_2439 ,csa_tree_add_7_25_groupi_n_593 ,csa_tree_add_7_25_groupi_n_596);
  nor csa_tree_add_7_25_groupi_g18707(csa_tree_add_7_25_groupi_n_2438 ,in1[10] ,in1[9]);
  and csa_tree_add_7_25_groupi_g18708(csa_tree_add_7_25_groupi_n_2437 ,in3[26] ,in2[24]);
  nor csa_tree_add_7_25_groupi_g18709(csa_tree_add_7_25_groupi_n_2436 ,in1[26] ,in1[25]);
  or csa_tree_add_7_25_groupi_g18710(csa_tree_add_7_25_groupi_n_2435 ,csa_tree_add_7_25_groupi_n_40 ,csa_tree_add_7_25_groupi_n_18);
  nor csa_tree_add_7_25_groupi_g18711(csa_tree_add_7_25_groupi_n_2434 ,in1[3] ,in1[2]);
  or csa_tree_add_7_25_groupi_g18712(csa_tree_add_7_25_groupi_n_2433 ,csa_tree_add_7_25_groupi_n_221 ,csa_tree_add_7_25_groupi_n_236);
  or csa_tree_add_7_25_groupi_g18713(csa_tree_add_7_25_groupi_n_2432 ,csa_tree_add_7_25_groupi_n_66 ,csa_tree_add_7_25_groupi_n_104);
  and csa_tree_add_7_25_groupi_g18714(csa_tree_add_7_25_groupi_n_2431 ,in3[29] ,in2[27]);
  or csa_tree_add_7_25_groupi_g18715(csa_tree_add_7_25_groupi_n_2430 ,csa_tree_add_7_25_groupi_n_32 ,csa_tree_add_7_25_groupi_n_58);
  or csa_tree_add_7_25_groupi_g18716(csa_tree_add_7_25_groupi_n_2429 ,csa_tree_add_7_25_groupi_n_218 ,csa_tree_add_7_25_groupi_n_539);
  or csa_tree_add_7_25_groupi_g18717(csa_tree_add_7_25_groupi_n_2428 ,csa_tree_add_7_25_groupi_n_566 ,csa_tree_add_7_25_groupi_n_572);
  or csa_tree_add_7_25_groupi_g18718(csa_tree_add_7_25_groupi_n_2427 ,in3[17] ,in2[15]);
  or csa_tree_add_7_25_groupi_g18719(csa_tree_add_7_25_groupi_n_2426 ,csa_tree_add_7_25_groupi_n_557 ,csa_tree_add_7_25_groupi_n_563);
  and csa_tree_add_7_25_groupi_g18720(csa_tree_add_7_25_groupi_n_2425 ,in3[17] ,in2[15]);
  or csa_tree_add_7_25_groupi_g18721(csa_tree_add_7_25_groupi_n_2424 ,csa_tree_add_7_25_groupi_n_20 ,csa_tree_add_7_25_groupi_n_24);
  or csa_tree_add_7_25_groupi_g18722(csa_tree_add_7_25_groupi_n_2423 ,csa_tree_add_7_25_groupi_n_36 ,csa_tree_add_7_25_groupi_n_106);
  nor csa_tree_add_7_25_groupi_g18723(csa_tree_add_7_25_groupi_n_2422 ,in1[13] ,in1[12]);
  nor csa_tree_add_7_25_groupi_g18724(csa_tree_add_7_25_groupi_n_2421 ,in1[12] ,in1[11]);
  or csa_tree_add_7_25_groupi_g18725(csa_tree_add_7_25_groupi_n_2420 ,csa_tree_add_7_25_groupi_n_14 ,csa_tree_add_7_25_groupi_n_34);
  or csa_tree_add_7_25_groupi_g18726(csa_tree_add_7_25_groupi_n_2419 ,in3[14] ,in2[12]);
  or csa_tree_add_7_25_groupi_g18727(csa_tree_add_7_25_groupi_n_2418 ,in3[26] ,in2[24]);
  nor csa_tree_add_7_25_groupi_g18728(csa_tree_add_7_25_groupi_n_2417 ,in1[6] ,in1[5]);
  or csa_tree_add_7_25_groupi_g18729(csa_tree_add_7_25_groupi_n_2416 ,csa_tree_add_7_25_groupi_n_16 ,csa_tree_add_7_25_groupi_n_10);
  or csa_tree_add_7_25_groupi_g18730(csa_tree_add_7_25_groupi_n_2415 ,csa_tree_add_7_25_groupi_n_540 ,csa_tree_add_7_25_groupi_n_560);
  or csa_tree_add_7_25_groupi_g18731(csa_tree_add_7_25_groupi_n_2475 ,csa_tree_add_7_25_groupi_n_22 ,csa_tree_add_7_25_groupi_n_546);
  not csa_tree_add_7_25_groupi_g18732(csa_tree_add_7_25_groupi_n_2414 ,in3[13]);
  not csa_tree_add_7_25_groupi_g18733(csa_tree_add_7_25_groupi_n_2413 ,in2[4]);
  not csa_tree_add_7_25_groupi_g18734(csa_tree_add_7_25_groupi_n_2412 ,in2[31]);
  not csa_tree_add_7_25_groupi_g18735(csa_tree_add_7_25_groupi_n_2411 ,in3[22]);
  not csa_tree_add_7_25_groupi_g18736(csa_tree_add_7_25_groupi_n_2410 ,in3[16]);
  not csa_tree_add_7_25_groupi_g18737(csa_tree_add_7_25_groupi_n_2409 ,in3[0]);
  not csa_tree_add_7_25_groupi_g18738(csa_tree_add_7_25_groupi_n_2408 ,in3[30]);
  not csa_tree_add_7_25_groupi_g18739(csa_tree_add_7_25_groupi_n_2407 ,in3[6]);
  not csa_tree_add_7_25_groupi_g18740(csa_tree_add_7_25_groupi_n_2406 ,in3[3]);
  not csa_tree_add_7_25_groupi_g18741(csa_tree_add_7_25_groupi_n_2405 ,in3[24]);
  not csa_tree_add_7_25_groupi_g18742(csa_tree_add_7_25_groupi_n_2404 ,in3[12]);
  not csa_tree_add_7_25_groupi_g18743(csa_tree_add_7_25_groupi_n_2403 ,in1[31]);
  not csa_tree_add_7_25_groupi_g18744(csa_tree_add_7_25_groupi_n_2402 ,in1[28]);
  not csa_tree_add_7_25_groupi_g18745(csa_tree_add_7_25_groupi_n_2401 ,in1[27]);
  not csa_tree_add_7_25_groupi_g18746(csa_tree_add_7_25_groupi_n_2400 ,in1[26]);
  not csa_tree_add_7_25_groupi_g18747(csa_tree_add_7_25_groupi_n_2399 ,in1[25]);
  not csa_tree_add_7_25_groupi_g18748(csa_tree_add_7_25_groupi_n_2398 ,in1[24]);
  not csa_tree_add_7_25_groupi_g18749(csa_tree_add_7_25_groupi_n_2397 ,in1[23]);
  not csa_tree_add_7_25_groupi_g18750(csa_tree_add_7_25_groupi_n_2396 ,in1[20]);
  not csa_tree_add_7_25_groupi_g18751(csa_tree_add_7_25_groupi_n_2395 ,in1[17]);
  not csa_tree_add_7_25_groupi_g18752(csa_tree_add_7_25_groupi_n_2394 ,in1[16]);
  not csa_tree_add_7_25_groupi_g18753(csa_tree_add_7_25_groupi_n_2393 ,in1[12]);
  not csa_tree_add_7_25_groupi_g18754(csa_tree_add_7_25_groupi_n_2392 ,in1[4]);
  not csa_tree_add_7_25_groupi_g18755(csa_tree_add_7_25_groupi_n_2391 ,in1[5]);
  not csa_tree_add_7_25_groupi_g18756(csa_tree_add_7_25_groupi_n_2390 ,in1[10]);
  not csa_tree_add_7_25_groupi_g18757(csa_tree_add_7_25_groupi_n_2389 ,in1[8]);
  not csa_tree_add_7_25_groupi_g18758(csa_tree_add_7_25_groupi_n_2388 ,in1[2]);
  not csa_tree_add_7_25_groupi_g18759(csa_tree_add_7_25_groupi_n_2387 ,in1[13]);
  not csa_tree_add_7_25_groupi_g18760(csa_tree_add_7_25_groupi_n_2386 ,in1[3]);
  not csa_tree_add_7_25_groupi_g18761(csa_tree_add_7_25_groupi_n_2385 ,in3[29]);
  not csa_tree_add_7_25_groupi_g18762(csa_tree_add_7_25_groupi_n_2384 ,in3[26]);
  not csa_tree_add_7_25_groupi_g18763(csa_tree_add_7_25_groupi_n_2383 ,in3[2]);
  not csa_tree_add_7_25_groupi_g18764(csa_tree_add_7_25_groupi_n_2382 ,in3[8]);
  not csa_tree_add_7_25_groupi_g18765(csa_tree_add_7_25_groupi_n_2381 ,in3[5]);
  not csa_tree_add_7_25_groupi_g18766(csa_tree_add_7_25_groupi_n_2380 ,in2[30]);
  not csa_tree_add_7_25_groupi_g18767(csa_tree_add_7_25_groupi_n_2379 ,in3[4]);
  not csa_tree_add_7_25_groupi_g18768(csa_tree_add_7_25_groupi_n_2378 ,in3[28]);
  not csa_tree_add_7_25_groupi_g18769(csa_tree_add_7_25_groupi_n_2377 ,in3[19]);
  not csa_tree_add_7_25_groupi_g18770(csa_tree_add_7_25_groupi_n_2376 ,in3[10]);
  not csa_tree_add_7_25_groupi_g18771(csa_tree_add_7_25_groupi_n_2375 ,in3[25]);
  not csa_tree_add_7_25_groupi_g18772(csa_tree_add_7_25_groupi_n_2374 ,in3[7]);
  not csa_tree_add_7_25_groupi_g18773(csa_tree_add_7_25_groupi_n_2373 ,in3[31]);
  not csa_tree_add_7_25_groupi_g18774(csa_tree_add_7_25_groupi_n_2372 ,in3[21]);
  not csa_tree_add_7_25_groupi_g18775(csa_tree_add_7_25_groupi_n_2371 ,in3[9]);
  not csa_tree_add_7_25_groupi_g18776(csa_tree_add_7_25_groupi_n_2370 ,in3[27]);
  not csa_tree_add_7_25_groupi_g18777(csa_tree_add_7_25_groupi_n_2369 ,in3[18]);
  not csa_tree_add_7_25_groupi_g18778(csa_tree_add_7_25_groupi_n_2368 ,in3[15]);
  not csa_tree_add_7_25_groupi_g18779(csa_tree_add_7_25_groupi_n_2367 ,in1[30]);
  not csa_tree_add_7_25_groupi_g18780(csa_tree_add_7_25_groupi_n_2366 ,in1[29]);
  not csa_tree_add_7_25_groupi_g18781(csa_tree_add_7_25_groupi_n_2365 ,in1[22]);
  not csa_tree_add_7_25_groupi_g18782(csa_tree_add_7_25_groupi_n_2364 ,in1[21]);
  not csa_tree_add_7_25_groupi_g18783(csa_tree_add_7_25_groupi_n_2363 ,in1[19]);
  not csa_tree_add_7_25_groupi_g18784(csa_tree_add_7_25_groupi_n_2362 ,in1[0]);
  not csa_tree_add_7_25_groupi_g18785(csa_tree_add_7_25_groupi_n_2361 ,in1[18]);
  not csa_tree_add_7_25_groupi_g18786(csa_tree_add_7_25_groupi_n_2360 ,in1[1]);
  not csa_tree_add_7_25_groupi_g18787(csa_tree_add_7_25_groupi_n_2359 ,in1[15]);
  not csa_tree_add_7_25_groupi_g18788(csa_tree_add_7_25_groupi_n_2358 ,in1[14]);
  not csa_tree_add_7_25_groupi_g18789(csa_tree_add_7_25_groupi_n_2357 ,in1[9]);
  not csa_tree_add_7_25_groupi_g18790(csa_tree_add_7_25_groupi_n_2356 ,in1[7]);
  not csa_tree_add_7_25_groupi_g18791(csa_tree_add_7_25_groupi_n_2355 ,in1[11]);
  not csa_tree_add_7_25_groupi_g18792(csa_tree_add_7_25_groupi_n_2354 ,in1[6]);
  not csa_tree_add_7_25_groupi_g18793(csa_tree_add_7_25_groupi_n_2353 ,in3[23]);
  not csa_tree_add_7_25_groupi_g18794(csa_tree_add_7_25_groupi_n_2352 ,in3[20]);
  not csa_tree_add_7_25_groupi_g18795(csa_tree_add_7_25_groupi_n_2351 ,in3[17]);
  not csa_tree_add_7_25_groupi_g18796(csa_tree_add_7_25_groupi_n_2350 ,in3[14]);
  not csa_tree_add_7_25_groupi_g18797(csa_tree_add_7_25_groupi_n_2349 ,in3[11]);
  not csa_tree_add_7_25_groupi_drc_bufs(csa_tree_add_7_25_groupi_n_2313 ,csa_tree_add_7_25_groupi_n_1195);
  not csa_tree_add_7_25_groupi_drc_bufs18798(csa_tree_add_7_25_groupi_n_2312 ,csa_tree_add_7_25_groupi_n_1196);
  not csa_tree_add_7_25_groupi_drc_bufs18799(csa_tree_add_7_25_groupi_n_2311 ,csa_tree_add_7_25_groupi_n_1195);
  not csa_tree_add_7_25_groupi_drc_bufs18800(csa_tree_add_7_25_groupi_n_2310 ,csa_tree_add_7_25_groupi_n_1196);
  not csa_tree_add_7_25_groupi_drc_bufs18805(csa_tree_add_7_25_groupi_n_2309 ,csa_tree_add_7_25_groupi_n_1169);
  not csa_tree_add_7_25_groupi_drc_bufs18806(csa_tree_add_7_25_groupi_n_2308 ,csa_tree_add_7_25_groupi_n_1170);
  not csa_tree_add_7_25_groupi_drc_bufs18807(csa_tree_add_7_25_groupi_n_2307 ,csa_tree_add_7_25_groupi_n_1169);
  not csa_tree_add_7_25_groupi_drc_bufs18808(csa_tree_add_7_25_groupi_n_2306 ,csa_tree_add_7_25_groupi_n_1170);
  not csa_tree_add_7_25_groupi_drc_bufs18813(csa_tree_add_7_25_groupi_n_2305 ,csa_tree_add_7_25_groupi_n_1171);
  not csa_tree_add_7_25_groupi_drc_bufs18814(csa_tree_add_7_25_groupi_n_2304 ,csa_tree_add_7_25_groupi_n_1172);
  not csa_tree_add_7_25_groupi_drc_bufs18815(csa_tree_add_7_25_groupi_n_2303 ,csa_tree_add_7_25_groupi_n_1171);
  not csa_tree_add_7_25_groupi_drc_bufs18816(csa_tree_add_7_25_groupi_n_2302 ,csa_tree_add_7_25_groupi_n_1172);
  not csa_tree_add_7_25_groupi_drc_bufs18821(csa_tree_add_7_25_groupi_n_2301 ,csa_tree_add_7_25_groupi_n_1219);
  not csa_tree_add_7_25_groupi_drc_bufs18822(csa_tree_add_7_25_groupi_n_2300 ,csa_tree_add_7_25_groupi_n_1220);
  not csa_tree_add_7_25_groupi_drc_bufs18823(csa_tree_add_7_25_groupi_n_2299 ,csa_tree_add_7_25_groupi_n_1219);
  not csa_tree_add_7_25_groupi_drc_bufs18824(csa_tree_add_7_25_groupi_n_2298 ,csa_tree_add_7_25_groupi_n_1220);
  not csa_tree_add_7_25_groupi_drc_bufs18829(csa_tree_add_7_25_groupi_n_2297 ,csa_tree_add_7_25_groupi_n_1201);
  not csa_tree_add_7_25_groupi_drc_bufs18830(csa_tree_add_7_25_groupi_n_2296 ,csa_tree_add_7_25_groupi_n_1202);
  not csa_tree_add_7_25_groupi_drc_bufs18831(csa_tree_add_7_25_groupi_n_2295 ,csa_tree_add_7_25_groupi_n_1201);
  not csa_tree_add_7_25_groupi_drc_bufs18832(csa_tree_add_7_25_groupi_n_2294 ,csa_tree_add_7_25_groupi_n_1202);
  not csa_tree_add_7_25_groupi_drc_bufs18837(csa_tree_add_7_25_groupi_n_2293 ,csa_tree_add_7_25_groupi_n_1187);
  not csa_tree_add_7_25_groupi_drc_bufs18838(csa_tree_add_7_25_groupi_n_2292 ,csa_tree_add_7_25_groupi_n_1188);
  not csa_tree_add_7_25_groupi_drc_bufs18839(csa_tree_add_7_25_groupi_n_2291 ,csa_tree_add_7_25_groupi_n_1187);
  not csa_tree_add_7_25_groupi_drc_bufs18840(csa_tree_add_7_25_groupi_n_2290 ,csa_tree_add_7_25_groupi_n_1188);
  not csa_tree_add_7_25_groupi_drc_bufs18845(csa_tree_add_7_25_groupi_n_2289 ,csa_tree_add_7_25_groupi_n_1213);
  not csa_tree_add_7_25_groupi_drc_bufs18846(csa_tree_add_7_25_groupi_n_2288 ,csa_tree_add_7_25_groupi_n_1214);
  not csa_tree_add_7_25_groupi_drc_bufs18847(csa_tree_add_7_25_groupi_n_2287 ,csa_tree_add_7_25_groupi_n_1213);
  not csa_tree_add_7_25_groupi_drc_bufs18848(csa_tree_add_7_25_groupi_n_2286 ,csa_tree_add_7_25_groupi_n_1214);
  not csa_tree_add_7_25_groupi_drc_bufs18853(csa_tree_add_7_25_groupi_n_2285 ,csa_tree_add_7_25_groupi_n_1215);
  not csa_tree_add_7_25_groupi_drc_bufs18854(csa_tree_add_7_25_groupi_n_2284 ,csa_tree_add_7_25_groupi_n_1216);
  not csa_tree_add_7_25_groupi_drc_bufs18855(csa_tree_add_7_25_groupi_n_2283 ,csa_tree_add_7_25_groupi_n_1215);
  not csa_tree_add_7_25_groupi_drc_bufs18856(csa_tree_add_7_25_groupi_n_2282 ,csa_tree_add_7_25_groupi_n_1216);
  not csa_tree_add_7_25_groupi_drc_bufs18861(csa_tree_add_7_25_groupi_n_2281 ,csa_tree_add_7_25_groupi_n_1207);
  not csa_tree_add_7_25_groupi_drc_bufs18862(csa_tree_add_7_25_groupi_n_2280 ,csa_tree_add_7_25_groupi_n_1208);
  not csa_tree_add_7_25_groupi_drc_bufs18863(csa_tree_add_7_25_groupi_n_2279 ,csa_tree_add_7_25_groupi_n_1207);
  not csa_tree_add_7_25_groupi_drc_bufs18864(csa_tree_add_7_25_groupi_n_2278 ,csa_tree_add_7_25_groupi_n_1208);
  not csa_tree_add_7_25_groupi_drc_bufs18869(csa_tree_add_7_25_groupi_n_2277 ,csa_tree_add_7_25_groupi_n_1203);
  not csa_tree_add_7_25_groupi_drc_bufs18870(csa_tree_add_7_25_groupi_n_2276 ,csa_tree_add_7_25_groupi_n_1204);
  not csa_tree_add_7_25_groupi_drc_bufs18871(csa_tree_add_7_25_groupi_n_2275 ,csa_tree_add_7_25_groupi_n_1203);
  not csa_tree_add_7_25_groupi_drc_bufs18872(csa_tree_add_7_25_groupi_n_2274 ,csa_tree_add_7_25_groupi_n_1204);
  not csa_tree_add_7_25_groupi_drc_bufs18877(csa_tree_add_7_25_groupi_n_2273 ,csa_tree_add_7_25_groupi_n_1185);
  not csa_tree_add_7_25_groupi_drc_bufs18878(csa_tree_add_7_25_groupi_n_2272 ,csa_tree_add_7_25_groupi_n_1186);
  not csa_tree_add_7_25_groupi_drc_bufs18879(csa_tree_add_7_25_groupi_n_2271 ,csa_tree_add_7_25_groupi_n_1185);
  not csa_tree_add_7_25_groupi_drc_bufs18880(csa_tree_add_7_25_groupi_n_2270 ,csa_tree_add_7_25_groupi_n_1186);
  not csa_tree_add_7_25_groupi_drc_bufs18885(csa_tree_add_7_25_groupi_n_2269 ,csa_tree_add_7_25_groupi_n_1199);
  not csa_tree_add_7_25_groupi_drc_bufs18886(csa_tree_add_7_25_groupi_n_2268 ,csa_tree_add_7_25_groupi_n_1200);
  not csa_tree_add_7_25_groupi_drc_bufs18887(csa_tree_add_7_25_groupi_n_2267 ,csa_tree_add_7_25_groupi_n_1199);
  not csa_tree_add_7_25_groupi_drc_bufs18888(csa_tree_add_7_25_groupi_n_2266 ,csa_tree_add_7_25_groupi_n_1200);
  not csa_tree_add_7_25_groupi_drc_bufs18893(csa_tree_add_7_25_groupi_n_2265 ,csa_tree_add_7_25_groupi_n_1183);
  not csa_tree_add_7_25_groupi_drc_bufs18894(csa_tree_add_7_25_groupi_n_2264 ,csa_tree_add_7_25_groupi_n_1184);
  not csa_tree_add_7_25_groupi_drc_bufs18895(csa_tree_add_7_25_groupi_n_2263 ,csa_tree_add_7_25_groupi_n_1183);
  not csa_tree_add_7_25_groupi_drc_bufs18896(csa_tree_add_7_25_groupi_n_2262 ,csa_tree_add_7_25_groupi_n_1184);
  not csa_tree_add_7_25_groupi_drc_bufs18901(csa_tree_add_7_25_groupi_n_2261 ,csa_tree_add_7_25_groupi_n_1191);
  not csa_tree_add_7_25_groupi_drc_bufs18902(csa_tree_add_7_25_groupi_n_2260 ,csa_tree_add_7_25_groupi_n_1192);
  not csa_tree_add_7_25_groupi_drc_bufs18903(csa_tree_add_7_25_groupi_n_2259 ,csa_tree_add_7_25_groupi_n_1191);
  not csa_tree_add_7_25_groupi_drc_bufs18904(csa_tree_add_7_25_groupi_n_2258 ,csa_tree_add_7_25_groupi_n_1192);
  not csa_tree_add_7_25_groupi_drc_bufs18909(csa_tree_add_7_25_groupi_n_2257 ,csa_tree_add_7_25_groupi_n_1223);
  not csa_tree_add_7_25_groupi_drc_bufs18910(csa_tree_add_7_25_groupi_n_2256 ,csa_tree_add_7_25_groupi_n_1224);
  not csa_tree_add_7_25_groupi_drc_bufs18911(csa_tree_add_7_25_groupi_n_2255 ,csa_tree_add_7_25_groupi_n_1223);
  not csa_tree_add_7_25_groupi_drc_bufs18912(csa_tree_add_7_25_groupi_n_2254 ,csa_tree_add_7_25_groupi_n_1224);
  not csa_tree_add_7_25_groupi_drc_bufs18917(csa_tree_add_7_25_groupi_n_2253 ,csa_tree_add_7_25_groupi_n_1217);
  not csa_tree_add_7_25_groupi_drc_bufs18918(csa_tree_add_7_25_groupi_n_2252 ,csa_tree_add_7_25_groupi_n_1218);
  not csa_tree_add_7_25_groupi_drc_bufs18919(csa_tree_add_7_25_groupi_n_2251 ,csa_tree_add_7_25_groupi_n_1217);
  not csa_tree_add_7_25_groupi_drc_bufs18920(csa_tree_add_7_25_groupi_n_2250 ,csa_tree_add_7_25_groupi_n_1218);
  not csa_tree_add_7_25_groupi_drc_bufs18925(csa_tree_add_7_25_groupi_n_2249 ,csa_tree_add_7_25_groupi_n_1221);
  not csa_tree_add_7_25_groupi_drc_bufs18926(csa_tree_add_7_25_groupi_n_2248 ,csa_tree_add_7_25_groupi_n_1222);
  not csa_tree_add_7_25_groupi_drc_bufs18927(csa_tree_add_7_25_groupi_n_2247 ,csa_tree_add_7_25_groupi_n_1221);
  not csa_tree_add_7_25_groupi_drc_bufs18928(csa_tree_add_7_25_groupi_n_2246 ,csa_tree_add_7_25_groupi_n_1222);
  not csa_tree_add_7_25_groupi_drc_bufs18933(csa_tree_add_7_25_groupi_n_2245 ,csa_tree_add_7_25_groupi_n_1209);
  not csa_tree_add_7_25_groupi_drc_bufs18934(csa_tree_add_7_25_groupi_n_2244 ,csa_tree_add_7_25_groupi_n_1210);
  not csa_tree_add_7_25_groupi_drc_bufs18935(csa_tree_add_7_25_groupi_n_2243 ,csa_tree_add_7_25_groupi_n_1209);
  not csa_tree_add_7_25_groupi_drc_bufs18936(csa_tree_add_7_25_groupi_n_2242 ,csa_tree_add_7_25_groupi_n_1210);
  not csa_tree_add_7_25_groupi_drc_bufs18941(csa_tree_add_7_25_groupi_n_2241 ,csa_tree_add_7_25_groupi_n_1205);
  not csa_tree_add_7_25_groupi_drc_bufs18942(csa_tree_add_7_25_groupi_n_2240 ,csa_tree_add_7_25_groupi_n_1206);
  not csa_tree_add_7_25_groupi_drc_bufs18943(csa_tree_add_7_25_groupi_n_2239 ,csa_tree_add_7_25_groupi_n_1205);
  not csa_tree_add_7_25_groupi_drc_bufs18944(csa_tree_add_7_25_groupi_n_2238 ,csa_tree_add_7_25_groupi_n_1206);
  not csa_tree_add_7_25_groupi_drc_bufs18949(csa_tree_add_7_25_groupi_n_2237 ,csa_tree_add_7_25_groupi_n_1175);
  not csa_tree_add_7_25_groupi_drc_bufs18950(csa_tree_add_7_25_groupi_n_2236 ,csa_tree_add_7_25_groupi_n_1176);
  not csa_tree_add_7_25_groupi_drc_bufs18951(csa_tree_add_7_25_groupi_n_2235 ,csa_tree_add_7_25_groupi_n_1175);
  not csa_tree_add_7_25_groupi_drc_bufs18952(csa_tree_add_7_25_groupi_n_2234 ,csa_tree_add_7_25_groupi_n_1176);
  not csa_tree_add_7_25_groupi_drc_bufs18957(csa_tree_add_7_25_groupi_n_2233 ,csa_tree_add_7_25_groupi_n_1211);
  not csa_tree_add_7_25_groupi_drc_bufs18958(csa_tree_add_7_25_groupi_n_2232 ,csa_tree_add_7_25_groupi_n_1212);
  not csa_tree_add_7_25_groupi_drc_bufs18959(csa_tree_add_7_25_groupi_n_2231 ,csa_tree_add_7_25_groupi_n_1211);
  not csa_tree_add_7_25_groupi_drc_bufs18960(csa_tree_add_7_25_groupi_n_2230 ,csa_tree_add_7_25_groupi_n_1212);
  not csa_tree_add_7_25_groupi_drc_bufs18965(csa_tree_add_7_25_groupi_n_2229 ,csa_tree_add_7_25_groupi_n_1167);
  not csa_tree_add_7_25_groupi_drc_bufs18966(csa_tree_add_7_25_groupi_n_2228 ,csa_tree_add_7_25_groupi_n_1168);
  not csa_tree_add_7_25_groupi_drc_bufs18967(csa_tree_add_7_25_groupi_n_2227 ,csa_tree_add_7_25_groupi_n_1167);
  not csa_tree_add_7_25_groupi_drc_bufs18968(csa_tree_add_7_25_groupi_n_2226 ,csa_tree_add_7_25_groupi_n_1168);
  not csa_tree_add_7_25_groupi_drc_bufs18973(csa_tree_add_7_25_groupi_n_2225 ,csa_tree_add_7_25_groupi_n_1189);
  not csa_tree_add_7_25_groupi_drc_bufs18974(csa_tree_add_7_25_groupi_n_2224 ,csa_tree_add_7_25_groupi_n_1190);
  not csa_tree_add_7_25_groupi_drc_bufs18975(csa_tree_add_7_25_groupi_n_2223 ,csa_tree_add_7_25_groupi_n_1189);
  not csa_tree_add_7_25_groupi_drc_bufs18976(csa_tree_add_7_25_groupi_n_2222 ,csa_tree_add_7_25_groupi_n_1190);
  not csa_tree_add_7_25_groupi_drc_bufs18981(csa_tree_add_7_25_groupi_n_2221 ,csa_tree_add_7_25_groupi_n_1179);
  not csa_tree_add_7_25_groupi_drc_bufs18982(csa_tree_add_7_25_groupi_n_2220 ,csa_tree_add_7_25_groupi_n_1180);
  not csa_tree_add_7_25_groupi_drc_bufs18983(csa_tree_add_7_25_groupi_n_2219 ,csa_tree_add_7_25_groupi_n_1179);
  not csa_tree_add_7_25_groupi_drc_bufs18984(csa_tree_add_7_25_groupi_n_2218 ,csa_tree_add_7_25_groupi_n_1180);
  not csa_tree_add_7_25_groupi_drc_bufs18989(csa_tree_add_7_25_groupi_n_2217 ,csa_tree_add_7_25_groupi_n_1181);
  not csa_tree_add_7_25_groupi_drc_bufs18990(csa_tree_add_7_25_groupi_n_2216 ,csa_tree_add_7_25_groupi_n_1182);
  not csa_tree_add_7_25_groupi_drc_bufs18991(csa_tree_add_7_25_groupi_n_2215 ,csa_tree_add_7_25_groupi_n_1181);
  not csa_tree_add_7_25_groupi_drc_bufs18992(csa_tree_add_7_25_groupi_n_2214 ,csa_tree_add_7_25_groupi_n_1182);
  not csa_tree_add_7_25_groupi_drc_bufs18997(csa_tree_add_7_25_groupi_n_2213 ,csa_tree_add_7_25_groupi_n_1177);
  not csa_tree_add_7_25_groupi_drc_bufs18998(csa_tree_add_7_25_groupi_n_2212 ,csa_tree_add_7_25_groupi_n_1178);
  not csa_tree_add_7_25_groupi_drc_bufs18999(csa_tree_add_7_25_groupi_n_2211 ,csa_tree_add_7_25_groupi_n_1177);
  not csa_tree_add_7_25_groupi_drc_bufs19000(csa_tree_add_7_25_groupi_n_2210 ,csa_tree_add_7_25_groupi_n_1178);
  not csa_tree_add_7_25_groupi_drc_bufs19005(csa_tree_add_7_25_groupi_n_2209 ,csa_tree_add_7_25_groupi_n_1197);
  not csa_tree_add_7_25_groupi_drc_bufs19006(csa_tree_add_7_25_groupi_n_2208 ,csa_tree_add_7_25_groupi_n_1198);
  not csa_tree_add_7_25_groupi_drc_bufs19007(csa_tree_add_7_25_groupi_n_2207 ,csa_tree_add_7_25_groupi_n_1197);
  not csa_tree_add_7_25_groupi_drc_bufs19008(csa_tree_add_7_25_groupi_n_2206 ,csa_tree_add_7_25_groupi_n_1198);
  not csa_tree_add_7_25_groupi_drc_bufs19013(csa_tree_add_7_25_groupi_n_2205 ,csa_tree_add_7_25_groupi_n_1173);
  not csa_tree_add_7_25_groupi_drc_bufs19014(csa_tree_add_7_25_groupi_n_2204 ,csa_tree_add_7_25_groupi_n_1174);
  not csa_tree_add_7_25_groupi_drc_bufs19015(csa_tree_add_7_25_groupi_n_2203 ,csa_tree_add_7_25_groupi_n_1173);
  not csa_tree_add_7_25_groupi_drc_bufs19016(csa_tree_add_7_25_groupi_n_2202 ,csa_tree_add_7_25_groupi_n_1174);
  not csa_tree_add_7_25_groupi_drc_bufs19021(csa_tree_add_7_25_groupi_n_2201 ,csa_tree_add_7_25_groupi_n_1193);
  not csa_tree_add_7_25_groupi_drc_bufs19022(csa_tree_add_7_25_groupi_n_2200 ,csa_tree_add_7_25_groupi_n_1194);
  not csa_tree_add_7_25_groupi_drc_bufs19023(csa_tree_add_7_25_groupi_n_2199 ,csa_tree_add_7_25_groupi_n_1193);
  not csa_tree_add_7_25_groupi_drc_bufs19024(csa_tree_add_7_25_groupi_n_2198 ,csa_tree_add_7_25_groupi_n_1194);
  not csa_tree_add_7_25_groupi_drc_bufs19787(csa_tree_add_7_25_groupi_n_2197 ,csa_tree_add_7_25_groupi_n_2196);
  not csa_tree_add_7_25_groupi_drc_bufs19788(csa_tree_add_7_25_groupi_n_2196 ,csa_tree_add_7_25_groupi_n_2792);
  not csa_tree_add_7_25_groupi_drc_bufs19791(csa_tree_add_7_25_groupi_n_2195 ,csa_tree_add_7_25_groupi_n_2194);
  not csa_tree_add_7_25_groupi_drc_bufs19792(csa_tree_add_7_25_groupi_n_2194 ,csa_tree_add_7_25_groupi_n_3523);
  not csa_tree_add_7_25_groupi_drc_bufs19794(csa_tree_add_7_25_groupi_n_2193 ,csa_tree_add_7_25_groupi_n_2191);
  not csa_tree_add_7_25_groupi_drc_bufs19795(csa_tree_add_7_25_groupi_n_2192 ,csa_tree_add_7_25_groupi_n_2191);
  not csa_tree_add_7_25_groupi_drc_bufs19796(csa_tree_add_7_25_groupi_n_2191 ,csa_tree_add_7_25_groupi_n_2322);
  not csa_tree_add_7_25_groupi_drc_bufs19798(csa_tree_add_7_25_groupi_n_2190 ,csa_tree_add_7_25_groupi_n_2188);
  not csa_tree_add_7_25_groupi_drc_bufs19799(csa_tree_add_7_25_groupi_n_2189 ,csa_tree_add_7_25_groupi_n_2188);
  not csa_tree_add_7_25_groupi_drc_bufs19800(csa_tree_add_7_25_groupi_n_2188 ,csa_tree_add_7_25_groupi_n_2323);
  not csa_tree_add_7_25_groupi_drc_bufs19802(csa_tree_add_7_25_groupi_n_2187 ,csa_tree_add_7_25_groupi_n_2185);
  not csa_tree_add_7_25_groupi_drc_bufs19803(csa_tree_add_7_25_groupi_n_2186 ,csa_tree_add_7_25_groupi_n_2185);
  not csa_tree_add_7_25_groupi_drc_bufs19804(csa_tree_add_7_25_groupi_n_2185 ,csa_tree_add_7_25_groupi_n_2839);
  not csa_tree_add_7_25_groupi_drc_bufs19806(csa_tree_add_7_25_groupi_n_2184 ,csa_tree_add_7_25_groupi_n_2182);
  not csa_tree_add_7_25_groupi_drc_bufs19807(csa_tree_add_7_25_groupi_n_2183 ,csa_tree_add_7_25_groupi_n_2182);
  not csa_tree_add_7_25_groupi_drc_bufs19808(csa_tree_add_7_25_groupi_n_2182 ,csa_tree_add_7_25_groupi_n_2838);
  not csa_tree_add_7_25_groupi_drc_bufs19810(csa_tree_add_7_25_groupi_n_2181 ,csa_tree_add_7_25_groupi_n_2179);
  not csa_tree_add_7_25_groupi_drc_bufs19811(csa_tree_add_7_25_groupi_n_2180 ,csa_tree_add_7_25_groupi_n_2179);
  not csa_tree_add_7_25_groupi_drc_bufs19812(csa_tree_add_7_25_groupi_n_2179 ,csa_tree_add_7_25_groupi_n_2337);
  not csa_tree_add_7_25_groupi_drc_bufs19814(csa_tree_add_7_25_groupi_n_2178 ,csa_tree_add_7_25_groupi_n_2176);
  not csa_tree_add_7_25_groupi_drc_bufs19815(csa_tree_add_7_25_groupi_n_2177 ,csa_tree_add_7_25_groupi_n_2176);
  not csa_tree_add_7_25_groupi_drc_bufs19816(csa_tree_add_7_25_groupi_n_2176 ,csa_tree_add_7_25_groupi_n_2336);
  not csa_tree_add_7_25_groupi_drc_bufs19818(csa_tree_add_7_25_groupi_n_2175 ,csa_tree_add_7_25_groupi_n_2173);
  not csa_tree_add_7_25_groupi_drc_bufs19819(csa_tree_add_7_25_groupi_n_2174 ,csa_tree_add_7_25_groupi_n_2173);
  not csa_tree_add_7_25_groupi_drc_bufs19820(csa_tree_add_7_25_groupi_n_2173 ,csa_tree_add_7_25_groupi_n_2335);
  not csa_tree_add_7_25_groupi_drc_bufs19822(csa_tree_add_7_25_groupi_n_2172 ,csa_tree_add_7_25_groupi_n_2170);
  not csa_tree_add_7_25_groupi_drc_bufs19823(csa_tree_add_7_25_groupi_n_2171 ,csa_tree_add_7_25_groupi_n_2170);
  not csa_tree_add_7_25_groupi_drc_bufs19824(csa_tree_add_7_25_groupi_n_2170 ,csa_tree_add_7_25_groupi_n_2337);
  not csa_tree_add_7_25_groupi_drc_bufs19826(csa_tree_add_7_25_groupi_n_2169 ,csa_tree_add_7_25_groupi_n_2167);
  not csa_tree_add_7_25_groupi_drc_bufs19827(csa_tree_add_7_25_groupi_n_2168 ,csa_tree_add_7_25_groupi_n_2167);
  not csa_tree_add_7_25_groupi_drc_bufs19828(csa_tree_add_7_25_groupi_n_2167 ,csa_tree_add_7_25_groupi_n_2336);
  not csa_tree_add_7_25_groupi_drc_bufs19830(csa_tree_add_7_25_groupi_n_2166 ,csa_tree_add_7_25_groupi_n_2164);
  not csa_tree_add_7_25_groupi_drc_bufs19831(csa_tree_add_7_25_groupi_n_2165 ,csa_tree_add_7_25_groupi_n_2164);
  not csa_tree_add_7_25_groupi_drc_bufs19832(csa_tree_add_7_25_groupi_n_2164 ,csa_tree_add_7_25_groupi_n_2321);
  not csa_tree_add_7_25_groupi_drc_bufs19834(csa_tree_add_7_25_groupi_n_2163 ,csa_tree_add_7_25_groupi_n_2161);
  not csa_tree_add_7_25_groupi_drc_bufs19835(csa_tree_add_7_25_groupi_n_2162 ,csa_tree_add_7_25_groupi_n_2161);
  not csa_tree_add_7_25_groupi_drc_bufs19836(csa_tree_add_7_25_groupi_n_2161 ,csa_tree_add_7_25_groupi_n_2316);
  not csa_tree_add_7_25_groupi_drc_bufs19838(csa_tree_add_7_25_groupi_n_2160 ,csa_tree_add_7_25_groupi_n_2158);
  not csa_tree_add_7_25_groupi_drc_bufs19839(csa_tree_add_7_25_groupi_n_2159 ,csa_tree_add_7_25_groupi_n_2158);
  not csa_tree_add_7_25_groupi_drc_bufs19840(csa_tree_add_7_25_groupi_n_2158 ,csa_tree_add_7_25_groupi_n_2753);
  not csa_tree_add_7_25_groupi_drc_bufs19842(csa_tree_add_7_25_groupi_n_2157 ,csa_tree_add_7_25_groupi_n_2155);
  not csa_tree_add_7_25_groupi_drc_bufs19843(csa_tree_add_7_25_groupi_n_2156 ,csa_tree_add_7_25_groupi_n_2155);
  not csa_tree_add_7_25_groupi_drc_bufs19844(csa_tree_add_7_25_groupi_n_2155 ,csa_tree_add_7_25_groupi_n_2752);
  not csa_tree_add_7_25_groupi_drc_bufs19846(csa_tree_add_7_25_groupi_n_2154 ,csa_tree_add_7_25_groupi_n_2152);
  not csa_tree_add_7_25_groupi_drc_bufs19847(csa_tree_add_7_25_groupi_n_2153 ,csa_tree_add_7_25_groupi_n_2152);
  not csa_tree_add_7_25_groupi_drc_bufs19848(csa_tree_add_7_25_groupi_n_2152 ,csa_tree_add_7_25_groupi_n_2325);
  not csa_tree_add_7_25_groupi_drc_bufs19850(csa_tree_add_7_25_groupi_n_2151 ,csa_tree_add_7_25_groupi_n_2149);
  not csa_tree_add_7_25_groupi_drc_bufs19851(csa_tree_add_7_25_groupi_n_2150 ,csa_tree_add_7_25_groupi_n_2149);
  not csa_tree_add_7_25_groupi_drc_bufs19852(csa_tree_add_7_25_groupi_n_2149 ,csa_tree_add_7_25_groupi_n_2324);
  not csa_tree_add_7_25_groupi_drc_bufs19854(csa_tree_add_7_25_groupi_n_2148 ,csa_tree_add_7_25_groupi_n_2146);
  not csa_tree_add_7_25_groupi_drc_bufs19855(csa_tree_add_7_25_groupi_n_2147 ,csa_tree_add_7_25_groupi_n_2146);
  not csa_tree_add_7_25_groupi_drc_bufs19856(csa_tree_add_7_25_groupi_n_2146 ,csa_tree_add_7_25_groupi_n_2325);
  not csa_tree_add_7_25_groupi_drc_bufs19858(csa_tree_add_7_25_groupi_n_2145 ,csa_tree_add_7_25_groupi_n_2143);
  not csa_tree_add_7_25_groupi_drc_bufs19859(csa_tree_add_7_25_groupi_n_2144 ,csa_tree_add_7_25_groupi_n_2143);
  not csa_tree_add_7_25_groupi_drc_bufs19860(csa_tree_add_7_25_groupi_n_2143 ,csa_tree_add_7_25_groupi_n_2324);
  not csa_tree_add_7_25_groupi_drc_bufs19862(csa_tree_add_7_25_groupi_n_2142 ,csa_tree_add_7_25_groupi_n_2140);
  not csa_tree_add_7_25_groupi_drc_bufs19863(csa_tree_add_7_25_groupi_n_2141 ,csa_tree_add_7_25_groupi_n_2140);
  not csa_tree_add_7_25_groupi_drc_bufs19864(csa_tree_add_7_25_groupi_n_2140 ,csa_tree_add_7_25_groupi_n_2748);
  not csa_tree_add_7_25_groupi_drc_bufs19866(csa_tree_add_7_25_groupi_n_2139 ,csa_tree_add_7_25_groupi_n_2137);
  not csa_tree_add_7_25_groupi_drc_bufs19867(csa_tree_add_7_25_groupi_n_2138 ,csa_tree_add_7_25_groupi_n_2137);
  not csa_tree_add_7_25_groupi_drc_bufs19868(csa_tree_add_7_25_groupi_n_2137 ,csa_tree_add_7_25_groupi_n_2749);
  not csa_tree_add_7_25_groupi_drc_bufs19870(csa_tree_add_7_25_groupi_n_2136 ,csa_tree_add_7_25_groupi_n_2134);
  not csa_tree_add_7_25_groupi_drc_bufs19871(csa_tree_add_7_25_groupi_n_2135 ,csa_tree_add_7_25_groupi_n_2134);
  not csa_tree_add_7_25_groupi_drc_bufs19872(csa_tree_add_7_25_groupi_n_2134 ,csa_tree_add_7_25_groupi_n_2321);
  not csa_tree_add_7_25_groupi_drc_bufs19874(csa_tree_add_7_25_groupi_n_2133 ,csa_tree_add_7_25_groupi_n_2131);
  not csa_tree_add_7_25_groupi_drc_bufs19875(csa_tree_add_7_25_groupi_n_2132 ,csa_tree_add_7_25_groupi_n_2131);
  not csa_tree_add_7_25_groupi_drc_bufs19876(csa_tree_add_7_25_groupi_n_2131 ,csa_tree_add_7_25_groupi_n_2320);
  not csa_tree_add_7_25_groupi_drc_bufs19878(csa_tree_add_7_25_groupi_n_2130 ,csa_tree_add_7_25_groupi_n_2128);
  not csa_tree_add_7_25_groupi_drc_bufs19879(csa_tree_add_7_25_groupi_n_2129 ,csa_tree_add_7_25_groupi_n_2128);
  not csa_tree_add_7_25_groupi_drc_bufs19880(csa_tree_add_7_25_groupi_n_2128 ,csa_tree_add_7_25_groupi_n_2322);
  not csa_tree_add_7_25_groupi_drc_bufs19882(csa_tree_add_7_25_groupi_n_2127 ,csa_tree_add_7_25_groupi_n_2125);
  not csa_tree_add_7_25_groupi_drc_bufs19883(csa_tree_add_7_25_groupi_n_2126 ,csa_tree_add_7_25_groupi_n_2125);
  not csa_tree_add_7_25_groupi_drc_bufs19884(csa_tree_add_7_25_groupi_n_2125 ,csa_tree_add_7_25_groupi_n_2745);
  not csa_tree_add_7_25_groupi_drc_bufs19886(csa_tree_add_7_25_groupi_n_2124 ,csa_tree_add_7_25_groupi_n_2122);
  not csa_tree_add_7_25_groupi_drc_bufs19887(csa_tree_add_7_25_groupi_n_2123 ,csa_tree_add_7_25_groupi_n_2122);
  not csa_tree_add_7_25_groupi_drc_bufs19888(csa_tree_add_7_25_groupi_n_2122 ,csa_tree_add_7_25_groupi_n_2744);
  not csa_tree_add_7_25_groupi_drc_bufs19890(csa_tree_add_7_25_groupi_n_2121 ,csa_tree_add_7_25_groupi_n_2119);
  not csa_tree_add_7_25_groupi_drc_bufs19891(csa_tree_add_7_25_groupi_n_2120 ,csa_tree_add_7_25_groupi_n_2119);
  not csa_tree_add_7_25_groupi_drc_bufs19892(csa_tree_add_7_25_groupi_n_2119 ,csa_tree_add_7_25_groupi_n_2318);
  not csa_tree_add_7_25_groupi_drc_bufs19894(csa_tree_add_7_25_groupi_n_2118 ,csa_tree_add_7_25_groupi_n_2116);
  not csa_tree_add_7_25_groupi_drc_bufs19895(csa_tree_add_7_25_groupi_n_2117 ,csa_tree_add_7_25_groupi_n_2116);
  not csa_tree_add_7_25_groupi_drc_bufs19896(csa_tree_add_7_25_groupi_n_2116 ,csa_tree_add_7_25_groupi_n_2317);
  not csa_tree_add_7_25_groupi_drc_bufs19898(csa_tree_add_7_25_groupi_n_2115 ,csa_tree_add_7_25_groupi_n_2113);
  not csa_tree_add_7_25_groupi_drc_bufs19899(csa_tree_add_7_25_groupi_n_2114 ,csa_tree_add_7_25_groupi_n_2113);
  not csa_tree_add_7_25_groupi_drc_bufs19900(csa_tree_add_7_25_groupi_n_2113 ,csa_tree_add_7_25_groupi_n_2319);
  not csa_tree_add_7_25_groupi_drc_bufs19902(csa_tree_add_7_25_groupi_n_2112 ,csa_tree_add_7_25_groupi_n_2110);
  not csa_tree_add_7_25_groupi_drc_bufs19903(csa_tree_add_7_25_groupi_n_2111 ,csa_tree_add_7_25_groupi_n_2110);
  not csa_tree_add_7_25_groupi_drc_bufs19904(csa_tree_add_7_25_groupi_n_2110 ,csa_tree_add_7_25_groupi_n_2318);
  not csa_tree_add_7_25_groupi_drc_bufs19906(csa_tree_add_7_25_groupi_n_2109 ,csa_tree_add_7_25_groupi_n_2107);
  not csa_tree_add_7_25_groupi_drc_bufs19907(csa_tree_add_7_25_groupi_n_2108 ,csa_tree_add_7_25_groupi_n_2107);
  not csa_tree_add_7_25_groupi_drc_bufs19908(csa_tree_add_7_25_groupi_n_2107 ,csa_tree_add_7_25_groupi_n_2319);
  not csa_tree_add_7_25_groupi_drc_bufs19910(csa_tree_add_7_25_groupi_n_2106 ,csa_tree_add_7_25_groupi_n_2104);
  not csa_tree_add_7_25_groupi_drc_bufs19911(csa_tree_add_7_25_groupi_n_2105 ,csa_tree_add_7_25_groupi_n_2104);
  not csa_tree_add_7_25_groupi_drc_bufs19912(csa_tree_add_7_25_groupi_n_2104 ,csa_tree_add_7_25_groupi_n_2741);
  not csa_tree_add_7_25_groupi_drc_bufs19914(csa_tree_add_7_25_groupi_n_2103 ,csa_tree_add_7_25_groupi_n_2101);
  not csa_tree_add_7_25_groupi_drc_bufs19915(csa_tree_add_7_25_groupi_n_2102 ,csa_tree_add_7_25_groupi_n_2101);
  not csa_tree_add_7_25_groupi_drc_bufs19916(csa_tree_add_7_25_groupi_n_2101 ,csa_tree_add_7_25_groupi_n_2740);
  not csa_tree_add_7_25_groupi_drc_bufs19918(csa_tree_add_7_25_groupi_n_2100 ,csa_tree_add_7_25_groupi_n_2098);
  not csa_tree_add_7_25_groupi_drc_bufs19919(csa_tree_add_7_25_groupi_n_2099 ,csa_tree_add_7_25_groupi_n_2098);
  not csa_tree_add_7_25_groupi_drc_bufs19920(csa_tree_add_7_25_groupi_n_2098 ,csa_tree_add_7_25_groupi_n_2315);
  not csa_tree_add_7_25_groupi_drc_bufs19922(csa_tree_add_7_25_groupi_n_2097 ,csa_tree_add_7_25_groupi_n_2095);
  not csa_tree_add_7_25_groupi_drc_bufs19923(csa_tree_add_7_25_groupi_n_2096 ,csa_tree_add_7_25_groupi_n_2095);
  not csa_tree_add_7_25_groupi_drc_bufs19924(csa_tree_add_7_25_groupi_n_2095 ,csa_tree_add_7_25_groupi_n_2314);
  not csa_tree_add_7_25_groupi_drc_bufs19926(csa_tree_add_7_25_groupi_n_2094 ,csa_tree_add_7_25_groupi_n_2092);
  not csa_tree_add_7_25_groupi_drc_bufs19927(csa_tree_add_7_25_groupi_n_2093 ,csa_tree_add_7_25_groupi_n_2092);
  not csa_tree_add_7_25_groupi_drc_bufs19928(csa_tree_add_7_25_groupi_n_2092 ,csa_tree_add_7_25_groupi_n_2316);
  not csa_tree_add_7_25_groupi_drc_bufs19930(csa_tree_add_7_25_groupi_n_2091 ,csa_tree_add_7_25_groupi_n_2089);
  not csa_tree_add_7_25_groupi_drc_bufs19931(csa_tree_add_7_25_groupi_n_2090 ,csa_tree_add_7_25_groupi_n_2089);
  not csa_tree_add_7_25_groupi_drc_bufs19932(csa_tree_add_7_25_groupi_n_2089 ,csa_tree_add_7_25_groupi_n_2315);
  not csa_tree_add_7_25_groupi_drc_bufs19934(csa_tree_add_7_25_groupi_n_2088 ,csa_tree_add_7_25_groupi_n_2086);
  not csa_tree_add_7_25_groupi_drc_bufs19935(csa_tree_add_7_25_groupi_n_2087 ,csa_tree_add_7_25_groupi_n_2086);
  not csa_tree_add_7_25_groupi_drc_bufs19936(csa_tree_add_7_25_groupi_n_2086 ,csa_tree_add_7_25_groupi_n_2748);
  not csa_tree_add_7_25_groupi_drc_bufs19938(csa_tree_add_7_25_groupi_n_2085 ,csa_tree_add_7_25_groupi_n_2083);
  not csa_tree_add_7_25_groupi_drc_bufs19939(csa_tree_add_7_25_groupi_n_2084 ,csa_tree_add_7_25_groupi_n_2083);
  not csa_tree_add_7_25_groupi_drc_bufs19940(csa_tree_add_7_25_groupi_n_2083 ,csa_tree_add_7_25_groupi_n_2838);
  not csa_tree_add_7_25_groupi_drc_bufs19942(csa_tree_add_7_25_groupi_n_2082 ,csa_tree_add_7_25_groupi_n_2080);
  not csa_tree_add_7_25_groupi_drc_bufs19943(csa_tree_add_7_25_groupi_n_2081 ,csa_tree_add_7_25_groupi_n_2080);
  not csa_tree_add_7_25_groupi_drc_bufs19944(csa_tree_add_7_25_groupi_n_2080 ,csa_tree_add_7_25_groupi_n_2752);
  not csa_tree_add_7_25_groupi_drc_bufs19946(csa_tree_add_7_25_groupi_n_2079 ,csa_tree_add_7_25_groupi_n_2077);
  not csa_tree_add_7_25_groupi_drc_bufs19947(csa_tree_add_7_25_groupi_n_2078 ,csa_tree_add_7_25_groupi_n_2077);
  not csa_tree_add_7_25_groupi_drc_bufs19948(csa_tree_add_7_25_groupi_n_2077 ,csa_tree_add_7_25_groupi_n_2744);
  not csa_tree_add_7_25_groupi_drc_bufs19950(csa_tree_add_7_25_groupi_n_2076 ,csa_tree_add_7_25_groupi_n_2074);
  not csa_tree_add_7_25_groupi_drc_bufs19951(csa_tree_add_7_25_groupi_n_2075 ,csa_tree_add_7_25_groupi_n_2074);
  not csa_tree_add_7_25_groupi_drc_bufs19952(csa_tree_add_7_25_groupi_n_2074 ,csa_tree_add_7_25_groupi_n_2740);
  not csa_tree_add_7_25_groupi_drc_bufs19954(csa_tree_add_7_25_groupi_n_2073 ,csa_tree_add_7_25_groupi_n_2071);
  not csa_tree_add_7_25_groupi_drc_bufs19955(csa_tree_add_7_25_groupi_n_2072 ,csa_tree_add_7_25_groupi_n_2071);
  not csa_tree_add_7_25_groupi_drc_bufs19956(csa_tree_add_7_25_groupi_n_2071 ,csa_tree_add_7_25_groupi_n_2779);
  not csa_tree_add_7_25_groupi_drc_bufs19958(csa_tree_add_7_25_groupi_n_2070 ,csa_tree_add_7_25_groupi_n_2068);
  not csa_tree_add_7_25_groupi_drc_bufs19959(csa_tree_add_7_25_groupi_n_2069 ,csa_tree_add_7_25_groupi_n_2068);
  not csa_tree_add_7_25_groupi_drc_bufs19960(csa_tree_add_7_25_groupi_n_2068 ,csa_tree_add_7_25_groupi_n_2781);
  not csa_tree_add_7_25_groupi_drc_bufs19962(csa_tree_add_7_25_groupi_n_2067 ,csa_tree_add_7_25_groupi_n_2065);
  not csa_tree_add_7_25_groupi_drc_bufs19963(csa_tree_add_7_25_groupi_n_2066 ,csa_tree_add_7_25_groupi_n_2065);
  not csa_tree_add_7_25_groupi_drc_bufs19964(csa_tree_add_7_25_groupi_n_2065 ,csa_tree_add_7_25_groupi_n_2327);
  not csa_tree_add_7_25_groupi_drc_bufs19966(csa_tree_add_7_25_groupi_n_2064 ,csa_tree_add_7_25_groupi_n_2062);
  not csa_tree_add_7_25_groupi_drc_bufs19967(csa_tree_add_7_25_groupi_n_2063 ,csa_tree_add_7_25_groupi_n_2062);
  not csa_tree_add_7_25_groupi_drc_bufs19968(csa_tree_add_7_25_groupi_n_2062 ,csa_tree_add_7_25_groupi_n_2326);
  not csa_tree_add_7_25_groupi_drc_bufs19970(csa_tree_add_7_25_groupi_n_2061 ,csa_tree_add_7_25_groupi_n_2059);
  not csa_tree_add_7_25_groupi_drc_bufs19971(csa_tree_add_7_25_groupi_n_2060 ,csa_tree_add_7_25_groupi_n_2059);
  not csa_tree_add_7_25_groupi_drc_bufs19972(csa_tree_add_7_25_groupi_n_2059 ,csa_tree_add_7_25_groupi_n_2327);
  not csa_tree_add_7_25_groupi_drc_bufs19974(csa_tree_add_7_25_groupi_n_2058 ,csa_tree_add_7_25_groupi_n_2056);
  not csa_tree_add_7_25_groupi_drc_bufs19975(csa_tree_add_7_25_groupi_n_2057 ,csa_tree_add_7_25_groupi_n_2056);
  not csa_tree_add_7_25_groupi_drc_bufs19976(csa_tree_add_7_25_groupi_n_2056 ,csa_tree_add_7_25_groupi_n_2326);
  not csa_tree_add_7_25_groupi_drc_bufs19978(csa_tree_add_7_25_groupi_n_2055 ,csa_tree_add_7_25_groupi_n_2053);
  not csa_tree_add_7_25_groupi_drc_bufs19979(csa_tree_add_7_25_groupi_n_2054 ,csa_tree_add_7_25_groupi_n_2053);
  not csa_tree_add_7_25_groupi_drc_bufs19980(csa_tree_add_7_25_groupi_n_2053 ,csa_tree_add_7_25_groupi_n_2781);
  not csa_tree_add_7_25_groupi_drc_bufs20010(csa_tree_add_7_25_groupi_n_2052 ,csa_tree_add_7_25_groupi_n_2050);
  not csa_tree_add_7_25_groupi_drc_bufs20011(csa_tree_add_7_25_groupi_n_2051 ,csa_tree_add_7_25_groupi_n_2050);
  not csa_tree_add_7_25_groupi_drc_bufs20012(csa_tree_add_7_25_groupi_n_2050 ,csa_tree_add_7_25_groupi_n_2329);
  not csa_tree_add_7_25_groupi_drc_bufs20014(csa_tree_add_7_25_groupi_n_2049 ,csa_tree_add_7_25_groupi_n_2047);
  not csa_tree_add_7_25_groupi_drc_bufs20015(csa_tree_add_7_25_groupi_n_2048 ,csa_tree_add_7_25_groupi_n_2047);
  not csa_tree_add_7_25_groupi_drc_bufs20016(csa_tree_add_7_25_groupi_n_2047 ,csa_tree_add_7_25_groupi_n_2783);
  not csa_tree_add_7_25_groupi_drc_bufs20018(csa_tree_add_7_25_groupi_n_2046 ,csa_tree_add_7_25_groupi_n_2044);
  not csa_tree_add_7_25_groupi_drc_bufs20019(csa_tree_add_7_25_groupi_n_2045 ,csa_tree_add_7_25_groupi_n_2044);
  not csa_tree_add_7_25_groupi_drc_bufs20020(csa_tree_add_7_25_groupi_n_2044 ,csa_tree_add_7_25_groupi_n_2329);
  not csa_tree_add_7_25_groupi_drc_bufs20022(csa_tree_add_7_25_groupi_n_2043 ,csa_tree_add_7_25_groupi_n_2041);
  not csa_tree_add_7_25_groupi_drc_bufs20023(csa_tree_add_7_25_groupi_n_2042 ,csa_tree_add_7_25_groupi_n_2041);
  not csa_tree_add_7_25_groupi_drc_bufs20024(csa_tree_add_7_25_groupi_n_2041 ,csa_tree_add_7_25_groupi_n_2328);
  not csa_tree_add_7_25_groupi_drc_bufs20026(csa_tree_add_7_25_groupi_n_2040 ,csa_tree_add_7_25_groupi_n_2038);
  not csa_tree_add_7_25_groupi_drc_bufs20027(csa_tree_add_7_25_groupi_n_2039 ,csa_tree_add_7_25_groupi_n_2038);
  not csa_tree_add_7_25_groupi_drc_bufs20028(csa_tree_add_7_25_groupi_n_2038 ,csa_tree_add_7_25_groupi_n_2330);
  not csa_tree_add_7_25_groupi_drc_bufs20030(csa_tree_add_7_25_groupi_n_2037 ,csa_tree_add_7_25_groupi_n_2035);
  not csa_tree_add_7_25_groupi_drc_bufs20031(csa_tree_add_7_25_groupi_n_2036 ,csa_tree_add_7_25_groupi_n_2035);
  not csa_tree_add_7_25_groupi_drc_bufs20032(csa_tree_add_7_25_groupi_n_2035 ,csa_tree_add_7_25_groupi_n_2783);
  not csa_tree_add_7_25_groupi_drc_bufs20034(csa_tree_add_7_25_groupi_n_2034 ,csa_tree_add_7_25_groupi_n_2032);
  not csa_tree_add_7_25_groupi_drc_bufs20035(csa_tree_add_7_25_groupi_n_2033 ,csa_tree_add_7_25_groupi_n_2032);
  not csa_tree_add_7_25_groupi_drc_bufs20036(csa_tree_add_7_25_groupi_n_2032 ,csa_tree_add_7_25_groupi_n_2330);
  not csa_tree_add_7_25_groupi_drc_bufs20038(csa_tree_add_7_25_groupi_n_2031 ,csa_tree_add_7_25_groupi_n_2029);
  not csa_tree_add_7_25_groupi_drc_bufs20039(csa_tree_add_7_25_groupi_n_2030 ,csa_tree_add_7_25_groupi_n_2029);
  not csa_tree_add_7_25_groupi_drc_bufs20040(csa_tree_add_7_25_groupi_n_2029 ,csa_tree_add_7_25_groupi_n_2334);
  not csa_tree_add_7_25_groupi_drc_bufs20042(csa_tree_add_7_25_groupi_n_2028 ,csa_tree_add_7_25_groupi_n_2026);
  not csa_tree_add_7_25_groupi_drc_bufs20043(csa_tree_add_7_25_groupi_n_2027 ,csa_tree_add_7_25_groupi_n_2026);
  not csa_tree_add_7_25_groupi_drc_bufs20044(csa_tree_add_7_25_groupi_n_2026 ,csa_tree_add_7_25_groupi_n_2790);
  not csa_tree_add_7_25_groupi_drc_bufs20046(csa_tree_add_7_25_groupi_n_2025 ,csa_tree_add_7_25_groupi_n_2023);
  not csa_tree_add_7_25_groupi_drc_bufs20047(csa_tree_add_7_25_groupi_n_2024 ,csa_tree_add_7_25_groupi_n_2023);
  not csa_tree_add_7_25_groupi_drc_bufs20048(csa_tree_add_7_25_groupi_n_2023 ,csa_tree_add_7_25_groupi_n_2334);
  not csa_tree_add_7_25_groupi_drc_bufs20050(csa_tree_add_7_25_groupi_n_2022 ,csa_tree_add_7_25_groupi_n_2020);
  not csa_tree_add_7_25_groupi_drc_bufs20051(csa_tree_add_7_25_groupi_n_2021 ,csa_tree_add_7_25_groupi_n_2020);
  not csa_tree_add_7_25_groupi_drc_bufs20052(csa_tree_add_7_25_groupi_n_2020 ,csa_tree_add_7_25_groupi_n_2332);
  not csa_tree_add_7_25_groupi_drc_bufs20054(csa_tree_add_7_25_groupi_n_2019 ,csa_tree_add_7_25_groupi_n_2017);
  not csa_tree_add_7_25_groupi_drc_bufs20055(csa_tree_add_7_25_groupi_n_2018 ,csa_tree_add_7_25_groupi_n_2017);
  not csa_tree_add_7_25_groupi_drc_bufs20056(csa_tree_add_7_25_groupi_n_2017 ,csa_tree_add_7_25_groupi_n_2333);
  not csa_tree_add_7_25_groupi_drc_bufs20058(csa_tree_add_7_25_groupi_n_2016 ,csa_tree_add_7_25_groupi_n_2014);
  not csa_tree_add_7_25_groupi_drc_bufs20059(csa_tree_add_7_25_groupi_n_2015 ,csa_tree_add_7_25_groupi_n_2014);
  not csa_tree_add_7_25_groupi_drc_bufs20060(csa_tree_add_7_25_groupi_n_2014 ,csa_tree_add_7_25_groupi_n_2789);
  not csa_tree_add_7_25_groupi_drc_bufs20062(csa_tree_add_7_25_groupi_n_2013 ,csa_tree_add_7_25_groupi_n_2011);
  not csa_tree_add_7_25_groupi_drc_bufs20063(csa_tree_add_7_25_groupi_n_2012 ,csa_tree_add_7_25_groupi_n_2011);
  not csa_tree_add_7_25_groupi_drc_bufs20064(csa_tree_add_7_25_groupi_n_2011 ,csa_tree_add_7_25_groupi_n_2788);
  not csa_tree_add_7_25_groupi_drc_bufs20066(csa_tree_add_7_25_groupi_n_2010 ,csa_tree_add_7_25_groupi_n_2008);
  not csa_tree_add_7_25_groupi_drc_bufs20067(csa_tree_add_7_25_groupi_n_2009 ,csa_tree_add_7_25_groupi_n_2008);
  not csa_tree_add_7_25_groupi_drc_bufs20068(csa_tree_add_7_25_groupi_n_2008 ,csa_tree_add_7_25_groupi_n_2339);
  not csa_tree_add_7_25_groupi_drc_bufs20070(csa_tree_add_7_25_groupi_n_2007 ,csa_tree_add_7_25_groupi_n_2005);
  not csa_tree_add_7_25_groupi_drc_bufs20071(csa_tree_add_7_25_groupi_n_2006 ,csa_tree_add_7_25_groupi_n_2005);
  not csa_tree_add_7_25_groupi_drc_bufs20072(csa_tree_add_7_25_groupi_n_2005 ,csa_tree_add_7_25_groupi_n_3522);
  not csa_tree_add_7_25_groupi_drc_bufs20074(csa_tree_add_7_25_groupi_n_2004 ,csa_tree_add_7_25_groupi_n_2002);
  not csa_tree_add_7_25_groupi_drc_bufs20075(csa_tree_add_7_25_groupi_n_2003 ,csa_tree_add_7_25_groupi_n_2002);
  not csa_tree_add_7_25_groupi_drc_bufs20076(csa_tree_add_7_25_groupi_n_2002 ,csa_tree_add_7_25_groupi_n_2338);
  not csa_tree_add_7_25_groupi_drc_bufs20078(csa_tree_add_7_25_groupi_n_2001 ,csa_tree_add_7_25_groupi_n_1999);
  not csa_tree_add_7_25_groupi_drc_bufs20079(csa_tree_add_7_25_groupi_n_2000 ,csa_tree_add_7_25_groupi_n_1999);
  not csa_tree_add_7_25_groupi_drc_bufs20080(csa_tree_add_7_25_groupi_n_1999 ,csa_tree_add_7_25_groupi_n_2868);
  not csa_tree_add_7_25_groupi_drc_bufs20082(csa_tree_add_7_25_groupi_n_1998 ,csa_tree_add_7_25_groupi_n_1996);
  not csa_tree_add_7_25_groupi_drc_bufs20083(csa_tree_add_7_25_groupi_n_1997 ,csa_tree_add_7_25_groupi_n_1996);
  not csa_tree_add_7_25_groupi_drc_bufs20084(csa_tree_add_7_25_groupi_n_1996 ,csa_tree_add_7_25_groupi_n_2331);
  not csa_tree_add_7_25_groupi_drc_bufs20086(csa_tree_add_7_25_groupi_n_1995 ,csa_tree_add_7_25_groupi_n_1993);
  not csa_tree_add_7_25_groupi_drc_bufs20087(csa_tree_add_7_25_groupi_n_1994 ,csa_tree_add_7_25_groupi_n_1993);
  not csa_tree_add_7_25_groupi_drc_bufs20088(csa_tree_add_7_25_groupi_n_1993 ,csa_tree_add_7_25_groupi_n_2340);
  not csa_tree_add_7_25_groupi_drc_bufs20639(csa_tree_add_7_25_groupi_n_1992 ,csa_tree_add_7_25_groupi_n_1991);
  not csa_tree_add_7_25_groupi_drc_bufs20641(csa_tree_add_7_25_groupi_n_1991 ,csa_tree_add_7_25_groupi_n_2782);
  not csa_tree_add_7_25_groupi_drc_bufs20644(csa_tree_add_7_25_groupi_n_1990 ,csa_tree_add_7_25_groupi_n_2340);
  not csa_tree_add_7_25_groupi_drc_bufs20645(csa_tree_add_7_25_groupi_n_2340 ,csa_tree_add_7_25_groupi_n_3526);
  not csa_tree_add_7_25_groupi_drc_bufs20648(csa_tree_add_7_25_groupi_n_1989 ,csa_tree_add_7_25_groupi_n_1988);
  not csa_tree_add_7_25_groupi_drc_bufs20649(csa_tree_add_7_25_groupi_n_1988 ,csa_tree_add_7_25_groupi_n_2862);
  not csa_tree_add_7_25_groupi_drc_bufs20652(csa_tree_add_7_25_groupi_n_1987 ,csa_tree_add_7_25_groupi_n_1986);
  not csa_tree_add_7_25_groupi_drc_bufs20653(csa_tree_add_7_25_groupi_n_1986 ,csa_tree_add_7_25_groupi_n_3516);
  not csa_tree_add_7_25_groupi_drc_bufs20656(csa_tree_add_7_25_groupi_n_1985 ,csa_tree_add_7_25_groupi_n_1984);
  not csa_tree_add_7_25_groupi_drc_bufs20657(csa_tree_add_7_25_groupi_n_1984 ,csa_tree_add_7_25_groupi_n_2857);
  not csa_tree_add_7_25_groupi_drc_bufs20660(csa_tree_add_7_25_groupi_n_1983 ,csa_tree_add_7_25_groupi_n_1982);
  not csa_tree_add_7_25_groupi_drc_bufs20661(csa_tree_add_7_25_groupi_n_1982 ,csa_tree_add_7_25_groupi_n_2852);
  not csa_tree_add_7_25_groupi_drc_bufs20664(csa_tree_add_7_25_groupi_n_1981 ,csa_tree_add_7_25_groupi_n_1980);
  not csa_tree_add_7_25_groupi_drc_bufs20665(csa_tree_add_7_25_groupi_n_1980 ,csa_tree_add_7_25_groupi_n_3511);
  not csa_tree_add_7_25_groupi_drc_bufs20668(csa_tree_add_7_25_groupi_n_1979 ,csa_tree_add_7_25_groupi_n_1978);
  not csa_tree_add_7_25_groupi_drc_bufs20669(csa_tree_add_7_25_groupi_n_1978 ,csa_tree_add_7_25_groupi_n_2847);
  not csa_tree_add_7_25_groupi_drc_bufs20672(csa_tree_add_7_25_groupi_n_1977 ,csa_tree_add_7_25_groupi_n_1976);
  not csa_tree_add_7_25_groupi_drc_bufs20673(csa_tree_add_7_25_groupi_n_1976 ,csa_tree_add_7_25_groupi_n_3506);
  not csa_tree_add_7_25_groupi_drc_bufs20676(csa_tree_add_7_25_groupi_n_1975 ,csa_tree_add_7_25_groupi_n_1974);
  not csa_tree_add_7_25_groupi_drc_bufs20677(csa_tree_add_7_25_groupi_n_1974 ,csa_tree_add_7_25_groupi_n_3501);
  not csa_tree_add_7_25_groupi_drc_bufs20680(csa_tree_add_7_25_groupi_n_1973 ,csa_tree_add_7_25_groupi_n_2346);
  not csa_tree_add_7_25_groupi_drc_bufs20681(csa_tree_add_7_25_groupi_n_2346 ,csa_tree_add_7_25_groupi_n_5386);
  not csa_tree_add_7_25_groupi_drc_bufs20684(csa_tree_add_7_25_groupi_n_1972 ,csa_tree_add_7_25_groupi_n_2341);
  not csa_tree_add_7_25_groupi_drc_bufs20685(csa_tree_add_7_25_groupi_n_2341 ,csa_tree_add_7_25_groupi_n_4369);
  not csa_tree_add_7_25_groupi_drc_bufs20691(csa_tree_add_7_25_groupi_n_1971 ,csa_tree_add_7_25_groupi_n_1970);
  not csa_tree_add_7_25_groupi_drc_bufs20692(csa_tree_add_7_25_groupi_n_1970 ,csa_tree_add_7_25_groupi_n_2684);
  not csa_tree_add_7_25_groupi_drc_bufs20695(csa_tree_add_7_25_groupi_n_1969 ,csa_tree_add_7_25_groupi_n_1968);
  not csa_tree_add_7_25_groupi_drc_bufs20696(csa_tree_add_7_25_groupi_n_1968 ,csa_tree_add_7_25_groupi_n_2520);
  not csa_tree_add_7_25_groupi_drc_bufs20699(csa_tree_add_7_25_groupi_n_1967 ,csa_tree_add_7_25_groupi_n_1966);
  not csa_tree_add_7_25_groupi_drc_bufs20700(csa_tree_add_7_25_groupi_n_1966 ,csa_tree_add_7_25_groupi_n_2842);
  not csa_tree_add_7_25_groupi_drc_bufs20703(csa_tree_add_7_25_groupi_n_1965 ,csa_tree_add_7_25_groupi_n_1964);
  not csa_tree_add_7_25_groupi_drc_bufs20704(csa_tree_add_7_25_groupi_n_1964 ,csa_tree_add_7_25_groupi_n_2776);
  not csa_tree_add_7_25_groupi_drc_bufs20707(csa_tree_add_7_25_groupi_n_1963 ,csa_tree_add_7_25_groupi_n_1962);
  not csa_tree_add_7_25_groupi_drc_bufs20708(csa_tree_add_7_25_groupi_n_1962 ,csa_tree_add_7_25_groupi_n_2771);
  not csa_tree_add_7_25_groupi_drc_bufs20711(csa_tree_add_7_25_groupi_n_1961 ,csa_tree_add_7_25_groupi_n_1960);
  not csa_tree_add_7_25_groupi_drc_bufs20712(csa_tree_add_7_25_groupi_n_1960 ,csa_tree_add_7_25_groupi_n_2766);
  not csa_tree_add_7_25_groupi_drc_bufs20715(csa_tree_add_7_25_groupi_n_1959 ,csa_tree_add_7_25_groupi_n_1958);
  not csa_tree_add_7_25_groupi_drc_bufs20716(csa_tree_add_7_25_groupi_n_1958 ,csa_tree_add_7_25_groupi_n_2761);
  not csa_tree_add_7_25_groupi_drc_bufs20719(csa_tree_add_7_25_groupi_n_1957 ,csa_tree_add_7_25_groupi_n_1956);
  not csa_tree_add_7_25_groupi_drc_bufs20720(csa_tree_add_7_25_groupi_n_1956 ,csa_tree_add_7_25_groupi_n_2756);
  not csa_tree_add_7_25_groupi_drc_bufs21184(csa_tree_add_7_25_groupi_n_1955 ,csa_tree_add_7_25_groupi_n_1953);
  not csa_tree_add_7_25_groupi_drc_bufs21185(csa_tree_add_7_25_groupi_n_1954 ,csa_tree_add_7_25_groupi_n_1953);
  not csa_tree_add_7_25_groupi_drc_bufs21186(csa_tree_add_7_25_groupi_n_1953 ,csa_tree_add_7_25_groupi_n_2366);
  not csa_tree_add_7_25_groupi_drc_bufs21204(csa_tree_add_7_25_groupi_n_1952 ,csa_tree_add_7_25_groupi_n_1950);
  not csa_tree_add_7_25_groupi_drc_bufs21205(csa_tree_add_7_25_groupi_n_1951 ,csa_tree_add_7_25_groupi_n_1950);
  not csa_tree_add_7_25_groupi_drc_bufs21206(csa_tree_add_7_25_groupi_n_1950 ,csa_tree_add_7_25_groupi_n_2367);
  not csa_tree_add_7_25_groupi_drc_bufs21219(csa_tree_add_7_25_groupi_n_1949 ,csa_tree_add_7_25_groupi_n_1947);
  not csa_tree_add_7_25_groupi_drc_bufs21220(csa_tree_add_7_25_groupi_n_1948 ,csa_tree_add_7_25_groupi_n_1947);
  not csa_tree_add_7_25_groupi_drc_bufs21221(csa_tree_add_7_25_groupi_n_1947 ,csa_tree_add_7_25_groupi_n_2887);
  not csa_tree_add_7_25_groupi_drc_bufs21379(csa_tree_add_7_25_groupi_n_1946 ,csa_tree_add_7_25_groupi_n_1945);
  not csa_tree_add_7_25_groupi_drc_bufs21381(csa_tree_add_7_25_groupi_n_1945 ,csa_tree_add_7_25_groupi_n_2403);
  not csa_tree_add_7_25_groupi_drc_bufs21389(csa_tree_add_7_25_groupi_n_1944 ,csa_tree_add_7_25_groupi_n_1943);
  not csa_tree_add_7_25_groupi_drc_bufs21391(csa_tree_add_7_25_groupi_n_1943 ,csa_tree_add_7_25_groupi_n_2888);
  not csa_tree_add_7_25_groupi_drc_bufs21394(csa_tree_add_7_25_groupi_n_1942 ,csa_tree_add_7_25_groupi_n_1941);
  not csa_tree_add_7_25_groupi_drc_bufs21396(csa_tree_add_7_25_groupi_n_1941 ,csa_tree_add_7_25_groupi_n_3535);
  not csa_tree_add_7_25_groupi_drc_bufs21409(csa_tree_add_7_25_groupi_n_1940 ,csa_tree_add_7_25_groupi_n_1939);
  not csa_tree_add_7_25_groupi_drc_bufs21411(csa_tree_add_7_25_groupi_n_1939 ,csa_tree_add_7_25_groupi_n_2889);
  not csa_tree_add_7_25_groupi_drc_bufs21478(csa_tree_add_7_25_groupi_n_1938 ,csa_tree_add_7_25_groupi_n_1936);
  not csa_tree_add_7_25_groupi_drc_bufs21479(csa_tree_add_7_25_groupi_n_1937 ,csa_tree_add_7_25_groupi_n_1936);
  not csa_tree_add_7_25_groupi_drc_bufs21480(csa_tree_add_7_25_groupi_n_1936 ,csa_tree_add_7_25_groupi_n_2801);
  not csa_tree_add_7_25_groupi_drc_bufs21482(csa_tree_add_7_25_groupi_n_1935 ,csa_tree_add_7_25_groupi_n_1933);
  not csa_tree_add_7_25_groupi_drc_bufs21483(csa_tree_add_7_25_groupi_n_1934 ,csa_tree_add_7_25_groupi_n_1933);
  not csa_tree_add_7_25_groupi_drc_bufs21484(csa_tree_add_7_25_groupi_n_1933 ,csa_tree_add_7_25_groupi_n_2801);
  not csa_tree_add_7_25_groupi_drc_bufs21486(csa_tree_add_7_25_groupi_n_1932 ,csa_tree_add_7_25_groupi_n_1930);
  not csa_tree_add_7_25_groupi_drc_bufs21487(csa_tree_add_7_25_groupi_n_1931 ,csa_tree_add_7_25_groupi_n_1930);
  not csa_tree_add_7_25_groupi_drc_bufs21488(csa_tree_add_7_25_groupi_n_1930 ,csa_tree_add_7_25_groupi_n_2798);
  not csa_tree_add_7_25_groupi_drc_bufs21490(csa_tree_add_7_25_groupi_n_1929 ,csa_tree_add_7_25_groupi_n_1927);
  not csa_tree_add_7_25_groupi_drc_bufs21491(csa_tree_add_7_25_groupi_n_1928 ,csa_tree_add_7_25_groupi_n_1927);
  not csa_tree_add_7_25_groupi_drc_bufs21492(csa_tree_add_7_25_groupi_n_1927 ,csa_tree_add_7_25_groupi_n_2879);
  not csa_tree_add_7_25_groupi_drc_bufs21494(csa_tree_add_7_25_groupi_n_1926 ,csa_tree_add_7_25_groupi_n_1924);
  not csa_tree_add_7_25_groupi_drc_bufs21495(csa_tree_add_7_25_groupi_n_1925 ,csa_tree_add_7_25_groupi_n_1924);
  not csa_tree_add_7_25_groupi_drc_bufs21496(csa_tree_add_7_25_groupi_n_1924 ,csa_tree_add_7_25_groupi_n_2803);
  not csa_tree_add_7_25_groupi_drc_bufs21498(csa_tree_add_7_25_groupi_n_1923 ,csa_tree_add_7_25_groupi_n_1921);
  not csa_tree_add_7_25_groupi_drc_bufs21499(csa_tree_add_7_25_groupi_n_1922 ,csa_tree_add_7_25_groupi_n_1921);
  not csa_tree_add_7_25_groupi_drc_bufs21500(csa_tree_add_7_25_groupi_n_1921 ,csa_tree_add_7_25_groupi_n_2798);
  not csa_tree_add_7_25_groupi_drc_bufs21506(csa_tree_add_7_25_groupi_n_1920 ,csa_tree_add_7_25_groupi_n_1918);
  not csa_tree_add_7_25_groupi_drc_bufs21507(csa_tree_add_7_25_groupi_n_1919 ,csa_tree_add_7_25_groupi_n_1918);
  not csa_tree_add_7_25_groupi_drc_bufs21508(csa_tree_add_7_25_groupi_n_1918 ,csa_tree_add_7_25_groupi_n_2687);
  not csa_tree_add_7_25_groupi_drc_bufs21618(csa_tree_add_7_25_groupi_n_1917 ,csa_tree_add_7_25_groupi_n_1915);
  not csa_tree_add_7_25_groupi_drc_bufs21619(csa_tree_add_7_25_groupi_n_1916 ,csa_tree_add_7_25_groupi_n_1915);
  not csa_tree_add_7_25_groupi_drc_bufs21620(csa_tree_add_7_25_groupi_n_1915 ,csa_tree_add_7_25_groupi_n_2885);
  not csa_tree_add_7_25_groupi_drc_bufs21638(csa_tree_add_7_25_groupi_n_1914 ,csa_tree_add_7_25_groupi_n_1912);
  not csa_tree_add_7_25_groupi_drc_bufs21639(csa_tree_add_7_25_groupi_n_1913 ,csa_tree_add_7_25_groupi_n_1912);
  not csa_tree_add_7_25_groupi_drc_bufs21640(csa_tree_add_7_25_groupi_n_1912 ,csa_tree_add_7_25_groupi_n_2873);
  not csa_tree_add_7_25_groupi_drc_bufs21642(csa_tree_add_7_25_groupi_n_1911 ,csa_tree_add_7_25_groupi_n_1909);
  not csa_tree_add_7_25_groupi_drc_bufs21643(csa_tree_add_7_25_groupi_n_1910 ,csa_tree_add_7_25_groupi_n_1909);
  not csa_tree_add_7_25_groupi_drc_bufs21644(csa_tree_add_7_25_groupi_n_1909 ,csa_tree_add_7_25_groupi_n_2879);
  not csa_tree_add_7_25_groupi_drc_bufs21646(csa_tree_add_7_25_groupi_n_1908 ,csa_tree_add_7_25_groupi_n_1906);
  not csa_tree_add_7_25_groupi_drc_bufs21647(csa_tree_add_7_25_groupi_n_1907 ,csa_tree_add_7_25_groupi_n_1906);
  not csa_tree_add_7_25_groupi_drc_bufs21648(csa_tree_add_7_25_groupi_n_1906 ,csa_tree_add_7_25_groupi_n_3533);
  not csa_tree_add_7_25_groupi_drc_bufs21650(csa_tree_add_7_25_groupi_n_1905 ,csa_tree_add_7_25_groupi_n_1903);
  not csa_tree_add_7_25_groupi_drc_bufs21651(csa_tree_add_7_25_groupi_n_1904 ,csa_tree_add_7_25_groupi_n_1903);
  not csa_tree_add_7_25_groupi_drc_bufs21652(csa_tree_add_7_25_groupi_n_1903 ,csa_tree_add_7_25_groupi_n_3533);
  not csa_tree_add_7_25_groupi_drc_bufs21654(csa_tree_add_7_25_groupi_n_1902 ,csa_tree_add_7_25_groupi_n_1900);
  not csa_tree_add_7_25_groupi_drc_bufs21655(csa_tree_add_7_25_groupi_n_1901 ,csa_tree_add_7_25_groupi_n_1900);
  not csa_tree_add_7_25_groupi_drc_bufs21656(csa_tree_add_7_25_groupi_n_1900 ,csa_tree_add_7_25_groupi_n_2882);
  not csa_tree_add_7_25_groupi_drc_bufs21659(csa_tree_add_7_25_groupi_n_1899 ,csa_tree_add_7_25_groupi_n_1898);
  not csa_tree_add_7_25_groupi_drc_bufs21660(csa_tree_add_7_25_groupi_n_1898 ,csa_tree_add_7_25_groupi_n_2207);
  not csa_tree_add_7_25_groupi_drc_bufs21663(csa_tree_add_7_25_groupi_n_1897 ,csa_tree_add_7_25_groupi_n_1896);
  not csa_tree_add_7_25_groupi_drc_bufs21664(csa_tree_add_7_25_groupi_n_1896 ,csa_tree_add_7_25_groupi_n_2206);
  not csa_tree_add_7_25_groupi_drc_bufs21667(csa_tree_add_7_25_groupi_n_1895 ,csa_tree_add_7_25_groupi_n_1894);
  not csa_tree_add_7_25_groupi_drc_bufs21668(csa_tree_add_7_25_groupi_n_1894 ,csa_tree_add_7_25_groupi_n_2205);
  not csa_tree_add_7_25_groupi_drc_bufs21671(csa_tree_add_7_25_groupi_n_1893 ,csa_tree_add_7_25_groupi_n_1892);
  not csa_tree_add_7_25_groupi_drc_bufs21672(csa_tree_add_7_25_groupi_n_1892 ,csa_tree_add_7_25_groupi_n_2204);
  not csa_tree_add_7_25_groupi_drc_bufs21675(csa_tree_add_7_25_groupi_n_1891 ,csa_tree_add_7_25_groupi_n_1890);
  not csa_tree_add_7_25_groupi_drc_bufs21676(csa_tree_add_7_25_groupi_n_1890 ,csa_tree_add_7_25_groupi_n_2203);
  not csa_tree_add_7_25_groupi_drc_bufs21679(csa_tree_add_7_25_groupi_n_1889 ,csa_tree_add_7_25_groupi_n_1888);
  not csa_tree_add_7_25_groupi_drc_bufs21680(csa_tree_add_7_25_groupi_n_1888 ,csa_tree_add_7_25_groupi_n_2201);
  not csa_tree_add_7_25_groupi_drc_bufs21683(csa_tree_add_7_25_groupi_n_1887 ,csa_tree_add_7_25_groupi_n_1886);
  not csa_tree_add_7_25_groupi_drc_bufs21684(csa_tree_add_7_25_groupi_n_1886 ,csa_tree_add_7_25_groupi_n_2200);
  not csa_tree_add_7_25_groupi_drc_bufs21687(csa_tree_add_7_25_groupi_n_1885 ,csa_tree_add_7_25_groupi_n_1884);
  not csa_tree_add_7_25_groupi_drc_bufs21688(csa_tree_add_7_25_groupi_n_1884 ,csa_tree_add_7_25_groupi_n_2210);
  not csa_tree_add_7_25_groupi_drc_bufs21691(csa_tree_add_7_25_groupi_n_1883 ,csa_tree_add_7_25_groupi_n_1882);
  not csa_tree_add_7_25_groupi_drc_bufs21692(csa_tree_add_7_25_groupi_n_1882 ,csa_tree_add_7_25_groupi_n_2199);
  not csa_tree_add_7_25_groupi_drc_bufs21695(csa_tree_add_7_25_groupi_n_1881 ,csa_tree_add_7_25_groupi_n_1880);
  not csa_tree_add_7_25_groupi_drc_bufs21696(csa_tree_add_7_25_groupi_n_1880 ,csa_tree_add_7_25_groupi_n_2198);
  not csa_tree_add_7_25_groupi_drc_bufs21698(csa_tree_add_7_25_groupi_n_1879 ,csa_tree_add_7_25_groupi_n_1877);
  not csa_tree_add_7_25_groupi_drc_bufs21699(csa_tree_add_7_25_groupi_n_1878 ,csa_tree_add_7_25_groupi_n_1877);
  not csa_tree_add_7_25_groupi_drc_bufs21700(csa_tree_add_7_25_groupi_n_1877 ,csa_tree_add_7_25_groupi_n_2885);
  not csa_tree_add_7_25_groupi_drc_bufs21702(csa_tree_add_7_25_groupi_n_1876 ,csa_tree_add_7_25_groupi_n_1874);
  not csa_tree_add_7_25_groupi_drc_bufs21703(csa_tree_add_7_25_groupi_n_1875 ,csa_tree_add_7_25_groupi_n_1874);
  not csa_tree_add_7_25_groupi_drc_bufs21704(csa_tree_add_7_25_groupi_n_1874 ,csa_tree_add_7_25_groupi_n_2614);
  not csa_tree_add_7_25_groupi_drc_bufs21706(csa_tree_add_7_25_groupi_n_1873 ,csa_tree_add_7_25_groupi_n_1871);
  not csa_tree_add_7_25_groupi_drc_bufs21707(csa_tree_add_7_25_groupi_n_1872 ,csa_tree_add_7_25_groupi_n_1871);
  not csa_tree_add_7_25_groupi_drc_bufs21708(csa_tree_add_7_25_groupi_n_1871 ,csa_tree_add_7_25_groupi_n_4198);
  not csa_tree_add_7_25_groupi_drc_bufs21711(csa_tree_add_7_25_groupi_n_1870 ,csa_tree_add_7_25_groupi_n_1869);
  not csa_tree_add_7_25_groupi_drc_bufs21712(csa_tree_add_7_25_groupi_n_1869 ,csa_tree_add_7_25_groupi_n_5533);
  not csa_tree_add_7_25_groupi_drc_bufs21714(csa_tree_add_7_25_groupi_n_1868 ,csa_tree_add_7_25_groupi_n_1866);
  not csa_tree_add_7_25_groupi_drc_bufs21715(csa_tree_add_7_25_groupi_n_1867 ,csa_tree_add_7_25_groupi_n_1866);
  not csa_tree_add_7_25_groupi_drc_bufs21716(csa_tree_add_7_25_groupi_n_1866 ,csa_tree_add_7_25_groupi_n_3742);
  not csa_tree_add_7_25_groupi_drc_bufs21718(csa_tree_add_7_25_groupi_n_1865 ,csa_tree_add_7_25_groupi_n_1863);
  not csa_tree_add_7_25_groupi_drc_bufs21719(csa_tree_add_7_25_groupi_n_1864 ,csa_tree_add_7_25_groupi_n_1863);
  not csa_tree_add_7_25_groupi_drc_bufs21720(csa_tree_add_7_25_groupi_n_1863 ,csa_tree_add_7_25_groupi_n_3199);
  not csa_tree_add_7_25_groupi_drc_bufs21722(csa_tree_add_7_25_groupi_n_1862 ,csa_tree_add_7_25_groupi_n_1860);
  not csa_tree_add_7_25_groupi_drc_bufs21723(csa_tree_add_7_25_groupi_n_1861 ,csa_tree_add_7_25_groupi_n_1860);
  not csa_tree_add_7_25_groupi_drc_bufs21724(csa_tree_add_7_25_groupi_n_1860 ,csa_tree_add_7_25_groupi_n_4792);
  not csa_tree_add_7_25_groupi_drc_bufs21726(csa_tree_add_7_25_groupi_n_1859 ,csa_tree_add_7_25_groupi_n_1857);
  not csa_tree_add_7_25_groupi_drc_bufs21727(csa_tree_add_7_25_groupi_n_1858 ,csa_tree_add_7_25_groupi_n_1857);
  not csa_tree_add_7_25_groupi_drc_bufs21728(csa_tree_add_7_25_groupi_n_1857 ,csa_tree_add_7_25_groupi_n_4676);
  not csa_tree_add_7_25_groupi_drc_bufs21731(csa_tree_add_7_25_groupi_n_1856 ,csa_tree_add_7_25_groupi_n_1855);
  not csa_tree_add_7_25_groupi_drc_bufs21732(csa_tree_add_7_25_groupi_n_1855 ,csa_tree_add_7_25_groupi_n_5423);
  not csa_tree_add_7_25_groupi_drc_bufs21734(csa_tree_add_7_25_groupi_n_1854 ,csa_tree_add_7_25_groupi_n_1853);
  not csa_tree_add_7_25_groupi_drc_bufs21736(csa_tree_add_7_25_groupi_n_1853 ,csa_tree_add_7_25_groupi_n_5648);
  not csa_tree_add_7_25_groupi_drc_bufs21738(csa_tree_add_7_25_groupi_n_1852 ,csa_tree_add_7_25_groupi_n_1850);
  not csa_tree_add_7_25_groupi_drc_bufs21739(csa_tree_add_7_25_groupi_n_1851 ,csa_tree_add_7_25_groupi_n_1850);
  not csa_tree_add_7_25_groupi_drc_bufs21740(csa_tree_add_7_25_groupi_n_1850 ,csa_tree_add_7_25_groupi_n_2873);
  not csa_tree_add_7_25_groupi_drc_bufs21742(csa_tree_add_7_25_groupi_n_1849 ,csa_tree_add_7_25_groupi_n_1847);
  not csa_tree_add_7_25_groupi_drc_bufs21743(csa_tree_add_7_25_groupi_n_1848 ,csa_tree_add_7_25_groupi_n_1847);
  not csa_tree_add_7_25_groupi_drc_bufs21744(csa_tree_add_7_25_groupi_n_1847 ,csa_tree_add_7_25_groupi_n_2882);
  not csa_tree_add_7_25_groupi_drc_bufs21746(csa_tree_add_7_25_groupi_n_1846 ,csa_tree_add_7_25_groupi_n_1844);
  not csa_tree_add_7_25_groupi_drc_bufs21747(csa_tree_add_7_25_groupi_n_1845 ,csa_tree_add_7_25_groupi_n_1844);
  not csa_tree_add_7_25_groupi_drc_bufs21748(csa_tree_add_7_25_groupi_n_1844 ,csa_tree_add_7_25_groupi_n_5188);
  not csa_tree_add_7_25_groupi_drc_bufs21750(csa_tree_add_7_25_groupi_n_1843 ,csa_tree_add_7_25_groupi_n_1841);
  not csa_tree_add_7_25_groupi_drc_bufs21751(csa_tree_add_7_25_groupi_n_1842 ,csa_tree_add_7_25_groupi_n_1841);
  not csa_tree_add_7_25_groupi_drc_bufs21752(csa_tree_add_7_25_groupi_n_1841 ,csa_tree_add_7_25_groupi_n_4460);
  not csa_tree_add_7_25_groupi_drc_bufs21754(csa_tree_add_7_25_groupi_n_1840 ,csa_tree_add_7_25_groupi_n_1838);
  not csa_tree_add_7_25_groupi_drc_bufs21755(csa_tree_add_7_25_groupi_n_1839 ,csa_tree_add_7_25_groupi_n_1838);
  not csa_tree_add_7_25_groupi_drc_bufs21756(csa_tree_add_7_25_groupi_n_1838 ,csa_tree_add_7_25_groupi_n_4351);
  not csa_tree_add_7_25_groupi_drc_bufs21758(csa_tree_add_7_25_groupi_n_1837 ,csa_tree_add_7_25_groupi_n_1835);
  not csa_tree_add_7_25_groupi_drc_bufs21759(csa_tree_add_7_25_groupi_n_1836 ,csa_tree_add_7_25_groupi_n_1835);
  not csa_tree_add_7_25_groupi_drc_bufs21760(csa_tree_add_7_25_groupi_n_1835 ,csa_tree_add_7_25_groupi_n_5303);
  not csa_tree_add_7_25_groupi_drc_bufs21762(csa_tree_add_7_25_groupi_n_1834 ,csa_tree_add_7_25_groupi_n_1832);
  not csa_tree_add_7_25_groupi_drc_bufs21763(csa_tree_add_7_25_groupi_n_1833 ,csa_tree_add_7_25_groupi_n_1832);
  not csa_tree_add_7_25_groupi_drc_bufs21764(csa_tree_add_7_25_groupi_n_1832 ,csa_tree_add_7_25_groupi_n_4110);
  not csa_tree_add_7_25_groupi_drc_bufs21766(csa_tree_add_7_25_groupi_n_1831 ,csa_tree_add_7_25_groupi_n_1829);
  not csa_tree_add_7_25_groupi_drc_bufs21767(csa_tree_add_7_25_groupi_n_1830 ,csa_tree_add_7_25_groupi_n_1829);
  not csa_tree_add_7_25_groupi_drc_bufs21768(csa_tree_add_7_25_groupi_n_1829 ,csa_tree_add_7_25_groupi_n_5093);
  not csa_tree_add_7_25_groupi_drc_bufs21770(csa_tree_add_7_25_groupi_n_1828 ,csa_tree_add_7_25_groupi_n_1826);
  not csa_tree_add_7_25_groupi_drc_bufs21771(csa_tree_add_7_25_groupi_n_1827 ,csa_tree_add_7_25_groupi_n_1826);
  not csa_tree_add_7_25_groupi_drc_bufs21772(csa_tree_add_7_25_groupi_n_1826 ,csa_tree_add_7_25_groupi_n_5007);
  not csa_tree_add_7_25_groupi_drc_bufs21774(csa_tree_add_7_25_groupi_n_1825 ,csa_tree_add_7_25_groupi_n_1823);
  not csa_tree_add_7_25_groupi_drc_bufs21775(csa_tree_add_7_25_groupi_n_1824 ,csa_tree_add_7_25_groupi_n_1823);
  not csa_tree_add_7_25_groupi_drc_bufs21776(csa_tree_add_7_25_groupi_n_1823 ,csa_tree_add_7_25_groupi_n_4903);
  not csa_tree_add_7_25_groupi_drc_bufs21778(csa_tree_add_7_25_groupi_n_1822 ,csa_tree_add_7_25_groupi_n_1820);
  not csa_tree_add_7_25_groupi_drc_bufs21779(csa_tree_add_7_25_groupi_n_1821 ,csa_tree_add_7_25_groupi_n_1820);
  not csa_tree_add_7_25_groupi_drc_bufs21780(csa_tree_add_7_25_groupi_n_1820 ,csa_tree_add_7_25_groupi_n_4573);
  not csa_tree_add_7_25_groupi_drc_bufs21782(csa_tree_add_7_25_groupi_n_1819 ,csa_tree_add_7_25_groupi_n_1817);
  not csa_tree_add_7_25_groupi_drc_bufs21783(csa_tree_add_7_25_groupi_n_1818 ,csa_tree_add_7_25_groupi_n_1817);
  not csa_tree_add_7_25_groupi_drc_bufs21784(csa_tree_add_7_25_groupi_n_1817 ,csa_tree_add_7_25_groupi_n_5423);
  not csa_tree_add_7_25_groupi_drc_bufs21786(csa_tree_add_7_25_groupi_n_1816 ,csa_tree_add_7_25_groupi_n_1814);
  not csa_tree_add_7_25_groupi_drc_bufs21787(csa_tree_add_7_25_groupi_n_1815 ,csa_tree_add_7_25_groupi_n_1814);
  not csa_tree_add_7_25_groupi_drc_bufs21788(csa_tree_add_7_25_groupi_n_1814 ,csa_tree_add_7_25_groupi_n_5648);
  not csa_tree_add_7_25_groupi_drc_bufs21790(csa_tree_add_7_25_groupi_n_1813 ,csa_tree_add_7_25_groupi_n_1811);
  not csa_tree_add_7_25_groupi_drc_bufs21791(csa_tree_add_7_25_groupi_n_1812 ,csa_tree_add_7_25_groupi_n_1811);
  not csa_tree_add_7_25_groupi_drc_bufs21792(csa_tree_add_7_25_groupi_n_1811 ,csa_tree_add_7_25_groupi_n_5533);
  not csa_tree_add_7_25_groupi_drc_bufs21795(csa_tree_add_7_25_groupi_n_1810 ,csa_tree_add_7_25_groupi_n_1809);
  not csa_tree_add_7_25_groupi_drc_bufs21796(csa_tree_add_7_25_groupi_n_1809 ,csa_tree_add_7_25_groupi_n_5979);
  not csa_tree_add_7_25_groupi_drc_bufs21799(csa_tree_add_7_25_groupi_n_1808 ,csa_tree_add_7_25_groupi_n_1807);
  not csa_tree_add_7_25_groupi_drc_bufs21800(csa_tree_add_7_25_groupi_n_1807 ,csa_tree_add_7_25_groupi_n_5864);
  not csa_tree_add_7_25_groupi_drc_bufs21803(csa_tree_add_7_25_groupi_n_1806 ,csa_tree_add_7_25_groupi_n_1805);
  not csa_tree_add_7_25_groupi_drc_bufs21804(csa_tree_add_7_25_groupi_n_1805 ,csa_tree_add_7_25_groupi_n_5763);
  not csa_tree_add_7_25_groupi_drc_bufs21808(csa_tree_add_7_25_groupi_n_1804 ,csa_tree_add_7_25_groupi_n_2837);
  not csa_tree_add_7_25_groupi_drc_bufs21812(csa_tree_add_7_25_groupi_n_1803 ,csa_tree_add_7_25_groupi_n_2747);
  not csa_tree_add_7_25_groupi_drc_bufs21816(csa_tree_add_7_25_groupi_n_1802 ,csa_tree_add_7_25_groupi_n_2743);
  not csa_tree_add_7_25_groupi_drc_bufs21820(csa_tree_add_7_25_groupi_n_1801 ,csa_tree_add_7_25_groupi_n_2739);
  not csa_tree_add_7_25_groupi_drc_bufs21824(csa_tree_add_7_25_groupi_n_1800 ,csa_tree_add_7_25_groupi_n_2751);
  not csa_tree_add_7_25_groupi_drc_bufs21826(csa_tree_add_7_25_groupi_n_1799 ,csa_tree_add_7_25_groupi_n_1797);
  not csa_tree_add_7_25_groupi_drc_bufs21827(csa_tree_add_7_25_groupi_n_1798 ,csa_tree_add_7_25_groupi_n_1797);
  not csa_tree_add_7_25_groupi_drc_bufs21828(csa_tree_add_7_25_groupi_n_1797 ,csa_tree_add_7_25_groupi_n_2796);
  not csa_tree_add_7_25_groupi_drc_bufs21830(csa_tree_add_7_25_groupi_n_1796 ,csa_tree_add_7_25_groupi_n_1794);
  not csa_tree_add_7_25_groupi_drc_bufs21831(csa_tree_add_7_25_groupi_n_1795 ,csa_tree_add_7_25_groupi_n_1794);
  not csa_tree_add_7_25_groupi_drc_bufs21832(csa_tree_add_7_25_groupi_n_1794 ,csa_tree_add_7_25_groupi_n_2802);
  not csa_tree_add_7_25_groupi_drc_bufs21834(csa_tree_add_7_25_groupi_n_1793 ,csa_tree_add_7_25_groupi_n_1791);
  not csa_tree_add_7_25_groupi_drc_bufs21835(csa_tree_add_7_25_groupi_n_1792 ,csa_tree_add_7_25_groupi_n_1791);
  not csa_tree_add_7_25_groupi_drc_bufs21836(csa_tree_add_7_25_groupi_n_1791 ,csa_tree_add_7_25_groupi_n_2786);
  not csa_tree_add_7_25_groupi_drc_bufs21838(csa_tree_add_7_25_groupi_n_1790 ,csa_tree_add_7_25_groupi_n_1788);
  not csa_tree_add_7_25_groupi_drc_bufs21839(csa_tree_add_7_25_groupi_n_1789 ,csa_tree_add_7_25_groupi_n_1788);
  not csa_tree_add_7_25_groupi_drc_bufs21840(csa_tree_add_7_25_groupi_n_1788 ,csa_tree_add_7_25_groupi_n_2786);
  not csa_tree_add_7_25_groupi_drc_bufs21842(csa_tree_add_7_25_groupi_n_1787 ,csa_tree_add_7_25_groupi_n_1785);
  not csa_tree_add_7_25_groupi_drc_bufs21843(csa_tree_add_7_25_groupi_n_1786 ,csa_tree_add_7_25_groupi_n_1785);
  not csa_tree_add_7_25_groupi_drc_bufs21844(csa_tree_add_7_25_groupi_n_1785 ,csa_tree_add_7_25_groupi_n_3520);
  not csa_tree_add_7_25_groupi_drc_bufs21846(csa_tree_add_7_25_groupi_n_1784 ,csa_tree_add_7_25_groupi_n_1782);
  not csa_tree_add_7_25_groupi_drc_bufs21847(csa_tree_add_7_25_groupi_n_1783 ,csa_tree_add_7_25_groupi_n_1782);
  not csa_tree_add_7_25_groupi_drc_bufs21848(csa_tree_add_7_25_groupi_n_1782 ,csa_tree_add_7_25_groupi_n_3520);
  not csa_tree_add_7_25_groupi_drc_bufs21850(csa_tree_add_7_25_groupi_n_1781 ,csa_tree_add_7_25_groupi_n_1779);
  not csa_tree_add_7_25_groupi_drc_bufs21851(csa_tree_add_7_25_groupi_n_1780 ,csa_tree_add_7_25_groupi_n_1779);
  not csa_tree_add_7_25_groupi_drc_bufs21852(csa_tree_add_7_25_groupi_n_1779 ,csa_tree_add_7_25_groupi_n_2866);
  not csa_tree_add_7_25_groupi_drc_bufs21854(csa_tree_add_7_25_groupi_n_1778 ,csa_tree_add_7_25_groupi_n_1776);
  not csa_tree_add_7_25_groupi_drc_bufs21855(csa_tree_add_7_25_groupi_n_1777 ,csa_tree_add_7_25_groupi_n_1776);
  not csa_tree_add_7_25_groupi_drc_bufs21856(csa_tree_add_7_25_groupi_n_1776 ,csa_tree_add_7_25_groupi_n_2866);
  not csa_tree_add_7_25_groupi_drc_bufs21858(csa_tree_add_7_25_groupi_n_1775 ,csa_tree_add_7_25_groupi_n_1773);
  not csa_tree_add_7_25_groupi_drc_bufs21859(csa_tree_add_7_25_groupi_n_1774 ,csa_tree_add_7_25_groupi_n_1773);
  not csa_tree_add_7_25_groupi_drc_bufs21860(csa_tree_add_7_25_groupi_n_1773 ,csa_tree_add_7_25_groupi_n_3529);
  not csa_tree_add_7_25_groupi_drc_bufs21862(csa_tree_add_7_25_groupi_n_1772 ,csa_tree_add_7_25_groupi_n_1770);
  not csa_tree_add_7_25_groupi_drc_bufs21863(csa_tree_add_7_25_groupi_n_1771 ,csa_tree_add_7_25_groupi_n_1770);
  not csa_tree_add_7_25_groupi_drc_bufs21864(csa_tree_add_7_25_groupi_n_1770 ,csa_tree_add_7_25_groupi_n_3531);
  not csa_tree_add_7_25_groupi_drc_bufs21866(csa_tree_add_7_25_groupi_n_1769 ,csa_tree_add_7_25_groupi_n_1767);
  not csa_tree_add_7_25_groupi_drc_bufs21867(csa_tree_add_7_25_groupi_n_1768 ,csa_tree_add_7_25_groupi_n_1767);
  not csa_tree_add_7_25_groupi_drc_bufs21868(csa_tree_add_7_25_groupi_n_1767 ,csa_tree_add_7_25_groupi_n_2877);
  not csa_tree_add_7_25_groupi_drc_bufs21870(csa_tree_add_7_25_groupi_n_1766 ,csa_tree_add_7_25_groupi_n_1764);
  not csa_tree_add_7_25_groupi_drc_bufs21871(csa_tree_add_7_25_groupi_n_1765 ,csa_tree_add_7_25_groupi_n_1764);
  not csa_tree_add_7_25_groupi_drc_bufs21872(csa_tree_add_7_25_groupi_n_1764 ,csa_tree_add_7_25_groupi_n_2876);
  not csa_tree_add_7_25_groupi_drc_bufs21874(csa_tree_add_7_25_groupi_n_1763 ,csa_tree_add_7_25_groupi_n_1761);
  not csa_tree_add_7_25_groupi_drc_bufs21875(csa_tree_add_7_25_groupi_n_1762 ,csa_tree_add_7_25_groupi_n_1761);
  not csa_tree_add_7_25_groupi_drc_bufs21876(csa_tree_add_7_25_groupi_n_1761 ,csa_tree_add_7_25_groupi_n_2876);
  not csa_tree_add_7_25_groupi_drc_bufs21878(csa_tree_add_7_25_groupi_n_1760 ,csa_tree_add_7_25_groupi_n_1758);
  not csa_tree_add_7_25_groupi_drc_bufs21879(csa_tree_add_7_25_groupi_n_1759 ,csa_tree_add_7_25_groupi_n_1758);
  not csa_tree_add_7_25_groupi_drc_bufs21880(csa_tree_add_7_25_groupi_n_1758 ,csa_tree_add_7_25_groupi_n_2794);
  not csa_tree_add_7_25_groupi_drc_bufs21882(csa_tree_add_7_25_groupi_n_1757 ,csa_tree_add_7_25_groupi_n_1755);
  not csa_tree_add_7_25_groupi_drc_bufs21883(csa_tree_add_7_25_groupi_n_1756 ,csa_tree_add_7_25_groupi_n_1755);
  not csa_tree_add_7_25_groupi_drc_bufs21884(csa_tree_add_7_25_groupi_n_1755 ,csa_tree_add_7_25_groupi_n_2875);
  not csa_tree_add_7_25_groupi_drc_bufs21886(csa_tree_add_7_25_groupi_n_1754 ,csa_tree_add_7_25_groupi_n_1752);
  not csa_tree_add_7_25_groupi_drc_bufs21887(csa_tree_add_7_25_groupi_n_1753 ,csa_tree_add_7_25_groupi_n_1752);
  not csa_tree_add_7_25_groupi_drc_bufs21888(csa_tree_add_7_25_groupi_n_1752 ,csa_tree_add_7_25_groupi_n_2795);
  not csa_tree_add_7_25_groupi_drc_bufs21890(csa_tree_add_7_25_groupi_n_1751 ,csa_tree_add_7_25_groupi_n_1749);
  not csa_tree_add_7_25_groupi_drc_bufs21891(csa_tree_add_7_25_groupi_n_1750 ,csa_tree_add_7_25_groupi_n_1749);
  not csa_tree_add_7_25_groupi_drc_bufs21892(csa_tree_add_7_25_groupi_n_1749 ,csa_tree_add_7_25_groupi_n_2795);
  not csa_tree_add_7_25_groupi_drc_bufs21894(csa_tree_add_7_25_groupi_n_1748 ,csa_tree_add_7_25_groupi_n_1746);
  not csa_tree_add_7_25_groupi_drc_bufs21895(csa_tree_add_7_25_groupi_n_1747 ,csa_tree_add_7_25_groupi_n_1746);
  not csa_tree_add_7_25_groupi_drc_bufs21896(csa_tree_add_7_25_groupi_n_1746 ,csa_tree_add_7_25_groupi_n_2794);
  not csa_tree_add_7_25_groupi_drc_bufs21898(csa_tree_add_7_25_groupi_n_1745 ,csa_tree_add_7_25_groupi_n_1743);
  not csa_tree_add_7_25_groupi_drc_bufs21899(csa_tree_add_7_25_groupi_n_1744 ,csa_tree_add_7_25_groupi_n_1743);
  not csa_tree_add_7_25_groupi_drc_bufs21900(csa_tree_add_7_25_groupi_n_1743 ,csa_tree_add_7_25_groupi_n_3530);
  not csa_tree_add_7_25_groupi_drc_bufs21902(csa_tree_add_7_25_groupi_n_1742 ,csa_tree_add_7_25_groupi_n_1740);
  not csa_tree_add_7_25_groupi_drc_bufs21903(csa_tree_add_7_25_groupi_n_1741 ,csa_tree_add_7_25_groupi_n_1740);
  not csa_tree_add_7_25_groupi_drc_bufs21904(csa_tree_add_7_25_groupi_n_1740 ,csa_tree_add_7_25_groupi_n_2877);
  not csa_tree_add_7_25_groupi_drc_bufs21906(csa_tree_add_7_25_groupi_n_1739 ,csa_tree_add_7_25_groupi_n_1737);
  not csa_tree_add_7_25_groupi_drc_bufs21907(csa_tree_add_7_25_groupi_n_1738 ,csa_tree_add_7_25_groupi_n_1737);
  not csa_tree_add_7_25_groupi_drc_bufs21908(csa_tree_add_7_25_groupi_n_1737 ,csa_tree_add_7_25_groupi_n_2871);
  not csa_tree_add_7_25_groupi_drc_bufs21910(csa_tree_add_7_25_groupi_n_1736 ,csa_tree_add_7_25_groupi_n_1734);
  not csa_tree_add_7_25_groupi_drc_bufs21911(csa_tree_add_7_25_groupi_n_1735 ,csa_tree_add_7_25_groupi_n_1734);
  not csa_tree_add_7_25_groupi_drc_bufs21912(csa_tree_add_7_25_groupi_n_1734 ,csa_tree_add_7_25_groupi_n_2872);
  not csa_tree_add_7_25_groupi_drc_bufs21914(csa_tree_add_7_25_groupi_n_1733 ,csa_tree_add_7_25_groupi_n_1731);
  not csa_tree_add_7_25_groupi_drc_bufs21915(csa_tree_add_7_25_groupi_n_1732 ,csa_tree_add_7_25_groupi_n_1731);
  not csa_tree_add_7_25_groupi_drc_bufs21916(csa_tree_add_7_25_groupi_n_1731 ,csa_tree_add_7_25_groupi_n_3530);
  not csa_tree_add_7_25_groupi_drc_bufs21918(csa_tree_add_7_25_groupi_n_1730 ,csa_tree_add_7_25_groupi_n_1728);
  not csa_tree_add_7_25_groupi_drc_bufs21919(csa_tree_add_7_25_groupi_n_1729 ,csa_tree_add_7_25_groupi_n_1728);
  not csa_tree_add_7_25_groupi_drc_bufs21920(csa_tree_add_7_25_groupi_n_1728 ,csa_tree_add_7_25_groupi_n_2871);
  not csa_tree_add_7_25_groupi_drc_bufs21922(csa_tree_add_7_25_groupi_n_1727 ,csa_tree_add_7_25_groupi_n_1725);
  not csa_tree_add_7_25_groupi_drc_bufs21923(csa_tree_add_7_25_groupi_n_1726 ,csa_tree_add_7_25_groupi_n_1725);
  not csa_tree_add_7_25_groupi_drc_bufs21924(csa_tree_add_7_25_groupi_n_1725 ,csa_tree_add_7_25_groupi_n_3529);
  not csa_tree_add_7_25_groupi_drc_bufs21926(csa_tree_add_7_25_groupi_n_1724 ,csa_tree_add_7_25_groupi_n_1722);
  not csa_tree_add_7_25_groupi_drc_bufs21927(csa_tree_add_7_25_groupi_n_1723 ,csa_tree_add_7_25_groupi_n_1722);
  not csa_tree_add_7_25_groupi_drc_bufs21928(csa_tree_add_7_25_groupi_n_1722 ,csa_tree_add_7_25_groupi_n_2875);
  not csa_tree_add_7_25_groupi_drc_bufs21930(csa_tree_add_7_25_groupi_n_1721 ,csa_tree_add_7_25_groupi_n_1719);
  not csa_tree_add_7_25_groupi_drc_bufs21931(csa_tree_add_7_25_groupi_n_1720 ,csa_tree_add_7_25_groupi_n_1719);
  not csa_tree_add_7_25_groupi_drc_bufs21932(csa_tree_add_7_25_groupi_n_1719 ,csa_tree_add_7_25_groupi_n_2796);
  not csa_tree_add_7_25_groupi_drc_bufs21934(csa_tree_add_7_25_groupi_n_1718 ,csa_tree_add_7_25_groupi_n_1716);
  not csa_tree_add_7_25_groupi_drc_bufs21935(csa_tree_add_7_25_groupi_n_1717 ,csa_tree_add_7_25_groupi_n_1716);
  not csa_tree_add_7_25_groupi_drc_bufs21936(csa_tree_add_7_25_groupi_n_1716 ,csa_tree_add_7_25_groupi_n_2872);
  not csa_tree_add_7_25_groupi_drc_bufs21938(csa_tree_add_7_25_groupi_n_1715 ,csa_tree_add_7_25_groupi_n_1713);
  not csa_tree_add_7_25_groupi_drc_bufs21939(csa_tree_add_7_25_groupi_n_1714 ,csa_tree_add_7_25_groupi_n_1713);
  not csa_tree_add_7_25_groupi_drc_bufs21940(csa_tree_add_7_25_groupi_n_1713 ,csa_tree_add_7_25_groupi_n_3518);
  not csa_tree_add_7_25_groupi_drc_bufs21942(csa_tree_add_7_25_groupi_n_1712 ,csa_tree_add_7_25_groupi_n_1710);
  not csa_tree_add_7_25_groupi_drc_bufs21943(csa_tree_add_7_25_groupi_n_1711 ,csa_tree_add_7_25_groupi_n_1710);
  not csa_tree_add_7_25_groupi_drc_bufs21944(csa_tree_add_7_25_groupi_n_1710 ,csa_tree_add_7_25_groupi_n_2865);
  not csa_tree_add_7_25_groupi_drc_bufs21946(csa_tree_add_7_25_groupi_n_1709 ,csa_tree_add_7_25_groupi_n_1707);
  not csa_tree_add_7_25_groupi_drc_bufs21947(csa_tree_add_7_25_groupi_n_1708 ,csa_tree_add_7_25_groupi_n_1707);
  not csa_tree_add_7_25_groupi_drc_bufs21948(csa_tree_add_7_25_groupi_n_1707 ,csa_tree_add_7_25_groupi_n_2685);
  not csa_tree_add_7_25_groupi_drc_bufs21950(csa_tree_add_7_25_groupi_n_1706 ,csa_tree_add_7_25_groupi_n_1704);
  not csa_tree_add_7_25_groupi_drc_bufs21951(csa_tree_add_7_25_groupi_n_1705 ,csa_tree_add_7_25_groupi_n_1704);
  not csa_tree_add_7_25_groupi_drc_bufs21952(csa_tree_add_7_25_groupi_n_1704 ,csa_tree_add_7_25_groupi_n_2685);
  not csa_tree_add_7_25_groupi_drc_bufs21954(csa_tree_add_7_25_groupi_n_1703 ,csa_tree_add_7_25_groupi_n_1701);
  not csa_tree_add_7_25_groupi_drc_bufs21955(csa_tree_add_7_25_groupi_n_1702 ,csa_tree_add_7_25_groupi_n_1701);
  not csa_tree_add_7_25_groupi_drc_bufs21956(csa_tree_add_7_25_groupi_n_1701 ,csa_tree_add_7_25_groupi_n_2683);
  not csa_tree_add_7_25_groupi_drc_bufs21958(csa_tree_add_7_25_groupi_n_1700 ,csa_tree_add_7_25_groupi_n_1698);
  not csa_tree_add_7_25_groupi_drc_bufs21959(csa_tree_add_7_25_groupi_n_1699 ,csa_tree_add_7_25_groupi_n_1698);
  not csa_tree_add_7_25_groupi_drc_bufs21960(csa_tree_add_7_25_groupi_n_1698 ,csa_tree_add_7_25_groupi_n_2859);
  not csa_tree_add_7_25_groupi_drc_bufs21962(csa_tree_add_7_25_groupi_n_1697 ,csa_tree_add_7_25_groupi_n_1695);
  not csa_tree_add_7_25_groupi_drc_bufs21963(csa_tree_add_7_25_groupi_n_1696 ,csa_tree_add_7_25_groupi_n_1695);
  not csa_tree_add_7_25_groupi_drc_bufs21964(csa_tree_add_7_25_groupi_n_1695 ,csa_tree_add_7_25_groupi_n_2683);
  not csa_tree_add_7_25_groupi_drc_bufs21966(csa_tree_add_7_25_groupi_n_1694 ,csa_tree_add_7_25_groupi_n_1692);
  not csa_tree_add_7_25_groupi_drc_bufs21967(csa_tree_add_7_25_groupi_n_1693 ,csa_tree_add_7_25_groupi_n_1692);
  not csa_tree_add_7_25_groupi_drc_bufs21968(csa_tree_add_7_25_groupi_n_1692 ,csa_tree_add_7_25_groupi_n_2682);
  not csa_tree_add_7_25_groupi_drc_bufs21970(csa_tree_add_7_25_groupi_n_1691 ,csa_tree_add_7_25_groupi_n_1689);
  not csa_tree_add_7_25_groupi_drc_bufs21971(csa_tree_add_7_25_groupi_n_1690 ,csa_tree_add_7_25_groupi_n_1689);
  not csa_tree_add_7_25_groupi_drc_bufs21972(csa_tree_add_7_25_groupi_n_1689 ,csa_tree_add_7_25_groupi_n_2682);
  not csa_tree_add_7_25_groupi_drc_bufs21974(csa_tree_add_7_25_groupi_n_1688 ,csa_tree_add_7_25_groupi_n_1686);
  not csa_tree_add_7_25_groupi_drc_bufs21975(csa_tree_add_7_25_groupi_n_1687 ,csa_tree_add_7_25_groupi_n_1686);
  not csa_tree_add_7_25_groupi_drc_bufs21976(csa_tree_add_7_25_groupi_n_1686 ,csa_tree_add_7_25_groupi_n_2686);
  not csa_tree_add_7_25_groupi_drc_bufs21978(csa_tree_add_7_25_groupi_n_1685 ,csa_tree_add_7_25_groupi_n_1683);
  not csa_tree_add_7_25_groupi_drc_bufs21979(csa_tree_add_7_25_groupi_n_1684 ,csa_tree_add_7_25_groupi_n_1683);
  not csa_tree_add_7_25_groupi_drc_bufs21980(csa_tree_add_7_25_groupi_n_1683 ,csa_tree_add_7_25_groupi_n_2843);
  not csa_tree_add_7_25_groupi_drc_bufs21982(csa_tree_add_7_25_groupi_n_1682 ,csa_tree_add_7_25_groupi_n_1680);
  not csa_tree_add_7_25_groupi_drc_bufs21983(csa_tree_add_7_25_groupi_n_1681 ,csa_tree_add_7_25_groupi_n_1680);
  not csa_tree_add_7_25_groupi_drc_bufs21984(csa_tree_add_7_25_groupi_n_1680 ,csa_tree_add_7_25_groupi_n_2843);
  not csa_tree_add_7_25_groupi_drc_bufs21986(csa_tree_add_7_25_groupi_n_1679 ,csa_tree_add_7_25_groupi_n_1677);
  not csa_tree_add_7_25_groupi_drc_bufs21987(csa_tree_add_7_25_groupi_n_1678 ,csa_tree_add_7_25_groupi_n_1677);
  not csa_tree_add_7_25_groupi_drc_bufs21988(csa_tree_add_7_25_groupi_n_1677 ,csa_tree_add_7_25_groupi_n_3499);
  not csa_tree_add_7_25_groupi_drc_bufs21990(csa_tree_add_7_25_groupi_n_1676 ,csa_tree_add_7_25_groupi_n_1674);
  not csa_tree_add_7_25_groupi_drc_bufs21991(csa_tree_add_7_25_groupi_n_1675 ,csa_tree_add_7_25_groupi_n_1674);
  not csa_tree_add_7_25_groupi_drc_bufs21992(csa_tree_add_7_25_groupi_n_1674 ,csa_tree_add_7_25_groupi_n_2860);
  not csa_tree_add_7_25_groupi_drc_bufs21994(csa_tree_add_7_25_groupi_n_1673 ,csa_tree_add_7_25_groupi_n_1671);
  not csa_tree_add_7_25_groupi_drc_bufs21995(csa_tree_add_7_25_groupi_n_1672 ,csa_tree_add_7_25_groupi_n_1671);
  not csa_tree_add_7_25_groupi_drc_bufs21996(csa_tree_add_7_25_groupi_n_1671 ,csa_tree_add_7_25_groupi_n_2841);
  not csa_tree_add_7_25_groupi_drc_bufs21998(csa_tree_add_7_25_groupi_n_1670 ,csa_tree_add_7_25_groupi_n_1668);
  not csa_tree_add_7_25_groupi_drc_bufs21999(csa_tree_add_7_25_groupi_n_1669 ,csa_tree_add_7_25_groupi_n_1668);
  not csa_tree_add_7_25_groupi_drc_bufs22000(csa_tree_add_7_25_groupi_n_1668 ,csa_tree_add_7_25_groupi_n_2840);
  not csa_tree_add_7_25_groupi_drc_bufs22002(csa_tree_add_7_25_groupi_n_1667 ,csa_tree_add_7_25_groupi_n_1665);
  not csa_tree_add_7_25_groupi_drc_bufs22003(csa_tree_add_7_25_groupi_n_1666 ,csa_tree_add_7_25_groupi_n_1665);
  not csa_tree_add_7_25_groupi_drc_bufs22004(csa_tree_add_7_25_groupi_n_1665 ,csa_tree_add_7_25_groupi_n_2840);
  not csa_tree_add_7_25_groupi_drc_bufs22006(csa_tree_add_7_25_groupi_n_1664 ,csa_tree_add_7_25_groupi_n_1662);
  not csa_tree_add_7_25_groupi_drc_bufs22007(csa_tree_add_7_25_groupi_n_1663 ,csa_tree_add_7_25_groupi_n_1662);
  not csa_tree_add_7_25_groupi_drc_bufs22008(csa_tree_add_7_25_groupi_n_1662 ,csa_tree_add_7_25_groupi_n_2777);
  not csa_tree_add_7_25_groupi_drc_bufs22010(csa_tree_add_7_25_groupi_n_1661 ,csa_tree_add_7_25_groupi_n_1659);
  not csa_tree_add_7_25_groupi_drc_bufs22011(csa_tree_add_7_25_groupi_n_1660 ,csa_tree_add_7_25_groupi_n_1659);
  not csa_tree_add_7_25_groupi_drc_bufs22012(csa_tree_add_7_25_groupi_n_1659 ,csa_tree_add_7_25_groupi_n_2775);
  not csa_tree_add_7_25_groupi_drc_bufs22014(csa_tree_add_7_25_groupi_n_1658 ,csa_tree_add_7_25_groupi_n_1656);
  not csa_tree_add_7_25_groupi_drc_bufs22015(csa_tree_add_7_25_groupi_n_1657 ,csa_tree_add_7_25_groupi_n_1656);
  not csa_tree_add_7_25_groupi_drc_bufs22016(csa_tree_add_7_25_groupi_n_1656 ,csa_tree_add_7_25_groupi_n_2775);
  not csa_tree_add_7_25_groupi_drc_bufs22018(csa_tree_add_7_25_groupi_n_1655 ,csa_tree_add_7_25_groupi_n_1653);
  not csa_tree_add_7_25_groupi_drc_bufs22019(csa_tree_add_7_25_groupi_n_1654 ,csa_tree_add_7_25_groupi_n_1653);
  not csa_tree_add_7_25_groupi_drc_bufs22020(csa_tree_add_7_25_groupi_n_1653 ,csa_tree_add_7_25_groupi_n_2774);
  not csa_tree_add_7_25_groupi_drc_bufs22022(csa_tree_add_7_25_groupi_n_1652 ,csa_tree_add_7_25_groupi_n_1650);
  not csa_tree_add_7_25_groupi_drc_bufs22023(csa_tree_add_7_25_groupi_n_1651 ,csa_tree_add_7_25_groupi_n_1650);
  not csa_tree_add_7_25_groupi_drc_bufs22024(csa_tree_add_7_25_groupi_n_1650 ,csa_tree_add_7_25_groupi_n_2772);
  not csa_tree_add_7_25_groupi_drc_bufs22026(csa_tree_add_7_25_groupi_n_1649 ,csa_tree_add_7_25_groupi_n_1647);
  not csa_tree_add_7_25_groupi_drc_bufs22027(csa_tree_add_7_25_groupi_n_1648 ,csa_tree_add_7_25_groupi_n_1647);
  not csa_tree_add_7_25_groupi_drc_bufs22028(csa_tree_add_7_25_groupi_n_1647 ,csa_tree_add_7_25_groupi_n_2772);
  not csa_tree_add_7_25_groupi_drc_bufs22030(csa_tree_add_7_25_groupi_n_1646 ,csa_tree_add_7_25_groupi_n_1644);
  not csa_tree_add_7_25_groupi_drc_bufs22031(csa_tree_add_7_25_groupi_n_1645 ,csa_tree_add_7_25_groupi_n_1644);
  not csa_tree_add_7_25_groupi_drc_bufs22032(csa_tree_add_7_25_groupi_n_1644 ,csa_tree_add_7_25_groupi_n_2770);
  not csa_tree_add_7_25_groupi_drc_bufs22034(csa_tree_add_7_25_groupi_n_1643 ,csa_tree_add_7_25_groupi_n_1641);
  not csa_tree_add_7_25_groupi_drc_bufs22035(csa_tree_add_7_25_groupi_n_1642 ,csa_tree_add_7_25_groupi_n_1641);
  not csa_tree_add_7_25_groupi_drc_bufs22036(csa_tree_add_7_25_groupi_n_1641 ,csa_tree_add_7_25_groupi_n_2769);
  not csa_tree_add_7_25_groupi_drc_bufs22038(csa_tree_add_7_25_groupi_n_1640 ,csa_tree_add_7_25_groupi_n_1638);
  not csa_tree_add_7_25_groupi_drc_bufs22039(csa_tree_add_7_25_groupi_n_1639 ,csa_tree_add_7_25_groupi_n_1638);
  not csa_tree_add_7_25_groupi_drc_bufs22040(csa_tree_add_7_25_groupi_n_1638 ,csa_tree_add_7_25_groupi_n_2769);
  not csa_tree_add_7_25_groupi_drc_bufs22042(csa_tree_add_7_25_groupi_n_1637 ,csa_tree_add_7_25_groupi_n_1635);
  not csa_tree_add_7_25_groupi_drc_bufs22043(csa_tree_add_7_25_groupi_n_1636 ,csa_tree_add_7_25_groupi_n_1635);
  not csa_tree_add_7_25_groupi_drc_bufs22044(csa_tree_add_7_25_groupi_n_1635 ,csa_tree_add_7_25_groupi_n_3517);
  not csa_tree_add_7_25_groupi_drc_bufs22046(csa_tree_add_7_25_groupi_n_1634 ,csa_tree_add_7_25_groupi_n_1632);
  not csa_tree_add_7_25_groupi_drc_bufs22047(csa_tree_add_7_25_groupi_n_1633 ,csa_tree_add_7_25_groupi_n_1632);
  not csa_tree_add_7_25_groupi_drc_bufs22048(csa_tree_add_7_25_groupi_n_1632 ,csa_tree_add_7_25_groupi_n_2767);
  not csa_tree_add_7_25_groupi_drc_bufs22050(csa_tree_add_7_25_groupi_n_1631 ,csa_tree_add_7_25_groupi_n_1629);
  not csa_tree_add_7_25_groupi_drc_bufs22051(csa_tree_add_7_25_groupi_n_1630 ,csa_tree_add_7_25_groupi_n_1629);
  not csa_tree_add_7_25_groupi_drc_bufs22052(csa_tree_add_7_25_groupi_n_1629 ,csa_tree_add_7_25_groupi_n_2765);
  not csa_tree_add_7_25_groupi_drc_bufs22054(csa_tree_add_7_25_groupi_n_1628 ,csa_tree_add_7_25_groupi_n_1626);
  not csa_tree_add_7_25_groupi_drc_bufs22055(csa_tree_add_7_25_groupi_n_1627 ,csa_tree_add_7_25_groupi_n_1626);
  not csa_tree_add_7_25_groupi_drc_bufs22056(csa_tree_add_7_25_groupi_n_1626 ,csa_tree_add_7_25_groupi_n_2765);
  not csa_tree_add_7_25_groupi_drc_bufs22058(csa_tree_add_7_25_groupi_n_1625 ,csa_tree_add_7_25_groupi_n_1623);
  not csa_tree_add_7_25_groupi_drc_bufs22059(csa_tree_add_7_25_groupi_n_1624 ,csa_tree_add_7_25_groupi_n_1623);
  not csa_tree_add_7_25_groupi_drc_bufs22060(csa_tree_add_7_25_groupi_n_1623 ,csa_tree_add_7_25_groupi_n_2764);
  not csa_tree_add_7_25_groupi_drc_bufs22062(csa_tree_add_7_25_groupi_n_1622 ,csa_tree_add_7_25_groupi_n_1620);
  not csa_tree_add_7_25_groupi_drc_bufs22063(csa_tree_add_7_25_groupi_n_1621 ,csa_tree_add_7_25_groupi_n_1620);
  not csa_tree_add_7_25_groupi_drc_bufs22064(csa_tree_add_7_25_groupi_n_1620 ,csa_tree_add_7_25_groupi_n_2764);
  not csa_tree_add_7_25_groupi_drc_bufs22066(csa_tree_add_7_25_groupi_n_1619 ,csa_tree_add_7_25_groupi_n_1617);
  not csa_tree_add_7_25_groupi_drc_bufs22067(csa_tree_add_7_25_groupi_n_1618 ,csa_tree_add_7_25_groupi_n_1617);
  not csa_tree_add_7_25_groupi_drc_bufs22068(csa_tree_add_7_25_groupi_n_1617 ,csa_tree_add_7_25_groupi_n_2762);
  not csa_tree_add_7_25_groupi_drc_bufs22070(csa_tree_add_7_25_groupi_n_1616 ,csa_tree_add_7_25_groupi_n_1614);
  not csa_tree_add_7_25_groupi_drc_bufs22071(csa_tree_add_7_25_groupi_n_1615 ,csa_tree_add_7_25_groupi_n_1614);
  not csa_tree_add_7_25_groupi_drc_bufs22072(csa_tree_add_7_25_groupi_n_1614 ,csa_tree_add_7_25_groupi_n_2762);
  not csa_tree_add_7_25_groupi_drc_bufs22074(csa_tree_add_7_25_groupi_n_1613 ,csa_tree_add_7_25_groupi_n_1611);
  not csa_tree_add_7_25_groupi_drc_bufs22075(csa_tree_add_7_25_groupi_n_1612 ,csa_tree_add_7_25_groupi_n_1611);
  not csa_tree_add_7_25_groupi_drc_bufs22076(csa_tree_add_7_25_groupi_n_1611 ,csa_tree_add_7_25_groupi_n_2759);
  not csa_tree_add_7_25_groupi_drc_bufs22078(csa_tree_add_7_25_groupi_n_1610 ,csa_tree_add_7_25_groupi_n_1608);
  not csa_tree_add_7_25_groupi_drc_bufs22079(csa_tree_add_7_25_groupi_n_1609 ,csa_tree_add_7_25_groupi_n_1608);
  not csa_tree_add_7_25_groupi_drc_bufs22080(csa_tree_add_7_25_groupi_n_1608 ,csa_tree_add_7_25_groupi_n_2757);
  not csa_tree_add_7_25_groupi_drc_bufs22082(csa_tree_add_7_25_groupi_n_1607 ,csa_tree_add_7_25_groupi_n_1605);
  not csa_tree_add_7_25_groupi_drc_bufs22083(csa_tree_add_7_25_groupi_n_1606 ,csa_tree_add_7_25_groupi_n_1605);
  not csa_tree_add_7_25_groupi_drc_bufs22084(csa_tree_add_7_25_groupi_n_1605 ,csa_tree_add_7_25_groupi_n_2757);
  not csa_tree_add_7_25_groupi_drc_bufs22086(csa_tree_add_7_25_groupi_n_1604 ,csa_tree_add_7_25_groupi_n_1602);
  not csa_tree_add_7_25_groupi_drc_bufs22087(csa_tree_add_7_25_groupi_n_1603 ,csa_tree_add_7_25_groupi_n_1602);
  not csa_tree_add_7_25_groupi_drc_bufs22088(csa_tree_add_7_25_groupi_n_1602 ,csa_tree_add_7_25_groupi_n_2754);
  not csa_tree_add_7_25_groupi_drc_bufs22090(csa_tree_add_7_25_groupi_n_1601 ,csa_tree_add_7_25_groupi_n_1599);
  not csa_tree_add_7_25_groupi_drc_bufs22091(csa_tree_add_7_25_groupi_n_1600 ,csa_tree_add_7_25_groupi_n_1599);
  not csa_tree_add_7_25_groupi_drc_bufs22092(csa_tree_add_7_25_groupi_n_1599 ,csa_tree_add_7_25_groupi_n_2755);
  not csa_tree_add_7_25_groupi_drc_bufs22094(csa_tree_add_7_25_groupi_n_1598 ,csa_tree_add_7_25_groupi_n_1596);
  not csa_tree_add_7_25_groupi_drc_bufs22095(csa_tree_add_7_25_groupi_n_1597 ,csa_tree_add_7_25_groupi_n_1596);
  not csa_tree_add_7_25_groupi_drc_bufs22096(csa_tree_add_7_25_groupi_n_1596 ,csa_tree_add_7_25_groupi_n_3502);
  not csa_tree_add_7_25_groupi_drc_bufs22098(csa_tree_add_7_25_groupi_n_1595 ,csa_tree_add_7_25_groupi_n_1593);
  not csa_tree_add_7_25_groupi_drc_bufs22099(csa_tree_add_7_25_groupi_n_1594 ,csa_tree_add_7_25_groupi_n_1593);
  not csa_tree_add_7_25_groupi_drc_bufs22100(csa_tree_add_7_25_groupi_n_1593 ,csa_tree_add_7_25_groupi_n_2760);
  not csa_tree_add_7_25_groupi_drc_bufs22102(csa_tree_add_7_25_groupi_n_1592 ,csa_tree_add_7_25_groupi_n_1590);
  not csa_tree_add_7_25_groupi_drc_bufs22103(csa_tree_add_7_25_groupi_n_1591 ,csa_tree_add_7_25_groupi_n_1590);
  not csa_tree_add_7_25_groupi_drc_bufs22104(csa_tree_add_7_25_groupi_n_1590 ,csa_tree_add_7_25_groupi_n_2521);
  not csa_tree_add_7_25_groupi_drc_bufs22106(csa_tree_add_7_25_groupi_n_1589 ,csa_tree_add_7_25_groupi_n_1587);
  not csa_tree_add_7_25_groupi_drc_bufs22107(csa_tree_add_7_25_groupi_n_1588 ,csa_tree_add_7_25_groupi_n_1587);
  not csa_tree_add_7_25_groupi_drc_bufs22108(csa_tree_add_7_25_groupi_n_1587 ,csa_tree_add_7_25_groupi_n_2521);
  not csa_tree_add_7_25_groupi_drc_bufs22110(csa_tree_add_7_25_groupi_n_1586 ,csa_tree_add_7_25_groupi_n_1584);
  not csa_tree_add_7_25_groupi_drc_bufs22111(csa_tree_add_7_25_groupi_n_1585 ,csa_tree_add_7_25_groupi_n_1584);
  not csa_tree_add_7_25_groupi_drc_bufs22112(csa_tree_add_7_25_groupi_n_1584 ,csa_tree_add_7_25_groupi_n_2519);
  not csa_tree_add_7_25_groupi_drc_bufs22114(csa_tree_add_7_25_groupi_n_1583 ,csa_tree_add_7_25_groupi_n_1581);
  not csa_tree_add_7_25_groupi_drc_bufs22115(csa_tree_add_7_25_groupi_n_1582 ,csa_tree_add_7_25_groupi_n_1581);
  not csa_tree_add_7_25_groupi_drc_bufs22116(csa_tree_add_7_25_groupi_n_1581 ,csa_tree_add_7_25_groupi_n_2519);
  not csa_tree_add_7_25_groupi_drc_bufs22118(csa_tree_add_7_25_groupi_n_1580 ,csa_tree_add_7_25_groupi_n_1578);
  not csa_tree_add_7_25_groupi_drc_bufs22119(csa_tree_add_7_25_groupi_n_1579 ,csa_tree_add_7_25_groupi_n_1578);
  not csa_tree_add_7_25_groupi_drc_bufs22120(csa_tree_add_7_25_groupi_n_1578 ,csa_tree_add_7_25_groupi_n_2518);
  not csa_tree_add_7_25_groupi_drc_bufs22122(csa_tree_add_7_25_groupi_n_1577 ,csa_tree_add_7_25_groupi_n_1575);
  not csa_tree_add_7_25_groupi_drc_bufs22123(csa_tree_add_7_25_groupi_n_1576 ,csa_tree_add_7_25_groupi_n_1575);
  not csa_tree_add_7_25_groupi_drc_bufs22124(csa_tree_add_7_25_groupi_n_1575 ,csa_tree_add_7_25_groupi_n_2518);
  not csa_tree_add_7_25_groupi_drc_bufs22126(csa_tree_add_7_25_groupi_n_1574 ,csa_tree_add_7_25_groupi_n_1572);
  not csa_tree_add_7_25_groupi_drc_bufs22127(csa_tree_add_7_25_groupi_n_1573 ,csa_tree_add_7_25_groupi_n_1572);
  not csa_tree_add_7_25_groupi_drc_bufs22128(csa_tree_add_7_25_groupi_n_1572 ,csa_tree_add_7_25_groupi_n_2522);
  not csa_tree_add_7_25_groupi_drc_bufs22130(csa_tree_add_7_25_groupi_n_1571 ,csa_tree_add_7_25_groupi_n_1569);
  not csa_tree_add_7_25_groupi_drc_bufs22131(csa_tree_add_7_25_groupi_n_1570 ,csa_tree_add_7_25_groupi_n_1569);
  not csa_tree_add_7_25_groupi_drc_bufs22132(csa_tree_add_7_25_groupi_n_1569 ,csa_tree_add_7_25_groupi_n_3524);
  not csa_tree_add_7_25_groupi_drc_bufs22134(csa_tree_add_7_25_groupi_n_1568 ,csa_tree_add_7_25_groupi_n_1566);
  not csa_tree_add_7_25_groupi_drc_bufs22135(csa_tree_add_7_25_groupi_n_1567 ,csa_tree_add_7_25_groupi_n_1566);
  not csa_tree_add_7_25_groupi_drc_bufs22136(csa_tree_add_7_25_groupi_n_1566 ,csa_tree_add_7_25_groupi_n_3524);
  not csa_tree_add_7_25_groupi_drc_bufs22138(csa_tree_add_7_25_groupi_n_1565 ,csa_tree_add_7_25_groupi_n_1563);
  not csa_tree_add_7_25_groupi_drc_bufs22139(csa_tree_add_7_25_groupi_n_1564 ,csa_tree_add_7_25_groupi_n_1563);
  not csa_tree_add_7_25_groupi_drc_bufs22140(csa_tree_add_7_25_groupi_n_1563 ,csa_tree_add_7_25_groupi_n_3518);
  not csa_tree_add_7_25_groupi_drc_bufs22142(csa_tree_add_7_25_groupi_n_1562 ,csa_tree_add_7_25_groupi_n_1560);
  not csa_tree_add_7_25_groupi_drc_bufs22143(csa_tree_add_7_25_groupi_n_1561 ,csa_tree_add_7_25_groupi_n_1560);
  not csa_tree_add_7_25_groupi_drc_bufs22144(csa_tree_add_7_25_groupi_n_1560 ,csa_tree_add_7_25_groupi_n_2846);
  not csa_tree_add_7_25_groupi_drc_bufs22146(csa_tree_add_7_25_groupi_n_1559 ,csa_tree_add_7_25_groupi_n_1557);
  not csa_tree_add_7_25_groupi_drc_bufs22147(csa_tree_add_7_25_groupi_n_1558 ,csa_tree_add_7_25_groupi_n_1557);
  not csa_tree_add_7_25_groupi_drc_bufs22148(csa_tree_add_7_25_groupi_n_1557 ,csa_tree_add_7_25_groupi_n_3525);
  not csa_tree_add_7_25_groupi_drc_bufs22150(csa_tree_add_7_25_groupi_n_1556 ,csa_tree_add_7_25_groupi_n_1554);
  not csa_tree_add_7_25_groupi_drc_bufs22151(csa_tree_add_7_25_groupi_n_1555 ,csa_tree_add_7_25_groupi_n_1554);
  not csa_tree_add_7_25_groupi_drc_bufs22152(csa_tree_add_7_25_groupi_n_1554 ,csa_tree_add_7_25_groupi_n_3525);
  not csa_tree_add_7_25_groupi_drc_bufs22154(csa_tree_add_7_25_groupi_n_1553 ,csa_tree_add_7_25_groupi_n_1551);
  not csa_tree_add_7_25_groupi_drc_bufs22155(csa_tree_add_7_25_groupi_n_1552 ,csa_tree_add_7_25_groupi_n_1551);
  not csa_tree_add_7_25_groupi_drc_bufs22156(csa_tree_add_7_25_groupi_n_1551 ,csa_tree_add_7_25_groupi_n_2686);
  not csa_tree_add_7_25_groupi_drc_bufs22158(csa_tree_add_7_25_groupi_n_1550 ,csa_tree_add_7_25_groupi_n_1548);
  not csa_tree_add_7_25_groupi_drc_bufs22159(csa_tree_add_7_25_groupi_n_1549 ,csa_tree_add_7_25_groupi_n_1548);
  not csa_tree_add_7_25_groupi_drc_bufs22160(csa_tree_add_7_25_groupi_n_1548 ,csa_tree_add_7_25_groupi_n_2855);
  not csa_tree_add_7_25_groupi_drc_bufs22162(csa_tree_add_7_25_groupi_n_1547 ,csa_tree_add_7_25_groupi_n_1545);
  not csa_tree_add_7_25_groupi_drc_bufs22163(csa_tree_add_7_25_groupi_n_1546 ,csa_tree_add_7_25_groupi_n_1545);
  not csa_tree_add_7_25_groupi_drc_bufs22164(csa_tree_add_7_25_groupi_n_1545 ,csa_tree_add_7_25_groupi_n_3517);
  not csa_tree_add_7_25_groupi_drc_bufs22166(csa_tree_add_7_25_groupi_n_1544 ,csa_tree_add_7_25_groupi_n_1542);
  not csa_tree_add_7_25_groupi_drc_bufs22167(csa_tree_add_7_25_groupi_n_1543 ,csa_tree_add_7_25_groupi_n_1542);
  not csa_tree_add_7_25_groupi_drc_bufs22168(csa_tree_add_7_25_groupi_n_1542 ,csa_tree_add_7_25_groupi_n_3514);
  not csa_tree_add_7_25_groupi_drc_bufs22170(csa_tree_add_7_25_groupi_n_1541 ,csa_tree_add_7_25_groupi_n_1539);
  not csa_tree_add_7_25_groupi_drc_bufs22171(csa_tree_add_7_25_groupi_n_1540 ,csa_tree_add_7_25_groupi_n_1539);
  not csa_tree_add_7_25_groupi_drc_bufs22172(csa_tree_add_7_25_groupi_n_1539 ,csa_tree_add_7_25_groupi_n_3514);
  not csa_tree_add_7_25_groupi_drc_bufs22174(csa_tree_add_7_25_groupi_n_1538 ,csa_tree_add_7_25_groupi_n_1536);
  not csa_tree_add_7_25_groupi_drc_bufs22175(csa_tree_add_7_25_groupi_n_1537 ,csa_tree_add_7_25_groupi_n_1536);
  not csa_tree_add_7_25_groupi_drc_bufs22176(csa_tree_add_7_25_groupi_n_1536 ,csa_tree_add_7_25_groupi_n_3513);
  not csa_tree_add_7_25_groupi_drc_bufs22178(csa_tree_add_7_25_groupi_n_1535 ,csa_tree_add_7_25_groupi_n_1533);
  not csa_tree_add_7_25_groupi_drc_bufs22179(csa_tree_add_7_25_groupi_n_1534 ,csa_tree_add_7_25_groupi_n_1533);
  not csa_tree_add_7_25_groupi_drc_bufs22180(csa_tree_add_7_25_groupi_n_1533 ,csa_tree_add_7_25_groupi_n_3512);
  not csa_tree_add_7_25_groupi_drc_bufs22182(csa_tree_add_7_25_groupi_n_1532 ,csa_tree_add_7_25_groupi_n_1530);
  not csa_tree_add_7_25_groupi_drc_bufs22183(csa_tree_add_7_25_groupi_n_1531 ,csa_tree_add_7_25_groupi_n_1530);
  not csa_tree_add_7_25_groupi_drc_bufs22184(csa_tree_add_7_25_groupi_n_1530 ,csa_tree_add_7_25_groupi_n_2846);
  not csa_tree_add_7_25_groupi_drc_bufs22186(csa_tree_add_7_25_groupi_n_1529 ,csa_tree_add_7_25_groupi_n_1527);
  not csa_tree_add_7_25_groupi_drc_bufs22187(csa_tree_add_7_25_groupi_n_1528 ,csa_tree_add_7_25_groupi_n_1527);
  not csa_tree_add_7_25_groupi_drc_bufs22188(csa_tree_add_7_25_groupi_n_1527 ,csa_tree_add_7_25_groupi_n_3512);
  not csa_tree_add_7_25_groupi_drc_bufs22190(csa_tree_add_7_25_groupi_n_1526 ,csa_tree_add_7_25_groupi_n_1524);
  not csa_tree_add_7_25_groupi_drc_bufs22191(csa_tree_add_7_25_groupi_n_1525 ,csa_tree_add_7_25_groupi_n_1524);
  not csa_tree_add_7_25_groupi_drc_bufs22192(csa_tree_add_7_25_groupi_n_1524 ,csa_tree_add_7_25_groupi_n_2849);
  not csa_tree_add_7_25_groupi_drc_bufs22194(csa_tree_add_7_25_groupi_n_1523 ,csa_tree_add_7_25_groupi_n_1521);
  not csa_tree_add_7_25_groupi_drc_bufs22195(csa_tree_add_7_25_groupi_n_1522 ,csa_tree_add_7_25_groupi_n_1521);
  not csa_tree_add_7_25_groupi_drc_bufs22196(csa_tree_add_7_25_groupi_n_1521 ,csa_tree_add_7_25_groupi_n_2850);
  not csa_tree_add_7_25_groupi_drc_bufs22198(csa_tree_add_7_25_groupi_n_1520 ,csa_tree_add_7_25_groupi_n_1518);
  not csa_tree_add_7_25_groupi_drc_bufs22199(csa_tree_add_7_25_groupi_n_1519 ,csa_tree_add_7_25_groupi_n_1518);
  not csa_tree_add_7_25_groupi_drc_bufs22200(csa_tree_add_7_25_groupi_n_1518 ,csa_tree_add_7_25_groupi_n_2851);
  not csa_tree_add_7_25_groupi_drc_bufs22202(csa_tree_add_7_25_groupi_n_1517 ,csa_tree_add_7_25_groupi_n_1515);
  not csa_tree_add_7_25_groupi_drc_bufs22203(csa_tree_add_7_25_groupi_n_1516 ,csa_tree_add_7_25_groupi_n_1515);
  not csa_tree_add_7_25_groupi_drc_bufs22204(csa_tree_add_7_25_groupi_n_1515 ,csa_tree_add_7_25_groupi_n_3510);
  not csa_tree_add_7_25_groupi_drc_bufs22206(csa_tree_add_7_25_groupi_n_1514 ,csa_tree_add_7_25_groupi_n_1512);
  not csa_tree_add_7_25_groupi_drc_bufs22207(csa_tree_add_7_25_groupi_n_1513 ,csa_tree_add_7_25_groupi_n_1512);
  not csa_tree_add_7_25_groupi_drc_bufs22208(csa_tree_add_7_25_groupi_n_1512 ,csa_tree_add_7_25_groupi_n_3509);
  not csa_tree_add_7_25_groupi_drc_bufs22210(csa_tree_add_7_25_groupi_n_1511 ,csa_tree_add_7_25_groupi_n_1509);
  not csa_tree_add_7_25_groupi_drc_bufs22211(csa_tree_add_7_25_groupi_n_1510 ,csa_tree_add_7_25_groupi_n_1509);
  not csa_tree_add_7_25_groupi_drc_bufs22212(csa_tree_add_7_25_groupi_n_1509 ,csa_tree_add_7_25_groupi_n_2855);
  not csa_tree_add_7_25_groupi_drc_bufs22214(csa_tree_add_7_25_groupi_n_1508 ,csa_tree_add_7_25_groupi_n_1506);
  not csa_tree_add_7_25_groupi_drc_bufs22215(csa_tree_add_7_25_groupi_n_1507 ,csa_tree_add_7_25_groupi_n_1506);
  not csa_tree_add_7_25_groupi_drc_bufs22216(csa_tree_add_7_25_groupi_n_1506 ,csa_tree_add_7_25_groupi_n_2856);
  not csa_tree_add_7_25_groupi_drc_bufs22218(csa_tree_add_7_25_groupi_n_1505 ,csa_tree_add_7_25_groupi_n_1503);
  not csa_tree_add_7_25_groupi_drc_bufs22219(csa_tree_add_7_25_groupi_n_1504 ,csa_tree_add_7_25_groupi_n_1503);
  not csa_tree_add_7_25_groupi_drc_bufs22220(csa_tree_add_7_25_groupi_n_1503 ,csa_tree_add_7_25_groupi_n_3509);
  not csa_tree_add_7_25_groupi_drc_bufs22222(csa_tree_add_7_25_groupi_n_1502 ,csa_tree_add_7_25_groupi_n_1500);
  not csa_tree_add_7_25_groupi_drc_bufs22223(csa_tree_add_7_25_groupi_n_1501 ,csa_tree_add_7_25_groupi_n_1500);
  not csa_tree_add_7_25_groupi_drc_bufs22224(csa_tree_add_7_25_groupi_n_1500 ,csa_tree_add_7_25_groupi_n_2859);
  not csa_tree_add_7_25_groupi_drc_bufs22226(csa_tree_add_7_25_groupi_n_1499 ,csa_tree_add_7_25_groupi_n_1497);
  not csa_tree_add_7_25_groupi_drc_bufs22227(csa_tree_add_7_25_groupi_n_1498 ,csa_tree_add_7_25_groupi_n_1497);
  not csa_tree_add_7_25_groupi_drc_bufs22228(csa_tree_add_7_25_groupi_n_1497 ,csa_tree_add_7_25_groupi_n_2860);
  not csa_tree_add_7_25_groupi_drc_bufs22230(csa_tree_add_7_25_groupi_n_1496 ,csa_tree_add_7_25_groupi_n_1494);
  not csa_tree_add_7_25_groupi_drc_bufs22231(csa_tree_add_7_25_groupi_n_1495 ,csa_tree_add_7_25_groupi_n_1494);
  not csa_tree_add_7_25_groupi_drc_bufs22232(csa_tree_add_7_25_groupi_n_1494 ,csa_tree_add_7_25_groupi_n_3508);
  not csa_tree_add_7_25_groupi_drc_bufs22234(csa_tree_add_7_25_groupi_n_1493 ,csa_tree_add_7_25_groupi_n_1491);
  not csa_tree_add_7_25_groupi_drc_bufs22235(csa_tree_add_7_25_groupi_n_1492 ,csa_tree_add_7_25_groupi_n_1491);
  not csa_tree_add_7_25_groupi_drc_bufs22236(csa_tree_add_7_25_groupi_n_1491 ,csa_tree_add_7_25_groupi_n_3515);
  not csa_tree_add_7_25_groupi_drc_bufs22238(csa_tree_add_7_25_groupi_n_1490 ,csa_tree_add_7_25_groupi_n_1488);
  not csa_tree_add_7_25_groupi_drc_bufs22239(csa_tree_add_7_25_groupi_n_1489 ,csa_tree_add_7_25_groupi_n_1488);
  not csa_tree_add_7_25_groupi_drc_bufs22240(csa_tree_add_7_25_groupi_n_1488 ,csa_tree_add_7_25_groupi_n_2864);
  not csa_tree_add_7_25_groupi_drc_bufs22242(csa_tree_add_7_25_groupi_n_1487 ,csa_tree_add_7_25_groupi_n_1485);
  not csa_tree_add_7_25_groupi_drc_bufs22243(csa_tree_add_7_25_groupi_n_1486 ,csa_tree_add_7_25_groupi_n_1485);
  not csa_tree_add_7_25_groupi_drc_bufs22244(csa_tree_add_7_25_groupi_n_1485 ,csa_tree_add_7_25_groupi_n_2864);
  not csa_tree_add_7_25_groupi_drc_bufs22246(csa_tree_add_7_25_groupi_n_1484 ,csa_tree_add_7_25_groupi_n_1482);
  not csa_tree_add_7_25_groupi_drc_bufs22247(csa_tree_add_7_25_groupi_n_1483 ,csa_tree_add_7_25_groupi_n_1482);
  not csa_tree_add_7_25_groupi_drc_bufs22248(csa_tree_add_7_25_groupi_n_1482 ,csa_tree_add_7_25_groupi_n_3500);
  not csa_tree_add_7_25_groupi_drc_bufs22250(csa_tree_add_7_25_groupi_n_1481 ,csa_tree_add_7_25_groupi_n_1479);
  not csa_tree_add_7_25_groupi_drc_bufs22251(csa_tree_add_7_25_groupi_n_1480 ,csa_tree_add_7_25_groupi_n_1479);
  not csa_tree_add_7_25_groupi_drc_bufs22252(csa_tree_add_7_25_groupi_n_1479 ,csa_tree_add_7_25_groupi_n_3515);
  not csa_tree_add_7_25_groupi_drc_bufs22254(csa_tree_add_7_25_groupi_n_1478 ,csa_tree_add_7_25_groupi_n_1476);
  not csa_tree_add_7_25_groupi_drc_bufs22255(csa_tree_add_7_25_groupi_n_1477 ,csa_tree_add_7_25_groupi_n_1476);
  not csa_tree_add_7_25_groupi_drc_bufs22256(csa_tree_add_7_25_groupi_n_1476 ,csa_tree_add_7_25_groupi_n_3507);
  not csa_tree_add_7_25_groupi_drc_bufs22258(csa_tree_add_7_25_groupi_n_1475 ,csa_tree_add_7_25_groupi_n_1473);
  not csa_tree_add_7_25_groupi_drc_bufs22259(csa_tree_add_7_25_groupi_n_1474 ,csa_tree_add_7_25_groupi_n_1473);
  not csa_tree_add_7_25_groupi_drc_bufs22260(csa_tree_add_7_25_groupi_n_1473 ,csa_tree_add_7_25_groupi_n_3505);
  not csa_tree_add_7_25_groupi_drc_bufs22262(csa_tree_add_7_25_groupi_n_1472 ,csa_tree_add_7_25_groupi_n_1470);
  not csa_tree_add_7_25_groupi_drc_bufs22263(csa_tree_add_7_25_groupi_n_1471 ,csa_tree_add_7_25_groupi_n_1470);
  not csa_tree_add_7_25_groupi_drc_bufs22264(csa_tree_add_7_25_groupi_n_1470 ,csa_tree_add_7_25_groupi_n_3505);
  not csa_tree_add_7_25_groupi_drc_bufs22266(csa_tree_add_7_25_groupi_n_1469 ,csa_tree_add_7_25_groupi_n_1467);
  not csa_tree_add_7_25_groupi_drc_bufs22267(csa_tree_add_7_25_groupi_n_1468 ,csa_tree_add_7_25_groupi_n_1467);
  not csa_tree_add_7_25_groupi_drc_bufs22268(csa_tree_add_7_25_groupi_n_1467 ,csa_tree_add_7_25_groupi_n_3504);
  not csa_tree_add_7_25_groupi_drc_bufs22270(csa_tree_add_7_25_groupi_n_1466 ,csa_tree_add_7_25_groupi_n_1464);
  not csa_tree_add_7_25_groupi_drc_bufs22271(csa_tree_add_7_25_groupi_n_1465 ,csa_tree_add_7_25_groupi_n_1464);
  not csa_tree_add_7_25_groupi_drc_bufs22272(csa_tree_add_7_25_groupi_n_1464 ,csa_tree_add_7_25_groupi_n_3503);
  not csa_tree_add_7_25_groupi_drc_bufs22274(csa_tree_add_7_25_groupi_n_1463 ,csa_tree_add_7_25_groupi_n_1461);
  not csa_tree_add_7_25_groupi_drc_bufs22275(csa_tree_add_7_25_groupi_n_1462 ,csa_tree_add_7_25_groupi_n_1461);
  not csa_tree_add_7_25_groupi_drc_bufs22276(csa_tree_add_7_25_groupi_n_1461 ,csa_tree_add_7_25_groupi_n_2844);
  not csa_tree_add_7_25_groupi_drc_bufs22278(csa_tree_add_7_25_groupi_n_1460 ,csa_tree_add_7_25_groupi_n_1458);
  not csa_tree_add_7_25_groupi_drc_bufs22279(csa_tree_add_7_25_groupi_n_1459 ,csa_tree_add_7_25_groupi_n_1458);
  not csa_tree_add_7_25_groupi_drc_bufs22280(csa_tree_add_7_25_groupi_n_1458 ,csa_tree_add_7_25_groupi_n_3502);
  not csa_tree_add_7_25_groupi_drc_bufs22282(csa_tree_add_7_25_groupi_n_1457 ,csa_tree_add_7_25_groupi_n_1455);
  not csa_tree_add_7_25_groupi_drc_bufs22283(csa_tree_add_7_25_groupi_n_1456 ,csa_tree_add_7_25_groupi_n_1455);
  not csa_tree_add_7_25_groupi_drc_bufs22284(csa_tree_add_7_25_groupi_n_1455 ,csa_tree_add_7_25_groupi_n_3500);
  not csa_tree_add_7_25_groupi_drc_bufs22286(csa_tree_add_7_25_groupi_n_1454 ,csa_tree_add_7_25_groupi_n_1452);
  not csa_tree_add_7_25_groupi_drc_bufs22287(csa_tree_add_7_25_groupi_n_1453 ,csa_tree_add_7_25_groupi_n_1452);
  not csa_tree_add_7_25_groupi_drc_bufs22288(csa_tree_add_7_25_groupi_n_1452 ,csa_tree_add_7_25_groupi_n_3499);
  not csa_tree_add_7_25_groupi_drc_bufs22290(csa_tree_add_7_25_groupi_n_1451 ,csa_tree_add_7_25_groupi_n_1449);
  not csa_tree_add_7_25_groupi_drc_bufs22291(csa_tree_add_7_25_groupi_n_1450 ,csa_tree_add_7_25_groupi_n_1449);
  not csa_tree_add_7_25_groupi_drc_bufs22292(csa_tree_add_7_25_groupi_n_1449 ,csa_tree_add_7_25_groupi_n_2863);
  not csa_tree_add_7_25_groupi_drc_bufs22294(csa_tree_add_7_25_groupi_n_1448 ,csa_tree_add_7_25_groupi_n_1446);
  not csa_tree_add_7_25_groupi_drc_bufs22295(csa_tree_add_7_25_groupi_n_1447 ,csa_tree_add_7_25_groupi_n_1446);
  not csa_tree_add_7_25_groupi_drc_bufs22296(csa_tree_add_7_25_groupi_n_1446 ,csa_tree_add_7_25_groupi_n_2861);
  not csa_tree_add_7_25_groupi_drc_bufs22298(csa_tree_add_7_25_groupi_n_1445 ,csa_tree_add_7_25_groupi_n_1443);
  not csa_tree_add_7_25_groupi_drc_bufs22299(csa_tree_add_7_25_groupi_n_1444 ,csa_tree_add_7_25_groupi_n_1443);
  not csa_tree_add_7_25_groupi_drc_bufs22300(csa_tree_add_7_25_groupi_n_1443 ,csa_tree_add_7_25_groupi_n_2861);
  not csa_tree_add_7_25_groupi_drc_bufs22302(csa_tree_add_7_25_groupi_n_1442 ,csa_tree_add_7_25_groupi_n_1440);
  not csa_tree_add_7_25_groupi_drc_bufs22303(csa_tree_add_7_25_groupi_n_1441 ,csa_tree_add_7_25_groupi_n_1440);
  not csa_tree_add_7_25_groupi_drc_bufs22304(csa_tree_add_7_25_groupi_n_1440 ,csa_tree_add_7_25_groupi_n_2854);
  not csa_tree_add_7_25_groupi_drc_bufs22306(csa_tree_add_7_25_groupi_n_1439 ,csa_tree_add_7_25_groupi_n_1437);
  not csa_tree_add_7_25_groupi_drc_bufs22307(csa_tree_add_7_25_groupi_n_1438 ,csa_tree_add_7_25_groupi_n_1437);
  not csa_tree_add_7_25_groupi_drc_bufs22308(csa_tree_add_7_25_groupi_n_1437 ,csa_tree_add_7_25_groupi_n_2854);
  not csa_tree_add_7_25_groupi_drc_bufs22310(csa_tree_add_7_25_groupi_n_1436 ,csa_tree_add_7_25_groupi_n_1434);
  not csa_tree_add_7_25_groupi_drc_bufs22311(csa_tree_add_7_25_groupi_n_1435 ,csa_tree_add_7_25_groupi_n_1434);
  not csa_tree_add_7_25_groupi_drc_bufs22312(csa_tree_add_7_25_groupi_n_1434 ,csa_tree_add_7_25_groupi_n_2858);
  not csa_tree_add_7_25_groupi_drc_bufs22314(csa_tree_add_7_25_groupi_n_1433 ,csa_tree_add_7_25_groupi_n_1431);
  not csa_tree_add_7_25_groupi_drc_bufs22315(csa_tree_add_7_25_groupi_n_1432 ,csa_tree_add_7_25_groupi_n_1431);
  not csa_tree_add_7_25_groupi_drc_bufs22316(csa_tree_add_7_25_groupi_n_1431 ,csa_tree_add_7_25_groupi_n_2856);
  not csa_tree_add_7_25_groupi_drc_bufs22318(csa_tree_add_7_25_groupi_n_1430 ,csa_tree_add_7_25_groupi_n_1428);
  not csa_tree_add_7_25_groupi_drc_bufs22319(csa_tree_add_7_25_groupi_n_1429 ,csa_tree_add_7_25_groupi_n_1428);
  not csa_tree_add_7_25_groupi_drc_bufs22320(csa_tree_add_7_25_groupi_n_1428 ,csa_tree_add_7_25_groupi_n_2522);
  not csa_tree_add_7_25_groupi_drc_bufs22322(csa_tree_add_7_25_groupi_n_1427 ,csa_tree_add_7_25_groupi_n_1425);
  not csa_tree_add_7_25_groupi_drc_bufs22323(csa_tree_add_7_25_groupi_n_1426 ,csa_tree_add_7_25_groupi_n_1425);
  not csa_tree_add_7_25_groupi_drc_bufs22324(csa_tree_add_7_25_groupi_n_1425 ,csa_tree_add_7_25_groupi_n_2858);
  not csa_tree_add_7_25_groupi_drc_bufs22326(csa_tree_add_7_25_groupi_n_1424 ,csa_tree_add_7_25_groupi_n_1422);
  not csa_tree_add_7_25_groupi_drc_bufs22327(csa_tree_add_7_25_groupi_n_1423 ,csa_tree_add_7_25_groupi_n_1422);
  not csa_tree_add_7_25_groupi_drc_bufs22328(csa_tree_add_7_25_groupi_n_1422 ,csa_tree_add_7_25_groupi_n_2853);
  not csa_tree_add_7_25_groupi_drc_bufs22330(csa_tree_add_7_25_groupi_n_1421 ,csa_tree_add_7_25_groupi_n_1419);
  not csa_tree_add_7_25_groupi_drc_bufs22331(csa_tree_add_7_25_groupi_n_1420 ,csa_tree_add_7_25_groupi_n_1419);
  not csa_tree_add_7_25_groupi_drc_bufs22332(csa_tree_add_7_25_groupi_n_1419 ,csa_tree_add_7_25_groupi_n_3503);
  not csa_tree_add_7_25_groupi_drc_bufs22334(csa_tree_add_7_25_groupi_n_1418 ,csa_tree_add_7_25_groupi_n_1416);
  not csa_tree_add_7_25_groupi_drc_bufs22335(csa_tree_add_7_25_groupi_n_1417 ,csa_tree_add_7_25_groupi_n_1416);
  not csa_tree_add_7_25_groupi_drc_bufs22336(csa_tree_add_7_25_groupi_n_1416 ,csa_tree_add_7_25_groupi_n_3513);
  not csa_tree_add_7_25_groupi_drc_bufs22338(csa_tree_add_7_25_groupi_n_1415 ,csa_tree_add_7_25_groupi_n_1413);
  not csa_tree_add_7_25_groupi_drc_bufs22339(csa_tree_add_7_25_groupi_n_1414 ,csa_tree_add_7_25_groupi_n_1413);
  not csa_tree_add_7_25_groupi_drc_bufs22340(csa_tree_add_7_25_groupi_n_1413 ,csa_tree_add_7_25_groupi_n_2848);
  not csa_tree_add_7_25_groupi_drc_bufs22342(csa_tree_add_7_25_groupi_n_1412 ,csa_tree_add_7_25_groupi_n_1410);
  not csa_tree_add_7_25_groupi_drc_bufs22343(csa_tree_add_7_25_groupi_n_1411 ,csa_tree_add_7_25_groupi_n_1410);
  not csa_tree_add_7_25_groupi_drc_bufs22344(csa_tree_add_7_25_groupi_n_1410 ,csa_tree_add_7_25_groupi_n_2768);
  not csa_tree_add_7_25_groupi_drc_bufs22346(csa_tree_add_7_25_groupi_n_1409 ,csa_tree_add_7_25_groupi_n_1407);
  not csa_tree_add_7_25_groupi_drc_bufs22347(csa_tree_add_7_25_groupi_n_1408 ,csa_tree_add_7_25_groupi_n_1407);
  not csa_tree_add_7_25_groupi_drc_bufs22348(csa_tree_add_7_25_groupi_n_1407 ,csa_tree_add_7_25_groupi_n_3519);
  not csa_tree_add_7_25_groupi_drc_bufs22350(csa_tree_add_7_25_groupi_n_1406 ,csa_tree_add_7_25_groupi_n_1404);
  not csa_tree_add_7_25_groupi_drc_bufs22351(csa_tree_add_7_25_groupi_n_1405 ,csa_tree_add_7_25_groupi_n_1404);
  not csa_tree_add_7_25_groupi_drc_bufs22352(csa_tree_add_7_25_groupi_n_1404 ,csa_tree_add_7_25_groupi_n_2763);
  not csa_tree_add_7_25_groupi_drc_bufs22354(csa_tree_add_7_25_groupi_n_1403 ,csa_tree_add_7_25_groupi_n_1401);
  not csa_tree_add_7_25_groupi_drc_bufs22355(csa_tree_add_7_25_groupi_n_1402 ,csa_tree_add_7_25_groupi_n_1401);
  not csa_tree_add_7_25_groupi_drc_bufs22356(csa_tree_add_7_25_groupi_n_1401 ,csa_tree_add_7_25_groupi_n_2758);
  not csa_tree_add_7_25_groupi_drc_bufs22358(csa_tree_add_7_25_groupi_n_1400 ,csa_tree_add_7_25_groupi_n_1398);
  not csa_tree_add_7_25_groupi_drc_bufs22359(csa_tree_add_7_25_groupi_n_1399 ,csa_tree_add_7_25_groupi_n_1398);
  not csa_tree_add_7_25_groupi_drc_bufs22360(csa_tree_add_7_25_groupi_n_1398 ,csa_tree_add_7_25_groupi_n_2759);
  not csa_tree_add_7_25_groupi_drc_bufs22362(csa_tree_add_7_25_groupi_n_1397 ,csa_tree_add_7_25_groupi_n_1395);
  not csa_tree_add_7_25_groupi_drc_bufs22363(csa_tree_add_7_25_groupi_n_1396 ,csa_tree_add_7_25_groupi_n_1395);
  not csa_tree_add_7_25_groupi_drc_bufs22364(csa_tree_add_7_25_groupi_n_1395 ,csa_tree_add_7_25_groupi_n_2754);
  not csa_tree_add_7_25_groupi_drc_bufs22366(csa_tree_add_7_25_groupi_n_1394 ,csa_tree_add_7_25_groupi_n_1392);
  not csa_tree_add_7_25_groupi_drc_bufs22367(csa_tree_add_7_25_groupi_n_1393 ,csa_tree_add_7_25_groupi_n_1392);
  not csa_tree_add_7_25_groupi_drc_bufs22368(csa_tree_add_7_25_groupi_n_1392 ,csa_tree_add_7_25_groupi_n_2841);
  not csa_tree_add_7_25_groupi_drc_bufs22370(csa_tree_add_7_25_groupi_n_1391 ,csa_tree_add_7_25_groupi_n_1389);
  not csa_tree_add_7_25_groupi_drc_bufs22371(csa_tree_add_7_25_groupi_n_1390 ,csa_tree_add_7_25_groupi_n_1389);
  not csa_tree_add_7_25_groupi_drc_bufs22372(csa_tree_add_7_25_groupi_n_1389 ,csa_tree_add_7_25_groupi_n_2760);
  not csa_tree_add_7_25_groupi_drc_bufs22374(csa_tree_add_7_25_groupi_n_1388 ,csa_tree_add_7_25_groupi_n_1386);
  not csa_tree_add_7_25_groupi_drc_bufs22375(csa_tree_add_7_25_groupi_n_1387 ,csa_tree_add_7_25_groupi_n_1386);
  not csa_tree_add_7_25_groupi_drc_bufs22376(csa_tree_add_7_25_groupi_n_1386 ,csa_tree_add_7_25_groupi_n_3508);
  not csa_tree_add_7_25_groupi_drc_bufs22378(csa_tree_add_7_25_groupi_n_1385 ,csa_tree_add_7_25_groupi_n_1383);
  not csa_tree_add_7_25_groupi_drc_bufs22379(csa_tree_add_7_25_groupi_n_1384 ,csa_tree_add_7_25_groupi_n_1383);
  not csa_tree_add_7_25_groupi_drc_bufs22380(csa_tree_add_7_25_groupi_n_1383 ,csa_tree_add_7_25_groupi_n_3504);
  not csa_tree_add_7_25_groupi_drc_bufs22382(csa_tree_add_7_25_groupi_n_1382 ,csa_tree_add_7_25_groupi_n_1380);
  not csa_tree_add_7_25_groupi_drc_bufs22383(csa_tree_add_7_25_groupi_n_1381 ,csa_tree_add_7_25_groupi_n_1380);
  not csa_tree_add_7_25_groupi_drc_bufs22384(csa_tree_add_7_25_groupi_n_1380 ,csa_tree_add_7_25_groupi_n_3510);
  not csa_tree_add_7_25_groupi_drc_bufs22386(csa_tree_add_7_25_groupi_n_1379 ,csa_tree_add_7_25_groupi_n_1377);
  not csa_tree_add_7_25_groupi_drc_bufs22387(csa_tree_add_7_25_groupi_n_1378 ,csa_tree_add_7_25_groupi_n_1377);
  not csa_tree_add_7_25_groupi_drc_bufs22388(csa_tree_add_7_25_groupi_n_1377 ,csa_tree_add_7_25_groupi_n_3507);
  not csa_tree_add_7_25_groupi_drc_bufs22390(csa_tree_add_7_25_groupi_n_1376 ,csa_tree_add_7_25_groupi_n_1374);
  not csa_tree_add_7_25_groupi_drc_bufs22391(csa_tree_add_7_25_groupi_n_1375 ,csa_tree_add_7_25_groupi_n_1374);
  not csa_tree_add_7_25_groupi_drc_bufs22392(csa_tree_add_7_25_groupi_n_1374 ,csa_tree_add_7_25_groupi_n_2845);
  not csa_tree_add_7_25_groupi_drc_bufs22394(csa_tree_add_7_25_groupi_n_1373 ,csa_tree_add_7_25_groupi_n_1371);
  not csa_tree_add_7_25_groupi_drc_bufs22395(csa_tree_add_7_25_groupi_n_1372 ,csa_tree_add_7_25_groupi_n_1371);
  not csa_tree_add_7_25_groupi_drc_bufs22396(csa_tree_add_7_25_groupi_n_1371 ,csa_tree_add_7_25_groupi_n_2773);
  not csa_tree_add_7_25_groupi_drc_bufs22398(csa_tree_add_7_25_groupi_n_1370 ,csa_tree_add_7_25_groupi_n_1368);
  not csa_tree_add_7_25_groupi_drc_bufs22399(csa_tree_add_7_25_groupi_n_1369 ,csa_tree_add_7_25_groupi_n_1368);
  not csa_tree_add_7_25_groupi_drc_bufs22400(csa_tree_add_7_25_groupi_n_1368 ,csa_tree_add_7_25_groupi_n_2845);
  not csa_tree_add_7_25_groupi_drc_bufs22402(csa_tree_add_7_25_groupi_n_1367 ,csa_tree_add_7_25_groupi_n_1365);
  not csa_tree_add_7_25_groupi_drc_bufs22403(csa_tree_add_7_25_groupi_n_1366 ,csa_tree_add_7_25_groupi_n_1365);
  not csa_tree_add_7_25_groupi_drc_bufs22404(csa_tree_add_7_25_groupi_n_1365 ,csa_tree_add_7_25_groupi_n_2849);
  not csa_tree_add_7_25_groupi_drc_bufs22406(csa_tree_add_7_25_groupi_n_1364 ,csa_tree_add_7_25_groupi_n_1362);
  not csa_tree_add_7_25_groupi_drc_bufs22407(csa_tree_add_7_25_groupi_n_1363 ,csa_tree_add_7_25_groupi_n_1362);
  not csa_tree_add_7_25_groupi_drc_bufs22408(csa_tree_add_7_25_groupi_n_1362 ,csa_tree_add_7_25_groupi_n_2770);
  not csa_tree_add_7_25_groupi_drc_bufs22410(csa_tree_add_7_25_groupi_n_1361 ,csa_tree_add_7_25_groupi_n_1359);
  not csa_tree_add_7_25_groupi_drc_bufs22411(csa_tree_add_7_25_groupi_n_1360 ,csa_tree_add_7_25_groupi_n_1359);
  not csa_tree_add_7_25_groupi_drc_bufs22412(csa_tree_add_7_25_groupi_n_1359 ,csa_tree_add_7_25_groupi_n_2755);
  not csa_tree_add_7_25_groupi_drc_bufs22414(csa_tree_add_7_25_groupi_n_1358 ,csa_tree_add_7_25_groupi_n_1356);
  not csa_tree_add_7_25_groupi_drc_bufs22415(csa_tree_add_7_25_groupi_n_1357 ,csa_tree_add_7_25_groupi_n_1356);
  not csa_tree_add_7_25_groupi_drc_bufs22416(csa_tree_add_7_25_groupi_n_1356 ,csa_tree_add_7_25_groupi_n_2767);
  not csa_tree_add_7_25_groupi_drc_bufs22418(csa_tree_add_7_25_groupi_n_1355 ,csa_tree_add_7_25_groupi_n_1353);
  not csa_tree_add_7_25_groupi_drc_bufs22419(csa_tree_add_7_25_groupi_n_1354 ,csa_tree_add_7_25_groupi_n_1353);
  not csa_tree_add_7_25_groupi_drc_bufs22420(csa_tree_add_7_25_groupi_n_1353 ,csa_tree_add_7_25_groupi_n_2848);
  not csa_tree_add_7_25_groupi_drc_bufs22422(csa_tree_add_7_25_groupi_n_1352 ,csa_tree_add_7_25_groupi_n_1350);
  not csa_tree_add_7_25_groupi_drc_bufs22423(csa_tree_add_7_25_groupi_n_1351 ,csa_tree_add_7_25_groupi_n_1350);
  not csa_tree_add_7_25_groupi_drc_bufs22424(csa_tree_add_7_25_groupi_n_1350 ,csa_tree_add_7_25_groupi_n_2774);
  not csa_tree_add_7_25_groupi_drc_bufs22426(csa_tree_add_7_25_groupi_n_1349 ,csa_tree_add_7_25_groupi_n_1347);
  not csa_tree_add_7_25_groupi_drc_bufs22427(csa_tree_add_7_25_groupi_n_1348 ,csa_tree_add_7_25_groupi_n_1347);
  not csa_tree_add_7_25_groupi_drc_bufs22428(csa_tree_add_7_25_groupi_n_1347 ,csa_tree_add_7_25_groupi_n_2863);
  not csa_tree_add_7_25_groupi_drc_bufs22430(csa_tree_add_7_25_groupi_n_1346 ,csa_tree_add_7_25_groupi_n_1344);
  not csa_tree_add_7_25_groupi_drc_bufs22431(csa_tree_add_7_25_groupi_n_1345 ,csa_tree_add_7_25_groupi_n_1344);
  not csa_tree_add_7_25_groupi_drc_bufs22432(csa_tree_add_7_25_groupi_n_1344 ,csa_tree_add_7_25_groupi_n_2865);
  not csa_tree_add_7_25_groupi_drc_bufs22434(csa_tree_add_7_25_groupi_n_1343 ,csa_tree_add_7_25_groupi_n_1341);
  not csa_tree_add_7_25_groupi_drc_bufs22435(csa_tree_add_7_25_groupi_n_1342 ,csa_tree_add_7_25_groupi_n_1341);
  not csa_tree_add_7_25_groupi_drc_bufs22436(csa_tree_add_7_25_groupi_n_1341 ,csa_tree_add_7_25_groupi_n_3519);
  not csa_tree_add_7_25_groupi_drc_bufs22438(csa_tree_add_7_25_groupi_n_1340 ,csa_tree_add_7_25_groupi_n_1338);
  not csa_tree_add_7_25_groupi_drc_bufs22439(csa_tree_add_7_25_groupi_n_1339 ,csa_tree_add_7_25_groupi_n_1338);
  not csa_tree_add_7_25_groupi_drc_bufs22440(csa_tree_add_7_25_groupi_n_1338 ,csa_tree_add_7_25_groupi_n_2851);
  not csa_tree_add_7_25_groupi_drc_bufs22442(csa_tree_add_7_25_groupi_n_1337 ,csa_tree_add_7_25_groupi_n_1335);
  not csa_tree_add_7_25_groupi_drc_bufs22443(csa_tree_add_7_25_groupi_n_1336 ,csa_tree_add_7_25_groupi_n_1335);
  not csa_tree_add_7_25_groupi_drc_bufs22444(csa_tree_add_7_25_groupi_n_1335 ,csa_tree_add_7_25_groupi_n_2785);
  not csa_tree_add_7_25_groupi_drc_bufs22446(csa_tree_add_7_25_groupi_n_1334 ,csa_tree_add_7_25_groupi_n_1332);
  not csa_tree_add_7_25_groupi_drc_bufs22447(csa_tree_add_7_25_groupi_n_1333 ,csa_tree_add_7_25_groupi_n_1332);
  not csa_tree_add_7_25_groupi_drc_bufs22448(csa_tree_add_7_25_groupi_n_1332 ,csa_tree_add_7_25_groupi_n_2850);
  not csa_tree_add_7_25_groupi_drc_bufs22450(csa_tree_add_7_25_groupi_n_1331 ,csa_tree_add_7_25_groupi_n_1329);
  not csa_tree_add_7_25_groupi_drc_bufs22451(csa_tree_add_7_25_groupi_n_1330 ,csa_tree_add_7_25_groupi_n_1329);
  not csa_tree_add_7_25_groupi_drc_bufs22452(csa_tree_add_7_25_groupi_n_1329 ,csa_tree_add_7_25_groupi_n_2785);
  not csa_tree_add_7_25_groupi_drc_bufs22454(csa_tree_add_7_25_groupi_n_1328 ,csa_tree_add_7_25_groupi_n_1326);
  not csa_tree_add_7_25_groupi_drc_bufs22455(csa_tree_add_7_25_groupi_n_1327 ,csa_tree_add_7_25_groupi_n_1326);
  not csa_tree_add_7_25_groupi_drc_bufs22456(csa_tree_add_7_25_groupi_n_1326 ,csa_tree_add_7_25_groupi_n_2853);
  not csa_tree_add_7_25_groupi_drc_bufs22458(csa_tree_add_7_25_groupi_n_1325 ,csa_tree_add_7_25_groupi_n_1323);
  not csa_tree_add_7_25_groupi_drc_bufs22459(csa_tree_add_7_25_groupi_n_1324 ,csa_tree_add_7_25_groupi_n_1323);
  not csa_tree_add_7_25_groupi_drc_bufs22460(csa_tree_add_7_25_groupi_n_1323 ,csa_tree_add_7_25_groupi_n_2777);
  not csa_tree_add_7_25_groupi_drc_bufs22462(csa_tree_add_7_25_groupi_n_1322 ,csa_tree_add_7_25_groupi_n_1320);
  not csa_tree_add_7_25_groupi_drc_bufs22463(csa_tree_add_7_25_groupi_n_1321 ,csa_tree_add_7_25_groupi_n_1320);
  not csa_tree_add_7_25_groupi_drc_bufs22464(csa_tree_add_7_25_groupi_n_1320 ,csa_tree_add_7_25_groupi_n_2886);
  not csa_tree_add_7_25_groupi_drc_bufs22466(csa_tree_add_7_25_groupi_n_1319 ,csa_tree_add_7_25_groupi_n_1317);
  not csa_tree_add_7_25_groupi_drc_bufs22467(csa_tree_add_7_25_groupi_n_1318 ,csa_tree_add_7_25_groupi_n_1317);
  not csa_tree_add_7_25_groupi_drc_bufs22468(csa_tree_add_7_25_groupi_n_1317 ,csa_tree_add_7_25_groupi_n_2886);
  not csa_tree_add_7_25_groupi_drc_bufs22470(csa_tree_add_7_25_groupi_n_1316 ,csa_tree_add_7_25_groupi_n_1314);
  not csa_tree_add_7_25_groupi_drc_bufs22471(csa_tree_add_7_25_groupi_n_1315 ,csa_tree_add_7_25_groupi_n_1314);
  not csa_tree_add_7_25_groupi_drc_bufs22472(csa_tree_add_7_25_groupi_n_1314 ,csa_tree_add_7_25_groupi_n_2883);
  not csa_tree_add_7_25_groupi_drc_bufs22474(csa_tree_add_7_25_groupi_n_1313 ,csa_tree_add_7_25_groupi_n_1311);
  not csa_tree_add_7_25_groupi_drc_bufs22475(csa_tree_add_7_25_groupi_n_1312 ,csa_tree_add_7_25_groupi_n_1311);
  not csa_tree_add_7_25_groupi_drc_bufs22476(csa_tree_add_7_25_groupi_n_1311 ,csa_tree_add_7_25_groupi_n_2799);
  not csa_tree_add_7_25_groupi_drc_bufs22478(csa_tree_add_7_25_groupi_n_1310 ,csa_tree_add_7_25_groupi_n_1308);
  not csa_tree_add_7_25_groupi_drc_bufs22479(csa_tree_add_7_25_groupi_n_1309 ,csa_tree_add_7_25_groupi_n_1308);
  not csa_tree_add_7_25_groupi_drc_bufs22480(csa_tree_add_7_25_groupi_n_1308 ,csa_tree_add_7_25_groupi_n_2802);
  not csa_tree_add_7_25_groupi_drc_bufs22482(csa_tree_add_7_25_groupi_n_1307 ,csa_tree_add_7_25_groupi_n_1305);
  not csa_tree_add_7_25_groupi_drc_bufs22483(csa_tree_add_7_25_groupi_n_1306 ,csa_tree_add_7_25_groupi_n_1305);
  not csa_tree_add_7_25_groupi_drc_bufs22484(csa_tree_add_7_25_groupi_n_1305 ,csa_tree_add_7_25_groupi_n_2883);
  not csa_tree_add_7_25_groupi_drc_bufs22486(csa_tree_add_7_25_groupi_n_1304 ,csa_tree_add_7_25_groupi_n_1302);
  not csa_tree_add_7_25_groupi_drc_bufs22487(csa_tree_add_7_25_groupi_n_1303 ,csa_tree_add_7_25_groupi_n_1302);
  not csa_tree_add_7_25_groupi_drc_bufs22488(csa_tree_add_7_25_groupi_n_1302 ,csa_tree_add_7_25_groupi_n_2799);
  not csa_tree_add_7_25_groupi_drc_bufs22490(csa_tree_add_7_25_groupi_n_1301 ,csa_tree_add_7_25_groupi_n_1299);
  not csa_tree_add_7_25_groupi_drc_bufs22491(csa_tree_add_7_25_groupi_n_1300 ,csa_tree_add_7_25_groupi_n_1299);
  not csa_tree_add_7_25_groupi_drc_bufs22492(csa_tree_add_7_25_groupi_n_1299 ,csa_tree_add_7_25_groupi_n_3534);
  not csa_tree_add_7_25_groupi_drc_bufs22494(csa_tree_add_7_25_groupi_n_1298 ,csa_tree_add_7_25_groupi_n_1296);
  not csa_tree_add_7_25_groupi_drc_bufs22495(csa_tree_add_7_25_groupi_n_1297 ,csa_tree_add_7_25_groupi_n_1296);
  not csa_tree_add_7_25_groupi_drc_bufs22496(csa_tree_add_7_25_groupi_n_1296 ,csa_tree_add_7_25_groupi_n_2880);
  not csa_tree_add_7_25_groupi_drc_bufs22498(csa_tree_add_7_25_groupi_n_1295 ,csa_tree_add_7_25_groupi_n_1293);
  not csa_tree_add_7_25_groupi_drc_bufs22499(csa_tree_add_7_25_groupi_n_1294 ,csa_tree_add_7_25_groupi_n_1293);
  not csa_tree_add_7_25_groupi_drc_bufs22500(csa_tree_add_7_25_groupi_n_1293 ,csa_tree_add_7_25_groupi_n_3534);
  not csa_tree_add_7_25_groupi_drc_bufs22502(csa_tree_add_7_25_groupi_n_1292 ,csa_tree_add_7_25_groupi_n_1290);
  not csa_tree_add_7_25_groupi_drc_bufs22503(csa_tree_add_7_25_groupi_n_1291 ,csa_tree_add_7_25_groupi_n_1290);
  not csa_tree_add_7_25_groupi_drc_bufs22504(csa_tree_add_7_25_groupi_n_1290 ,csa_tree_add_7_25_groupi_n_2880);
  not csa_tree_add_7_25_groupi_drc_bufs22506(csa_tree_add_7_25_groupi_n_1289 ,csa_tree_add_7_25_groupi_n_1287);
  not csa_tree_add_7_25_groupi_drc_bufs22507(csa_tree_add_7_25_groupi_n_1288 ,csa_tree_add_7_25_groupi_n_1287);
  not csa_tree_add_7_25_groupi_drc_bufs22508(csa_tree_add_7_25_groupi_n_1287 ,csa_tree_add_7_25_groupi_n_6463);
  not csa_tree_add_7_25_groupi_drc_bufs22510(csa_tree_add_7_25_groupi_n_1286 ,csa_tree_add_7_25_groupi_n_1284);
  not csa_tree_add_7_25_groupi_drc_bufs22511(csa_tree_add_7_25_groupi_n_1285 ,csa_tree_add_7_25_groupi_n_1284);
  not csa_tree_add_7_25_groupi_drc_bufs22512(csa_tree_add_7_25_groupi_n_1284 ,csa_tree_add_7_25_groupi_n_5763);
  not csa_tree_add_7_25_groupi_drc_bufs22514(csa_tree_add_7_25_groupi_n_1283 ,csa_tree_add_7_25_groupi_n_1281);
  not csa_tree_add_7_25_groupi_drc_bufs22515(csa_tree_add_7_25_groupi_n_1282 ,csa_tree_add_7_25_groupi_n_1281);
  not csa_tree_add_7_25_groupi_drc_bufs22516(csa_tree_add_7_25_groupi_n_1281 ,csa_tree_add_7_25_groupi_n_6178);
  not csa_tree_add_7_25_groupi_drc_bufs22518(csa_tree_add_7_25_groupi_n_1280 ,csa_tree_add_7_25_groupi_n_1278);
  not csa_tree_add_7_25_groupi_drc_bufs22519(csa_tree_add_7_25_groupi_n_1279 ,csa_tree_add_7_25_groupi_n_1278);
  not csa_tree_add_7_25_groupi_drc_bufs22520(csa_tree_add_7_25_groupi_n_1278 ,csa_tree_add_7_25_groupi_n_6087);
  not csa_tree_add_7_25_groupi_drc_bufs22522(csa_tree_add_7_25_groupi_n_1277 ,csa_tree_add_7_25_groupi_n_1275);
  not csa_tree_add_7_25_groupi_drc_bufs22523(csa_tree_add_7_25_groupi_n_1276 ,csa_tree_add_7_25_groupi_n_1275);
  not csa_tree_add_7_25_groupi_drc_bufs22524(csa_tree_add_7_25_groupi_n_1275 ,csa_tree_add_7_25_groupi_n_6284);
  not csa_tree_add_7_25_groupi_drc_bufs22526(csa_tree_add_7_25_groupi_n_1274 ,csa_tree_add_7_25_groupi_n_1272);
  not csa_tree_add_7_25_groupi_drc_bufs22527(csa_tree_add_7_25_groupi_n_1273 ,csa_tree_add_7_25_groupi_n_1272);
  not csa_tree_add_7_25_groupi_drc_bufs22528(csa_tree_add_7_25_groupi_n_1272 ,csa_tree_add_7_25_groupi_n_6087);
  not csa_tree_add_7_25_groupi_drc_bufs22530(csa_tree_add_7_25_groupi_n_1271 ,csa_tree_add_7_25_groupi_n_1269);
  not csa_tree_add_7_25_groupi_drc_bufs22531(csa_tree_add_7_25_groupi_n_1270 ,csa_tree_add_7_25_groupi_n_1269);
  not csa_tree_add_7_25_groupi_drc_bufs22532(csa_tree_add_7_25_groupi_n_1269 ,csa_tree_add_7_25_groupi_n_6178);
  not csa_tree_add_7_25_groupi_drc_bufs22534(csa_tree_add_7_25_groupi_n_1268 ,csa_tree_add_7_25_groupi_n_1266);
  not csa_tree_add_7_25_groupi_drc_bufs22535(csa_tree_add_7_25_groupi_n_1267 ,csa_tree_add_7_25_groupi_n_1266);
  not csa_tree_add_7_25_groupi_drc_bufs22536(csa_tree_add_7_25_groupi_n_1266 ,csa_tree_add_7_25_groupi_n_6284);
  not csa_tree_add_7_25_groupi_drc_bufs22538(csa_tree_add_7_25_groupi_n_1265 ,csa_tree_add_7_25_groupi_n_1263);
  not csa_tree_add_7_25_groupi_drc_bufs22539(csa_tree_add_7_25_groupi_n_1264 ,csa_tree_add_7_25_groupi_n_1263);
  not csa_tree_add_7_25_groupi_drc_bufs22540(csa_tree_add_7_25_groupi_n_1263 ,csa_tree_add_7_25_groupi_n_6382);
  not csa_tree_add_7_25_groupi_drc_bufs22542(csa_tree_add_7_25_groupi_n_1262 ,csa_tree_add_7_25_groupi_n_1260);
  not csa_tree_add_7_25_groupi_drc_bufs22543(csa_tree_add_7_25_groupi_n_1261 ,csa_tree_add_7_25_groupi_n_1260);
  not csa_tree_add_7_25_groupi_drc_bufs22544(csa_tree_add_7_25_groupi_n_1260 ,csa_tree_add_7_25_groupi_n_5979);
  not csa_tree_add_7_25_groupi_drc_bufs22546(csa_tree_add_7_25_groupi_n_1259 ,csa_tree_add_7_25_groupi_n_1257);
  not csa_tree_add_7_25_groupi_drc_bufs22547(csa_tree_add_7_25_groupi_n_1258 ,csa_tree_add_7_25_groupi_n_1257);
  not csa_tree_add_7_25_groupi_drc_bufs22548(csa_tree_add_7_25_groupi_n_1257 ,csa_tree_add_7_25_groupi_n_6560);
  not csa_tree_add_7_25_groupi_drc_bufs22550(csa_tree_add_7_25_groupi_n_1256 ,csa_tree_add_7_25_groupi_n_1254);
  not csa_tree_add_7_25_groupi_drc_bufs22551(csa_tree_add_7_25_groupi_n_1255 ,csa_tree_add_7_25_groupi_n_1254);
  not csa_tree_add_7_25_groupi_drc_bufs22552(csa_tree_add_7_25_groupi_n_1254 ,csa_tree_add_7_25_groupi_n_5864);
  not csa_tree_add_7_25_groupi_drc_bufs22554(csa_tree_add_7_25_groupi_n_1253 ,csa_tree_add_7_25_groupi_n_1803);
  not csa_tree_add_7_25_groupi_drc_bufs22558(csa_tree_add_7_25_groupi_n_1252 ,csa_tree_add_7_25_groupi_n_1802);
  not csa_tree_add_7_25_groupi_drc_bufs22562(csa_tree_add_7_25_groupi_n_1251 ,csa_tree_add_7_25_groupi_n_1250);
  not csa_tree_add_7_25_groupi_drc_bufs22564(csa_tree_add_7_25_groupi_n_1250 ,csa_tree_add_7_25_groupi_n_2780);
  not csa_tree_add_7_25_groupi_drc_bufs22566(csa_tree_add_7_25_groupi_n_1249 ,csa_tree_add_7_25_groupi_n_1250);
  not csa_tree_add_7_25_groupi_drc_bufs22574(csa_tree_add_7_25_groupi_n_1248 ,csa_tree_add_7_25_groupi_n_1804);
  not csa_tree_add_7_25_groupi_drc_bufs22578(csa_tree_add_7_25_groupi_n_1247 ,csa_tree_add_7_25_groupi_n_1801);
  not csa_tree_add_7_25_groupi_drc_bufs22582(csa_tree_add_7_25_groupi_n_1246 ,csa_tree_add_7_25_groupi_n_1800);
  not csa_tree_add_7_25_groupi_drc_bufs22586(csa_tree_add_7_25_groupi_n_1245 ,csa_tree_add_7_25_groupi_n_1243);
  not csa_tree_add_7_25_groupi_drc_bufs22587(csa_tree_add_7_25_groupi_n_1244 ,csa_tree_add_7_25_groupi_n_1243);
  not csa_tree_add_7_25_groupi_drc_bufs22588(csa_tree_add_7_25_groupi_n_1243 ,csa_tree_add_7_25_groupi_n_2773);
  not csa_tree_add_7_25_groupi_drc_bufs22590(csa_tree_add_7_25_groupi_n_1242 ,csa_tree_add_7_25_groupi_n_1240);
  not csa_tree_add_7_25_groupi_drc_bufs22591(csa_tree_add_7_25_groupi_n_1241 ,csa_tree_add_7_25_groupi_n_1240);
  not csa_tree_add_7_25_groupi_drc_bufs22592(csa_tree_add_7_25_groupi_n_1240 ,csa_tree_add_7_25_groupi_n_2758);
  not csa_tree_add_7_25_groupi_drc_bufs22594(csa_tree_add_7_25_groupi_n_1239 ,csa_tree_add_7_25_groupi_n_1237);
  not csa_tree_add_7_25_groupi_drc_bufs22595(csa_tree_add_7_25_groupi_n_1238 ,csa_tree_add_7_25_groupi_n_1237);
  not csa_tree_add_7_25_groupi_drc_bufs22596(csa_tree_add_7_25_groupi_n_1237 ,csa_tree_add_7_25_groupi_n_2778);
  not csa_tree_add_7_25_groupi_drc_bufs22598(csa_tree_add_7_25_groupi_n_1236 ,csa_tree_add_7_25_groupi_n_1234);
  not csa_tree_add_7_25_groupi_drc_bufs22599(csa_tree_add_7_25_groupi_n_1235 ,csa_tree_add_7_25_groupi_n_1234);
  not csa_tree_add_7_25_groupi_drc_bufs22600(csa_tree_add_7_25_groupi_n_1234 ,csa_tree_add_7_25_groupi_n_2768);
  not csa_tree_add_7_25_groupi_drc_bufs22602(csa_tree_add_7_25_groupi_n_1233 ,csa_tree_add_7_25_groupi_n_1231);
  not csa_tree_add_7_25_groupi_drc_bufs22603(csa_tree_add_7_25_groupi_n_1232 ,csa_tree_add_7_25_groupi_n_1231);
  not csa_tree_add_7_25_groupi_drc_bufs22604(csa_tree_add_7_25_groupi_n_1231 ,csa_tree_add_7_25_groupi_n_2844);
  not csa_tree_add_7_25_groupi_drc_bufs22606(csa_tree_add_7_25_groupi_n_1230 ,csa_tree_add_7_25_groupi_n_1228);
  not csa_tree_add_7_25_groupi_drc_bufs22607(csa_tree_add_7_25_groupi_n_1229 ,csa_tree_add_7_25_groupi_n_1228);
  not csa_tree_add_7_25_groupi_drc_bufs22608(csa_tree_add_7_25_groupi_n_1228 ,csa_tree_add_7_25_groupi_n_2763);
  not csa_tree_add_7_25_groupi_drc_bufs22610(csa_tree_add_7_25_groupi_n_1227 ,csa_tree_add_7_25_groupi_n_1225);
  not csa_tree_add_7_25_groupi_drc_bufs22611(csa_tree_add_7_25_groupi_n_1226 ,csa_tree_add_7_25_groupi_n_1225);
  not csa_tree_add_7_25_groupi_drc_bufs22612(csa_tree_add_7_25_groupi_n_1225 ,csa_tree_add_7_25_groupi_n_2383);
  not csa_tree_add_7_25_groupi_drc_bufs22614(csa_tree_add_7_25_groupi_n_1224 ,csa_tree_add_7_25_groupi_n_2362);
  not csa_tree_add_7_25_groupi_drc_bufs22615(csa_tree_add_7_25_groupi_n_1223 ,csa_tree_add_7_25_groupi_n_2362);
  not csa_tree_add_7_25_groupi_drc_bufs22618(csa_tree_add_7_25_groupi_n_1222 ,csa_tree_add_7_25_groupi_n_2394);
  not csa_tree_add_7_25_groupi_drc_bufs22619(csa_tree_add_7_25_groupi_n_1221 ,csa_tree_add_7_25_groupi_n_2394);
  not csa_tree_add_7_25_groupi_drc_bufs22622(csa_tree_add_7_25_groupi_n_1220 ,csa_tree_add_7_25_groupi_n_2392);
  not csa_tree_add_7_25_groupi_drc_bufs22623(csa_tree_add_7_25_groupi_n_1219 ,csa_tree_add_7_25_groupi_n_2392);
  not csa_tree_add_7_25_groupi_drc_bufs22626(csa_tree_add_7_25_groupi_n_1218 ,csa_tree_add_7_25_groupi_n_2359);
  not csa_tree_add_7_25_groupi_drc_bufs22627(csa_tree_add_7_25_groupi_n_1217 ,csa_tree_add_7_25_groupi_n_2359);
  not csa_tree_add_7_25_groupi_drc_bufs22630(csa_tree_add_7_25_groupi_n_1216 ,csa_tree_add_7_25_groupi_n_2360);
  not csa_tree_add_7_25_groupi_drc_bufs22631(csa_tree_add_7_25_groupi_n_1215 ,csa_tree_add_7_25_groupi_n_2360);
  not csa_tree_add_7_25_groupi_drc_bufs22634(csa_tree_add_7_25_groupi_n_1214 ,csa_tree_add_7_25_groupi_n_2386);
  not csa_tree_add_7_25_groupi_drc_bufs22635(csa_tree_add_7_25_groupi_n_1213 ,csa_tree_add_7_25_groupi_n_2386);
  not csa_tree_add_7_25_groupi_drc_bufs22638(csa_tree_add_7_25_groupi_n_1212 ,csa_tree_add_7_25_groupi_n_2396);
  not csa_tree_add_7_25_groupi_drc_bufs22639(csa_tree_add_7_25_groupi_n_1211 ,csa_tree_add_7_25_groupi_n_2396);
  not csa_tree_add_7_25_groupi_drc_bufs22642(csa_tree_add_7_25_groupi_n_1210 ,csa_tree_add_7_25_groupi_n_2395);
  not csa_tree_add_7_25_groupi_drc_bufs22643(csa_tree_add_7_25_groupi_n_1209 ,csa_tree_add_7_25_groupi_n_2395);
  not csa_tree_add_7_25_groupi_drc_bufs22646(csa_tree_add_7_25_groupi_n_1208 ,csa_tree_add_7_25_groupi_n_2357);
  not csa_tree_add_7_25_groupi_drc_bufs22647(csa_tree_add_7_25_groupi_n_1207 ,csa_tree_add_7_25_groupi_n_2357);
  not csa_tree_add_7_25_groupi_drc_bufs22650(csa_tree_add_7_25_groupi_n_1206 ,csa_tree_add_7_25_groupi_n_2361);
  not csa_tree_add_7_25_groupi_drc_bufs22651(csa_tree_add_7_25_groupi_n_1205 ,csa_tree_add_7_25_groupi_n_2361);
  not csa_tree_add_7_25_groupi_drc_bufs22654(csa_tree_add_7_25_groupi_n_1204 ,csa_tree_add_7_25_groupi_n_2388);
  not csa_tree_add_7_25_groupi_drc_bufs22655(csa_tree_add_7_25_groupi_n_1203 ,csa_tree_add_7_25_groupi_n_2388);
  not csa_tree_add_7_25_groupi_drc_bufs22658(csa_tree_add_7_25_groupi_n_1202 ,csa_tree_add_7_25_groupi_n_2390);
  not csa_tree_add_7_25_groupi_drc_bufs22659(csa_tree_add_7_25_groupi_n_1201 ,csa_tree_add_7_25_groupi_n_2390);
  not csa_tree_add_7_25_groupi_drc_bufs22662(csa_tree_add_7_25_groupi_n_1200 ,csa_tree_add_7_25_groupi_n_2355);
  not csa_tree_add_7_25_groupi_drc_bufs22663(csa_tree_add_7_25_groupi_n_1199 ,csa_tree_add_7_25_groupi_n_2355);
  not csa_tree_add_7_25_groupi_drc_bufs22666(csa_tree_add_7_25_groupi_n_1198 ,csa_tree_add_7_25_groupi_n_2400);
  not csa_tree_add_7_25_groupi_drc_bufs22667(csa_tree_add_7_25_groupi_n_1197 ,csa_tree_add_7_25_groupi_n_2400);
  not csa_tree_add_7_25_groupi_drc_bufs22670(csa_tree_add_7_25_groupi_n_1196 ,csa_tree_add_7_25_groupi_n_2387);
  not csa_tree_add_7_25_groupi_drc_bufs22671(csa_tree_add_7_25_groupi_n_1195 ,csa_tree_add_7_25_groupi_n_2387);
  not csa_tree_add_7_25_groupi_drc_bufs22674(csa_tree_add_7_25_groupi_n_1194 ,csa_tree_add_7_25_groupi_n_2402);
  not csa_tree_add_7_25_groupi_drc_bufs22675(csa_tree_add_7_25_groupi_n_1193 ,csa_tree_add_7_25_groupi_n_2402);
  not csa_tree_add_7_25_groupi_drc_bufs22678(csa_tree_add_7_25_groupi_n_1192 ,csa_tree_add_7_25_groupi_n_2358);
  not csa_tree_add_7_25_groupi_drc_bufs22679(csa_tree_add_7_25_groupi_n_1191 ,csa_tree_add_7_25_groupi_n_2358);
  not csa_tree_add_7_25_groupi_drc_bufs22682(csa_tree_add_7_25_groupi_n_1190 ,csa_tree_add_7_25_groupi_n_2365);
  not csa_tree_add_7_25_groupi_drc_bufs22683(csa_tree_add_7_25_groupi_n_1189 ,csa_tree_add_7_25_groupi_n_2365);
  not csa_tree_add_7_25_groupi_drc_bufs22686(csa_tree_add_7_25_groupi_n_1188 ,csa_tree_add_7_25_groupi_n_2389);
  not csa_tree_add_7_25_groupi_drc_bufs22687(csa_tree_add_7_25_groupi_n_1187 ,csa_tree_add_7_25_groupi_n_2389);
  not csa_tree_add_7_25_groupi_drc_bufs22690(csa_tree_add_7_25_groupi_n_1186 ,csa_tree_add_7_25_groupi_n_2356);
  not csa_tree_add_7_25_groupi_drc_bufs22691(csa_tree_add_7_25_groupi_n_1185 ,csa_tree_add_7_25_groupi_n_2356);
  not csa_tree_add_7_25_groupi_drc_bufs22694(csa_tree_add_7_25_groupi_n_1184 ,csa_tree_add_7_25_groupi_n_2391);
  not csa_tree_add_7_25_groupi_drc_bufs22695(csa_tree_add_7_25_groupi_n_1183 ,csa_tree_add_7_25_groupi_n_2391);
  not csa_tree_add_7_25_groupi_drc_bufs22698(csa_tree_add_7_25_groupi_n_1182 ,csa_tree_add_7_25_groupi_n_2398);
  not csa_tree_add_7_25_groupi_drc_bufs22699(csa_tree_add_7_25_groupi_n_1181 ,csa_tree_add_7_25_groupi_n_2398);
  not csa_tree_add_7_25_groupi_drc_bufs22702(csa_tree_add_7_25_groupi_n_1180 ,csa_tree_add_7_25_groupi_n_2397);
  not csa_tree_add_7_25_groupi_drc_bufs22703(csa_tree_add_7_25_groupi_n_1179 ,csa_tree_add_7_25_groupi_n_2397);
  not csa_tree_add_7_25_groupi_drc_bufs22706(csa_tree_add_7_25_groupi_n_1178 ,csa_tree_add_7_25_groupi_n_2399);
  not csa_tree_add_7_25_groupi_drc_bufs22707(csa_tree_add_7_25_groupi_n_1177 ,csa_tree_add_7_25_groupi_n_2399);
  not csa_tree_add_7_25_groupi_drc_bufs22710(csa_tree_add_7_25_groupi_n_1176 ,csa_tree_add_7_25_groupi_n_2363);
  not csa_tree_add_7_25_groupi_drc_bufs22711(csa_tree_add_7_25_groupi_n_1175 ,csa_tree_add_7_25_groupi_n_2363);
  not csa_tree_add_7_25_groupi_drc_bufs22714(csa_tree_add_7_25_groupi_n_1174 ,csa_tree_add_7_25_groupi_n_2401);
  not csa_tree_add_7_25_groupi_drc_bufs22715(csa_tree_add_7_25_groupi_n_1173 ,csa_tree_add_7_25_groupi_n_2401);
  not csa_tree_add_7_25_groupi_drc_bufs22718(csa_tree_add_7_25_groupi_n_1172 ,csa_tree_add_7_25_groupi_n_2393);
  not csa_tree_add_7_25_groupi_drc_bufs22719(csa_tree_add_7_25_groupi_n_1171 ,csa_tree_add_7_25_groupi_n_2393);
  not csa_tree_add_7_25_groupi_drc_bufs22722(csa_tree_add_7_25_groupi_n_1170 ,csa_tree_add_7_25_groupi_n_2354);
  not csa_tree_add_7_25_groupi_drc_bufs22723(csa_tree_add_7_25_groupi_n_1169 ,csa_tree_add_7_25_groupi_n_2354);
  not csa_tree_add_7_25_groupi_drc_bufs22726(csa_tree_add_7_25_groupi_n_1168 ,csa_tree_add_7_25_groupi_n_2364);
  not csa_tree_add_7_25_groupi_drc_bufs22727(csa_tree_add_7_25_groupi_n_1167 ,csa_tree_add_7_25_groupi_n_2364);
  not csa_tree_add_7_25_groupi_drc_bufs22730(csa_tree_add_7_25_groupi_n_1166 ,csa_tree_add_7_25_groupi_n_1164);
  not csa_tree_add_7_25_groupi_drc_bufs22731(csa_tree_add_7_25_groupi_n_1165 ,csa_tree_add_7_25_groupi_n_1164);
  not csa_tree_add_7_25_groupi_drc_bufs22732(csa_tree_add_7_25_groupi_n_1164 ,csa_tree_add_7_25_groupi_n_2869);
  not csa_tree_add_7_25_groupi_drc_bufs22734(csa_tree_add_7_25_groupi_n_1163 ,csa_tree_add_7_25_groupi_n_1161);
  not csa_tree_add_7_25_groupi_drc_bufs22735(csa_tree_add_7_25_groupi_n_1162 ,csa_tree_add_7_25_groupi_n_1161);
  not csa_tree_add_7_25_groupi_drc_bufs22736(csa_tree_add_7_25_groupi_n_1161 ,csa_tree_add_7_25_groupi_n_3523);
  not csa_tree_add_7_25_groupi_drc_bufs22738(csa_tree_add_7_25_groupi_n_1160 ,csa_tree_add_7_25_groupi_n_1158);
  not csa_tree_add_7_25_groupi_drc_bufs22739(csa_tree_add_7_25_groupi_n_1159 ,csa_tree_add_7_25_groupi_n_1158);
  not csa_tree_add_7_25_groupi_drc_bufs22740(csa_tree_add_7_25_groupi_n_1158 ,csa_tree_add_7_25_groupi_n_2869);
  not csa_tree_add_7_25_groupi_drc_bufs22742(csa_tree_add_7_25_groupi_n_1157 ,csa_tree_add_7_25_groupi_n_1155);
  not csa_tree_add_7_25_groupi_drc_bufs22743(csa_tree_add_7_25_groupi_n_1156 ,csa_tree_add_7_25_groupi_n_1155);
  not csa_tree_add_7_25_groupi_drc_bufs22744(csa_tree_add_7_25_groupi_n_1155 ,csa_tree_add_7_25_groupi_n_3531);
  not csa_tree_add_7_25_groupi_drc_bufs22746(csa_tree_add_7_25_groupi_n_1154 ,csa_tree_add_7_25_groupi_n_1152);
  not csa_tree_add_7_25_groupi_drc_bufs22747(csa_tree_add_7_25_groupi_n_1153 ,csa_tree_add_7_25_groupi_n_1152);
  not csa_tree_add_7_25_groupi_drc_bufs22748(csa_tree_add_7_25_groupi_n_1152 ,csa_tree_add_7_25_groupi_n_3527);
  not csa_tree_add_7_25_groupi_drc_bufs22750(csa_tree_add_7_25_groupi_n_1151 ,csa_tree_add_7_25_groupi_n_1149);
  not csa_tree_add_7_25_groupi_drc_bufs22751(csa_tree_add_7_25_groupi_n_1150 ,csa_tree_add_7_25_groupi_n_1149);
  not csa_tree_add_7_25_groupi_drc_bufs22752(csa_tree_add_7_25_groupi_n_1149 ,csa_tree_add_7_25_groupi_n_3527);
  not csa_tree_add_7_25_groupi_drc_bufs22754(csa_tree_add_7_25_groupi_n_1148 ,csa_tree_add_7_25_groupi_n_1146);
  not csa_tree_add_7_25_groupi_drc_bufs22755(csa_tree_add_7_25_groupi_n_1147 ,csa_tree_add_7_25_groupi_n_1146);
  not csa_tree_add_7_25_groupi_drc_bufs22756(csa_tree_add_7_25_groupi_n_1146 ,csa_tree_add_7_25_groupi_n_2778);
  not csa_tree_add_7_25_groupi_drc_bufs22758(csa_tree_add_7_25_groupi_n_1145 ,csa_tree_add_7_25_groupi_n_2347);
  not csa_tree_add_7_25_groupi_drc_bufs22760(csa_tree_add_7_25_groupi_n_2347 ,csa_tree_add_7_25_groupi_n_6938);
  not csa_tree_add_7_25_groupi_drc_bufs22762(csa_tree_add_7_25_groupi_n_1144 ,csa_tree_add_7_25_groupi_n_1143);
  not csa_tree_add_7_25_groupi_drc_bufs22764(csa_tree_add_7_25_groupi_n_1143 ,csa_tree_add_7_25_groupi_n_6560);
  not csa_tree_add_7_25_groupi_drc_bufs22766(csa_tree_add_7_25_groupi_n_1142 ,csa_tree_add_7_25_groupi_n_1140);
  not csa_tree_add_7_25_groupi_drc_bufs22767(csa_tree_add_7_25_groupi_n_1141 ,csa_tree_add_7_25_groupi_n_1140);
  not csa_tree_add_7_25_groupi_drc_bufs22768(csa_tree_add_7_25_groupi_n_1140 ,csa_tree_add_7_25_groupi_n_6884);
  not csa_tree_add_7_25_groupi_drc_bufs22770(csa_tree_add_7_25_groupi_n_1139 ,csa_tree_add_7_25_groupi_n_1138);
  not csa_tree_add_7_25_groupi_drc_bufs22772(csa_tree_add_7_25_groupi_n_1138 ,csa_tree_add_7_25_groupi_n_6718);
  not csa_tree_add_7_25_groupi_drc_bufs22774(csa_tree_add_7_25_groupi_n_1137 ,csa_tree_add_7_25_groupi_n_1136);
  not csa_tree_add_7_25_groupi_drc_bufs22776(csa_tree_add_7_25_groupi_n_1136 ,csa_tree_add_7_25_groupi_n_6382);
  not csa_tree_add_7_25_groupi_drc_bufs22778(csa_tree_add_7_25_groupi_n_1135 ,csa_tree_add_7_25_groupi_n_1134);
  not csa_tree_add_7_25_groupi_drc_bufs22780(csa_tree_add_7_25_groupi_n_1134 ,csa_tree_add_7_25_groupi_n_6463);
  not csa_tree_add_7_25_groupi_drc_bufs22782(csa_tree_add_7_25_groupi_n_1133 ,csa_tree_add_7_25_groupi_n_1132);
  not csa_tree_add_7_25_groupi_drc_bufs22784(csa_tree_add_7_25_groupi_n_1132 ,csa_tree_add_7_25_groupi_n_6806);
  not csa_tree_add_7_25_groupi_drc_bufs22786(csa_tree_add_7_25_groupi_n_1131 ,csa_tree_add_7_25_groupi_n_1129);
  not csa_tree_add_7_25_groupi_drc_bufs22787(csa_tree_add_7_25_groupi_n_1130 ,csa_tree_add_7_25_groupi_n_1129);
  not csa_tree_add_7_25_groupi_drc_bufs22788(csa_tree_add_7_25_groupi_n_1129 ,csa_tree_add_7_25_groupi_n_6806);
  not csa_tree_add_7_25_groupi_drc_bufs22790(csa_tree_add_7_25_groupi_n_1128 ,csa_tree_add_7_25_groupi_n_1126);
  not csa_tree_add_7_25_groupi_drc_bufs22791(csa_tree_add_7_25_groupi_n_1127 ,csa_tree_add_7_25_groupi_n_1126);
  not csa_tree_add_7_25_groupi_drc_bufs22792(csa_tree_add_7_25_groupi_n_1126 ,csa_tree_add_7_25_groupi_n_6718);
  not csa_tree_add_7_25_groupi_drc_bufs22794(csa_tree_add_7_25_groupi_n_1125 ,csa_tree_add_7_25_groupi_n_1124);
  not csa_tree_add_7_25_groupi_drc_bufs22796(csa_tree_add_7_25_groupi_n_1124 ,csa_tree_add_7_25_groupi_n_6647);
  not csa_tree_add_7_25_groupi_drc_bufs22798(csa_tree_add_7_25_groupi_n_1123 ,csa_tree_add_7_25_groupi_n_1121);
  not csa_tree_add_7_25_groupi_drc_bufs22799(csa_tree_add_7_25_groupi_n_1122 ,csa_tree_add_7_25_groupi_n_1121);
  not csa_tree_add_7_25_groupi_drc_bufs22800(csa_tree_add_7_25_groupi_n_1121 ,csa_tree_add_7_25_groupi_n_6938);
  not csa_tree_add_7_25_groupi_drc_bufs22802(csa_tree_add_7_25_groupi_n_1120 ,csa_tree_add_7_25_groupi_n_1118);
  not csa_tree_add_7_25_groupi_drc_bufs22803(csa_tree_add_7_25_groupi_n_1119 ,csa_tree_add_7_25_groupi_n_1118);
  not csa_tree_add_7_25_groupi_drc_bufs22804(csa_tree_add_7_25_groupi_n_1118 ,csa_tree_add_7_25_groupi_n_6647);
  not csa_tree_add_7_25_groupi_drc_bufs22806(csa_tree_add_7_25_groupi_n_1117 ,csa_tree_add_7_25_groupi_n_2339);
  not csa_tree_add_7_25_groupi_drc_bufs22808(csa_tree_add_7_25_groupi_n_2339 ,csa_tree_add_7_25_groupi_n_3521);
  not csa_tree_add_7_25_groupi_drc_bufs22810(csa_tree_add_7_25_groupi_n_1116 ,csa_tree_add_7_25_groupi_n_2338);
  not csa_tree_add_7_25_groupi_drc_bufs22812(csa_tree_add_7_25_groupi_n_2338 ,csa_tree_add_7_25_groupi_n_2867);
  not csa_tree_add_7_25_groupi_drc_bufs22814(csa_tree_add_7_25_groupi_n_1115 ,csa_tree_add_7_25_groupi_n_1113);
  not csa_tree_add_7_25_groupi_drc_bufs22815(csa_tree_add_7_25_groupi_n_1114 ,csa_tree_add_7_25_groupi_n_1113);
  not csa_tree_add_7_25_groupi_drc_bufs22816(csa_tree_add_7_25_groupi_n_1113 ,csa_tree_add_7_25_groupi_n_6949);
  not csa_tree_add_7_25_groupi_drc_bufs22818(csa_tree_add_7_25_groupi_n_1112 ,csa_tree_add_7_25_groupi_n_2328);
  not csa_tree_add_7_25_groupi_drc_bufs22820(csa_tree_add_7_25_groupi_n_2328 ,csa_tree_add_7_25_groupi_n_2784);
  not csa_tree_add_7_25_groupi_drc_bufs22822(csa_tree_add_7_25_groupi_n_1111 ,csa_tree_add_7_25_groupi_n_2332);
  not csa_tree_add_7_25_groupi_drc_bufs22824(csa_tree_add_7_25_groupi_n_2332 ,csa_tree_add_7_25_groupi_n_2791);
  not csa_tree_add_7_25_groupi_drc_bufs22826(csa_tree_add_7_25_groupi_n_1110 ,csa_tree_add_7_25_groupi_n_2331);
  not csa_tree_add_7_25_groupi_drc_bufs22828(csa_tree_add_7_25_groupi_n_2331 ,csa_tree_add_7_25_groupi_n_2787);
  not csa_tree_add_7_25_groupi_drc_bufs22832(csa_tree_add_7_25_groupi_n_2333 ,csa_tree_add_7_25_groupi_n_2791);
  not csa_tree_add_7_25_groupi_drc_bufs22834(csa_tree_add_7_25_groupi_n_1109 ,csa_tree_add_7_25_groupi_n_2343);
  not csa_tree_add_7_25_groupi_drc_bufs22836(csa_tree_add_7_25_groupi_n_2343 ,csa_tree_add_7_25_groupi_n_4554);
  not csa_tree_add_7_25_groupi_drc_bufs22838(csa_tree_add_7_25_groupi_n_1108 ,csa_tree_add_7_25_groupi_n_2345);
  not csa_tree_add_7_25_groupi_drc_bufs22840(csa_tree_add_7_25_groupi_n_2345 ,csa_tree_add_7_25_groupi_n_5156);
  not csa_tree_add_7_25_groupi_drc_bufs22842(csa_tree_add_7_25_groupi_n_1107 ,csa_tree_add_7_25_groupi_n_2344);
  not csa_tree_add_7_25_groupi_drc_bufs22844(csa_tree_add_7_25_groupi_n_2344 ,csa_tree_add_7_25_groupi_n_4883);
  not csa_tree_add_7_25_groupi_drc_bufs22846(csa_tree_add_7_25_groupi_n_1106 ,csa_tree_add_7_25_groupi_n_1105);
  not csa_tree_add_7_25_groupi_drc_bufs22848(csa_tree_add_7_25_groupi_n_1105 ,csa_tree_add_7_25_groupi_n_2792);
  not csa_tree_add_7_25_groupi_drc_bufs22851(csa_tree_add_7_25_groupi_n_1104 ,csa_tree_add_7_25_groupi_n_1103);
  not csa_tree_add_7_25_groupi_drc_bufs22852(csa_tree_add_7_25_groupi_n_1103 ,csa_tree_add_7_25_groupi_n_5074);
  not csa_tree_add_7_25_groupi_drc_bufs22855(csa_tree_add_7_25_groupi_n_1102 ,csa_tree_add_7_25_groupi_n_1101);
  not csa_tree_add_7_25_groupi_drc_bufs22856(csa_tree_add_7_25_groupi_n_1101 ,csa_tree_add_7_25_groupi_n_4771);
  not csa_tree_add_7_25_groupi_drc_bufs22859(csa_tree_add_7_25_groupi_n_1100 ,csa_tree_add_7_25_groupi_n_1099);
  not csa_tree_add_7_25_groupi_drc_bufs22860(csa_tree_add_7_25_groupi_n_1099 ,csa_tree_add_7_25_groupi_n_4554);
  not csa_tree_add_7_25_groupi_drc_bufs22863(csa_tree_add_7_25_groupi_n_1098 ,csa_tree_add_7_25_groupi_n_1097);
  not csa_tree_add_7_25_groupi_drc_bufs22864(csa_tree_add_7_25_groupi_n_1097 ,csa_tree_add_7_25_groupi_n_4883);
  not csa_tree_add_7_25_groupi_drc_bufs22867(csa_tree_add_7_25_groupi_n_1096 ,csa_tree_add_7_25_groupi_n_1095);
  not csa_tree_add_7_25_groupi_drc_bufs22868(csa_tree_add_7_25_groupi_n_1095 ,csa_tree_add_7_25_groupi_n_5156);
  not csa_tree_add_7_25_groupi_drc_bufs22871(csa_tree_add_7_25_groupi_n_1094 ,csa_tree_add_7_25_groupi_n_1093);
  not csa_tree_add_7_25_groupi_drc_bufs22872(csa_tree_add_7_25_groupi_n_1093 ,csa_tree_add_7_25_groupi_n_4442);
  not csa_tree_add_7_25_groupi_drc_bufs22875(csa_tree_add_7_25_groupi_n_1092 ,csa_tree_add_7_25_groupi_n_1091);
  not csa_tree_add_7_25_groupi_drc_bufs22876(csa_tree_add_7_25_groupi_n_1091 ,csa_tree_add_7_25_groupi_n_2383);
  not csa_tree_add_7_25_groupi_drc_bufs22886(csa_tree_add_7_25_groupi_n_1090 ,csa_tree_add_7_25_groupi_n_2342);
  not csa_tree_add_7_25_groupi_drc_bufs22887(csa_tree_add_7_25_groupi_n_2342 ,csa_tree_add_7_25_groupi_n_4442);
  not csa_tree_add_7_25_groupi_drc_bufs22892(csa_tree_add_7_25_groupi_n_1089 ,csa_tree_add_7_25_groupi_n_1088);
  not csa_tree_add_7_25_groupi_drc_bufs22893(csa_tree_add_7_25_groupi_n_1088 ,csa_tree_add_7_25_groupi_n_1955);
  not csa_tree_add_7_25_groupi_drc_bufs22895(csa_tree_add_7_25_groupi_n_1087 ,csa_tree_add_7_25_groupi_n_1085);
  not csa_tree_add_7_25_groupi_drc_bufs22896(csa_tree_add_7_25_groupi_n_1086 ,csa_tree_add_7_25_groupi_n_1085);
  not csa_tree_add_7_25_groupi_drc_bufs22897(csa_tree_add_7_25_groupi_n_1085 ,csa_tree_add_7_25_groupi_n_2313);
  not csa_tree_add_7_25_groupi_drc_bufs22899(csa_tree_add_7_25_groupi_n_1084 ,csa_tree_add_7_25_groupi_n_1082);
  not csa_tree_add_7_25_groupi_drc_bufs22900(csa_tree_add_7_25_groupi_n_1083 ,csa_tree_add_7_25_groupi_n_1082);
  not csa_tree_add_7_25_groupi_drc_bufs22901(csa_tree_add_7_25_groupi_n_1082 ,csa_tree_add_7_25_groupi_n_2269);
  not csa_tree_add_7_25_groupi_drc_bufs22903(csa_tree_add_7_25_groupi_n_1081 ,csa_tree_add_7_25_groupi_n_1079);
  not csa_tree_add_7_25_groupi_drc_bufs22904(csa_tree_add_7_25_groupi_n_1080 ,csa_tree_add_7_25_groupi_n_1079);
  not csa_tree_add_7_25_groupi_drc_bufs22905(csa_tree_add_7_25_groupi_n_1079 ,csa_tree_add_7_25_groupi_n_2292);
  not csa_tree_add_7_25_groupi_drc_bufs22907(csa_tree_add_7_25_groupi_n_1078 ,csa_tree_add_7_25_groupi_n_1076);
  not csa_tree_add_7_25_groupi_drc_bufs22908(csa_tree_add_7_25_groupi_n_1077 ,csa_tree_add_7_25_groupi_n_1076);
  not csa_tree_add_7_25_groupi_drc_bufs22909(csa_tree_add_7_25_groupi_n_1076 ,csa_tree_add_7_25_groupi_n_2289);
  not csa_tree_add_7_25_groupi_drc_bufs22911(csa_tree_add_7_25_groupi_n_1075 ,csa_tree_add_7_25_groupi_n_1073);
  not csa_tree_add_7_25_groupi_drc_bufs22912(csa_tree_add_7_25_groupi_n_1074 ,csa_tree_add_7_25_groupi_n_1073);
  not csa_tree_add_7_25_groupi_drc_bufs22913(csa_tree_add_7_25_groupi_n_1073 ,csa_tree_add_7_25_groupi_n_2268);
  not csa_tree_add_7_25_groupi_drc_bufs22915(csa_tree_add_7_25_groupi_n_1072 ,csa_tree_add_7_25_groupi_n_1070);
  not csa_tree_add_7_25_groupi_drc_bufs22916(csa_tree_add_7_25_groupi_n_1071 ,csa_tree_add_7_25_groupi_n_1070);
  not csa_tree_add_7_25_groupi_drc_bufs22917(csa_tree_add_7_25_groupi_n_1070 ,csa_tree_add_7_25_groupi_n_2288);
  not csa_tree_add_7_25_groupi_drc_bufs22919(csa_tree_add_7_25_groupi_n_1069 ,csa_tree_add_7_25_groupi_n_1067);
  not csa_tree_add_7_25_groupi_drc_bufs22920(csa_tree_add_7_25_groupi_n_1068 ,csa_tree_add_7_25_groupi_n_1067);
  not csa_tree_add_7_25_groupi_drc_bufs22921(csa_tree_add_7_25_groupi_n_1067 ,csa_tree_add_7_25_groupi_n_2312);
  not csa_tree_add_7_25_groupi_drc_bufs22923(csa_tree_add_7_25_groupi_n_1066 ,csa_tree_add_7_25_groupi_n_1064);
  not csa_tree_add_7_25_groupi_drc_bufs22924(csa_tree_add_7_25_groupi_n_1065 ,csa_tree_add_7_25_groupi_n_1064);
  not csa_tree_add_7_25_groupi_drc_bufs22925(csa_tree_add_7_25_groupi_n_1064 ,csa_tree_add_7_25_groupi_n_2297);
  not csa_tree_add_7_25_groupi_drc_bufs22927(csa_tree_add_7_25_groupi_n_1063 ,csa_tree_add_7_25_groupi_n_1061);
  not csa_tree_add_7_25_groupi_drc_bufs22928(csa_tree_add_7_25_groupi_n_1062 ,csa_tree_add_7_25_groupi_n_1061);
  not csa_tree_add_7_25_groupi_drc_bufs22929(csa_tree_add_7_25_groupi_n_1061 ,csa_tree_add_7_25_groupi_n_2293);
  not csa_tree_add_7_25_groupi_drc_bufs22931(csa_tree_add_7_25_groupi_n_1060 ,csa_tree_add_7_25_groupi_n_1058);
  not csa_tree_add_7_25_groupi_drc_bufs22932(csa_tree_add_7_25_groupi_n_1059 ,csa_tree_add_7_25_groupi_n_1058);
  not csa_tree_add_7_25_groupi_drc_bufs22933(csa_tree_add_7_25_groupi_n_1058 ,csa_tree_add_7_25_groupi_n_2305);
  not csa_tree_add_7_25_groupi_drc_bufs22935(csa_tree_add_7_25_groupi_n_1057 ,csa_tree_add_7_25_groupi_n_1055);
  not csa_tree_add_7_25_groupi_drc_bufs22936(csa_tree_add_7_25_groupi_n_1056 ,csa_tree_add_7_25_groupi_n_1055);
  not csa_tree_add_7_25_groupi_drc_bufs22937(csa_tree_add_7_25_groupi_n_1055 ,csa_tree_add_7_25_groupi_n_2304);
  not csa_tree_add_7_25_groupi_drc_bufs22939(csa_tree_add_7_25_groupi_n_1054 ,csa_tree_add_7_25_groupi_n_1052);
  not csa_tree_add_7_25_groupi_drc_bufs22940(csa_tree_add_7_25_groupi_n_1053 ,csa_tree_add_7_25_groupi_n_1052);
  not csa_tree_add_7_25_groupi_drc_bufs22941(csa_tree_add_7_25_groupi_n_1052 ,csa_tree_add_7_25_groupi_n_2273);
  not csa_tree_add_7_25_groupi_drc_bufs22943(csa_tree_add_7_25_groupi_n_1051 ,csa_tree_add_7_25_groupi_n_1049);
  not csa_tree_add_7_25_groupi_drc_bufs22944(csa_tree_add_7_25_groupi_n_1050 ,csa_tree_add_7_25_groupi_n_1049);
  not csa_tree_add_7_25_groupi_drc_bufs22945(csa_tree_add_7_25_groupi_n_1049 ,csa_tree_add_7_25_groupi_n_2265);
  not csa_tree_add_7_25_groupi_drc_bufs22947(csa_tree_add_7_25_groupi_n_1048 ,csa_tree_add_7_25_groupi_n_1046);
  not csa_tree_add_7_25_groupi_drc_bufs22948(csa_tree_add_7_25_groupi_n_1047 ,csa_tree_add_7_25_groupi_n_1046);
  not csa_tree_add_7_25_groupi_drc_bufs22949(csa_tree_add_7_25_groupi_n_1046 ,csa_tree_add_7_25_groupi_n_2285);
  not csa_tree_add_7_25_groupi_drc_bufs22951(csa_tree_add_7_25_groupi_n_1045 ,csa_tree_add_7_25_groupi_n_1043);
  not csa_tree_add_7_25_groupi_drc_bufs22952(csa_tree_add_7_25_groupi_n_1044 ,csa_tree_add_7_25_groupi_n_1043);
  not csa_tree_add_7_25_groupi_drc_bufs22953(csa_tree_add_7_25_groupi_n_1043 ,csa_tree_add_7_25_groupi_n_2284);
  not csa_tree_add_7_25_groupi_drc_bufs22955(csa_tree_add_7_25_groupi_n_1042 ,csa_tree_add_7_25_groupi_n_1040);
  not csa_tree_add_7_25_groupi_drc_bufs22956(csa_tree_add_7_25_groupi_n_1041 ,csa_tree_add_7_25_groupi_n_1040);
  not csa_tree_add_7_25_groupi_drc_bufs22957(csa_tree_add_7_25_groupi_n_1040 ,csa_tree_add_7_25_groupi_n_2309);
  not csa_tree_add_7_25_groupi_drc_bufs22959(csa_tree_add_7_25_groupi_n_1039 ,csa_tree_add_7_25_groupi_n_1037);
  not csa_tree_add_7_25_groupi_drc_bufs22960(csa_tree_add_7_25_groupi_n_1038 ,csa_tree_add_7_25_groupi_n_1037);
  not csa_tree_add_7_25_groupi_drc_bufs22961(csa_tree_add_7_25_groupi_n_1037 ,csa_tree_add_7_25_groupi_n_2272);
  not csa_tree_add_7_25_groupi_drc_bufs22963(csa_tree_add_7_25_groupi_n_1036 ,csa_tree_add_7_25_groupi_n_1034);
  not csa_tree_add_7_25_groupi_drc_bufs22964(csa_tree_add_7_25_groupi_n_1035 ,csa_tree_add_7_25_groupi_n_1034);
  not csa_tree_add_7_25_groupi_drc_bufs22965(csa_tree_add_7_25_groupi_n_1034 ,csa_tree_add_7_25_groupi_n_2261);
  not csa_tree_add_7_25_groupi_drc_bufs22967(csa_tree_add_7_25_groupi_n_1033 ,csa_tree_add_7_25_groupi_n_1031);
  not csa_tree_add_7_25_groupi_drc_bufs22968(csa_tree_add_7_25_groupi_n_1032 ,csa_tree_add_7_25_groupi_n_1031);
  not csa_tree_add_7_25_groupi_drc_bufs22969(csa_tree_add_7_25_groupi_n_1031 ,csa_tree_add_7_25_groupi_n_2281);
  not csa_tree_add_7_25_groupi_drc_bufs22971(csa_tree_add_7_25_groupi_n_1030 ,csa_tree_add_7_25_groupi_n_1028);
  not csa_tree_add_7_25_groupi_drc_bufs22972(csa_tree_add_7_25_groupi_n_1029 ,csa_tree_add_7_25_groupi_n_1028);
  not csa_tree_add_7_25_groupi_drc_bufs22973(csa_tree_add_7_25_groupi_n_1028 ,csa_tree_add_7_25_groupi_n_2280);
  not csa_tree_add_7_25_groupi_drc_bufs22975(csa_tree_add_7_25_groupi_n_1027 ,csa_tree_add_7_25_groupi_n_1025);
  not csa_tree_add_7_25_groupi_drc_bufs22976(csa_tree_add_7_25_groupi_n_1026 ,csa_tree_add_7_25_groupi_n_1025);
  not csa_tree_add_7_25_groupi_drc_bufs22977(csa_tree_add_7_25_groupi_n_1025 ,csa_tree_add_7_25_groupi_n_2311);
  not csa_tree_add_7_25_groupi_drc_bufs22979(csa_tree_add_7_25_groupi_n_1024 ,csa_tree_add_7_25_groupi_n_1022);
  not csa_tree_add_7_25_groupi_drc_bufs22980(csa_tree_add_7_25_groupi_n_1023 ,csa_tree_add_7_25_groupi_n_1022);
  not csa_tree_add_7_25_groupi_drc_bufs22981(csa_tree_add_7_25_groupi_n_1022 ,csa_tree_add_7_25_groupi_n_2301);
  not csa_tree_add_7_25_groupi_drc_bufs22983(csa_tree_add_7_25_groupi_n_1021 ,csa_tree_add_7_25_groupi_n_1019);
  not csa_tree_add_7_25_groupi_drc_bufs22984(csa_tree_add_7_25_groupi_n_1020 ,csa_tree_add_7_25_groupi_n_1019);
  not csa_tree_add_7_25_groupi_drc_bufs22985(csa_tree_add_7_25_groupi_n_1019 ,csa_tree_add_7_25_groupi_n_2277);
  not csa_tree_add_7_25_groupi_drc_bufs22987(csa_tree_add_7_25_groupi_n_1018 ,csa_tree_add_7_25_groupi_n_1016);
  not csa_tree_add_7_25_groupi_drc_bufs22988(csa_tree_add_7_25_groupi_n_1017 ,csa_tree_add_7_25_groupi_n_1016);
  not csa_tree_add_7_25_groupi_drc_bufs22989(csa_tree_add_7_25_groupi_n_1016 ,csa_tree_add_7_25_groupi_n_2296);
  not csa_tree_add_7_25_groupi_drc_bufs22991(csa_tree_add_7_25_groupi_n_1015 ,csa_tree_add_7_25_groupi_n_1013);
  not csa_tree_add_7_25_groupi_drc_bufs22992(csa_tree_add_7_25_groupi_n_1014 ,csa_tree_add_7_25_groupi_n_1013);
  not csa_tree_add_7_25_groupi_drc_bufs22993(csa_tree_add_7_25_groupi_n_1013 ,csa_tree_add_7_25_groupi_n_2308);
  not csa_tree_add_7_25_groupi_drc_bufs22995(csa_tree_add_7_25_groupi_n_1012 ,csa_tree_add_7_25_groupi_n_1010);
  not csa_tree_add_7_25_groupi_drc_bufs22996(csa_tree_add_7_25_groupi_n_1011 ,csa_tree_add_7_25_groupi_n_1010);
  not csa_tree_add_7_25_groupi_drc_bufs22997(csa_tree_add_7_25_groupi_n_1010 ,csa_tree_add_7_25_groupi_n_2300);
  not csa_tree_add_7_25_groupi_drc_bufs22999(csa_tree_add_7_25_groupi_n_1009 ,csa_tree_add_7_25_groupi_n_1007);
  not csa_tree_add_7_25_groupi_drc_bufs23000(csa_tree_add_7_25_groupi_n_1008 ,csa_tree_add_7_25_groupi_n_1007);
  not csa_tree_add_7_25_groupi_drc_bufs23001(csa_tree_add_7_25_groupi_n_1007 ,csa_tree_add_7_25_groupi_n_2276);
  not csa_tree_add_7_25_groupi_drc_bufs23003(csa_tree_add_7_25_groupi_n_1006 ,csa_tree_add_7_25_groupi_n_1004);
  not csa_tree_add_7_25_groupi_drc_bufs23004(csa_tree_add_7_25_groupi_n_1005 ,csa_tree_add_7_25_groupi_n_1004);
  not csa_tree_add_7_25_groupi_drc_bufs23005(csa_tree_add_7_25_groupi_n_1004 ,csa_tree_add_7_25_groupi_n_2307);
  not csa_tree_add_7_25_groupi_drc_bufs23007(csa_tree_add_7_25_groupi_n_1003 ,csa_tree_add_7_25_groupi_n_1001);
  not csa_tree_add_7_25_groupi_drc_bufs23008(csa_tree_add_7_25_groupi_n_1002 ,csa_tree_add_7_25_groupi_n_1001);
  not csa_tree_add_7_25_groupi_drc_bufs23009(csa_tree_add_7_25_groupi_n_1001 ,csa_tree_add_7_25_groupi_n_2366);
  not csa_tree_add_7_25_groupi_drc_bufs23011(csa_tree_add_7_25_groupi_n_1000 ,csa_tree_add_7_25_groupi_n_998);
  not csa_tree_add_7_25_groupi_drc_bufs23012(csa_tree_add_7_25_groupi_n_999 ,csa_tree_add_7_25_groupi_n_998);
  not csa_tree_add_7_25_groupi_drc_bufs23013(csa_tree_add_7_25_groupi_n_998 ,csa_tree_add_7_25_groupi_n_2367);
  not csa_tree_add_7_25_groupi_drc_bufs23015(csa_tree_add_7_25_groupi_n_997 ,csa_tree_add_7_25_groupi_n_995);
  not csa_tree_add_7_25_groupi_drc_bufs23016(csa_tree_add_7_25_groupi_n_996 ,csa_tree_add_7_25_groupi_n_995);
  not csa_tree_add_7_25_groupi_drc_bufs23017(csa_tree_add_7_25_groupi_n_995 ,csa_tree_add_7_25_groupi_n_2366);
  not csa_tree_add_7_25_groupi_drc_bufs23020(csa_tree_add_7_25_groupi_n_994 ,csa_tree_add_7_25_groupi_n_993);
  not csa_tree_add_7_25_groupi_drc_bufs23021(csa_tree_add_7_25_groupi_n_993 ,csa_tree_add_7_25_groupi_n_1952);
  not csa_tree_add_7_25_groupi_drc_bufs23023(csa_tree_add_7_25_groupi_n_992 ,csa_tree_add_7_25_groupi_n_990);
  not csa_tree_add_7_25_groupi_drc_bufs23024(csa_tree_add_7_25_groupi_n_991 ,csa_tree_add_7_25_groupi_n_990);
  not csa_tree_add_7_25_groupi_drc_bufs23025(csa_tree_add_7_25_groupi_n_990 ,csa_tree_add_7_25_groupi_n_2887);
  not csa_tree_add_7_25_groupi_drc_bufs23028(csa_tree_add_7_25_groupi_n_989 ,csa_tree_add_7_25_groupi_n_988);
  not csa_tree_add_7_25_groupi_drc_bufs23029(csa_tree_add_7_25_groupi_n_988 ,csa_tree_add_7_25_groupi_n_1949);
  not csa_tree_add_7_25_groupi_drc_bufs23031(csa_tree_add_7_25_groupi_n_987 ,csa_tree_add_7_25_groupi_n_985);
  not csa_tree_add_7_25_groupi_drc_bufs23032(csa_tree_add_7_25_groupi_n_986 ,csa_tree_add_7_25_groupi_n_985);
  not csa_tree_add_7_25_groupi_drc_bufs23033(csa_tree_add_7_25_groupi_n_985 ,csa_tree_add_7_25_groupi_n_2266);
  not csa_tree_add_7_25_groupi_drc_bufs23035(csa_tree_add_7_25_groupi_n_984 ,csa_tree_add_7_25_groupi_n_982);
  not csa_tree_add_7_25_groupi_drc_bufs23036(csa_tree_add_7_25_groupi_n_983 ,csa_tree_add_7_25_groupi_n_982);
  not csa_tree_add_7_25_groupi_drc_bufs23037(csa_tree_add_7_25_groupi_n_982 ,csa_tree_add_7_25_groupi_n_2263);
  not csa_tree_add_7_25_groupi_drc_bufs23039(csa_tree_add_7_25_groupi_n_981 ,csa_tree_add_7_25_groupi_n_979);
  not csa_tree_add_7_25_groupi_drc_bufs23040(csa_tree_add_7_25_groupi_n_980 ,csa_tree_add_7_25_groupi_n_979);
  not csa_tree_add_7_25_groupi_drc_bufs23041(csa_tree_add_7_25_groupi_n_979 ,csa_tree_add_7_25_groupi_n_2262);
  not csa_tree_add_7_25_groupi_drc_bufs23043(csa_tree_add_7_25_groupi_n_978 ,csa_tree_add_7_25_groupi_n_976);
  not csa_tree_add_7_25_groupi_drc_bufs23044(csa_tree_add_7_25_groupi_n_977 ,csa_tree_add_7_25_groupi_n_976);
  not csa_tree_add_7_25_groupi_drc_bufs23045(csa_tree_add_7_25_groupi_n_976 ,csa_tree_add_7_25_groupi_n_2294);
  not csa_tree_add_7_25_groupi_drc_bufs23047(csa_tree_add_7_25_groupi_n_975 ,csa_tree_add_7_25_groupi_n_973);
  not csa_tree_add_7_25_groupi_drc_bufs23048(csa_tree_add_7_25_groupi_n_974 ,csa_tree_add_7_25_groupi_n_973);
  not csa_tree_add_7_25_groupi_drc_bufs23049(csa_tree_add_7_25_groupi_n_973 ,csa_tree_add_7_25_groupi_n_2258);
  not csa_tree_add_7_25_groupi_drc_bufs23051(csa_tree_add_7_25_groupi_n_972 ,csa_tree_add_7_25_groupi_n_970);
  not csa_tree_add_7_25_groupi_drc_bufs23052(csa_tree_add_7_25_groupi_n_971 ,csa_tree_add_7_25_groupi_n_970);
  not csa_tree_add_7_25_groupi_drc_bufs23053(csa_tree_add_7_25_groupi_n_970 ,csa_tree_add_7_25_groupi_n_2290);
  not csa_tree_add_7_25_groupi_drc_bufs23055(csa_tree_add_7_25_groupi_n_969 ,csa_tree_add_7_25_groupi_n_967);
  not csa_tree_add_7_25_groupi_drc_bufs23056(csa_tree_add_7_25_groupi_n_968 ,csa_tree_add_7_25_groupi_n_967);
  not csa_tree_add_7_25_groupi_drc_bufs23057(csa_tree_add_7_25_groupi_n_967 ,csa_tree_add_7_25_groupi_n_2286);
  not csa_tree_add_7_25_groupi_drc_bufs23059(csa_tree_add_7_25_groupi_n_966 ,csa_tree_add_7_25_groupi_n_964);
  not csa_tree_add_7_25_groupi_drc_bufs23060(csa_tree_add_7_25_groupi_n_965 ,csa_tree_add_7_25_groupi_n_964);
  not csa_tree_add_7_25_groupi_drc_bufs23061(csa_tree_add_7_25_groupi_n_964 ,csa_tree_add_7_25_groupi_n_2250);
  not csa_tree_add_7_25_groupi_drc_bufs23063(csa_tree_add_7_25_groupi_n_963 ,csa_tree_add_7_25_groupi_n_961);
  not csa_tree_add_7_25_groupi_drc_bufs23064(csa_tree_add_7_25_groupi_n_962 ,csa_tree_add_7_25_groupi_n_961);
  not csa_tree_add_7_25_groupi_drc_bufs23065(csa_tree_add_7_25_groupi_n_961 ,csa_tree_add_7_25_groupi_n_2282);
  not csa_tree_add_7_25_groupi_drc_bufs23067(csa_tree_add_7_25_groupi_n_960 ,csa_tree_add_7_25_groupi_n_958);
  not csa_tree_add_7_25_groupi_drc_bufs23068(csa_tree_add_7_25_groupi_n_959 ,csa_tree_add_7_25_groupi_n_958);
  not csa_tree_add_7_25_groupi_drc_bufs23069(csa_tree_add_7_25_groupi_n_958 ,csa_tree_add_7_25_groupi_n_2302);
  not csa_tree_add_7_25_groupi_drc_bufs23071(csa_tree_add_7_25_groupi_n_957 ,csa_tree_add_7_25_groupi_n_955);
  not csa_tree_add_7_25_groupi_drc_bufs23072(csa_tree_add_7_25_groupi_n_956 ,csa_tree_add_7_25_groupi_n_955);
  not csa_tree_add_7_25_groupi_drc_bufs23073(csa_tree_add_7_25_groupi_n_955 ,csa_tree_add_7_25_groupi_n_2278);
  not csa_tree_add_7_25_groupi_drc_bufs23075(csa_tree_add_7_25_groupi_n_954 ,csa_tree_add_7_25_groupi_n_952);
  not csa_tree_add_7_25_groupi_drc_bufs23076(csa_tree_add_7_25_groupi_n_953 ,csa_tree_add_7_25_groupi_n_952);
  not csa_tree_add_7_25_groupi_drc_bufs23077(csa_tree_add_7_25_groupi_n_952 ,csa_tree_add_7_25_groupi_n_2274);
  not csa_tree_add_7_25_groupi_drc_bufs23079(csa_tree_add_7_25_groupi_n_951 ,csa_tree_add_7_25_groupi_n_949);
  not csa_tree_add_7_25_groupi_drc_bufs23080(csa_tree_add_7_25_groupi_n_950 ,csa_tree_add_7_25_groupi_n_949);
  not csa_tree_add_7_25_groupi_drc_bufs23081(csa_tree_add_7_25_groupi_n_949 ,csa_tree_add_7_25_groupi_n_2403);
  not csa_tree_add_7_25_groupi_drc_bufs23083(csa_tree_add_7_25_groupi_n_948 ,csa_tree_add_7_25_groupi_n_946);
  not csa_tree_add_7_25_groupi_drc_bufs23084(csa_tree_add_7_25_groupi_n_947 ,csa_tree_add_7_25_groupi_n_946);
  not csa_tree_add_7_25_groupi_drc_bufs23085(csa_tree_add_7_25_groupi_n_946 ,csa_tree_add_7_25_groupi_n_2270);
  not csa_tree_add_7_25_groupi_drc_bufs23087(csa_tree_add_7_25_groupi_n_945 ,csa_tree_add_7_25_groupi_n_943);
  not csa_tree_add_7_25_groupi_drc_bufs23088(csa_tree_add_7_25_groupi_n_944 ,csa_tree_add_7_25_groupi_n_943);
  not csa_tree_add_7_25_groupi_drc_bufs23089(csa_tree_add_7_25_groupi_n_943 ,csa_tree_add_7_25_groupi_n_2298);
  not csa_tree_add_7_25_groupi_drc_bufs23091(csa_tree_add_7_25_groupi_n_942 ,csa_tree_add_7_25_groupi_n_940);
  not csa_tree_add_7_25_groupi_drc_bufs23092(csa_tree_add_7_25_groupi_n_941 ,csa_tree_add_7_25_groupi_n_940);
  not csa_tree_add_7_25_groupi_drc_bufs23093(csa_tree_add_7_25_groupi_n_940 ,csa_tree_add_7_25_groupi_n_3535);
  not csa_tree_add_7_25_groupi_drc_bufs23095(csa_tree_add_7_25_groupi_n_939 ,csa_tree_add_7_25_groupi_n_937);
  not csa_tree_add_7_25_groupi_drc_bufs23096(csa_tree_add_7_25_groupi_n_938 ,csa_tree_add_7_25_groupi_n_937);
  not csa_tree_add_7_25_groupi_drc_bufs23097(csa_tree_add_7_25_groupi_n_937 ,csa_tree_add_7_25_groupi_n_2257);
  not csa_tree_add_7_25_groupi_drc_bufs23099(csa_tree_add_7_25_groupi_n_936 ,csa_tree_add_7_25_groupi_n_934);
  not csa_tree_add_7_25_groupi_drc_bufs23100(csa_tree_add_7_25_groupi_n_935 ,csa_tree_add_7_25_groupi_n_934);
  not csa_tree_add_7_25_groupi_drc_bufs23101(csa_tree_add_7_25_groupi_n_934 ,csa_tree_add_7_25_groupi_n_2256);
  not csa_tree_add_7_25_groupi_drc_bufs23103(csa_tree_add_7_25_groupi_n_933 ,csa_tree_add_7_25_groupi_n_931);
  not csa_tree_add_7_25_groupi_drc_bufs23104(csa_tree_add_7_25_groupi_n_932 ,csa_tree_add_7_25_groupi_n_931);
  not csa_tree_add_7_25_groupi_drc_bufs23105(csa_tree_add_7_25_groupi_n_931 ,csa_tree_add_7_25_groupi_n_2283);
  not csa_tree_add_7_25_groupi_drc_bufs23107(csa_tree_add_7_25_groupi_n_930 ,csa_tree_add_7_25_groupi_n_928);
  not csa_tree_add_7_25_groupi_drc_bufs23108(csa_tree_add_7_25_groupi_n_929 ,csa_tree_add_7_25_groupi_n_928);
  not csa_tree_add_7_25_groupi_drc_bufs23109(csa_tree_add_7_25_groupi_n_928 ,csa_tree_add_7_25_groupi_n_2283);
  not csa_tree_add_7_25_groupi_drc_bufs23111(csa_tree_add_7_25_groupi_n_927 ,csa_tree_add_7_25_groupi_n_925);
  not csa_tree_add_7_25_groupi_drc_bufs23112(csa_tree_add_7_25_groupi_n_926 ,csa_tree_add_7_25_groupi_n_925);
  not csa_tree_add_7_25_groupi_drc_bufs23113(csa_tree_add_7_25_groupi_n_925 ,csa_tree_add_7_25_groupi_n_2266);
  not csa_tree_add_7_25_groupi_drc_bufs23115(csa_tree_add_7_25_groupi_n_924 ,csa_tree_add_7_25_groupi_n_922);
  not csa_tree_add_7_25_groupi_drc_bufs23116(csa_tree_add_7_25_groupi_n_923 ,csa_tree_add_7_25_groupi_n_922);
  not csa_tree_add_7_25_groupi_drc_bufs23117(csa_tree_add_7_25_groupi_n_922 ,csa_tree_add_7_25_groupi_n_2303);
  not csa_tree_add_7_25_groupi_drc_bufs23119(csa_tree_add_7_25_groupi_n_921 ,csa_tree_add_7_25_groupi_n_919);
  not csa_tree_add_7_25_groupi_drc_bufs23120(csa_tree_add_7_25_groupi_n_920 ,csa_tree_add_7_25_groupi_n_919);
  not csa_tree_add_7_25_groupi_drc_bufs23121(csa_tree_add_7_25_groupi_n_919 ,csa_tree_add_7_25_groupi_n_2303);
  not csa_tree_add_7_25_groupi_drc_bufs23123(csa_tree_add_7_25_groupi_n_918 ,csa_tree_add_7_25_groupi_n_916);
  not csa_tree_add_7_25_groupi_drc_bufs23124(csa_tree_add_7_25_groupi_n_917 ,csa_tree_add_7_25_groupi_n_916);
  not csa_tree_add_7_25_groupi_drc_bufs23125(csa_tree_add_7_25_groupi_n_916 ,csa_tree_add_7_25_groupi_n_2263);
  not csa_tree_add_7_25_groupi_drc_bufs23127(csa_tree_add_7_25_groupi_n_915 ,csa_tree_add_7_25_groupi_n_913);
  not csa_tree_add_7_25_groupi_drc_bufs23128(csa_tree_add_7_25_groupi_n_914 ,csa_tree_add_7_25_groupi_n_913);
  not csa_tree_add_7_25_groupi_drc_bufs23129(csa_tree_add_7_25_groupi_n_913 ,csa_tree_add_7_25_groupi_n_2279);
  not csa_tree_add_7_25_groupi_drc_bufs23131(csa_tree_add_7_25_groupi_n_912 ,csa_tree_add_7_25_groupi_n_910);
  not csa_tree_add_7_25_groupi_drc_bufs23132(csa_tree_add_7_25_groupi_n_911 ,csa_tree_add_7_25_groupi_n_910);
  not csa_tree_add_7_25_groupi_drc_bufs23133(csa_tree_add_7_25_groupi_n_910 ,csa_tree_add_7_25_groupi_n_2279);
  not csa_tree_add_7_25_groupi_drc_bufs23135(csa_tree_add_7_25_groupi_n_909 ,csa_tree_add_7_25_groupi_n_907);
  not csa_tree_add_7_25_groupi_drc_bufs23136(csa_tree_add_7_25_groupi_n_908 ,csa_tree_add_7_25_groupi_n_907);
  not csa_tree_add_7_25_groupi_drc_bufs23137(csa_tree_add_7_25_groupi_n_907 ,csa_tree_add_7_25_groupi_n_2292);
  not csa_tree_add_7_25_groupi_drc_bufs23139(csa_tree_add_7_25_groupi_n_906 ,csa_tree_add_7_25_groupi_n_904);
  not csa_tree_add_7_25_groupi_drc_bufs23140(csa_tree_add_7_25_groupi_n_905 ,csa_tree_add_7_25_groupi_n_904);
  not csa_tree_add_7_25_groupi_drc_bufs23141(csa_tree_add_7_25_groupi_n_904 ,csa_tree_add_7_25_groupi_n_2275);
  not csa_tree_add_7_25_groupi_drc_bufs23143(csa_tree_add_7_25_groupi_n_903 ,csa_tree_add_7_25_groupi_n_901);
  not csa_tree_add_7_25_groupi_drc_bufs23144(csa_tree_add_7_25_groupi_n_902 ,csa_tree_add_7_25_groupi_n_901);
  not csa_tree_add_7_25_groupi_drc_bufs23145(csa_tree_add_7_25_groupi_n_901 ,csa_tree_add_7_25_groupi_n_2275);
  not csa_tree_add_7_25_groupi_drc_bufs23147(csa_tree_add_7_25_groupi_n_900 ,csa_tree_add_7_25_groupi_n_898);
  not csa_tree_add_7_25_groupi_drc_bufs23148(csa_tree_add_7_25_groupi_n_899 ,csa_tree_add_7_25_groupi_n_898);
  not csa_tree_add_7_25_groupi_drc_bufs23149(csa_tree_add_7_25_groupi_n_898 ,csa_tree_add_7_25_groupi_n_2262);
  not csa_tree_add_7_25_groupi_drc_bufs23151(csa_tree_add_7_25_groupi_n_897 ,csa_tree_add_7_25_groupi_n_895);
  not csa_tree_add_7_25_groupi_drc_bufs23152(csa_tree_add_7_25_groupi_n_896 ,csa_tree_add_7_25_groupi_n_895);
  not csa_tree_add_7_25_groupi_drc_bufs23153(csa_tree_add_7_25_groupi_n_895 ,csa_tree_add_7_25_groupi_n_2299);
  not csa_tree_add_7_25_groupi_drc_bufs23155(csa_tree_add_7_25_groupi_n_894 ,csa_tree_add_7_25_groupi_n_892);
  not csa_tree_add_7_25_groupi_drc_bufs23156(csa_tree_add_7_25_groupi_n_893 ,csa_tree_add_7_25_groupi_n_892);
  not csa_tree_add_7_25_groupi_drc_bufs23157(csa_tree_add_7_25_groupi_n_892 ,csa_tree_add_7_25_groupi_n_2299);
  not csa_tree_add_7_25_groupi_drc_bufs23159(csa_tree_add_7_25_groupi_n_891 ,csa_tree_add_7_25_groupi_n_889);
  not csa_tree_add_7_25_groupi_drc_bufs23160(csa_tree_add_7_25_groupi_n_890 ,csa_tree_add_7_25_groupi_n_889);
  not csa_tree_add_7_25_groupi_drc_bufs23161(csa_tree_add_7_25_groupi_n_889 ,csa_tree_add_7_25_groupi_n_2269);
  not csa_tree_add_7_25_groupi_drc_bufs23163(csa_tree_add_7_25_groupi_n_888 ,csa_tree_add_7_25_groupi_n_886);
  not csa_tree_add_7_25_groupi_drc_bufs23164(csa_tree_add_7_25_groupi_n_887 ,csa_tree_add_7_25_groupi_n_886);
  not csa_tree_add_7_25_groupi_drc_bufs23165(csa_tree_add_7_25_groupi_n_886 ,csa_tree_add_7_25_groupi_n_2271);
  not csa_tree_add_7_25_groupi_drc_bufs23167(csa_tree_add_7_25_groupi_n_885 ,csa_tree_add_7_25_groupi_n_883);
  not csa_tree_add_7_25_groupi_drc_bufs23168(csa_tree_add_7_25_groupi_n_884 ,csa_tree_add_7_25_groupi_n_883);
  not csa_tree_add_7_25_groupi_drc_bufs23169(csa_tree_add_7_25_groupi_n_883 ,csa_tree_add_7_25_groupi_n_2271);
  not csa_tree_add_7_25_groupi_drc_bufs23171(csa_tree_add_7_25_groupi_n_882 ,csa_tree_add_7_25_groupi_n_880);
  not csa_tree_add_7_25_groupi_drc_bufs23172(csa_tree_add_7_25_groupi_n_881 ,csa_tree_add_7_25_groupi_n_880);
  not csa_tree_add_7_25_groupi_drc_bufs23173(csa_tree_add_7_25_groupi_n_880 ,csa_tree_add_7_25_groupi_n_2294);
  not csa_tree_add_7_25_groupi_drc_bufs23175(csa_tree_add_7_25_groupi_n_879 ,csa_tree_add_7_25_groupi_n_877);
  not csa_tree_add_7_25_groupi_drc_bufs23176(csa_tree_add_7_25_groupi_n_878 ,csa_tree_add_7_25_groupi_n_877);
  not csa_tree_add_7_25_groupi_drc_bufs23177(csa_tree_add_7_25_groupi_n_877 ,csa_tree_add_7_25_groupi_n_2259);
  not csa_tree_add_7_25_groupi_drc_bufs23179(csa_tree_add_7_25_groupi_n_876 ,csa_tree_add_7_25_groupi_n_874);
  not csa_tree_add_7_25_groupi_drc_bufs23180(csa_tree_add_7_25_groupi_n_875 ,csa_tree_add_7_25_groupi_n_874);
  not csa_tree_add_7_25_groupi_drc_bufs23181(csa_tree_add_7_25_groupi_n_874 ,csa_tree_add_7_25_groupi_n_2289);
  not csa_tree_add_7_25_groupi_drc_bufs23183(csa_tree_add_7_25_groupi_n_873 ,csa_tree_add_7_25_groupi_n_871);
  not csa_tree_add_7_25_groupi_drc_bufs23184(csa_tree_add_7_25_groupi_n_872 ,csa_tree_add_7_25_groupi_n_871);
  not csa_tree_add_7_25_groupi_drc_bufs23185(csa_tree_add_7_25_groupi_n_871 ,csa_tree_add_7_25_groupi_n_2291);
  not csa_tree_add_7_25_groupi_drc_bufs23187(csa_tree_add_7_25_groupi_n_870 ,csa_tree_add_7_25_groupi_n_868);
  not csa_tree_add_7_25_groupi_drc_bufs23188(csa_tree_add_7_25_groupi_n_869 ,csa_tree_add_7_25_groupi_n_868);
  not csa_tree_add_7_25_groupi_drc_bufs23189(csa_tree_add_7_25_groupi_n_868 ,csa_tree_add_7_25_groupi_n_2291);
  not csa_tree_add_7_25_groupi_drc_bufs23191(csa_tree_add_7_25_groupi_n_867 ,csa_tree_add_7_25_groupi_n_865);
  not csa_tree_add_7_25_groupi_drc_bufs23192(csa_tree_add_7_25_groupi_n_866 ,csa_tree_add_7_25_groupi_n_865);
  not csa_tree_add_7_25_groupi_drc_bufs23193(csa_tree_add_7_25_groupi_n_865 ,csa_tree_add_7_25_groupi_n_2258);
  not csa_tree_add_7_25_groupi_drc_bufs23195(csa_tree_add_7_25_groupi_n_864 ,csa_tree_add_7_25_groupi_n_862);
  not csa_tree_add_7_25_groupi_drc_bufs23196(csa_tree_add_7_25_groupi_n_863 ,csa_tree_add_7_25_groupi_n_862);
  not csa_tree_add_7_25_groupi_drc_bufs23197(csa_tree_add_7_25_groupi_n_862 ,csa_tree_add_7_25_groupi_n_2253);
  not csa_tree_add_7_25_groupi_drc_bufs23199(csa_tree_add_7_25_groupi_n_861 ,csa_tree_add_7_25_groupi_n_859);
  not csa_tree_add_7_25_groupi_drc_bufs23200(csa_tree_add_7_25_groupi_n_860 ,csa_tree_add_7_25_groupi_n_859);
  not csa_tree_add_7_25_groupi_drc_bufs23201(csa_tree_add_7_25_groupi_n_859 ,csa_tree_add_7_25_groupi_n_2297);
  not csa_tree_add_7_25_groupi_drc_bufs23203(csa_tree_add_7_25_groupi_n_858 ,csa_tree_add_7_25_groupi_n_856);
  not csa_tree_add_7_25_groupi_drc_bufs23204(csa_tree_add_7_25_groupi_n_857 ,csa_tree_add_7_25_groupi_n_856);
  not csa_tree_add_7_25_groupi_drc_bufs23205(csa_tree_add_7_25_groupi_n_856 ,csa_tree_add_7_25_groupi_n_2306);
  not csa_tree_add_7_25_groupi_drc_bufs23207(csa_tree_add_7_25_groupi_n_855 ,csa_tree_add_7_25_groupi_n_853);
  not csa_tree_add_7_25_groupi_drc_bufs23208(csa_tree_add_7_25_groupi_n_854 ,csa_tree_add_7_25_groupi_n_853);
  not csa_tree_add_7_25_groupi_drc_bufs23209(csa_tree_add_7_25_groupi_n_853 ,csa_tree_add_7_25_groupi_n_2290);
  not csa_tree_add_7_25_groupi_drc_bufs23211(csa_tree_add_7_25_groupi_n_852 ,csa_tree_add_7_25_groupi_n_850);
  not csa_tree_add_7_25_groupi_drc_bufs23212(csa_tree_add_7_25_groupi_n_851 ,csa_tree_add_7_25_groupi_n_850);
  not csa_tree_add_7_25_groupi_drc_bufs23213(csa_tree_add_7_25_groupi_n_850 ,csa_tree_add_7_25_groupi_n_2246);
  not csa_tree_add_7_25_groupi_drc_bufs23215(csa_tree_add_7_25_groupi_n_849 ,csa_tree_add_7_25_groupi_n_847);
  not csa_tree_add_7_25_groupi_drc_bufs23216(csa_tree_add_7_25_groupi_n_848 ,csa_tree_add_7_25_groupi_n_847);
  not csa_tree_add_7_25_groupi_drc_bufs23217(csa_tree_add_7_25_groupi_n_847 ,csa_tree_add_7_25_groupi_n_2288);
  not csa_tree_add_7_25_groupi_drc_bufs23219(csa_tree_add_7_25_groupi_n_846 ,csa_tree_add_7_25_groupi_n_844);
  not csa_tree_add_7_25_groupi_drc_bufs23220(csa_tree_add_7_25_groupi_n_845 ,csa_tree_add_7_25_groupi_n_844);
  not csa_tree_add_7_25_groupi_drc_bufs23221(csa_tree_add_7_25_groupi_n_844 ,csa_tree_add_7_25_groupi_n_2244);
  not csa_tree_add_7_25_groupi_drc_bufs23223(csa_tree_add_7_25_groupi_n_843 ,csa_tree_add_7_25_groupi_n_841);
  not csa_tree_add_7_25_groupi_drc_bufs23224(csa_tree_add_7_25_groupi_n_842 ,csa_tree_add_7_25_groupi_n_841);
  not csa_tree_add_7_25_groupi_drc_bufs23225(csa_tree_add_7_25_groupi_n_841 ,csa_tree_add_7_25_groupi_n_2286);
  not csa_tree_add_7_25_groupi_drc_bufs23227(csa_tree_add_7_25_groupi_n_840 ,csa_tree_add_7_25_groupi_n_838);
  not csa_tree_add_7_25_groupi_drc_bufs23228(csa_tree_add_7_25_groupi_n_839 ,csa_tree_add_7_25_groupi_n_838);
  not csa_tree_add_7_25_groupi_drc_bufs23229(csa_tree_add_7_25_groupi_n_838 ,csa_tree_add_7_25_groupi_n_2241);
  not csa_tree_add_7_25_groupi_drc_bufs23231(csa_tree_add_7_25_groupi_n_837 ,csa_tree_add_7_25_groupi_n_835);
  not csa_tree_add_7_25_groupi_drc_bufs23232(csa_tree_add_7_25_groupi_n_836 ,csa_tree_add_7_25_groupi_n_835);
  not csa_tree_add_7_25_groupi_drc_bufs23233(csa_tree_add_7_25_groupi_n_835 ,csa_tree_add_7_25_groupi_n_2268);
  not csa_tree_add_7_25_groupi_drc_bufs23235(csa_tree_add_7_25_groupi_n_834 ,csa_tree_add_7_25_groupi_n_832);
  not csa_tree_add_7_25_groupi_drc_bufs23236(csa_tree_add_7_25_groupi_n_833 ,csa_tree_add_7_25_groupi_n_832);
  not csa_tree_add_7_25_groupi_drc_bufs23237(csa_tree_add_7_25_groupi_n_832 ,csa_tree_add_7_25_groupi_n_2240);
  not csa_tree_add_7_25_groupi_drc_bufs23239(csa_tree_add_7_25_groupi_n_831 ,csa_tree_add_7_25_groupi_n_829);
  not csa_tree_add_7_25_groupi_drc_bufs23240(csa_tree_add_7_25_groupi_n_830 ,csa_tree_add_7_25_groupi_n_829);
  not csa_tree_add_7_25_groupi_drc_bufs23241(csa_tree_add_7_25_groupi_n_829 ,csa_tree_add_7_25_groupi_n_2250);
  not csa_tree_add_7_25_groupi_drc_bufs23243(csa_tree_add_7_25_groupi_n_828 ,csa_tree_add_7_25_groupi_n_826);
  not csa_tree_add_7_25_groupi_drc_bufs23244(csa_tree_add_7_25_groupi_n_827 ,csa_tree_add_7_25_groupi_n_826);
  not csa_tree_add_7_25_groupi_drc_bufs23245(csa_tree_add_7_25_groupi_n_826 ,csa_tree_add_7_25_groupi_n_2247);
  not csa_tree_add_7_25_groupi_drc_bufs23247(csa_tree_add_7_25_groupi_n_825 ,csa_tree_add_7_25_groupi_n_823);
  not csa_tree_add_7_25_groupi_drc_bufs23248(csa_tree_add_7_25_groupi_n_824 ,csa_tree_add_7_25_groupi_n_823);
  not csa_tree_add_7_25_groupi_drc_bufs23249(csa_tree_add_7_25_groupi_n_823 ,csa_tree_add_7_25_groupi_n_2312);
  not csa_tree_add_7_25_groupi_drc_bufs23251(csa_tree_add_7_25_groupi_n_822 ,csa_tree_add_7_25_groupi_n_820);
  not csa_tree_add_7_25_groupi_drc_bufs23252(csa_tree_add_7_25_groupi_n_821 ,csa_tree_add_7_25_groupi_n_820);
  not csa_tree_add_7_25_groupi_drc_bufs23253(csa_tree_add_7_25_groupi_n_820 ,csa_tree_add_7_25_groupi_n_2282);
  not csa_tree_add_7_25_groupi_drc_bufs23255(csa_tree_add_7_25_groupi_n_819 ,csa_tree_add_7_25_groupi_n_817);
  not csa_tree_add_7_25_groupi_drc_bufs23256(csa_tree_add_7_25_groupi_n_818 ,csa_tree_add_7_25_groupi_n_817);
  not csa_tree_add_7_25_groupi_drc_bufs23257(csa_tree_add_7_25_groupi_n_817 ,csa_tree_add_7_25_groupi_n_2313);
  not csa_tree_add_7_25_groupi_drc_bufs23259(csa_tree_add_7_25_groupi_n_816 ,csa_tree_add_7_25_groupi_n_814);
  not csa_tree_add_7_25_groupi_drc_bufs23260(csa_tree_add_7_25_groupi_n_815 ,csa_tree_add_7_25_groupi_n_814);
  not csa_tree_add_7_25_groupi_drc_bufs23261(csa_tree_add_7_25_groupi_n_814 ,csa_tree_add_7_25_groupi_n_2302);
  not csa_tree_add_7_25_groupi_drc_bufs23263(csa_tree_add_7_25_groupi_n_813 ,csa_tree_add_7_25_groupi_n_811);
  not csa_tree_add_7_25_groupi_drc_bufs23264(csa_tree_add_7_25_groupi_n_812 ,csa_tree_add_7_25_groupi_n_811);
  not csa_tree_add_7_25_groupi_drc_bufs23265(csa_tree_add_7_25_groupi_n_811 ,csa_tree_add_7_25_groupi_n_2305);
  not csa_tree_add_7_25_groupi_drc_bufs23267(csa_tree_add_7_25_groupi_n_810 ,csa_tree_add_7_25_groupi_n_808);
  not csa_tree_add_7_25_groupi_drc_bufs23268(csa_tree_add_7_25_groupi_n_809 ,csa_tree_add_7_25_groupi_n_808);
  not csa_tree_add_7_25_groupi_drc_bufs23269(csa_tree_add_7_25_groupi_n_808 ,csa_tree_add_7_25_groupi_n_2278);
  not csa_tree_add_7_25_groupi_drc_bufs23271(csa_tree_add_7_25_groupi_n_807 ,csa_tree_add_7_25_groupi_n_805);
  not csa_tree_add_7_25_groupi_drc_bufs23272(csa_tree_add_7_25_groupi_n_806 ,csa_tree_add_7_25_groupi_n_805);
  not csa_tree_add_7_25_groupi_drc_bufs23273(csa_tree_add_7_25_groupi_n_805 ,csa_tree_add_7_25_groupi_n_2293);
  not csa_tree_add_7_25_groupi_drc_bufs23275(csa_tree_add_7_25_groupi_n_804 ,csa_tree_add_7_25_groupi_n_802);
  not csa_tree_add_7_25_groupi_drc_bufs23276(csa_tree_add_7_25_groupi_n_803 ,csa_tree_add_7_25_groupi_n_802);
  not csa_tree_add_7_25_groupi_drc_bufs23277(csa_tree_add_7_25_groupi_n_802 ,csa_tree_add_7_25_groupi_n_2274);
  not csa_tree_add_7_25_groupi_drc_bufs23279(csa_tree_add_7_25_groupi_n_801 ,csa_tree_add_7_25_groupi_n_799);
  not csa_tree_add_7_25_groupi_drc_bufs23280(csa_tree_add_7_25_groupi_n_800 ,csa_tree_add_7_25_groupi_n_799);
  not csa_tree_add_7_25_groupi_drc_bufs23281(csa_tree_add_7_25_groupi_n_799 ,csa_tree_add_7_25_groupi_n_2304);
  not csa_tree_add_7_25_groupi_drc_bufs23283(csa_tree_add_7_25_groupi_n_798 ,csa_tree_add_7_25_groupi_n_796);
  not csa_tree_add_7_25_groupi_drc_bufs23284(csa_tree_add_7_25_groupi_n_797 ,csa_tree_add_7_25_groupi_n_796);
  not csa_tree_add_7_25_groupi_drc_bufs23285(csa_tree_add_7_25_groupi_n_796 ,csa_tree_add_7_25_groupi_n_2273);
  not csa_tree_add_7_25_groupi_drc_bufs23287(csa_tree_add_7_25_groupi_n_795 ,csa_tree_add_7_25_groupi_n_793);
  not csa_tree_add_7_25_groupi_drc_bufs23288(csa_tree_add_7_25_groupi_n_794 ,csa_tree_add_7_25_groupi_n_793);
  not csa_tree_add_7_25_groupi_drc_bufs23289(csa_tree_add_7_25_groupi_n_793 ,csa_tree_add_7_25_groupi_n_2242);
  not csa_tree_add_7_25_groupi_drc_bufs23291(csa_tree_add_7_25_groupi_n_792 ,csa_tree_add_7_25_groupi_n_790);
  not csa_tree_add_7_25_groupi_drc_bufs23292(csa_tree_add_7_25_groupi_n_791 ,csa_tree_add_7_25_groupi_n_790);
  not csa_tree_add_7_25_groupi_drc_bufs23293(csa_tree_add_7_25_groupi_n_790 ,csa_tree_add_7_25_groupi_n_2285);
  not csa_tree_add_7_25_groupi_drc_bufs23295(csa_tree_add_7_25_groupi_n_789 ,csa_tree_add_7_25_groupi_n_787);
  not csa_tree_add_7_25_groupi_drc_bufs23296(csa_tree_add_7_25_groupi_n_788 ,csa_tree_add_7_25_groupi_n_787);
  not csa_tree_add_7_25_groupi_drc_bufs23297(csa_tree_add_7_25_groupi_n_787 ,csa_tree_add_7_25_groupi_n_2239);
  not csa_tree_add_7_25_groupi_drc_bufs23299(csa_tree_add_7_25_groupi_n_786 ,csa_tree_add_7_25_groupi_n_784);
  not csa_tree_add_7_25_groupi_drc_bufs23300(csa_tree_add_7_25_groupi_n_785 ,csa_tree_add_7_25_groupi_n_784);
  not csa_tree_add_7_25_groupi_drc_bufs23301(csa_tree_add_7_25_groupi_n_784 ,csa_tree_add_7_25_groupi_n_2238);
  not csa_tree_add_7_25_groupi_drc_bufs23303(csa_tree_add_7_25_groupi_n_783 ,csa_tree_add_7_25_groupi_n_781);
  not csa_tree_add_7_25_groupi_drc_bufs23304(csa_tree_add_7_25_groupi_n_782 ,csa_tree_add_7_25_groupi_n_781);
  not csa_tree_add_7_25_groupi_drc_bufs23305(csa_tree_add_7_25_groupi_n_781 ,csa_tree_add_7_25_groupi_n_2265);
  not csa_tree_add_7_25_groupi_drc_bufs23307(csa_tree_add_7_25_groupi_n_780 ,csa_tree_add_7_25_groupi_n_778);
  not csa_tree_add_7_25_groupi_drc_bufs23308(csa_tree_add_7_25_groupi_n_779 ,csa_tree_add_7_25_groupi_n_778);
  not csa_tree_add_7_25_groupi_drc_bufs23309(csa_tree_add_7_25_groupi_n_778 ,csa_tree_add_7_25_groupi_n_2237);
  not csa_tree_add_7_25_groupi_drc_bufs23311(csa_tree_add_7_25_groupi_n_777 ,csa_tree_add_7_25_groupi_n_775);
  not csa_tree_add_7_25_groupi_drc_bufs23312(csa_tree_add_7_25_groupi_n_776 ,csa_tree_add_7_25_groupi_n_775);
  not csa_tree_add_7_25_groupi_drc_bufs23313(csa_tree_add_7_25_groupi_n_775 ,csa_tree_add_7_25_groupi_n_2284);
  not csa_tree_add_7_25_groupi_drc_bufs23315(csa_tree_add_7_25_groupi_n_774 ,csa_tree_add_7_25_groupi_n_772);
  not csa_tree_add_7_25_groupi_drc_bufs23316(csa_tree_add_7_25_groupi_n_773 ,csa_tree_add_7_25_groupi_n_772);
  not csa_tree_add_7_25_groupi_drc_bufs23317(csa_tree_add_7_25_groupi_n_772 ,csa_tree_add_7_25_groupi_n_2236);
  not csa_tree_add_7_25_groupi_drc_bufs23319(csa_tree_add_7_25_groupi_n_771 ,csa_tree_add_7_25_groupi_n_769);
  not csa_tree_add_7_25_groupi_drc_bufs23320(csa_tree_add_7_25_groupi_n_770 ,csa_tree_add_7_25_groupi_n_769);
  not csa_tree_add_7_25_groupi_drc_bufs23321(csa_tree_add_7_25_groupi_n_769 ,csa_tree_add_7_25_groupi_n_2235);
  not csa_tree_add_7_25_groupi_drc_bufs23323(csa_tree_add_7_25_groupi_n_768 ,csa_tree_add_7_25_groupi_n_766);
  not csa_tree_add_7_25_groupi_drc_bufs23324(csa_tree_add_7_25_groupi_n_767 ,csa_tree_add_7_25_groupi_n_766);
  not csa_tree_add_7_25_groupi_drc_bufs23325(csa_tree_add_7_25_groupi_n_766 ,csa_tree_add_7_25_groupi_n_2233);
  not csa_tree_add_7_25_groupi_drc_bufs23327(csa_tree_add_7_25_groupi_n_765 ,csa_tree_add_7_25_groupi_n_763);
  not csa_tree_add_7_25_groupi_drc_bufs23328(csa_tree_add_7_25_groupi_n_764 ,csa_tree_add_7_25_groupi_n_763);
  not csa_tree_add_7_25_groupi_drc_bufs23329(csa_tree_add_7_25_groupi_n_763 ,csa_tree_add_7_25_groupi_n_2232);
  not csa_tree_add_7_25_groupi_drc_bufs23331(csa_tree_add_7_25_groupi_n_762 ,csa_tree_add_7_25_groupi_n_760);
  not csa_tree_add_7_25_groupi_drc_bufs23332(csa_tree_add_7_25_groupi_n_761 ,csa_tree_add_7_25_groupi_n_760);
  not csa_tree_add_7_25_groupi_drc_bufs23333(csa_tree_add_7_25_groupi_n_760 ,csa_tree_add_7_25_groupi_n_2229);
  not csa_tree_add_7_25_groupi_drc_bufs23335(csa_tree_add_7_25_groupi_n_759 ,csa_tree_add_7_25_groupi_n_757);
  not csa_tree_add_7_25_groupi_drc_bufs23336(csa_tree_add_7_25_groupi_n_758 ,csa_tree_add_7_25_groupi_n_757);
  not csa_tree_add_7_25_groupi_drc_bufs23337(csa_tree_add_7_25_groupi_n_757 ,csa_tree_add_7_25_groupi_n_2281);
  not csa_tree_add_7_25_groupi_drc_bufs23339(csa_tree_add_7_25_groupi_n_756 ,csa_tree_add_7_25_groupi_n_754);
  not csa_tree_add_7_25_groupi_drc_bufs23340(csa_tree_add_7_25_groupi_n_755 ,csa_tree_add_7_25_groupi_n_754);
  not csa_tree_add_7_25_groupi_drc_bufs23341(csa_tree_add_7_25_groupi_n_754 ,csa_tree_add_7_25_groupi_n_2261);
  not csa_tree_add_7_25_groupi_drc_bufs23343(csa_tree_add_7_25_groupi_n_753 ,csa_tree_add_7_25_groupi_n_751);
  not csa_tree_add_7_25_groupi_drc_bufs23344(csa_tree_add_7_25_groupi_n_752 ,csa_tree_add_7_25_groupi_n_751);
  not csa_tree_add_7_25_groupi_drc_bufs23345(csa_tree_add_7_25_groupi_n_751 ,csa_tree_add_7_25_groupi_n_2280);
  not csa_tree_add_7_25_groupi_drc_bufs23347(csa_tree_add_7_25_groupi_n_750 ,csa_tree_add_7_25_groupi_n_748);
  not csa_tree_add_7_25_groupi_drc_bufs23348(csa_tree_add_7_25_groupi_n_749 ,csa_tree_add_7_25_groupi_n_748);
  not csa_tree_add_7_25_groupi_drc_bufs23349(csa_tree_add_7_25_groupi_n_748 ,csa_tree_add_7_25_groupi_n_2272);
  not csa_tree_add_7_25_groupi_drc_bufs23351(csa_tree_add_7_25_groupi_n_747 ,csa_tree_add_7_25_groupi_n_745);
  not csa_tree_add_7_25_groupi_drc_bufs23352(csa_tree_add_7_25_groupi_n_746 ,csa_tree_add_7_25_groupi_n_745);
  not csa_tree_add_7_25_groupi_drc_bufs23353(csa_tree_add_7_25_groupi_n_745 ,csa_tree_add_7_25_groupi_n_2301);
  not csa_tree_add_7_25_groupi_drc_bufs23355(csa_tree_add_7_25_groupi_n_744 ,csa_tree_add_7_25_groupi_n_742);
  not csa_tree_add_7_25_groupi_drc_bufs23356(csa_tree_add_7_25_groupi_n_743 ,csa_tree_add_7_25_groupi_n_742);
  not csa_tree_add_7_25_groupi_drc_bufs23357(csa_tree_add_7_25_groupi_n_742 ,csa_tree_add_7_25_groupi_n_2267);
  not csa_tree_add_7_25_groupi_drc_bufs23359(csa_tree_add_7_25_groupi_n_741 ,csa_tree_add_7_25_groupi_n_739);
  not csa_tree_add_7_25_groupi_drc_bufs23360(csa_tree_add_7_25_groupi_n_740 ,csa_tree_add_7_25_groupi_n_739);
  not csa_tree_add_7_25_groupi_drc_bufs23361(csa_tree_add_7_25_groupi_n_739 ,csa_tree_add_7_25_groupi_n_1938);
  not csa_tree_add_7_25_groupi_drc_bufs23363(csa_tree_add_7_25_groupi_n_738 ,csa_tree_add_7_25_groupi_n_736);
  not csa_tree_add_7_25_groupi_drc_bufs23364(csa_tree_add_7_25_groupi_n_737 ,csa_tree_add_7_25_groupi_n_736);
  not csa_tree_add_7_25_groupi_drc_bufs23365(csa_tree_add_7_25_groupi_n_736 ,csa_tree_add_7_25_groupi_n_2267);
  not csa_tree_add_7_25_groupi_drc_bufs23367(csa_tree_add_7_25_groupi_n_735 ,csa_tree_add_7_25_groupi_n_733);
  not csa_tree_add_7_25_groupi_drc_bufs23368(csa_tree_add_7_25_groupi_n_734 ,csa_tree_add_7_25_groupi_n_733);
  not csa_tree_add_7_25_groupi_drc_bufs23369(csa_tree_add_7_25_groupi_n_733 ,csa_tree_add_7_25_groupi_n_2311);
  not csa_tree_add_7_25_groupi_drc_bufs23371(csa_tree_add_7_25_groupi_n_732 ,csa_tree_add_7_25_groupi_n_730);
  not csa_tree_add_7_25_groupi_drc_bufs23372(csa_tree_add_7_25_groupi_n_731 ,csa_tree_add_7_25_groupi_n_730);
  not csa_tree_add_7_25_groupi_drc_bufs23373(csa_tree_add_7_25_groupi_n_730 ,csa_tree_add_7_25_groupi_n_2310);
  not csa_tree_add_7_25_groupi_drc_bufs23375(csa_tree_add_7_25_groupi_n_729 ,csa_tree_add_7_25_groupi_n_727);
  not csa_tree_add_7_25_groupi_drc_bufs23376(csa_tree_add_7_25_groupi_n_728 ,csa_tree_add_7_25_groupi_n_727);
  not csa_tree_add_7_25_groupi_drc_bufs23377(csa_tree_add_7_25_groupi_n_727 ,csa_tree_add_7_25_groupi_n_2310);
  not csa_tree_add_7_25_groupi_drc_bufs23379(csa_tree_add_7_25_groupi_n_726 ,csa_tree_add_7_25_groupi_n_724);
  not csa_tree_add_7_25_groupi_drc_bufs23380(csa_tree_add_7_25_groupi_n_725 ,csa_tree_add_7_25_groupi_n_724);
  not csa_tree_add_7_25_groupi_drc_bufs23381(csa_tree_add_7_25_groupi_n_724 ,csa_tree_add_7_25_groupi_n_2277);
  not csa_tree_add_7_25_groupi_drc_bufs23383(csa_tree_add_7_25_groupi_n_723 ,csa_tree_add_7_25_groupi_n_721);
  not csa_tree_add_7_25_groupi_drc_bufs23384(csa_tree_add_7_25_groupi_n_722 ,csa_tree_add_7_25_groupi_n_721);
  not csa_tree_add_7_25_groupi_drc_bufs23385(csa_tree_add_7_25_groupi_n_721 ,csa_tree_add_7_25_groupi_n_2295);
  not csa_tree_add_7_25_groupi_drc_bufs23387(csa_tree_add_7_25_groupi_n_720 ,csa_tree_add_7_25_groupi_n_718);
  not csa_tree_add_7_25_groupi_drc_bufs23388(csa_tree_add_7_25_groupi_n_719 ,csa_tree_add_7_25_groupi_n_718);
  not csa_tree_add_7_25_groupi_drc_bufs23389(csa_tree_add_7_25_groupi_n_718 ,csa_tree_add_7_25_groupi_n_2295);
  not csa_tree_add_7_25_groupi_drc_bufs23391(csa_tree_add_7_25_groupi_n_717 ,csa_tree_add_7_25_groupi_n_715);
  not csa_tree_add_7_25_groupi_drc_bufs23392(csa_tree_add_7_25_groupi_n_716 ,csa_tree_add_7_25_groupi_n_715);
  not csa_tree_add_7_25_groupi_drc_bufs23393(csa_tree_add_7_25_groupi_n_715 ,csa_tree_add_7_25_groupi_n_2309);
  not csa_tree_add_7_25_groupi_drc_bufs23395(csa_tree_add_7_25_groupi_n_714 ,csa_tree_add_7_25_groupi_n_712);
  not csa_tree_add_7_25_groupi_drc_bufs23396(csa_tree_add_7_25_groupi_n_713 ,csa_tree_add_7_25_groupi_n_712);
  not csa_tree_add_7_25_groupi_drc_bufs23397(csa_tree_add_7_25_groupi_n_712 ,csa_tree_add_7_25_groupi_n_2264);
  not csa_tree_add_7_25_groupi_drc_bufs23399(csa_tree_add_7_25_groupi_n_711 ,csa_tree_add_7_25_groupi_n_709);
  not csa_tree_add_7_25_groupi_drc_bufs23400(csa_tree_add_7_25_groupi_n_710 ,csa_tree_add_7_25_groupi_n_709);
  not csa_tree_add_7_25_groupi_drc_bufs23401(csa_tree_add_7_25_groupi_n_709 ,csa_tree_add_7_25_groupi_n_2264);
  not csa_tree_add_7_25_groupi_drc_bufs23403(csa_tree_add_7_25_groupi_n_708 ,csa_tree_add_7_25_groupi_n_706);
  not csa_tree_add_7_25_groupi_drc_bufs23404(csa_tree_add_7_25_groupi_n_707 ,csa_tree_add_7_25_groupi_n_706);
  not csa_tree_add_7_25_groupi_drc_bufs23405(csa_tree_add_7_25_groupi_n_706 ,csa_tree_add_7_25_groupi_n_2300);
  not csa_tree_add_7_25_groupi_drc_bufs23407(csa_tree_add_7_25_groupi_n_705 ,csa_tree_add_7_25_groupi_n_703);
  not csa_tree_add_7_25_groupi_drc_bufs23408(csa_tree_add_7_25_groupi_n_704 ,csa_tree_add_7_25_groupi_n_703);
  not csa_tree_add_7_25_groupi_drc_bufs23409(csa_tree_add_7_25_groupi_n_703 ,csa_tree_add_7_25_groupi_n_2260);
  not csa_tree_add_7_25_groupi_drc_bufs23411(csa_tree_add_7_25_groupi_n_702 ,csa_tree_add_7_25_groupi_n_700);
  not csa_tree_add_7_25_groupi_drc_bufs23412(csa_tree_add_7_25_groupi_n_701 ,csa_tree_add_7_25_groupi_n_700);
  not csa_tree_add_7_25_groupi_drc_bufs23413(csa_tree_add_7_25_groupi_n_700 ,csa_tree_add_7_25_groupi_n_2260);
  not csa_tree_add_7_25_groupi_drc_bufs23415(csa_tree_add_7_25_groupi_n_699 ,csa_tree_add_7_25_groupi_n_697);
  not csa_tree_add_7_25_groupi_drc_bufs23416(csa_tree_add_7_25_groupi_n_698 ,csa_tree_add_7_25_groupi_n_697);
  not csa_tree_add_7_25_groupi_drc_bufs23417(csa_tree_add_7_25_groupi_n_697 ,csa_tree_add_7_25_groupi_n_2308);
  not csa_tree_add_7_25_groupi_drc_bufs23419(csa_tree_add_7_25_groupi_n_696 ,csa_tree_add_7_25_groupi_n_694);
  not csa_tree_add_7_25_groupi_drc_bufs23420(csa_tree_add_7_25_groupi_n_695 ,csa_tree_add_7_25_groupi_n_694);
  not csa_tree_add_7_25_groupi_drc_bufs23421(csa_tree_add_7_25_groupi_n_694 ,csa_tree_add_7_25_groupi_n_2252);
  not csa_tree_add_7_25_groupi_drc_bufs23423(csa_tree_add_7_25_groupi_n_693 ,csa_tree_add_7_25_groupi_n_691);
  not csa_tree_add_7_25_groupi_drc_bufs23424(csa_tree_add_7_25_groupi_n_692 ,csa_tree_add_7_25_groupi_n_691);
  not csa_tree_add_7_25_groupi_drc_bufs23425(csa_tree_add_7_25_groupi_n_691 ,csa_tree_add_7_25_groupi_n_2252);
  not csa_tree_add_7_25_groupi_drc_bufs23427(csa_tree_add_7_25_groupi_n_690 ,csa_tree_add_7_25_groupi_n_688);
  not csa_tree_add_7_25_groupi_drc_bufs23428(csa_tree_add_7_25_groupi_n_689 ,csa_tree_add_7_25_groupi_n_688);
  not csa_tree_add_7_25_groupi_drc_bufs23429(csa_tree_add_7_25_groupi_n_688 ,csa_tree_add_7_25_groupi_n_2276);
  not csa_tree_add_7_25_groupi_drc_bufs23431(csa_tree_add_7_25_groupi_n_687 ,csa_tree_add_7_25_groupi_n_685);
  not csa_tree_add_7_25_groupi_drc_bufs23432(csa_tree_add_7_25_groupi_n_686 ,csa_tree_add_7_25_groupi_n_685);
  not csa_tree_add_7_25_groupi_drc_bufs23433(csa_tree_add_7_25_groupi_n_685 ,csa_tree_add_7_25_groupi_n_2251);
  not csa_tree_add_7_25_groupi_drc_bufs23435(csa_tree_add_7_25_groupi_n_684 ,csa_tree_add_7_25_groupi_n_682);
  not csa_tree_add_7_25_groupi_drc_bufs23436(csa_tree_add_7_25_groupi_n_683 ,csa_tree_add_7_25_groupi_n_682);
  not csa_tree_add_7_25_groupi_drc_bufs23437(csa_tree_add_7_25_groupi_n_682 ,csa_tree_add_7_25_groupi_n_2251);
  not csa_tree_add_7_25_groupi_drc_bufs23439(csa_tree_add_7_25_groupi_n_681 ,csa_tree_add_7_25_groupi_n_679);
  not csa_tree_add_7_25_groupi_drc_bufs23440(csa_tree_add_7_25_groupi_n_680 ,csa_tree_add_7_25_groupi_n_679);
  not csa_tree_add_7_25_groupi_drc_bufs23441(csa_tree_add_7_25_groupi_n_679 ,csa_tree_add_7_25_groupi_n_2270);
  not csa_tree_add_7_25_groupi_drc_bufs23443(csa_tree_add_7_25_groupi_n_678 ,csa_tree_add_7_25_groupi_n_676);
  not csa_tree_add_7_25_groupi_drc_bufs23444(csa_tree_add_7_25_groupi_n_677 ,csa_tree_add_7_25_groupi_n_676);
  not csa_tree_add_7_25_groupi_drc_bufs23445(csa_tree_add_7_25_groupi_n_676 ,csa_tree_add_7_25_groupi_n_2287);
  not csa_tree_add_7_25_groupi_drc_bufs23447(csa_tree_add_7_25_groupi_n_675 ,csa_tree_add_7_25_groupi_n_673);
  not csa_tree_add_7_25_groupi_drc_bufs23448(csa_tree_add_7_25_groupi_n_674 ,csa_tree_add_7_25_groupi_n_673);
  not csa_tree_add_7_25_groupi_drc_bufs23449(csa_tree_add_7_25_groupi_n_673 ,csa_tree_add_7_25_groupi_n_2287);
  not csa_tree_add_7_25_groupi_drc_bufs23451(csa_tree_add_7_25_groupi_n_672 ,csa_tree_add_7_25_groupi_n_670);
  not csa_tree_add_7_25_groupi_drc_bufs23452(csa_tree_add_7_25_groupi_n_671 ,csa_tree_add_7_25_groupi_n_670);
  not csa_tree_add_7_25_groupi_drc_bufs23453(csa_tree_add_7_25_groupi_n_670 ,csa_tree_add_7_25_groupi_n_2296);
  not csa_tree_add_7_25_groupi_drc_bufs23455(csa_tree_add_7_25_groupi_n_669 ,csa_tree_add_7_25_groupi_n_667);
  not csa_tree_add_7_25_groupi_drc_bufs23456(csa_tree_add_7_25_groupi_n_668 ,csa_tree_add_7_25_groupi_n_667);
  not csa_tree_add_7_25_groupi_drc_bufs23457(csa_tree_add_7_25_groupi_n_667 ,csa_tree_add_7_25_groupi_n_2249);
  not csa_tree_add_7_25_groupi_drc_bufs23459(csa_tree_add_7_25_groupi_n_666 ,csa_tree_add_7_25_groupi_n_664);
  not csa_tree_add_7_25_groupi_drc_bufs23460(csa_tree_add_7_25_groupi_n_665 ,csa_tree_add_7_25_groupi_n_664);
  not csa_tree_add_7_25_groupi_drc_bufs23461(csa_tree_add_7_25_groupi_n_664 ,csa_tree_add_7_25_groupi_n_2249);
  not csa_tree_add_7_25_groupi_drc_bufs23463(csa_tree_add_7_25_groupi_n_663 ,csa_tree_add_7_25_groupi_n_661);
  not csa_tree_add_7_25_groupi_drc_bufs23464(csa_tree_add_7_25_groupi_n_662 ,csa_tree_add_7_25_groupi_n_661);
  not csa_tree_add_7_25_groupi_drc_bufs23465(csa_tree_add_7_25_groupi_n_661 ,csa_tree_add_7_25_groupi_n_2298);
  not csa_tree_add_7_25_groupi_drc_bufs23467(csa_tree_add_7_25_groupi_n_660 ,csa_tree_add_7_25_groupi_n_658);
  not csa_tree_add_7_25_groupi_drc_bufs23468(csa_tree_add_7_25_groupi_n_659 ,csa_tree_add_7_25_groupi_n_658);
  not csa_tree_add_7_25_groupi_drc_bufs23469(csa_tree_add_7_25_groupi_n_658 ,csa_tree_add_7_25_groupi_n_2248);
  not csa_tree_add_7_25_groupi_drc_bufs23471(csa_tree_add_7_25_groupi_n_657 ,csa_tree_add_7_25_groupi_n_655);
  not csa_tree_add_7_25_groupi_drc_bufs23472(csa_tree_add_7_25_groupi_n_656 ,csa_tree_add_7_25_groupi_n_655);
  not csa_tree_add_7_25_groupi_drc_bufs23473(csa_tree_add_7_25_groupi_n_655 ,csa_tree_add_7_25_groupi_n_2248);
  not csa_tree_add_7_25_groupi_drc_bufs23475(csa_tree_add_7_25_groupi_n_654 ,csa_tree_add_7_25_groupi_n_652);
  not csa_tree_add_7_25_groupi_drc_bufs23476(csa_tree_add_7_25_groupi_n_653 ,csa_tree_add_7_25_groupi_n_652);
  not csa_tree_add_7_25_groupi_drc_bufs23477(csa_tree_add_7_25_groupi_n_652 ,csa_tree_add_7_25_groupi_n_2307);
  not csa_tree_add_7_25_groupi_drc_bufs23479(csa_tree_add_7_25_groupi_n_651 ,csa_tree_add_7_25_groupi_n_649);
  not csa_tree_add_7_25_groupi_drc_bufs23480(csa_tree_add_7_25_groupi_n_650 ,csa_tree_add_7_25_groupi_n_649);
  not csa_tree_add_7_25_groupi_drc_bufs23481(csa_tree_add_7_25_groupi_n_649 ,csa_tree_add_7_25_groupi_n_2245);
  not csa_tree_add_7_25_groupi_drc_bufs23483(csa_tree_add_7_25_groupi_n_648 ,csa_tree_add_7_25_groupi_n_646);
  not csa_tree_add_7_25_groupi_drc_bufs23484(csa_tree_add_7_25_groupi_n_647 ,csa_tree_add_7_25_groupi_n_646);
  not csa_tree_add_7_25_groupi_drc_bufs23485(csa_tree_add_7_25_groupi_n_646 ,csa_tree_add_7_25_groupi_n_2245);
  not csa_tree_add_7_25_groupi_drc_bufs23487(csa_tree_add_7_25_groupi_n_645 ,csa_tree_add_7_25_groupi_n_643);
  not csa_tree_add_7_25_groupi_drc_bufs23488(csa_tree_add_7_25_groupi_n_644 ,csa_tree_add_7_25_groupi_n_643);
  not csa_tree_add_7_25_groupi_drc_bufs23489(csa_tree_add_7_25_groupi_n_643 ,csa_tree_add_7_25_groupi_n_1946);
  not csa_tree_add_7_25_groupi_drc_bufs23491(csa_tree_add_7_25_groupi_n_642 ,csa_tree_add_7_25_groupi_n_640);
  not csa_tree_add_7_25_groupi_drc_bufs23492(csa_tree_add_7_25_groupi_n_641 ,csa_tree_add_7_25_groupi_n_640);
  not csa_tree_add_7_25_groupi_drc_bufs23493(csa_tree_add_7_25_groupi_n_640 ,csa_tree_add_7_25_groupi_n_1946);
  not csa_tree_add_7_25_groupi_drc_bufs23495(csa_tree_add_7_25_groupi_n_639 ,csa_tree_add_7_25_groupi_n_637);
  not csa_tree_add_7_25_groupi_drc_bufs23496(csa_tree_add_7_25_groupi_n_638 ,csa_tree_add_7_25_groupi_n_637);
  not csa_tree_add_7_25_groupi_drc_bufs23497(csa_tree_add_7_25_groupi_n_637 ,csa_tree_add_7_25_groupi_n_2888);
  not csa_tree_add_7_25_groupi_drc_bufs23499(csa_tree_add_7_25_groupi_n_636 ,csa_tree_add_7_25_groupi_n_634);
  not csa_tree_add_7_25_groupi_drc_bufs23500(csa_tree_add_7_25_groupi_n_635 ,csa_tree_add_7_25_groupi_n_634);
  not csa_tree_add_7_25_groupi_drc_bufs23501(csa_tree_add_7_25_groupi_n_634 ,csa_tree_add_7_25_groupi_n_1944);
  not csa_tree_add_7_25_groupi_drc_bufs23503(csa_tree_add_7_25_groupi_n_633 ,csa_tree_add_7_25_groupi_n_631);
  not csa_tree_add_7_25_groupi_drc_bufs23504(csa_tree_add_7_25_groupi_n_632 ,csa_tree_add_7_25_groupi_n_631);
  not csa_tree_add_7_25_groupi_drc_bufs23505(csa_tree_add_7_25_groupi_n_631 ,csa_tree_add_7_25_groupi_n_1954);
  not csa_tree_add_7_25_groupi_drc_bufs23507(csa_tree_add_7_25_groupi_n_630 ,csa_tree_add_7_25_groupi_n_628);
  not csa_tree_add_7_25_groupi_drc_bufs23508(csa_tree_add_7_25_groupi_n_629 ,csa_tree_add_7_25_groupi_n_628);
  not csa_tree_add_7_25_groupi_drc_bufs23509(csa_tree_add_7_25_groupi_n_628 ,csa_tree_add_7_25_groupi_n_2367);
  not csa_tree_add_7_25_groupi_drc_bufs23511(csa_tree_add_7_25_groupi_n_627 ,csa_tree_add_7_25_groupi_n_625);
  not csa_tree_add_7_25_groupi_drc_bufs23512(csa_tree_add_7_25_groupi_n_626 ,csa_tree_add_7_25_groupi_n_625);
  not csa_tree_add_7_25_groupi_drc_bufs23513(csa_tree_add_7_25_groupi_n_625 ,csa_tree_add_7_25_groupi_n_1951);
  not csa_tree_add_7_25_groupi_drc_bufs23515(csa_tree_add_7_25_groupi_n_624 ,csa_tree_add_7_25_groupi_n_622);
  not csa_tree_add_7_25_groupi_drc_bufs23516(csa_tree_add_7_25_groupi_n_623 ,csa_tree_add_7_25_groupi_n_622);
  not csa_tree_add_7_25_groupi_drc_bufs23517(csa_tree_add_7_25_groupi_n_622 ,csa_tree_add_7_25_groupi_n_2403);
  not csa_tree_add_7_25_groupi_drc_bufs23519(csa_tree_add_7_25_groupi_n_621 ,csa_tree_add_7_25_groupi_n_619);
  not csa_tree_add_7_25_groupi_drc_bufs23520(csa_tree_add_7_25_groupi_n_620 ,csa_tree_add_7_25_groupi_n_619);
  not csa_tree_add_7_25_groupi_drc_bufs23521(csa_tree_add_7_25_groupi_n_619 ,csa_tree_add_7_25_groupi_n_2259);
  not csa_tree_add_7_25_groupi_drc_bufs23523(csa_tree_add_7_25_groupi_n_618 ,csa_tree_add_7_25_groupi_n_616);
  not csa_tree_add_7_25_groupi_drc_bufs23524(csa_tree_add_7_25_groupi_n_617 ,csa_tree_add_7_25_groupi_n_616);
  not csa_tree_add_7_25_groupi_drc_bufs23525(csa_tree_add_7_25_groupi_n_616 ,csa_tree_add_7_25_groupi_n_2253);
  not csa_tree_add_7_25_groupi_drc_bufs23527(csa_tree_add_7_25_groupi_n_615 ,csa_tree_add_7_25_groupi_n_613);
  not csa_tree_add_7_25_groupi_drc_bufs23528(csa_tree_add_7_25_groupi_n_614 ,csa_tree_add_7_25_groupi_n_613);
  not csa_tree_add_7_25_groupi_drc_bufs23529(csa_tree_add_7_25_groupi_n_613 ,csa_tree_add_7_25_groupi_n_2306);
  not csa_tree_add_7_25_groupi_drc_bufs23531(csa_tree_add_7_25_groupi_n_612 ,csa_tree_add_7_25_groupi_n_610);
  not csa_tree_add_7_25_groupi_drc_bufs23532(csa_tree_add_7_25_groupi_n_611 ,csa_tree_add_7_25_groupi_n_610);
  not csa_tree_add_7_25_groupi_drc_bufs23533(csa_tree_add_7_25_groupi_n_610 ,csa_tree_add_7_25_groupi_n_2243);
  not csa_tree_add_7_25_groupi_drc_bufs23535(csa_tree_add_7_25_groupi_n_609 ,csa_tree_add_7_25_groupi_n_607);
  not csa_tree_add_7_25_groupi_drc_bufs23536(csa_tree_add_7_25_groupi_n_608 ,csa_tree_add_7_25_groupi_n_607);
  not csa_tree_add_7_25_groupi_drc_bufs23537(csa_tree_add_7_25_groupi_n_607 ,csa_tree_add_7_25_groupi_n_2246);
  not csa_tree_add_7_25_groupi_drc_bufs23539(csa_tree_add_7_25_groupi_n_606 ,csa_tree_add_7_25_groupi_n_604);
  not csa_tree_add_7_25_groupi_drc_bufs23540(csa_tree_add_7_25_groupi_n_605 ,csa_tree_add_7_25_groupi_n_604);
  not csa_tree_add_7_25_groupi_drc_bufs23541(csa_tree_add_7_25_groupi_n_604 ,csa_tree_add_7_25_groupi_n_2244);
  not csa_tree_add_7_25_groupi_drc_bufs23543(csa_tree_add_7_25_groupi_n_603 ,csa_tree_add_7_25_groupi_n_601);
  not csa_tree_add_7_25_groupi_drc_bufs23544(csa_tree_add_7_25_groupi_n_602 ,csa_tree_add_7_25_groupi_n_601);
  not csa_tree_add_7_25_groupi_drc_bufs23545(csa_tree_add_7_25_groupi_n_601 ,csa_tree_add_7_25_groupi_n_2241);
  not csa_tree_add_7_25_groupi_drc_bufs23547(csa_tree_add_7_25_groupi_n_600 ,csa_tree_add_7_25_groupi_n_598);
  not csa_tree_add_7_25_groupi_drc_bufs23548(csa_tree_add_7_25_groupi_n_599 ,csa_tree_add_7_25_groupi_n_598);
  not csa_tree_add_7_25_groupi_drc_bufs23549(csa_tree_add_7_25_groupi_n_598 ,csa_tree_add_7_25_groupi_n_2240);
  not csa_tree_add_7_25_groupi_drc_bufs23551(csa_tree_add_7_25_groupi_n_597 ,csa_tree_add_7_25_groupi_n_595);
  not csa_tree_add_7_25_groupi_drc_bufs23552(csa_tree_add_7_25_groupi_n_596 ,csa_tree_add_7_25_groupi_n_595);
  not csa_tree_add_7_25_groupi_drc_bufs23553(csa_tree_add_7_25_groupi_n_595 ,csa_tree_add_7_25_groupi_n_2247);
  not csa_tree_add_7_25_groupi_drc_bufs23555(csa_tree_add_7_25_groupi_n_594 ,csa_tree_add_7_25_groupi_n_592);
  not csa_tree_add_7_25_groupi_drc_bufs23556(csa_tree_add_7_25_groupi_n_593 ,csa_tree_add_7_25_groupi_n_592);
  not csa_tree_add_7_25_groupi_drc_bufs23557(csa_tree_add_7_25_groupi_n_592 ,csa_tree_add_7_25_groupi_n_2243);
  not csa_tree_add_7_25_groupi_drc_bufs23559(csa_tree_add_7_25_groupi_n_591 ,csa_tree_add_7_25_groupi_n_589);
  not csa_tree_add_7_25_groupi_drc_bufs23560(csa_tree_add_7_25_groupi_n_590 ,csa_tree_add_7_25_groupi_n_589);
  not csa_tree_add_7_25_groupi_drc_bufs23561(csa_tree_add_7_25_groupi_n_589 ,csa_tree_add_7_25_groupi_n_2234);
  not csa_tree_add_7_25_groupi_drc_bufs23563(csa_tree_add_7_25_groupi_n_588 ,csa_tree_add_7_25_groupi_n_586);
  not csa_tree_add_7_25_groupi_drc_bufs23564(csa_tree_add_7_25_groupi_n_587 ,csa_tree_add_7_25_groupi_n_586);
  not csa_tree_add_7_25_groupi_drc_bufs23565(csa_tree_add_7_25_groupi_n_586 ,csa_tree_add_7_25_groupi_n_2234);
  not csa_tree_add_7_25_groupi_drc_bufs23567(csa_tree_add_7_25_groupi_n_585 ,csa_tree_add_7_25_groupi_n_583);
  not csa_tree_add_7_25_groupi_drc_bufs23568(csa_tree_add_7_25_groupi_n_584 ,csa_tree_add_7_25_groupi_n_583);
  not csa_tree_add_7_25_groupi_drc_bufs23569(csa_tree_add_7_25_groupi_n_583 ,csa_tree_add_7_25_groupi_n_2255);
  not csa_tree_add_7_25_groupi_drc_bufs23571(csa_tree_add_7_25_groupi_n_582 ,csa_tree_add_7_25_groupi_n_580);
  not csa_tree_add_7_25_groupi_drc_bufs23572(csa_tree_add_7_25_groupi_n_581 ,csa_tree_add_7_25_groupi_n_580);
  not csa_tree_add_7_25_groupi_drc_bufs23573(csa_tree_add_7_25_groupi_n_580 ,csa_tree_add_7_25_groupi_n_2254);
  not csa_tree_add_7_25_groupi_drc_bufs23575(csa_tree_add_7_25_groupi_n_579 ,csa_tree_add_7_25_groupi_n_577);
  not csa_tree_add_7_25_groupi_drc_bufs23576(csa_tree_add_7_25_groupi_n_578 ,csa_tree_add_7_25_groupi_n_577);
  not csa_tree_add_7_25_groupi_drc_bufs23577(csa_tree_add_7_25_groupi_n_577 ,csa_tree_add_7_25_groupi_n_2257);
  not csa_tree_add_7_25_groupi_drc_bufs23579(csa_tree_add_7_25_groupi_n_576 ,csa_tree_add_7_25_groupi_n_574);
  not csa_tree_add_7_25_groupi_drc_bufs23580(csa_tree_add_7_25_groupi_n_575 ,csa_tree_add_7_25_groupi_n_574);
  not csa_tree_add_7_25_groupi_drc_bufs23581(csa_tree_add_7_25_groupi_n_574 ,csa_tree_add_7_25_groupi_n_2256);
  not csa_tree_add_7_25_groupi_drc_bufs23583(csa_tree_add_7_25_groupi_n_573 ,csa_tree_add_7_25_groupi_n_571);
  not csa_tree_add_7_25_groupi_drc_bufs23584(csa_tree_add_7_25_groupi_n_572 ,csa_tree_add_7_25_groupi_n_571);
  not csa_tree_add_7_25_groupi_drc_bufs23585(csa_tree_add_7_25_groupi_n_571 ,csa_tree_add_7_25_groupi_n_2231);
  not csa_tree_add_7_25_groupi_drc_bufs23587(csa_tree_add_7_25_groupi_n_570 ,csa_tree_add_7_25_groupi_n_568);
  not csa_tree_add_7_25_groupi_drc_bufs23588(csa_tree_add_7_25_groupi_n_569 ,csa_tree_add_7_25_groupi_n_568);
  not csa_tree_add_7_25_groupi_drc_bufs23589(csa_tree_add_7_25_groupi_n_568 ,csa_tree_add_7_25_groupi_n_2230);
  not csa_tree_add_7_25_groupi_drc_bufs23591(csa_tree_add_7_25_groupi_n_567 ,csa_tree_add_7_25_groupi_n_565);
  not csa_tree_add_7_25_groupi_drc_bufs23592(csa_tree_add_7_25_groupi_n_566 ,csa_tree_add_7_25_groupi_n_565);
  not csa_tree_add_7_25_groupi_drc_bufs23593(csa_tree_add_7_25_groupi_n_565 ,csa_tree_add_7_25_groupi_n_2228);
  not csa_tree_add_7_25_groupi_drc_bufs23595(csa_tree_add_7_25_groupi_n_564 ,csa_tree_add_7_25_groupi_n_562);
  not csa_tree_add_7_25_groupi_drc_bufs23596(csa_tree_add_7_25_groupi_n_563 ,csa_tree_add_7_25_groupi_n_562);
  not csa_tree_add_7_25_groupi_drc_bufs23597(csa_tree_add_7_25_groupi_n_562 ,csa_tree_add_7_25_groupi_n_2227);
  not csa_tree_add_7_25_groupi_drc_bufs23599(csa_tree_add_7_25_groupi_n_561 ,csa_tree_add_7_25_groupi_n_559);
  not csa_tree_add_7_25_groupi_drc_bufs23600(csa_tree_add_7_25_groupi_n_560 ,csa_tree_add_7_25_groupi_n_559);
  not csa_tree_add_7_25_groupi_drc_bufs23601(csa_tree_add_7_25_groupi_n_559 ,csa_tree_add_7_25_groupi_n_2225);
  not csa_tree_add_7_25_groupi_drc_bufs23603(csa_tree_add_7_25_groupi_n_558 ,csa_tree_add_7_25_groupi_n_556);
  not csa_tree_add_7_25_groupi_drc_bufs23604(csa_tree_add_7_25_groupi_n_557 ,csa_tree_add_7_25_groupi_n_556);
  not csa_tree_add_7_25_groupi_drc_bufs23605(csa_tree_add_7_25_groupi_n_556 ,csa_tree_add_7_25_groupi_n_2224);
  not csa_tree_add_7_25_groupi_drc_bufs23607(csa_tree_add_7_25_groupi_n_555 ,csa_tree_add_7_25_groupi_n_553);
  not csa_tree_add_7_25_groupi_drc_bufs23608(csa_tree_add_7_25_groupi_n_554 ,csa_tree_add_7_25_groupi_n_553);
  not csa_tree_add_7_25_groupi_drc_bufs23609(csa_tree_add_7_25_groupi_n_553 ,csa_tree_add_7_25_groupi_n_1935);
  not csa_tree_add_7_25_groupi_drc_bufs23611(csa_tree_add_7_25_groupi_n_552 ,csa_tree_add_7_25_groupi_n_550);
  not csa_tree_add_7_25_groupi_drc_bufs23612(csa_tree_add_7_25_groupi_n_551 ,csa_tree_add_7_25_groupi_n_550);
  not csa_tree_add_7_25_groupi_drc_bufs23613(csa_tree_add_7_25_groupi_n_550 ,csa_tree_add_7_25_groupi_n_2888);
  not csa_tree_add_7_25_groupi_drc_bufs23615(csa_tree_add_7_25_groupi_n_549 ,csa_tree_add_7_25_groupi_n_547);
  not csa_tree_add_7_25_groupi_drc_bufs23616(csa_tree_add_7_25_groupi_n_548 ,csa_tree_add_7_25_groupi_n_547);
  not csa_tree_add_7_25_groupi_drc_bufs23617(csa_tree_add_7_25_groupi_n_547 ,csa_tree_add_7_25_groupi_n_1944);
  not csa_tree_add_7_25_groupi_drc_bufs23619(csa_tree_add_7_25_groupi_n_546 ,csa_tree_add_7_25_groupi_n_544);
  not csa_tree_add_7_25_groupi_drc_bufs23620(csa_tree_add_7_25_groupi_n_545 ,csa_tree_add_7_25_groupi_n_544);
  not csa_tree_add_7_25_groupi_drc_bufs23621(csa_tree_add_7_25_groupi_n_544 ,csa_tree_add_7_25_groupi_n_2255);
  not csa_tree_add_7_25_groupi_drc_bufs23623(csa_tree_add_7_25_groupi_n_543 ,csa_tree_add_7_25_groupi_n_541);
  not csa_tree_add_7_25_groupi_drc_bufs23624(csa_tree_add_7_25_groupi_n_542 ,csa_tree_add_7_25_groupi_n_541);
  not csa_tree_add_7_25_groupi_drc_bufs23625(csa_tree_add_7_25_groupi_n_541 ,csa_tree_add_7_25_groupi_n_2254);
  not csa_tree_add_7_25_groupi_drc_bufs23627(csa_tree_add_7_25_groupi_n_540 ,csa_tree_add_7_25_groupi_n_538);
  not csa_tree_add_7_25_groupi_drc_bufs23628(csa_tree_add_7_25_groupi_n_539 ,csa_tree_add_7_25_groupi_n_538);
  not csa_tree_add_7_25_groupi_drc_bufs23629(csa_tree_add_7_25_groupi_n_538 ,csa_tree_add_7_25_groupi_n_2218);
  not csa_tree_add_7_25_groupi_drc_bufs23631(csa_tree_add_7_25_groupi_n_537 ,csa_tree_add_7_25_groupi_n_535);
  not csa_tree_add_7_25_groupi_drc_bufs23632(csa_tree_add_7_25_groupi_n_536 ,csa_tree_add_7_25_groupi_n_535);
  not csa_tree_add_7_25_groupi_drc_bufs23633(csa_tree_add_7_25_groupi_n_535 ,csa_tree_add_7_25_groupi_n_1942);
  not csa_tree_add_7_25_groupi_drc_bufs23635(csa_tree_add_7_25_groupi_n_534 ,csa_tree_add_7_25_groupi_n_532);
  not csa_tree_add_7_25_groupi_drc_bufs23636(csa_tree_add_7_25_groupi_n_533 ,csa_tree_add_7_25_groupi_n_532);
  not csa_tree_add_7_25_groupi_drc_bufs23637(csa_tree_add_7_25_groupi_n_532 ,csa_tree_add_7_25_groupi_n_1942);
  not csa_tree_add_7_25_groupi_drc_bufs23639(csa_tree_add_7_25_groupi_n_531 ,csa_tree_add_7_25_groupi_n_529);
  not csa_tree_add_7_25_groupi_drc_bufs23640(csa_tree_add_7_25_groupi_n_530 ,csa_tree_add_7_25_groupi_n_529);
  not csa_tree_add_7_25_groupi_drc_bufs23641(csa_tree_add_7_25_groupi_n_529 ,csa_tree_add_7_25_groupi_n_2887);
  not csa_tree_add_7_25_groupi_drc_bufs23643(csa_tree_add_7_25_groupi_n_528 ,csa_tree_add_7_25_groupi_n_526);
  not csa_tree_add_7_25_groupi_drc_bufs23644(csa_tree_add_7_25_groupi_n_527 ,csa_tree_add_7_25_groupi_n_526);
  not csa_tree_add_7_25_groupi_drc_bufs23645(csa_tree_add_7_25_groupi_n_526 ,csa_tree_add_7_25_groupi_n_3535);
  not csa_tree_add_7_25_groupi_drc_bufs23647(csa_tree_add_7_25_groupi_n_525 ,csa_tree_add_7_25_groupi_n_523);
  not csa_tree_add_7_25_groupi_drc_bufs23648(csa_tree_add_7_25_groupi_n_524 ,csa_tree_add_7_25_groupi_n_523);
  not csa_tree_add_7_25_groupi_drc_bufs23649(csa_tree_add_7_25_groupi_n_523 ,csa_tree_add_7_25_groupi_n_1932);
  not csa_tree_add_7_25_groupi_drc_bufs23651(csa_tree_add_7_25_groupi_n_522 ,csa_tree_add_7_25_groupi_n_520);
  not csa_tree_add_7_25_groupi_drc_bufs23652(csa_tree_add_7_25_groupi_n_521 ,csa_tree_add_7_25_groupi_n_520);
  not csa_tree_add_7_25_groupi_drc_bufs23653(csa_tree_add_7_25_groupi_n_520 ,csa_tree_add_7_25_groupi_n_1929);
  not csa_tree_add_7_25_groupi_drc_bufs23655(csa_tree_add_7_25_groupi_n_519 ,csa_tree_add_7_25_groupi_n_517);
  not csa_tree_add_7_25_groupi_drc_bufs23656(csa_tree_add_7_25_groupi_n_518 ,csa_tree_add_7_25_groupi_n_517);
  not csa_tree_add_7_25_groupi_drc_bufs23657(csa_tree_add_7_25_groupi_n_517 ,csa_tree_add_7_25_groupi_n_1926);
  not csa_tree_add_7_25_groupi_drc_bufs23659(csa_tree_add_7_25_groupi_n_516 ,csa_tree_add_7_25_groupi_n_514);
  not csa_tree_add_7_25_groupi_drc_bufs23660(csa_tree_add_7_25_groupi_n_515 ,csa_tree_add_7_25_groupi_n_514);
  not csa_tree_add_7_25_groupi_drc_bufs23661(csa_tree_add_7_25_groupi_n_514 ,csa_tree_add_7_25_groupi_n_1948);
  not csa_tree_add_7_25_groupi_drc_bufs23663(csa_tree_add_7_25_groupi_n_513 ,csa_tree_add_7_25_groupi_n_511);
  not csa_tree_add_7_25_groupi_drc_bufs23664(csa_tree_add_7_25_groupi_n_512 ,csa_tree_add_7_25_groupi_n_511);
  not csa_tree_add_7_25_groupi_drc_bufs23665(csa_tree_add_7_25_groupi_n_511 ,csa_tree_add_7_25_groupi_n_2803);
  not csa_tree_add_7_25_groupi_drc_bufs23667(csa_tree_add_7_25_groupi_n_510 ,csa_tree_add_7_25_groupi_n_508);
  not csa_tree_add_7_25_groupi_drc_bufs23668(csa_tree_add_7_25_groupi_n_509 ,csa_tree_add_7_25_groupi_n_508);
  not csa_tree_add_7_25_groupi_drc_bufs23669(csa_tree_add_7_25_groupi_n_508 ,csa_tree_add_7_25_groupi_n_2803);
  not csa_tree_add_7_25_groupi_drc_bufs23671(csa_tree_add_7_25_groupi_n_507 ,csa_tree_add_7_25_groupi_n_505);
  not csa_tree_add_7_25_groupi_drc_bufs23672(csa_tree_add_7_25_groupi_n_506 ,csa_tree_add_7_25_groupi_n_505);
  not csa_tree_add_7_25_groupi_drc_bufs23673(csa_tree_add_7_25_groupi_n_505 ,csa_tree_add_7_25_groupi_n_1923);
  not csa_tree_add_7_25_groupi_drc_bufs23675(csa_tree_add_7_25_groupi_n_504 ,csa_tree_add_7_25_groupi_n_502);
  not csa_tree_add_7_25_groupi_drc_bufs23676(csa_tree_add_7_25_groupi_n_503 ,csa_tree_add_7_25_groupi_n_502);
  not csa_tree_add_7_25_groupi_drc_bufs23677(csa_tree_add_7_25_groupi_n_502 ,csa_tree_add_7_25_groupi_n_2889);
  not csa_tree_add_7_25_groupi_drc_bufs23679(csa_tree_add_7_25_groupi_n_501 ,csa_tree_add_7_25_groupi_n_499);
  not csa_tree_add_7_25_groupi_drc_bufs23680(csa_tree_add_7_25_groupi_n_500 ,csa_tree_add_7_25_groupi_n_499);
  not csa_tree_add_7_25_groupi_drc_bufs23681(csa_tree_add_7_25_groupi_n_499 ,csa_tree_add_7_25_groupi_n_1940);
  not csa_tree_add_7_25_groupi_drc_bufs23683(csa_tree_add_7_25_groupi_n_498 ,csa_tree_add_7_25_groupi_n_496);
  not csa_tree_add_7_25_groupi_drc_bufs23684(csa_tree_add_7_25_groupi_n_497 ,csa_tree_add_7_25_groupi_n_496);
  not csa_tree_add_7_25_groupi_drc_bufs23685(csa_tree_add_7_25_groupi_n_496 ,csa_tree_add_7_25_groupi_n_2889);
  not csa_tree_add_7_25_groupi_drc_bufs23687(csa_tree_add_7_25_groupi_n_495 ,csa_tree_add_7_25_groupi_n_493);
  not csa_tree_add_7_25_groupi_drc_bufs23688(csa_tree_add_7_25_groupi_n_494 ,csa_tree_add_7_25_groupi_n_493);
  not csa_tree_add_7_25_groupi_drc_bufs23689(csa_tree_add_7_25_groupi_n_493 ,csa_tree_add_7_25_groupi_n_1940);
  not csa_tree_add_7_25_groupi_drc_bufs23691(csa_tree_add_7_25_groupi_n_492 ,csa_tree_add_7_25_groupi_n_490);
  not csa_tree_add_7_25_groupi_drc_bufs23692(csa_tree_add_7_25_groupi_n_491 ,csa_tree_add_7_25_groupi_n_490);
  not csa_tree_add_7_25_groupi_drc_bufs23693(csa_tree_add_7_25_groupi_n_490 ,csa_tree_add_7_25_groupi_n_2687);
  not csa_tree_add_7_25_groupi_drc_bufs23695(csa_tree_add_7_25_groupi_n_489 ,csa_tree_add_7_25_groupi_n_487);
  not csa_tree_add_7_25_groupi_drc_bufs23696(csa_tree_add_7_25_groupi_n_488 ,csa_tree_add_7_25_groupi_n_487);
  not csa_tree_add_7_25_groupi_drc_bufs23697(csa_tree_add_7_25_groupi_n_487 ,csa_tree_add_7_25_groupi_n_1920);
  not csa_tree_add_7_25_groupi_drc_bufs23699(csa_tree_add_7_25_groupi_n_486 ,csa_tree_add_7_25_groupi_n_484);
  not csa_tree_add_7_25_groupi_drc_bufs23700(csa_tree_add_7_25_groupi_n_485 ,csa_tree_add_7_25_groupi_n_484);
  not csa_tree_add_7_25_groupi_drc_bufs23701(csa_tree_add_7_25_groupi_n_484 ,csa_tree_add_7_25_groupi_n_2208);
  not csa_tree_add_7_25_groupi_drc_bufs23703(csa_tree_add_7_25_groupi_n_483 ,csa_tree_add_7_25_groupi_n_482);
  not csa_tree_add_7_25_groupi_drc_bufs23705(csa_tree_add_7_25_groupi_n_482 ,csa_tree_add_7_25_groupi_n_1917);
  not csa_tree_add_7_25_groupi_drc_bufs23707(csa_tree_add_7_25_groupi_n_481 ,csa_tree_add_7_25_groupi_n_479);
  not csa_tree_add_7_25_groupi_drc_bufs23708(csa_tree_add_7_25_groupi_n_480 ,csa_tree_add_7_25_groupi_n_479);
  not csa_tree_add_7_25_groupi_drc_bufs23709(csa_tree_add_7_25_groupi_n_479 ,csa_tree_add_7_25_groupi_n_2200);
  not csa_tree_add_7_25_groupi_drc_bufs23711(csa_tree_add_7_25_groupi_n_478 ,csa_tree_add_7_25_groupi_n_476);
  not csa_tree_add_7_25_groupi_drc_bufs23712(csa_tree_add_7_25_groupi_n_477 ,csa_tree_add_7_25_groupi_n_476);
  not csa_tree_add_7_25_groupi_drc_bufs23713(csa_tree_add_7_25_groupi_n_476 ,csa_tree_add_7_25_groupi_n_2204);
  not csa_tree_add_7_25_groupi_drc_bufs23715(csa_tree_add_7_25_groupi_n_475 ,csa_tree_add_7_25_groupi_n_473);
  not csa_tree_add_7_25_groupi_drc_bufs23716(csa_tree_add_7_25_groupi_n_474 ,csa_tree_add_7_25_groupi_n_473);
  not csa_tree_add_7_25_groupi_drc_bufs23717(csa_tree_add_7_25_groupi_n_473 ,csa_tree_add_7_25_groupi_n_2237);
  not csa_tree_add_7_25_groupi_drc_bufs23719(csa_tree_add_7_25_groupi_n_472 ,csa_tree_add_7_25_groupi_n_470);
  not csa_tree_add_7_25_groupi_drc_bufs23720(csa_tree_add_7_25_groupi_n_471 ,csa_tree_add_7_25_groupi_n_470);
  not csa_tree_add_7_25_groupi_drc_bufs23721(csa_tree_add_7_25_groupi_n_470 ,csa_tree_add_7_25_groupi_n_2235);
  not csa_tree_add_7_25_groupi_drc_bufs23723(csa_tree_add_7_25_groupi_n_469 ,csa_tree_add_7_25_groupi_n_467);
  not csa_tree_add_7_25_groupi_drc_bufs23724(csa_tree_add_7_25_groupi_n_468 ,csa_tree_add_7_25_groupi_n_467);
  not csa_tree_add_7_25_groupi_drc_bufs23725(csa_tree_add_7_25_groupi_n_467 ,csa_tree_add_7_25_groupi_n_2205);
  not csa_tree_add_7_25_groupi_drc_bufs23727(csa_tree_add_7_25_groupi_n_466 ,csa_tree_add_7_25_groupi_n_464);
  not csa_tree_add_7_25_groupi_drc_bufs23728(csa_tree_add_7_25_groupi_n_465 ,csa_tree_add_7_25_groupi_n_464);
  not csa_tree_add_7_25_groupi_drc_bufs23729(csa_tree_add_7_25_groupi_n_464 ,csa_tree_add_7_25_groupi_n_2203);
  not csa_tree_add_7_25_groupi_drc_bufs23731(csa_tree_add_7_25_groupi_n_463 ,csa_tree_add_7_25_groupi_n_461);
  not csa_tree_add_7_25_groupi_drc_bufs23732(csa_tree_add_7_25_groupi_n_462 ,csa_tree_add_7_25_groupi_n_461);
  not csa_tree_add_7_25_groupi_drc_bufs23733(csa_tree_add_7_25_groupi_n_461 ,csa_tree_add_7_25_groupi_n_2201);
  not csa_tree_add_7_25_groupi_drc_bufs23735(csa_tree_add_7_25_groupi_n_460 ,csa_tree_add_7_25_groupi_n_458);
  not csa_tree_add_7_25_groupi_drc_bufs23736(csa_tree_add_7_25_groupi_n_459 ,csa_tree_add_7_25_groupi_n_458);
  not csa_tree_add_7_25_groupi_drc_bufs23737(csa_tree_add_7_25_groupi_n_458 ,csa_tree_add_7_25_groupi_n_2213);
  not csa_tree_add_7_25_groupi_drc_bufs23739(csa_tree_add_7_25_groupi_n_457 ,csa_tree_add_7_25_groupi_n_455);
  not csa_tree_add_7_25_groupi_drc_bufs23740(csa_tree_add_7_25_groupi_n_456 ,csa_tree_add_7_25_groupi_n_455);
  not csa_tree_add_7_25_groupi_drc_bufs23741(csa_tree_add_7_25_groupi_n_455 ,csa_tree_add_7_25_groupi_n_2211);
  not csa_tree_add_7_25_groupi_drc_bufs23743(csa_tree_add_7_25_groupi_n_454 ,csa_tree_add_7_25_groupi_n_452);
  not csa_tree_add_7_25_groupi_drc_bufs23744(csa_tree_add_7_25_groupi_n_453 ,csa_tree_add_7_25_groupi_n_452);
  not csa_tree_add_7_25_groupi_drc_bufs23745(csa_tree_add_7_25_groupi_n_452 ,csa_tree_add_7_25_groupi_n_2212);
  not csa_tree_add_7_25_groupi_drc_bufs23747(csa_tree_add_7_25_groupi_n_451 ,csa_tree_add_7_25_groupi_n_449);
  not csa_tree_add_7_25_groupi_drc_bufs23748(csa_tree_add_7_25_groupi_n_450 ,csa_tree_add_7_25_groupi_n_449);
  not csa_tree_add_7_25_groupi_drc_bufs23749(csa_tree_add_7_25_groupi_n_449 ,csa_tree_add_7_25_groupi_n_2213);
  not csa_tree_add_7_25_groupi_drc_bufs23751(csa_tree_add_7_25_groupi_n_448 ,csa_tree_add_7_25_groupi_n_446);
  not csa_tree_add_7_25_groupi_drc_bufs23752(csa_tree_add_7_25_groupi_n_447 ,csa_tree_add_7_25_groupi_n_446);
  not csa_tree_add_7_25_groupi_drc_bufs23753(csa_tree_add_7_25_groupi_n_446 ,csa_tree_add_7_25_groupi_n_2209);
  not csa_tree_add_7_25_groupi_drc_bufs23755(csa_tree_add_7_25_groupi_n_445 ,csa_tree_add_7_25_groupi_n_443);
  not csa_tree_add_7_25_groupi_drc_bufs23756(csa_tree_add_7_25_groupi_n_444 ,csa_tree_add_7_25_groupi_n_443);
  not csa_tree_add_7_25_groupi_drc_bufs23757(csa_tree_add_7_25_groupi_n_443 ,csa_tree_add_7_25_groupi_n_2207);
  not csa_tree_add_7_25_groupi_drc_bufs23759(csa_tree_add_7_25_groupi_n_442 ,csa_tree_add_7_25_groupi_n_440);
  not csa_tree_add_7_25_groupi_drc_bufs23760(csa_tree_add_7_25_groupi_n_441 ,csa_tree_add_7_25_groupi_n_440);
  not csa_tree_add_7_25_groupi_drc_bufs23761(csa_tree_add_7_25_groupi_n_440 ,csa_tree_add_7_25_groupi_n_2206);
  not csa_tree_add_7_25_groupi_drc_bufs23763(csa_tree_add_7_25_groupi_n_439 ,csa_tree_add_7_25_groupi_n_437);
  not csa_tree_add_7_25_groupi_drc_bufs23764(csa_tree_add_7_25_groupi_n_438 ,csa_tree_add_7_25_groupi_n_437);
  not csa_tree_add_7_25_groupi_drc_bufs23765(csa_tree_add_7_25_groupi_n_437 ,csa_tree_add_7_25_groupi_n_2217);
  not csa_tree_add_7_25_groupi_drc_bufs23767(csa_tree_add_7_25_groupi_n_436 ,csa_tree_add_7_25_groupi_n_434);
  not csa_tree_add_7_25_groupi_drc_bufs23768(csa_tree_add_7_25_groupi_n_435 ,csa_tree_add_7_25_groupi_n_434);
  not csa_tree_add_7_25_groupi_drc_bufs23769(csa_tree_add_7_25_groupi_n_434 ,csa_tree_add_7_25_groupi_n_2242);
  not csa_tree_add_7_25_groupi_drc_bufs23771(csa_tree_add_7_25_groupi_n_433 ,csa_tree_add_7_25_groupi_n_431);
  not csa_tree_add_7_25_groupi_drc_bufs23772(csa_tree_add_7_25_groupi_n_432 ,csa_tree_add_7_25_groupi_n_431);
  not csa_tree_add_7_25_groupi_drc_bufs23773(csa_tree_add_7_25_groupi_n_431 ,csa_tree_add_7_25_groupi_n_2239);
  not csa_tree_add_7_25_groupi_drc_bufs23775(csa_tree_add_7_25_groupi_n_430 ,csa_tree_add_7_25_groupi_n_428);
  not csa_tree_add_7_25_groupi_drc_bufs23776(csa_tree_add_7_25_groupi_n_429 ,csa_tree_add_7_25_groupi_n_428);
  not csa_tree_add_7_25_groupi_drc_bufs23777(csa_tree_add_7_25_groupi_n_428 ,csa_tree_add_7_25_groupi_n_2222);
  not csa_tree_add_7_25_groupi_drc_bufs23779(csa_tree_add_7_25_groupi_n_427 ,csa_tree_add_7_25_groupi_n_425);
  not csa_tree_add_7_25_groupi_drc_bufs23780(csa_tree_add_7_25_groupi_n_426 ,csa_tree_add_7_25_groupi_n_425);
  not csa_tree_add_7_25_groupi_drc_bufs23781(csa_tree_add_7_25_groupi_n_425 ,csa_tree_add_7_25_groupi_n_2238);
  not csa_tree_add_7_25_groupi_drc_bufs23783(csa_tree_add_7_25_groupi_n_424 ,csa_tree_add_7_25_groupi_n_422);
  not csa_tree_add_7_25_groupi_drc_bufs23784(csa_tree_add_7_25_groupi_n_423 ,csa_tree_add_7_25_groupi_n_422);
  not csa_tree_add_7_25_groupi_drc_bufs23785(csa_tree_add_7_25_groupi_n_422 ,csa_tree_add_7_25_groupi_n_2215);
  not csa_tree_add_7_25_groupi_drc_bufs23787(csa_tree_add_7_25_groupi_n_421 ,csa_tree_add_7_25_groupi_n_419);
  not csa_tree_add_7_25_groupi_drc_bufs23788(csa_tree_add_7_25_groupi_n_420 ,csa_tree_add_7_25_groupi_n_419);
  not csa_tree_add_7_25_groupi_drc_bufs23789(csa_tree_add_7_25_groupi_n_419 ,csa_tree_add_7_25_groupi_n_2223);
  not csa_tree_add_7_25_groupi_drc_bufs23791(csa_tree_add_7_25_groupi_n_418 ,csa_tree_add_7_25_groupi_n_416);
  not csa_tree_add_7_25_groupi_drc_bufs23792(csa_tree_add_7_25_groupi_n_417 ,csa_tree_add_7_25_groupi_n_416);
  not csa_tree_add_7_25_groupi_drc_bufs23793(csa_tree_add_7_25_groupi_n_416 ,csa_tree_add_7_25_groupi_n_2226);
  not csa_tree_add_7_25_groupi_drc_bufs23795(csa_tree_add_7_25_groupi_n_415 ,csa_tree_add_7_25_groupi_n_413);
  not csa_tree_add_7_25_groupi_drc_bufs23796(csa_tree_add_7_25_groupi_n_414 ,csa_tree_add_7_25_groupi_n_413);
  not csa_tree_add_7_25_groupi_drc_bufs23797(csa_tree_add_7_25_groupi_n_413 ,csa_tree_add_7_25_groupi_n_2222);
  not csa_tree_add_7_25_groupi_drc_bufs23799(csa_tree_add_7_25_groupi_n_412 ,csa_tree_add_7_25_groupi_n_410);
  not csa_tree_add_7_25_groupi_drc_bufs23800(csa_tree_add_7_25_groupi_n_411 ,csa_tree_add_7_25_groupi_n_410);
  not csa_tree_add_7_25_groupi_drc_bufs23801(csa_tree_add_7_25_groupi_n_410 ,csa_tree_add_7_25_groupi_n_2223);
  not csa_tree_add_7_25_groupi_drc_bufs23803(csa_tree_add_7_25_groupi_n_409 ,csa_tree_add_7_25_groupi_n_407);
  not csa_tree_add_7_25_groupi_drc_bufs23804(csa_tree_add_7_25_groupi_n_408 ,csa_tree_add_7_25_groupi_n_407);
  not csa_tree_add_7_25_groupi_drc_bufs23805(csa_tree_add_7_25_groupi_n_407 ,csa_tree_add_7_25_groupi_n_2216);
  not csa_tree_add_7_25_groupi_drc_bufs23807(csa_tree_add_7_25_groupi_n_406 ,csa_tree_add_7_25_groupi_n_404);
  not csa_tree_add_7_25_groupi_drc_bufs23808(csa_tree_add_7_25_groupi_n_405 ,csa_tree_add_7_25_groupi_n_404);
  not csa_tree_add_7_25_groupi_drc_bufs23809(csa_tree_add_7_25_groupi_n_404 ,csa_tree_add_7_25_groupi_n_2233);
  not csa_tree_add_7_25_groupi_drc_bufs23811(csa_tree_add_7_25_groupi_n_403 ,csa_tree_add_7_25_groupi_n_401);
  not csa_tree_add_7_25_groupi_drc_bufs23812(csa_tree_add_7_25_groupi_n_402 ,csa_tree_add_7_25_groupi_n_401);
  not csa_tree_add_7_25_groupi_drc_bufs23813(csa_tree_add_7_25_groupi_n_401 ,csa_tree_add_7_25_groupi_n_2232);
  not csa_tree_add_7_25_groupi_drc_bufs23815(csa_tree_add_7_25_groupi_n_400 ,csa_tree_add_7_25_groupi_n_398);
  not csa_tree_add_7_25_groupi_drc_bufs23816(csa_tree_add_7_25_groupi_n_399 ,csa_tree_add_7_25_groupi_n_398);
  not csa_tree_add_7_25_groupi_drc_bufs23817(csa_tree_add_7_25_groupi_n_398 ,csa_tree_add_7_25_groupi_n_2229);
  not csa_tree_add_7_25_groupi_drc_bufs23819(csa_tree_add_7_25_groupi_n_397 ,csa_tree_add_7_25_groupi_n_395);
  not csa_tree_add_7_25_groupi_drc_bufs23820(csa_tree_add_7_25_groupi_n_396 ,csa_tree_add_7_25_groupi_n_395);
  not csa_tree_add_7_25_groupi_drc_bufs23821(csa_tree_add_7_25_groupi_n_395 ,csa_tree_add_7_25_groupi_n_2217);
  not csa_tree_add_7_25_groupi_drc_bufs23823(csa_tree_add_7_25_groupi_n_394 ,csa_tree_add_7_25_groupi_n_392);
  not csa_tree_add_7_25_groupi_drc_bufs23824(csa_tree_add_7_25_groupi_n_393 ,csa_tree_add_7_25_groupi_n_392);
  not csa_tree_add_7_25_groupi_drc_bufs23825(csa_tree_add_7_25_groupi_n_392 ,csa_tree_add_7_25_groupi_n_2230);
  not csa_tree_add_7_25_groupi_drc_bufs23827(csa_tree_add_7_25_groupi_n_391 ,csa_tree_add_7_25_groupi_n_389);
  not csa_tree_add_7_25_groupi_drc_bufs23828(csa_tree_add_7_25_groupi_n_390 ,csa_tree_add_7_25_groupi_n_389);
  not csa_tree_add_7_25_groupi_drc_bufs23829(csa_tree_add_7_25_groupi_n_389 ,csa_tree_add_7_25_groupi_n_2216);
  not csa_tree_add_7_25_groupi_drc_bufs23831(csa_tree_add_7_25_groupi_n_388 ,csa_tree_add_7_25_groupi_n_386);
  not csa_tree_add_7_25_groupi_drc_bufs23832(csa_tree_add_7_25_groupi_n_387 ,csa_tree_add_7_25_groupi_n_386);
  not csa_tree_add_7_25_groupi_drc_bufs23833(csa_tree_add_7_25_groupi_n_386 ,csa_tree_add_7_25_groupi_n_2236);
  not csa_tree_add_7_25_groupi_drc_bufs23835(csa_tree_add_7_25_groupi_n_385 ,csa_tree_add_7_25_groupi_n_383);
  not csa_tree_add_7_25_groupi_drc_bufs23836(csa_tree_add_7_25_groupi_n_384 ,csa_tree_add_7_25_groupi_n_383);
  not csa_tree_add_7_25_groupi_drc_bufs23837(csa_tree_add_7_25_groupi_n_383 ,csa_tree_add_7_25_groupi_n_2224);
  not csa_tree_add_7_25_groupi_drc_bufs23839(csa_tree_add_7_25_groupi_n_382 ,csa_tree_add_7_25_groupi_n_380);
  not csa_tree_add_7_25_groupi_drc_bufs23840(csa_tree_add_7_25_groupi_n_381 ,csa_tree_add_7_25_groupi_n_380);
  not csa_tree_add_7_25_groupi_drc_bufs23841(csa_tree_add_7_25_groupi_n_380 ,csa_tree_add_7_25_groupi_n_2219);
  not csa_tree_add_7_25_groupi_drc_bufs23843(csa_tree_add_7_25_groupi_n_379 ,csa_tree_add_7_25_groupi_n_378);
  not csa_tree_add_7_25_groupi_drc_bufs23845(csa_tree_add_7_25_groupi_n_378 ,csa_tree_add_7_25_groupi_n_1937);
  not csa_tree_add_7_25_groupi_drc_bufs23847(csa_tree_add_7_25_groupi_n_377 ,csa_tree_add_7_25_groupi_n_375);
  not csa_tree_add_7_25_groupi_drc_bufs23848(csa_tree_add_7_25_groupi_n_376 ,csa_tree_add_7_25_groupi_n_375);
  not csa_tree_add_7_25_groupi_drc_bufs23849(csa_tree_add_7_25_groupi_n_375 ,csa_tree_add_7_25_groupi_n_2220);
  not csa_tree_add_7_25_groupi_drc_bufs23851(csa_tree_add_7_25_groupi_n_374 ,csa_tree_add_7_25_groupi_n_372);
  not csa_tree_add_7_25_groupi_drc_bufs23852(csa_tree_add_7_25_groupi_n_373 ,csa_tree_add_7_25_groupi_n_372);
  not csa_tree_add_7_25_groupi_drc_bufs23853(csa_tree_add_7_25_groupi_n_372 ,csa_tree_add_7_25_groupi_n_2221);
  not csa_tree_add_7_25_groupi_drc_bufs23855(csa_tree_add_7_25_groupi_n_371 ,csa_tree_add_7_25_groupi_n_369);
  not csa_tree_add_7_25_groupi_drc_bufs23856(csa_tree_add_7_25_groupi_n_370 ,csa_tree_add_7_25_groupi_n_369);
  not csa_tree_add_7_25_groupi_drc_bufs23857(csa_tree_add_7_25_groupi_n_369 ,csa_tree_add_7_25_groupi_n_2221);
  not csa_tree_add_7_25_groupi_drc_bufs23859(csa_tree_add_7_25_groupi_n_368 ,csa_tree_add_7_25_groupi_n_366);
  not csa_tree_add_7_25_groupi_drc_bufs23860(csa_tree_add_7_25_groupi_n_367 ,csa_tree_add_7_25_groupi_n_366);
  not csa_tree_add_7_25_groupi_drc_bufs23861(csa_tree_add_7_25_groupi_n_366 ,csa_tree_add_7_25_groupi_n_2220);
  not csa_tree_add_7_25_groupi_drc_bufs23863(csa_tree_add_7_25_groupi_n_365 ,csa_tree_add_7_25_groupi_n_363);
  not csa_tree_add_7_25_groupi_drc_bufs23864(csa_tree_add_7_25_groupi_n_364 ,csa_tree_add_7_25_groupi_n_363);
  not csa_tree_add_7_25_groupi_drc_bufs23865(csa_tree_add_7_25_groupi_n_363 ,csa_tree_add_7_25_groupi_n_2219);
  not csa_tree_add_7_25_groupi_drc_bufs23867(csa_tree_add_7_25_groupi_n_362 ,csa_tree_add_7_25_groupi_n_361);
  not csa_tree_add_7_25_groupi_drc_bufs23869(csa_tree_add_7_25_groupi_n_361 ,csa_tree_add_7_25_groupi_n_1934);
  not csa_tree_add_7_25_groupi_drc_bufs23871(csa_tree_add_7_25_groupi_n_360 ,csa_tree_add_7_25_groupi_n_358);
  not csa_tree_add_7_25_groupi_drc_bufs23872(csa_tree_add_7_25_groupi_n_359 ,csa_tree_add_7_25_groupi_n_358);
  not csa_tree_add_7_25_groupi_drc_bufs23873(csa_tree_add_7_25_groupi_n_358 ,csa_tree_add_7_25_groupi_n_2231);
  not csa_tree_add_7_25_groupi_drc_bufs23875(csa_tree_add_7_25_groupi_n_357 ,csa_tree_add_7_25_groupi_n_355);
  not csa_tree_add_7_25_groupi_drc_bufs23876(csa_tree_add_7_25_groupi_n_356 ,csa_tree_add_7_25_groupi_n_355);
  not csa_tree_add_7_25_groupi_drc_bufs23877(csa_tree_add_7_25_groupi_n_355 ,csa_tree_add_7_25_groupi_n_2218);
  not csa_tree_add_7_25_groupi_drc_bufs23879(csa_tree_add_7_25_groupi_n_354 ,csa_tree_add_7_25_groupi_n_352);
  not csa_tree_add_7_25_groupi_drc_bufs23880(csa_tree_add_7_25_groupi_n_353 ,csa_tree_add_7_25_groupi_n_352);
  not csa_tree_add_7_25_groupi_drc_bufs23881(csa_tree_add_7_25_groupi_n_352 ,csa_tree_add_7_25_groupi_n_2226);
  not csa_tree_add_7_25_groupi_drc_bufs23883(csa_tree_add_7_25_groupi_n_351 ,csa_tree_add_7_25_groupi_n_349);
  not csa_tree_add_7_25_groupi_drc_bufs23884(csa_tree_add_7_25_groupi_n_350 ,csa_tree_add_7_25_groupi_n_349);
  not csa_tree_add_7_25_groupi_drc_bufs23885(csa_tree_add_7_25_groupi_n_349 ,csa_tree_add_7_25_groupi_n_2225);
  not csa_tree_add_7_25_groupi_drc_bufs23887(csa_tree_add_7_25_groupi_n_348 ,csa_tree_add_7_25_groupi_n_346);
  not csa_tree_add_7_25_groupi_drc_bufs23888(csa_tree_add_7_25_groupi_n_347 ,csa_tree_add_7_25_groupi_n_346);
  not csa_tree_add_7_25_groupi_drc_bufs23889(csa_tree_add_7_25_groupi_n_346 ,csa_tree_add_7_25_groupi_n_2214);
  not csa_tree_add_7_25_groupi_drc_bufs23891(csa_tree_add_7_25_groupi_n_345 ,csa_tree_add_7_25_groupi_n_343);
  not csa_tree_add_7_25_groupi_drc_bufs23892(csa_tree_add_7_25_groupi_n_344 ,csa_tree_add_7_25_groupi_n_343);
  not csa_tree_add_7_25_groupi_drc_bufs23893(csa_tree_add_7_25_groupi_n_343 ,csa_tree_add_7_25_groupi_n_2227);
  not csa_tree_add_7_25_groupi_drc_bufs23895(csa_tree_add_7_25_groupi_n_342 ,csa_tree_add_7_25_groupi_n_340);
  not csa_tree_add_7_25_groupi_drc_bufs23896(csa_tree_add_7_25_groupi_n_341 ,csa_tree_add_7_25_groupi_n_340);
  not csa_tree_add_7_25_groupi_drc_bufs23897(csa_tree_add_7_25_groupi_n_340 ,csa_tree_add_7_25_groupi_n_2228);
  not csa_tree_add_7_25_groupi_drc_bufs23899(csa_tree_add_7_25_groupi_n_339 ,csa_tree_add_7_25_groupi_n_337);
  not csa_tree_add_7_25_groupi_drc_bufs23900(csa_tree_add_7_25_groupi_n_338 ,csa_tree_add_7_25_groupi_n_337);
  not csa_tree_add_7_25_groupi_drc_bufs23901(csa_tree_add_7_25_groupi_n_337 ,csa_tree_add_7_25_groupi_n_5188);
  not csa_tree_add_7_25_groupi_drc_bufs23903(csa_tree_add_7_25_groupi_n_336 ,csa_tree_add_7_25_groupi_n_334);
  not csa_tree_add_7_25_groupi_drc_bufs23904(csa_tree_add_7_25_groupi_n_335 ,csa_tree_add_7_25_groupi_n_334);
  not csa_tree_add_7_25_groupi_drc_bufs23905(csa_tree_add_7_25_groupi_n_334 ,csa_tree_add_7_25_groupi_n_5188);
  not csa_tree_add_7_25_groupi_drc_bufs23907(csa_tree_add_7_25_groupi_n_333 ,csa_tree_add_7_25_groupi_n_331);
  not csa_tree_add_7_25_groupi_drc_bufs23908(csa_tree_add_7_25_groupi_n_332 ,csa_tree_add_7_25_groupi_n_331);
  not csa_tree_add_7_25_groupi_drc_bufs23909(csa_tree_add_7_25_groupi_n_331 ,csa_tree_add_7_25_groupi_n_4676);
  not csa_tree_add_7_25_groupi_drc_bufs23911(csa_tree_add_7_25_groupi_n_330 ,csa_tree_add_7_25_groupi_n_328);
  not csa_tree_add_7_25_groupi_drc_bufs23912(csa_tree_add_7_25_groupi_n_329 ,csa_tree_add_7_25_groupi_n_328);
  not csa_tree_add_7_25_groupi_drc_bufs23913(csa_tree_add_7_25_groupi_n_328 ,csa_tree_add_7_25_groupi_n_4460);
  not csa_tree_add_7_25_groupi_drc_bufs23915(csa_tree_add_7_25_groupi_n_327 ,csa_tree_add_7_25_groupi_n_325);
  not csa_tree_add_7_25_groupi_drc_bufs23916(csa_tree_add_7_25_groupi_n_326 ,csa_tree_add_7_25_groupi_n_325);
  not csa_tree_add_7_25_groupi_drc_bufs23917(csa_tree_add_7_25_groupi_n_325 ,csa_tree_add_7_25_groupi_n_4198);
  not csa_tree_add_7_25_groupi_drc_bufs23919(csa_tree_add_7_25_groupi_n_324 ,csa_tree_add_7_25_groupi_n_322);
  not csa_tree_add_7_25_groupi_drc_bufs23920(csa_tree_add_7_25_groupi_n_323 ,csa_tree_add_7_25_groupi_n_322);
  not csa_tree_add_7_25_groupi_drc_bufs23921(csa_tree_add_7_25_groupi_n_322 ,csa_tree_add_7_25_groupi_n_4110);
  not csa_tree_add_7_25_groupi_drc_bufs23923(csa_tree_add_7_25_groupi_n_321 ,csa_tree_add_7_25_groupi_n_319);
  not csa_tree_add_7_25_groupi_drc_bufs23924(csa_tree_add_7_25_groupi_n_320 ,csa_tree_add_7_25_groupi_n_319);
  not csa_tree_add_7_25_groupi_drc_bufs23925(csa_tree_add_7_25_groupi_n_319 ,csa_tree_add_7_25_groupi_n_4573);
  not csa_tree_add_7_25_groupi_drc_bufs23927(csa_tree_add_7_25_groupi_n_318 ,csa_tree_add_7_25_groupi_n_316);
  not csa_tree_add_7_25_groupi_drc_bufs23928(csa_tree_add_7_25_groupi_n_317 ,csa_tree_add_7_25_groupi_n_316);
  not csa_tree_add_7_25_groupi_drc_bufs23929(csa_tree_add_7_25_groupi_n_316 ,csa_tree_add_7_25_groupi_n_3742);
  not csa_tree_add_7_25_groupi_drc_bufs23931(csa_tree_add_7_25_groupi_n_315 ,csa_tree_add_7_25_groupi_n_313);
  not csa_tree_add_7_25_groupi_drc_bufs23932(csa_tree_add_7_25_groupi_n_314 ,csa_tree_add_7_25_groupi_n_313);
  not csa_tree_add_7_25_groupi_drc_bufs23933(csa_tree_add_7_25_groupi_n_313 ,csa_tree_add_7_25_groupi_n_5007);
  not csa_tree_add_7_25_groupi_drc_bufs23935(csa_tree_add_7_25_groupi_n_312 ,csa_tree_add_7_25_groupi_n_310);
  not csa_tree_add_7_25_groupi_drc_bufs23936(csa_tree_add_7_25_groupi_n_311 ,csa_tree_add_7_25_groupi_n_310);
  not csa_tree_add_7_25_groupi_drc_bufs23937(csa_tree_add_7_25_groupi_n_310 ,csa_tree_add_7_25_groupi_n_3199);
  not csa_tree_add_7_25_groupi_drc_bufs23939(csa_tree_add_7_25_groupi_n_309 ,csa_tree_add_7_25_groupi_n_307);
  not csa_tree_add_7_25_groupi_drc_bufs23940(csa_tree_add_7_25_groupi_n_308 ,csa_tree_add_7_25_groupi_n_307);
  not csa_tree_add_7_25_groupi_drc_bufs23941(csa_tree_add_7_25_groupi_n_307 ,csa_tree_add_7_25_groupi_n_4676);
  not csa_tree_add_7_25_groupi_drc_bufs23943(csa_tree_add_7_25_groupi_n_306 ,csa_tree_add_7_25_groupi_n_304);
  not csa_tree_add_7_25_groupi_drc_bufs23944(csa_tree_add_7_25_groupi_n_305 ,csa_tree_add_7_25_groupi_n_304);
  not csa_tree_add_7_25_groupi_drc_bufs23945(csa_tree_add_7_25_groupi_n_304 ,csa_tree_add_7_25_groupi_n_4792);
  not csa_tree_add_7_25_groupi_drc_bufs23947(csa_tree_add_7_25_groupi_n_303 ,csa_tree_add_7_25_groupi_n_301);
  not csa_tree_add_7_25_groupi_drc_bufs23948(csa_tree_add_7_25_groupi_n_302 ,csa_tree_add_7_25_groupi_n_301);
  not csa_tree_add_7_25_groupi_drc_bufs23949(csa_tree_add_7_25_groupi_n_301 ,csa_tree_add_7_25_groupi_n_5093);
  not csa_tree_add_7_25_groupi_drc_bufs23951(csa_tree_add_7_25_groupi_n_300 ,csa_tree_add_7_25_groupi_n_299);
  not csa_tree_add_7_25_groupi_drc_bufs23953(csa_tree_add_7_25_groupi_n_299 ,csa_tree_add_7_25_groupi_n_1876);
  not csa_tree_add_7_25_groupi_drc_bufs23955(csa_tree_add_7_25_groupi_n_298 ,csa_tree_add_7_25_groupi_n_296);
  not csa_tree_add_7_25_groupi_drc_bufs23956(csa_tree_add_7_25_groupi_n_297 ,csa_tree_add_7_25_groupi_n_296);
  not csa_tree_add_7_25_groupi_drc_bufs23957(csa_tree_add_7_25_groupi_n_296 ,csa_tree_add_7_25_groupi_n_2210);
  not csa_tree_add_7_25_groupi_drc_bufs23959(csa_tree_add_7_25_groupi_n_295 ,csa_tree_add_7_25_groupi_n_293);
  not csa_tree_add_7_25_groupi_drc_bufs23960(csa_tree_add_7_25_groupi_n_294 ,csa_tree_add_7_25_groupi_n_293);
  not csa_tree_add_7_25_groupi_drc_bufs23961(csa_tree_add_7_25_groupi_n_293 ,csa_tree_add_7_25_groupi_n_4351);
  not csa_tree_add_7_25_groupi_drc_bufs23963(csa_tree_add_7_25_groupi_n_292 ,csa_tree_add_7_25_groupi_n_290);
  not csa_tree_add_7_25_groupi_drc_bufs23964(csa_tree_add_7_25_groupi_n_291 ,csa_tree_add_7_25_groupi_n_290);
  not csa_tree_add_7_25_groupi_drc_bufs23965(csa_tree_add_7_25_groupi_n_290 ,csa_tree_add_7_25_groupi_n_3742);
  not csa_tree_add_7_25_groupi_drc_bufs23967(csa_tree_add_7_25_groupi_n_289 ,csa_tree_add_7_25_groupi_n_287);
  not csa_tree_add_7_25_groupi_drc_bufs23968(csa_tree_add_7_25_groupi_n_288 ,csa_tree_add_7_25_groupi_n_287);
  not csa_tree_add_7_25_groupi_drc_bufs23969(csa_tree_add_7_25_groupi_n_287 ,csa_tree_add_7_25_groupi_n_4792);
  not csa_tree_add_7_25_groupi_drc_bufs23971(csa_tree_add_7_25_groupi_n_286 ,csa_tree_add_7_25_groupi_n_284);
  not csa_tree_add_7_25_groupi_drc_bufs23972(csa_tree_add_7_25_groupi_n_285 ,csa_tree_add_7_25_groupi_n_284);
  not csa_tree_add_7_25_groupi_drc_bufs23973(csa_tree_add_7_25_groupi_n_284 ,csa_tree_add_7_25_groupi_n_3199);
  not csa_tree_add_7_25_groupi_drc_bufs23975(csa_tree_add_7_25_groupi_n_283 ,csa_tree_add_7_25_groupi_n_281);
  not csa_tree_add_7_25_groupi_drc_bufs23976(csa_tree_add_7_25_groupi_n_282 ,csa_tree_add_7_25_groupi_n_281);
  not csa_tree_add_7_25_groupi_drc_bufs23977(csa_tree_add_7_25_groupi_n_281 ,csa_tree_add_7_25_groupi_n_5007);
  not csa_tree_add_7_25_groupi_drc_bufs23979(csa_tree_add_7_25_groupi_n_280 ,csa_tree_add_7_25_groupi_n_278);
  not csa_tree_add_7_25_groupi_drc_bufs23980(csa_tree_add_7_25_groupi_n_279 ,csa_tree_add_7_25_groupi_n_278);
  not csa_tree_add_7_25_groupi_drc_bufs23981(csa_tree_add_7_25_groupi_n_278 ,csa_tree_add_7_25_groupi_n_5093);
  not csa_tree_add_7_25_groupi_drc_bufs23983(csa_tree_add_7_25_groupi_n_277 ,csa_tree_add_7_25_groupi_n_275);
  not csa_tree_add_7_25_groupi_drc_bufs23984(csa_tree_add_7_25_groupi_n_276 ,csa_tree_add_7_25_groupi_n_275);
  not csa_tree_add_7_25_groupi_drc_bufs23985(csa_tree_add_7_25_groupi_n_275 ,csa_tree_add_7_25_groupi_n_2614);
  not csa_tree_add_7_25_groupi_drc_bufs23987(csa_tree_add_7_25_groupi_n_274 ,csa_tree_add_7_25_groupi_n_272);
  not csa_tree_add_7_25_groupi_drc_bufs23988(csa_tree_add_7_25_groupi_n_273 ,csa_tree_add_7_25_groupi_n_272);
  not csa_tree_add_7_25_groupi_drc_bufs23989(csa_tree_add_7_25_groupi_n_272 ,csa_tree_add_7_25_groupi_n_4198);
  not csa_tree_add_7_25_groupi_drc_bufs23991(csa_tree_add_7_25_groupi_n_271 ,csa_tree_add_7_25_groupi_n_269);
  not csa_tree_add_7_25_groupi_drc_bufs23992(csa_tree_add_7_25_groupi_n_270 ,csa_tree_add_7_25_groupi_n_269);
  not csa_tree_add_7_25_groupi_drc_bufs23993(csa_tree_add_7_25_groupi_n_269 ,csa_tree_add_7_25_groupi_n_4573);
  not csa_tree_add_7_25_groupi_drc_bufs23995(csa_tree_add_7_25_groupi_n_268 ,csa_tree_add_7_25_groupi_n_267);
  not csa_tree_add_7_25_groupi_drc_bufs23997(csa_tree_add_7_25_groupi_n_267 ,csa_tree_add_7_25_groupi_n_4351);
  not csa_tree_add_7_25_groupi_drc_bufs23999(csa_tree_add_7_25_groupi_n_266 ,csa_tree_add_7_25_groupi_n_265);
  not csa_tree_add_7_25_groupi_drc_bufs24001(csa_tree_add_7_25_groupi_n_265 ,csa_tree_add_7_25_groupi_n_1879);
  not csa_tree_add_7_25_groupi_drc_bufs24003(csa_tree_add_7_25_groupi_n_264 ,csa_tree_add_7_25_groupi_n_262);
  not csa_tree_add_7_25_groupi_drc_bufs24004(csa_tree_add_7_25_groupi_n_263 ,csa_tree_add_7_25_groupi_n_262);
  not csa_tree_add_7_25_groupi_drc_bufs24005(csa_tree_add_7_25_groupi_n_262 ,csa_tree_add_7_25_groupi_n_5303);
  not csa_tree_add_7_25_groupi_drc_bufs24007(csa_tree_add_7_25_groupi_n_261 ,csa_tree_add_7_25_groupi_n_259);
  not csa_tree_add_7_25_groupi_drc_bufs24008(csa_tree_add_7_25_groupi_n_260 ,csa_tree_add_7_25_groupi_n_259);
  not csa_tree_add_7_25_groupi_drc_bufs24009(csa_tree_add_7_25_groupi_n_259 ,csa_tree_add_7_25_groupi_n_5303);
  not csa_tree_add_7_25_groupi_drc_bufs24011(csa_tree_add_7_25_groupi_n_258 ,csa_tree_add_7_25_groupi_n_256);
  not csa_tree_add_7_25_groupi_drc_bufs24012(csa_tree_add_7_25_groupi_n_257 ,csa_tree_add_7_25_groupi_n_256);
  not csa_tree_add_7_25_groupi_drc_bufs24013(csa_tree_add_7_25_groupi_n_256 ,csa_tree_add_7_25_groupi_n_4460);
  not csa_tree_add_7_25_groupi_drc_bufs24015(csa_tree_add_7_25_groupi_n_255 ,csa_tree_add_7_25_groupi_n_253);
  not csa_tree_add_7_25_groupi_drc_bufs24016(csa_tree_add_7_25_groupi_n_254 ,csa_tree_add_7_25_groupi_n_253);
  not csa_tree_add_7_25_groupi_drc_bufs24017(csa_tree_add_7_25_groupi_n_253 ,csa_tree_add_7_25_groupi_n_4903);
  not csa_tree_add_7_25_groupi_drc_bufs24019(csa_tree_add_7_25_groupi_n_252 ,csa_tree_add_7_25_groupi_n_250);
  not csa_tree_add_7_25_groupi_drc_bufs24020(csa_tree_add_7_25_groupi_n_251 ,csa_tree_add_7_25_groupi_n_250);
  not csa_tree_add_7_25_groupi_drc_bufs24021(csa_tree_add_7_25_groupi_n_250 ,csa_tree_add_7_25_groupi_n_4903);
  not csa_tree_add_7_25_groupi_drc_bufs24023(csa_tree_add_7_25_groupi_n_249 ,csa_tree_add_7_25_groupi_n_247);
  not csa_tree_add_7_25_groupi_drc_bufs24024(csa_tree_add_7_25_groupi_n_248 ,csa_tree_add_7_25_groupi_n_247);
  not csa_tree_add_7_25_groupi_drc_bufs24025(csa_tree_add_7_25_groupi_n_247 ,csa_tree_add_7_25_groupi_n_4110);
  not csa_tree_add_7_25_groupi_drc_bufs24027(csa_tree_add_7_25_groupi_n_246 ,csa_tree_add_7_25_groupi_n_245);
  not csa_tree_add_7_25_groupi_drc_bufs24029(csa_tree_add_7_25_groupi_n_245 ,csa_tree_add_7_25_groupi_n_1914);
  not csa_tree_add_7_25_groupi_drc_bufs24031(csa_tree_add_7_25_groupi_n_244 ,csa_tree_add_7_25_groupi_n_242);
  not csa_tree_add_7_25_groupi_drc_bufs24032(csa_tree_add_7_25_groupi_n_243 ,csa_tree_add_7_25_groupi_n_242);
  not csa_tree_add_7_25_groupi_drc_bufs24033(csa_tree_add_7_25_groupi_n_242 ,csa_tree_add_7_25_groupi_n_2214);
  not csa_tree_add_7_25_groupi_drc_bufs24035(csa_tree_add_7_25_groupi_n_241 ,csa_tree_add_7_25_groupi_n_240);
  not csa_tree_add_7_25_groupi_drc_bufs24037(csa_tree_add_7_25_groupi_n_240 ,csa_tree_add_7_25_groupi_n_1916);
  not csa_tree_add_7_25_groupi_drc_bufs24039(csa_tree_add_7_25_groupi_n_239 ,csa_tree_add_7_25_groupi_n_237);
  not csa_tree_add_7_25_groupi_drc_bufs24040(csa_tree_add_7_25_groupi_n_238 ,csa_tree_add_7_25_groupi_n_237);
  not csa_tree_add_7_25_groupi_drc_bufs24041(csa_tree_add_7_25_groupi_n_237 ,csa_tree_add_7_25_groupi_n_2199);
  not csa_tree_add_7_25_groupi_drc_bufs24043(csa_tree_add_7_25_groupi_n_236 ,csa_tree_add_7_25_groupi_n_234);
  not csa_tree_add_7_25_groupi_drc_bufs24044(csa_tree_add_7_25_groupi_n_235 ,csa_tree_add_7_25_groupi_n_234);
  not csa_tree_add_7_25_groupi_drc_bufs24045(csa_tree_add_7_25_groupi_n_234 ,csa_tree_add_7_25_groupi_n_2209);
  not csa_tree_add_7_25_groupi_drc_bufs24047(csa_tree_add_7_25_groupi_n_233 ,csa_tree_add_7_25_groupi_n_231);
  not csa_tree_add_7_25_groupi_drc_bufs24048(csa_tree_add_7_25_groupi_n_232 ,csa_tree_add_7_25_groupi_n_231);
  not csa_tree_add_7_25_groupi_drc_bufs24049(csa_tree_add_7_25_groupi_n_231 ,csa_tree_add_7_25_groupi_n_2202);
  not csa_tree_add_7_25_groupi_drc_bufs24051(csa_tree_add_7_25_groupi_n_230 ,csa_tree_add_7_25_groupi_n_228);
  not csa_tree_add_7_25_groupi_drc_bufs24052(csa_tree_add_7_25_groupi_n_229 ,csa_tree_add_7_25_groupi_n_228);
  not csa_tree_add_7_25_groupi_drc_bufs24053(csa_tree_add_7_25_groupi_n_228 ,csa_tree_add_7_25_groupi_n_2208);
  not csa_tree_add_7_25_groupi_drc_bufs24055(csa_tree_add_7_25_groupi_n_227 ,csa_tree_add_7_25_groupi_n_225);
  not csa_tree_add_7_25_groupi_drc_bufs24056(csa_tree_add_7_25_groupi_n_226 ,csa_tree_add_7_25_groupi_n_225);
  not csa_tree_add_7_25_groupi_drc_bufs24057(csa_tree_add_7_25_groupi_n_225 ,csa_tree_add_7_25_groupi_n_2212);
  not csa_tree_add_7_25_groupi_drc_bufs24059(csa_tree_add_7_25_groupi_n_224 ,csa_tree_add_7_25_groupi_n_222);
  not csa_tree_add_7_25_groupi_drc_bufs24060(csa_tree_add_7_25_groupi_n_223 ,csa_tree_add_7_25_groupi_n_222);
  not csa_tree_add_7_25_groupi_drc_bufs24061(csa_tree_add_7_25_groupi_n_222 ,csa_tree_add_7_25_groupi_n_2211);
  not csa_tree_add_7_25_groupi_drc_bufs24063(csa_tree_add_7_25_groupi_n_221 ,csa_tree_add_7_25_groupi_n_219);
  not csa_tree_add_7_25_groupi_drc_bufs24064(csa_tree_add_7_25_groupi_n_220 ,csa_tree_add_7_25_groupi_n_219);
  not csa_tree_add_7_25_groupi_drc_bufs24065(csa_tree_add_7_25_groupi_n_219 ,csa_tree_add_7_25_groupi_n_2202);
  not csa_tree_add_7_25_groupi_drc_bufs24067(csa_tree_add_7_25_groupi_n_218 ,csa_tree_add_7_25_groupi_n_216);
  not csa_tree_add_7_25_groupi_drc_bufs24068(csa_tree_add_7_25_groupi_n_217 ,csa_tree_add_7_25_groupi_n_216);
  not csa_tree_add_7_25_groupi_drc_bufs24069(csa_tree_add_7_25_groupi_n_216 ,csa_tree_add_7_25_groupi_n_2215);
  not csa_tree_add_7_25_groupi_drc_bufs24071(csa_tree_add_7_25_groupi_n_215 ,csa_tree_add_7_25_groupi_n_213);
  not csa_tree_add_7_25_groupi_drc_bufs24072(csa_tree_add_7_25_groupi_n_214 ,csa_tree_add_7_25_groupi_n_213);
  not csa_tree_add_7_25_groupi_drc_bufs24073(csa_tree_add_7_25_groupi_n_213 ,csa_tree_add_7_25_groupi_n_2198);
  not csa_tree_add_7_25_groupi_drc_bufs24075(csa_tree_add_7_25_groupi_n_212 ,csa_tree_add_7_25_groupi_n_210);
  not csa_tree_add_7_25_groupi_drc_bufs24076(csa_tree_add_7_25_groupi_n_211 ,csa_tree_add_7_25_groupi_n_210);
  not csa_tree_add_7_25_groupi_drc_bufs24077(csa_tree_add_7_25_groupi_n_210 ,csa_tree_add_7_25_groupi_n_2614);
  not csa_tree_add_7_25_groupi_drc_bufs24079(csa_tree_add_7_25_groupi_n_209 ,csa_tree_add_7_25_groupi_n_207);
  not csa_tree_add_7_25_groupi_drc_bufs24080(csa_tree_add_7_25_groupi_n_208 ,csa_tree_add_7_25_groupi_n_207);
  not csa_tree_add_7_25_groupi_drc_bufs24081(csa_tree_add_7_25_groupi_n_207 ,csa_tree_add_7_25_groupi_n_5533);
  not csa_tree_add_7_25_groupi_drc_bufs24083(csa_tree_add_7_25_groupi_n_206 ,csa_tree_add_7_25_groupi_n_205);
  not csa_tree_add_7_25_groupi_drc_bufs24085(csa_tree_add_7_25_groupi_n_205 ,csa_tree_add_7_25_groupi_n_1872);
  not csa_tree_add_7_25_groupi_drc_bufs24087(csa_tree_add_7_25_groupi_n_204 ,csa_tree_add_7_25_groupi_n_203);
  not csa_tree_add_7_25_groupi_drc_bufs24089(csa_tree_add_7_25_groupi_n_203 ,csa_tree_add_7_25_groupi_n_1840);
  not csa_tree_add_7_25_groupi_drc_bufs24091(csa_tree_add_7_25_groupi_n_202 ,csa_tree_add_7_25_groupi_n_201);
  not csa_tree_add_7_25_groupi_drc_bufs24093(csa_tree_add_7_25_groupi_n_201 ,csa_tree_add_7_25_groupi_n_1908);
  not csa_tree_add_7_25_groupi_drc_bufs24095(csa_tree_add_7_25_groupi_n_200 ,csa_tree_add_7_25_groupi_n_199);
  not csa_tree_add_7_25_groupi_drc_bufs24097(csa_tree_add_7_25_groupi_n_199 ,csa_tree_add_7_25_groupi_n_1931);
  not csa_tree_add_7_25_groupi_drc_bufs24099(csa_tree_add_7_25_groupi_n_198 ,csa_tree_add_7_25_groupi_n_197);
  not csa_tree_add_7_25_groupi_drc_bufs24101(csa_tree_add_7_25_groupi_n_197 ,csa_tree_add_7_25_groupi_n_1904);
  not csa_tree_add_7_25_groupi_drc_bufs24103(csa_tree_add_7_25_groupi_n_196 ,csa_tree_add_7_25_groupi_n_194);
  not csa_tree_add_7_25_groupi_drc_bufs24104(csa_tree_add_7_25_groupi_n_195 ,csa_tree_add_7_25_groupi_n_194);
  not csa_tree_add_7_25_groupi_drc_bufs24105(csa_tree_add_7_25_groupi_n_194 ,csa_tree_add_7_25_groupi_n_5763);
  not csa_tree_add_7_25_groupi_drc_bufs24107(csa_tree_add_7_25_groupi_n_193 ,csa_tree_add_7_25_groupi_n_191);
  not csa_tree_add_7_25_groupi_drc_bufs24108(csa_tree_add_7_25_groupi_n_192 ,csa_tree_add_7_25_groupi_n_191);
  not csa_tree_add_7_25_groupi_drc_bufs24109(csa_tree_add_7_25_groupi_n_191 ,csa_tree_add_7_25_groupi_n_5648);
  not csa_tree_add_7_25_groupi_drc_bufs24111(csa_tree_add_7_25_groupi_n_190 ,csa_tree_add_7_25_groupi_n_188);
  not csa_tree_add_7_25_groupi_drc_bufs24112(csa_tree_add_7_25_groupi_n_189 ,csa_tree_add_7_25_groupi_n_188);
  not csa_tree_add_7_25_groupi_drc_bufs24113(csa_tree_add_7_25_groupi_n_188 ,csa_tree_add_7_25_groupi_n_5423);
  not csa_tree_add_7_25_groupi_drc_bufs24115(csa_tree_add_7_25_groupi_n_187 ,csa_tree_add_7_25_groupi_n_186);
  not csa_tree_add_7_25_groupi_drc_bufs24117(csa_tree_add_7_25_groupi_n_186 ,csa_tree_add_7_25_groupi_n_1828);
  not csa_tree_add_7_25_groupi_drc_bufs24119(csa_tree_add_7_25_groupi_n_185 ,csa_tree_add_7_25_groupi_n_184);
  not csa_tree_add_7_25_groupi_drc_bufs24121(csa_tree_add_7_25_groupi_n_184 ,csa_tree_add_7_25_groupi_n_1819);
  not csa_tree_add_7_25_groupi_drc_bufs24123(csa_tree_add_7_25_groupi_n_183 ,csa_tree_add_7_25_groupi_n_182);
  not csa_tree_add_7_25_groupi_drc_bufs24125(csa_tree_add_7_25_groupi_n_182 ,csa_tree_add_7_25_groupi_n_1902);
  not csa_tree_add_7_25_groupi_drc_bufs24127(csa_tree_add_7_25_groupi_n_181 ,csa_tree_add_7_25_groupi_n_180);
  not csa_tree_add_7_25_groupi_drc_bufs24129(csa_tree_add_7_25_groupi_n_180 ,csa_tree_add_7_25_groupi_n_1837);
  not csa_tree_add_7_25_groupi_drc_bufs24131(csa_tree_add_7_25_groupi_n_179 ,csa_tree_add_7_25_groupi_n_178);
  not csa_tree_add_7_25_groupi_drc_bufs24133(csa_tree_add_7_25_groupi_n_178 ,csa_tree_add_7_25_groupi_n_1813);
  not csa_tree_add_7_25_groupi_drc_bufs24135(csa_tree_add_7_25_groupi_n_177 ,csa_tree_add_7_25_groupi_n_175);
  not csa_tree_add_7_25_groupi_drc_bufs24136(csa_tree_add_7_25_groupi_n_176 ,csa_tree_add_7_25_groupi_n_175);
  not csa_tree_add_7_25_groupi_drc_bufs24137(csa_tree_add_7_25_groupi_n_175 ,csa_tree_add_7_25_groupi_n_5979);
  not csa_tree_add_7_25_groupi_drc_bufs24139(csa_tree_add_7_25_groupi_n_174 ,csa_tree_add_7_25_groupi_n_173);
  not csa_tree_add_7_25_groupi_drc_bufs24141(csa_tree_add_7_25_groupi_n_173 ,csa_tree_add_7_25_groupi_n_1822);
  not csa_tree_add_7_25_groupi_drc_bufs24143(csa_tree_add_7_25_groupi_n_172 ,csa_tree_add_7_25_groupi_n_171);
  not csa_tree_add_7_25_groupi_drc_bufs24145(csa_tree_add_7_25_groupi_n_171 ,csa_tree_add_7_25_groupi_n_1816);
  not csa_tree_add_7_25_groupi_drc_bufs24147(csa_tree_add_7_25_groupi_n_170 ,csa_tree_add_7_25_groupi_n_169);
  not csa_tree_add_7_25_groupi_drc_bufs24149(csa_tree_add_7_25_groupi_n_169 ,csa_tree_add_7_25_groupi_n_1911);
  not csa_tree_add_7_25_groupi_drc_bufs24151(csa_tree_add_7_25_groupi_n_168 ,csa_tree_add_7_25_groupi_n_167);
  not csa_tree_add_7_25_groupi_drc_bufs24153(csa_tree_add_7_25_groupi_n_167 ,csa_tree_add_7_25_groupi_n_1905);
  not csa_tree_add_7_25_groupi_drc_bufs24155(csa_tree_add_7_25_groupi_n_166 ,csa_tree_add_7_25_groupi_n_165);
  not csa_tree_add_7_25_groupi_drc_bufs24157(csa_tree_add_7_25_groupi_n_165 ,csa_tree_add_7_25_groupi_n_1864);
  not csa_tree_add_7_25_groupi_drc_bufs24159(csa_tree_add_7_25_groupi_n_164 ,csa_tree_add_7_25_groupi_n_163);
  not csa_tree_add_7_25_groupi_drc_bufs24161(csa_tree_add_7_25_groupi_n_163 ,csa_tree_add_7_25_groupi_n_1928);
  not csa_tree_add_7_25_groupi_drc_bufs24163(csa_tree_add_7_25_groupi_n_162 ,csa_tree_add_7_25_groupi_n_161);
  not csa_tree_add_7_25_groupi_drc_bufs24165(csa_tree_add_7_25_groupi_n_161 ,csa_tree_add_7_25_groupi_n_1913);
  not csa_tree_add_7_25_groupi_drc_bufs24167(csa_tree_add_7_25_groupi_n_160 ,csa_tree_add_7_25_groupi_n_2335);
  not csa_tree_add_7_25_groupi_drc_bufs24169(csa_tree_add_7_25_groupi_n_2335 ,csa_tree_add_7_25_groupi_n_2837);
  not csa_tree_add_7_25_groupi_drc_bufs24171(csa_tree_add_7_25_groupi_n_159 ,csa_tree_add_7_25_groupi_n_158);
  not csa_tree_add_7_25_groupi_drc_bufs24173(csa_tree_add_7_25_groupi_n_158 ,csa_tree_add_7_25_groupi_n_1834);
  not csa_tree_add_7_25_groupi_drc_bufs24175(csa_tree_add_7_25_groupi_n_157 ,csa_tree_add_7_25_groupi_n_156);
  not csa_tree_add_7_25_groupi_drc_bufs24177(csa_tree_add_7_25_groupi_n_156 ,csa_tree_add_7_25_groupi_n_1843);
  not csa_tree_add_7_25_groupi_drc_bufs24179(csa_tree_add_7_25_groupi_n_155 ,csa_tree_add_7_25_groupi_n_153);
  not csa_tree_add_7_25_groupi_drc_bufs24180(csa_tree_add_7_25_groupi_n_154 ,csa_tree_add_7_25_groupi_n_153);
  not csa_tree_add_7_25_groupi_drc_bufs24181(csa_tree_add_7_25_groupi_n_153 ,csa_tree_add_7_25_groupi_n_5864);
  not csa_tree_add_7_25_groupi_drc_bufs24183(csa_tree_add_7_25_groupi_n_152 ,csa_tree_add_7_25_groupi_n_151);
  not csa_tree_add_7_25_groupi_drc_bufs24185(csa_tree_add_7_25_groupi_n_151 ,csa_tree_add_7_25_groupi_n_1922);
  not csa_tree_add_7_25_groupi_drc_bufs24187(csa_tree_add_7_25_groupi_n_150 ,csa_tree_add_7_25_groupi_n_149);
  not csa_tree_add_7_25_groupi_drc_bufs24189(csa_tree_add_7_25_groupi_n_149 ,csa_tree_add_7_25_groupi_n_1858);
  not csa_tree_add_7_25_groupi_drc_bufs24191(csa_tree_add_7_25_groupi_n_148 ,csa_tree_add_7_25_groupi_n_147);
  not csa_tree_add_7_25_groupi_drc_bufs24193(csa_tree_add_7_25_groupi_n_147 ,csa_tree_add_7_25_groupi_n_1825);
  not csa_tree_add_7_25_groupi_drc_bufs24195(csa_tree_add_7_25_groupi_n_146 ,csa_tree_add_7_25_groupi_n_2317);
  not csa_tree_add_7_25_groupi_drc_bufs24197(csa_tree_add_7_25_groupi_n_2317 ,csa_tree_add_7_25_groupi_n_2743);
  not csa_tree_add_7_25_groupi_drc_bufs24199(csa_tree_add_7_25_groupi_n_145 ,csa_tree_add_7_25_groupi_n_144);
  not csa_tree_add_7_25_groupi_drc_bufs24201(csa_tree_add_7_25_groupi_n_144 ,csa_tree_add_7_25_groupi_n_1862);
  not csa_tree_add_7_25_groupi_drc_bufs24203(csa_tree_add_7_25_groupi_n_143 ,csa_tree_add_7_25_groupi_n_142);
  not csa_tree_add_7_25_groupi_drc_bufs24205(csa_tree_add_7_25_groupi_n_142 ,csa_tree_add_7_25_groupi_n_1867);
  not csa_tree_add_7_25_groupi_drc_bufs24207(csa_tree_add_7_25_groupi_n_141 ,csa_tree_add_7_25_groupi_n_140);
  not csa_tree_add_7_25_groupi_drc_bufs24209(csa_tree_add_7_25_groupi_n_140 ,csa_tree_add_7_25_groupi_n_1831);
  not csa_tree_add_7_25_groupi_drc_bufs24211(csa_tree_add_7_25_groupi_n_139 ,csa_tree_add_7_25_groupi_n_138);
  not csa_tree_add_7_25_groupi_drc_bufs24213(csa_tree_add_7_25_groupi_n_138 ,csa_tree_add_7_25_groupi_n_1910);
  not csa_tree_add_7_25_groupi_drc_bufs24215(csa_tree_add_7_25_groupi_n_137 ,csa_tree_add_7_25_groupi_n_2314);
  not csa_tree_add_7_25_groupi_drc_bufs24217(csa_tree_add_7_25_groupi_n_2314 ,csa_tree_add_7_25_groupi_n_2739);
  not csa_tree_add_7_25_groupi_drc_bufs24219(csa_tree_add_7_25_groupi_n_136 ,csa_tree_add_7_25_groupi_n_135);
  not csa_tree_add_7_25_groupi_drc_bufs24221(csa_tree_add_7_25_groupi_n_135 ,csa_tree_add_7_25_groupi_n_1852);
  not csa_tree_add_7_25_groupi_drc_bufs24223(csa_tree_add_7_25_groupi_n_134 ,csa_tree_add_7_25_groupi_n_133);
  not csa_tree_add_7_25_groupi_drc_bufs24225(csa_tree_add_7_25_groupi_n_133 ,csa_tree_add_7_25_groupi_n_1907);
  not csa_tree_add_7_25_groupi_drc_bufs24227(csa_tree_add_7_25_groupi_n_132 ,csa_tree_add_7_25_groupi_n_131);
  not csa_tree_add_7_25_groupi_drc_bufs24229(csa_tree_add_7_25_groupi_n_131 ,csa_tree_add_7_25_groupi_n_1846);
  not csa_tree_add_7_25_groupi_drc_bufs24231(csa_tree_add_7_25_groupi_n_130 ,csa_tree_add_7_25_groupi_n_2320);
  not csa_tree_add_7_25_groupi_drc_bufs24233(csa_tree_add_7_25_groupi_n_2320 ,csa_tree_add_7_25_groupi_n_2747);
  not csa_tree_add_7_25_groupi_drc_bufs24235(csa_tree_add_7_25_groupi_n_129 ,csa_tree_add_7_25_groupi_n_128);
  not csa_tree_add_7_25_groupi_drc_bufs24237(csa_tree_add_7_25_groupi_n_128 ,csa_tree_add_7_25_groupi_n_1849);
  not csa_tree_add_7_25_groupi_drc_bufs24239(csa_tree_add_7_25_groupi_n_127 ,csa_tree_add_7_25_groupi_n_2323);
  not csa_tree_add_7_25_groupi_drc_bufs24241(csa_tree_add_7_25_groupi_n_2323 ,csa_tree_add_7_25_groupi_n_2751);
  not csa_tree_add_7_25_groupi_drc_bufs24243(csa_tree_add_7_25_groupi_n_126 ,csa_tree_add_7_25_groupi_n_125);
  not csa_tree_add_7_25_groupi_drc_bufs24245(csa_tree_add_7_25_groupi_n_125 ,csa_tree_add_7_25_groupi_n_1925);
  not csa_tree_add_7_25_groupi_drc_bufs24247(csa_tree_add_7_25_groupi_n_124 ,csa_tree_add_7_25_groupi_n_123);
  not csa_tree_add_7_25_groupi_drc_bufs24249(csa_tree_add_7_25_groupi_n_123 ,csa_tree_add_7_25_groupi_n_1799);
  not csa_tree_add_7_25_groupi_drc_bufs24251(csa_tree_add_7_25_groupi_n_122 ,csa_tree_add_7_25_groupi_n_121);
  not csa_tree_add_7_25_groupi_drc_bufs24253(csa_tree_add_7_25_groupi_n_121 ,csa_tree_add_7_25_groupi_n_1901);
  not csa_tree_add_7_25_groupi_drc_bufs24255(csa_tree_add_7_25_groupi_n_120 ,csa_tree_add_7_25_groupi_n_118);
  not csa_tree_add_7_25_groupi_drc_bufs24256(csa_tree_add_7_25_groupi_n_119 ,csa_tree_add_7_25_groupi_n_118);
  not csa_tree_add_7_25_groupi_drc_bufs24257(csa_tree_add_7_25_groupi_n_118 ,csa_tree_add_7_25_groupi_n_2687);
  not csa_tree_add_7_25_groupi_drc_bufs24259(csa_tree_add_7_25_groupi_n_117 ,csa_tree_add_7_25_groupi_n_116);
  not csa_tree_add_7_25_groupi_drc_bufs24261(csa_tree_add_7_25_groupi_n_116 ,csa_tree_add_7_25_groupi_n_1919);
  not csa_tree_add_7_25_groupi_drc_bufs24263(csa_tree_add_7_25_groupi_n_115 ,csa_tree_add_7_25_groupi_n_113);
  not csa_tree_add_7_25_groupi_drc_bufs24264(csa_tree_add_7_25_groupi_n_114 ,csa_tree_add_7_25_groupi_n_113);
  not csa_tree_add_7_25_groupi_drc_bufs24265(csa_tree_add_7_25_groupi_n_113 ,csa_tree_add_7_25_groupi_n_1955);
  not csa_tree_add_7_25_groupi_drc_bufs24267(csa_tree_add_7_25_groupi_n_112 ,csa_tree_add_7_25_groupi_n_111);
  not csa_tree_add_7_25_groupi_drc_bufs24269(csa_tree_add_7_25_groupi_n_111 ,csa_tree_add_7_25_groupi_n_1087);
  not csa_tree_add_7_25_groupi_drc_bufs24271(csa_tree_add_7_25_groupi_n_110 ,csa_tree_add_7_25_groupi_n_109);
  not csa_tree_add_7_25_groupi_drc_bufs24273(csa_tree_add_7_25_groupi_n_109 ,csa_tree_add_7_25_groupi_n_1081);
  not csa_tree_add_7_25_groupi_drc_bufs24275(csa_tree_add_7_25_groupi_n_108 ,csa_tree_add_7_25_groupi_n_107);
  not csa_tree_add_7_25_groupi_drc_bufs24277(csa_tree_add_7_25_groupi_n_107 ,csa_tree_add_7_25_groupi_n_1069);
  not csa_tree_add_7_25_groupi_drc_bufs24279(csa_tree_add_7_25_groupi_n_106 ,csa_tree_add_7_25_groupi_n_105);
  not csa_tree_add_7_25_groupi_drc_bufs24281(csa_tree_add_7_25_groupi_n_105 ,csa_tree_add_7_25_groupi_n_1045);
  not csa_tree_add_7_25_groupi_drc_bufs24283(csa_tree_add_7_25_groupi_n_104 ,csa_tree_add_7_25_groupi_n_103);
  not csa_tree_add_7_25_groupi_drc_bufs24285(csa_tree_add_7_25_groupi_n_103 ,csa_tree_add_7_25_groupi_n_997);
  not csa_tree_add_7_25_groupi_drc_bufs24287(csa_tree_add_7_25_groupi_n_102 ,csa_tree_add_7_25_groupi_n_100);
  not csa_tree_add_7_25_groupi_drc_bufs24288(csa_tree_add_7_25_groupi_n_101 ,csa_tree_add_7_25_groupi_n_100);
  not csa_tree_add_7_25_groupi_drc_bufs24289(csa_tree_add_7_25_groupi_n_100 ,csa_tree_add_7_25_groupi_n_1952);
  not csa_tree_add_7_25_groupi_drc_bufs24291(csa_tree_add_7_25_groupi_n_99 ,csa_tree_add_7_25_groupi_n_98);
  not csa_tree_add_7_25_groupi_drc_bufs24293(csa_tree_add_7_25_groupi_n_98 ,csa_tree_add_7_25_groupi_n_1042);
  not csa_tree_add_7_25_groupi_drc_bufs24295(csa_tree_add_7_25_groupi_n_97 ,csa_tree_add_7_25_groupi_n_96);
  not csa_tree_add_7_25_groupi_drc_bufs24297(csa_tree_add_7_25_groupi_n_96 ,csa_tree_add_7_25_groupi_n_992);
  not csa_tree_add_7_25_groupi_drc_bufs24299(csa_tree_add_7_25_groupi_n_95 ,csa_tree_add_7_25_groupi_n_93);
  not csa_tree_add_7_25_groupi_drc_bufs24300(csa_tree_add_7_25_groupi_n_94 ,csa_tree_add_7_25_groupi_n_93);
  not csa_tree_add_7_25_groupi_drc_bufs24301(csa_tree_add_7_25_groupi_n_93 ,csa_tree_add_7_25_groupi_n_1949);
  not csa_tree_add_7_25_groupi_drc_bufs24303(csa_tree_add_7_25_groupi_n_92 ,csa_tree_add_7_25_groupi_n_91);
  not csa_tree_add_7_25_groupi_drc_bufs24305(csa_tree_add_7_25_groupi_n_91 ,csa_tree_add_7_25_groupi_n_1066);
  not csa_tree_add_7_25_groupi_drc_bufs24307(csa_tree_add_7_25_groupi_n_90 ,csa_tree_add_7_25_groupi_n_89);
  not csa_tree_add_7_25_groupi_drc_bufs24309(csa_tree_add_7_25_groupi_n_89 ,csa_tree_add_7_25_groupi_n_1039);
  not csa_tree_add_7_25_groupi_drc_bufs24311(csa_tree_add_7_25_groupi_n_88 ,csa_tree_add_7_25_groupi_n_87);
  not csa_tree_add_7_25_groupi_drc_bufs24313(csa_tree_add_7_25_groupi_n_87 ,csa_tree_add_7_25_groupi_n_1036);
  not csa_tree_add_7_25_groupi_drc_bufs24315(csa_tree_add_7_25_groupi_n_86 ,csa_tree_add_7_25_groupi_n_85);
  not csa_tree_add_7_25_groupi_drc_bufs24317(csa_tree_add_7_25_groupi_n_85 ,csa_tree_add_7_25_groupi_n_1078);
  not csa_tree_add_7_25_groupi_drc_bufs24319(csa_tree_add_7_25_groupi_n_84 ,csa_tree_add_7_25_groupi_n_83);
  not csa_tree_add_7_25_groupi_drc_bufs24321(csa_tree_add_7_25_groupi_n_83 ,csa_tree_add_7_25_groupi_n_1063);
  not csa_tree_add_7_25_groupi_drc_bufs24323(csa_tree_add_7_25_groupi_n_82 ,csa_tree_add_7_25_groupi_n_81);
  not csa_tree_add_7_25_groupi_drc_bufs24325(csa_tree_add_7_25_groupi_n_81 ,csa_tree_add_7_25_groupi_n_1033);
  not csa_tree_add_7_25_groupi_drc_bufs24327(csa_tree_add_7_25_groupi_n_80 ,csa_tree_add_7_25_groupi_n_79);
  not csa_tree_add_7_25_groupi_drc_bufs24329(csa_tree_add_7_25_groupi_n_79 ,csa_tree_add_7_25_groupi_n_1030);
  not csa_tree_add_7_25_groupi_drc_bufs24331(csa_tree_add_7_25_groupi_n_78 ,csa_tree_add_7_25_groupi_n_77);
  not csa_tree_add_7_25_groupi_drc_bufs24333(csa_tree_add_7_25_groupi_n_77 ,csa_tree_add_7_25_groupi_n_1060);
  not csa_tree_add_7_25_groupi_drc_bufs24335(csa_tree_add_7_25_groupi_n_76 ,csa_tree_add_7_25_groupi_n_75);
  not csa_tree_add_7_25_groupi_drc_bufs24337(csa_tree_add_7_25_groupi_n_75 ,csa_tree_add_7_25_groupi_n_1027);
  not csa_tree_add_7_25_groupi_drc_bufs24339(csa_tree_add_7_25_groupi_n_74 ,csa_tree_add_7_25_groupi_n_73);
  not csa_tree_add_7_25_groupi_drc_bufs24341(csa_tree_add_7_25_groupi_n_73 ,csa_tree_add_7_25_groupi_n_1024);
  not csa_tree_add_7_25_groupi_drc_bufs24343(csa_tree_add_7_25_groupi_n_72 ,csa_tree_add_7_25_groupi_n_71);
  not csa_tree_add_7_25_groupi_drc_bufs24345(csa_tree_add_7_25_groupi_n_71 ,csa_tree_add_7_25_groupi_n_1084);
  not csa_tree_add_7_25_groupi_drc_bufs24347(csa_tree_add_7_25_groupi_n_70 ,csa_tree_add_7_25_groupi_n_69);
  not csa_tree_add_7_25_groupi_drc_bufs24349(csa_tree_add_7_25_groupi_n_69 ,csa_tree_add_7_25_groupi_n_1075);
  not csa_tree_add_7_25_groupi_drc_bufs24351(csa_tree_add_7_25_groupi_n_68 ,csa_tree_add_7_25_groupi_n_67);
  not csa_tree_add_7_25_groupi_drc_bufs24353(csa_tree_add_7_25_groupi_n_67 ,csa_tree_add_7_25_groupi_n_1057);
  not csa_tree_add_7_25_groupi_drc_bufs24355(csa_tree_add_7_25_groupi_n_66 ,csa_tree_add_7_25_groupi_n_65);
  not csa_tree_add_7_25_groupi_drc_bufs24357(csa_tree_add_7_25_groupi_n_65 ,csa_tree_add_7_25_groupi_n_1000);
  not csa_tree_add_7_25_groupi_drc_bufs24359(csa_tree_add_7_25_groupi_n_64 ,csa_tree_add_7_25_groupi_n_63);
  not csa_tree_add_7_25_groupi_drc_bufs24361(csa_tree_add_7_25_groupi_n_63 ,csa_tree_add_7_25_groupi_n_1003);
  not csa_tree_add_7_25_groupi_drc_bufs24363(csa_tree_add_7_25_groupi_n_62 ,csa_tree_add_7_25_groupi_n_61);
  not csa_tree_add_7_25_groupi_drc_bufs24365(csa_tree_add_7_25_groupi_n_61 ,csa_tree_add_7_25_groupi_n_1006);
  not csa_tree_add_7_25_groupi_drc_bufs24367(csa_tree_add_7_25_groupi_n_60 ,csa_tree_add_7_25_groupi_n_59);
  not csa_tree_add_7_25_groupi_drc_bufs24369(csa_tree_add_7_25_groupi_n_59 ,csa_tree_add_7_25_groupi_n_1009);
  not csa_tree_add_7_25_groupi_drc_bufs24371(csa_tree_add_7_25_groupi_n_58 ,csa_tree_add_7_25_groupi_n_57);
  not csa_tree_add_7_25_groupi_drc_bufs24373(csa_tree_add_7_25_groupi_n_57 ,csa_tree_add_7_25_groupi_n_1012);
  not csa_tree_add_7_25_groupi_drc_bufs24375(csa_tree_add_7_25_groupi_n_56 ,csa_tree_add_7_25_groupi_n_55);
  not csa_tree_add_7_25_groupi_drc_bufs24377(csa_tree_add_7_25_groupi_n_55 ,csa_tree_add_7_25_groupi_n_1015);
  not csa_tree_add_7_25_groupi_drc_bufs24379(csa_tree_add_7_25_groupi_n_54 ,csa_tree_add_7_25_groupi_n_53);
  not csa_tree_add_7_25_groupi_drc_bufs24381(csa_tree_add_7_25_groupi_n_53 ,csa_tree_add_7_25_groupi_n_1021);
  not csa_tree_add_7_25_groupi_drc_bufs24383(csa_tree_add_7_25_groupi_n_52 ,csa_tree_add_7_25_groupi_n_51);
  not csa_tree_add_7_25_groupi_drc_bufs24385(csa_tree_add_7_25_groupi_n_51 ,csa_tree_add_7_25_groupi_n_1018);
  not csa_tree_add_7_25_groupi_drc_bufs24387(csa_tree_add_7_25_groupi_n_50 ,csa_tree_add_7_25_groupi_n_49);
  not csa_tree_add_7_25_groupi_drc_bufs24389(csa_tree_add_7_25_groupi_n_49 ,csa_tree_add_7_25_groupi_n_1054);
  not csa_tree_add_7_25_groupi_drc_bufs24391(csa_tree_add_7_25_groupi_n_48 ,csa_tree_add_7_25_groupi_n_47);
  not csa_tree_add_7_25_groupi_drc_bufs24393(csa_tree_add_7_25_groupi_n_47 ,csa_tree_add_7_25_groupi_n_1072);
  not csa_tree_add_7_25_groupi_drc_bufs24395(csa_tree_add_7_25_groupi_n_46 ,csa_tree_add_7_25_groupi_n_45);
  not csa_tree_add_7_25_groupi_drc_bufs24397(csa_tree_add_7_25_groupi_n_45 ,csa_tree_add_7_25_groupi_n_1051);
  not csa_tree_add_7_25_groupi_drc_bufs24399(csa_tree_add_7_25_groupi_n_44 ,csa_tree_add_7_25_groupi_n_43);
  not csa_tree_add_7_25_groupi_drc_bufs24401(csa_tree_add_7_25_groupi_n_43 ,csa_tree_add_7_25_groupi_n_1048);
  not csa_tree_add_7_25_groupi_drc_bufs24403(csa_tree_add_7_25_groupi_n_42 ,csa_tree_add_7_25_groupi_n_41);
  not csa_tree_add_7_25_groupi_drc_bufs24405(csa_tree_add_7_25_groupi_n_41 ,csa_tree_add_7_25_groupi_n_942);
  not csa_tree_add_7_25_groupi_drc_bufs24408(csa_tree_add_7_25_groupi_n_40 ,csa_tree_add_7_25_groupi_n_39);
  not csa_tree_add_7_25_groupi_drc_bufs24409(csa_tree_add_7_25_groupi_n_39 ,csa_tree_add_7_25_groupi_n_956);
  not csa_tree_add_7_25_groupi_drc_bufs24412(csa_tree_add_7_25_groupi_n_38 ,csa_tree_add_7_25_groupi_n_37);
  not csa_tree_add_7_25_groupi_drc_bufs24413(csa_tree_add_7_25_groupi_n_37 ,csa_tree_add_7_25_groupi_n_950);
  not csa_tree_add_7_25_groupi_drc_bufs24416(csa_tree_add_7_25_groupi_n_36 ,csa_tree_add_7_25_groupi_n_35);
  not csa_tree_add_7_25_groupi_drc_bufs24417(csa_tree_add_7_25_groupi_n_35 ,csa_tree_add_7_25_groupi_n_953);
  not csa_tree_add_7_25_groupi_drc_bufs24420(csa_tree_add_7_25_groupi_n_34 ,csa_tree_add_7_25_groupi_n_33);
  not csa_tree_add_7_25_groupi_drc_bufs24421(csa_tree_add_7_25_groupi_n_33 ,csa_tree_add_7_25_groupi_n_977);
  not csa_tree_add_7_25_groupi_drc_bufs24424(csa_tree_add_7_25_groupi_n_32 ,csa_tree_add_7_25_groupi_n_31);
  not csa_tree_add_7_25_groupi_drc_bufs24425(csa_tree_add_7_25_groupi_n_31 ,csa_tree_add_7_25_groupi_n_980);
  not csa_tree_add_7_25_groupi_drc_bufs24428(csa_tree_add_7_25_groupi_n_30 ,csa_tree_add_7_25_groupi_n_29);
  not csa_tree_add_7_25_groupi_drc_bufs24429(csa_tree_add_7_25_groupi_n_29 ,csa_tree_add_7_25_groupi_n_939);
  not csa_tree_add_7_25_groupi_drc_bufs24432(csa_tree_add_7_25_groupi_n_28 ,csa_tree_add_7_25_groupi_n_27);
  not csa_tree_add_7_25_groupi_drc_bufs24433(csa_tree_add_7_25_groupi_n_27 ,csa_tree_add_7_25_groupi_n_936);
  not csa_tree_add_7_25_groupi_drc_bufs24436(csa_tree_add_7_25_groupi_n_26 ,csa_tree_add_7_25_groupi_n_25);
  not csa_tree_add_7_25_groupi_drc_bufs24437(csa_tree_add_7_25_groupi_n_25 ,csa_tree_add_7_25_groupi_n_983);
  not csa_tree_add_7_25_groupi_drc_bufs24440(csa_tree_add_7_25_groupi_n_24 ,csa_tree_add_7_25_groupi_n_23);
  not csa_tree_add_7_25_groupi_drc_bufs24441(csa_tree_add_7_25_groupi_n_23 ,csa_tree_add_7_25_groupi_n_974);
  not csa_tree_add_7_25_groupi_drc_bufs24444(csa_tree_add_7_25_groupi_n_22 ,csa_tree_add_7_25_groupi_n_21);
  not csa_tree_add_7_25_groupi_drc_bufs24445(csa_tree_add_7_25_groupi_n_21 ,csa_tree_add_7_25_groupi_n_962);
  not csa_tree_add_7_25_groupi_drc_bufs24448(csa_tree_add_7_25_groupi_n_20 ,csa_tree_add_7_25_groupi_n_19);
  not csa_tree_add_7_25_groupi_drc_bufs24449(csa_tree_add_7_25_groupi_n_19 ,csa_tree_add_7_25_groupi_n_965);
  not csa_tree_add_7_25_groupi_drc_bufs24452(csa_tree_add_7_25_groupi_n_18 ,csa_tree_add_7_25_groupi_n_17);
  not csa_tree_add_7_25_groupi_drc_bufs24453(csa_tree_add_7_25_groupi_n_17 ,csa_tree_add_7_25_groupi_n_971);
  not csa_tree_add_7_25_groupi_drc_bufs24456(csa_tree_add_7_25_groupi_n_16 ,csa_tree_add_7_25_groupi_n_15);
  not csa_tree_add_7_25_groupi_drc_bufs24457(csa_tree_add_7_25_groupi_n_15 ,csa_tree_add_7_25_groupi_n_944);
  not csa_tree_add_7_25_groupi_drc_bufs24460(csa_tree_add_7_25_groupi_n_14 ,csa_tree_add_7_25_groupi_n_13);
  not csa_tree_add_7_25_groupi_drc_bufs24461(csa_tree_add_7_25_groupi_n_13 ,csa_tree_add_7_25_groupi_n_986);
  not csa_tree_add_7_25_groupi_drc_bufs24464(csa_tree_add_7_25_groupi_n_12 ,csa_tree_add_7_25_groupi_n_11);
  not csa_tree_add_7_25_groupi_drc_bufs24465(csa_tree_add_7_25_groupi_n_11 ,csa_tree_add_7_25_groupi_n_947);
  not csa_tree_add_7_25_groupi_drc_bufs24468(csa_tree_add_7_25_groupi_n_10 ,csa_tree_add_7_25_groupi_n_9);
  not csa_tree_add_7_25_groupi_drc_bufs24469(csa_tree_add_7_25_groupi_n_9 ,csa_tree_add_7_25_groupi_n_968);
  not csa_tree_add_7_25_groupi_drc_bufs24472(csa_tree_add_7_25_groupi_n_8 ,csa_tree_add_7_25_groupi_n_7);
  not csa_tree_add_7_25_groupi_drc_bufs24473(csa_tree_add_7_25_groupi_n_7 ,csa_tree_add_7_25_groupi_n_959);
  xor csa_tree_add_7_25_groupi_g2(out2[38] ,csa_tree_add_7_25_groupi_n_7245 ,csa_tree_add_7_25_groupi_n_7212);
  xor csa_tree_add_7_25_groupi_g24475(out2[37] ,csa_tree_add_7_25_groupi_n_7243 ,csa_tree_add_7_25_groupi_n_7210);
  xor csa_tree_add_7_25_groupi_g24476(out2[35] ,csa_tree_add_7_25_groupi_n_7238 ,csa_tree_add_7_25_groupi_n_7209);
  xor csa_tree_add_7_25_groupi_g24477(out2[34] ,csa_tree_add_7_25_groupi_n_7236 ,csa_tree_add_7_25_groupi_n_7208);
  and csa_tree_add_7_25_groupi_g24478(csa_tree_add_7_25_groupi_n_2 ,csa_tree_add_7_25_groupi_n_267 ,csa_tree_add_7_25_groupi_n_1105);
  xor csa_tree_add_7_25_groupi_g24479(csa_tree_add_7_25_groupi_n_1 ,csa_tree_add_7_25_groupi_n_5077 ,csa_tree_add_7_25_groupi_n_1103);
  xor csa_tree_add_7_25_groupi_g24480(csa_tree_add_7_25_groupi_n_0 ,csa_tree_add_7_25_groupi_n_4774 ,csa_tree_add_7_25_groupi_n_1101);
  buf g24481(csa_tree_add_7_25_groupi_n_2660 ,csa_tree_add_7_25_groupi_n_2475);
endmodule
