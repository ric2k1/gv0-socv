module cmos_demo(input a, b, output [1:0] y);
assign y = a + b;
endmodule
