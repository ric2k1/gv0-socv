module top( n1 , n4 , n10 , n13 , n26 , n27 , n32 , n34 , n46 , n52 , n54 , n58 , n61 , n64 , n65 , n66 );
    input n1 , n4 , n10 , n13 , n27 , n32 , n46 , n58 , n61 , n64 , n65 , n66 ;
    output n26 , n34 , n52 , n54 ;
    wire n0 , n2 , n3 , n5 , n6 , n7 , n8 , n9 , n11 , n12 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n28 , n29 , n30 , n31 , n33 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n47 , n48 , n49 , n50 , n51 , n53 , n55 , n56 , n57 , n59 , n60 , n62 , n63 , n67 , n68 , n69 , n70 ;
assign n33 = ~n46;
assign n17 = n8 & n40;
assign n23 = ~(n14 ^ n64);
assign n47 = ~(n17 | n49);
assign n29 = n61 | n33;
assign n69 = ~(n19 | n36);
assign n34 = ~(n49 ^ n0);
assign n18 = ~(n40 | n8);
assign n7 = ~n58;
assign n16 = ~(n20 ^ n1);
assign n37 = ~n70;
assign n8 = ~(n70 ^ n44);
assign n53 = ~n24;
assign n40 = ~n27;
assign n14 = ~(n18 | n47);
assign n24 = n41 & n2;
assign n12 = ~(n48 | n69);
assign n35 = ~(n29 ^ n63);
assign n60 = ~n55;
assign n63 = n66 | n7;
assign n55 = n67 & n11;
assign n68 = n11 | n67;
assign n22 = n1 | n60;
assign n25 = ~(n57 | n12);
assign n19 = ~n53;
assign n51 = ~(n13 | n66);
assign n39 = ~(n25 ^ n50);
assign n41 = ~n13;
assign n50 = ~(n70 | n44);
assign n43 = ~(n39 ^ n23);
assign n38 = ~(n24 ^ n48);
assign n20 = n9 | n37;
assign n70 = n53 | n28;
assign n28 = ~n67;
assign n11 = ~n4;
assign n31 = ~n55;
assign n44 = ~(n36 ^ n38);
assign n9 = ~(n56 | n51);
assign n15 = n42 | n20;
assign n67 = n62 & n3;
assign n21 = n13 | n30;
assign n49 = n15 & n22;
assign n30 = ~n10;
assign n48 = n66 | n5;
assign n52 = ~(n59 ^ n43);
assign n0 = ~(n8 ^ n27);
assign n45 = ~(n6 ^ n21);
assign n54 = n60 & n68;
assign n57 = n36 & n19;
assign n5 = ~n65;
assign n62 = ~n61;
assign n3 = ~n66;
assign n2 = ~n32;
assign n56 = ~(n61 | n32);
assign n59 = ~(n35 ^ n45);
assign n26 = ~(n55 ^ n16);
assign n36 = n62 & n10;
assign n42 = n31 & n1;
assign n6 = ~(n32 | n5);
endmodule
