module top;
	rand const reg rx;
	const reg ry;
	rand reg rz;
	rand const integer ix;
	const integer iy;
	rand integer iz;
endmodule
