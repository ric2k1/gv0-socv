module a;
wire [3]x;
endmodule

