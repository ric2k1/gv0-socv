module top( n19 , n24 , n29 , n32 , n36 , n49 , n52 , n58 , n59 , n60 , n69 , n73 , n76 , n96 , n97 , n100 , n108 , n117 , n123 , n143 , n149 , n151 , n152 , n158 , n167 , n189 , n194 , n196 , n197 , n198 , n206 , n209 , n210 , n217 , n218 , n222 , n224 , n226 , n233 , n242 , n245 , n248 , n258 );
    input n19 , n24 , n32 , n36 , n49 , n52 , n58 , n59 , n60 , n69 , n73 , n96 , n97 , n100 , n108 , n117 , n123 , n143 , n149 , n151 , n158 , n167 , n189 , n196 , n197 , n198 , n206 , n209 , n210 , n217 , n218 , n222 , n226 , n233 , n242 , n258 ;
    output n29 , n76 , n152 , n194 , n224 , n245 , n248 ;
    wire n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n20 , n21 , n22 , n23 , n25 , n26 , n27 , n28 , n30 , n31 , n33 , n34 , n35 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n50 , n51 , n53 , n54 , n55 , n56 , n57 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n70 , n71 , n72 , n74 , n75 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n98 , n99 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n118 , n119 , n120 , n121 , n122 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n144 , n145 , n146 , n147 , n148 , n150 , n153 , n154 , n155 , n156 , n157 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n190 , n191 , n192 , n193 , n195 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n207 , n208 , n211 , n212 , n213 , n214 , n215 , n216 , n219 , n220 , n221 , n223 , n225 , n227 , n228 , n229 , n230 , n231 , n232 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n243 , n244 , n246 , n247 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n259 , n260 , n261 , n262 ;
assign n95 = ~(n29 ^ n40);
assign n43 = ~n218;
assign n141 = ~(n87 | n5);
assign n216 = n123 & n179;
assign n180 = n253 | n88;
assign n2 = n245 ^ n190;
assign n88 = ~n213;
assign n191 = n185 & n114;
assign n199 = n250 | n157;
assign n129 = n109 & n214;
assign n236 = n21 & n10;
assign n40 = ~n184;
assign n168 = n117 & n137;
assign n27 = n117;
assign n9 = ~(n220 | n42);
assign n7 = n129 | n34;
assign n41 = ~n168;
assign n257 = ~n210;
assign n70 = ~n197;
assign n156 = n150 & n141;
assign n173 = n68 | n11;
assign n223 = ~(n29 ^ n35);
assign n219 = n120 | n131;
assign n262 = n70 & n55;
assign n28 = ~n149;
assign n122 = n243 | n238;
assign n120 = n69 & n29;
assign n94 = n245 ^ n31;
assign n137 = ~n233;
assign n237 = ~n222;
assign n75 = n59 & n204;
assign n205 = n99 | n126;
assign n215 = n245 ^ n154;
assign n155 = n70 | n88;
assign n99 = n12 & n33;
assign n239 = ~(n145 | n234);
assign n111 = n28 | n49;
assign n104 = n163 & n208;
assign n224 = n85 | n56;
assign n193 = ~n190;
assign n175 = n192 | n20;
assign n0 = n223 | n215;
assign n47 = n204 | n72;
assign n102 = ~n209;
assign n170 = n149 & n202;
assign n203 = n3 | n46;
assign n183 = ~(n166 | n223);
assign n55 = ~(n93 | n68);
assign n246 = ~(n102 | n225);
assign n89 = ~(n195 | n95);
assign n184 = n100 & n64;
assign n166 = ~n123;
assign n110 = ~n79;
assign n153 = ~n117;
assign n34 = n44 & n105;
assign n234 = ~n18;
assign n61 = n65;
assign n82 = ~(n227 | n165);
assign n221 = ~n188;
assign n130 = n75 | n13;
assign n18 = n26 & n106;
assign n152 = n6 | n207;
assign n65 = n191 & n216;
assign n144 = n245 ^ n241;
assign n12 = n47 & n155;
assign n243 = ~(n164 | n212);
assign n150 = n128 | n69;
assign n211 = n122 | n30;
assign n86 = n188 | n110;
assign n6 = n99 | n112;
assign n78 = n100 & n25;
assign n83 = n128 | n136;
assign n192 = ~n19;
assign n42 = n225 | n228;
assign n79 = n186 & n71;
assign n53 = ~(n61 | n86);
assign n62 = n251 | n135;
assign n164 = n50 | n32;
assign n71 = n149 & n54;
assign n163 = n64 | n72;
assign n169 = ~n49;
assign n3 = n258 & n43;
assign n76 = ~(n17 | n63);
assign n101 = n43 | n72;
assign n136 = n198 & n194;
assign n4 = n245 ^ n178;
assign n20 = ~n194;
assign n67 = n77 & n180;
assign n204 = ~n151;
assign n85 = n99 | n188;
assign n35 = ~n46;
assign n29 = ~n156;
assign n248 = n171 | n205;
assign n148 = n188 | n236;
assign n107 = ~n170;
assign n31 = n237 & n51;
assign n252 = ~n194;
assign n146 = ~(n230 | n16);
assign n51 = ~(n28 | n200);
assign n1 = n257 | n45;
assign n244 = n80 | n146;
assign n124 = n202 | n45;
assign n250 = ~n158;
assign n231 = n245 ^ n34;
assign n213 = ~n15;
assign n45 = ~n38;
assign n17 = ~(n148 | n62);
assign n38 = ~n156;
assign n121 = n166 | n226;
assign n15 = n193 & n82;
assign n139 = n237 | n88;
assign n177 = n260 | n244;
assign n253 = ~n52;
assign n214 = ~(n50 | n39);
assign n93 = ~n59;
assign n112 = n159 & n239;
assign n109 = ~n189;
assign n178 = n250 & n127;
assign n21 = n1 & n199;
assign n77 = n91 | n72;
assign n57 = ~n75;
assign n13 = n209 & n91;
assign n235 = ~(n29 ^ n150);
assign n165 = n22 | n7;
assign n232 = ~n160;
assign n200 = ~(n29 ^ n107);
assign n174 = ~(n236 | n240);
assign n159 = ~(n188 | n236);
assign n14 = ~n60;
assign n128 = ~n73;
assign n181 = ~n242;
assign n72 = ~n38;
assign n81 = n99 | n27;
assign n254 = ~n206;
assign n125 = ~n96;
assign n256 = n245 ^ n129;
assign n5 = n203 | n116;
assign n132 = n209 & n8;
assign n154 = n254 & n183;
assign n176 = n128 | n198;
assign n80 = ~(n172 | n74);
assign n16 = n95 | n144;
assign n119 = ~n217;
assign n185 = n48 | n45;
assign n44 = ~n196;
assign n227 = n103 | n187;
assign n140 = n109 | n157;
assign n228 = n245 ^ n255;
assign n54 = n169 | n20;
assign n201 = n177 | n211;
assign n145 = n104 & n78;
assign n74 = n142 | n4;
assign n8 = n125 | n20;
assign n207 = n126 | n53;
assign n10 = n217 & n175;
assign n229 = ~n167;
assign n133 = ~n143;
assign n212 = n39 | n256;
assign n230 = n195 | n167;
assign n25 = n229 | n20;
assign n98 = ~(n29 ^ n41);
assign n171 = n188 | n145;
assign n247 = ~n65;
assign n238 = ~(n121 | n0);
assign n105 = ~(n153 | n98);
assign n113 = n261 | n252;
assign n103 = n255 | n178;
assign n249 = n160 | n184;
assign n106 = n258 & n113;
assign n179 = n134 | n252;
assign n116 = n170 | n168;
assign n225 = ~(n29 ^ n138);
assign n142 = ~(n29 ^ n232);
assign n63 = ~(n219 | n83);
assign n134 = ~n226;
assign n259 = ~n3;
assign n50 = ~n258;
assign n30 = n66 | n92;
assign n147 = n18 | n79;
assign n157 = ~n213;
assign n11 = n245 ^ n262;
assign n64 = ~n24;
assign n37 = n93 | n143;
assign n240 = n145 | n247;
assign n39 = ~(n29 ^ n259);
assign n245 = ~n15;
assign n115 = ~(n37 | n173);
assign n87 = n130 | n249;
assign n261 = ~n32;
assign n22 = n241 | n154;
assign n172 = n119 | n19;
assign n26 = n101 & n140;
assign n48 = ~n97;
assign n194 = n84 | n201;
assign n33 = n59 & n90;
assign n186 = n124 & n139;
assign n187 = n262 | n31;
assign n188 = n67 & n132;
assign n195 = ~n100;
assign n160 = n217 & n257;
assign n162 = n200 | n94;
assign n114 = n254 | n157;
assign n182 = ~(n128 | n235);
assign n220 = n102 | n96;
assign n92 = ~(n118 | n161);
assign n90 = n133 | n252;
assign n66 = ~(n111 | n162);
assign n91 = ~n108;
assign n84 = ~(n176 | n23);
assign n56 = n174 | n112;
assign n241 = n14 & n89;
assign n202 = ~n58;
assign n190 = n181 & n182;
assign n46 = n123 & n48;
assign n260 = n115 | n9;
assign n208 = n14 | n88;
assign n251 = n145 | n65;
assign n118 = n153 | n36;
assign n255 = n253 & n246;
assign n135 = n147 | n81;
assign n68 = ~(n29 ^ n57);
assign n161 = n98 | n231;
assign n138 = ~n13;
assign n23 = n235 | n2;
assign n131 = n242 & n245;
assign n126 = n221 & n236;
assign n127 = ~(n119 | n142);
endmodule
