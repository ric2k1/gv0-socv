module top(in1, in2, in3, out1, out2, out3, out4, out5, out6);
  input [30:0] in1;
  input [31:0] in2, in3;
  output [32:0] out1, out4;
  output out2, out3, out5, out6;
  wire [30:0] in1;
  wire [31:0] in2, in3;
  wire [32:0] out1, out4;
  wire out2, out3, out5, out6;
  wire w__1, w__2, w__3, w__4, w__5, w__6, w__7, w__8;
  wire w__9, w__10, w__11, w__12, w__13, w__14, w__15, w__16;
  wire w__17, w__18, w__19, w__20, w__21, w__22, w__23, w__24;
  wire w__25, w__26, w__27, w__28, w__29, w__30, w__31, w__32;
  wire w__33, w__34, w__35, w__36, w__37, w__38, w__39, w__40;
  wire w__41, w__42, w__43, w__44, w__45, w__46, w__47, w__48;
  wire w__49, w__50, w__51, w__52, w__53, w__54, w__55, w__56;
  wire w__57, w__58, w__59, w__60, w__61, w__62, w__63, w__64;
  wire w__65, w__66, w__67, w__68, w__69, w__70, w__71, w__72;
  wire w__73, w__74, w__75, w__76, w__77, w__78, w__79, w__80;
  wire w__81, w__82, w__83, w__84, w__85, w__86, w__87, w__88;
  wire w__89, w__90, w__91, w__92, w__93, w__94, w__95, w__96;
  wire w__97, w__98, w__99, w__100, w__101, w__102, w__103, w__104;
  wire w__105, w__106, w__107, w__108, w__109, w__110, w__111, w__112;
  wire w__113, w__114, w__115, w__116, w__117, w__118, w__119, w__120;
  wire w__121, w__122, w__123, w__124, w__125, w__126, w__127, w__128;
  wire w__129, w__130, w__131, w__132, w__133, w__134, w__135, w__136;
  wire w__137, w__138, w__139, w__140, w__141, w__142, w__143, w__144;
  wire w__145, w__146, w__147, w__148, w__149, w__150, w__151, w__152;
  wire w__153, w__154, w__155, w__156, w__157, w__158, w__159, w__160;
  wire w__161, w__162, w__163, w__164, w__165, w__166, w__167, w__168;
  wire w__169, w__170, w__171, w__172, w__173, w__174, w__175, w__176;
  wire w__177, w__178, w__179, w__180, w__181, w__182, w__183, w__184;
  wire w__185, w__186, w__187, w__188, w__189, w__190, w__191, w__192;
  wire w__193, w__194, w__195, w__196, w__197, w__198, w__199, w__200;
  wire w__201, w__202, w__203, w__204, w__205, w__206, w__207, w__208;
  wire w__209, w__210, w__211, w__212, w__213, w__214, w__215, w__216;
  wire w__217, w__218, w__219, w__220, w__221, w__222, w__223, w__224;
  wire w__225, w__226, w__227, w__228, w__229, w__230, w__231, w__232;
  wire w__233, w__234, w__235, w__236, w__237, w__238, w__239, w__240;
  wire w__241, w__242, w__243, w__244, w__245, w__246, w__247, w__248;
  wire w__249, w__250, w__251, w__252, w__253, w__254, w__255, w__256;
  wire w__257, w__258, w__259, w__260, w__261, w__262, w__263, w__264;
  wire w__265, w__266, w__267, w__268, w__269, w__270, w__271, w__272;
  wire w__273, w__274, w__275, w__276, w__277, w__278, w__279, w__280;
  wire w__281, w__282, w__283, w__284, w__285, w__286, w__287, w__288;
  wire w__289, w__290, w__291, w__292, w__293, w__294, w__295, w__296;
  wire w__297, w__298, w__299, w__300, w__301, w__302, w__303, w__304;
  wire w__305, w__306, w__307, w__308, w__309, w__310, w__311, w__312;
  wire w__313, w__314, w__315, w__316, w__317, w__318, w__319, w__320;
  wire w__321, w__322, w__323, w__324, w__325, w__326, w__327, w__328;
  wire w__329, w__330, w__331, w__332, w__333, w__334, w__335, w__336;
  wire w__337, w__338, w__339, w__340, w__341, w__342, w__343, w__344;
  wire w__345, w__346, w__347, w__348, w__349, w__350, w__351, w__352;
  wire w__353, w__354, w__355, w__356, w__357, w__358, w__359, w__360;
  wire w__361, w__362, w__363, w__364, w__365, w__366, w__367, w__368;
  wire w__369, w__370, w__371, w__372, w__373, w__374, w__375, w__376;
  wire w__377, w__378, w__379, w__380, w__381, w__382, w__383, w__384;
  wire w__385, w__386, w__387, w__388, w__389, w__390, w__391, w__392;
  wire w__393, w__394, w__395, w__396, w__397, w__398, w__399, w__400;
  wire w__401, w__402, w__403, w__404, w__405, w__406, w__407, w__408;
  wire w__409, w__410, w__411, w__412, w__413, w__414, w__415, w__416;
  wire w__417, w__418, w__419, w__420, w__421, w__422, w__423, w__424;
  wire w__425, w__426, w__427, w__428, w__429, w__430, w__431, w__432;
  wire w__433, w__434, w__435, w__436, w__437, w__438, w__439, w__440;
  wire w__441, w__442, w__443, w__444, w__445, w__446, w__447, w__448;
  wire w__449, w__450, w__451, w__452, w__453, w__454, w__455, w__456;
  wire w__457, w__458, w__459, w__460, w__461, w__462, w__463, w__464;
  wire w__465, w__466, w__467, w__468, w__469, w__470, w__471, w__472;
  wire w__473, w__474, w__475, w__476, w__477, w__478, w__479, w__480;
  wire w__481, w__482, w__483, w__484, w__485, w__486, w__487, w__488;
  wire w__489, w__490, w__491, w__492, w__493, w__494, w__495, w__496;
  wire w__497, w__498, w__499, w__500, w__501, w__502, w__503, w__504;
  wire w__505, w__506, w__507, w__508, w__509, w__510, w__511, w__512;
  wire w__513, w__514, w__515, w__516, w__517, w__518, w__519, w__520;
  wire w__521, w__522, w__523, w__524, w__525, w__526, w__527, w__528;
  wire w__529, w__530, w__531, w__532, w__533, w__534, w__535, w__536;
  wire w__537, w__538, w__539, w__540, w__541, w__542, w__543, w__544;
  wire w__545, w__546, w__547, w__548, w__549, w__550, w__551, w__552;
  wire w__553, w__554, w__555, w__556, w__557, w__558, w__559, w__560;
  wire w__561, w__562, w__563, w__564, w__565, w__566, w__567, w__568;
  wire w__569, w__570, w__571, w__572, w__573, w__574, w__575, w__576;
  wire w__577, w__578, w__579, w__580, w__581, w__582, w__583, w__584;
  wire w__585, w__586, w__587, w__588, w__589, w__590, w__591, w__592;
  wire w__593, w__594, w__595, w__596, w__597, w__598, w__599, w__600;
  wire w__601, w__602, w__603, w__604, w__605, w__606, w__607, w__608;
  wire w__609, w__610, w__611, w__612, w__613, w__614, w__615, w__616;
  wire w__617, w__618, w__619, w__620, w__621, w__622, w__623, w__624;
  wire w__625, w__626, w__627, w__628, w__629, w__630, w__631, w__632;
  wire w__633, w__634, w__635, w__636, w__637, w__638, w__639, w__640;
  wire w__641, w__642, w__643, w__644, w__645, w__646, w__647, w__648;
  wire w__649, w__650, w__651, w__652, w__653, w__654, w__655, w__656;
  wire w__657, w__658, w__659, w__660, w__661, w__662, w__663, w__664;
  wire w__665, w__666, w__667, w__668, w__669, w__670, w__671, w__672;
  wire w__673, w__674, w__675, w__676, w__677, w__678, w__679, w__680;
  wire w__681, w__682, w__683, w__684, w__685, w__686, w__687, w__688;
  wire w__689, w__690, w__691, w__692, w__693, w__694, w__695, w__696;
  wire w__697, w__698, w__699, w__700, w__701, w__702, w__703, w__704;
  wire w__705, w__706, w__707, w__708, w__709, w__710, w__711, w__712;
  wire w__713, w__714, w__715, w__716, w__717, w__718, w__719, w__720;
  wire w__721, w__722, w__723, w__724, w__725, w__726, w__727, w__728;
  wire w__729, w__730, w__731, w__732, w__733, w__734, w__735, w__736;
  wire w__737, w__738, w__739, w__740, w__741, w__742, w__743, w__744;
  wire w__745, w__746, w__747, w__748, w__749, w__750, w__751, w__752;
  wire w__753, w__754, w__755, w__756, w__757, w__758, w__759, w__760;
  wire w__761, w__762, w__763, w__764, w__765, w__766, w__767, w__768;
  wire w__769, w__770, w__771, w__772, w__773, w__774, w__775, w__776;
  wire w__777, w__778, w__779, w__780, w__781, w__782, w__783, w__784;
  wire w__785, w__786, w__787, w__788, w__789, w__790, w__791, w__792;
  wire w__793, w__794, w__795, w__796, w__797, w__798, w__799, w__800;
  wire w__801, w__802, w__803, w__804, w__805, w__806, w__807, w__808;
  wire w__809, w__810, w__811, w__812, w__813, w__814, w__815, w__816;
  wire w__817, w__818, w__819, w__820, w__821, w__822, w__823, w__824;
  wire w__825, w__826, w__827, w__828, w__829, w__830, w__831, w__832;
  wire w__833, w__834, w__835, w__836, w__837, w__838, w__839, w__840;
  wire w__841, w__842, w__843, w__844, w__845, w__846, w__847, w__848;
  wire w__849, w__850, w__851, w__852, w__853, w__854, w__855, w__856;
  wire w__857, w__858, w__859, w__860, w__861, w__862, w__863, w__864;
  wire w__865, w__866, w__867, w__868;
  not g__1(w__264 ,in1[1]);
  xnor g__2(w__293 ,w__87 ,in1[30]);
  and g__3(w__294 ,in1[30] ,w__86);
  and g__4(w__292 ,w__85 ,w__87);
  not g__5(w__86 ,w__87);
  or g__6(w__87 ,w__15 ,w__84);
  or g__7(w__85 ,in1[29] ,w__83);
  xnor g__8(w__291 ,w__81 ,in1[28]);
  not g__9(w__84 ,w__83);
  and g__10(w__83 ,in1[28] ,w__80);
  and g__11(w__290 ,w__82 ,w__81);
  or g__12(w__82 ,in1[27] ,w__78);
  not g__13(w__80 ,w__81);
  or g__14(w__81 ,w__5 ,w__79);
  xnor g__15(w__289 ,w__76 ,in1[26]);
  not g__16(w__79 ,w__78);
  and g__17(w__78 ,in1[26] ,w__75);
  and g__18(w__288 ,w__77 ,w__76);
  or g__19(w__77 ,in1[25] ,w__73);
  not g__20(w__75 ,w__76);
  or g__21(w__76 ,w__3 ,w__74);
  xnor g__22(w__287 ,w__71 ,in1[24]);
  not g__23(w__74 ,w__73);
  and g__24(w__73 ,in1[24] ,w__70);
  and g__25(w__286 ,w__72 ,w__71);
  or g__26(w__72 ,in1[23] ,w__68);
  not g__27(w__70 ,w__71);
  or g__28(w__71 ,w__8 ,w__69);
  xnor g__29(w__285 ,w__67 ,in1[22]);
  not g__30(w__69 ,w__68);
  and g__31(w__68 ,in1[22] ,w__66);
  and g__32(w__284 ,w__65 ,w__67);
  not g__33(w__66 ,w__67);
  or g__34(w__67 ,w__4 ,w__64);
  or g__35(w__65 ,in1[21] ,w__63);
  xnor g__36(w__283 ,w__61 ,in1[20]);
  not g__37(w__64 ,w__63);
  and g__38(w__63 ,in1[20] ,w__60);
  and g__39(w__282 ,w__62 ,w__61);
  or g__40(w__62 ,in1[19] ,w__58);
  not g__41(w__60 ,w__61);
  or g__42(w__61 ,w__11 ,w__59);
  xnor g__43(w__281 ,w__56 ,in1[18]);
  not g__44(w__59 ,w__58);
  and g__45(w__58 ,in1[18] ,w__55);
  and g__46(w__280 ,w__57 ,w__56);
  or g__47(w__57 ,in1[17] ,w__53);
  not g__48(w__55 ,w__56);
  or g__49(w__56 ,w__16 ,w__54);
  xnor g__50(w__279 ,w__51 ,in1[16]);
  not g__51(w__54 ,w__53);
  and g__52(w__53 ,in1[16] ,w__50);
  and g__53(w__278 ,w__52 ,w__51);
  or g__54(w__52 ,in1[15] ,w__48);
  not g__55(w__50 ,w__51);
  or g__56(w__51 ,w__2 ,w__49);
  xnor g__57(w__277 ,w__47 ,in1[14]);
  not g__58(w__49 ,w__48);
  and g__59(w__48 ,in1[14] ,w__46);
  and g__60(w__276 ,w__45 ,w__47);
  not g__61(w__46 ,w__47);
  or g__62(w__47 ,w__9 ,w__44);
  or g__63(w__45 ,in1[13] ,w__43);
  xnor g__64(w__275 ,w__42 ,in1[12]);
  not g__65(w__44 ,w__43);
  and g__66(w__43 ,in1[12] ,w__41);
  and g__67(w__274 ,w__40 ,w__42);
  not g__68(w__41 ,w__42);
  or g__69(w__42 ,w__14 ,w__39);
  or g__70(w__40 ,in1[11] ,w__38);
  xnor g__71(w__273 ,w__36 ,in1[10]);
  not g__72(w__39 ,w__38);
  and g__73(w__38 ,in1[10] ,w__35);
  and g__74(w__272 ,w__37 ,w__36);
  or g__75(w__37 ,in1[9] ,w__33);
  not g__76(w__35 ,w__36);
  or g__77(w__36 ,w__1 ,w__34);
  xnor g__78(w__271 ,w__31 ,in1[8]);
  not g__79(w__34 ,w__33);
  and g__80(w__33 ,in1[8] ,w__30);
  and g__81(w__270 ,w__32 ,w__31);
  or g__82(w__32 ,in1[7] ,w__28);
  not g__83(w__30 ,w__31);
  or g__84(w__31 ,w__7 ,w__29);
  xnor g__85(w__269 ,w__26 ,in1[6]);
  not g__86(w__29 ,w__28);
  and g__87(w__28 ,in1[6] ,w__25);
  and g__88(w__268 ,w__27 ,w__26);
  or g__89(w__27 ,in1[5] ,w__23);
  not g__90(w__25 ,w__26);
  or g__91(w__26 ,w__13 ,w__24);
  xnor g__92(w__267 ,w__22 ,in1[4]);
  not g__93(w__24 ,w__23);
  and g__94(w__23 ,in1[4] ,w__21);
  and g__95(w__266 ,w__20 ,w__22);
  not g__96(w__21 ,w__22);
  or g__97(w__22 ,w__6 ,w__19);
  or g__98(w__20 ,in1[3] ,w__18);
  and g__99(w__265 ,w__19 ,w__17);
  not g__100(w__18 ,w__19);
  or g__101(w__19 ,w__10 ,w__12);
  or g__102(w__17 ,in1[2] ,in1[1]);
  not g__103(w__16 ,in1[17]);
  not g__104(w__15 ,in1[29]);
  not g__105(w__14 ,in1[11]);
  not g__106(w__13 ,in1[5]);
  not g__107(w__12 ,in1[1]);
  not g__108(w__11 ,in1[19]);
  not g__109(w__10 ,in1[2]);
  not g__110(w__9 ,in1[13]);
  not g__111(w__8 ,in1[23]);
  not g__112(w__7 ,in1[7]);
  not g__113(w__6 ,in1[3]);
  not g__114(w__5 ,in1[27]);
  not g__115(w__4 ,in1[21]);
  not g__116(w__3 ,in1[25]);
  not g__117(w__2 ,in1[15]);
  not g__118(w__1 ,in1[9]);
  nor g__119(w__116 ,out1[32] ,w__115);
  and g__120(w__115 ,w__99 ,w__114);
  nor g__121(w__114 ,out1[29] ,w__113);
  or g__122(w__113 ,w__102 ,w__112);
  or g__123(w__112 ,out1[24] ,w__111);
  or g__124(w__111 ,w__104 ,w__110);
  or g__125(w__110 ,out1[19] ,w__109);
  or g__126(w__109 ,w__100 ,w__108);
  or g__127(w__108 ,out1[14] ,w__107);
  or g__128(w__107 ,w__103 ,w__106);
  or g__129(w__106 ,out1[9] ,w__105);
  or g__130(w__105 ,w__93 ,w__101);
  or g__131(w__104 ,w__96 ,w__92);
  or g__132(w__103 ,w__97 ,w__95);
  or g__133(w__102 ,w__94 ,w__89);
  or g__134(w__101 ,w__91 ,w__90);
  or g__135(w__100 ,w__88 ,w__98);
  nor g__136(w__99 ,out1[31] ,out1[30]);
  or g__137(w__98 ,out1[16] ,out1[15]);
  or g__138(w__97 ,out1[13] ,out1[12]);
  or g__139(w__96 ,out1[23] ,out1[22]);
  or g__140(w__95 ,out1[11] ,out1[10]);
  or g__141(w__94 ,out1[28] ,out1[27]);
  or g__142(w__93 ,out1[4] ,out1[3]);
  or g__143(w__92 ,out1[21] ,out1[20]);
  or g__144(w__91 ,out1[8] ,out1[7]);
  or g__145(w__90 ,out1[6] ,out1[5]);
  or g__146(w__89 ,out1[26] ,out1[25]);
  or g__147(w__88 ,out1[18] ,out1[17]);
  buf g__148(out2 ,w__116);
  and g__149(out3 ,out1[32] ,w__175);
  or g__150(w__175 ,w__164 ,w__174);
  or g__151(w__174 ,w__126 ,w__173);
  or g__152(w__173 ,w__160 ,w__172);
  or g__153(w__172 ,w__120 ,w__171);
  or g__154(w__171 ,w__161 ,w__170);
  or g__155(w__170 ,w__143 ,w__169);
  or g__156(w__169 ,w__163 ,w__168);
  or g__157(w__168 ,w__132 ,w__167);
  or g__158(w__167 ,w__162 ,w__166);
  or g__159(w__166 ,w__146 ,w__165);
  or g__160(w__165 ,w__151 ,w__159);
  or g__161(w__164 ,w__136 ,w__152);
  or g__162(w__163 ,w__157 ,w__156);
  or g__163(w__162 ,w__155 ,w__153);
  or g__164(w__161 ,w__154 ,w__150);
  or g__165(w__160 ,w__149 ,w__158);
  or g__166(w__159 ,w__148 ,w__147);
  or g__167(w__158 ,w__131 ,w__129);
  or g__168(w__157 ,w__118 ,w__122);
  or g__169(w__156 ,w__121 ,w__128);
  or g__170(w__155 ,w__119 ,w__124);
  or g__171(w__154 ,w__125 ,w__130);
  or g__172(w__153 ,w__127 ,w__123);
  or g__173(w__152 ,w__141 ,w__145);
  or g__174(w__151 ,w__138 ,w__140);
  or g__175(w__150 ,w__135 ,w__139);
  or g__176(w__149 ,w__137 ,w__144);
  or g__177(w__148 ,w__142 ,w__117);
  or g__178(w__147 ,w__133 ,w__134);
  not g__179(w__146 ,out1[8]);
  not g__180(w__145 ,out1[30]);
  not g__181(w__144 ,out1[26]);
  not g__182(w__143 ,out1[18]);
  not g__183(w__142 ,out1[7]);
  not g__184(w__141 ,out1[31]);
  not g__185(w__140 ,out1[2]);
  not g__186(w__139 ,out1[19]);
  not g__187(w__138 ,out1[3]);
  not g__188(w__137 ,out1[27]);
  not g__189(w__136 ,out1[28]);
  not g__190(w__135 ,out1[20]);
  not g__191(w__134 ,out1[4]);
  not g__192(w__133 ,out1[5]);
  not g__193(w__132 ,out1[13]);
  not g__194(w__131 ,out1[25]);
  not g__195(w__130 ,out1[21]);
  not g__196(w__129 ,out1[24]);
  not g__197(w__128 ,out1[14]);
  not g__198(w__127 ,out1[10]);
  not g__199(w__126 ,out1[29]);
  not g__200(w__125 ,out1[22]);
  not g__201(w__124 ,out1[11]);
  not g__202(w__123 ,out1[9]);
  not g__203(w__122 ,out1[16]);
  not g__204(w__121 ,out1[15]);
  not g__205(w__120 ,out1[23]);
  not g__206(w__119 ,out1[12]);
  not g__207(w__118 ,out1[17]);
  not g__208(w__117 ,out1[6]);
  nor g__209(w__204 ,out4[32] ,w__203);
  and g__210(w__203 ,w__187 ,w__202);
  nor g__211(w__202 ,out4[29] ,w__201);
  or g__212(w__201 ,w__190 ,w__200);
  or g__213(w__200 ,out4[24] ,w__199);
  or g__214(w__199 ,w__192 ,w__198);
  or g__215(w__198 ,out4[19] ,w__197);
  or g__216(w__197 ,w__188 ,w__196);
  or g__217(w__196 ,out4[14] ,w__195);
  or g__218(w__195 ,w__191 ,w__194);
  or g__219(w__194 ,out4[9] ,w__193);
  or g__220(w__193 ,w__181 ,w__189);
  or g__221(w__192 ,w__184 ,w__180);
  or g__222(w__191 ,w__185 ,w__183);
  or g__223(w__190 ,w__182 ,w__177);
  or g__224(w__189 ,w__179 ,w__178);
  or g__225(w__188 ,w__176 ,w__186);
  nor g__226(w__187 ,out4[31] ,out4[30]);
  or g__227(w__186 ,out4[16] ,out4[15]);
  or g__228(w__185 ,out4[13] ,out4[12]);
  or g__229(w__184 ,out4[23] ,out4[22]);
  or g__230(w__183 ,out4[11] ,out4[10]);
  or g__231(w__182 ,out4[28] ,out4[27]);
  or g__232(w__181 ,out4[4] ,out4[3]);
  or g__233(w__180 ,out4[21] ,out4[20]);
  or g__234(w__179 ,out4[8] ,out4[7]);
  or g__235(w__178 ,out4[6] ,out4[5]);
  or g__236(w__177 ,out4[26] ,out4[25]);
  or g__237(w__176 ,out4[18] ,out4[17]);
  buf g__238(out5 ,w__204);
  and g__239(out6 ,out4[32] ,w__263);
  or g__240(w__263 ,w__252 ,w__262);
  or g__241(w__262 ,w__214 ,w__261);
  or g__242(w__261 ,w__248 ,w__260);
  or g__243(w__260 ,w__208 ,w__259);
  or g__244(w__259 ,w__249 ,w__258);
  or g__245(w__258 ,w__231 ,w__257);
  or g__246(w__257 ,w__251 ,w__256);
  or g__247(w__256 ,w__220 ,w__255);
  or g__248(w__255 ,w__250 ,w__254);
  or g__249(w__254 ,w__234 ,w__253);
  or g__250(w__253 ,w__239 ,w__247);
  or g__251(w__252 ,w__224 ,w__240);
  or g__252(w__251 ,w__245 ,w__244);
  or g__253(w__250 ,w__243 ,w__241);
  or g__254(w__249 ,w__242 ,w__238);
  or g__255(w__248 ,w__237 ,w__246);
  or g__256(w__247 ,w__236 ,w__235);
  or g__257(w__246 ,w__219 ,w__217);
  or g__258(w__245 ,w__206 ,w__210);
  or g__259(w__244 ,w__209 ,w__216);
  or g__260(w__243 ,w__207 ,w__212);
  or g__261(w__242 ,w__213 ,w__218);
  or g__262(w__241 ,w__215 ,w__211);
  or g__263(w__240 ,w__229 ,w__233);
  or g__264(w__239 ,w__226 ,w__228);
  or g__265(w__238 ,w__223 ,w__227);
  or g__266(w__237 ,w__225 ,w__232);
  or g__267(w__236 ,w__230 ,w__205);
  or g__268(w__235 ,w__221 ,w__222);
  not g__269(w__234 ,out4[8]);
  not g__270(w__233 ,out4[30]);
  not g__271(w__232 ,out4[26]);
  not g__272(w__231 ,out4[18]);
  not g__273(w__230 ,out4[7]);
  not g__274(w__229 ,out4[31]);
  not g__275(w__228 ,out4[2]);
  not g__276(w__227 ,out4[19]);
  not g__277(w__226 ,out4[3]);
  not g__278(w__225 ,out4[27]);
  not g__279(w__224 ,out4[28]);
  not g__280(w__223 ,out4[20]);
  not g__281(w__222 ,out4[4]);
  not g__282(w__221 ,out4[5]);
  not g__283(w__220 ,out4[13]);
  not g__284(w__219 ,out4[25]);
  not g__285(w__218 ,out4[21]);
  not g__286(w__217 ,out4[24]);
  not g__287(w__216 ,out4[14]);
  not g__288(w__215 ,out4[10]);
  not g__289(w__214 ,out4[29]);
  not g__290(w__213 ,out4[22]);
  not g__291(w__212 ,out4[11]);
  not g__292(w__211 ,out4[9]);
  not g__293(w__210 ,out4[16]);
  not g__294(w__209 ,out4[15]);
  not g__295(w__208 ,out4[23]);
  not g__296(w__207 ,out4[12]);
  not g__297(w__206 ,out4[17]);
  not g__298(w__205 ,out4[6]);
  or g__299(w__581 ,w__425 ,w__579);
  xnor g__300(w__580 ,w__578 ,w__470);
  and g__301(w__579 ,w__404 ,w__578);
  and g__302(w__578 ,w__449 ,w__576);
  xnor g__303(w__577 ,w__575 ,w__469);
  or g__304(w__576 ,w__415 ,w__575);
  and g__305(w__575 ,w__403 ,w__573);
  xnor g__306(w__574 ,w__572 ,w__468);
  or g__307(w__573 ,w__441 ,w__572);
  and g__308(w__572 ,w__437 ,w__570);
  xnor g__309(w__571 ,w__569 ,w__467);
  or g__310(w__570 ,w__420 ,w__569);
  and g__311(w__569 ,w__414 ,w__567);
  xnor g__312(w__568 ,w__566 ,w__466);
  or g__313(w__567 ,w__398 ,w__566);
  and g__314(w__566 ,w__457 ,w__564);
  xnor g__315(w__565 ,w__563 ,w__465);
  or g__316(w__564 ,w__444 ,w__563);
  and g__317(w__563 ,w__433 ,w__561);
  xnor g__318(w__562 ,w__560 ,w__464);
  or g__319(w__561 ,w__434 ,w__560);
  and g__320(w__560 ,w__432 ,w__558);
  xnor g__321(w__559 ,w__557 ,w__463);
  or g__322(w__558 ,w__421 ,w__557);
  and g__323(w__557 ,w__419 ,w__555);
  xnor g__324(w__556 ,w__554 ,w__462);
  or g__325(w__555 ,w__459 ,w__554);
  and g__326(w__554 ,w__409 ,w__552);
  xnor g__327(w__553 ,w__551 ,w__461);
  or g__328(w__552 ,w__400 ,w__551);
  and g__329(w__551 ,w__397 ,w__549);
  xnor g__330(w__550 ,w__548 ,w__460);
  or g__331(w__549 ,w__438 ,w__548);
  and g__332(w__548 ,w__453 ,w__546);
  xnor g__333(w__547 ,w__545 ,w__490);
  or g__334(w__546 ,w__443 ,w__545);
  and g__335(w__545 ,w__448 ,w__543);
  xnor g__336(w__544 ,w__542 ,w__489);
  or g__337(w__543 ,w__442 ,w__542);
  and g__338(w__542 ,w__439 ,w__540);
  xnor g__339(w__541 ,w__539 ,w__488);
  or g__340(w__540 ,w__413 ,w__539);
  and g__341(w__539 ,w__430 ,w__537);
  xnor g__342(w__538 ,w__536 ,w__487);
  or g__343(w__537 ,w__456 ,w__536);
  and g__344(w__536 ,w__429 ,w__534);
  xnor g__345(w__535 ,w__533 ,w__486);
  or g__346(w__534 ,w__423 ,w__533);
  and g__347(w__533 ,w__422 ,w__531);
  xnor g__348(w__532 ,w__530 ,w__485);
  or g__349(w__531 ,w__418 ,w__530);
  and g__350(w__530 ,w__417 ,w__528);
  xnor g__351(w__529 ,w__527 ,w__484);
  or g__352(w__528 ,w__412 ,w__527);
  and g__353(w__527 ,w__427 ,w__525);
  xnor g__354(w__526 ,w__524 ,w__483);
  or g__355(w__525 ,w__406 ,w__524);
  and g__356(w__524 ,w__405 ,w__522);
  xnor g__357(w__523 ,w__521 ,w__482);
  or g__358(w__522 ,w__402 ,w__521);
  and g__359(w__521 ,w__401 ,w__519);
  xnor g__360(w__520 ,w__518 ,w__481);
  or g__361(w__519 ,w__426 ,w__518);
  and g__362(w__518 ,w__458 ,w__516);
  xnor g__363(w__517 ,w__515 ,w__480);
  or g__364(w__516 ,w__455 ,w__515);
  and g__365(w__515 ,w__454 ,w__513);
  xnor g__366(w__514 ,w__512 ,w__479);
  or g__367(w__513 ,w__452 ,w__512);
  and g__368(w__512 ,w__451 ,w__510);
  xnor g__369(w__511 ,w__509 ,w__478);
  or g__370(w__510 ,w__447 ,w__509);
  and g__371(w__509 ,w__446 ,w__507);
  xnor g__372(w__508 ,w__506 ,w__477);
  or g__373(w__507 ,w__450 ,w__506);
  and g__374(w__506 ,w__431 ,w__504);
  xnor g__375(w__505 ,w__503 ,w__476);
  or g__376(w__504 ,w__440 ,w__503);
  and g__377(w__503 ,w__445 ,w__501);
  xnor g__378(w__502 ,w__500 ,w__475);
  or g__379(w__501 ,w__407 ,w__500);
  and g__380(w__500 ,w__399 ,w__498);
  xnor g__381(w__499 ,w__497 ,w__474);
  or g__382(w__498 ,w__410 ,w__497);
  and g__383(w__497 ,w__435 ,w__495);
  xnor g__384(w__496 ,w__494 ,w__473);
  or g__385(w__495 ,w__408 ,w__494);
  and g__386(w__494 ,w__424 ,w__493);
  xnor g__387(out1[2] ,w__492 ,w__472);
  or g__388(w__493 ,w__416 ,w__492);
  xnor g__389(out1[1] ,w__428 ,w__471);
  and g__390(w__492 ,w__436 ,w__491);
  xor g__391(out1[0] ,in2[0] ,in1[0]);
  or g__392(w__491 ,w__411 ,w__428);
  xnor g__393(w__490 ,w__338 ,in2[20]);
  xnor g__394(w__489 ,w__329 ,in2[19]);
  xnor g__395(w__488 ,w__315 ,in2[18]);
  xnor g__396(w__487 ,w__331 ,in2[17]);
  xnor g__397(w__486 ,w__318 ,in2[16]);
  xnor g__398(w__485 ,w__320 ,in2[15]);
  xnor g__399(w__484 ,w__333 ,in2[14]);
  xnor g__400(w__483 ,w__324 ,in2[13]);
  xnor g__401(w__482 ,w__335 ,in2[12]);
  xnor g__402(w__481 ,w__327 ,in2[11]);
  xnor g__403(w__480 ,w__339 ,in2[10]);
  xnor g__404(w__479 ,w__330 ,in2[9]);
  xnor g__405(w__478 ,w__340 ,in2[8]);
  xnor g__406(w__477 ,w__322 ,in2[7]);
  xnor g__407(w__476 ,w__336 ,in2[6]);
  xnor g__408(w__475 ,w__303 ,in2[5]);
  xnor g__409(w__474 ,w__341 ,in2[4]);
  xnor g__410(w__473 ,w__300 ,in2[3]);
  xnor g__411(w__472 ,w__332 ,in2[2]);
  xnor g__412(w__471 ,w__297 ,in2[1]);
  xnor g__413(w__470 ,w__319 ,in2[31]);
  xnor g__414(w__469 ,w__306 ,in2[30]);
  xnor g__415(w__468 ,w__321 ,in2[29]);
  xnor g__416(w__467 ,w__309 ,in2[28]);
  xnor g__417(w__466 ,w__323 ,in2[27]);
  xnor g__418(w__465 ,w__334 ,in2[26]);
  xnor g__419(w__464 ,w__325 ,in2[25]);
  xnor g__420(w__463 ,w__312 ,in2[24]);
  xnor g__421(w__462 ,w__326 ,in2[23]);
  xnor g__422(w__461 ,w__337 ,in2[22]);
  xnor g__423(w__460 ,w__328 ,in2[21]);
  nor g__424(w__459 ,w__345 ,in2[23]);
  or g__425(w__458 ,w__375 ,w__339);
  or g__426(w__457 ,w__368 ,w__334);
  nor g__427(w__456 ,w__355 ,in2[17]);
  nor g__428(w__455 ,w__350 ,in2[10]);
  or g__429(w__454 ,w__395 ,w__330);
  or g__430(w__453 ,w__388 ,w__338);
  nor g__431(w__452 ,w__342 ,in2[9]);
  or g__432(w__451 ,w__390 ,w__340);
  nor g__433(w__450 ,w__348 ,in2[7]);
  or g__434(w__449 ,w__369 ,w__305);
  or g__435(w__448 ,w__383 ,w__329);
  nor g__436(w__447 ,w__354 ,in2[8]);
  or g__437(w__446 ,w__373 ,w__322);
  or g__438(w__445 ,w__394 ,w__302);
  nor g__439(w__444 ,w__364 ,in2[26]);
  nor g__440(w__443 ,w__357 ,in2[20]);
  nor g__441(w__442 ,w__347 ,in2[19]);
  nor g__442(w__441 ,w__359 ,in2[29]);
  nor g__443(w__440 ,w__358 ,in2[6]);
  or g__444(w__439 ,w__387 ,w__314);
  nor g__445(w__438 ,w__349 ,in2[21]);
  or g__446(w__437 ,w__376 ,w__308);
  or g__447(w__436 ,w__386 ,w__296);
  or g__448(w__435 ,w__380 ,w__299);
  nor g__449(w__434 ,w__351 ,in2[25]);
  or g__450(w__433 ,w__367 ,w__325);
  or g__451(w__432 ,w__382 ,w__311);
  or g__452(w__431 ,w__372 ,w__336);
  or g__453(w__430 ,w__370 ,w__331);
  or g__454(w__429 ,w__366 ,w__317);
  or g__455(w__427 ,w__393 ,w__324);
  nor g__456(w__426 ,w__360 ,in2[11]);
  nor g__457(w__425 ,w__343 ,in2[31]);
  or g__458(w__424 ,w__374 ,w__332);
  and g__459(w__423 ,w__318 ,w__366);
  or g__460(w__422 ,w__379 ,w__320);
  and g__461(w__421 ,w__312 ,w__382);
  and g__462(w__420 ,w__309 ,w__376);
  or g__463(w__419 ,w__371 ,w__326);
  nor g__464(w__418 ,w__344 ,in2[15]);
  or g__465(w__417 ,w__389 ,w__333);
  nor g__466(w__416 ,w__353 ,in2[2]);
  and g__467(w__415 ,w__306 ,w__369);
  or g__468(w__414 ,w__391 ,w__323);
  and g__469(w__413 ,w__315 ,w__387);
  nor g__470(w__412 ,w__352 ,in2[14]);
  and g__471(w__411 ,w__297 ,w__386);
  nor g__472(w__410 ,w__361 ,in2[4]);
  or g__473(w__409 ,w__365 ,w__337);
  and g__474(w__408 ,w__300 ,w__380);
  and g__475(w__407 ,w__303 ,w__394);
  nor g__476(w__406 ,w__363 ,in2[13]);
  or g__477(w__405 ,w__396 ,w__335);
  or g__478(w__404 ,w__384 ,w__319);
  or g__479(w__403 ,w__381 ,w__321);
  nor g__480(w__402 ,w__356 ,in2[12]);
  or g__481(w__401 ,w__385 ,w__327);
  nor g__482(w__400 ,w__362 ,in2[22]);
  or g__483(w__399 ,w__378 ,w__341);
  nor g__484(w__398 ,w__346 ,in2[27]);
  or g__485(w__397 ,w__392 ,w__328);
  and g__486(w__428 ,in1[0] ,w__377);
  not g__487(w__396 ,in2[12]);
  not g__488(w__395 ,in2[9]);
  not g__489(w__394 ,in2[5]);
  not g__490(w__393 ,in2[13]);
  not g__491(w__392 ,in2[21]);
  not g__492(w__391 ,in2[27]);
  not g__493(w__390 ,in2[8]);
  not g__494(w__389 ,in2[14]);
  not g__495(w__388 ,in2[20]);
  not g__496(w__387 ,in2[18]);
  not g__497(w__386 ,in2[1]);
  not g__498(w__385 ,in2[11]);
  not g__499(w__384 ,in2[31]);
  not g__500(w__383 ,in2[19]);
  not g__501(w__382 ,in2[24]);
  not g__502(w__381 ,in2[29]);
  not g__503(w__380 ,in2[3]);
  not g__504(w__379 ,in2[15]);
  not g__505(w__378 ,in2[4]);
  not g__506(w__377 ,in2[0]);
  not g__507(w__376 ,in2[28]);
  not g__508(w__375 ,in2[10]);
  not g__509(w__374 ,in2[2]);
  not g__510(w__373 ,in2[7]);
  not g__511(w__372 ,in2[6]);
  not g__512(w__371 ,in2[23]);
  not g__513(w__370 ,in2[17]);
  not g__514(w__369 ,in2[30]);
  not g__515(w__368 ,in2[26]);
  not g__516(w__367 ,in2[25]);
  not g__517(w__366 ,in2[16]);
  not g__518(w__365 ,in2[22]);
  not g__519(w__341 ,w__361);
  not g__520(w__361 ,w__267);
  not g__521(w__340 ,w__354);
  not g__522(w__354 ,w__271);
  not g__523(w__339 ,w__350);
  not g__524(w__350 ,w__273);
  not g__525(w__338 ,w__357);
  not g__526(w__357 ,w__283);
  not g__527(w__337 ,w__362);
  not g__528(w__362 ,w__285);
  not g__529(w__336 ,w__358);
  not g__530(w__358 ,w__269);
  not g__531(w__335 ,w__356);
  not g__532(w__356 ,w__275);
  not g__533(w__334 ,w__364);
  not g__534(w__364 ,w__289);
  not g__535(w__333 ,w__352);
  not g__536(w__352 ,w__277);
  not g__537(w__332 ,w__353);
  not g__538(w__353 ,w__265);
  not g__539(w__331 ,w__355);
  not g__540(w__355 ,w__280);
  not g__541(w__330 ,w__342);
  not g__542(w__342 ,w__272);
  not g__543(w__329 ,w__347);
  not g__544(w__347 ,w__282);
  not g__545(w__328 ,w__349);
  not g__546(w__349 ,w__284);
  not g__547(w__327 ,w__360);
  not g__548(w__360 ,w__274);
  not g__549(w__326 ,w__345);
  not g__550(w__345 ,w__286);
  not g__551(w__325 ,w__351);
  not g__552(w__351 ,w__288);
  not g__553(w__324 ,w__363);
  not g__554(w__363 ,w__276);
  not g__555(w__323 ,w__346);
  not g__556(w__346 ,w__290);
  not g__557(w__322 ,w__348);
  not g__558(w__348 ,w__270);
  not g__559(w__321 ,w__359);
  not g__560(w__359 ,w__292);
  not g__561(w__320 ,w__344);
  not g__562(w__344 ,w__278);
  not g__563(w__319 ,w__343);
  not g__564(w__343 ,w__294);
  not g__565(w__318 ,w__316);
  not g__566(w__317 ,w__316);
  not g__567(w__316 ,w__279);
  not g__568(w__315 ,w__313);
  not g__569(w__314 ,w__313);
  not g__570(w__313 ,w__281);
  not g__571(w__312 ,w__310);
  not g__572(w__311 ,w__310);
  not g__573(w__310 ,w__287);
  not g__574(w__309 ,w__307);
  not g__575(w__308 ,w__307);
  not g__576(w__307 ,w__291);
  not g__577(w__306 ,w__304);
  not g__578(w__305 ,w__304);
  not g__579(w__304 ,w__293);
  not g__580(w__303 ,w__301);
  not g__581(w__302 ,w__301);
  not g__582(w__301 ,w__268);
  not g__583(w__300 ,w__298);
  not g__584(w__299 ,w__298);
  not g__585(w__298 ,w__266);
  not g__586(w__297 ,w__295);
  not g__587(w__296 ,w__295);
  not g__588(w__295 ,w__264);
  buf g__589(out1[31] ,w__580);
  buf g__590(out1[29] ,w__574);
  buf g__591(out1[30] ,w__577);
  buf g__592(out1[32] ,w__581);
  buf g__593(out1[10] ,w__517);
  buf g__594(out1[7] ,w__508);
  buf g__595(out1[8] ,w__511);
  buf g__596(out1[19] ,w__544);
  buf g__597(out1[14] ,w__529);
  buf g__598(out1[4] ,w__499);
  buf g__599(out1[3] ,w__496);
  buf g__600(out1[5] ,w__502);
  buf g__601(out1[11] ,w__520);
  buf g__602(out1[12] ,w__523);
  buf g__603(out1[25] ,w__562);
  buf g__604(out1[21] ,w__550);
  buf g__605(out1[27] ,w__568);
  buf g__606(out1[23] ,w__556);
  buf g__607(out1[18] ,w__541);
  buf g__608(out1[24] ,w__559);
  buf g__609(out1[15] ,w__532);
  buf g__610(out1[16] ,w__535);
  buf g__611(out1[17] ,w__538);
  buf g__612(out1[22] ,w__553);
  buf g__613(out1[28] ,w__571);
  buf g__614(out1[6] ,w__505);
  buf g__615(out1[26] ,w__565);
  buf g__616(out1[9] ,w__514);
  buf g__617(out1[13] ,w__526);
  buf g__618(out1[20] ,w__547);
  or g__619(w__868 ,w__712 ,w__866);
  xnor g__620(w__867 ,w__865 ,w__757);
  and g__621(w__866 ,w__691 ,w__865);
  and g__622(w__865 ,w__736 ,w__863);
  xnor g__623(w__864 ,w__862 ,w__756);
  or g__624(w__863 ,w__702 ,w__862);
  and g__625(w__862 ,w__690 ,w__860);
  xnor g__626(w__861 ,w__859 ,w__755);
  or g__627(w__860 ,w__728 ,w__859);
  and g__628(w__859 ,w__724 ,w__857);
  xnor g__629(w__858 ,w__856 ,w__754);
  or g__630(w__857 ,w__707 ,w__856);
  and g__631(w__856 ,w__701 ,w__854);
  xnor g__632(w__855 ,w__853 ,w__753);
  or g__633(w__854 ,w__685 ,w__853);
  and g__634(w__853 ,w__744 ,w__851);
  xnor g__635(w__852 ,w__850 ,w__752);
  or g__636(w__851 ,w__731 ,w__850);
  and g__637(w__850 ,w__720 ,w__848);
  xnor g__638(w__849 ,w__847 ,w__751);
  or g__639(w__848 ,w__721 ,w__847);
  and g__640(w__847 ,w__719 ,w__845);
  xnor g__641(w__846 ,w__844 ,w__750);
  or g__642(w__845 ,w__708 ,w__844);
  and g__643(w__844 ,w__706 ,w__842);
  xnor g__644(w__843 ,w__841 ,w__749);
  or g__645(w__842 ,w__746 ,w__841);
  and g__646(w__841 ,w__696 ,w__839);
  xnor g__647(w__840 ,w__838 ,w__748);
  or g__648(w__839 ,w__687 ,w__838);
  and g__649(w__838 ,w__684 ,w__836);
  xnor g__650(w__837 ,w__835 ,w__747);
  or g__651(w__836 ,w__725 ,w__835);
  and g__652(w__835 ,w__740 ,w__833);
  xnor g__653(w__834 ,w__832 ,w__777);
  or g__654(w__833 ,w__730 ,w__832);
  and g__655(w__832 ,w__735 ,w__830);
  xnor g__656(w__831 ,w__829 ,w__776);
  or g__657(w__830 ,w__729 ,w__829);
  and g__658(w__829 ,w__726 ,w__827);
  xnor g__659(w__828 ,w__826 ,w__775);
  or g__660(w__827 ,w__700 ,w__826);
  and g__661(w__826 ,w__717 ,w__824);
  xnor g__662(w__825 ,w__823 ,w__774);
  or g__663(w__824 ,w__743 ,w__823);
  and g__664(w__823 ,w__716 ,w__821);
  xnor g__665(w__822 ,w__820 ,w__773);
  or g__666(w__821 ,w__710 ,w__820);
  and g__667(w__820 ,w__709 ,w__818);
  xnor g__668(w__819 ,w__817 ,w__772);
  or g__669(w__818 ,w__705 ,w__817);
  and g__670(w__817 ,w__704 ,w__815);
  xnor g__671(w__816 ,w__814 ,w__771);
  or g__672(w__815 ,w__699 ,w__814);
  and g__673(w__814 ,w__714 ,w__812);
  xnor g__674(w__813 ,w__811 ,w__770);
  or g__675(w__812 ,w__693 ,w__811);
  and g__676(w__811 ,w__692 ,w__809);
  xnor g__677(w__810 ,w__808 ,w__769);
  or g__678(w__809 ,w__689 ,w__808);
  and g__679(w__808 ,w__688 ,w__806);
  xnor g__680(w__807 ,w__805 ,w__768);
  or g__681(w__806 ,w__713 ,w__805);
  and g__682(w__805 ,w__745 ,w__803);
  xnor g__683(w__804 ,w__802 ,w__767);
  or g__684(w__803 ,w__742 ,w__802);
  and g__685(w__802 ,w__741 ,w__800);
  xnor g__686(w__801 ,w__799 ,w__766);
  or g__687(w__800 ,w__739 ,w__799);
  and g__688(w__799 ,w__738 ,w__797);
  xnor g__689(w__798 ,w__796 ,w__765);
  or g__690(w__797 ,w__734 ,w__796);
  and g__691(w__796 ,w__733 ,w__794);
  xnor g__692(w__795 ,w__793 ,w__764);
  or g__693(w__794 ,w__737 ,w__793);
  and g__694(w__793 ,w__718 ,w__791);
  xnor g__695(w__792 ,w__790 ,w__763);
  or g__696(w__791 ,w__727 ,w__790);
  and g__697(w__790 ,w__732 ,w__788);
  xnor g__698(w__789 ,w__787 ,w__762);
  or g__699(w__788 ,w__694 ,w__787);
  and g__700(w__787 ,w__686 ,w__785);
  xnor g__701(w__786 ,w__784 ,w__761);
  or g__702(w__785 ,w__697 ,w__784);
  and g__703(w__784 ,w__722 ,w__782);
  xnor g__704(w__783 ,w__781 ,w__760);
  or g__705(w__782 ,w__695 ,w__781);
  and g__706(w__781 ,w__711 ,w__780);
  xnor g__707(out4[2] ,w__779 ,w__759);
  or g__708(w__780 ,w__703 ,w__779);
  xnor g__709(out4[1] ,w__715 ,w__758);
  and g__710(w__779 ,w__723 ,w__778);
  xor g__711(out4[0] ,in3[0] ,in1[0]);
  or g__712(w__778 ,w__698 ,w__715);
  xnor g__713(w__777 ,w__625 ,in3[20]);
  xnor g__714(w__776 ,w__616 ,in3[19]);
  xnor g__715(w__775 ,w__602 ,in3[18]);
  xnor g__716(w__774 ,w__618 ,in3[17]);
  xnor g__717(w__773 ,w__605 ,in3[16]);
  xnor g__718(w__772 ,w__607 ,in3[15]);
  xnor g__719(w__771 ,w__620 ,in3[14]);
  xnor g__720(w__770 ,w__611 ,in3[13]);
  xnor g__721(w__769 ,w__622 ,in3[12]);
  xnor g__722(w__768 ,w__614 ,in3[11]);
  xnor g__723(w__767 ,w__626 ,in3[10]);
  xnor g__724(w__766 ,w__617 ,in3[9]);
  xnor g__725(w__765 ,w__627 ,in3[8]);
  xnor g__726(w__764 ,w__609 ,in3[7]);
  xnor g__727(w__763 ,w__623 ,in3[6]);
  xnor g__728(w__762 ,w__590 ,in3[5]);
  xnor g__729(w__761 ,w__628 ,in3[4]);
  xnor g__730(w__760 ,w__587 ,in3[3]);
  xnor g__731(w__759 ,w__619 ,in3[2]);
  xnor g__732(w__758 ,w__584 ,in3[1]);
  xnor g__733(w__757 ,w__606 ,in3[31]);
  xnor g__734(w__756 ,w__593 ,in3[30]);
  xnor g__735(w__755 ,w__608 ,in3[29]);
  xnor g__736(w__754 ,w__596 ,in3[28]);
  xnor g__737(w__753 ,w__610 ,in3[27]);
  xnor g__738(w__752 ,w__621 ,in3[26]);
  xnor g__739(w__751 ,w__612 ,in3[25]);
  xnor g__740(w__750 ,w__599 ,in3[24]);
  xnor g__741(w__749 ,w__613 ,in3[23]);
  xnor g__742(w__748 ,w__624 ,in3[22]);
  xnor g__743(w__747 ,w__615 ,in3[21]);
  nor g__744(w__746 ,w__632 ,in3[23]);
  or g__745(w__745 ,w__662 ,w__626);
  or g__746(w__744 ,w__655 ,w__621);
  nor g__747(w__743 ,w__642 ,in3[17]);
  nor g__748(w__742 ,w__637 ,in3[10]);
  or g__749(w__741 ,w__682 ,w__617);
  or g__750(w__740 ,w__675 ,w__625);
  nor g__751(w__739 ,w__629 ,in3[9]);
  or g__752(w__738 ,w__677 ,w__627);
  nor g__753(w__737 ,w__635 ,in3[7]);
  or g__754(w__736 ,w__656 ,w__592);
  or g__755(w__735 ,w__670 ,w__616);
  nor g__756(w__734 ,w__641 ,in3[8]);
  or g__757(w__733 ,w__660 ,w__609);
  or g__758(w__732 ,w__681 ,w__589);
  nor g__759(w__731 ,w__651 ,in3[26]);
  nor g__760(w__730 ,w__644 ,in3[20]);
  nor g__761(w__729 ,w__634 ,in3[19]);
  nor g__762(w__728 ,w__646 ,in3[29]);
  nor g__763(w__727 ,w__645 ,in3[6]);
  or g__764(w__726 ,w__674 ,w__601);
  nor g__765(w__725 ,w__636 ,in3[21]);
  or g__766(w__724 ,w__663 ,w__595);
  or g__767(w__723 ,w__673 ,w__583);
  or g__768(w__722 ,w__667 ,w__586);
  nor g__769(w__721 ,w__638 ,in3[25]);
  or g__770(w__720 ,w__654 ,w__612);
  or g__771(w__719 ,w__669 ,w__598);
  or g__772(w__718 ,w__659 ,w__623);
  or g__773(w__717 ,w__657 ,w__618);
  or g__774(w__716 ,w__653 ,w__604);
  or g__775(w__714 ,w__680 ,w__611);
  nor g__776(w__713 ,w__647 ,in3[11]);
  nor g__777(w__712 ,w__630 ,in3[31]);
  or g__778(w__711 ,w__661 ,w__619);
  and g__779(w__710 ,w__605 ,w__653);
  or g__780(w__709 ,w__666 ,w__607);
  and g__781(w__708 ,w__599 ,w__669);
  and g__782(w__707 ,w__596 ,w__663);
  or g__783(w__706 ,w__658 ,w__613);
  nor g__784(w__705 ,w__631 ,in3[15]);
  or g__785(w__704 ,w__676 ,w__620);
  nor g__786(w__703 ,w__640 ,in3[2]);
  and g__787(w__702 ,w__593 ,w__656);
  or g__788(w__701 ,w__678 ,w__610);
  and g__789(w__700 ,w__602 ,w__674);
  nor g__790(w__699 ,w__639 ,in3[14]);
  and g__791(w__698 ,w__584 ,w__673);
  nor g__792(w__697 ,w__648 ,in3[4]);
  or g__793(w__696 ,w__652 ,w__624);
  and g__794(w__695 ,w__587 ,w__667);
  and g__795(w__694 ,w__590 ,w__681);
  nor g__796(w__693 ,w__650 ,in3[13]);
  or g__797(w__692 ,w__683 ,w__622);
  or g__798(w__691 ,w__671 ,w__606);
  or g__799(w__690 ,w__668 ,w__608);
  nor g__800(w__689 ,w__643 ,in3[12]);
  or g__801(w__688 ,w__672 ,w__614);
  nor g__802(w__687 ,w__649 ,in3[22]);
  or g__803(w__686 ,w__665 ,w__628);
  nor g__804(w__685 ,w__633 ,in3[27]);
  or g__805(w__684 ,w__679 ,w__615);
  and g__806(w__715 ,in1[0] ,w__664);
  not g__807(w__683 ,in3[12]);
  not g__808(w__682 ,in3[9]);
  not g__809(w__681 ,in3[5]);
  not g__810(w__680 ,in3[13]);
  not g__811(w__679 ,in3[21]);
  not g__812(w__678 ,in3[27]);
  not g__813(w__677 ,in3[8]);
  not g__814(w__676 ,in3[14]);
  not g__815(w__675 ,in3[20]);
  not g__816(w__674 ,in3[18]);
  not g__817(w__673 ,in3[1]);
  not g__818(w__672 ,in3[11]);
  not g__819(w__671 ,in3[31]);
  not g__820(w__670 ,in3[19]);
  not g__821(w__669 ,in3[24]);
  not g__822(w__668 ,in3[29]);
  not g__823(w__667 ,in3[3]);
  not g__824(w__666 ,in3[15]);
  not g__825(w__665 ,in3[4]);
  not g__826(w__664 ,in3[0]);
  not g__827(w__663 ,in3[28]);
  not g__828(w__662 ,in3[10]);
  not g__829(w__661 ,in3[2]);
  not g__830(w__660 ,in3[7]);
  not g__831(w__659 ,in3[6]);
  not g__832(w__658 ,in3[23]);
  not g__833(w__657 ,in3[17]);
  not g__834(w__656 ,in3[30]);
  not g__835(w__655 ,in3[26]);
  not g__836(w__654 ,in3[25]);
  not g__837(w__653 ,in3[16]);
  not g__838(w__652 ,in3[22]);
  not g__839(w__628 ,w__648);
  not g__840(w__648 ,w__267);
  not g__841(w__627 ,w__641);
  not g__842(w__641 ,w__271);
  not g__843(w__626 ,w__637);
  not g__844(w__637 ,w__273);
  not g__845(w__625 ,w__644);
  not g__846(w__644 ,w__283);
  not g__847(w__624 ,w__649);
  not g__848(w__649 ,w__285);
  not g__849(w__623 ,w__645);
  not g__850(w__645 ,w__269);
  not g__851(w__622 ,w__643);
  not g__852(w__643 ,w__275);
  not g__853(w__621 ,w__651);
  not g__854(w__651 ,w__289);
  not g__855(w__620 ,w__639);
  not g__856(w__639 ,w__277);
  not g__857(w__619 ,w__640);
  not g__858(w__640 ,w__265);
  not g__859(w__618 ,w__642);
  not g__860(w__642 ,w__280);
  not g__861(w__617 ,w__629);
  not g__862(w__629 ,w__272);
  not g__863(w__616 ,w__634);
  not g__864(w__634 ,w__282);
  not g__865(w__615 ,w__636);
  not g__866(w__636 ,w__284);
  not g__867(w__614 ,w__647);
  not g__868(w__647 ,w__274);
  not g__869(w__613 ,w__632);
  not g__870(w__632 ,w__286);
  not g__871(w__612 ,w__638);
  not g__872(w__638 ,w__288);
  not g__873(w__611 ,w__650);
  not g__874(w__650 ,w__276);
  not g__875(w__610 ,w__633);
  not g__876(w__633 ,w__290);
  not g__877(w__609 ,w__635);
  not g__878(w__635 ,w__270);
  not g__879(w__608 ,w__646);
  not g__880(w__646 ,w__292);
  not g__881(w__607 ,w__631);
  not g__882(w__631 ,w__278);
  not g__883(w__606 ,w__630);
  not g__884(w__630 ,w__294);
  not g__885(w__605 ,w__603);
  not g__886(w__604 ,w__603);
  not g__887(w__603 ,w__279);
  not g__888(w__602 ,w__600);
  not g__889(w__601 ,w__600);
  not g__890(w__600 ,w__281);
  not g__891(w__599 ,w__597);
  not g__892(w__598 ,w__597);
  not g__893(w__597 ,w__287);
  not g__894(w__596 ,w__594);
  not g__895(w__595 ,w__594);
  not g__896(w__594 ,w__291);
  not g__897(w__593 ,w__591);
  not g__898(w__592 ,w__591);
  not g__899(w__591 ,w__293);
  not g__900(w__590 ,w__588);
  not g__901(w__589 ,w__588);
  not g__902(w__588 ,w__268);
  not g__903(w__587 ,w__585);
  not g__904(w__586 ,w__585);
  not g__905(w__585 ,w__266);
  not g__906(w__584 ,w__582);
  not g__907(w__583 ,w__582);
  not g__908(w__582 ,w__264);
  buf g__909(out4[31] ,w__867);
  buf g__910(out4[29] ,w__861);
  buf g__911(out4[30] ,w__864);
  buf g__912(out4[32] ,w__868);
  buf g__913(out4[10] ,w__804);
  buf g__914(out4[7] ,w__795);
  buf g__915(out4[8] ,w__798);
  buf g__916(out4[19] ,w__831);
  buf g__917(out4[14] ,w__816);
  buf g__918(out4[4] ,w__786);
  buf g__919(out4[3] ,w__783);
  buf g__920(out4[5] ,w__789);
  buf g__921(out4[11] ,w__807);
  buf g__922(out4[12] ,w__810);
  buf g__923(out4[25] ,w__849);
  buf g__924(out4[21] ,w__837);
  buf g__925(out4[27] ,w__855);
  buf g__926(out4[23] ,w__843);
  buf g__927(out4[18] ,w__828);
  buf g__928(out4[24] ,w__846);
  buf g__929(out4[15] ,w__819);
  buf g__930(out4[16] ,w__822);
  buf g__931(out4[17] ,w__825);
  buf g__932(out4[22] ,w__840);
  buf g__933(out4[28] ,w__858);
  buf g__934(out4[6] ,w__792);
  buf g__935(out4[26] ,w__852);
  buf g__936(out4[9] ,w__801);
  buf g__937(out4[13] ,w__813);
  buf g__938(out4[20] ,w__834);
endmodule
