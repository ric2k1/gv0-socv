module top( 2_n5 , 2_n13 , 2_n17 , 2_n20 , 2_n27 , 2_n36 , 2_n37 , 2_n53 , 2_n62 , 2_n75 , 2_n80 , 2_n86 , 2_n93 , 2_n105 , 2_n106 , 2_n111 , 2_n117 , 2_n139 , 2_n145 , 2_n147 , 2_n157 , 2_n161 , 2_n175 , 2_n176 , 2_n182 , 2_n190 , 2_n198 , 2_n204 , 2_n208 , 2_n214 , 2_n217 , 2_n219 , 2_n224 , 2_n225 , 2_n226 , 2_n229 , 2_n235 , 2_n241 , 2_n244 , 2_n249 , 2_n256 , 2_n281 , 2_n287 , 2_n289 , 2_n294 , 2_n300 , 2_n303 , 2_n319 , 2_n345 , 2_n346 , 2_n364 , 2_n365 , 2_n368 , 2_n384 , 2_n387 , 2_n389 , 2_n393 , 2_n403 , 2_n409 , 2_n410 , 2_n417 , 2_n430 , 2_n439 , 2_n442 , 2_n457 , 2_n465 , 2_n473 , 2_n477 , 2_n489 , 2_n491 , 2_n493 , 2_n503 , 2_n506 , 2_n511 , 2_n515 , 2_n518 , 2_n521 , 2_n532 , 2_n537 , 2_n587 , 2_n588 , 2_n593 , 2_n594 , 2_n595 , 2_n606 , 2_n618 , 2_n630 , 2_n642 , 2_n648 , 2_n656 , 2_n671 , 2_n680 , 2_n684 , 2_n690 , 2_n691 , 2_n693 , 2_n699 , 2_n702 , 2_n703 , 2_n704 , 2_n706 , 2_n716 , 2_n741 , 2_n742 , 2_n743 , 2_n746 , 2_n753 , 2_n756 , 2_n765 , 2_n777 , 2_n782 , 2_n788 );
    input 2_n5 , 2_n13 , 2_n17 , 2_n20 , 2_n36 , 2_n37 , 2_n53 , 2_n75 , 2_n80 , 2_n86 , 2_n93 , 2_n105 , 2_n106 , 2_n111 , 2_n117 , 2_n139 , 2_n147 , 2_n157 , 2_n161 , 2_n182 , 2_n190 , 2_n198 , 2_n204 , 2_n208 , 2_n214 , 2_n217 , 2_n219 , 2_n224 , 2_n226 , 2_n229 , 2_n235 , 2_n244 , 2_n249 , 2_n281 , 2_n287 , 2_n289 , 2_n300 , 2_n303 , 2_n319 , 2_n346 , 2_n364 , 2_n365 , 2_n368 , 2_n384 , 2_n393 , 2_n403 , 2_n409 , 2_n410 , 2_n417 , 2_n439 , 2_n457 , 2_n465 , 2_n473 , 2_n477 , 2_n503 , 2_n506 , 2_n511 , 2_n518 , 2_n521 , 2_n532 , 2_n537 , 2_n587 , 2_n588 , 2_n593 , 2_n594 , 2_n595 , 2_n606 , 2_n642 , 2_n648 , 2_n656 , 2_n671 , 2_n680 , 2_n684 , 2_n690 , 2_n693 , 2_n699 , 2_n702 , 2_n706 , 2_n716 , 2_n741 , 2_n742 , 2_n743 , 2_n746 , 2_n777 , 2_n782 , 2_n788 ;
    output 2_n27 , 2_n62 , 2_n145 , 2_n175 , 2_n176 , 2_n225 , 2_n241 , 2_n256 , 2_n294 , 2_n345 , 2_n387 , 2_n389 , 2_n430 , 2_n442 , 2_n489 , 2_n491 , 2_n493 , 2_n515 , 2_n618 , 2_n630 , 2_n691 , 2_n703 , 2_n704 , 2_n753 , 2_n756 , 2_n765 ;
    wire 2_n0 , 2_n1 , 2_n2 , 2_n3 , 2_n4 , 2_n6 , 2_n7 , 2_n8 , 2_n9 , 2_n10 , 2_n11 , 2_n12 , 2_n14 , 2_n15 , 2_n16 , 2_n18 , 2_n19 , 2_n21 , 2_n22 , 2_n23 , 2_n24 , 2_n25 , 2_n26 , 2_n28 , 2_n29 , 2_n30 , 2_n31 , 2_n32 , 2_n33 , 2_n34 , 2_n35 , 2_n38 , 2_n39 , 2_n40 , 2_n41 , 2_n42 , 2_n43 , 2_n44 , 2_n45 , 2_n46 , 2_n47 , 2_n48 , 2_n49 , 2_n50 , 2_n51 , 2_n52 , 2_n54 , 2_n55 , 2_n56 , 2_n57 , 2_n58 , 2_n59 , 2_n60 , 2_n61 , 2_n63 , 2_n64 , 2_n65 , 2_n66 , 2_n67 , 2_n68 , 2_n69 , 2_n70 , 2_n71 , 2_n72 , 2_n73 , 2_n74 , 2_n76 , 2_n77 , 2_n78 , 2_n79 , 2_n81 , 2_n82 , 2_n83 , 2_n84 , 2_n85 , 2_n87 , 2_n88 , 2_n89 , 2_n90 , 2_n91 , 2_n92 , 2_n94 , 2_n95 , 2_n96 , 2_n97 , 2_n98 , 2_n99 , 2_n100 , 2_n101 , 2_n102 , 2_n103 , 2_n104 , 2_n107 , 2_n108 , 2_n109 , 2_n110 , 2_n112 , 2_n113 , 2_n114 , 2_n115 , 2_n116 , 2_n118 , 2_n119 , 2_n120 , 2_n121 , 2_n122 , 2_n123 , 2_n124 , 2_n125 , 2_n126 , 2_n127 , 2_n128 , 2_n129 , 2_n130 , 2_n131 , 2_n132 , 2_n133 , 2_n134 , 2_n135 , 2_n136 , 2_n137 , 2_n138 , 2_n140 , 2_n141 , 2_n142 , 2_n143 , 2_n144 , 2_n146 , 2_n148 , 2_n149 , 2_n150 , 2_n151 , 2_n152 , 2_n153 , 2_n154 , 2_n155 , 2_n156 , 2_n158 , 2_n159 , 2_n160 , 2_n162 , 2_n163 , 2_n164 , 2_n165 , 2_n166 , 2_n167 , 2_n168 , 2_n169 , 2_n170 , 2_n171 , 2_n172 , 2_n173 , 2_n174 , 2_n177 , 2_n178 , 2_n179 , 2_n180 , 2_n181 , 2_n183 , 2_n184 , 2_n185 , 2_n186 , 2_n187 , 2_n188 , 2_n189 , 2_n191 , 2_n192 , 2_n193 , 2_n194 , 2_n195 , 2_n196 , 2_n197 , 2_n199 , 2_n200 , 2_n201 , 2_n202 , 2_n203 , 2_n205 , 2_n206 , 2_n207 , 2_n209 , 2_n210 , 2_n211 , 2_n212 , 2_n213 , 2_n215 , 2_n216 , 2_n218 , 2_n220 , 2_n221 , 2_n222 , 2_n223 , 2_n227 , 2_n228 , 2_n230 , 2_n231 , 2_n232 , 2_n233 , 2_n234 , 2_n236 , 2_n237 , 2_n238 , 2_n239 , 2_n240 , 2_n242 , 2_n243 , 2_n245 , 2_n246 , 2_n247 , 2_n248 , 2_n250 , 2_n251 , 2_n252 , 2_n253 , 2_n254 , 2_n255 , 2_n257 , 2_n258 , 2_n259 , 2_n260 , 2_n261 , 2_n262 , 2_n263 , 2_n264 , 2_n265 , 2_n266 , 2_n267 , 2_n268 , 2_n269 , 2_n270 , 2_n271 , 2_n272 , 2_n273 , 2_n274 , 2_n275 , 2_n276 , 2_n277 , 2_n278 , 2_n279 , 2_n280 , 2_n282 , 2_n283 , 2_n284 , 2_n285 , 2_n286 , 2_n288 , 2_n290 , 2_n291 , 2_n292 , 2_n293 , 2_n295 , 2_n296 , 2_n297 , 2_n298 , 2_n299 , 2_n301 , 2_n302 , 2_n304 , 2_n305 , 2_n306 , 2_n307 , 2_n308 , 2_n309 , 2_n310 , 2_n311 , 2_n312 , 2_n313 , 2_n314 , 2_n315 , 2_n316 , 2_n317 , 2_n318 , 2_n320 , 2_n321 , 2_n322 , 2_n323 , 2_n324 , 2_n325 , 2_n326 , 2_n327 , 2_n328 , 2_n329 , 2_n330 , 2_n331 , 2_n332 , 2_n333 , 2_n334 , 2_n335 , 2_n336 , 2_n337 , 2_n338 , 2_n339 , 2_n340 , 2_n341 , 2_n342 , 2_n343 , 2_n344 , 2_n347 , 2_n348 , 2_n349 , 2_n350 , 2_n351 , 2_n352 , 2_n353 , 2_n354 , 2_n355 , 2_n356 , 2_n357 , 2_n358 , 2_n359 , 2_n360 , 2_n361 , 2_n362 , 2_n363 , 2_n366 , 2_n367 , 2_n369 , 2_n370 , 2_n371 , 2_n372 , 2_n373 , 2_n374 , 2_n375 , 2_n376 , 2_n377 , 2_n378 , 2_n379 , 2_n380 , 2_n381 , 2_n382 , 2_n383 , 2_n385 , 2_n386 , 2_n388 , 2_n390 , 2_n391 , 2_n392 , 2_n394 , 2_n395 , 2_n396 , 2_n397 , 2_n398 , 2_n399 , 2_n400 , 2_n401 , 2_n402 , 2_n404 , 2_n405 , 2_n406 , 2_n407 , 2_n408 , 2_n411 , 2_n412 , 2_n413 , 2_n414 , 2_n415 , 2_n416 , 2_n418 , 2_n419 , 2_n420 , 2_n421 , 2_n422 , 2_n423 , 2_n424 , 2_n425 , 2_n426 , 2_n427 , 2_n428 , 2_n429 , 2_n431 , 2_n432 , 2_n433 , 2_n434 , 2_n435 , 2_n436 , 2_n437 , 2_n438 , 2_n440 , 2_n441 , 2_n443 , 2_n444 , 2_n445 , 2_n446 , 2_n447 , 2_n448 , 2_n449 , 2_n450 , 2_n451 , 2_n452 , 2_n453 , 2_n454 , 2_n455 , 2_n456 , 2_n458 , 2_n459 , 2_n460 , 2_n461 , 2_n462 , 2_n463 , 2_n464 , 2_n466 , 2_n467 , 2_n468 , 2_n469 , 2_n470 , 2_n471 , 2_n472 , 2_n474 , 2_n475 , 2_n476 , 2_n478 , 2_n479 , 2_n480 , 2_n481 , 2_n482 , 2_n483 , 2_n484 , 2_n485 , 2_n486 , 2_n487 , 2_n488 , 2_n490 , 2_n492 , 2_n494 , 2_n495 , 2_n496 , 2_n497 , 2_n498 , 2_n499 , 2_n500 , 2_n501 , 2_n502 , 2_n504 , 2_n505 , 2_n507 , 2_n508 , 2_n509 , 2_n510 , 2_n512 , 2_n513 , 2_n514 , 2_n516 , 2_n517 , 2_n519 , 2_n520 , 2_n522 , 2_n523 , 2_n524 , 2_n525 , 2_n526 , 2_n527 , 2_n528 , 2_n529 , 2_n530 , 2_n531 , 2_n533 , 2_n534 , 2_n535 , 2_n536 , 2_n538 , 2_n539 , 2_n540 , 2_n541 , 2_n542 , 2_n543 , 2_n544 , 2_n545 , 2_n546 , 2_n547 , 2_n548 , 2_n549 , 2_n550 , 2_n551 , 2_n552 , 2_n553 , 2_n554 , 2_n555 , 2_n556 , 2_n557 , 2_n558 , 2_n559 , 2_n560 , 2_n561 , 2_n562 , 2_n563 , 2_n564 , 2_n565 , 2_n566 , 2_n567 , 2_n568 , 2_n569 , 2_n570 , 2_n571 , 2_n572 , 2_n573 , 2_n574 , 2_n575 , 2_n576 , 2_n577 , 2_n578 , 2_n579 , 2_n580 , 2_n581 , 2_n582 , 2_n583 , 2_n584 , 2_n585 , 2_n586 , 2_n589 , 2_n590 , 2_n591 , 2_n592 , 2_n596 , 2_n597 , 2_n598 , 2_n599 , 2_n600 , 2_n601 , 2_n602 , 2_n603 , 2_n604 , 2_n605 , 2_n607 , 2_n608 , 2_n609 , 2_n610 , 2_n611 , 2_n612 , 2_n613 , 2_n614 , 2_n615 , 2_n616 , 2_n617 , 2_n619 , 2_n620 , 2_n621 , 2_n622 , 2_n623 , 2_n624 , 2_n625 , 2_n626 , 2_n627 , 2_n628 , 2_n629 , 2_n631 , 2_n632 , 2_n633 , 2_n634 , 2_n635 , 2_n636 , 2_n637 , 2_n638 , 2_n639 , 2_n640 , 2_n641 , 2_n643 , 2_n644 , 2_n645 , 2_n646 , 2_n647 , 2_n649 , 2_n650 , 2_n651 , 2_n652 , 2_n653 , 2_n654 , 2_n655 , 2_n657 , 2_n658 , 2_n659 , 2_n660 , 2_n661 , 2_n662 , 2_n663 , 2_n664 , 2_n665 , 2_n666 , 2_n667 , 2_n668 , 2_n669 , 2_n670 , 2_n672 , 2_n673 , 2_n674 , 2_n675 , 2_n676 , 2_n677 , 2_n678 , 2_n679 , 2_n681 , 2_n682 , 2_n683 , 2_n685 , 2_n686 , 2_n687 , 2_n688 , 2_n689 , 2_n692 , 2_n694 , 2_n695 , 2_n696 , 2_n697 , 2_n698 , 2_n700 , 2_n701 , 2_n705 , 2_n707 , 2_n708 , 2_n709 , 2_n710 , 2_n711 , 2_n712 , 2_n713 , 2_n714 , 2_n715 , 2_n717 , 2_n718 , 2_n719 , 2_n720 , 2_n721 , 2_n722 , 2_n723 , 2_n724 , 2_n725 , 2_n726 , 2_n727 , 2_n728 , 2_n729 , 2_n730 , 2_n731 , 2_n732 , 2_n733 , 2_n734 , 2_n735 , 2_n736 , 2_n737 , 2_n738 , 2_n739 , 2_n740 , 2_n744 , 2_n745 , 2_n747 , 2_n748 , 2_n749 , 2_n750 , 2_n751 , 2_n752 , 2_n754 , 2_n755 , 2_n757 , 2_n758 , 2_n759 , 2_n760 , 2_n761 , 2_n762 , 2_n763 , 2_n764 , 2_n766 , 2_n767 , 2_n768 , 2_n769 , 2_n770 , 2_n771 , 2_n772 , 2_n773 , 2_n774 , 2_n775 , 2_n776 , 2_n778 , 2_n779 , 2_n780 , 2_n781 , 2_n783 , 2_n784 , 2_n785 , 2_n786 , 2_n787 , 2_n789 ;
assign 2_n8 = 2_n559 | 2_n136;
assign 2_n676 = 2_n578 & 2_n778;
assign 2_n683 = ~(2_n403 | 2_n783);
assign 2_n213 = 2_n293 | 2_n774;
assign 2_n273 = ~(2_n300 | 2_n250);
assign 2_n34 = ~(2_n196 | 2_n40);
assign 2_n109 = 2_n787 & 2_n405;
assign 2_n122 = 2_n114 & 2_n600;
assign 2_n645 = ~(2_n452 | 2_n488);
assign 2_n621 = 2_n433 | 2_n106;
assign 2_n312 = 2_n381 | 2_n296;
assign 2_n534 = ~2_n226;
assign 2_n657 = 2_n341 | 2_n59;
assign 2_n6 = ~(2_n393 | 2_n447);
assign 2_n778 = ~2_n268;
assign 2_n673 = 2_n717 | 2_n737;
assign 2_n634 = 2_n692 & 2_n597;
assign 2_n719 = ~(2_n452 | 2_n655);
assign 2_n644 = ~(2_n475 ^ 2_n716);
assign 2_n323 = ~(2_n648 | 2_n223);
assign 2_n646 = ~2_n5;
assign 2_n369 = 2_n46 & 2_n230;
assign 2_n681 = ~2_n521;
assign 2_n411 = 2_n760 & 2_n88;
assign 2_n600 = ~(2_n656 | 2_n155);
assign 2_n698 = ~(2_n452 | 2_n552);
assign 2_n774 = 2_n656 & 2_n695;
assign 2_n311 = ~(2_n751 ^ 2_n680);
assign 2_n586 = 2_n391 | 2_n652;
assign 2_n206 = 2_n165 | 2_n153;
assign 2_n760 = ~2_n202;
assign 2_n628 = ~2_n157;
assign 2_n91 = 2_n165 & 2_n153;
assign 2_n493 = 2_n309 | 2_n12;
assign 2_n203 = 2_n38 | 2_n697;
assign 2_n375 = 2_n686 | 2_n772;
assign 2_n288 = 2_n150 | 2_n598;
assign 2_n268 = 2_n522 & 2_n443;
assign 2_n31 = 2_n459 | 2_n656;
assign 2_n415 = ~(2_n98 | 2_n363);
assign 2_n685 = 2_n546 | 2_n276;
assign 2_n63 = 2_n131 & 2_n627;
assign 2_n764 = 2_n656 & 2_n135;
assign 2_n707 = 2_n452 | 2_n761;
assign 2_n450 = 2_n666 & 2_n257;
assign 2_n52 = 2_n391 & 2_n767;
assign 2_n772 = 2_n452 | 2_n270;
assign 2_n252 = ~(2_n166 | 2_n189);
assign 2_n466 = 2_n75 & 2_n452;
assign 2_n399 = ~2_n603;
assign 2_n16 = 2_n42 & 2_n29;
assign 2_n207 = ~(2_n537 | 2_n212);
assign 2_n277 = 2_n581 & 2_n248;
assign 2_n407 = ~2_n749;
assign 2_n574 = 2_n607 | 2_n264;
assign 2_n383 = ~2_n520;
assign 2_n169 = ~2_n236;
assign 2_n97 = 2_n537 | 2_n300;
assign 2_n559 = ~2_n393;
assign 2_n14 = ~(2_n440 ^ 2_n19);
assign 2_n762 = ~(2_n484 | 2_n635);
assign 2_n589 = ~(2_n656 | 2_n568);
assign 2_n462 = 2_n42 | 2_n29;
assign 2_n110 = ~(2_n403 | 2_n590);
assign 2_n258 = 2_n331 | 2_n121;
assign 2_n257 = 2_n546 & 2_n757;
assign 2_n639 = 2_n16 | 2_n752;
assign 2_n661 = ~2_n351;
assign 2_n127 = ~2_n106;
assign 2_n655 = ~(2_n749 ^ 2_n163);
assign 2_n48 = ~(2_n656 | 2_n674);
assign 2_n678 = ~(2_n417 | 2_n550);
assign 2_n381 = ~2_n439;
assign 2_n65 = ~(2_n582 ^ 2_n788);
assign 2_n153 = 2_n609 & 2_n81;
assign 2_n615 = ~(2_n409 ^ 2_n642);
assign 2_n264 = ~2_n584;
assign 2_n452 = ~2_n656;
assign 2_n177 = ~(2_n643 ^ 2_n780);
assign 2_n200 = 2_n728 | 2_n694;
assign 2_n42 = 2_n591 & 2_n288;
assign 2_n173 = 2_n330 & 2_n599;
assign 2_n533 = ~(2_n452 | 2_n676);
assign 2_n269 = ~(2_n439 | 2_n117);
assign 2_n233 = 2_n559 | 2_n779;
assign 2_n167 = ~2_n300;
assign 2_n552 = ~(2_n228 ^ 2_n487);
assign 2_n76 = 2_n766 | 2_n158;
assign 2_n664 = ~2_n642;
assign 2_n471 = 2_n559 | 2_n436;
assign 2_n186 = ~2_n713;
assign 2_n456 = 2_n300 | 2_n106;
assign 2_n604 = ~(2_n656 | 2_n3);
assign 2_n557 = 2_n37 & 2_n501;
assign 2_n643 = 2_n460 | 2_n7;
assign 2_n56 = ~(2_n656 | 2_n140);
assign 2_n688 = ~2_n700;
assign 2_n519 = ~2_n17;
assign 2_n199 = 2_n362 & 2_n397;
assign 2_n602 = ~2_n786;
assign 2_n251 = 2_n127 | 2_n74;
assign 2_n766 = 2_n503 & 2_n182;
assign 2_n126 = ~2_n657;
assign 2_n185 = 2_n660 & 2_n441;
assign 2_n755 = 2_n202 | 2_n560;
assign 2_n154 = ~(2_n384 | 2_n129);
assign 2_n133 = ~(2_n693 | 2_n17);
assign 2_n659 = 2_n746 & 2_n127;
assign 2_n163 = 2_n152 & 2_n596;
assign 2_n274 = 2_n656 & 2_n776;
assign 2_n733 = ~(2_n214 | 2_n69);
assign 2_n514 = ~(2_n355 | 2_n536);
assign 2_n77 = 2_n656 & 2_n71;
assign 2_n336 = ~(2_n228 | 2_n372);
assign 2_n115 = ~(2_n452 | 2_n544);
assign 2_n376 = 2_n656 | 2_n563;
assign 2_n222 = ~2_n148;
assign 2_n597 = 2_n393 | 2_n454;
assign 2_n360 = 2_n356 | 2_n299;
assign 2_n228 = 2_n535 | 2_n274;
assign 2_n391 = ~2_n680;
assign 2_n636 = 2_n626 | 2_n641;
assign 2_n350 = 2_n458 | 2_n613;
assign 2_n170 = ~(2_n649 | 2_n376);
assign 2_n461 = ~(2_n350 | 2_n0);
assign 2_n181 = 2_n595 & 2_n452;
assign 2_n526 = 2_n767 ^ 2_n453;
assign 2_n316 = 2_n393 | 2_n508;
assign 2_n516 = ~(2_n439 ^ 2_n742);
assign 2_n686 = ~(2_n513 | 2_n28);
assign 2_n50 = 2_n218 & 2_n396;
assign 2_n168 = 2_n656 & 2_n444;
assign 2_n480 = ~2_n592;
assign 2_n70 = ~(2_n656 | 2_n631);
assign 2_n441 = ~2_n19;
assign 2_n549 = 2_n628 | 2_n340;
assign 2_n490 = 2_n228 & 2_n372;
assign 2_n497 = 2_n656 & 2_n408;
assign 2_n267 = 2_n403 & 2_n311;
assign 2_n174 = 2_n23 | 2_n520;
assign 2_n581 = ~2_n159;
assign 2_n30 = 2_n519 | 2_n423;
assign 2_n143 = 2_n366 & 2_n369;
assign 2_n502 = ~(2_n705 | 2_n251);
assign 2_n582 = 2_n125 | 2_n353;
assign 2_n380 = 2_n462 & 2_n639;
assign 2_n529 = ~(2_n656 | 2_n388);
assign 2_n736 = 2_n621 | 2_n553;
assign 2_n540 = ~(2_n759 | 2_n246);
assign 2_n607 = 2_n690 & 2_n217;
assign 2_n58 = 2_n687 | 2_n148;
assign 2_n404 = ~(2_n189 ^ 2_n61);
assign 2_n618 = 2_n589 | 2_n576;
assign 2_n763 = ~(2_n300 | 2_n789);
assign 2_n753 = 2_n47 | 2_n395;
assign 2_n561 = 2_n547 & 2_n260;
assign 2_n102 = ~(2_n452 | 2_n385);
assign 2_n29 = ~2_n68;
assign 2_n39 = ~(2_n452 | 2_n33);
assign 2_n292 = ~2_n287;
assign 2_n573 = ~(2_n440 | 2_n441);
assign 2_n354 = ~2_n330;
assign 2_n262 = 2_n525 | 2_n524;
assign 2_n197 = ~(2_n157 | 2_n303);
assign 2_n332 = 2_n174 & 2_n509;
assign 2_n396 = 2_n549 | 2_n374;
assign 2_n114 = 2_n297 | 2_n60;
assign 2_n520 = ~(2_n574 ^ 2_n690);
assign 2_n339 = ~(2_n527 | 2_n667);
assign 2_n25 = ~(2_n537 | 2_n286);
assign 2_n494 = ~(2_n724 | 2_n35);
assign 2_n592 = 2_n506 & 2_n169;
assign 2_n155 = ~(2_n495 | 2_n556);
assign 2_n241 = 2_n731 | 2_n698;
assign 2_n130 = ~(2_n76 ^ 2_n777);
assign 2_n270 = 2_n513 & 2_n28;
assign 2_n221 = 2_n518 & 2_n452;
assign 2_n717 = 2_n352 & 2_n516;
assign 2_n507 = ~(2_n726 | 2_n193);
assign 2_n726 = 2_n754 | 2_n497;
assign 2_n230 = 2_n608 & 2_n237;
assign 2_n385 = ~(2_n213 ^ 2_n230);
assign 2_n555 = ~(2_n17 ^ 2_n13);
assign 2_n340 = ~2_n303;
assign 2_n756 = 2_n386 | 2_n172;
assign 2_n560 = 2_n688 & 2_n314;
assign 2_n98 = ~(2_n78 | 2_n470);
assign 2_n322 = 2_n656 & 2_n344;
assign 2_n697 = 2_n403 | 2_n537;
assign 2_n565 = 2_n73 | 2_n446;
assign 2_n119 = ~(2_n787 | 2_n405);
assign 2_n663 = 2_n735 | 2_n200;
assign 2_n370 = ~(2_n185 | 2_n727);
assign 2_n256 = 2_n160 | 2_n321;
assign 2_n749 = 2_n632 | 2_n476;
assign 2_n694 = ~2_n76;
assign 2_n327 = 2_n127 | 2_n714;
assign 2_n735 = ~2_n281;
assign 2_n486 = ~(2_n452 | 2_n432);
assign 2_n132 = ~2_n200;
assign 2_n296 = ~2_n742;
assign 2_n525 = ~2_n648;
assign 2_n499 = ~(2_n300 | 2_n485);
assign 2_n227 = 2_n15 | 2_n668;
assign 2_n695 = ~(2_n236 ^ 2_n506);
assign 2_n725 = 2_n373 & 2_n101;
assign 2_n331 = ~2_n417;
assign 2_n438 = 2_n368 & 2_n452;
assign 2_n547 = ~2_n549;
assign 2_n400 = 2_n292 | 2_n656;
assign 2_n246 = ~(2_n355 ^ 2_n141);
assign 2_n701 = 2_n660 | 2_n19;
assign 2_n189 = 2_n32 | 2_n658;
assign 2_n476 = 2_n656 & 2_n770;
assign 2_n583 = 2_n44 | 2_n380;
assign 2_n566 = ~2_n636;
assign 2_n131 = 2_n412 | 2_n787;
assign 2_n530 = ~2_n299;
assign 2_n687 = ~2_n672;
assign 2_n789 = 2_n137 & 2_n327;
assign 2_n239 = 2_n608 | 2_n636;
assign 2_n348 = 2_n20 & 2_n57;
assign 2_n669 = 2_n666 | 2_n685;
assign 2_n46 = ~2_n213;
assign 2_n341 = 2_n161 & 2_n452;
assign 2_n286 = ~(2_n313 | 2_n763);
assign 2_n108 = ~(2_n350 ^ 2_n369);
assign 2_n771 = 2_n78 & 2_n470;
assign 2_n430 = 2_n494 | 2_n307;
assign 2_n609 = 2_n688 | 2_n164;
assign 2_n148 = 2_n407 | 2_n232;
assign 2_n775 = ~(2_n5 ^ 2_n157);
assign 2_n692 = 2_n559 | 2_n418;
assign 2_n32 = 2_n439 & 2_n117;
assign 2_n263 = ~(2_n258 ^ 2_n20);
assign 2_n454 = ~(2_n358 | 2_n482);
assign 2_n479 = ~2_n606;
assign 2_n255 = ~2_n490;
assign 2_n62 = 2_n604 | 2_n87;
assign 2_n489 = 2_n56 | 2_n102;
assign 2_n142 = 2_n559 | 2_n722;
assign 2_n193 = 2_n687 & 2_n392;
assign 2_n548 = ~(2_n759 | 2_n615);
assign 2_n278 = ~(2_n64 | 2_n625);
assign 2_n470 = 2_n495 | 2_n778;
assign 2_n202 = 2_n700 & 2_n164;
assign 2_n55 = 2_n244 & 2_n452;
assign 2_n469 = 2_n656 & 2_n65;
assign 2_n247 = 2_n547 | 2_n197;
assign 2_n144 = ~(2_n656 | 2_n496);
assign 2_n553 = 2_n272 | 2_n97;
assign 2_n750 = 2_n24 & 2_n193;
assign 2_n329 = 2_n532 & 2_n452;
assign 2_n632 = 2_n743 & 2_n452;
assign 2_n611 = 2_n715 & 2_n623;
assign 2_n220 = 2_n702 & 2_n452;
assign 2_n405 = ~(2_n184 ^ 2_n422);
assign 2_n759 = ~2_n537;
assign 2_n343 = 2_n116 | 2_n603;
assign 2_n483 = ~(2_n159 ^ 2_n248);
assign 2_n345 = 2_n144 | 2_n696;
assign 2_n712 = 2_n14 & 2_n173;
assign 2_n95 = 2_n429 | 2_n539;
assign 2_n183 = ~2_n706;
assign 2_n458 = 2_n224 & 2_n452;
assign 2_n783 = ~(2_n577 | 2_n207);
assign 2_n603 = 2_n24 | 2_n58;
assign 2_n758 = ~2_n384;
assign 2_n211 = ~(2_n94 | 2_n169);
assign 2_n652 = ~2_n594;
assign 2_n382 = 2_n455 | 2_n747;
assign 2_n569 = ~(2_n452 | 2_n10);
assign 2_n429 = 2_n235 & 2_n452;
assign 2_n721 = 2_n46 | 2_n239;
assign 2_n242 = ~(2_n540 | 2_n191);
assign 2_n492 = 2_n300 & 2_n404;
assign 2_n445 = ~(2_n439 ^ 2_n117);
assign 2_n435 = ~(2_n700 ^ 2_n314);
assign 2_n640 = 2_n412 & 2_n787;
assign 2_n41 = 2_n662 | 2_n480;
assign 2_n402 = 2_n400 & 2_n375;
assign 2_n201 = ~(2_n377 | 2_n647);
assign 2_n421 = ~(2_n284 | 2_n380);
assign 2_n724 = 2_n617 & 2_n638;
assign 2_n428 = 2_n184 & 2_n240;
assign 2_n413 = ~(2_n349 ^ 2_n445);
assign 2_n243 = 2_n452 | 2_n379;
assign 2_n660 = ~2_n440;
assign 2_n424 = 2_n620 | 2_n178;
assign 2_n146 = ~2_n190;
assign 2_n704 = 2_n624 | 2_n533;
assign 2_n362 = 2_n472 | 2_n335;
assign 2_n158 = ~(2_n720 | 2_n28);
assign 2_n614 = ~2_n582;
assign 2_n123 = ~(2_n217 ^ 2_n365);
assign 2_n770 = ~(2_n154 | 2_n661);
assign 2_n718 = ~2_n663;
assign 2_n576 = 2_n206 & 2_n134;
assign 2_n527 = ~2_n382;
assign 2_n45 = ~(2_n298 | 2_n718);
assign 2_n24 = ~2_n726;
assign 2_n658 = ~(2_n349 | 2_n269);
assign 2_n769 = 2_n610 | 2_n650;
assign 2_n113 = ~2_n685;
assign 2_n28 = 2_n586 & 2_n781;
assign 2_n1 = ~(2_n452 | 2_n177);
assign 2_n596 = 2_n185 | 2_n173;
assign 2_n196 = ~(2_n741 | 2_n713);
assign 2_n440 = 2_n221 | 2_n261;
assign 2_n408 = ~(2_n323 | 2_n390);
assign 2_n612 = ~(2_n36 | 2_n348);
assign 2_n460 = 2_n587 & 2_n452;
assign 2_n482 = ~(2_n403 | 2_n242);
assign 2_n103 = ~2_n669;
assign 2_n238 = 2_n249 & 2_n439;
assign 2_n394 = ~2_n564;
assign 2_n558 = ~2_n214;
assign 2_n500 = 2_n120 & 2_n748;
assign 2_n578 = 2_n522 | 2_n443;
assign 2_n156 = 2_n336 | 2_n490;
assign 2_n554 = ~2_n741;
assign 2_n416 = ~(2_n367 | 2_n171);
assign 2_n0 = ~2_n721;
assign 2_n101 = 2_n478 | 2_n290;
assign 2_n727 = ~2_n152;
assign 2_n314 = 2_n481 & 2_n85;
assign 2_n129 = 2_n699 & 2_n718;
assign 2_n512 = 2_n364 & 2_n452;
assign 2_n508 = ~(2_n267 | 2_n110);
assign 2_n317 = ~(2_n619 ^ 2_n503);
assign 2_n149 = ~(2_n656 | 2_n538);
assign 2_n23 = ~2_n503;
assign 2_n682 = ~(2_n700 | 2_n314);
assign 2_n544 = ~(2_n505 ^ 2_n257);
assign 2_n635 = 2_n656 | 2_n2;
assign 2_n517 = ~(2_n359 | 2_n128);
assign 2_n780 = 2_n179 & 2_n487;
assign 2_n89 = 2_n628 | 2_n739;
assign 2_n225 = 2_n271 | 2_n531;
assign 2_n351 = 2_n758 | 2_n320;
assign 2_n356 = ~2_n245;
assign 2_n309 = ~(2_n461 | 2_n670);
assign 2_n218 = 2_n646 | 2_n107;
assign 2_n231 = ~2_n402;
assign 2_n412 = ~2_n184;
assign 2_n324 = ~2_n69;
assign 2_n371 = ~(2_n657 ^ 2_n567);
assign 2_n732 = 2_n537 & 2_n304;
assign 2_n359 = 2_n473 & 2_n127;
assign 2_n484 = 2_n435 & 2_n285;
assign 2_n54 = ~(2_n495 ^ 2_n268);
assign 2_n118 = ~(2_n749 ^ 2_n49);
assign 2_n605 = 2_n428 | 2_n580;
assign 2_n487 = 2_n116 & 2_n750;
assign 2_n398 = 2_n416 | 2_n113;
assign 2_n357 = ~(2_n334 | 2_n354);
assign 2_n740 = 2_n157 & 2_n393;
assign 2_n84 = 2_n343 & 2_n529;
assign 2_n307 = ~(2_n452 | 2_n26);
assign 2_n786 = 2_n558 | 2_n324;
assign 2_n776 = ~(2_n678 | 2_n57);
assign 2_n297 = ~2_n495;
assign 2_n443 = 2_n356 & 2_n143;
assign 2_n590 = ~(2_n732 | 2_n572);
assign 2_n510 = 2_n229 & 2_n452;
assign 2_n260 = 2_n5 ^ 2_n671;
assign 2_n531 = ~(2_n452 | 2_n679);
assign 2_n501 = 2_n53 & 2_n602;
assign 2_n74 = 2_n30 & 2_n729;
assign 2_n620 = 2_n503 & 2_n611;
assign 2_n389 = 2_n72 | 2_n543;
assign 2_n321 = ~(2_n452 | 2_n483);
assign 2_n768 = ~2_n240;
assign 2_n22 = 2_n55 | 2_n708;
assign 2_n236 = 2_n681 | 2_n4;
assign 2_n378 = 2_n14 | 2_n173;
assign 2_n349 = 2_n664 | 2_n479;
assign 2_n495 = 2_n310 | 2_n83;
assign 2_n641 = ~2_n446;
assign 2_n67 = ~(2_n284 | 2_n420);
assign 2_n172 = ~(2_n452 | 2_n371);
assign 2_n432 = ~(2_n629 ^ 2_n755);
assign 2_n81 = 2_n682 | 2_n21;
assign 2_n474 = ~(2_n78 ^ 2_n114);
assign 2_n747 = ~(2_n452 | 2_n247);
assign 2_n290 = 2_n51 & 2_n504;
assign 2_n209 = ~(2_n672 | 2_n222);
assign 2_n73 = ~(2_n159 | 2_n318);
assign 2_n406 = ~(2_n663 ^ 2_n699);
assign 2_n3 = ~(2_n290 ^ 2_n67);
assign 2_n59 = 2_n656 & 2_n644;
assign 2_n505 = 2_n512 | 2_n469;
assign 2_n308 = ~(2_n672 ^ 2_n392);
assign 2_n444 = ~(2_n612 | 2_n614);
assign 2_n35 = 2_n656 | 2_n11;
assign 2_n546 = ~2_n367;
assign 2_n737 = 2_n127 | 2_n315;
assign 2_n386 = 2_n419 & 2_n434;
assign 2_n330 = 2_n472 | 2_n677;
assign 2_n134 = ~(2_n452 | 2_n91);
assign 2_n730 = ~2_n41;
assign 2_n773 = ~(2_n452 | 2_n130);
assign 2_n467 = ~(2_n657 | 2_n563);
assign 2_n622 = ~(2_n452 | 2_n712);
assign 2_n223 = 2_n457 & 2_n661;
assign 2_n591 = 2_n183 | 2_n656;
assign 2_n691 = 2_n9 | 2_n415;
assign 2_n302 = 2_n42 & 2_n68;
assign 2_n434 = ~(2_n656 | 2_n467);
assign 2_n138 = 2_n656 | 2_n556;
assign 2_n145 = 2_n84 | 2_n39;
assign 2_n675 = ~(2_n505 ^ 2_n113);
assign 2_n433 = ~2_n319;
assign 2_n472 = ~2_n283;
assign 2_n563 = ~2_n333;
assign 2_n51 = 2_n42 | 2_n68;
assign 2_n187 = 2_n220 | 2_n99;
assign 2_n668 = 2_n347 | 2_n266;
assign 2_n723 = ~(2_n95 ^ 2_n450);
assign 2_n535 = 2_n465 & 2_n452;
assign 2_n9 = ~(2_n656 | 2_n474);
assign 2_n191 = ~(2_n537 | 2_n431);
assign 2_n387 = 2_n170 | 2_n637;
assign 2_n475 = 2_n554 | 2_n186;
assign 2_n513 = ~(2_n503 ^ 2_n182);
assign 2_n528 = ~2_n574;
assign 2_n192 = ~(2_n167 | 2_n413);
assign 2_n667 = 2_n740 | 2_n295;
assign 2_n250 = 2_n90 & 2_n673;
assign 2_n66 = 2_n534 | 2_n656;
assign 2_n305 = 2_n522 & 2_n360;
assign 2_n100 = 2_n785 & 2_n424;
assign 2_n585 = 2_n656 & 2_n45;
assign 2_n254 = ~(2_n187 | 2_n566);
assign 2_n333 = 2_n275 | 2_n669;
assign 2_n104 = ~(2_n680 ^ 2_n594);
assign 2_n551 = ~(2_n786 ^ 2_n53);
assign 2_n754 = 2_n588 & 2_n452;
assign 2_n152 = 2_n660 | 2_n441;
assign 2_n69 = 2_n208 & 2_n730;
assign 2_n784 = ~2_n111;
assign 2_n447 = ~(2_n403 | 2_n18);
assign 2_n64 = 2_n693 & 2_n17;
assign 2_n781 = 2_n280 | 2_n50;
assign 2_n194 = ~2_n210;
assign 2_n373 = 2_n402 | 2_n210;
assign 2_n463 = ~(2_n367 ^ 2_n757);
assign 2_n175 = 2_n768 | 2_n339;
assign 2_n377 = ~(2_n17 | 2_n782);
assign 2_n610 = ~(2_n37 | 2_n501);
assign 2_n779 = ~(2_n332 ^ 2_n43);
assign 2_n26 = ~(2_n605 ^ 2_n616);
assign 2_n488 = 2_n44 & 2_n380;
assign 2_n99 = 2_n656 & 2_n211;
assign 2_n347 = 2_n393 | 2_n403;
assign 2_n283 = 2_n151 | 2_n585;
assign 2_n353 = ~2_n348;
assign 2_n703 = 2_n48 | 2_n1;
assign 2_n729 = 2_n312 & 2_n326;
assign 2_n291 = ~(2_n642 ^ 2_n606);
assign 2_n638 = ~(2_n42 ^ 2_n29);
assign 2_n448 = ~(2_n283 | 2_n677);
assign 2_n248 = 2_n126 & 2_n567;
assign 2_n679 = ~(2_n245 ^ 2_n143);
assign 2_n395 = ~(2_n452 | 2_n451);
assign 2_n625 = 2_n238 | 2_n514;
assign 2_n71 = ~(2_n162 ^ 2_n147);
assign 2_n731 = ~(2_n656 | 2_n156);
assign 2_n38 = ~2_n93;
assign 2_n363 = 2_n452 | 2_n771;
assign 2_n124 = ~(2_n739 | 2_n279);
assign 2_n374 = ~(2_n5 | 2_n671);
assign 2_n538 = ~(2_n188 ^ 2_n446);
assign 2_n426 = ~(2_n555 | 2_n729);
assign 2_n579 = 2_n656 | 2_n109;
assign 2_n295 = 2_n89 & 2_n6;
assign 2_n584 = 2_n449 | 2_n265;
assign 2_n650 = 2_n452 | 2_n557;
assign 2_n15 = 2_n711 | 2_n106;
assign 2_n313 = ~(2_n167 | 2_n291);
assign 2_n82 = ~(2_n184 | 2_n240);
assign 2_n536 = ~(2_n249 | 2_n439);
assign 2_n710 = ~(2_n633 | 2_n730);
assign 2_n361 = 2_n573 | 2_n199;
assign 2_n564 = 2_n716 & 2_n40;
assign 2_n392 = 2_n407 & 2_n163;
assign 2_n121 = ~2_n550;
assign 2_n491 = 2_n70 | 2_n498;
assign 2_n179 = ~2_n228;
assign 2_n562 = ~(2_n452 | 2_n54);
assign 2_n623 = 2_n52 | 2_n123;
assign 2_n33 = ~(2_n22 ^ 2_n750);
assign 2_n180 = 2_n147 & 2_n523;
assign 2_n285 = ~2_n725;
assign 2_n68 = 2_n112 & 2_n316;
assign 2_n478 = ~(2_n231 | 2_n194);
assign 2_n498 = ~(2_n507 | 2_n243);
assign 2_n715 = 2_n391 | 2_n767;
assign 2_n320 = ~2_n129;
assign 2_n677 = ~2_n335;
assign 2_n92 = ~2_n511;
assign 2_n79 = 2_n104 & 2_n50;
assign 2_n212 = ~(2_n201 | 2_n499);
assign 2_n575 = ~(2_n188 ^ 2_n277);
assign 2_n326 = 2_n352 | 2_n216;
assign 2_n713 = 2_n788 & 2_n614;
assign 2_n709 = ~2_n643;
assign 2_n437 = 2_n393 | 2_n651;
assign 2_n379 = 2_n726 & 2_n193;
assign 2_n275 = ~2_n95;
assign 2_n116 = ~2_n22;
assign 2_n388 = ~(2_n22 | 2_n399);
assign 2_n310 = 2_n410 & 2_n452;
assign 2_n556 = ~2_n60;
assign 2_n651 = ~(2_n601 | 2_n683);
assign 2_n601 = 2_n403 & 2_n317;
assign 2_n335 = 2_n736 & 2_n233;
assign 2_n739 = ~2_n403;
assign 2_n276 = 2_n709 | 2_n255;
assign 2_n515 = 2_n653 | 2_n719;
assign 2_n481 = 2_n393 | 2_n427;
assign 2_n571 = 2_n656 & 2_n195;
assign 2_n617 = ~2_n63;
assign 2_n696 = 2_n378 & 2_n622;
assign 2_n464 = ~(2_n452 | 2_n575);
assign 2_n245 = 2_n466 | 2_n571;
assign 2_n672 = 2_n438 | 2_n322;
assign 2_n504 = 2_n302 | 2_n63;
assign 2_n176 = 2_n762 | 2_n486;
assign 2_n271 = ~(2_n656 | 2_n541);
assign 2_n419 = 2_n126 | 2_n333;
assign 2_n522 = 2_n31 & 2_n707;
assign 2_n165 = ~(2_n283 ^ 2_n335);
assign 2_n670 = 2_n656 | 2_n530;
assign 2_n11 = ~(2_n617 | 2_n638);
assign 2_n261 = 2_n656 & 2_n406;
assign 2_n568 = ~(2_n411 ^ 2_n357);
assign 2_n150 = ~(2_n104 | 2_n50);
assign 2_n141 = ~(2_n249 ^ 2_n439);
assign 2_n662 = ~2_n86;
assign 2_n734 = ~2_n58;
assign 2_n40 = ~2_n475;
assign 2_n401 = ~(2_n262 ^ 2_n204);
assign 2_n397 = 2_n448 | 2_n411;
assign 2_n112 = 2_n559 | 2_n526;
assign 2_n334 = 2_n472 & 2_n677;
assign 2_n567 = 2_n275 & 2_n450;
assign 2_n572 = ~(2_n537 | 2_n328);
assign 2_n171 = ~2_n276;
assign 2_n294 = 2_n342 | 2_n115;
assign 2_n748 = ~(2_n452 | 2_n561);
assign 2_n509 = 2_n205 | 2_n100;
assign 2_n159 = 2_n329 | 2_n764;
assign 2_n272 = 2_n393 | 2_n403;
assign 2_n352 = 2_n664 | 2_n784;
assign 2_n282 = ~(2_n456 | 2_n203);
assign 2_n19 = 2_n227 & 2_n142;
assign 2_n94 = ~(2_n521 | 2_n180);
assign 2_n580 = ~(2_n82 | 2_n422);
assign 2_n279 = 2_n23 | 2_n619;
assign 2_n280 = ~(2_n680 | 2_n594);
assign 2_n7 = 2_n656 & 2_n263;
assign 2_n616 = ~(2_n42 ^ 2_n68);
assign 2_n265 = ~2_n365;
assign 2_n423 = ~2_n13;
assign 2_n751 = 2_n646 | 2_n628;
assign 2_n523 = ~2_n162;
assign 2_n425 = ~(2_n452 | 2_n463);
assign 2_n125 = ~2_n36;
assign 2_n372 = ~2_n343;
assign 2_n253 = 2_n346 & 2_n452;
assign 2_n665 = ~(2_n693 ^ 2_n17);
assign 2_n160 = ~(2_n656 | 2_n565);
assign 2_n633 = ~(2_n86 | 2_n592);
assign 2_n627 = 2_n640 | 2_n634;
assign 2_n195 = ~(2_n41 ^ 2_n208);
assign 2_n390 = ~2_n262;
assign 2_n446 = 2_n159 & 2_n318;
assign 2_n631 = ~(2_n726 ^ 2_n734);
assign 2_n542 = ~2_n239;
assign 2_n711 = ~2_n139;
assign 2_n577 = ~(2_n133 | 2_n325);
assign 2_n87 = 2_n583 & 2_n645;
assign 2_n708 = 2_n656 & 2_n401;
assign 2_n744 = ~(2_n178 ^ 2_n503);
assign 2_n599 = 2_n334 | 2_n153;
assign 2_n598 = 2_n452 | 2_n79;
assign 2_n43 = 2_n215 | 2_n528;
assign 2_n761 = 2_n733 | 2_n602;
assign 2_n422 = ~2_n634;
assign 2_n78 = 2_n66 & 2_n769;
assign 2_n366 = ~2_n350;
assign 2_n757 = 2_n709 & 2_n780;
assign 2_n418 = ~(2_n5 ^ 2_n365);
assign 2_n649 = ~(2_n95 | 2_n103);
assign 2_n284 = 2_n402 & 2_n194;
assign 2_n215 = ~2_n690;
assign 2_n414 = ~2_n409;
assign 2_n720 = ~(2_n503 | 2_n182);
assign 2_n451 = ~(2_n240 ^ 2_n405);
assign 2_n442 = 2_n122 | 2_n562;
assign 2_n325 = 2_n759 | 2_n278;
assign 2_n745 = ~(2_n300 | 2_n517);
assign 2_n107 = ~2_n671;
assign 2_n626 = ~2_n188;
assign 2_n240 = 2_n382 | 2_n689;
assign 2_n420 = 2_n231 & 2_n210;
assign 2_n135 = ~(2_n545 | 2_n523);
assign 2_n301 = 2_n127 | 2_n738;
assign 2_n674 = ~(2_n643 ^ 2_n490);
assign 2_n44 = ~(2_n231 ^ 2_n210);
assign 2_n96 = ~(2_n306 | 2_n100);
assign 2_n205 = ~(2_n503 | 2_n383);
assign 2_n315 = ~(2_n352 | 2_n516);
assign 2_n367 = 2_n181 | 2_n168;
assign 2_n57 = ~2_n258;
assign 2_n705 = ~(2_n17 | 2_n13);
assign 2_n61 = ~(2_n17 ^ 2_n782);
assign 2_n550 = 2_n204 & 2_n390;
assign 2_n624 = ~(2_n305 | 2_n138);
assign 2_n164 = ~2_n314;
assign 2_n714 = ~(2_n642 ^ 2_n111);
assign 2_n468 = ~2_n289;
assign 2_n47 = ~(2_n119 | 2_n579);
assign 2_n608 = ~2_n187;
assign 2_n647 = 2_n167 | 2_n252;
assign 2_n629 = 2_n420 | 2_n421;
assign 2_n700 = 2_n253 | 2_n773;
assign 2_n630 = 2_n234 | 2_n425;
assign 2_n654 = ~(2_n209 | 2_n734);
assign 2_n216 = ~(2_n439 | 2_n742);
assign 2_n293 = 2_n80 & 2_n452;
assign 2_n266 = 2_n537 | 2_n300;
assign 2_n728 = ~2_n777;
assign 2_n128 = ~(2_n426 | 2_n301);
assign 2_n449 = ~2_n217;
assign 2_n689 = ~2_n667;
assign 2_n337 = 2_n593 & 2_n452;
assign 2_n2 = ~(2_n435 | 2_n285);
assign 2_n765 = 2_n338 | 2_n569;
assign 2_n162 = 2_n146 | 2_n394;
assign 2_n140 = ~(2_n213 ^ 2_n542);
assign 2_n436 = 2_n306 & 2_n100;
assign 2_n338 = ~(2_n656 | 2_n570);
assign 2_n237 = 2_n626 & 2_n277;
assign 2_n136 = ~(2_n611 ^ 2_n744);
assign 2_n752 = ~2_n605;
assign 2_n619 = 2_n391 | 2_n751;
assign 2_n18 = 2_n548 | 2_n25;
assign 2_n485 = ~(2_n659 | 2_n502);
assign 2_n543 = ~(2_n452 | 2_n308);
assign 2_n342 = ~(2_n656 | 2_n675);
assign 2_n4 = ~2_n180;
assign 2_n539 = 2_n656 & 2_n34;
assign 2_n431 = ~(2_n192 | 2_n273);
assign 2_n455 = 2_n684 & 2_n452;
assign 2_n90 = 2_n92 | 2_n106;
assign 2_n137 = 2_n468 | 2_n106;
assign 2_n304 = ~(2_n625 ^ 2_n665);
assign 2_n232 = 2_n701 & 2_n361;
assign 2_n85 = 2_n96 | 2_n471;
assign 2_n785 = 2_n503 | 2_n611;
assign 2_n27 = 2_n149 | 2_n464;
assign 2_n666 = ~2_n505;
assign 2_n210 = 2_n437 & 2_n8;
assign 2_n358 = ~(2_n739 | 2_n775);
assign 2_n496 = ~(2_n199 ^ 2_n370);
assign 2_n21 = ~2_n629;
assign 2_n184 = 2_n337 | 2_n500;
assign 2_n259 = ~(2_n584 ^ 2_n217);
assign 2_n541 = ~(2_n245 ^ 2_n530);
assign 2_n298 = ~(2_n281 | 2_n132);
assign 2_n49 = ~2_n232;
assign 2_n10 = ~(2_n187 ^ 2_n237);
assign 2_n299 = 2_n366 | 2_n721;
assign 2_n722 = 2_n43 | 2_n332;
assign 2_n88 = 2_n560 | 2_n725;
assign 2_n344 = ~(2_n351 ^ 2_n457);
assign 2_n12 = ~(2_n452 | 2_n108);
assign 2_n188 = 2_n510 | 2_n77;
assign 2_n653 = ~(2_n656 | 2_n118);
assign 2_n459 = ~2_n105;
assign 2_n178 = ~(2_n259 ^ 2_n690);
assign 2_n427 = ~(2_n124 | 2_n282);
assign 2_n328 = ~(2_n492 | 2_n745);
assign 2_n355 = 2_n414 | 2_n664;
assign 2_n545 = ~(2_n190 | 2_n564);
assign 2_n767 = 2_n646 | 2_n265;
assign 2_n613 = 2_n656 & 2_n710;
assign 2_n120 = 2_n547 | 2_n260;
assign 2_n570 = 2_n254 | 2_n542;
assign 2_n318 = ~2_n419;
assign 2_n151 = 2_n219 & 2_n452;
assign 2_n637 = ~(2_n452 | 2_n723);
assign 2_n306 = ~(2_n383 ^ 2_n503);
assign 2_n453 = ~(2_n123 ^ 2_n680);
assign 2_n524 = ~2_n223;
assign 2_n787 = 2_n527 | 2_n689;
assign 2_n72 = 2_n452 & 2_n654;
assign 2_n234 = ~(2_n656 | 2_n398);
assign 2_n166 = 2_n17 & 2_n782;
assign 2_n60 = 2_n522 | 2_n360;
assign 2_n738 = 2_n555 & 2_n729;
assign 2_n83 = 2_n656 & 2_n551;
endmodule
