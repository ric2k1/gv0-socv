module top(in1, in2, in3, out1);
  input [31:0] in1, in2, in3;
  output [64:0] out1;
  wire [31:0] in1, in2, in3;
  wire [64:0] out1;
  wire csa_tree_add_6_33_groupi_n_0, csa_tree_add_6_33_groupi_n_1, csa_tree_add_6_33_groupi_n_17, csa_tree_add_6_33_groupi_n_18, csa_tree_add_6_33_groupi_n_19, csa_tree_add_6_33_groupi_n_20, csa_tree_add_6_33_groupi_n_21, csa_tree_add_6_33_groupi_n_22;
  wire csa_tree_add_6_33_groupi_n_23, csa_tree_add_6_33_groupi_n_24, csa_tree_add_6_33_groupi_n_25, csa_tree_add_6_33_groupi_n_26, csa_tree_add_6_33_groupi_n_27, csa_tree_add_6_33_groupi_n_28, csa_tree_add_6_33_groupi_n_29, csa_tree_add_6_33_groupi_n_30;
  wire csa_tree_add_6_33_groupi_n_31, csa_tree_add_6_33_groupi_n_32, csa_tree_add_6_33_groupi_n_33, csa_tree_add_6_33_groupi_n_34, csa_tree_add_6_33_groupi_n_35, csa_tree_add_6_33_groupi_n_36, csa_tree_add_6_33_groupi_n_37, csa_tree_add_6_33_groupi_n_38;
  wire csa_tree_add_6_33_groupi_n_39, csa_tree_add_6_33_groupi_n_40, csa_tree_add_6_33_groupi_n_41, csa_tree_add_6_33_groupi_n_42, csa_tree_add_6_33_groupi_n_43, csa_tree_add_6_33_groupi_n_44, csa_tree_add_6_33_groupi_n_45, csa_tree_add_6_33_groupi_n_46;
  wire csa_tree_add_6_33_groupi_n_47, csa_tree_add_6_33_groupi_n_48, csa_tree_add_6_33_groupi_n_49, csa_tree_add_6_33_groupi_n_50, csa_tree_add_6_33_groupi_n_51, csa_tree_add_6_33_groupi_n_52, csa_tree_add_6_33_groupi_n_53, csa_tree_add_6_33_groupi_n_54;
  wire csa_tree_add_6_33_groupi_n_55, csa_tree_add_6_33_groupi_n_56, csa_tree_add_6_33_groupi_n_57, csa_tree_add_6_33_groupi_n_58, csa_tree_add_6_33_groupi_n_59, csa_tree_add_6_33_groupi_n_60, csa_tree_add_6_33_groupi_n_61, csa_tree_add_6_33_groupi_n_62;
  wire csa_tree_add_6_33_groupi_n_63, csa_tree_add_6_33_groupi_n_64, csa_tree_add_6_33_groupi_n_65, csa_tree_add_6_33_groupi_n_66, csa_tree_add_6_33_groupi_n_67, csa_tree_add_6_33_groupi_n_68, csa_tree_add_6_33_groupi_n_69, csa_tree_add_6_33_groupi_n_70;
  wire csa_tree_add_6_33_groupi_n_71, csa_tree_add_6_33_groupi_n_72, csa_tree_add_6_33_groupi_n_73, csa_tree_add_6_33_groupi_n_74, csa_tree_add_6_33_groupi_n_75, csa_tree_add_6_33_groupi_n_76, csa_tree_add_6_33_groupi_n_77, csa_tree_add_6_33_groupi_n_78;
  wire csa_tree_add_6_33_groupi_n_79, csa_tree_add_6_33_groupi_n_80, csa_tree_add_6_33_groupi_n_81, csa_tree_add_6_33_groupi_n_82, csa_tree_add_6_33_groupi_n_83, csa_tree_add_6_33_groupi_n_84, csa_tree_add_6_33_groupi_n_85, csa_tree_add_6_33_groupi_n_86;
  wire csa_tree_add_6_33_groupi_n_87, csa_tree_add_6_33_groupi_n_88, csa_tree_add_6_33_groupi_n_89, csa_tree_add_6_33_groupi_n_90, csa_tree_add_6_33_groupi_n_91, csa_tree_add_6_33_groupi_n_92, csa_tree_add_6_33_groupi_n_93, csa_tree_add_6_33_groupi_n_94;
  wire csa_tree_add_6_33_groupi_n_95, csa_tree_add_6_33_groupi_n_96, csa_tree_add_6_33_groupi_n_97, csa_tree_add_6_33_groupi_n_98, csa_tree_add_6_33_groupi_n_99, csa_tree_add_6_33_groupi_n_100, csa_tree_add_6_33_groupi_n_101, csa_tree_add_6_33_groupi_n_102;
  wire csa_tree_add_6_33_groupi_n_103, csa_tree_add_6_33_groupi_n_104, csa_tree_add_6_33_groupi_n_105, csa_tree_add_6_33_groupi_n_106, csa_tree_add_6_33_groupi_n_107, csa_tree_add_6_33_groupi_n_108, csa_tree_add_6_33_groupi_n_109, csa_tree_add_6_33_groupi_n_110;
  wire csa_tree_add_6_33_groupi_n_111, csa_tree_add_6_33_groupi_n_112, csa_tree_add_6_33_groupi_n_113, csa_tree_add_6_33_groupi_n_114, csa_tree_add_6_33_groupi_n_115, csa_tree_add_6_33_groupi_n_116, csa_tree_add_6_33_groupi_n_117, csa_tree_add_6_33_groupi_n_118;
  wire csa_tree_add_6_33_groupi_n_119, csa_tree_add_6_33_groupi_n_120, csa_tree_add_6_33_groupi_n_121, csa_tree_add_6_33_groupi_n_122, csa_tree_add_6_33_groupi_n_123, csa_tree_add_6_33_groupi_n_124, csa_tree_add_6_33_groupi_n_125, csa_tree_add_6_33_groupi_n_126;
  wire csa_tree_add_6_33_groupi_n_127, csa_tree_add_6_33_groupi_n_128, csa_tree_add_6_33_groupi_n_129, csa_tree_add_6_33_groupi_n_130, csa_tree_add_6_33_groupi_n_131, csa_tree_add_6_33_groupi_n_132, csa_tree_add_6_33_groupi_n_133, csa_tree_add_6_33_groupi_n_134;
  wire csa_tree_add_6_33_groupi_n_135, csa_tree_add_6_33_groupi_n_136, csa_tree_add_6_33_groupi_n_137, csa_tree_add_6_33_groupi_n_138, csa_tree_add_6_33_groupi_n_139, csa_tree_add_6_33_groupi_n_140, csa_tree_add_6_33_groupi_n_141, csa_tree_add_6_33_groupi_n_142;
  wire csa_tree_add_6_33_groupi_n_143, csa_tree_add_6_33_groupi_n_144, csa_tree_add_6_33_groupi_n_145, csa_tree_add_6_33_groupi_n_146, csa_tree_add_6_33_groupi_n_147, csa_tree_add_6_33_groupi_n_148, csa_tree_add_6_33_groupi_n_149, csa_tree_add_6_33_groupi_n_150;
  wire csa_tree_add_6_33_groupi_n_151, csa_tree_add_6_33_groupi_n_152, csa_tree_add_6_33_groupi_n_153, csa_tree_add_6_33_groupi_n_154, csa_tree_add_6_33_groupi_n_155, csa_tree_add_6_33_groupi_n_156, csa_tree_add_6_33_groupi_n_157, csa_tree_add_6_33_groupi_n_158;
  wire csa_tree_add_6_33_groupi_n_159, csa_tree_add_6_33_groupi_n_160, csa_tree_add_6_33_groupi_n_161, csa_tree_add_6_33_groupi_n_162, csa_tree_add_6_33_groupi_n_163, csa_tree_add_6_33_groupi_n_164, csa_tree_add_6_33_groupi_n_165, csa_tree_add_6_33_groupi_n_166;
  wire csa_tree_add_6_33_groupi_n_167, csa_tree_add_6_33_groupi_n_168, csa_tree_add_6_33_groupi_n_169, csa_tree_add_6_33_groupi_n_170, csa_tree_add_6_33_groupi_n_171, csa_tree_add_6_33_groupi_n_172, csa_tree_add_6_33_groupi_n_173, csa_tree_add_6_33_groupi_n_174;
  wire csa_tree_add_6_33_groupi_n_175, csa_tree_add_6_33_groupi_n_176, csa_tree_add_6_33_groupi_n_177, csa_tree_add_6_33_groupi_n_178, csa_tree_add_6_33_groupi_n_179, csa_tree_add_6_33_groupi_n_180, csa_tree_add_6_33_groupi_n_181, csa_tree_add_6_33_groupi_n_182;
  wire csa_tree_add_6_33_groupi_n_183, csa_tree_add_6_33_groupi_n_184, csa_tree_add_6_33_groupi_n_185, csa_tree_add_6_33_groupi_n_186, csa_tree_add_6_33_groupi_n_187, csa_tree_add_6_33_groupi_n_188, csa_tree_add_6_33_groupi_n_189, csa_tree_add_6_33_groupi_n_190;
  wire csa_tree_add_6_33_groupi_n_191, csa_tree_add_6_33_groupi_n_192, csa_tree_add_6_33_groupi_n_193, csa_tree_add_6_33_groupi_n_194, csa_tree_add_6_33_groupi_n_195, csa_tree_add_6_33_groupi_n_196, csa_tree_add_6_33_groupi_n_197, csa_tree_add_6_33_groupi_n_198;
  wire csa_tree_add_6_33_groupi_n_199, csa_tree_add_6_33_groupi_n_200, csa_tree_add_6_33_groupi_n_201, csa_tree_add_6_33_groupi_n_202, csa_tree_add_6_33_groupi_n_203, csa_tree_add_6_33_groupi_n_204, csa_tree_add_6_33_groupi_n_205, csa_tree_add_6_33_groupi_n_206;
  wire csa_tree_add_6_33_groupi_n_207, csa_tree_add_6_33_groupi_n_208, csa_tree_add_6_33_groupi_n_209, csa_tree_add_6_33_groupi_n_210, csa_tree_add_6_33_groupi_n_211, csa_tree_add_6_33_groupi_n_212, csa_tree_add_6_33_groupi_n_213, csa_tree_add_6_33_groupi_n_214;
  wire csa_tree_add_6_33_groupi_n_215, csa_tree_add_6_33_groupi_n_216, csa_tree_add_6_33_groupi_n_217, csa_tree_add_6_33_groupi_n_218, csa_tree_add_6_33_groupi_n_219, csa_tree_add_6_33_groupi_n_220, csa_tree_add_6_33_groupi_n_221, csa_tree_add_6_33_groupi_n_222;
  wire csa_tree_add_6_33_groupi_n_223, csa_tree_add_6_33_groupi_n_224, csa_tree_add_6_33_groupi_n_225, csa_tree_add_6_33_groupi_n_226, csa_tree_add_6_33_groupi_n_227, csa_tree_add_6_33_groupi_n_228, csa_tree_add_6_33_groupi_n_229, csa_tree_add_6_33_groupi_n_230;
  wire csa_tree_add_6_33_groupi_n_231, csa_tree_add_6_33_groupi_n_232, csa_tree_add_6_33_groupi_n_233, csa_tree_add_6_33_groupi_n_234, csa_tree_add_6_33_groupi_n_235, csa_tree_add_6_33_groupi_n_236, csa_tree_add_6_33_groupi_n_237, csa_tree_add_6_33_groupi_n_238;
  wire csa_tree_add_6_33_groupi_n_239, csa_tree_add_6_33_groupi_n_240, csa_tree_add_6_33_groupi_n_241, csa_tree_add_6_33_groupi_n_242, csa_tree_add_6_33_groupi_n_243, csa_tree_add_6_33_groupi_n_244, csa_tree_add_6_33_groupi_n_245, csa_tree_add_6_33_groupi_n_246;
  wire csa_tree_add_6_33_groupi_n_247, csa_tree_add_6_33_groupi_n_248, csa_tree_add_6_33_groupi_n_249, csa_tree_add_6_33_groupi_n_250, csa_tree_add_6_33_groupi_n_251, csa_tree_add_6_33_groupi_n_252, csa_tree_add_6_33_groupi_n_253, csa_tree_add_6_33_groupi_n_254;
  wire csa_tree_add_6_33_groupi_n_255, csa_tree_add_6_33_groupi_n_256, csa_tree_add_6_33_groupi_n_257, csa_tree_add_6_33_groupi_n_258, csa_tree_add_6_33_groupi_n_259, csa_tree_add_6_33_groupi_n_260, csa_tree_add_6_33_groupi_n_261, csa_tree_add_6_33_groupi_n_262;
  wire csa_tree_add_6_33_groupi_n_263, csa_tree_add_6_33_groupi_n_264, csa_tree_add_6_33_groupi_n_265, csa_tree_add_6_33_groupi_n_266, csa_tree_add_6_33_groupi_n_267, csa_tree_add_6_33_groupi_n_268, csa_tree_add_6_33_groupi_n_269, csa_tree_add_6_33_groupi_n_270;
  wire csa_tree_add_6_33_groupi_n_271, csa_tree_add_6_33_groupi_n_272, csa_tree_add_6_33_groupi_n_273, csa_tree_add_6_33_groupi_n_274, csa_tree_add_6_33_groupi_n_275, csa_tree_add_6_33_groupi_n_276, csa_tree_add_6_33_groupi_n_277, csa_tree_add_6_33_groupi_n_278;
  wire csa_tree_add_6_33_groupi_n_279, csa_tree_add_6_33_groupi_n_280, csa_tree_add_6_33_groupi_n_281, csa_tree_add_6_33_groupi_n_282, csa_tree_add_6_33_groupi_n_283, csa_tree_add_6_33_groupi_n_284, csa_tree_add_6_33_groupi_n_285, csa_tree_add_6_33_groupi_n_286;
  wire csa_tree_add_6_33_groupi_n_287, csa_tree_add_6_33_groupi_n_288, csa_tree_add_6_33_groupi_n_289, csa_tree_add_6_33_groupi_n_290, csa_tree_add_6_33_groupi_n_291, csa_tree_add_6_33_groupi_n_292, csa_tree_add_6_33_groupi_n_293, csa_tree_add_6_33_groupi_n_294;
  wire csa_tree_add_6_33_groupi_n_295, csa_tree_add_6_33_groupi_n_296, csa_tree_add_6_33_groupi_n_297, csa_tree_add_6_33_groupi_n_298, csa_tree_add_6_33_groupi_n_299, csa_tree_add_6_33_groupi_n_300, csa_tree_add_6_33_groupi_n_301, csa_tree_add_6_33_groupi_n_302;
  wire csa_tree_add_6_33_groupi_n_303, csa_tree_add_6_33_groupi_n_304, csa_tree_add_6_33_groupi_n_305, csa_tree_add_6_33_groupi_n_306, csa_tree_add_6_33_groupi_n_307, csa_tree_add_6_33_groupi_n_308, csa_tree_add_6_33_groupi_n_309, csa_tree_add_6_33_groupi_n_310;
  wire csa_tree_add_6_33_groupi_n_311, csa_tree_add_6_33_groupi_n_312, csa_tree_add_6_33_groupi_n_313, csa_tree_add_6_33_groupi_n_314, csa_tree_add_6_33_groupi_n_315, csa_tree_add_6_33_groupi_n_316, csa_tree_add_6_33_groupi_n_317, csa_tree_add_6_33_groupi_n_318;
  wire csa_tree_add_6_33_groupi_n_319, csa_tree_add_6_33_groupi_n_320, csa_tree_add_6_33_groupi_n_321, csa_tree_add_6_33_groupi_n_322, csa_tree_add_6_33_groupi_n_323, csa_tree_add_6_33_groupi_n_324, csa_tree_add_6_33_groupi_n_325, csa_tree_add_6_33_groupi_n_326;
  wire csa_tree_add_6_33_groupi_n_327, csa_tree_add_6_33_groupi_n_328, csa_tree_add_6_33_groupi_n_329, csa_tree_add_6_33_groupi_n_330, csa_tree_add_6_33_groupi_n_331, csa_tree_add_6_33_groupi_n_332, csa_tree_add_6_33_groupi_n_333, csa_tree_add_6_33_groupi_n_334;
  wire csa_tree_add_6_33_groupi_n_335, csa_tree_add_6_33_groupi_n_336, csa_tree_add_6_33_groupi_n_337, csa_tree_add_6_33_groupi_n_338, csa_tree_add_6_33_groupi_n_339, csa_tree_add_6_33_groupi_n_340, csa_tree_add_6_33_groupi_n_341, csa_tree_add_6_33_groupi_n_342;
  wire csa_tree_add_6_33_groupi_n_343, csa_tree_add_6_33_groupi_n_344, csa_tree_add_6_33_groupi_n_345, csa_tree_add_6_33_groupi_n_346, csa_tree_add_6_33_groupi_n_347, csa_tree_add_6_33_groupi_n_348, csa_tree_add_6_33_groupi_n_349, csa_tree_add_6_33_groupi_n_350;
  wire csa_tree_add_6_33_groupi_n_351, csa_tree_add_6_33_groupi_n_352, csa_tree_add_6_33_groupi_n_353, csa_tree_add_6_33_groupi_n_354, csa_tree_add_6_33_groupi_n_355, csa_tree_add_6_33_groupi_n_356, csa_tree_add_6_33_groupi_n_357, csa_tree_add_6_33_groupi_n_358;
  wire csa_tree_add_6_33_groupi_n_359, csa_tree_add_6_33_groupi_n_360, csa_tree_add_6_33_groupi_n_361, csa_tree_add_6_33_groupi_n_362, csa_tree_add_6_33_groupi_n_363, csa_tree_add_6_33_groupi_n_364, csa_tree_add_6_33_groupi_n_365, csa_tree_add_6_33_groupi_n_366;
  wire csa_tree_add_6_33_groupi_n_367, csa_tree_add_6_33_groupi_n_368, csa_tree_add_6_33_groupi_n_369, csa_tree_add_6_33_groupi_n_370, csa_tree_add_6_33_groupi_n_371, csa_tree_add_6_33_groupi_n_372, csa_tree_add_6_33_groupi_n_373, csa_tree_add_6_33_groupi_n_374;
  wire csa_tree_add_6_33_groupi_n_375, csa_tree_add_6_33_groupi_n_376, csa_tree_add_6_33_groupi_n_377, csa_tree_add_6_33_groupi_n_378, csa_tree_add_6_33_groupi_n_379, csa_tree_add_6_33_groupi_n_380, csa_tree_add_6_33_groupi_n_381, csa_tree_add_6_33_groupi_n_382;
  wire csa_tree_add_6_33_groupi_n_383, csa_tree_add_6_33_groupi_n_384, csa_tree_add_6_33_groupi_n_385, csa_tree_add_6_33_groupi_n_386, csa_tree_add_6_33_groupi_n_387, csa_tree_add_6_33_groupi_n_388, csa_tree_add_6_33_groupi_n_389, csa_tree_add_6_33_groupi_n_390;
  wire csa_tree_add_6_33_groupi_n_391, csa_tree_add_6_33_groupi_n_392, csa_tree_add_6_33_groupi_n_393, csa_tree_add_6_33_groupi_n_394, csa_tree_add_6_33_groupi_n_395, csa_tree_add_6_33_groupi_n_396, csa_tree_add_6_33_groupi_n_397, csa_tree_add_6_33_groupi_n_398;
  wire csa_tree_add_6_33_groupi_n_399, csa_tree_add_6_33_groupi_n_400, csa_tree_add_6_33_groupi_n_401, csa_tree_add_6_33_groupi_n_402, csa_tree_add_6_33_groupi_n_403, csa_tree_add_6_33_groupi_n_404, csa_tree_add_6_33_groupi_n_405, csa_tree_add_6_33_groupi_n_406;
  wire csa_tree_add_6_33_groupi_n_407, csa_tree_add_6_33_groupi_n_408, csa_tree_add_6_33_groupi_n_409, csa_tree_add_6_33_groupi_n_410, csa_tree_add_6_33_groupi_n_411, csa_tree_add_6_33_groupi_n_412, csa_tree_add_6_33_groupi_n_413, csa_tree_add_6_33_groupi_n_414;
  wire csa_tree_add_6_33_groupi_n_415, csa_tree_add_6_33_groupi_n_416, csa_tree_add_6_33_groupi_n_417, csa_tree_add_6_33_groupi_n_418, csa_tree_add_6_33_groupi_n_419, csa_tree_add_6_33_groupi_n_420, csa_tree_add_6_33_groupi_n_421, csa_tree_add_6_33_groupi_n_422;
  wire csa_tree_add_6_33_groupi_n_423, csa_tree_add_6_33_groupi_n_424, csa_tree_add_6_33_groupi_n_425, csa_tree_add_6_33_groupi_n_426, csa_tree_add_6_33_groupi_n_427, csa_tree_add_6_33_groupi_n_428, csa_tree_add_6_33_groupi_n_429, csa_tree_add_6_33_groupi_n_430;
  wire csa_tree_add_6_33_groupi_n_431, csa_tree_add_6_33_groupi_n_432, csa_tree_add_6_33_groupi_n_433, csa_tree_add_6_33_groupi_n_434, csa_tree_add_6_33_groupi_n_435, csa_tree_add_6_33_groupi_n_436, csa_tree_add_6_33_groupi_n_437, csa_tree_add_6_33_groupi_n_438;
  wire csa_tree_add_6_33_groupi_n_439, csa_tree_add_6_33_groupi_n_440, csa_tree_add_6_33_groupi_n_441, csa_tree_add_6_33_groupi_n_442, csa_tree_add_6_33_groupi_n_443, csa_tree_add_6_33_groupi_n_444, csa_tree_add_6_33_groupi_n_445, csa_tree_add_6_33_groupi_n_446;
  wire csa_tree_add_6_33_groupi_n_447, csa_tree_add_6_33_groupi_n_448, csa_tree_add_6_33_groupi_n_449, csa_tree_add_6_33_groupi_n_450, csa_tree_add_6_33_groupi_n_451, csa_tree_add_6_33_groupi_n_452, csa_tree_add_6_33_groupi_n_453, csa_tree_add_6_33_groupi_n_454;
  wire csa_tree_add_6_33_groupi_n_455, csa_tree_add_6_33_groupi_n_456, csa_tree_add_6_33_groupi_n_457, csa_tree_add_6_33_groupi_n_458, csa_tree_add_6_33_groupi_n_459, csa_tree_add_6_33_groupi_n_460, csa_tree_add_6_33_groupi_n_461, csa_tree_add_6_33_groupi_n_462;
  wire csa_tree_add_6_33_groupi_n_463, csa_tree_add_6_33_groupi_n_464, csa_tree_add_6_33_groupi_n_465, csa_tree_add_6_33_groupi_n_466, csa_tree_add_6_33_groupi_n_467, csa_tree_add_6_33_groupi_n_468, csa_tree_add_6_33_groupi_n_469, csa_tree_add_6_33_groupi_n_470;
  wire csa_tree_add_6_33_groupi_n_471, csa_tree_add_6_33_groupi_n_472, csa_tree_add_6_33_groupi_n_473, csa_tree_add_6_33_groupi_n_474, csa_tree_add_6_33_groupi_n_475, csa_tree_add_6_33_groupi_n_476, csa_tree_add_6_33_groupi_n_477, csa_tree_add_6_33_groupi_n_478;
  wire csa_tree_add_6_33_groupi_n_479, csa_tree_add_6_33_groupi_n_480, csa_tree_add_6_33_groupi_n_481, csa_tree_add_6_33_groupi_n_482, csa_tree_add_6_33_groupi_n_483, csa_tree_add_6_33_groupi_n_484, csa_tree_add_6_33_groupi_n_485, csa_tree_add_6_33_groupi_n_486;
  wire csa_tree_add_6_33_groupi_n_487, csa_tree_add_6_33_groupi_n_488, csa_tree_add_6_33_groupi_n_489, csa_tree_add_6_33_groupi_n_490, csa_tree_add_6_33_groupi_n_491, csa_tree_add_6_33_groupi_n_492, csa_tree_add_6_33_groupi_n_493, csa_tree_add_6_33_groupi_n_494;
  wire csa_tree_add_6_33_groupi_n_495, csa_tree_add_6_33_groupi_n_496, csa_tree_add_6_33_groupi_n_497, csa_tree_add_6_33_groupi_n_498, csa_tree_add_6_33_groupi_n_499, csa_tree_add_6_33_groupi_n_500, csa_tree_add_6_33_groupi_n_501, csa_tree_add_6_33_groupi_n_502;
  wire csa_tree_add_6_33_groupi_n_503, csa_tree_add_6_33_groupi_n_504, csa_tree_add_6_33_groupi_n_505, csa_tree_add_6_33_groupi_n_506, csa_tree_add_6_33_groupi_n_507, csa_tree_add_6_33_groupi_n_508, csa_tree_add_6_33_groupi_n_509, csa_tree_add_6_33_groupi_n_510;
  wire csa_tree_add_6_33_groupi_n_511, csa_tree_add_6_33_groupi_n_512, csa_tree_add_6_33_groupi_n_513, csa_tree_add_6_33_groupi_n_514, csa_tree_add_6_33_groupi_n_515, csa_tree_add_6_33_groupi_n_516, csa_tree_add_6_33_groupi_n_517, csa_tree_add_6_33_groupi_n_518;
  wire csa_tree_add_6_33_groupi_n_519, csa_tree_add_6_33_groupi_n_520, csa_tree_add_6_33_groupi_n_521, csa_tree_add_6_33_groupi_n_522, csa_tree_add_6_33_groupi_n_523, csa_tree_add_6_33_groupi_n_524, csa_tree_add_6_33_groupi_n_525, csa_tree_add_6_33_groupi_n_526;
  wire csa_tree_add_6_33_groupi_n_527, csa_tree_add_6_33_groupi_n_528, csa_tree_add_6_33_groupi_n_529, csa_tree_add_6_33_groupi_n_530, csa_tree_add_6_33_groupi_n_531, csa_tree_add_6_33_groupi_n_532, csa_tree_add_6_33_groupi_n_533, csa_tree_add_6_33_groupi_n_534;
  wire csa_tree_add_6_33_groupi_n_535, csa_tree_add_6_33_groupi_n_536, csa_tree_add_6_33_groupi_n_537, csa_tree_add_6_33_groupi_n_538, csa_tree_add_6_33_groupi_n_539, csa_tree_add_6_33_groupi_n_540, csa_tree_add_6_33_groupi_n_541, csa_tree_add_6_33_groupi_n_542;
  wire csa_tree_add_6_33_groupi_n_543, csa_tree_add_6_33_groupi_n_544, csa_tree_add_6_33_groupi_n_545, csa_tree_add_6_33_groupi_n_546, csa_tree_add_6_33_groupi_n_547, csa_tree_add_6_33_groupi_n_548, csa_tree_add_6_33_groupi_n_549, csa_tree_add_6_33_groupi_n_550;
  wire csa_tree_add_6_33_groupi_n_551, csa_tree_add_6_33_groupi_n_552, csa_tree_add_6_33_groupi_n_553, csa_tree_add_6_33_groupi_n_554, csa_tree_add_6_33_groupi_n_555, csa_tree_add_6_33_groupi_n_556, csa_tree_add_6_33_groupi_n_557, csa_tree_add_6_33_groupi_n_558;
  wire csa_tree_add_6_33_groupi_n_559, csa_tree_add_6_33_groupi_n_560, csa_tree_add_6_33_groupi_n_561, csa_tree_add_6_33_groupi_n_562, csa_tree_add_6_33_groupi_n_563, csa_tree_add_6_33_groupi_n_564, csa_tree_add_6_33_groupi_n_565, csa_tree_add_6_33_groupi_n_566;
  wire csa_tree_add_6_33_groupi_n_567, csa_tree_add_6_33_groupi_n_568, csa_tree_add_6_33_groupi_n_569, csa_tree_add_6_33_groupi_n_570, csa_tree_add_6_33_groupi_n_571, csa_tree_add_6_33_groupi_n_572, csa_tree_add_6_33_groupi_n_573, csa_tree_add_6_33_groupi_n_574;
  wire csa_tree_add_6_33_groupi_n_575, csa_tree_add_6_33_groupi_n_576, csa_tree_add_6_33_groupi_n_577, csa_tree_add_6_33_groupi_n_578, csa_tree_add_6_33_groupi_n_579, csa_tree_add_6_33_groupi_n_580, csa_tree_add_6_33_groupi_n_581, csa_tree_add_6_33_groupi_n_582;
  wire csa_tree_add_6_33_groupi_n_583, csa_tree_add_6_33_groupi_n_584, csa_tree_add_6_33_groupi_n_585, csa_tree_add_6_33_groupi_n_586, csa_tree_add_6_33_groupi_n_587, csa_tree_add_6_33_groupi_n_588, csa_tree_add_6_33_groupi_n_589, csa_tree_add_6_33_groupi_n_590;
  wire csa_tree_add_6_33_groupi_n_591, csa_tree_add_6_33_groupi_n_592, csa_tree_add_6_33_groupi_n_593, csa_tree_add_6_33_groupi_n_594, csa_tree_add_6_33_groupi_n_595, csa_tree_add_6_33_groupi_n_596, csa_tree_add_6_33_groupi_n_597, csa_tree_add_6_33_groupi_n_598;
  wire csa_tree_add_6_33_groupi_n_599, csa_tree_add_6_33_groupi_n_600, csa_tree_add_6_33_groupi_n_601, csa_tree_add_6_33_groupi_n_602, csa_tree_add_6_33_groupi_n_603, csa_tree_add_6_33_groupi_n_604, csa_tree_add_6_33_groupi_n_605, csa_tree_add_6_33_groupi_n_606;
  wire csa_tree_add_6_33_groupi_n_607, csa_tree_add_6_33_groupi_n_608, csa_tree_add_6_33_groupi_n_609, csa_tree_add_6_33_groupi_n_610, csa_tree_add_6_33_groupi_n_611, csa_tree_add_6_33_groupi_n_612, csa_tree_add_6_33_groupi_n_613, csa_tree_add_6_33_groupi_n_614;
  wire csa_tree_add_6_33_groupi_n_615, csa_tree_add_6_33_groupi_n_616, csa_tree_add_6_33_groupi_n_617, csa_tree_add_6_33_groupi_n_618, csa_tree_add_6_33_groupi_n_619, csa_tree_add_6_33_groupi_n_620, csa_tree_add_6_33_groupi_n_621, csa_tree_add_6_33_groupi_n_622;
  wire csa_tree_add_6_33_groupi_n_623, csa_tree_add_6_33_groupi_n_624, csa_tree_add_6_33_groupi_n_625, csa_tree_add_6_33_groupi_n_626, csa_tree_add_6_33_groupi_n_627, csa_tree_add_6_33_groupi_n_628, csa_tree_add_6_33_groupi_n_629, csa_tree_add_6_33_groupi_n_630;
  wire csa_tree_add_6_33_groupi_n_631, csa_tree_add_6_33_groupi_n_632, csa_tree_add_6_33_groupi_n_633, csa_tree_add_6_33_groupi_n_634, csa_tree_add_6_33_groupi_n_635, csa_tree_add_6_33_groupi_n_636, csa_tree_add_6_33_groupi_n_637, csa_tree_add_6_33_groupi_n_638;
  wire csa_tree_add_6_33_groupi_n_639, csa_tree_add_6_33_groupi_n_640, csa_tree_add_6_33_groupi_n_641, csa_tree_add_6_33_groupi_n_642, csa_tree_add_6_33_groupi_n_643, csa_tree_add_6_33_groupi_n_644, csa_tree_add_6_33_groupi_n_645, csa_tree_add_6_33_groupi_n_646;
  wire csa_tree_add_6_33_groupi_n_647, csa_tree_add_6_33_groupi_n_648, csa_tree_add_6_33_groupi_n_649, csa_tree_add_6_33_groupi_n_650, csa_tree_add_6_33_groupi_n_651, csa_tree_add_6_33_groupi_n_652, csa_tree_add_6_33_groupi_n_653, csa_tree_add_6_33_groupi_n_654;
  wire csa_tree_add_6_33_groupi_n_655, csa_tree_add_6_33_groupi_n_656, csa_tree_add_6_33_groupi_n_657, csa_tree_add_6_33_groupi_n_658, csa_tree_add_6_33_groupi_n_659, csa_tree_add_6_33_groupi_n_660, csa_tree_add_6_33_groupi_n_661, csa_tree_add_6_33_groupi_n_662;
  wire csa_tree_add_6_33_groupi_n_663, csa_tree_add_6_33_groupi_n_664, csa_tree_add_6_33_groupi_n_665, csa_tree_add_6_33_groupi_n_666, csa_tree_add_6_33_groupi_n_667, csa_tree_add_6_33_groupi_n_668, csa_tree_add_6_33_groupi_n_669, csa_tree_add_6_33_groupi_n_670;
  wire csa_tree_add_6_33_groupi_n_671, csa_tree_add_6_33_groupi_n_672, csa_tree_add_6_33_groupi_n_673, csa_tree_add_6_33_groupi_n_674, csa_tree_add_6_33_groupi_n_675, csa_tree_add_6_33_groupi_n_676, csa_tree_add_6_33_groupi_n_677, csa_tree_add_6_33_groupi_n_678;
  wire csa_tree_add_6_33_groupi_n_679, csa_tree_add_6_33_groupi_n_680, csa_tree_add_6_33_groupi_n_681, csa_tree_add_6_33_groupi_n_682, csa_tree_add_6_33_groupi_n_683, csa_tree_add_6_33_groupi_n_684, csa_tree_add_6_33_groupi_n_685, csa_tree_add_6_33_groupi_n_686;
  wire csa_tree_add_6_33_groupi_n_687, csa_tree_add_6_33_groupi_n_688, csa_tree_add_6_33_groupi_n_689, csa_tree_add_6_33_groupi_n_690, csa_tree_add_6_33_groupi_n_691, csa_tree_add_6_33_groupi_n_692, csa_tree_add_6_33_groupi_n_693, csa_tree_add_6_33_groupi_n_694;
  wire csa_tree_add_6_33_groupi_n_695, csa_tree_add_6_33_groupi_n_696, csa_tree_add_6_33_groupi_n_697, csa_tree_add_6_33_groupi_n_698, csa_tree_add_6_33_groupi_n_699, csa_tree_add_6_33_groupi_n_700, csa_tree_add_6_33_groupi_n_701, csa_tree_add_6_33_groupi_n_702;
  wire csa_tree_add_6_33_groupi_n_703, csa_tree_add_6_33_groupi_n_704, csa_tree_add_6_33_groupi_n_705, csa_tree_add_6_33_groupi_n_706, csa_tree_add_6_33_groupi_n_707, csa_tree_add_6_33_groupi_n_708, csa_tree_add_6_33_groupi_n_709, csa_tree_add_6_33_groupi_n_710;
  wire csa_tree_add_6_33_groupi_n_711, csa_tree_add_6_33_groupi_n_712, csa_tree_add_6_33_groupi_n_713, csa_tree_add_6_33_groupi_n_714, csa_tree_add_6_33_groupi_n_715, csa_tree_add_6_33_groupi_n_716, csa_tree_add_6_33_groupi_n_717, csa_tree_add_6_33_groupi_n_718;
  wire csa_tree_add_6_33_groupi_n_719, csa_tree_add_6_33_groupi_n_720, csa_tree_add_6_33_groupi_n_721, csa_tree_add_6_33_groupi_n_722, csa_tree_add_6_33_groupi_n_723, csa_tree_add_6_33_groupi_n_724, csa_tree_add_6_33_groupi_n_725, csa_tree_add_6_33_groupi_n_726;
  wire csa_tree_add_6_33_groupi_n_727, csa_tree_add_6_33_groupi_n_728, csa_tree_add_6_33_groupi_n_729, csa_tree_add_6_33_groupi_n_730, csa_tree_add_6_33_groupi_n_731, csa_tree_add_6_33_groupi_n_732, csa_tree_add_6_33_groupi_n_733, csa_tree_add_6_33_groupi_n_734;
  wire csa_tree_add_6_33_groupi_n_735, csa_tree_add_6_33_groupi_n_736, csa_tree_add_6_33_groupi_n_737, csa_tree_add_6_33_groupi_n_738, csa_tree_add_6_33_groupi_n_739, csa_tree_add_6_33_groupi_n_740, csa_tree_add_6_33_groupi_n_741, csa_tree_add_6_33_groupi_n_742;
  wire csa_tree_add_6_33_groupi_n_743, csa_tree_add_6_33_groupi_n_744, csa_tree_add_6_33_groupi_n_745, csa_tree_add_6_33_groupi_n_746, csa_tree_add_6_33_groupi_n_747, csa_tree_add_6_33_groupi_n_748, csa_tree_add_6_33_groupi_n_749, csa_tree_add_6_33_groupi_n_750;
  wire csa_tree_add_6_33_groupi_n_751, csa_tree_add_6_33_groupi_n_752, csa_tree_add_6_33_groupi_n_753, csa_tree_add_6_33_groupi_n_754, csa_tree_add_6_33_groupi_n_755, csa_tree_add_6_33_groupi_n_756, csa_tree_add_6_33_groupi_n_757, csa_tree_add_6_33_groupi_n_758;
  wire csa_tree_add_6_33_groupi_n_759, csa_tree_add_6_33_groupi_n_760, csa_tree_add_6_33_groupi_n_761, csa_tree_add_6_33_groupi_n_762, csa_tree_add_6_33_groupi_n_763, csa_tree_add_6_33_groupi_n_764, csa_tree_add_6_33_groupi_n_765, csa_tree_add_6_33_groupi_n_766;
  wire csa_tree_add_6_33_groupi_n_767, csa_tree_add_6_33_groupi_n_768, csa_tree_add_6_33_groupi_n_769, csa_tree_add_6_33_groupi_n_770, csa_tree_add_6_33_groupi_n_771, csa_tree_add_6_33_groupi_n_772, csa_tree_add_6_33_groupi_n_773, csa_tree_add_6_33_groupi_n_774;
  wire csa_tree_add_6_33_groupi_n_775, csa_tree_add_6_33_groupi_n_776, csa_tree_add_6_33_groupi_n_777, csa_tree_add_6_33_groupi_n_778, csa_tree_add_6_33_groupi_n_779, csa_tree_add_6_33_groupi_n_780, csa_tree_add_6_33_groupi_n_781, csa_tree_add_6_33_groupi_n_782;
  wire csa_tree_add_6_33_groupi_n_783, csa_tree_add_6_33_groupi_n_784, csa_tree_add_6_33_groupi_n_785, csa_tree_add_6_33_groupi_n_786, csa_tree_add_6_33_groupi_n_787, csa_tree_add_6_33_groupi_n_788, csa_tree_add_6_33_groupi_n_789, csa_tree_add_6_33_groupi_n_790;
  wire csa_tree_add_6_33_groupi_n_791, csa_tree_add_6_33_groupi_n_792, csa_tree_add_6_33_groupi_n_793, csa_tree_add_6_33_groupi_n_794, csa_tree_add_6_33_groupi_n_795, csa_tree_add_6_33_groupi_n_796, csa_tree_add_6_33_groupi_n_797, csa_tree_add_6_33_groupi_n_798;
  wire csa_tree_add_6_33_groupi_n_799, csa_tree_add_6_33_groupi_n_800, csa_tree_add_6_33_groupi_n_801, csa_tree_add_6_33_groupi_n_802, csa_tree_add_6_33_groupi_n_803, csa_tree_add_6_33_groupi_n_804, csa_tree_add_6_33_groupi_n_805, csa_tree_add_6_33_groupi_n_806;
  wire csa_tree_add_6_33_groupi_n_807, csa_tree_add_6_33_groupi_n_808, csa_tree_add_6_33_groupi_n_809, csa_tree_add_6_33_groupi_n_810, csa_tree_add_6_33_groupi_n_811, csa_tree_add_6_33_groupi_n_812, csa_tree_add_6_33_groupi_n_813, csa_tree_add_6_33_groupi_n_814;
  wire csa_tree_add_6_33_groupi_n_815, csa_tree_add_6_33_groupi_n_816, csa_tree_add_6_33_groupi_n_817, csa_tree_add_6_33_groupi_n_818, csa_tree_add_6_33_groupi_n_819, csa_tree_add_6_33_groupi_n_820, csa_tree_add_6_33_groupi_n_821, csa_tree_add_6_33_groupi_n_822;
  wire csa_tree_add_6_33_groupi_n_823, csa_tree_add_6_33_groupi_n_824, csa_tree_add_6_33_groupi_n_825, csa_tree_add_6_33_groupi_n_826, csa_tree_add_6_33_groupi_n_827, csa_tree_add_6_33_groupi_n_828, csa_tree_add_6_33_groupi_n_829, csa_tree_add_6_33_groupi_n_830;
  wire csa_tree_add_6_33_groupi_n_831, csa_tree_add_6_33_groupi_n_832, csa_tree_add_6_33_groupi_n_833, csa_tree_add_6_33_groupi_n_834, csa_tree_add_6_33_groupi_n_835, csa_tree_add_6_33_groupi_n_836, csa_tree_add_6_33_groupi_n_837, csa_tree_add_6_33_groupi_n_838;
  wire csa_tree_add_6_33_groupi_n_839, csa_tree_add_6_33_groupi_n_840, csa_tree_add_6_33_groupi_n_841, csa_tree_add_6_33_groupi_n_842, csa_tree_add_6_33_groupi_n_843, csa_tree_add_6_33_groupi_n_844, csa_tree_add_6_33_groupi_n_845, csa_tree_add_6_33_groupi_n_846;
  wire csa_tree_add_6_33_groupi_n_847, csa_tree_add_6_33_groupi_n_848, csa_tree_add_6_33_groupi_n_849, csa_tree_add_6_33_groupi_n_850, csa_tree_add_6_33_groupi_n_851, csa_tree_add_6_33_groupi_n_852, csa_tree_add_6_33_groupi_n_853, csa_tree_add_6_33_groupi_n_854;
  wire csa_tree_add_6_33_groupi_n_855, csa_tree_add_6_33_groupi_n_856, csa_tree_add_6_33_groupi_n_857, csa_tree_add_6_33_groupi_n_858, csa_tree_add_6_33_groupi_n_859, csa_tree_add_6_33_groupi_n_860, csa_tree_add_6_33_groupi_n_861, csa_tree_add_6_33_groupi_n_862;
  wire csa_tree_add_6_33_groupi_n_863, csa_tree_add_6_33_groupi_n_864, csa_tree_add_6_33_groupi_n_865, csa_tree_add_6_33_groupi_n_866, csa_tree_add_6_33_groupi_n_867, csa_tree_add_6_33_groupi_n_868, csa_tree_add_6_33_groupi_n_869, csa_tree_add_6_33_groupi_n_870;
  wire csa_tree_add_6_33_groupi_n_871, csa_tree_add_6_33_groupi_n_872, csa_tree_add_6_33_groupi_n_873, csa_tree_add_6_33_groupi_n_874, csa_tree_add_6_33_groupi_n_875, csa_tree_add_6_33_groupi_n_876, csa_tree_add_6_33_groupi_n_877, csa_tree_add_6_33_groupi_n_878;
  wire csa_tree_add_6_33_groupi_n_879, csa_tree_add_6_33_groupi_n_880, csa_tree_add_6_33_groupi_n_881, csa_tree_add_6_33_groupi_n_882, csa_tree_add_6_33_groupi_n_883, csa_tree_add_6_33_groupi_n_884, csa_tree_add_6_33_groupi_n_885, csa_tree_add_6_33_groupi_n_886;
  wire csa_tree_add_6_33_groupi_n_887, csa_tree_add_6_33_groupi_n_888, csa_tree_add_6_33_groupi_n_889, csa_tree_add_6_33_groupi_n_890, csa_tree_add_6_33_groupi_n_891, csa_tree_add_6_33_groupi_n_892, csa_tree_add_6_33_groupi_n_893, csa_tree_add_6_33_groupi_n_894;
  wire csa_tree_add_6_33_groupi_n_895, csa_tree_add_6_33_groupi_n_896, csa_tree_add_6_33_groupi_n_897, csa_tree_add_6_33_groupi_n_898, csa_tree_add_6_33_groupi_n_899, csa_tree_add_6_33_groupi_n_900, csa_tree_add_6_33_groupi_n_901, csa_tree_add_6_33_groupi_n_902;
  wire csa_tree_add_6_33_groupi_n_903, csa_tree_add_6_33_groupi_n_904, csa_tree_add_6_33_groupi_n_905, csa_tree_add_6_33_groupi_n_906, csa_tree_add_6_33_groupi_n_907, csa_tree_add_6_33_groupi_n_908, csa_tree_add_6_33_groupi_n_909, csa_tree_add_6_33_groupi_n_910;
  wire csa_tree_add_6_33_groupi_n_911, csa_tree_add_6_33_groupi_n_912, csa_tree_add_6_33_groupi_n_913, csa_tree_add_6_33_groupi_n_914, csa_tree_add_6_33_groupi_n_915, csa_tree_add_6_33_groupi_n_916, csa_tree_add_6_33_groupi_n_917, csa_tree_add_6_33_groupi_n_918;
  wire csa_tree_add_6_33_groupi_n_919, csa_tree_add_6_33_groupi_n_920, csa_tree_add_6_33_groupi_n_921, csa_tree_add_6_33_groupi_n_922, csa_tree_add_6_33_groupi_n_923, csa_tree_add_6_33_groupi_n_924, csa_tree_add_6_33_groupi_n_925, csa_tree_add_6_33_groupi_n_926;
  wire csa_tree_add_6_33_groupi_n_927, csa_tree_add_6_33_groupi_n_928, csa_tree_add_6_33_groupi_n_929, csa_tree_add_6_33_groupi_n_930, csa_tree_add_6_33_groupi_n_931, csa_tree_add_6_33_groupi_n_932, csa_tree_add_6_33_groupi_n_933, csa_tree_add_6_33_groupi_n_934;
  wire csa_tree_add_6_33_groupi_n_935, csa_tree_add_6_33_groupi_n_936, csa_tree_add_6_33_groupi_n_937, csa_tree_add_6_33_groupi_n_938, csa_tree_add_6_33_groupi_n_939, csa_tree_add_6_33_groupi_n_940, csa_tree_add_6_33_groupi_n_941, csa_tree_add_6_33_groupi_n_942;
  wire csa_tree_add_6_33_groupi_n_943, csa_tree_add_6_33_groupi_n_944, csa_tree_add_6_33_groupi_n_945, csa_tree_add_6_33_groupi_n_946, csa_tree_add_6_33_groupi_n_947, csa_tree_add_6_33_groupi_n_948, csa_tree_add_6_33_groupi_n_949, csa_tree_add_6_33_groupi_n_950;
  wire csa_tree_add_6_33_groupi_n_951, csa_tree_add_6_33_groupi_n_952, csa_tree_add_6_33_groupi_n_953, csa_tree_add_6_33_groupi_n_954, csa_tree_add_6_33_groupi_n_955, csa_tree_add_6_33_groupi_n_956, csa_tree_add_6_33_groupi_n_957, csa_tree_add_6_33_groupi_n_958;
  wire csa_tree_add_6_33_groupi_n_959, csa_tree_add_6_33_groupi_n_960, csa_tree_add_6_33_groupi_n_961, csa_tree_add_6_33_groupi_n_962, csa_tree_add_6_33_groupi_n_963, csa_tree_add_6_33_groupi_n_964, csa_tree_add_6_33_groupi_n_965, csa_tree_add_6_33_groupi_n_966;
  wire csa_tree_add_6_33_groupi_n_967, csa_tree_add_6_33_groupi_n_968, csa_tree_add_6_33_groupi_n_969, csa_tree_add_6_33_groupi_n_970, csa_tree_add_6_33_groupi_n_971, csa_tree_add_6_33_groupi_n_972, csa_tree_add_6_33_groupi_n_973, csa_tree_add_6_33_groupi_n_974;
  wire csa_tree_add_6_33_groupi_n_975, csa_tree_add_6_33_groupi_n_976, csa_tree_add_6_33_groupi_n_977, csa_tree_add_6_33_groupi_n_978, csa_tree_add_6_33_groupi_n_979, csa_tree_add_6_33_groupi_n_980, csa_tree_add_6_33_groupi_n_981, csa_tree_add_6_33_groupi_n_982;
  wire csa_tree_add_6_33_groupi_n_983, csa_tree_add_6_33_groupi_n_984, csa_tree_add_6_33_groupi_n_985, csa_tree_add_6_33_groupi_n_986, csa_tree_add_6_33_groupi_n_987, csa_tree_add_6_33_groupi_n_988, csa_tree_add_6_33_groupi_n_989, csa_tree_add_6_33_groupi_n_990;
  wire csa_tree_add_6_33_groupi_n_991, csa_tree_add_6_33_groupi_n_992, csa_tree_add_6_33_groupi_n_993, csa_tree_add_6_33_groupi_n_994, csa_tree_add_6_33_groupi_n_995, csa_tree_add_6_33_groupi_n_996, csa_tree_add_6_33_groupi_n_997, csa_tree_add_6_33_groupi_n_998;
  wire csa_tree_add_6_33_groupi_n_999, csa_tree_add_6_33_groupi_n_1000, csa_tree_add_6_33_groupi_n_1001, csa_tree_add_6_33_groupi_n_1002, csa_tree_add_6_33_groupi_n_1003, csa_tree_add_6_33_groupi_n_1004, csa_tree_add_6_33_groupi_n_1005, csa_tree_add_6_33_groupi_n_1006;
  wire csa_tree_add_6_33_groupi_n_1007, csa_tree_add_6_33_groupi_n_1008, csa_tree_add_6_33_groupi_n_1009, csa_tree_add_6_33_groupi_n_1010, csa_tree_add_6_33_groupi_n_1011, csa_tree_add_6_33_groupi_n_1012, csa_tree_add_6_33_groupi_n_1013, csa_tree_add_6_33_groupi_n_1014;
  wire csa_tree_add_6_33_groupi_n_1015, csa_tree_add_6_33_groupi_n_1016, csa_tree_add_6_33_groupi_n_1017, csa_tree_add_6_33_groupi_n_1018, csa_tree_add_6_33_groupi_n_1019, csa_tree_add_6_33_groupi_n_1020, csa_tree_add_6_33_groupi_n_1021, csa_tree_add_6_33_groupi_n_1022;
  wire csa_tree_add_6_33_groupi_n_1023, csa_tree_add_6_33_groupi_n_1024, csa_tree_add_6_33_groupi_n_1025, csa_tree_add_6_33_groupi_n_1026, csa_tree_add_6_33_groupi_n_1027, csa_tree_add_6_33_groupi_n_1028, csa_tree_add_6_33_groupi_n_1029, csa_tree_add_6_33_groupi_n_1030;
  wire csa_tree_add_6_33_groupi_n_1031, csa_tree_add_6_33_groupi_n_1032, csa_tree_add_6_33_groupi_n_1033, csa_tree_add_6_33_groupi_n_1034, csa_tree_add_6_33_groupi_n_1035, csa_tree_add_6_33_groupi_n_1036, csa_tree_add_6_33_groupi_n_1037, csa_tree_add_6_33_groupi_n_1038;
  wire csa_tree_add_6_33_groupi_n_1039, csa_tree_add_6_33_groupi_n_1040, csa_tree_add_6_33_groupi_n_1041, csa_tree_add_6_33_groupi_n_1042, csa_tree_add_6_33_groupi_n_1043, csa_tree_add_6_33_groupi_n_1044, csa_tree_add_6_33_groupi_n_1045, csa_tree_add_6_33_groupi_n_1046;
  wire csa_tree_add_6_33_groupi_n_1047, csa_tree_add_6_33_groupi_n_1048, csa_tree_add_6_33_groupi_n_1049, csa_tree_add_6_33_groupi_n_1050, csa_tree_add_6_33_groupi_n_1051, csa_tree_add_6_33_groupi_n_1052, csa_tree_add_6_33_groupi_n_1053, csa_tree_add_6_33_groupi_n_1054;
  wire csa_tree_add_6_33_groupi_n_1055, csa_tree_add_6_33_groupi_n_1056, csa_tree_add_6_33_groupi_n_1057, csa_tree_add_6_33_groupi_n_1058, csa_tree_add_6_33_groupi_n_1059, csa_tree_add_6_33_groupi_n_1060, csa_tree_add_6_33_groupi_n_1061, csa_tree_add_6_33_groupi_n_1062;
  wire csa_tree_add_6_33_groupi_n_1063, csa_tree_add_6_33_groupi_n_1064, csa_tree_add_6_33_groupi_n_1065, csa_tree_add_6_33_groupi_n_1066, csa_tree_add_6_33_groupi_n_1067, csa_tree_add_6_33_groupi_n_1068, csa_tree_add_6_33_groupi_n_1069, csa_tree_add_6_33_groupi_n_1070;
  wire csa_tree_add_6_33_groupi_n_1071, csa_tree_add_6_33_groupi_n_1072, csa_tree_add_6_33_groupi_n_1073, csa_tree_add_6_33_groupi_n_1074, csa_tree_add_6_33_groupi_n_1075, csa_tree_add_6_33_groupi_n_1076, csa_tree_add_6_33_groupi_n_1077, csa_tree_add_6_33_groupi_n_1078;
  wire csa_tree_add_6_33_groupi_n_1079, csa_tree_add_6_33_groupi_n_1080, csa_tree_add_6_33_groupi_n_1081, csa_tree_add_6_33_groupi_n_1082, csa_tree_add_6_33_groupi_n_1083, csa_tree_add_6_33_groupi_n_1084, csa_tree_add_6_33_groupi_n_1085, csa_tree_add_6_33_groupi_n_1086;
  wire csa_tree_add_6_33_groupi_n_1087, csa_tree_add_6_33_groupi_n_1088, csa_tree_add_6_33_groupi_n_1089, csa_tree_add_6_33_groupi_n_1090, csa_tree_add_6_33_groupi_n_1091, csa_tree_add_6_33_groupi_n_1092, csa_tree_add_6_33_groupi_n_1093, csa_tree_add_6_33_groupi_n_1094;
  wire csa_tree_add_6_33_groupi_n_1095, csa_tree_add_6_33_groupi_n_1096, csa_tree_add_6_33_groupi_n_1097, csa_tree_add_6_33_groupi_n_1098, csa_tree_add_6_33_groupi_n_1099, csa_tree_add_6_33_groupi_n_1100, csa_tree_add_6_33_groupi_n_1101, csa_tree_add_6_33_groupi_n_1102;
  wire csa_tree_add_6_33_groupi_n_1103, csa_tree_add_6_33_groupi_n_1104, csa_tree_add_6_33_groupi_n_1105, csa_tree_add_6_33_groupi_n_1106, csa_tree_add_6_33_groupi_n_1107, csa_tree_add_6_33_groupi_n_1108, csa_tree_add_6_33_groupi_n_1109, csa_tree_add_6_33_groupi_n_1110;
  wire csa_tree_add_6_33_groupi_n_1111, csa_tree_add_6_33_groupi_n_1112, csa_tree_add_6_33_groupi_n_1113, csa_tree_add_6_33_groupi_n_1114, csa_tree_add_6_33_groupi_n_1115, csa_tree_add_6_33_groupi_n_1116, csa_tree_add_6_33_groupi_n_1117, csa_tree_add_6_33_groupi_n_1118;
  wire csa_tree_add_6_33_groupi_n_1119, csa_tree_add_6_33_groupi_n_1120, csa_tree_add_6_33_groupi_n_1121, csa_tree_add_6_33_groupi_n_1122, csa_tree_add_6_33_groupi_n_1123, csa_tree_add_6_33_groupi_n_1124, csa_tree_add_6_33_groupi_n_1125, csa_tree_add_6_33_groupi_n_1126;
  wire csa_tree_add_6_33_groupi_n_1127, csa_tree_add_6_33_groupi_n_1128, csa_tree_add_6_33_groupi_n_1129, csa_tree_add_6_33_groupi_n_1130, csa_tree_add_6_33_groupi_n_1131, csa_tree_add_6_33_groupi_n_1132, csa_tree_add_6_33_groupi_n_1133, csa_tree_add_6_33_groupi_n_1134;
  wire csa_tree_add_6_33_groupi_n_1135, csa_tree_add_6_33_groupi_n_1136, csa_tree_add_6_33_groupi_n_1137, csa_tree_add_6_33_groupi_n_1138, csa_tree_add_6_33_groupi_n_1139, csa_tree_add_6_33_groupi_n_1140, csa_tree_add_6_33_groupi_n_1141, csa_tree_add_6_33_groupi_n_1142;
  wire csa_tree_add_6_33_groupi_n_1143, csa_tree_add_6_33_groupi_n_1144, csa_tree_add_6_33_groupi_n_1145, csa_tree_add_6_33_groupi_n_1146, csa_tree_add_6_33_groupi_n_1147, csa_tree_add_6_33_groupi_n_1148, csa_tree_add_6_33_groupi_n_1149, csa_tree_add_6_33_groupi_n_1150;
  wire csa_tree_add_6_33_groupi_n_1151, csa_tree_add_6_33_groupi_n_1152, csa_tree_add_6_33_groupi_n_1153, csa_tree_add_6_33_groupi_n_1154, csa_tree_add_6_33_groupi_n_1155, csa_tree_add_6_33_groupi_n_1156, csa_tree_add_6_33_groupi_n_1157, csa_tree_add_6_33_groupi_n_1158;
  wire csa_tree_add_6_33_groupi_n_1159, csa_tree_add_6_33_groupi_n_1160, csa_tree_add_6_33_groupi_n_1161, csa_tree_add_6_33_groupi_n_1162, csa_tree_add_6_33_groupi_n_1163, csa_tree_add_6_33_groupi_n_1164, csa_tree_add_6_33_groupi_n_1165, csa_tree_add_6_33_groupi_n_1166;
  wire csa_tree_add_6_33_groupi_n_1167, csa_tree_add_6_33_groupi_n_1168, csa_tree_add_6_33_groupi_n_1169, csa_tree_add_6_33_groupi_n_1170, csa_tree_add_6_33_groupi_n_1171, csa_tree_add_6_33_groupi_n_1172, csa_tree_add_6_33_groupi_n_1173, csa_tree_add_6_33_groupi_n_1174;
  wire csa_tree_add_6_33_groupi_n_1175, csa_tree_add_6_33_groupi_n_1176, csa_tree_add_6_33_groupi_n_1177, csa_tree_add_6_33_groupi_n_1178, csa_tree_add_6_33_groupi_n_1179, csa_tree_add_6_33_groupi_n_1180, csa_tree_add_6_33_groupi_n_1181, csa_tree_add_6_33_groupi_n_1182;
  wire csa_tree_add_6_33_groupi_n_1183, csa_tree_add_6_33_groupi_n_1184, csa_tree_add_6_33_groupi_n_1185, csa_tree_add_6_33_groupi_n_1186, csa_tree_add_6_33_groupi_n_1187, csa_tree_add_6_33_groupi_n_1188, csa_tree_add_6_33_groupi_n_1189, csa_tree_add_6_33_groupi_n_1190;
  wire csa_tree_add_6_33_groupi_n_1191, csa_tree_add_6_33_groupi_n_1192, csa_tree_add_6_33_groupi_n_1193, csa_tree_add_6_33_groupi_n_1194, csa_tree_add_6_33_groupi_n_1195, csa_tree_add_6_33_groupi_n_1196, csa_tree_add_6_33_groupi_n_1197, csa_tree_add_6_33_groupi_n_1198;
  wire csa_tree_add_6_33_groupi_n_1199, csa_tree_add_6_33_groupi_n_1200, csa_tree_add_6_33_groupi_n_1201, csa_tree_add_6_33_groupi_n_1202, csa_tree_add_6_33_groupi_n_1203, csa_tree_add_6_33_groupi_n_1204, csa_tree_add_6_33_groupi_n_1205, csa_tree_add_6_33_groupi_n_1206;
  wire csa_tree_add_6_33_groupi_n_1207, csa_tree_add_6_33_groupi_n_1208, csa_tree_add_6_33_groupi_n_1209, csa_tree_add_6_33_groupi_n_1210, csa_tree_add_6_33_groupi_n_1211, csa_tree_add_6_33_groupi_n_1212, csa_tree_add_6_33_groupi_n_1213, csa_tree_add_6_33_groupi_n_1214;
  wire csa_tree_add_6_33_groupi_n_1215, csa_tree_add_6_33_groupi_n_1216, csa_tree_add_6_33_groupi_n_1217, csa_tree_add_6_33_groupi_n_1218, csa_tree_add_6_33_groupi_n_1219, csa_tree_add_6_33_groupi_n_1220, csa_tree_add_6_33_groupi_n_1221, csa_tree_add_6_33_groupi_n_1222;
  wire csa_tree_add_6_33_groupi_n_1223, csa_tree_add_6_33_groupi_n_1224, csa_tree_add_6_33_groupi_n_1225, csa_tree_add_6_33_groupi_n_1226, csa_tree_add_6_33_groupi_n_1227, csa_tree_add_6_33_groupi_n_1228, csa_tree_add_6_33_groupi_n_1229, csa_tree_add_6_33_groupi_n_1230;
  wire csa_tree_add_6_33_groupi_n_1231, csa_tree_add_6_33_groupi_n_1232, csa_tree_add_6_33_groupi_n_1233, csa_tree_add_6_33_groupi_n_1234, csa_tree_add_6_33_groupi_n_1235, csa_tree_add_6_33_groupi_n_1236, csa_tree_add_6_33_groupi_n_1237, csa_tree_add_6_33_groupi_n_1238;
  wire csa_tree_add_6_33_groupi_n_1239, csa_tree_add_6_33_groupi_n_1240, csa_tree_add_6_33_groupi_n_1241, csa_tree_add_6_33_groupi_n_1242, csa_tree_add_6_33_groupi_n_1243, csa_tree_add_6_33_groupi_n_1244, csa_tree_add_6_33_groupi_n_1245, csa_tree_add_6_33_groupi_n_1246;
  wire csa_tree_add_6_33_groupi_n_1247, csa_tree_add_6_33_groupi_n_1248, csa_tree_add_6_33_groupi_n_1249, csa_tree_add_6_33_groupi_n_1250, csa_tree_add_6_33_groupi_n_1251, csa_tree_add_6_33_groupi_n_1252, csa_tree_add_6_33_groupi_n_1253, csa_tree_add_6_33_groupi_n_1254;
  wire csa_tree_add_6_33_groupi_n_1255, csa_tree_add_6_33_groupi_n_1256, csa_tree_add_6_33_groupi_n_1257, csa_tree_add_6_33_groupi_n_1258, csa_tree_add_6_33_groupi_n_1259, csa_tree_add_6_33_groupi_n_1260, csa_tree_add_6_33_groupi_n_1261, csa_tree_add_6_33_groupi_n_1262;
  wire csa_tree_add_6_33_groupi_n_1263, csa_tree_add_6_33_groupi_n_1264, csa_tree_add_6_33_groupi_n_1265, csa_tree_add_6_33_groupi_n_1266, csa_tree_add_6_33_groupi_n_1267, csa_tree_add_6_33_groupi_n_1268, csa_tree_add_6_33_groupi_n_1269, csa_tree_add_6_33_groupi_n_1270;
  wire csa_tree_add_6_33_groupi_n_1271, csa_tree_add_6_33_groupi_n_1272, csa_tree_add_6_33_groupi_n_1273, csa_tree_add_6_33_groupi_n_1274, csa_tree_add_6_33_groupi_n_1275, csa_tree_add_6_33_groupi_n_1276, csa_tree_add_6_33_groupi_n_1277, csa_tree_add_6_33_groupi_n_1278;
  wire csa_tree_add_6_33_groupi_n_1279, csa_tree_add_6_33_groupi_n_1280, csa_tree_add_6_33_groupi_n_1281, csa_tree_add_6_33_groupi_n_1282, csa_tree_add_6_33_groupi_n_1283, csa_tree_add_6_33_groupi_n_1284, csa_tree_add_6_33_groupi_n_1285, csa_tree_add_6_33_groupi_n_1286;
  wire csa_tree_add_6_33_groupi_n_1287, csa_tree_add_6_33_groupi_n_1288, csa_tree_add_6_33_groupi_n_1289, csa_tree_add_6_33_groupi_n_1290, csa_tree_add_6_33_groupi_n_1291, csa_tree_add_6_33_groupi_n_1292, csa_tree_add_6_33_groupi_n_1293, csa_tree_add_6_33_groupi_n_1294;
  wire csa_tree_add_6_33_groupi_n_1295, csa_tree_add_6_33_groupi_n_1296, csa_tree_add_6_33_groupi_n_1297, csa_tree_add_6_33_groupi_n_1298, csa_tree_add_6_33_groupi_n_1299, csa_tree_add_6_33_groupi_n_1300, csa_tree_add_6_33_groupi_n_1301, csa_tree_add_6_33_groupi_n_1302;
  wire csa_tree_add_6_33_groupi_n_1303, csa_tree_add_6_33_groupi_n_1304, csa_tree_add_6_33_groupi_n_1305, csa_tree_add_6_33_groupi_n_1306, csa_tree_add_6_33_groupi_n_1307, csa_tree_add_6_33_groupi_n_1308, csa_tree_add_6_33_groupi_n_1309, csa_tree_add_6_33_groupi_n_1310;
  wire csa_tree_add_6_33_groupi_n_1311, csa_tree_add_6_33_groupi_n_1312, csa_tree_add_6_33_groupi_n_1313, csa_tree_add_6_33_groupi_n_1314, csa_tree_add_6_33_groupi_n_1315, csa_tree_add_6_33_groupi_n_1316, csa_tree_add_6_33_groupi_n_1317, csa_tree_add_6_33_groupi_n_1318;
  wire csa_tree_add_6_33_groupi_n_1319, csa_tree_add_6_33_groupi_n_1320, csa_tree_add_6_33_groupi_n_1321, csa_tree_add_6_33_groupi_n_1322, csa_tree_add_6_33_groupi_n_1323, csa_tree_add_6_33_groupi_n_1324, csa_tree_add_6_33_groupi_n_1325, csa_tree_add_6_33_groupi_n_1326;
  wire csa_tree_add_6_33_groupi_n_1327, csa_tree_add_6_33_groupi_n_1328, csa_tree_add_6_33_groupi_n_1329, csa_tree_add_6_33_groupi_n_1330, csa_tree_add_6_33_groupi_n_1331, csa_tree_add_6_33_groupi_n_1332, csa_tree_add_6_33_groupi_n_1333, csa_tree_add_6_33_groupi_n_1334;
  wire csa_tree_add_6_33_groupi_n_1335, csa_tree_add_6_33_groupi_n_1336, csa_tree_add_6_33_groupi_n_1337, csa_tree_add_6_33_groupi_n_1338, csa_tree_add_6_33_groupi_n_1339, csa_tree_add_6_33_groupi_n_1340, csa_tree_add_6_33_groupi_n_1341, csa_tree_add_6_33_groupi_n_1342;
  wire csa_tree_add_6_33_groupi_n_1343, csa_tree_add_6_33_groupi_n_1344, csa_tree_add_6_33_groupi_n_1345, csa_tree_add_6_33_groupi_n_1346, csa_tree_add_6_33_groupi_n_1347, csa_tree_add_6_33_groupi_n_1348, csa_tree_add_6_33_groupi_n_1349, csa_tree_add_6_33_groupi_n_1350;
  wire csa_tree_add_6_33_groupi_n_1351, csa_tree_add_6_33_groupi_n_1352, csa_tree_add_6_33_groupi_n_1353, csa_tree_add_6_33_groupi_n_1354, csa_tree_add_6_33_groupi_n_1355, csa_tree_add_6_33_groupi_n_1356, csa_tree_add_6_33_groupi_n_1357, csa_tree_add_6_33_groupi_n_1358;
  wire csa_tree_add_6_33_groupi_n_1359, csa_tree_add_6_33_groupi_n_1360, csa_tree_add_6_33_groupi_n_1361, csa_tree_add_6_33_groupi_n_1362, csa_tree_add_6_33_groupi_n_1363, csa_tree_add_6_33_groupi_n_1364, csa_tree_add_6_33_groupi_n_1365, csa_tree_add_6_33_groupi_n_1366;
  wire csa_tree_add_6_33_groupi_n_1367, csa_tree_add_6_33_groupi_n_1368, csa_tree_add_6_33_groupi_n_1369, csa_tree_add_6_33_groupi_n_1370, csa_tree_add_6_33_groupi_n_1371, csa_tree_add_6_33_groupi_n_1372, csa_tree_add_6_33_groupi_n_1373, csa_tree_add_6_33_groupi_n_1374;
  wire csa_tree_add_6_33_groupi_n_1375, csa_tree_add_6_33_groupi_n_1376, csa_tree_add_6_33_groupi_n_1377, csa_tree_add_6_33_groupi_n_1378, csa_tree_add_6_33_groupi_n_1379, csa_tree_add_6_33_groupi_n_1380, csa_tree_add_6_33_groupi_n_1381, csa_tree_add_6_33_groupi_n_1382;
  wire csa_tree_add_6_33_groupi_n_1383, csa_tree_add_6_33_groupi_n_1384, csa_tree_add_6_33_groupi_n_1385, csa_tree_add_6_33_groupi_n_1386, csa_tree_add_6_33_groupi_n_1387, csa_tree_add_6_33_groupi_n_1388, csa_tree_add_6_33_groupi_n_1389, csa_tree_add_6_33_groupi_n_1390;
  wire csa_tree_add_6_33_groupi_n_1391, csa_tree_add_6_33_groupi_n_1392, csa_tree_add_6_33_groupi_n_1393, csa_tree_add_6_33_groupi_n_1394, csa_tree_add_6_33_groupi_n_1395, csa_tree_add_6_33_groupi_n_1396, csa_tree_add_6_33_groupi_n_1397, csa_tree_add_6_33_groupi_n_1398;
  wire csa_tree_add_6_33_groupi_n_1399, csa_tree_add_6_33_groupi_n_1400, csa_tree_add_6_33_groupi_n_1401, csa_tree_add_6_33_groupi_n_1402, csa_tree_add_6_33_groupi_n_1403, csa_tree_add_6_33_groupi_n_1404, csa_tree_add_6_33_groupi_n_1405, csa_tree_add_6_33_groupi_n_1406;
  wire csa_tree_add_6_33_groupi_n_1407, csa_tree_add_6_33_groupi_n_1408, csa_tree_add_6_33_groupi_n_1409, csa_tree_add_6_33_groupi_n_1410, csa_tree_add_6_33_groupi_n_1411, csa_tree_add_6_33_groupi_n_1412, csa_tree_add_6_33_groupi_n_1413, csa_tree_add_6_33_groupi_n_1414;
  wire csa_tree_add_6_33_groupi_n_1415, csa_tree_add_6_33_groupi_n_1416, csa_tree_add_6_33_groupi_n_1417, csa_tree_add_6_33_groupi_n_1418, csa_tree_add_6_33_groupi_n_1419, csa_tree_add_6_33_groupi_n_1420, csa_tree_add_6_33_groupi_n_1421, csa_tree_add_6_33_groupi_n_1422;
  wire csa_tree_add_6_33_groupi_n_1423, csa_tree_add_6_33_groupi_n_1424, csa_tree_add_6_33_groupi_n_1425, csa_tree_add_6_33_groupi_n_1426, csa_tree_add_6_33_groupi_n_1427, csa_tree_add_6_33_groupi_n_1428, csa_tree_add_6_33_groupi_n_1429, csa_tree_add_6_33_groupi_n_1430;
  wire csa_tree_add_6_33_groupi_n_1431, csa_tree_add_6_33_groupi_n_1432, csa_tree_add_6_33_groupi_n_1433, csa_tree_add_6_33_groupi_n_1434, csa_tree_add_6_33_groupi_n_1435, csa_tree_add_6_33_groupi_n_1436, csa_tree_add_6_33_groupi_n_1437, csa_tree_add_6_33_groupi_n_1438;
  wire csa_tree_add_6_33_groupi_n_1439, csa_tree_add_6_33_groupi_n_1440, csa_tree_add_6_33_groupi_n_1441, csa_tree_add_6_33_groupi_n_1442, csa_tree_add_6_33_groupi_n_1443, csa_tree_add_6_33_groupi_n_1444, csa_tree_add_6_33_groupi_n_1445, csa_tree_add_6_33_groupi_n_1446;
  wire csa_tree_add_6_33_groupi_n_1447, csa_tree_add_6_33_groupi_n_1448, csa_tree_add_6_33_groupi_n_1449, csa_tree_add_6_33_groupi_n_1450, csa_tree_add_6_33_groupi_n_1451, csa_tree_add_6_33_groupi_n_1452, csa_tree_add_6_33_groupi_n_1453, csa_tree_add_6_33_groupi_n_1454;
  wire csa_tree_add_6_33_groupi_n_1455, csa_tree_add_6_33_groupi_n_1456, csa_tree_add_6_33_groupi_n_1457, csa_tree_add_6_33_groupi_n_1458, csa_tree_add_6_33_groupi_n_1459, csa_tree_add_6_33_groupi_n_1460, csa_tree_add_6_33_groupi_n_1461, csa_tree_add_6_33_groupi_n_1462;
  wire csa_tree_add_6_33_groupi_n_1463, csa_tree_add_6_33_groupi_n_1464, csa_tree_add_6_33_groupi_n_1465, csa_tree_add_6_33_groupi_n_1466, csa_tree_add_6_33_groupi_n_1467, csa_tree_add_6_33_groupi_n_1468, csa_tree_add_6_33_groupi_n_1469, csa_tree_add_6_33_groupi_n_1470;
  wire csa_tree_add_6_33_groupi_n_1471, csa_tree_add_6_33_groupi_n_1472, csa_tree_add_6_33_groupi_n_1473, csa_tree_add_6_33_groupi_n_1474, csa_tree_add_6_33_groupi_n_1475, csa_tree_add_6_33_groupi_n_1476, csa_tree_add_6_33_groupi_n_1477, csa_tree_add_6_33_groupi_n_1478;
  wire csa_tree_add_6_33_groupi_n_1479, csa_tree_add_6_33_groupi_n_1480, csa_tree_add_6_33_groupi_n_1481, csa_tree_add_6_33_groupi_n_1482, csa_tree_add_6_33_groupi_n_1483, csa_tree_add_6_33_groupi_n_1484, csa_tree_add_6_33_groupi_n_1485, csa_tree_add_6_33_groupi_n_1486;
  wire csa_tree_add_6_33_groupi_n_1487, csa_tree_add_6_33_groupi_n_1488, csa_tree_add_6_33_groupi_n_1489, csa_tree_add_6_33_groupi_n_1490, csa_tree_add_6_33_groupi_n_1491, csa_tree_add_6_33_groupi_n_1492, csa_tree_add_6_33_groupi_n_1493, csa_tree_add_6_33_groupi_n_1494;
  wire csa_tree_add_6_33_groupi_n_1495, csa_tree_add_6_33_groupi_n_1496, csa_tree_add_6_33_groupi_n_1497, csa_tree_add_6_33_groupi_n_1498, csa_tree_add_6_33_groupi_n_1499, csa_tree_add_6_33_groupi_n_1500, csa_tree_add_6_33_groupi_n_1501, csa_tree_add_6_33_groupi_n_1502;
  wire csa_tree_add_6_33_groupi_n_1503, csa_tree_add_6_33_groupi_n_1504, csa_tree_add_6_33_groupi_n_1505, csa_tree_add_6_33_groupi_n_1506, csa_tree_add_6_33_groupi_n_1507, csa_tree_add_6_33_groupi_n_1508, csa_tree_add_6_33_groupi_n_1509, csa_tree_add_6_33_groupi_n_1510;
  wire csa_tree_add_6_33_groupi_n_1511, csa_tree_add_6_33_groupi_n_1512, csa_tree_add_6_33_groupi_n_1513, csa_tree_add_6_33_groupi_n_1514, csa_tree_add_6_33_groupi_n_1515, csa_tree_add_6_33_groupi_n_1516, csa_tree_add_6_33_groupi_n_1517, csa_tree_add_6_33_groupi_n_1518;
  wire csa_tree_add_6_33_groupi_n_1519, csa_tree_add_6_33_groupi_n_1520, csa_tree_add_6_33_groupi_n_1521, csa_tree_add_6_33_groupi_n_1522, csa_tree_add_6_33_groupi_n_1523, csa_tree_add_6_33_groupi_n_1524, csa_tree_add_6_33_groupi_n_1525, csa_tree_add_6_33_groupi_n_1526;
  wire csa_tree_add_6_33_groupi_n_1527, csa_tree_add_6_33_groupi_n_1528, csa_tree_add_6_33_groupi_n_1529, csa_tree_add_6_33_groupi_n_1530, csa_tree_add_6_33_groupi_n_1531, csa_tree_add_6_33_groupi_n_1532, csa_tree_add_6_33_groupi_n_1533, csa_tree_add_6_33_groupi_n_1534;
  wire csa_tree_add_6_33_groupi_n_1535, csa_tree_add_6_33_groupi_n_1536, csa_tree_add_6_33_groupi_n_1537, csa_tree_add_6_33_groupi_n_1538, csa_tree_add_6_33_groupi_n_1539, csa_tree_add_6_33_groupi_n_1540, csa_tree_add_6_33_groupi_n_1541, csa_tree_add_6_33_groupi_n_1542;
  wire csa_tree_add_6_33_groupi_n_1543, csa_tree_add_6_33_groupi_n_1544, csa_tree_add_6_33_groupi_n_1545, csa_tree_add_6_33_groupi_n_1546, csa_tree_add_6_33_groupi_n_1547, csa_tree_add_6_33_groupi_n_1548, csa_tree_add_6_33_groupi_n_1549, csa_tree_add_6_33_groupi_n_1550;
  wire csa_tree_add_6_33_groupi_n_1551, csa_tree_add_6_33_groupi_n_1552, csa_tree_add_6_33_groupi_n_1553, csa_tree_add_6_33_groupi_n_1554, csa_tree_add_6_33_groupi_n_1555, csa_tree_add_6_33_groupi_n_1556, csa_tree_add_6_33_groupi_n_1557, csa_tree_add_6_33_groupi_n_1558;
  wire csa_tree_add_6_33_groupi_n_1559, csa_tree_add_6_33_groupi_n_1560, csa_tree_add_6_33_groupi_n_1561, csa_tree_add_6_33_groupi_n_1562, csa_tree_add_6_33_groupi_n_1563, csa_tree_add_6_33_groupi_n_1564, csa_tree_add_6_33_groupi_n_1565, csa_tree_add_6_33_groupi_n_1566;
  wire csa_tree_add_6_33_groupi_n_1567, csa_tree_add_6_33_groupi_n_1568, csa_tree_add_6_33_groupi_n_1569, csa_tree_add_6_33_groupi_n_1570, csa_tree_add_6_33_groupi_n_1571, csa_tree_add_6_33_groupi_n_1572, csa_tree_add_6_33_groupi_n_1573, csa_tree_add_6_33_groupi_n_1574;
  wire csa_tree_add_6_33_groupi_n_1575, csa_tree_add_6_33_groupi_n_1576, csa_tree_add_6_33_groupi_n_1577, csa_tree_add_6_33_groupi_n_1578, csa_tree_add_6_33_groupi_n_1579, csa_tree_add_6_33_groupi_n_1580, csa_tree_add_6_33_groupi_n_1581, csa_tree_add_6_33_groupi_n_1582;
  wire csa_tree_add_6_33_groupi_n_1583, csa_tree_add_6_33_groupi_n_1584, csa_tree_add_6_33_groupi_n_1585, csa_tree_add_6_33_groupi_n_1586, csa_tree_add_6_33_groupi_n_1587, csa_tree_add_6_33_groupi_n_1588, csa_tree_add_6_33_groupi_n_1589, csa_tree_add_6_33_groupi_n_1590;
  wire csa_tree_add_6_33_groupi_n_1591, csa_tree_add_6_33_groupi_n_1592, csa_tree_add_6_33_groupi_n_1593, csa_tree_add_6_33_groupi_n_1594, csa_tree_add_6_33_groupi_n_1595, csa_tree_add_6_33_groupi_n_1596, csa_tree_add_6_33_groupi_n_1597, csa_tree_add_6_33_groupi_n_1598;
  wire csa_tree_add_6_33_groupi_n_1599, csa_tree_add_6_33_groupi_n_1600, csa_tree_add_6_33_groupi_n_1601, csa_tree_add_6_33_groupi_n_1602, csa_tree_add_6_33_groupi_n_1603, csa_tree_add_6_33_groupi_n_1604, csa_tree_add_6_33_groupi_n_1605, csa_tree_add_6_33_groupi_n_1606;
  wire csa_tree_add_6_33_groupi_n_1607, csa_tree_add_6_33_groupi_n_1608, csa_tree_add_6_33_groupi_n_1609, csa_tree_add_6_33_groupi_n_1610, csa_tree_add_6_33_groupi_n_1611, csa_tree_add_6_33_groupi_n_1612, csa_tree_add_6_33_groupi_n_1613, csa_tree_add_6_33_groupi_n_1614;
  wire csa_tree_add_6_33_groupi_n_1615, csa_tree_add_6_33_groupi_n_1616, csa_tree_add_6_33_groupi_n_1617, csa_tree_add_6_33_groupi_n_1618, csa_tree_add_6_33_groupi_n_1619, csa_tree_add_6_33_groupi_n_1620, csa_tree_add_6_33_groupi_n_1621, csa_tree_add_6_33_groupi_n_1622;
  wire csa_tree_add_6_33_groupi_n_1623, csa_tree_add_6_33_groupi_n_1624, csa_tree_add_6_33_groupi_n_1625, csa_tree_add_6_33_groupi_n_1626, csa_tree_add_6_33_groupi_n_1627, csa_tree_add_6_33_groupi_n_1628, csa_tree_add_6_33_groupi_n_1629, csa_tree_add_6_33_groupi_n_1630;
  wire csa_tree_add_6_33_groupi_n_1631, csa_tree_add_6_33_groupi_n_1632, csa_tree_add_6_33_groupi_n_1633, csa_tree_add_6_33_groupi_n_1634, csa_tree_add_6_33_groupi_n_1635, csa_tree_add_6_33_groupi_n_1636, csa_tree_add_6_33_groupi_n_1637, csa_tree_add_6_33_groupi_n_1638;
  wire csa_tree_add_6_33_groupi_n_1639, csa_tree_add_6_33_groupi_n_1640, csa_tree_add_6_33_groupi_n_1641, csa_tree_add_6_33_groupi_n_1642, csa_tree_add_6_33_groupi_n_1643, csa_tree_add_6_33_groupi_n_1644, csa_tree_add_6_33_groupi_n_1645, csa_tree_add_6_33_groupi_n_1646;
  wire csa_tree_add_6_33_groupi_n_1647, csa_tree_add_6_33_groupi_n_1648, csa_tree_add_6_33_groupi_n_1649, csa_tree_add_6_33_groupi_n_1650, csa_tree_add_6_33_groupi_n_1651, csa_tree_add_6_33_groupi_n_1652, csa_tree_add_6_33_groupi_n_1653, csa_tree_add_6_33_groupi_n_1654;
  wire csa_tree_add_6_33_groupi_n_1655, csa_tree_add_6_33_groupi_n_1656, csa_tree_add_6_33_groupi_n_1657, csa_tree_add_6_33_groupi_n_1658, csa_tree_add_6_33_groupi_n_1659, csa_tree_add_6_33_groupi_n_1660, csa_tree_add_6_33_groupi_n_1661, csa_tree_add_6_33_groupi_n_1662;
  wire csa_tree_add_6_33_groupi_n_1663, csa_tree_add_6_33_groupi_n_1664, csa_tree_add_6_33_groupi_n_1665, csa_tree_add_6_33_groupi_n_1666, csa_tree_add_6_33_groupi_n_1667, csa_tree_add_6_33_groupi_n_1668, csa_tree_add_6_33_groupi_n_1669, csa_tree_add_6_33_groupi_n_1670;
  wire csa_tree_add_6_33_groupi_n_1671, csa_tree_add_6_33_groupi_n_1673, csa_tree_add_6_33_groupi_n_1674, csa_tree_add_6_33_groupi_n_1675, csa_tree_add_6_33_groupi_n_1676, csa_tree_add_6_33_groupi_n_1677, csa_tree_add_6_33_groupi_n_1678, csa_tree_add_6_33_groupi_n_1679;
  wire csa_tree_add_6_33_groupi_n_1680, csa_tree_add_6_33_groupi_n_1681, csa_tree_add_6_33_groupi_n_1682, csa_tree_add_6_33_groupi_n_1683, csa_tree_add_6_33_groupi_n_1684, csa_tree_add_6_33_groupi_n_1685, csa_tree_add_6_33_groupi_n_1686, csa_tree_add_6_33_groupi_n_1687;
  wire csa_tree_add_6_33_groupi_n_1688, csa_tree_add_6_33_groupi_n_1689, csa_tree_add_6_33_groupi_n_1690, csa_tree_add_6_33_groupi_n_1691, csa_tree_add_6_33_groupi_n_1692, csa_tree_add_6_33_groupi_n_1693, csa_tree_add_6_33_groupi_n_1694, csa_tree_add_6_33_groupi_n_1695;
  wire csa_tree_add_6_33_groupi_n_1696, csa_tree_add_6_33_groupi_n_1697, csa_tree_add_6_33_groupi_n_1698, csa_tree_add_6_33_groupi_n_1699, csa_tree_add_6_33_groupi_n_1700, csa_tree_add_6_33_groupi_n_1701, csa_tree_add_6_33_groupi_n_1702, csa_tree_add_6_33_groupi_n_1703;
  wire csa_tree_add_6_33_groupi_n_1704, csa_tree_add_6_33_groupi_n_1705, csa_tree_add_6_33_groupi_n_1706, csa_tree_add_6_33_groupi_n_1707, csa_tree_add_6_33_groupi_n_1709, csa_tree_add_6_33_groupi_n_1710, csa_tree_add_6_33_groupi_n_1711, csa_tree_add_6_33_groupi_n_1712;
  wire csa_tree_add_6_33_groupi_n_1713, csa_tree_add_6_33_groupi_n_1714, csa_tree_add_6_33_groupi_n_1715, csa_tree_add_6_33_groupi_n_1716, csa_tree_add_6_33_groupi_n_1717, csa_tree_add_6_33_groupi_n_1718, csa_tree_add_6_33_groupi_n_1719, csa_tree_add_6_33_groupi_n_1720;
  wire csa_tree_add_6_33_groupi_n_1721, csa_tree_add_6_33_groupi_n_1722, csa_tree_add_6_33_groupi_n_1723, csa_tree_add_6_33_groupi_n_1724, csa_tree_add_6_33_groupi_n_1725, csa_tree_add_6_33_groupi_n_1726, csa_tree_add_6_33_groupi_n_1727, csa_tree_add_6_33_groupi_n_1728;
  wire csa_tree_add_6_33_groupi_n_1729, csa_tree_add_6_33_groupi_n_1730, csa_tree_add_6_33_groupi_n_1731, csa_tree_add_6_33_groupi_n_1732, csa_tree_add_6_33_groupi_n_1733, csa_tree_add_6_33_groupi_n_1734, csa_tree_add_6_33_groupi_n_1735, csa_tree_add_6_33_groupi_n_1736;
  wire csa_tree_add_6_33_groupi_n_1737, csa_tree_add_6_33_groupi_n_1738, csa_tree_add_6_33_groupi_n_1739, csa_tree_add_6_33_groupi_n_1740, csa_tree_add_6_33_groupi_n_1741, csa_tree_add_6_33_groupi_n_1742, csa_tree_add_6_33_groupi_n_1743, csa_tree_add_6_33_groupi_n_1744;
  wire csa_tree_add_6_33_groupi_n_1745, csa_tree_add_6_33_groupi_n_1746, csa_tree_add_6_33_groupi_n_1747, csa_tree_add_6_33_groupi_n_1748, csa_tree_add_6_33_groupi_n_1749, csa_tree_add_6_33_groupi_n_1750, csa_tree_add_6_33_groupi_n_1751, csa_tree_add_6_33_groupi_n_1752;
  wire csa_tree_add_6_33_groupi_n_1753, csa_tree_add_6_33_groupi_n_1754, csa_tree_add_6_33_groupi_n_1755, csa_tree_add_6_33_groupi_n_1756, csa_tree_add_6_33_groupi_n_1757, csa_tree_add_6_33_groupi_n_1758, csa_tree_add_6_33_groupi_n_1759, csa_tree_add_6_33_groupi_n_1760;
  wire csa_tree_add_6_33_groupi_n_1761, csa_tree_add_6_33_groupi_n_1762, csa_tree_add_6_33_groupi_n_1763, csa_tree_add_6_33_groupi_n_1764, csa_tree_add_6_33_groupi_n_1765, csa_tree_add_6_33_groupi_n_1766, csa_tree_add_6_33_groupi_n_1767, csa_tree_add_6_33_groupi_n_1768;
  wire csa_tree_add_6_33_groupi_n_1769, csa_tree_add_6_33_groupi_n_1770, csa_tree_add_6_33_groupi_n_1771, csa_tree_add_6_33_groupi_n_1772, csa_tree_add_6_33_groupi_n_1773, csa_tree_add_6_33_groupi_n_1774, csa_tree_add_6_33_groupi_n_1775, csa_tree_add_6_33_groupi_n_1776;
  wire csa_tree_add_6_33_groupi_n_1777, csa_tree_add_6_33_groupi_n_1778, csa_tree_add_6_33_groupi_n_1779, csa_tree_add_6_33_groupi_n_1780, csa_tree_add_6_33_groupi_n_1781, csa_tree_add_6_33_groupi_n_1782, csa_tree_add_6_33_groupi_n_1783, csa_tree_add_6_33_groupi_n_1784;
  wire csa_tree_add_6_33_groupi_n_1785, csa_tree_add_6_33_groupi_n_1786, csa_tree_add_6_33_groupi_n_1787, csa_tree_add_6_33_groupi_n_1788, csa_tree_add_6_33_groupi_n_1789, csa_tree_add_6_33_groupi_n_1790, csa_tree_add_6_33_groupi_n_1791, csa_tree_add_6_33_groupi_n_1792;
  wire csa_tree_add_6_33_groupi_n_1793, csa_tree_add_6_33_groupi_n_1794, csa_tree_add_6_33_groupi_n_1795, csa_tree_add_6_33_groupi_n_1796, csa_tree_add_6_33_groupi_n_1797, csa_tree_add_6_33_groupi_n_1798, csa_tree_add_6_33_groupi_n_1799, csa_tree_add_6_33_groupi_n_1800;
  wire csa_tree_add_6_33_groupi_n_1801, csa_tree_add_6_33_groupi_n_1802, csa_tree_add_6_33_groupi_n_1803, csa_tree_add_6_33_groupi_n_1804, csa_tree_add_6_33_groupi_n_1805, csa_tree_add_6_33_groupi_n_1806, csa_tree_add_6_33_groupi_n_1807, csa_tree_add_6_33_groupi_n_1808;
  wire csa_tree_add_6_33_groupi_n_1809, csa_tree_add_6_33_groupi_n_1810, csa_tree_add_6_33_groupi_n_1811, csa_tree_add_6_33_groupi_n_1812, csa_tree_add_6_33_groupi_n_1813, csa_tree_add_6_33_groupi_n_1814, csa_tree_add_6_33_groupi_n_1815, csa_tree_add_6_33_groupi_n_1816;
  wire csa_tree_add_6_33_groupi_n_1817, csa_tree_add_6_33_groupi_n_1818, csa_tree_add_6_33_groupi_n_1819, csa_tree_add_6_33_groupi_n_1820, csa_tree_add_6_33_groupi_n_1821, csa_tree_add_6_33_groupi_n_1822, csa_tree_add_6_33_groupi_n_1823, csa_tree_add_6_33_groupi_n_1824;
  wire csa_tree_add_6_33_groupi_n_1825, csa_tree_add_6_33_groupi_n_1826, csa_tree_add_6_33_groupi_n_1827, csa_tree_add_6_33_groupi_n_1828, csa_tree_add_6_33_groupi_n_1829, csa_tree_add_6_33_groupi_n_1830, csa_tree_add_6_33_groupi_n_1831, csa_tree_add_6_33_groupi_n_1832;
  wire csa_tree_add_6_33_groupi_n_1833, csa_tree_add_6_33_groupi_n_1834, csa_tree_add_6_33_groupi_n_1835, csa_tree_add_6_33_groupi_n_1836, csa_tree_add_6_33_groupi_n_1837, csa_tree_add_6_33_groupi_n_1838, csa_tree_add_6_33_groupi_n_1839, csa_tree_add_6_33_groupi_n_1840;
  wire csa_tree_add_6_33_groupi_n_1841, csa_tree_add_6_33_groupi_n_1842, csa_tree_add_6_33_groupi_n_1843, csa_tree_add_6_33_groupi_n_1844, csa_tree_add_6_33_groupi_n_1845, csa_tree_add_6_33_groupi_n_1846, csa_tree_add_6_33_groupi_n_1847, csa_tree_add_6_33_groupi_n_1848;
  wire csa_tree_add_6_33_groupi_n_1849, csa_tree_add_6_33_groupi_n_1850, csa_tree_add_6_33_groupi_n_1851, csa_tree_add_6_33_groupi_n_1852, csa_tree_add_6_33_groupi_n_1853, csa_tree_add_6_33_groupi_n_1854, csa_tree_add_6_33_groupi_n_1855, csa_tree_add_6_33_groupi_n_1856;
  wire csa_tree_add_6_33_groupi_n_1857, csa_tree_add_6_33_groupi_n_1858, csa_tree_add_6_33_groupi_n_1859, csa_tree_add_6_33_groupi_n_1860, csa_tree_add_6_33_groupi_n_1861, csa_tree_add_6_33_groupi_n_1862, csa_tree_add_6_33_groupi_n_1863, csa_tree_add_6_33_groupi_n_1864;
  wire csa_tree_add_6_33_groupi_n_1866, csa_tree_add_6_33_groupi_n_1867, csa_tree_add_6_33_groupi_n_1868, csa_tree_add_6_33_groupi_n_1869, csa_tree_add_6_33_groupi_n_1870, csa_tree_add_6_33_groupi_n_1871, csa_tree_add_6_33_groupi_n_1872, csa_tree_add_6_33_groupi_n_1873;
  wire csa_tree_add_6_33_groupi_n_1874, csa_tree_add_6_33_groupi_n_1875, csa_tree_add_6_33_groupi_n_1876, csa_tree_add_6_33_groupi_n_1877, csa_tree_add_6_33_groupi_n_1878, csa_tree_add_6_33_groupi_n_1879, csa_tree_add_6_33_groupi_n_1880, csa_tree_add_6_33_groupi_n_1881;
  wire csa_tree_add_6_33_groupi_n_1882, csa_tree_add_6_33_groupi_n_1883, csa_tree_add_6_33_groupi_n_1884, csa_tree_add_6_33_groupi_n_1885, csa_tree_add_6_33_groupi_n_1886, csa_tree_add_6_33_groupi_n_1887, csa_tree_add_6_33_groupi_n_1888, csa_tree_add_6_33_groupi_n_1889;
  wire csa_tree_add_6_33_groupi_n_1890, csa_tree_add_6_33_groupi_n_1891, csa_tree_add_6_33_groupi_n_1892, csa_tree_add_6_33_groupi_n_1893, csa_tree_add_6_33_groupi_n_1894, csa_tree_add_6_33_groupi_n_1896, csa_tree_add_6_33_groupi_n_1897, csa_tree_add_6_33_groupi_n_1898;
  wire csa_tree_add_6_33_groupi_n_1899, csa_tree_add_6_33_groupi_n_1900, csa_tree_add_6_33_groupi_n_1901, csa_tree_add_6_33_groupi_n_1902, csa_tree_add_6_33_groupi_n_1903, csa_tree_add_6_33_groupi_n_1904, csa_tree_add_6_33_groupi_n_1905, csa_tree_add_6_33_groupi_n_1906;
  wire csa_tree_add_6_33_groupi_n_1907, csa_tree_add_6_33_groupi_n_1908, csa_tree_add_6_33_groupi_n_1909, csa_tree_add_6_33_groupi_n_1910, csa_tree_add_6_33_groupi_n_1911, csa_tree_add_6_33_groupi_n_1912, csa_tree_add_6_33_groupi_n_1913, csa_tree_add_6_33_groupi_n_1914;
  wire csa_tree_add_6_33_groupi_n_1915, csa_tree_add_6_33_groupi_n_1916, csa_tree_add_6_33_groupi_n_1917, csa_tree_add_6_33_groupi_n_1918, csa_tree_add_6_33_groupi_n_1919, csa_tree_add_6_33_groupi_n_1920, csa_tree_add_6_33_groupi_n_1921, csa_tree_add_6_33_groupi_n_1922;
  wire csa_tree_add_6_33_groupi_n_1923, csa_tree_add_6_33_groupi_n_1924, csa_tree_add_6_33_groupi_n_1925, csa_tree_add_6_33_groupi_n_1926, csa_tree_add_6_33_groupi_n_1927, csa_tree_add_6_33_groupi_n_1928, csa_tree_add_6_33_groupi_n_1929, csa_tree_add_6_33_groupi_n_1930;
  wire csa_tree_add_6_33_groupi_n_1931, csa_tree_add_6_33_groupi_n_1932, csa_tree_add_6_33_groupi_n_1933, csa_tree_add_6_33_groupi_n_1934, csa_tree_add_6_33_groupi_n_1935, csa_tree_add_6_33_groupi_n_1936, csa_tree_add_6_33_groupi_n_1937, csa_tree_add_6_33_groupi_n_1938;
  wire csa_tree_add_6_33_groupi_n_1939, csa_tree_add_6_33_groupi_n_1941, csa_tree_add_6_33_groupi_n_1942, csa_tree_add_6_33_groupi_n_1943, csa_tree_add_6_33_groupi_n_1944, csa_tree_add_6_33_groupi_n_1945, csa_tree_add_6_33_groupi_n_1946, csa_tree_add_6_33_groupi_n_1947;
  wire csa_tree_add_6_33_groupi_n_1948, csa_tree_add_6_33_groupi_n_1949, csa_tree_add_6_33_groupi_n_1950, csa_tree_add_6_33_groupi_n_1951, csa_tree_add_6_33_groupi_n_1952, csa_tree_add_6_33_groupi_n_1953, csa_tree_add_6_33_groupi_n_1954, csa_tree_add_6_33_groupi_n_1955;
  wire csa_tree_add_6_33_groupi_n_1956, csa_tree_add_6_33_groupi_n_1958, csa_tree_add_6_33_groupi_n_1959, csa_tree_add_6_33_groupi_n_1960, csa_tree_add_6_33_groupi_n_1961, csa_tree_add_6_33_groupi_n_1962, csa_tree_add_6_33_groupi_n_1963, csa_tree_add_6_33_groupi_n_1964;
  wire csa_tree_add_6_33_groupi_n_1965, csa_tree_add_6_33_groupi_n_1966, csa_tree_add_6_33_groupi_n_1967, csa_tree_add_6_33_groupi_n_1968, csa_tree_add_6_33_groupi_n_1969, csa_tree_add_6_33_groupi_n_1970, csa_tree_add_6_33_groupi_n_1971, csa_tree_add_6_33_groupi_n_1972;
  wire csa_tree_add_6_33_groupi_n_1973, csa_tree_add_6_33_groupi_n_1975, csa_tree_add_6_33_groupi_n_1976, csa_tree_add_6_33_groupi_n_1978, csa_tree_add_6_33_groupi_n_1979, csa_tree_add_6_33_groupi_n_1980, csa_tree_add_6_33_groupi_n_1981, csa_tree_add_6_33_groupi_n_1982;
  wire csa_tree_add_6_33_groupi_n_1983, csa_tree_add_6_33_groupi_n_1984, csa_tree_add_6_33_groupi_n_1985, csa_tree_add_6_33_groupi_n_1986, csa_tree_add_6_33_groupi_n_1987, csa_tree_add_6_33_groupi_n_1988, csa_tree_add_6_33_groupi_n_1989, csa_tree_add_6_33_groupi_n_1990;
  wire csa_tree_add_6_33_groupi_n_1992, csa_tree_add_6_33_groupi_n_1993, csa_tree_add_6_33_groupi_n_1994, csa_tree_add_6_33_groupi_n_1995, csa_tree_add_6_33_groupi_n_1996, csa_tree_add_6_33_groupi_n_1997, csa_tree_add_6_33_groupi_n_1998, csa_tree_add_6_33_groupi_n_1999;
  wire csa_tree_add_6_33_groupi_n_2000, csa_tree_add_6_33_groupi_n_2001, csa_tree_add_6_33_groupi_n_2002, csa_tree_add_6_33_groupi_n_2003, csa_tree_add_6_33_groupi_n_2004, csa_tree_add_6_33_groupi_n_2005, csa_tree_add_6_33_groupi_n_2006, csa_tree_add_6_33_groupi_n_2007;
  wire csa_tree_add_6_33_groupi_n_2008, csa_tree_add_6_33_groupi_n_2009, csa_tree_add_6_33_groupi_n_2010, csa_tree_add_6_33_groupi_n_2011, csa_tree_add_6_33_groupi_n_2012, csa_tree_add_6_33_groupi_n_2013, csa_tree_add_6_33_groupi_n_2014, csa_tree_add_6_33_groupi_n_2015;
  wire csa_tree_add_6_33_groupi_n_2016, csa_tree_add_6_33_groupi_n_2017, csa_tree_add_6_33_groupi_n_2018, csa_tree_add_6_33_groupi_n_2019, csa_tree_add_6_33_groupi_n_2020, csa_tree_add_6_33_groupi_n_2021, csa_tree_add_6_33_groupi_n_2022, csa_tree_add_6_33_groupi_n_2023;
  wire csa_tree_add_6_33_groupi_n_2024, csa_tree_add_6_33_groupi_n_2025, csa_tree_add_6_33_groupi_n_2026, csa_tree_add_6_33_groupi_n_2027, csa_tree_add_6_33_groupi_n_2028, csa_tree_add_6_33_groupi_n_2029, csa_tree_add_6_33_groupi_n_2030, csa_tree_add_6_33_groupi_n_2031;
  wire csa_tree_add_6_33_groupi_n_2032, csa_tree_add_6_33_groupi_n_2033, csa_tree_add_6_33_groupi_n_2034, csa_tree_add_6_33_groupi_n_2035, csa_tree_add_6_33_groupi_n_2036, csa_tree_add_6_33_groupi_n_2037, csa_tree_add_6_33_groupi_n_2038, csa_tree_add_6_33_groupi_n_2039;
  wire csa_tree_add_6_33_groupi_n_2040, csa_tree_add_6_33_groupi_n_2041, csa_tree_add_6_33_groupi_n_2042, csa_tree_add_6_33_groupi_n_2043, csa_tree_add_6_33_groupi_n_2044, csa_tree_add_6_33_groupi_n_2045, csa_tree_add_6_33_groupi_n_2046, csa_tree_add_6_33_groupi_n_2047;
  wire csa_tree_add_6_33_groupi_n_2048, csa_tree_add_6_33_groupi_n_2049, csa_tree_add_6_33_groupi_n_2050, csa_tree_add_6_33_groupi_n_2051, csa_tree_add_6_33_groupi_n_2052, csa_tree_add_6_33_groupi_n_2053, csa_tree_add_6_33_groupi_n_2054, csa_tree_add_6_33_groupi_n_2055;
  wire csa_tree_add_6_33_groupi_n_2056, csa_tree_add_6_33_groupi_n_2057, csa_tree_add_6_33_groupi_n_2058, csa_tree_add_6_33_groupi_n_2059, csa_tree_add_6_33_groupi_n_2060, csa_tree_add_6_33_groupi_n_2061, csa_tree_add_6_33_groupi_n_2062, csa_tree_add_6_33_groupi_n_2063;
  wire csa_tree_add_6_33_groupi_n_2064, csa_tree_add_6_33_groupi_n_2065, csa_tree_add_6_33_groupi_n_2066, csa_tree_add_6_33_groupi_n_2067, csa_tree_add_6_33_groupi_n_2068, csa_tree_add_6_33_groupi_n_2069, csa_tree_add_6_33_groupi_n_2070, csa_tree_add_6_33_groupi_n_2071;
  wire csa_tree_add_6_33_groupi_n_2072, csa_tree_add_6_33_groupi_n_2073, csa_tree_add_6_33_groupi_n_2074, csa_tree_add_6_33_groupi_n_2075, csa_tree_add_6_33_groupi_n_2076, csa_tree_add_6_33_groupi_n_2077, csa_tree_add_6_33_groupi_n_2078, csa_tree_add_6_33_groupi_n_2079;
  wire csa_tree_add_6_33_groupi_n_2080, csa_tree_add_6_33_groupi_n_2081, csa_tree_add_6_33_groupi_n_2082, csa_tree_add_6_33_groupi_n_2083, csa_tree_add_6_33_groupi_n_2084, csa_tree_add_6_33_groupi_n_2085, csa_tree_add_6_33_groupi_n_2086, csa_tree_add_6_33_groupi_n_2087;
  wire csa_tree_add_6_33_groupi_n_2088, csa_tree_add_6_33_groupi_n_2089, csa_tree_add_6_33_groupi_n_2090, csa_tree_add_6_33_groupi_n_2091, csa_tree_add_6_33_groupi_n_2092, csa_tree_add_6_33_groupi_n_2093, csa_tree_add_6_33_groupi_n_2094, csa_tree_add_6_33_groupi_n_2095;
  wire csa_tree_add_6_33_groupi_n_2096, csa_tree_add_6_33_groupi_n_2097, csa_tree_add_6_33_groupi_n_2098, csa_tree_add_6_33_groupi_n_2099, csa_tree_add_6_33_groupi_n_2100, csa_tree_add_6_33_groupi_n_2101, csa_tree_add_6_33_groupi_n_2102, csa_tree_add_6_33_groupi_n_2103;
  wire csa_tree_add_6_33_groupi_n_2104, csa_tree_add_6_33_groupi_n_2105, csa_tree_add_6_33_groupi_n_2106, csa_tree_add_6_33_groupi_n_2107, csa_tree_add_6_33_groupi_n_2108, csa_tree_add_6_33_groupi_n_2109, csa_tree_add_6_33_groupi_n_2110, csa_tree_add_6_33_groupi_n_2111;
  wire csa_tree_add_6_33_groupi_n_2112, csa_tree_add_6_33_groupi_n_2113, csa_tree_add_6_33_groupi_n_2114, csa_tree_add_6_33_groupi_n_2115, csa_tree_add_6_33_groupi_n_2116, csa_tree_add_6_33_groupi_n_2117, csa_tree_add_6_33_groupi_n_2118, csa_tree_add_6_33_groupi_n_2119;
  wire csa_tree_add_6_33_groupi_n_2120, csa_tree_add_6_33_groupi_n_2121, csa_tree_add_6_33_groupi_n_2122, csa_tree_add_6_33_groupi_n_2123, csa_tree_add_6_33_groupi_n_2124, csa_tree_add_6_33_groupi_n_2125, csa_tree_add_6_33_groupi_n_2126, csa_tree_add_6_33_groupi_n_2127;
  wire csa_tree_add_6_33_groupi_n_2128, csa_tree_add_6_33_groupi_n_2129, csa_tree_add_6_33_groupi_n_2130, csa_tree_add_6_33_groupi_n_2131, csa_tree_add_6_33_groupi_n_2132, csa_tree_add_6_33_groupi_n_2133, csa_tree_add_6_33_groupi_n_2134, csa_tree_add_6_33_groupi_n_2135;
  wire csa_tree_add_6_33_groupi_n_2136, csa_tree_add_6_33_groupi_n_2137, csa_tree_add_6_33_groupi_n_2138, csa_tree_add_6_33_groupi_n_2139, csa_tree_add_6_33_groupi_n_2140, csa_tree_add_6_33_groupi_n_2141, csa_tree_add_6_33_groupi_n_2142, csa_tree_add_6_33_groupi_n_2143;
  wire csa_tree_add_6_33_groupi_n_2144, csa_tree_add_6_33_groupi_n_2145, csa_tree_add_6_33_groupi_n_2146, csa_tree_add_6_33_groupi_n_2147, csa_tree_add_6_33_groupi_n_2148, csa_tree_add_6_33_groupi_n_2149, csa_tree_add_6_33_groupi_n_2150, csa_tree_add_6_33_groupi_n_2151;
  wire csa_tree_add_6_33_groupi_n_2152, csa_tree_add_6_33_groupi_n_2153, csa_tree_add_6_33_groupi_n_2154, csa_tree_add_6_33_groupi_n_2155, csa_tree_add_6_33_groupi_n_2156, csa_tree_add_6_33_groupi_n_2157, csa_tree_add_6_33_groupi_n_2158, csa_tree_add_6_33_groupi_n_2159;
  wire csa_tree_add_6_33_groupi_n_2160, csa_tree_add_6_33_groupi_n_2161, csa_tree_add_6_33_groupi_n_2162, csa_tree_add_6_33_groupi_n_2163, csa_tree_add_6_33_groupi_n_2164, csa_tree_add_6_33_groupi_n_2165, csa_tree_add_6_33_groupi_n_2166, csa_tree_add_6_33_groupi_n_2167;
  wire csa_tree_add_6_33_groupi_n_2168, csa_tree_add_6_33_groupi_n_2169, csa_tree_add_6_33_groupi_n_2170, csa_tree_add_6_33_groupi_n_2171, csa_tree_add_6_33_groupi_n_2172, csa_tree_add_6_33_groupi_n_2173, csa_tree_add_6_33_groupi_n_2174, csa_tree_add_6_33_groupi_n_2175;
  wire csa_tree_add_6_33_groupi_n_2176, csa_tree_add_6_33_groupi_n_2177, csa_tree_add_6_33_groupi_n_2178, csa_tree_add_6_33_groupi_n_2179, csa_tree_add_6_33_groupi_n_2180, csa_tree_add_6_33_groupi_n_2181, csa_tree_add_6_33_groupi_n_2182, csa_tree_add_6_33_groupi_n_2183;
  wire csa_tree_add_6_33_groupi_n_2184, csa_tree_add_6_33_groupi_n_2185, csa_tree_add_6_33_groupi_n_2186, csa_tree_add_6_33_groupi_n_2187, csa_tree_add_6_33_groupi_n_2188, csa_tree_add_6_33_groupi_n_2189, csa_tree_add_6_33_groupi_n_2190, csa_tree_add_6_33_groupi_n_2191;
  wire csa_tree_add_6_33_groupi_n_2192, csa_tree_add_6_33_groupi_n_2193, csa_tree_add_6_33_groupi_n_2194, csa_tree_add_6_33_groupi_n_2195, csa_tree_add_6_33_groupi_n_2196, csa_tree_add_6_33_groupi_n_2197, csa_tree_add_6_33_groupi_n_2198, csa_tree_add_6_33_groupi_n_2199;
  wire csa_tree_add_6_33_groupi_n_2200, csa_tree_add_6_33_groupi_n_2201, csa_tree_add_6_33_groupi_n_2202, csa_tree_add_6_33_groupi_n_2203, csa_tree_add_6_33_groupi_n_2204, csa_tree_add_6_33_groupi_n_2205, csa_tree_add_6_33_groupi_n_2206, csa_tree_add_6_33_groupi_n_2207;
  wire csa_tree_add_6_33_groupi_n_2208, csa_tree_add_6_33_groupi_n_2209, csa_tree_add_6_33_groupi_n_2210, csa_tree_add_6_33_groupi_n_2211, csa_tree_add_6_33_groupi_n_2212, csa_tree_add_6_33_groupi_n_2213, csa_tree_add_6_33_groupi_n_2214, csa_tree_add_6_33_groupi_n_2215;
  wire csa_tree_add_6_33_groupi_n_2216, csa_tree_add_6_33_groupi_n_2217, csa_tree_add_6_33_groupi_n_2218, csa_tree_add_6_33_groupi_n_2219, csa_tree_add_6_33_groupi_n_2220, csa_tree_add_6_33_groupi_n_2221, csa_tree_add_6_33_groupi_n_2222, csa_tree_add_6_33_groupi_n_2223;
  wire csa_tree_add_6_33_groupi_n_2224, csa_tree_add_6_33_groupi_n_2225, csa_tree_add_6_33_groupi_n_2226, csa_tree_add_6_33_groupi_n_2227, csa_tree_add_6_33_groupi_n_2228, csa_tree_add_6_33_groupi_n_2229, csa_tree_add_6_33_groupi_n_2230, csa_tree_add_6_33_groupi_n_2231;
  wire csa_tree_add_6_33_groupi_n_2232, csa_tree_add_6_33_groupi_n_2233, csa_tree_add_6_33_groupi_n_2234, csa_tree_add_6_33_groupi_n_2235, csa_tree_add_6_33_groupi_n_2236, csa_tree_add_6_33_groupi_n_2237, csa_tree_add_6_33_groupi_n_2238, csa_tree_add_6_33_groupi_n_2239;
  wire csa_tree_add_6_33_groupi_n_2240, csa_tree_add_6_33_groupi_n_2241, csa_tree_add_6_33_groupi_n_2242, csa_tree_add_6_33_groupi_n_2243, csa_tree_add_6_33_groupi_n_2244, csa_tree_add_6_33_groupi_n_2245, csa_tree_add_6_33_groupi_n_2246, csa_tree_add_6_33_groupi_n_2247;
  wire csa_tree_add_6_33_groupi_n_2248, csa_tree_add_6_33_groupi_n_2249, csa_tree_add_6_33_groupi_n_2250, csa_tree_add_6_33_groupi_n_2251, csa_tree_add_6_33_groupi_n_2252, csa_tree_add_6_33_groupi_n_2253, csa_tree_add_6_33_groupi_n_2254, csa_tree_add_6_33_groupi_n_2255;
  wire csa_tree_add_6_33_groupi_n_2256, csa_tree_add_6_33_groupi_n_2257, csa_tree_add_6_33_groupi_n_2258, csa_tree_add_6_33_groupi_n_2259, csa_tree_add_6_33_groupi_n_2260, csa_tree_add_6_33_groupi_n_2261, csa_tree_add_6_33_groupi_n_2262, csa_tree_add_6_33_groupi_n_2263;
  wire csa_tree_add_6_33_groupi_n_2264, csa_tree_add_6_33_groupi_n_2265, csa_tree_add_6_33_groupi_n_2266, csa_tree_add_6_33_groupi_n_2267, csa_tree_add_6_33_groupi_n_2268, csa_tree_add_6_33_groupi_n_2269, csa_tree_add_6_33_groupi_n_2270, csa_tree_add_6_33_groupi_n_2271;
  wire csa_tree_add_6_33_groupi_n_2272, csa_tree_add_6_33_groupi_n_2273, csa_tree_add_6_33_groupi_n_2274, csa_tree_add_6_33_groupi_n_2275, csa_tree_add_6_33_groupi_n_2276, csa_tree_add_6_33_groupi_n_2277, csa_tree_add_6_33_groupi_n_2278, csa_tree_add_6_33_groupi_n_2279;
  wire csa_tree_add_6_33_groupi_n_2280, csa_tree_add_6_33_groupi_n_2281, csa_tree_add_6_33_groupi_n_2282, csa_tree_add_6_33_groupi_n_2283, csa_tree_add_6_33_groupi_n_2284, csa_tree_add_6_33_groupi_n_2285, csa_tree_add_6_33_groupi_n_2286, csa_tree_add_6_33_groupi_n_2287;
  wire csa_tree_add_6_33_groupi_n_2288, csa_tree_add_6_33_groupi_n_2289, csa_tree_add_6_33_groupi_n_2290, csa_tree_add_6_33_groupi_n_2291, csa_tree_add_6_33_groupi_n_2292, csa_tree_add_6_33_groupi_n_2293, csa_tree_add_6_33_groupi_n_2294, csa_tree_add_6_33_groupi_n_2295;
  wire csa_tree_add_6_33_groupi_n_2296, csa_tree_add_6_33_groupi_n_2297, csa_tree_add_6_33_groupi_n_2298, csa_tree_add_6_33_groupi_n_2299, csa_tree_add_6_33_groupi_n_2300, csa_tree_add_6_33_groupi_n_2301, csa_tree_add_6_33_groupi_n_2302, csa_tree_add_6_33_groupi_n_2303;
  wire csa_tree_add_6_33_groupi_n_2304, csa_tree_add_6_33_groupi_n_2305, csa_tree_add_6_33_groupi_n_2306, csa_tree_add_6_33_groupi_n_2307, csa_tree_add_6_33_groupi_n_2308, csa_tree_add_6_33_groupi_n_2309, csa_tree_add_6_33_groupi_n_2310, csa_tree_add_6_33_groupi_n_2311;
  wire csa_tree_add_6_33_groupi_n_2312, csa_tree_add_6_33_groupi_n_2313, csa_tree_add_6_33_groupi_n_2314, csa_tree_add_6_33_groupi_n_2315, csa_tree_add_6_33_groupi_n_2316, csa_tree_add_6_33_groupi_n_2317, csa_tree_add_6_33_groupi_n_2318, csa_tree_add_6_33_groupi_n_2319;
  wire csa_tree_add_6_33_groupi_n_2320, csa_tree_add_6_33_groupi_n_2321, csa_tree_add_6_33_groupi_n_2322, csa_tree_add_6_33_groupi_n_2323, csa_tree_add_6_33_groupi_n_2324, csa_tree_add_6_33_groupi_n_2325, csa_tree_add_6_33_groupi_n_2326, csa_tree_add_6_33_groupi_n_2327;
  wire csa_tree_add_6_33_groupi_n_2328, csa_tree_add_6_33_groupi_n_2329, csa_tree_add_6_33_groupi_n_2330, csa_tree_add_6_33_groupi_n_2331, csa_tree_add_6_33_groupi_n_2332, csa_tree_add_6_33_groupi_n_2333, csa_tree_add_6_33_groupi_n_2334, csa_tree_add_6_33_groupi_n_2335;
  wire csa_tree_add_6_33_groupi_n_2336, csa_tree_add_6_33_groupi_n_2337, csa_tree_add_6_33_groupi_n_2338, csa_tree_add_6_33_groupi_n_2339, csa_tree_add_6_33_groupi_n_2340, csa_tree_add_6_33_groupi_n_2341, csa_tree_add_6_33_groupi_n_2342, csa_tree_add_6_33_groupi_n_2343;
  wire csa_tree_add_6_33_groupi_n_2344, csa_tree_add_6_33_groupi_n_2345, csa_tree_add_6_33_groupi_n_2346, csa_tree_add_6_33_groupi_n_2347, csa_tree_add_6_33_groupi_n_2348, csa_tree_add_6_33_groupi_n_2349, csa_tree_add_6_33_groupi_n_2350, csa_tree_add_6_33_groupi_n_2351;
  wire csa_tree_add_6_33_groupi_n_2352, csa_tree_add_6_33_groupi_n_2353, csa_tree_add_6_33_groupi_n_2354, csa_tree_add_6_33_groupi_n_2355, csa_tree_add_6_33_groupi_n_2356, csa_tree_add_6_33_groupi_n_2357, csa_tree_add_6_33_groupi_n_2358, csa_tree_add_6_33_groupi_n_2359;
  wire csa_tree_add_6_33_groupi_n_2360, csa_tree_add_6_33_groupi_n_2361, csa_tree_add_6_33_groupi_n_2362, csa_tree_add_6_33_groupi_n_2363, csa_tree_add_6_33_groupi_n_2364, csa_tree_add_6_33_groupi_n_2365, csa_tree_add_6_33_groupi_n_2366, csa_tree_add_6_33_groupi_n_2367;
  wire csa_tree_add_6_33_groupi_n_2368, csa_tree_add_6_33_groupi_n_2369, csa_tree_add_6_33_groupi_n_2370, csa_tree_add_6_33_groupi_n_2371, csa_tree_add_6_33_groupi_n_2372, csa_tree_add_6_33_groupi_n_2373, csa_tree_add_6_33_groupi_n_2374, csa_tree_add_6_33_groupi_n_2376;
  wire csa_tree_add_6_33_groupi_n_2377, csa_tree_add_6_33_groupi_n_2378, csa_tree_add_6_33_groupi_n_2379, csa_tree_add_6_33_groupi_n_2380, csa_tree_add_6_33_groupi_n_2381, csa_tree_add_6_33_groupi_n_2382, csa_tree_add_6_33_groupi_n_2383, csa_tree_add_6_33_groupi_n_2384;
  wire csa_tree_add_6_33_groupi_n_2385, csa_tree_add_6_33_groupi_n_2386, csa_tree_add_6_33_groupi_n_2387, csa_tree_add_6_33_groupi_n_2388, csa_tree_add_6_33_groupi_n_2389, csa_tree_add_6_33_groupi_n_2390, csa_tree_add_6_33_groupi_n_2391, csa_tree_add_6_33_groupi_n_2392;
  wire csa_tree_add_6_33_groupi_n_2393, csa_tree_add_6_33_groupi_n_2394, csa_tree_add_6_33_groupi_n_2395, csa_tree_add_6_33_groupi_n_2396, csa_tree_add_6_33_groupi_n_2397, csa_tree_add_6_33_groupi_n_2398, csa_tree_add_6_33_groupi_n_2399, csa_tree_add_6_33_groupi_n_2400;
  wire csa_tree_add_6_33_groupi_n_2401, csa_tree_add_6_33_groupi_n_2402, csa_tree_add_6_33_groupi_n_2403, csa_tree_add_6_33_groupi_n_2404, csa_tree_add_6_33_groupi_n_2405, csa_tree_add_6_33_groupi_n_2406, csa_tree_add_6_33_groupi_n_2407, csa_tree_add_6_33_groupi_n_2408;
  wire csa_tree_add_6_33_groupi_n_2409, csa_tree_add_6_33_groupi_n_2410, csa_tree_add_6_33_groupi_n_2411, csa_tree_add_6_33_groupi_n_2412, csa_tree_add_6_33_groupi_n_2413, csa_tree_add_6_33_groupi_n_2414, csa_tree_add_6_33_groupi_n_2415, csa_tree_add_6_33_groupi_n_2416;
  wire csa_tree_add_6_33_groupi_n_2417, csa_tree_add_6_33_groupi_n_2418, csa_tree_add_6_33_groupi_n_2419, csa_tree_add_6_33_groupi_n_2420, csa_tree_add_6_33_groupi_n_2421, csa_tree_add_6_33_groupi_n_2422, csa_tree_add_6_33_groupi_n_2423, csa_tree_add_6_33_groupi_n_2424;
  wire csa_tree_add_6_33_groupi_n_2425, csa_tree_add_6_33_groupi_n_2426, csa_tree_add_6_33_groupi_n_2427, csa_tree_add_6_33_groupi_n_2428, csa_tree_add_6_33_groupi_n_2429, csa_tree_add_6_33_groupi_n_2430, csa_tree_add_6_33_groupi_n_2431, csa_tree_add_6_33_groupi_n_2432;
  wire csa_tree_add_6_33_groupi_n_2433, csa_tree_add_6_33_groupi_n_2434, csa_tree_add_6_33_groupi_n_2435, csa_tree_add_6_33_groupi_n_2436, csa_tree_add_6_33_groupi_n_2437, csa_tree_add_6_33_groupi_n_2438, csa_tree_add_6_33_groupi_n_2439, csa_tree_add_6_33_groupi_n_2440;
  wire csa_tree_add_6_33_groupi_n_2441, csa_tree_add_6_33_groupi_n_2442, csa_tree_add_6_33_groupi_n_2443, csa_tree_add_6_33_groupi_n_2444, csa_tree_add_6_33_groupi_n_2445, csa_tree_add_6_33_groupi_n_2446, csa_tree_add_6_33_groupi_n_2447, csa_tree_add_6_33_groupi_n_2448;
  wire csa_tree_add_6_33_groupi_n_2449, csa_tree_add_6_33_groupi_n_2450, csa_tree_add_6_33_groupi_n_2451, csa_tree_add_6_33_groupi_n_2452, csa_tree_add_6_33_groupi_n_2453, csa_tree_add_6_33_groupi_n_2454, csa_tree_add_6_33_groupi_n_2455, csa_tree_add_6_33_groupi_n_2456;
  wire csa_tree_add_6_33_groupi_n_2457, csa_tree_add_6_33_groupi_n_2458, csa_tree_add_6_33_groupi_n_2459, csa_tree_add_6_33_groupi_n_2460, csa_tree_add_6_33_groupi_n_2461, csa_tree_add_6_33_groupi_n_2462, csa_tree_add_6_33_groupi_n_2463, csa_tree_add_6_33_groupi_n_2464;
  wire csa_tree_add_6_33_groupi_n_2465, csa_tree_add_6_33_groupi_n_2466, csa_tree_add_6_33_groupi_n_2467, csa_tree_add_6_33_groupi_n_2468, csa_tree_add_6_33_groupi_n_2469, csa_tree_add_6_33_groupi_n_2470, csa_tree_add_6_33_groupi_n_2471, csa_tree_add_6_33_groupi_n_2472;
  wire csa_tree_add_6_33_groupi_n_2473, csa_tree_add_6_33_groupi_n_2474, csa_tree_add_6_33_groupi_n_2475, csa_tree_add_6_33_groupi_n_2476, csa_tree_add_6_33_groupi_n_2477, csa_tree_add_6_33_groupi_n_2478, csa_tree_add_6_33_groupi_n_2479, csa_tree_add_6_33_groupi_n_2480;
  wire csa_tree_add_6_33_groupi_n_2481, csa_tree_add_6_33_groupi_n_2482, csa_tree_add_6_33_groupi_n_2483, csa_tree_add_6_33_groupi_n_2484, csa_tree_add_6_33_groupi_n_2485, csa_tree_add_6_33_groupi_n_2486, csa_tree_add_6_33_groupi_n_2487, csa_tree_add_6_33_groupi_n_2488;
  wire csa_tree_add_6_33_groupi_n_2489, csa_tree_add_6_33_groupi_n_2490, csa_tree_add_6_33_groupi_n_2491, csa_tree_add_6_33_groupi_n_2492, csa_tree_add_6_33_groupi_n_2493, csa_tree_add_6_33_groupi_n_2494, csa_tree_add_6_33_groupi_n_2495, csa_tree_add_6_33_groupi_n_2496;
  wire csa_tree_add_6_33_groupi_n_2497, csa_tree_add_6_33_groupi_n_2498, csa_tree_add_6_33_groupi_n_2499, csa_tree_add_6_33_groupi_n_2500, csa_tree_add_6_33_groupi_n_2501, csa_tree_add_6_33_groupi_n_2502, csa_tree_add_6_33_groupi_n_2503, csa_tree_add_6_33_groupi_n_2504;
  wire csa_tree_add_6_33_groupi_n_2505, csa_tree_add_6_33_groupi_n_2506, csa_tree_add_6_33_groupi_n_2507, csa_tree_add_6_33_groupi_n_2508, csa_tree_add_6_33_groupi_n_2509, csa_tree_add_6_33_groupi_n_2510, csa_tree_add_6_33_groupi_n_2511, csa_tree_add_6_33_groupi_n_2512;
  wire csa_tree_add_6_33_groupi_n_2513, csa_tree_add_6_33_groupi_n_2514, csa_tree_add_6_33_groupi_n_2515, csa_tree_add_6_33_groupi_n_2516, csa_tree_add_6_33_groupi_n_2517, csa_tree_add_6_33_groupi_n_2518, csa_tree_add_6_33_groupi_n_2519, csa_tree_add_6_33_groupi_n_2520;
  wire csa_tree_add_6_33_groupi_n_2521, csa_tree_add_6_33_groupi_n_2522, csa_tree_add_6_33_groupi_n_2523, csa_tree_add_6_33_groupi_n_2524, csa_tree_add_6_33_groupi_n_2525, csa_tree_add_6_33_groupi_n_2526, csa_tree_add_6_33_groupi_n_2527, csa_tree_add_6_33_groupi_n_2528;
  wire csa_tree_add_6_33_groupi_n_2529, csa_tree_add_6_33_groupi_n_2530, csa_tree_add_6_33_groupi_n_2531, csa_tree_add_6_33_groupi_n_2532, csa_tree_add_6_33_groupi_n_2533, csa_tree_add_6_33_groupi_n_2534, csa_tree_add_6_33_groupi_n_2535, csa_tree_add_6_33_groupi_n_2536;
  wire csa_tree_add_6_33_groupi_n_2537, csa_tree_add_6_33_groupi_n_2538, csa_tree_add_6_33_groupi_n_2539, csa_tree_add_6_33_groupi_n_2540, csa_tree_add_6_33_groupi_n_2541, csa_tree_add_6_33_groupi_n_2542, csa_tree_add_6_33_groupi_n_2543, csa_tree_add_6_33_groupi_n_2544;
  wire csa_tree_add_6_33_groupi_n_2545, csa_tree_add_6_33_groupi_n_2546, csa_tree_add_6_33_groupi_n_2547, csa_tree_add_6_33_groupi_n_2548, csa_tree_add_6_33_groupi_n_2549, csa_tree_add_6_33_groupi_n_2550, csa_tree_add_6_33_groupi_n_2551, csa_tree_add_6_33_groupi_n_2552;
  wire csa_tree_add_6_33_groupi_n_2553, csa_tree_add_6_33_groupi_n_2554, csa_tree_add_6_33_groupi_n_2555, csa_tree_add_6_33_groupi_n_2556, csa_tree_add_6_33_groupi_n_2557, csa_tree_add_6_33_groupi_n_2558, csa_tree_add_6_33_groupi_n_2559, csa_tree_add_6_33_groupi_n_2560;
  wire csa_tree_add_6_33_groupi_n_2561, csa_tree_add_6_33_groupi_n_2562, csa_tree_add_6_33_groupi_n_2563, csa_tree_add_6_33_groupi_n_2564, csa_tree_add_6_33_groupi_n_2565, csa_tree_add_6_33_groupi_n_2566, csa_tree_add_6_33_groupi_n_2567, csa_tree_add_6_33_groupi_n_2568;
  wire csa_tree_add_6_33_groupi_n_2569, csa_tree_add_6_33_groupi_n_2570, csa_tree_add_6_33_groupi_n_2571, csa_tree_add_6_33_groupi_n_2572, csa_tree_add_6_33_groupi_n_2573, csa_tree_add_6_33_groupi_n_2574, csa_tree_add_6_33_groupi_n_2575, csa_tree_add_6_33_groupi_n_2576;
  wire csa_tree_add_6_33_groupi_n_2577, csa_tree_add_6_33_groupi_n_2578, csa_tree_add_6_33_groupi_n_2579, csa_tree_add_6_33_groupi_n_2580, csa_tree_add_6_33_groupi_n_2581, csa_tree_add_6_33_groupi_n_2582, csa_tree_add_6_33_groupi_n_2583, csa_tree_add_6_33_groupi_n_2584;
  wire csa_tree_add_6_33_groupi_n_2585, csa_tree_add_6_33_groupi_n_2586, csa_tree_add_6_33_groupi_n_2588, csa_tree_add_6_33_groupi_n_2589, csa_tree_add_6_33_groupi_n_2590, csa_tree_add_6_33_groupi_n_2591, csa_tree_add_6_33_groupi_n_2592, csa_tree_add_6_33_groupi_n_2593;
  wire csa_tree_add_6_33_groupi_n_2594, csa_tree_add_6_33_groupi_n_2595, csa_tree_add_6_33_groupi_n_2596, csa_tree_add_6_33_groupi_n_2597, csa_tree_add_6_33_groupi_n_2598, csa_tree_add_6_33_groupi_n_2599, csa_tree_add_6_33_groupi_n_2600, csa_tree_add_6_33_groupi_n_2601;
  wire csa_tree_add_6_33_groupi_n_2602, csa_tree_add_6_33_groupi_n_2603, csa_tree_add_6_33_groupi_n_2604, csa_tree_add_6_33_groupi_n_2605, csa_tree_add_6_33_groupi_n_2606, csa_tree_add_6_33_groupi_n_2607, csa_tree_add_6_33_groupi_n_2608, csa_tree_add_6_33_groupi_n_2609;
  wire csa_tree_add_6_33_groupi_n_2610, csa_tree_add_6_33_groupi_n_2611, csa_tree_add_6_33_groupi_n_2612, csa_tree_add_6_33_groupi_n_2613, csa_tree_add_6_33_groupi_n_2614, csa_tree_add_6_33_groupi_n_2615, csa_tree_add_6_33_groupi_n_2616, csa_tree_add_6_33_groupi_n_2617;
  wire csa_tree_add_6_33_groupi_n_2618, csa_tree_add_6_33_groupi_n_2619, csa_tree_add_6_33_groupi_n_2620, csa_tree_add_6_33_groupi_n_2621, csa_tree_add_6_33_groupi_n_2622, csa_tree_add_6_33_groupi_n_2623, csa_tree_add_6_33_groupi_n_2624, csa_tree_add_6_33_groupi_n_2625;
  wire csa_tree_add_6_33_groupi_n_2626, csa_tree_add_6_33_groupi_n_2627, csa_tree_add_6_33_groupi_n_2628, csa_tree_add_6_33_groupi_n_2629, csa_tree_add_6_33_groupi_n_2630, csa_tree_add_6_33_groupi_n_2631, csa_tree_add_6_33_groupi_n_2632, csa_tree_add_6_33_groupi_n_2633;
  wire csa_tree_add_6_33_groupi_n_2634, csa_tree_add_6_33_groupi_n_2635, csa_tree_add_6_33_groupi_n_2636, csa_tree_add_6_33_groupi_n_2637, csa_tree_add_6_33_groupi_n_2638, csa_tree_add_6_33_groupi_n_2639, csa_tree_add_6_33_groupi_n_2640, csa_tree_add_6_33_groupi_n_2641;
  wire csa_tree_add_6_33_groupi_n_2642, csa_tree_add_6_33_groupi_n_2643, csa_tree_add_6_33_groupi_n_2644, csa_tree_add_6_33_groupi_n_2645, csa_tree_add_6_33_groupi_n_2646, csa_tree_add_6_33_groupi_n_2647, csa_tree_add_6_33_groupi_n_2648, csa_tree_add_6_33_groupi_n_2649;
  wire csa_tree_add_6_33_groupi_n_2650, csa_tree_add_6_33_groupi_n_2651, csa_tree_add_6_33_groupi_n_2652, csa_tree_add_6_33_groupi_n_2653, csa_tree_add_6_33_groupi_n_2654, csa_tree_add_6_33_groupi_n_2655, csa_tree_add_6_33_groupi_n_2656, csa_tree_add_6_33_groupi_n_2657;
  wire csa_tree_add_6_33_groupi_n_2658, csa_tree_add_6_33_groupi_n_2659, csa_tree_add_6_33_groupi_n_2660, csa_tree_add_6_33_groupi_n_2661, csa_tree_add_6_33_groupi_n_2662, csa_tree_add_6_33_groupi_n_2663, csa_tree_add_6_33_groupi_n_2664, csa_tree_add_6_33_groupi_n_2665;
  wire csa_tree_add_6_33_groupi_n_2666, csa_tree_add_6_33_groupi_n_2667, csa_tree_add_6_33_groupi_n_2668, csa_tree_add_6_33_groupi_n_2669, csa_tree_add_6_33_groupi_n_2670, csa_tree_add_6_33_groupi_n_2671, csa_tree_add_6_33_groupi_n_2672, csa_tree_add_6_33_groupi_n_2673;
  wire csa_tree_add_6_33_groupi_n_2674, csa_tree_add_6_33_groupi_n_2675, csa_tree_add_6_33_groupi_n_2676, csa_tree_add_6_33_groupi_n_2677, csa_tree_add_6_33_groupi_n_2678, csa_tree_add_6_33_groupi_n_2679, csa_tree_add_6_33_groupi_n_2680, csa_tree_add_6_33_groupi_n_2681;
  wire csa_tree_add_6_33_groupi_n_2682, csa_tree_add_6_33_groupi_n_2683, csa_tree_add_6_33_groupi_n_2684, csa_tree_add_6_33_groupi_n_2685, csa_tree_add_6_33_groupi_n_2686, csa_tree_add_6_33_groupi_n_2687, csa_tree_add_6_33_groupi_n_2688, csa_tree_add_6_33_groupi_n_2689;
  wire csa_tree_add_6_33_groupi_n_2690, csa_tree_add_6_33_groupi_n_2691, csa_tree_add_6_33_groupi_n_2692, csa_tree_add_6_33_groupi_n_2693, csa_tree_add_6_33_groupi_n_2694, csa_tree_add_6_33_groupi_n_2695, csa_tree_add_6_33_groupi_n_2696, csa_tree_add_6_33_groupi_n_2697;
  wire csa_tree_add_6_33_groupi_n_2698, csa_tree_add_6_33_groupi_n_2699, csa_tree_add_6_33_groupi_n_2700, csa_tree_add_6_33_groupi_n_2701, csa_tree_add_6_33_groupi_n_2702, csa_tree_add_6_33_groupi_n_2703, csa_tree_add_6_33_groupi_n_2704, csa_tree_add_6_33_groupi_n_2705;
  wire csa_tree_add_6_33_groupi_n_2706, csa_tree_add_6_33_groupi_n_2707, csa_tree_add_6_33_groupi_n_2708, csa_tree_add_6_33_groupi_n_2709, csa_tree_add_6_33_groupi_n_2710, csa_tree_add_6_33_groupi_n_2711, csa_tree_add_6_33_groupi_n_2712, csa_tree_add_6_33_groupi_n_2713;
  wire csa_tree_add_6_33_groupi_n_2714, csa_tree_add_6_33_groupi_n_2715, csa_tree_add_6_33_groupi_n_2716, csa_tree_add_6_33_groupi_n_2717, csa_tree_add_6_33_groupi_n_2718, csa_tree_add_6_33_groupi_n_2719, csa_tree_add_6_33_groupi_n_2720, csa_tree_add_6_33_groupi_n_2721;
  wire csa_tree_add_6_33_groupi_n_2722, csa_tree_add_6_33_groupi_n_2723, csa_tree_add_6_33_groupi_n_2724, csa_tree_add_6_33_groupi_n_2725, csa_tree_add_6_33_groupi_n_2726, csa_tree_add_6_33_groupi_n_2727, csa_tree_add_6_33_groupi_n_2728, csa_tree_add_6_33_groupi_n_2729;
  wire csa_tree_add_6_33_groupi_n_2730, csa_tree_add_6_33_groupi_n_2731, csa_tree_add_6_33_groupi_n_2732, csa_tree_add_6_33_groupi_n_2733, csa_tree_add_6_33_groupi_n_2734, csa_tree_add_6_33_groupi_n_2735, csa_tree_add_6_33_groupi_n_2736, csa_tree_add_6_33_groupi_n_2737;
  wire csa_tree_add_6_33_groupi_n_2738, csa_tree_add_6_33_groupi_n_2739, csa_tree_add_6_33_groupi_n_2740, csa_tree_add_6_33_groupi_n_2741, csa_tree_add_6_33_groupi_n_2742, csa_tree_add_6_33_groupi_n_2743, csa_tree_add_6_33_groupi_n_2744, csa_tree_add_6_33_groupi_n_2745;
  wire csa_tree_add_6_33_groupi_n_2746, csa_tree_add_6_33_groupi_n_2747, csa_tree_add_6_33_groupi_n_2748, csa_tree_add_6_33_groupi_n_2749, csa_tree_add_6_33_groupi_n_2750, csa_tree_add_6_33_groupi_n_2751, csa_tree_add_6_33_groupi_n_2752, csa_tree_add_6_33_groupi_n_2753;
  wire csa_tree_add_6_33_groupi_n_2754, csa_tree_add_6_33_groupi_n_2755, csa_tree_add_6_33_groupi_n_2756, csa_tree_add_6_33_groupi_n_2757, csa_tree_add_6_33_groupi_n_2758, csa_tree_add_6_33_groupi_n_2759, csa_tree_add_6_33_groupi_n_2760, csa_tree_add_6_33_groupi_n_2761;
  wire csa_tree_add_6_33_groupi_n_2762, csa_tree_add_6_33_groupi_n_2763, csa_tree_add_6_33_groupi_n_2764, csa_tree_add_6_33_groupi_n_2765, csa_tree_add_6_33_groupi_n_2766, csa_tree_add_6_33_groupi_n_2767, csa_tree_add_6_33_groupi_n_2768, csa_tree_add_6_33_groupi_n_2769;
  wire csa_tree_add_6_33_groupi_n_2770, csa_tree_add_6_33_groupi_n_2771, csa_tree_add_6_33_groupi_n_2772, csa_tree_add_6_33_groupi_n_2773, csa_tree_add_6_33_groupi_n_2774, csa_tree_add_6_33_groupi_n_2775, csa_tree_add_6_33_groupi_n_2776, csa_tree_add_6_33_groupi_n_2777;
  wire csa_tree_add_6_33_groupi_n_2778, csa_tree_add_6_33_groupi_n_2779, csa_tree_add_6_33_groupi_n_2780, csa_tree_add_6_33_groupi_n_2781, csa_tree_add_6_33_groupi_n_2782, csa_tree_add_6_33_groupi_n_2783, csa_tree_add_6_33_groupi_n_2784, csa_tree_add_6_33_groupi_n_2785;
  wire csa_tree_add_6_33_groupi_n_2786, csa_tree_add_6_33_groupi_n_2787, csa_tree_add_6_33_groupi_n_2788, csa_tree_add_6_33_groupi_n_2789, csa_tree_add_6_33_groupi_n_2790, csa_tree_add_6_33_groupi_n_2791, csa_tree_add_6_33_groupi_n_2792, csa_tree_add_6_33_groupi_n_2793;
  wire csa_tree_add_6_33_groupi_n_2794, csa_tree_add_6_33_groupi_n_2795, csa_tree_add_6_33_groupi_n_2796, csa_tree_add_6_33_groupi_n_2797, csa_tree_add_6_33_groupi_n_2798, csa_tree_add_6_33_groupi_n_2799, csa_tree_add_6_33_groupi_n_2800, csa_tree_add_6_33_groupi_n_2801;
  wire csa_tree_add_6_33_groupi_n_2802, csa_tree_add_6_33_groupi_n_2803, csa_tree_add_6_33_groupi_n_2804, csa_tree_add_6_33_groupi_n_2805, csa_tree_add_6_33_groupi_n_2806, csa_tree_add_6_33_groupi_n_2807, csa_tree_add_6_33_groupi_n_2808, csa_tree_add_6_33_groupi_n_2809;
  wire csa_tree_add_6_33_groupi_n_2810, csa_tree_add_6_33_groupi_n_2811, csa_tree_add_6_33_groupi_n_2812, csa_tree_add_6_33_groupi_n_2813, csa_tree_add_6_33_groupi_n_2814, csa_tree_add_6_33_groupi_n_2815, csa_tree_add_6_33_groupi_n_2816, csa_tree_add_6_33_groupi_n_2817;
  wire csa_tree_add_6_33_groupi_n_2818, csa_tree_add_6_33_groupi_n_2819, csa_tree_add_6_33_groupi_n_2820, csa_tree_add_6_33_groupi_n_2821, csa_tree_add_6_33_groupi_n_2822, csa_tree_add_6_33_groupi_n_2823, csa_tree_add_6_33_groupi_n_2824, csa_tree_add_6_33_groupi_n_2825;
  wire csa_tree_add_6_33_groupi_n_2826, csa_tree_add_6_33_groupi_n_2827, csa_tree_add_6_33_groupi_n_2828, csa_tree_add_6_33_groupi_n_2829, csa_tree_add_6_33_groupi_n_2830, csa_tree_add_6_33_groupi_n_2831, csa_tree_add_6_33_groupi_n_2832, csa_tree_add_6_33_groupi_n_2833;
  wire csa_tree_add_6_33_groupi_n_2834, csa_tree_add_6_33_groupi_n_2835, csa_tree_add_6_33_groupi_n_2836, csa_tree_add_6_33_groupi_n_2837, csa_tree_add_6_33_groupi_n_2838, csa_tree_add_6_33_groupi_n_2839, csa_tree_add_6_33_groupi_n_2840, csa_tree_add_6_33_groupi_n_2841;
  wire csa_tree_add_6_33_groupi_n_2842, csa_tree_add_6_33_groupi_n_2843, csa_tree_add_6_33_groupi_n_2844, csa_tree_add_6_33_groupi_n_2845, csa_tree_add_6_33_groupi_n_2846, csa_tree_add_6_33_groupi_n_2847, csa_tree_add_6_33_groupi_n_2848, csa_tree_add_6_33_groupi_n_2849;
  wire csa_tree_add_6_33_groupi_n_2850, csa_tree_add_6_33_groupi_n_2851, csa_tree_add_6_33_groupi_n_2852, csa_tree_add_6_33_groupi_n_2853, csa_tree_add_6_33_groupi_n_2854, csa_tree_add_6_33_groupi_n_2855, csa_tree_add_6_33_groupi_n_2856, csa_tree_add_6_33_groupi_n_2857;
  wire csa_tree_add_6_33_groupi_n_2858, csa_tree_add_6_33_groupi_n_2859, csa_tree_add_6_33_groupi_n_2860, csa_tree_add_6_33_groupi_n_2861, csa_tree_add_6_33_groupi_n_2862, csa_tree_add_6_33_groupi_n_2863, csa_tree_add_6_33_groupi_n_2864, csa_tree_add_6_33_groupi_n_2865;
  wire csa_tree_add_6_33_groupi_n_2866, csa_tree_add_6_33_groupi_n_2867, csa_tree_add_6_33_groupi_n_2868, csa_tree_add_6_33_groupi_n_2869, csa_tree_add_6_33_groupi_n_2870, csa_tree_add_6_33_groupi_n_2871, csa_tree_add_6_33_groupi_n_2872, csa_tree_add_6_33_groupi_n_2873;
  wire csa_tree_add_6_33_groupi_n_2874, csa_tree_add_6_33_groupi_n_2875, csa_tree_add_6_33_groupi_n_2876, csa_tree_add_6_33_groupi_n_2877, csa_tree_add_6_33_groupi_n_2878, csa_tree_add_6_33_groupi_n_2879, csa_tree_add_6_33_groupi_n_2880, csa_tree_add_6_33_groupi_n_2881;
  wire csa_tree_add_6_33_groupi_n_2882, csa_tree_add_6_33_groupi_n_2883, csa_tree_add_6_33_groupi_n_2884, csa_tree_add_6_33_groupi_n_2885, csa_tree_add_6_33_groupi_n_2886, csa_tree_add_6_33_groupi_n_2887, csa_tree_add_6_33_groupi_n_2888, csa_tree_add_6_33_groupi_n_2889;
  wire csa_tree_add_6_33_groupi_n_2890, csa_tree_add_6_33_groupi_n_2891, csa_tree_add_6_33_groupi_n_2892, csa_tree_add_6_33_groupi_n_2893, csa_tree_add_6_33_groupi_n_2894, csa_tree_add_6_33_groupi_n_2895, csa_tree_add_6_33_groupi_n_2896, csa_tree_add_6_33_groupi_n_2897;
  wire csa_tree_add_6_33_groupi_n_2898, csa_tree_add_6_33_groupi_n_2899, csa_tree_add_6_33_groupi_n_2900, csa_tree_add_6_33_groupi_n_2901, csa_tree_add_6_33_groupi_n_2902, csa_tree_add_6_33_groupi_n_2903, csa_tree_add_6_33_groupi_n_2904, csa_tree_add_6_33_groupi_n_2905;
  wire csa_tree_add_6_33_groupi_n_2906, csa_tree_add_6_33_groupi_n_2907, csa_tree_add_6_33_groupi_n_2908, csa_tree_add_6_33_groupi_n_2909, csa_tree_add_6_33_groupi_n_2910, csa_tree_add_6_33_groupi_n_2911, csa_tree_add_6_33_groupi_n_2912, csa_tree_add_6_33_groupi_n_2913;
  wire csa_tree_add_6_33_groupi_n_2914, csa_tree_add_6_33_groupi_n_2915, csa_tree_add_6_33_groupi_n_2916, csa_tree_add_6_33_groupi_n_2917, csa_tree_add_6_33_groupi_n_2918, csa_tree_add_6_33_groupi_n_2919, csa_tree_add_6_33_groupi_n_2920, csa_tree_add_6_33_groupi_n_2921;
  wire csa_tree_add_6_33_groupi_n_2922, csa_tree_add_6_33_groupi_n_2923, csa_tree_add_6_33_groupi_n_2924, csa_tree_add_6_33_groupi_n_2925, csa_tree_add_6_33_groupi_n_2926, csa_tree_add_6_33_groupi_n_2927, csa_tree_add_6_33_groupi_n_2928, csa_tree_add_6_33_groupi_n_2929;
  wire csa_tree_add_6_33_groupi_n_2930, csa_tree_add_6_33_groupi_n_2931, csa_tree_add_6_33_groupi_n_2932, csa_tree_add_6_33_groupi_n_2933, csa_tree_add_6_33_groupi_n_2934, csa_tree_add_6_33_groupi_n_2935, csa_tree_add_6_33_groupi_n_2936, csa_tree_add_6_33_groupi_n_2937;
  wire csa_tree_add_6_33_groupi_n_2938, csa_tree_add_6_33_groupi_n_2939, csa_tree_add_6_33_groupi_n_2940, csa_tree_add_6_33_groupi_n_2941, csa_tree_add_6_33_groupi_n_2942, csa_tree_add_6_33_groupi_n_2943, csa_tree_add_6_33_groupi_n_2944, csa_tree_add_6_33_groupi_n_2945;
  wire csa_tree_add_6_33_groupi_n_2946, csa_tree_add_6_33_groupi_n_2947, csa_tree_add_6_33_groupi_n_2948, csa_tree_add_6_33_groupi_n_2949, csa_tree_add_6_33_groupi_n_2950, csa_tree_add_6_33_groupi_n_2951, csa_tree_add_6_33_groupi_n_2952, csa_tree_add_6_33_groupi_n_2953;
  wire csa_tree_add_6_33_groupi_n_2954, csa_tree_add_6_33_groupi_n_2955, csa_tree_add_6_33_groupi_n_2956, csa_tree_add_6_33_groupi_n_2957, csa_tree_add_6_33_groupi_n_2958, csa_tree_add_6_33_groupi_n_2959, csa_tree_add_6_33_groupi_n_2960, csa_tree_add_6_33_groupi_n_2961;
  wire csa_tree_add_6_33_groupi_n_2962, csa_tree_add_6_33_groupi_n_2963, csa_tree_add_6_33_groupi_n_2964, csa_tree_add_6_33_groupi_n_2965, csa_tree_add_6_33_groupi_n_2966, csa_tree_add_6_33_groupi_n_2967, csa_tree_add_6_33_groupi_n_2968, csa_tree_add_6_33_groupi_n_2969;
  wire csa_tree_add_6_33_groupi_n_2970, csa_tree_add_6_33_groupi_n_2971, csa_tree_add_6_33_groupi_n_2972, csa_tree_add_6_33_groupi_n_2973, csa_tree_add_6_33_groupi_n_2974, csa_tree_add_6_33_groupi_n_2975, csa_tree_add_6_33_groupi_n_2976, csa_tree_add_6_33_groupi_n_2977;
  wire csa_tree_add_6_33_groupi_n_2978, csa_tree_add_6_33_groupi_n_2979, csa_tree_add_6_33_groupi_n_2980, csa_tree_add_6_33_groupi_n_2981, csa_tree_add_6_33_groupi_n_2982, csa_tree_add_6_33_groupi_n_2983, csa_tree_add_6_33_groupi_n_2984, csa_tree_add_6_33_groupi_n_2985;
  wire csa_tree_add_6_33_groupi_n_2986, csa_tree_add_6_33_groupi_n_2987, csa_tree_add_6_33_groupi_n_2988, csa_tree_add_6_33_groupi_n_2989, csa_tree_add_6_33_groupi_n_2990, csa_tree_add_6_33_groupi_n_2991, csa_tree_add_6_33_groupi_n_2992, csa_tree_add_6_33_groupi_n_2993;
  wire csa_tree_add_6_33_groupi_n_2994, csa_tree_add_6_33_groupi_n_2995, csa_tree_add_6_33_groupi_n_2996, csa_tree_add_6_33_groupi_n_2997, csa_tree_add_6_33_groupi_n_2998, csa_tree_add_6_33_groupi_n_2999, csa_tree_add_6_33_groupi_n_3000, csa_tree_add_6_33_groupi_n_3001;
  wire csa_tree_add_6_33_groupi_n_3002, csa_tree_add_6_33_groupi_n_3003, csa_tree_add_6_33_groupi_n_3004, csa_tree_add_6_33_groupi_n_3005, csa_tree_add_6_33_groupi_n_3006, csa_tree_add_6_33_groupi_n_3007, csa_tree_add_6_33_groupi_n_3008, csa_tree_add_6_33_groupi_n_3009;
  wire csa_tree_add_6_33_groupi_n_3010, csa_tree_add_6_33_groupi_n_3011, csa_tree_add_6_33_groupi_n_3012, csa_tree_add_6_33_groupi_n_3013, csa_tree_add_6_33_groupi_n_3014, csa_tree_add_6_33_groupi_n_3015, csa_tree_add_6_33_groupi_n_3016, csa_tree_add_6_33_groupi_n_3017;
  wire csa_tree_add_6_33_groupi_n_3018, csa_tree_add_6_33_groupi_n_3019, csa_tree_add_6_33_groupi_n_3020, csa_tree_add_6_33_groupi_n_3021, csa_tree_add_6_33_groupi_n_3022, csa_tree_add_6_33_groupi_n_3023, csa_tree_add_6_33_groupi_n_3024, csa_tree_add_6_33_groupi_n_3025;
  wire csa_tree_add_6_33_groupi_n_3026, csa_tree_add_6_33_groupi_n_3027, csa_tree_add_6_33_groupi_n_3028, csa_tree_add_6_33_groupi_n_3029, csa_tree_add_6_33_groupi_n_3030, csa_tree_add_6_33_groupi_n_3031, csa_tree_add_6_33_groupi_n_3032, csa_tree_add_6_33_groupi_n_3033;
  wire csa_tree_add_6_33_groupi_n_3034, csa_tree_add_6_33_groupi_n_3035, csa_tree_add_6_33_groupi_n_3036, csa_tree_add_6_33_groupi_n_3037, csa_tree_add_6_33_groupi_n_3038, csa_tree_add_6_33_groupi_n_3039, csa_tree_add_6_33_groupi_n_3040, csa_tree_add_6_33_groupi_n_3041;
  wire csa_tree_add_6_33_groupi_n_3042, csa_tree_add_6_33_groupi_n_3043, csa_tree_add_6_33_groupi_n_3044, csa_tree_add_6_33_groupi_n_3045, csa_tree_add_6_33_groupi_n_3046, csa_tree_add_6_33_groupi_n_3047, csa_tree_add_6_33_groupi_n_3048, csa_tree_add_6_33_groupi_n_3049;
  wire csa_tree_add_6_33_groupi_n_3050, csa_tree_add_6_33_groupi_n_3051, csa_tree_add_6_33_groupi_n_3052, csa_tree_add_6_33_groupi_n_3053, csa_tree_add_6_33_groupi_n_3054, csa_tree_add_6_33_groupi_n_3055, csa_tree_add_6_33_groupi_n_3056, csa_tree_add_6_33_groupi_n_3057;
  wire csa_tree_add_6_33_groupi_n_3058, csa_tree_add_6_33_groupi_n_3059, csa_tree_add_6_33_groupi_n_3060, csa_tree_add_6_33_groupi_n_3061, csa_tree_add_6_33_groupi_n_3062, csa_tree_add_6_33_groupi_n_3063, csa_tree_add_6_33_groupi_n_3064, csa_tree_add_6_33_groupi_n_3065;
  wire csa_tree_add_6_33_groupi_n_3066, csa_tree_add_6_33_groupi_n_3067, csa_tree_add_6_33_groupi_n_3068, csa_tree_add_6_33_groupi_n_3069, csa_tree_add_6_33_groupi_n_3070, csa_tree_add_6_33_groupi_n_3071, csa_tree_add_6_33_groupi_n_3072, csa_tree_add_6_33_groupi_n_3073;
  wire csa_tree_add_6_33_groupi_n_3074, csa_tree_add_6_33_groupi_n_3075, csa_tree_add_6_33_groupi_n_3076, csa_tree_add_6_33_groupi_n_3077, csa_tree_add_6_33_groupi_n_3078, csa_tree_add_6_33_groupi_n_3079, csa_tree_add_6_33_groupi_n_3080, csa_tree_add_6_33_groupi_n_3081;
  wire csa_tree_add_6_33_groupi_n_3082, csa_tree_add_6_33_groupi_n_3083, csa_tree_add_6_33_groupi_n_3084, csa_tree_add_6_33_groupi_n_3085, csa_tree_add_6_33_groupi_n_3086, csa_tree_add_6_33_groupi_n_3087, csa_tree_add_6_33_groupi_n_3088, csa_tree_add_6_33_groupi_n_3089;
  wire csa_tree_add_6_33_groupi_n_3090, csa_tree_add_6_33_groupi_n_3091, csa_tree_add_6_33_groupi_n_3092, csa_tree_add_6_33_groupi_n_3093, csa_tree_add_6_33_groupi_n_3094, csa_tree_add_6_33_groupi_n_3095, csa_tree_add_6_33_groupi_n_3096, csa_tree_add_6_33_groupi_n_3097;
  wire csa_tree_add_6_33_groupi_n_3098, csa_tree_add_6_33_groupi_n_3099, csa_tree_add_6_33_groupi_n_3100, csa_tree_add_6_33_groupi_n_3101, csa_tree_add_6_33_groupi_n_3102, csa_tree_add_6_33_groupi_n_3103, csa_tree_add_6_33_groupi_n_3104, csa_tree_add_6_33_groupi_n_3105;
  wire csa_tree_add_6_33_groupi_n_3106, csa_tree_add_6_33_groupi_n_3107, csa_tree_add_6_33_groupi_n_3108, csa_tree_add_6_33_groupi_n_3109, csa_tree_add_6_33_groupi_n_3110, csa_tree_add_6_33_groupi_n_3111, csa_tree_add_6_33_groupi_n_3112, csa_tree_add_6_33_groupi_n_3113;
  wire csa_tree_add_6_33_groupi_n_3114, csa_tree_add_6_33_groupi_n_3115, csa_tree_add_6_33_groupi_n_3116, csa_tree_add_6_33_groupi_n_3117, csa_tree_add_6_33_groupi_n_3118, csa_tree_add_6_33_groupi_n_3119, csa_tree_add_6_33_groupi_n_3120, csa_tree_add_6_33_groupi_n_3121;
  wire csa_tree_add_6_33_groupi_n_3122, csa_tree_add_6_33_groupi_n_3123, csa_tree_add_6_33_groupi_n_3124, csa_tree_add_6_33_groupi_n_3125, csa_tree_add_6_33_groupi_n_3126, csa_tree_add_6_33_groupi_n_3127, csa_tree_add_6_33_groupi_n_3128, csa_tree_add_6_33_groupi_n_3129;
  wire csa_tree_add_6_33_groupi_n_3130, csa_tree_add_6_33_groupi_n_3131, csa_tree_add_6_33_groupi_n_3132, csa_tree_add_6_33_groupi_n_3133, csa_tree_add_6_33_groupi_n_3134, csa_tree_add_6_33_groupi_n_3135, csa_tree_add_6_33_groupi_n_3136, csa_tree_add_6_33_groupi_n_3137;
  wire csa_tree_add_6_33_groupi_n_3138, csa_tree_add_6_33_groupi_n_3139, csa_tree_add_6_33_groupi_n_3140, csa_tree_add_6_33_groupi_n_3141, csa_tree_add_6_33_groupi_n_3142, csa_tree_add_6_33_groupi_n_3143, csa_tree_add_6_33_groupi_n_3144, csa_tree_add_6_33_groupi_n_3145;
  wire csa_tree_add_6_33_groupi_n_3146, csa_tree_add_6_33_groupi_n_3147, csa_tree_add_6_33_groupi_n_3148, csa_tree_add_6_33_groupi_n_3149, csa_tree_add_6_33_groupi_n_3150, csa_tree_add_6_33_groupi_n_3151, csa_tree_add_6_33_groupi_n_3152, csa_tree_add_6_33_groupi_n_3153;
  wire csa_tree_add_6_33_groupi_n_3154, csa_tree_add_6_33_groupi_n_3155, csa_tree_add_6_33_groupi_n_3156, csa_tree_add_6_33_groupi_n_3157, csa_tree_add_6_33_groupi_n_3158, csa_tree_add_6_33_groupi_n_3159, csa_tree_add_6_33_groupi_n_3160, csa_tree_add_6_33_groupi_n_3161;
  wire csa_tree_add_6_33_groupi_n_3162, csa_tree_add_6_33_groupi_n_3163, csa_tree_add_6_33_groupi_n_3164, csa_tree_add_6_33_groupi_n_3165, csa_tree_add_6_33_groupi_n_3166, csa_tree_add_6_33_groupi_n_3167, csa_tree_add_6_33_groupi_n_3168, csa_tree_add_6_33_groupi_n_3169;
  wire csa_tree_add_6_33_groupi_n_3170, csa_tree_add_6_33_groupi_n_3171, csa_tree_add_6_33_groupi_n_3172, csa_tree_add_6_33_groupi_n_3173, csa_tree_add_6_33_groupi_n_3174, csa_tree_add_6_33_groupi_n_3175, csa_tree_add_6_33_groupi_n_3176, csa_tree_add_6_33_groupi_n_3177;
  wire csa_tree_add_6_33_groupi_n_3178, csa_tree_add_6_33_groupi_n_3179, csa_tree_add_6_33_groupi_n_3180, csa_tree_add_6_33_groupi_n_3181, csa_tree_add_6_33_groupi_n_3182, csa_tree_add_6_33_groupi_n_3183, csa_tree_add_6_33_groupi_n_3184, csa_tree_add_6_33_groupi_n_3185;
  wire csa_tree_add_6_33_groupi_n_3186, csa_tree_add_6_33_groupi_n_3187, csa_tree_add_6_33_groupi_n_3188, csa_tree_add_6_33_groupi_n_3189, csa_tree_add_6_33_groupi_n_3190, csa_tree_add_6_33_groupi_n_3191, csa_tree_add_6_33_groupi_n_3192, csa_tree_add_6_33_groupi_n_3193;
  wire csa_tree_add_6_33_groupi_n_3194, csa_tree_add_6_33_groupi_n_3195, csa_tree_add_6_33_groupi_n_3196, csa_tree_add_6_33_groupi_n_3197, csa_tree_add_6_33_groupi_n_3198, csa_tree_add_6_33_groupi_n_3199, csa_tree_add_6_33_groupi_n_3200, csa_tree_add_6_33_groupi_n_3201;
  wire csa_tree_add_6_33_groupi_n_3202, csa_tree_add_6_33_groupi_n_3203, csa_tree_add_6_33_groupi_n_3204, csa_tree_add_6_33_groupi_n_3205, csa_tree_add_6_33_groupi_n_3206, csa_tree_add_6_33_groupi_n_3207, csa_tree_add_6_33_groupi_n_3208, csa_tree_add_6_33_groupi_n_3209;
  wire csa_tree_add_6_33_groupi_n_3210, csa_tree_add_6_33_groupi_n_3211, csa_tree_add_6_33_groupi_n_3212, csa_tree_add_6_33_groupi_n_3213, csa_tree_add_6_33_groupi_n_3214, csa_tree_add_6_33_groupi_n_3215, csa_tree_add_6_33_groupi_n_3216, csa_tree_add_6_33_groupi_n_3217;
  wire csa_tree_add_6_33_groupi_n_3218, csa_tree_add_6_33_groupi_n_3219, csa_tree_add_6_33_groupi_n_3220, csa_tree_add_6_33_groupi_n_3221, csa_tree_add_6_33_groupi_n_3222, csa_tree_add_6_33_groupi_n_3223, csa_tree_add_6_33_groupi_n_3224, csa_tree_add_6_33_groupi_n_3225;
  wire csa_tree_add_6_33_groupi_n_3226, csa_tree_add_6_33_groupi_n_3227, csa_tree_add_6_33_groupi_n_3228, csa_tree_add_6_33_groupi_n_3229, csa_tree_add_6_33_groupi_n_3230, csa_tree_add_6_33_groupi_n_3231, csa_tree_add_6_33_groupi_n_3232, csa_tree_add_6_33_groupi_n_3233;
  wire csa_tree_add_6_33_groupi_n_3234, csa_tree_add_6_33_groupi_n_3235, csa_tree_add_6_33_groupi_n_3236, csa_tree_add_6_33_groupi_n_3237, csa_tree_add_6_33_groupi_n_3238, csa_tree_add_6_33_groupi_n_3239, csa_tree_add_6_33_groupi_n_3240, csa_tree_add_6_33_groupi_n_3241;
  wire csa_tree_add_6_33_groupi_n_3242, csa_tree_add_6_33_groupi_n_3243, csa_tree_add_6_33_groupi_n_3244, csa_tree_add_6_33_groupi_n_3245, csa_tree_add_6_33_groupi_n_3246, csa_tree_add_6_33_groupi_n_3247, csa_tree_add_6_33_groupi_n_3248, csa_tree_add_6_33_groupi_n_3249;
  wire csa_tree_add_6_33_groupi_n_3250, csa_tree_add_6_33_groupi_n_3251, csa_tree_add_6_33_groupi_n_3252, csa_tree_add_6_33_groupi_n_3253, csa_tree_add_6_33_groupi_n_3254, csa_tree_add_6_33_groupi_n_3255, csa_tree_add_6_33_groupi_n_3256, csa_tree_add_6_33_groupi_n_3257;
  wire csa_tree_add_6_33_groupi_n_3258, csa_tree_add_6_33_groupi_n_3259, csa_tree_add_6_33_groupi_n_3260, csa_tree_add_6_33_groupi_n_3261, csa_tree_add_6_33_groupi_n_3262, csa_tree_add_6_33_groupi_n_3263, csa_tree_add_6_33_groupi_n_3264, csa_tree_add_6_33_groupi_n_3265;
  wire csa_tree_add_6_33_groupi_n_3266, csa_tree_add_6_33_groupi_n_3267, csa_tree_add_6_33_groupi_n_3268, csa_tree_add_6_33_groupi_n_3269, csa_tree_add_6_33_groupi_n_3270, csa_tree_add_6_33_groupi_n_3271, csa_tree_add_6_33_groupi_n_3272, csa_tree_add_6_33_groupi_n_3273;
  wire csa_tree_add_6_33_groupi_n_3274, csa_tree_add_6_33_groupi_n_3275, csa_tree_add_6_33_groupi_n_3276, csa_tree_add_6_33_groupi_n_3277, csa_tree_add_6_33_groupi_n_3278, csa_tree_add_6_33_groupi_n_3279, csa_tree_add_6_33_groupi_n_3280, csa_tree_add_6_33_groupi_n_3281;
  wire csa_tree_add_6_33_groupi_n_3282, csa_tree_add_6_33_groupi_n_3283, csa_tree_add_6_33_groupi_n_3284, csa_tree_add_6_33_groupi_n_3285, csa_tree_add_6_33_groupi_n_3286, csa_tree_add_6_33_groupi_n_3287, csa_tree_add_6_33_groupi_n_3288, csa_tree_add_6_33_groupi_n_3289;
  wire csa_tree_add_6_33_groupi_n_3290, csa_tree_add_6_33_groupi_n_3291, csa_tree_add_6_33_groupi_n_3292, csa_tree_add_6_33_groupi_n_3293, csa_tree_add_6_33_groupi_n_3294, csa_tree_add_6_33_groupi_n_3295, csa_tree_add_6_33_groupi_n_3296, csa_tree_add_6_33_groupi_n_3297;
  wire csa_tree_add_6_33_groupi_n_3298, csa_tree_add_6_33_groupi_n_3299, csa_tree_add_6_33_groupi_n_3300, csa_tree_add_6_33_groupi_n_3301, csa_tree_add_6_33_groupi_n_3302, csa_tree_add_6_33_groupi_n_3303, csa_tree_add_6_33_groupi_n_3304, csa_tree_add_6_33_groupi_n_3305;
  wire csa_tree_add_6_33_groupi_n_3306, csa_tree_add_6_33_groupi_n_3307, csa_tree_add_6_33_groupi_n_3308, csa_tree_add_6_33_groupi_n_3309, csa_tree_add_6_33_groupi_n_3310, csa_tree_add_6_33_groupi_n_3311, csa_tree_add_6_33_groupi_n_3312, csa_tree_add_6_33_groupi_n_3313;
  wire csa_tree_add_6_33_groupi_n_3314, csa_tree_add_6_33_groupi_n_3315, csa_tree_add_6_33_groupi_n_3316, csa_tree_add_6_33_groupi_n_3317, csa_tree_add_6_33_groupi_n_3318, csa_tree_add_6_33_groupi_n_3319, csa_tree_add_6_33_groupi_n_3320, csa_tree_add_6_33_groupi_n_3321;
  wire csa_tree_add_6_33_groupi_n_3322, csa_tree_add_6_33_groupi_n_3323, csa_tree_add_6_33_groupi_n_3324, csa_tree_add_6_33_groupi_n_3325, csa_tree_add_6_33_groupi_n_3326, csa_tree_add_6_33_groupi_n_3327, csa_tree_add_6_33_groupi_n_3328, csa_tree_add_6_33_groupi_n_3329;
  wire csa_tree_add_6_33_groupi_n_3330, csa_tree_add_6_33_groupi_n_3331, csa_tree_add_6_33_groupi_n_3332, csa_tree_add_6_33_groupi_n_3333, csa_tree_add_6_33_groupi_n_3334, csa_tree_add_6_33_groupi_n_3335, csa_tree_add_6_33_groupi_n_3336, csa_tree_add_6_33_groupi_n_3337;
  wire csa_tree_add_6_33_groupi_n_3338, csa_tree_add_6_33_groupi_n_3339, csa_tree_add_6_33_groupi_n_3340, csa_tree_add_6_33_groupi_n_3341, csa_tree_add_6_33_groupi_n_3342, csa_tree_add_6_33_groupi_n_3343, csa_tree_add_6_33_groupi_n_3344, csa_tree_add_6_33_groupi_n_3345;
  wire csa_tree_add_6_33_groupi_n_3346, csa_tree_add_6_33_groupi_n_3347, csa_tree_add_6_33_groupi_n_3348, csa_tree_add_6_33_groupi_n_3349, csa_tree_add_6_33_groupi_n_3350, csa_tree_add_6_33_groupi_n_3351, csa_tree_add_6_33_groupi_n_3352, csa_tree_add_6_33_groupi_n_3353;
  wire csa_tree_add_6_33_groupi_n_3354, csa_tree_add_6_33_groupi_n_3355, csa_tree_add_6_33_groupi_n_3356, csa_tree_add_6_33_groupi_n_3357, csa_tree_add_6_33_groupi_n_3358, csa_tree_add_6_33_groupi_n_3359, csa_tree_add_6_33_groupi_n_3360, csa_tree_add_6_33_groupi_n_3361;
  wire csa_tree_add_6_33_groupi_n_3362, csa_tree_add_6_33_groupi_n_3363, csa_tree_add_6_33_groupi_n_3364, csa_tree_add_6_33_groupi_n_3365, csa_tree_add_6_33_groupi_n_3366, csa_tree_add_6_33_groupi_n_3367, csa_tree_add_6_33_groupi_n_3368, csa_tree_add_6_33_groupi_n_3369;
  wire csa_tree_add_6_33_groupi_n_3370, csa_tree_add_6_33_groupi_n_3371, csa_tree_add_6_33_groupi_n_3372, csa_tree_add_6_33_groupi_n_3373, csa_tree_add_6_33_groupi_n_3374, csa_tree_add_6_33_groupi_n_3375, csa_tree_add_6_33_groupi_n_3376, csa_tree_add_6_33_groupi_n_3377;
  wire csa_tree_add_6_33_groupi_n_3378, csa_tree_add_6_33_groupi_n_3379, csa_tree_add_6_33_groupi_n_3380, csa_tree_add_6_33_groupi_n_3381, csa_tree_add_6_33_groupi_n_3382, csa_tree_add_6_33_groupi_n_3383, csa_tree_add_6_33_groupi_n_3384, csa_tree_add_6_33_groupi_n_3385;
  wire csa_tree_add_6_33_groupi_n_3386, csa_tree_add_6_33_groupi_n_3387, csa_tree_add_6_33_groupi_n_3388, csa_tree_add_6_33_groupi_n_3389, csa_tree_add_6_33_groupi_n_3390, csa_tree_add_6_33_groupi_n_3391, csa_tree_add_6_33_groupi_n_3392, csa_tree_add_6_33_groupi_n_3393;
  wire csa_tree_add_6_33_groupi_n_3394, csa_tree_add_6_33_groupi_n_3395, csa_tree_add_6_33_groupi_n_3396, csa_tree_add_6_33_groupi_n_3397, csa_tree_add_6_33_groupi_n_3398, csa_tree_add_6_33_groupi_n_3399, csa_tree_add_6_33_groupi_n_3400, csa_tree_add_6_33_groupi_n_3401;
  wire csa_tree_add_6_33_groupi_n_3402, csa_tree_add_6_33_groupi_n_3403, csa_tree_add_6_33_groupi_n_3405, csa_tree_add_6_33_groupi_n_3406, csa_tree_add_6_33_groupi_n_3407, csa_tree_add_6_33_groupi_n_3408, csa_tree_add_6_33_groupi_n_3409, csa_tree_add_6_33_groupi_n_3410;
  wire csa_tree_add_6_33_groupi_n_3411, csa_tree_add_6_33_groupi_n_3412, csa_tree_add_6_33_groupi_n_3413, csa_tree_add_6_33_groupi_n_3414, csa_tree_add_6_33_groupi_n_3415, csa_tree_add_6_33_groupi_n_3416, csa_tree_add_6_33_groupi_n_3417, csa_tree_add_6_33_groupi_n_3418;
  wire csa_tree_add_6_33_groupi_n_3419, csa_tree_add_6_33_groupi_n_3420, csa_tree_add_6_33_groupi_n_3421, csa_tree_add_6_33_groupi_n_3422, csa_tree_add_6_33_groupi_n_3423, csa_tree_add_6_33_groupi_n_3424, csa_tree_add_6_33_groupi_n_3425, csa_tree_add_6_33_groupi_n_3426;
  wire csa_tree_add_6_33_groupi_n_3427, csa_tree_add_6_33_groupi_n_3428, csa_tree_add_6_33_groupi_n_3429, csa_tree_add_6_33_groupi_n_3430, csa_tree_add_6_33_groupi_n_3431, csa_tree_add_6_33_groupi_n_3432, csa_tree_add_6_33_groupi_n_3433, csa_tree_add_6_33_groupi_n_3434;
  wire csa_tree_add_6_33_groupi_n_3435, csa_tree_add_6_33_groupi_n_3436, csa_tree_add_6_33_groupi_n_3437, csa_tree_add_6_33_groupi_n_3438, csa_tree_add_6_33_groupi_n_3439, csa_tree_add_6_33_groupi_n_3440, csa_tree_add_6_33_groupi_n_3441, csa_tree_add_6_33_groupi_n_3442;
  wire csa_tree_add_6_33_groupi_n_3443, csa_tree_add_6_33_groupi_n_3444, csa_tree_add_6_33_groupi_n_3445, csa_tree_add_6_33_groupi_n_3446, csa_tree_add_6_33_groupi_n_3447, csa_tree_add_6_33_groupi_n_3448, csa_tree_add_6_33_groupi_n_3449, csa_tree_add_6_33_groupi_n_3450;
  wire csa_tree_add_6_33_groupi_n_3451, csa_tree_add_6_33_groupi_n_3452, csa_tree_add_6_33_groupi_n_3453, csa_tree_add_6_33_groupi_n_3454, csa_tree_add_6_33_groupi_n_3455, csa_tree_add_6_33_groupi_n_3456, csa_tree_add_6_33_groupi_n_3457, csa_tree_add_6_33_groupi_n_3458;
  wire csa_tree_add_6_33_groupi_n_3459, csa_tree_add_6_33_groupi_n_3460, csa_tree_add_6_33_groupi_n_3461, csa_tree_add_6_33_groupi_n_3462, csa_tree_add_6_33_groupi_n_3463, csa_tree_add_6_33_groupi_n_3464, csa_tree_add_6_33_groupi_n_3465, csa_tree_add_6_33_groupi_n_3466;
  wire csa_tree_add_6_33_groupi_n_3467, csa_tree_add_6_33_groupi_n_3468, csa_tree_add_6_33_groupi_n_3469, csa_tree_add_6_33_groupi_n_3470, csa_tree_add_6_33_groupi_n_3471, csa_tree_add_6_33_groupi_n_3472, csa_tree_add_6_33_groupi_n_3473, csa_tree_add_6_33_groupi_n_3474;
  wire csa_tree_add_6_33_groupi_n_3475, csa_tree_add_6_33_groupi_n_3476, csa_tree_add_6_33_groupi_n_3477, csa_tree_add_6_33_groupi_n_3478, csa_tree_add_6_33_groupi_n_3479, csa_tree_add_6_33_groupi_n_3480, csa_tree_add_6_33_groupi_n_3481, csa_tree_add_6_33_groupi_n_3482;
  wire csa_tree_add_6_33_groupi_n_3483, csa_tree_add_6_33_groupi_n_3484, csa_tree_add_6_33_groupi_n_3485, csa_tree_add_6_33_groupi_n_3486, csa_tree_add_6_33_groupi_n_3487, csa_tree_add_6_33_groupi_n_3488, csa_tree_add_6_33_groupi_n_3489, csa_tree_add_6_33_groupi_n_3490;
  wire csa_tree_add_6_33_groupi_n_3491, csa_tree_add_6_33_groupi_n_3492, csa_tree_add_6_33_groupi_n_3493, csa_tree_add_6_33_groupi_n_3494, csa_tree_add_6_33_groupi_n_3495, csa_tree_add_6_33_groupi_n_3496, csa_tree_add_6_33_groupi_n_3497, csa_tree_add_6_33_groupi_n_3498;
  wire csa_tree_add_6_33_groupi_n_3499, csa_tree_add_6_33_groupi_n_3500, csa_tree_add_6_33_groupi_n_3501, csa_tree_add_6_33_groupi_n_3502, csa_tree_add_6_33_groupi_n_3503, csa_tree_add_6_33_groupi_n_3504, csa_tree_add_6_33_groupi_n_3505, csa_tree_add_6_33_groupi_n_3506;
  wire csa_tree_add_6_33_groupi_n_3507, csa_tree_add_6_33_groupi_n_3508, csa_tree_add_6_33_groupi_n_3509, csa_tree_add_6_33_groupi_n_3510, csa_tree_add_6_33_groupi_n_3511, csa_tree_add_6_33_groupi_n_3512, csa_tree_add_6_33_groupi_n_3513, csa_tree_add_6_33_groupi_n_3514;
  wire csa_tree_add_6_33_groupi_n_3515, csa_tree_add_6_33_groupi_n_3516, csa_tree_add_6_33_groupi_n_3517, csa_tree_add_6_33_groupi_n_3518, csa_tree_add_6_33_groupi_n_3519, csa_tree_add_6_33_groupi_n_3520, csa_tree_add_6_33_groupi_n_3521, csa_tree_add_6_33_groupi_n_3522;
  wire csa_tree_add_6_33_groupi_n_3523, csa_tree_add_6_33_groupi_n_3524, csa_tree_add_6_33_groupi_n_3525, csa_tree_add_6_33_groupi_n_3526, csa_tree_add_6_33_groupi_n_3527, csa_tree_add_6_33_groupi_n_3528, csa_tree_add_6_33_groupi_n_3529, csa_tree_add_6_33_groupi_n_3530;
  wire csa_tree_add_6_33_groupi_n_3531, csa_tree_add_6_33_groupi_n_3532, csa_tree_add_6_33_groupi_n_3533, csa_tree_add_6_33_groupi_n_3534, csa_tree_add_6_33_groupi_n_3535, csa_tree_add_6_33_groupi_n_3536, csa_tree_add_6_33_groupi_n_3537, csa_tree_add_6_33_groupi_n_3538;
  wire csa_tree_add_6_33_groupi_n_3539, csa_tree_add_6_33_groupi_n_3540, csa_tree_add_6_33_groupi_n_3541, csa_tree_add_6_33_groupi_n_3542, csa_tree_add_6_33_groupi_n_3543, csa_tree_add_6_33_groupi_n_3544, csa_tree_add_6_33_groupi_n_3545, csa_tree_add_6_33_groupi_n_3546;
  wire csa_tree_add_6_33_groupi_n_3547, csa_tree_add_6_33_groupi_n_3548, csa_tree_add_6_33_groupi_n_3549, csa_tree_add_6_33_groupi_n_3550, csa_tree_add_6_33_groupi_n_3551, csa_tree_add_6_33_groupi_n_3552, csa_tree_add_6_33_groupi_n_3553, csa_tree_add_6_33_groupi_n_3554;
  wire csa_tree_add_6_33_groupi_n_3555, csa_tree_add_6_33_groupi_n_3556, csa_tree_add_6_33_groupi_n_3557, csa_tree_add_6_33_groupi_n_3558, csa_tree_add_6_33_groupi_n_3559, csa_tree_add_6_33_groupi_n_3560, csa_tree_add_6_33_groupi_n_3561, csa_tree_add_6_33_groupi_n_3562;
  wire csa_tree_add_6_33_groupi_n_3563, csa_tree_add_6_33_groupi_n_3564, csa_tree_add_6_33_groupi_n_3565, csa_tree_add_6_33_groupi_n_3566, csa_tree_add_6_33_groupi_n_3567, csa_tree_add_6_33_groupi_n_3568, csa_tree_add_6_33_groupi_n_3569, csa_tree_add_6_33_groupi_n_3570;
  wire csa_tree_add_6_33_groupi_n_3571, csa_tree_add_6_33_groupi_n_3572, csa_tree_add_6_33_groupi_n_3573, csa_tree_add_6_33_groupi_n_3574, csa_tree_add_6_33_groupi_n_3575, csa_tree_add_6_33_groupi_n_3576, csa_tree_add_6_33_groupi_n_3577, csa_tree_add_6_33_groupi_n_3578;
  wire csa_tree_add_6_33_groupi_n_3579, csa_tree_add_6_33_groupi_n_3580, csa_tree_add_6_33_groupi_n_3581, csa_tree_add_6_33_groupi_n_3582, csa_tree_add_6_33_groupi_n_3583, csa_tree_add_6_33_groupi_n_3584, csa_tree_add_6_33_groupi_n_3585, csa_tree_add_6_33_groupi_n_3586;
  wire csa_tree_add_6_33_groupi_n_3587, csa_tree_add_6_33_groupi_n_3588, csa_tree_add_6_33_groupi_n_3589, csa_tree_add_6_33_groupi_n_3590, csa_tree_add_6_33_groupi_n_3591, csa_tree_add_6_33_groupi_n_3592, csa_tree_add_6_33_groupi_n_3593, csa_tree_add_6_33_groupi_n_3594;
  wire csa_tree_add_6_33_groupi_n_3596, csa_tree_add_6_33_groupi_n_3597, csa_tree_add_6_33_groupi_n_3598, csa_tree_add_6_33_groupi_n_3599, csa_tree_add_6_33_groupi_n_3600, csa_tree_add_6_33_groupi_n_3601, csa_tree_add_6_33_groupi_n_3602, csa_tree_add_6_33_groupi_n_3603;
  wire csa_tree_add_6_33_groupi_n_3604, csa_tree_add_6_33_groupi_n_3605, csa_tree_add_6_33_groupi_n_3606, csa_tree_add_6_33_groupi_n_3607, csa_tree_add_6_33_groupi_n_3608, csa_tree_add_6_33_groupi_n_3609, csa_tree_add_6_33_groupi_n_3610, csa_tree_add_6_33_groupi_n_3611;
  wire csa_tree_add_6_33_groupi_n_3612, csa_tree_add_6_33_groupi_n_3613, csa_tree_add_6_33_groupi_n_3614, csa_tree_add_6_33_groupi_n_3615, csa_tree_add_6_33_groupi_n_3616, csa_tree_add_6_33_groupi_n_3617, csa_tree_add_6_33_groupi_n_3618, csa_tree_add_6_33_groupi_n_3619;
  wire csa_tree_add_6_33_groupi_n_3620, csa_tree_add_6_33_groupi_n_3621, csa_tree_add_6_33_groupi_n_3622, csa_tree_add_6_33_groupi_n_3623, csa_tree_add_6_33_groupi_n_3624, csa_tree_add_6_33_groupi_n_3625, csa_tree_add_6_33_groupi_n_3626, csa_tree_add_6_33_groupi_n_3627;
  wire csa_tree_add_6_33_groupi_n_3628, csa_tree_add_6_33_groupi_n_3629, csa_tree_add_6_33_groupi_n_3630, csa_tree_add_6_33_groupi_n_3631, csa_tree_add_6_33_groupi_n_3632, csa_tree_add_6_33_groupi_n_3633, csa_tree_add_6_33_groupi_n_3634, csa_tree_add_6_33_groupi_n_3635;
  wire csa_tree_add_6_33_groupi_n_3636, csa_tree_add_6_33_groupi_n_3637, csa_tree_add_6_33_groupi_n_3638, csa_tree_add_6_33_groupi_n_3639, csa_tree_add_6_33_groupi_n_3640, csa_tree_add_6_33_groupi_n_3641, csa_tree_add_6_33_groupi_n_3642, csa_tree_add_6_33_groupi_n_3643;
  wire csa_tree_add_6_33_groupi_n_3644, csa_tree_add_6_33_groupi_n_3645, csa_tree_add_6_33_groupi_n_3646, csa_tree_add_6_33_groupi_n_3647, csa_tree_add_6_33_groupi_n_3648, csa_tree_add_6_33_groupi_n_3649, csa_tree_add_6_33_groupi_n_3650, csa_tree_add_6_33_groupi_n_3651;
  wire csa_tree_add_6_33_groupi_n_3652, csa_tree_add_6_33_groupi_n_3653, csa_tree_add_6_33_groupi_n_3654, csa_tree_add_6_33_groupi_n_3655, csa_tree_add_6_33_groupi_n_3656, csa_tree_add_6_33_groupi_n_3657, csa_tree_add_6_33_groupi_n_3658, csa_tree_add_6_33_groupi_n_3659;
  wire csa_tree_add_6_33_groupi_n_3660, csa_tree_add_6_33_groupi_n_3661, csa_tree_add_6_33_groupi_n_3662, csa_tree_add_6_33_groupi_n_3663, csa_tree_add_6_33_groupi_n_3664, csa_tree_add_6_33_groupi_n_3665, csa_tree_add_6_33_groupi_n_3666, csa_tree_add_6_33_groupi_n_3667;
  wire csa_tree_add_6_33_groupi_n_3668, csa_tree_add_6_33_groupi_n_3669, csa_tree_add_6_33_groupi_n_3670, csa_tree_add_6_33_groupi_n_3671, csa_tree_add_6_33_groupi_n_3672, csa_tree_add_6_33_groupi_n_3673, csa_tree_add_6_33_groupi_n_3674, csa_tree_add_6_33_groupi_n_3675;
  wire csa_tree_add_6_33_groupi_n_3676, csa_tree_add_6_33_groupi_n_3677, csa_tree_add_6_33_groupi_n_3678, csa_tree_add_6_33_groupi_n_3679, csa_tree_add_6_33_groupi_n_3680, csa_tree_add_6_33_groupi_n_3681, csa_tree_add_6_33_groupi_n_3682, csa_tree_add_6_33_groupi_n_3683;
  wire csa_tree_add_6_33_groupi_n_3684, csa_tree_add_6_33_groupi_n_3685, csa_tree_add_6_33_groupi_n_3686, csa_tree_add_6_33_groupi_n_3687, csa_tree_add_6_33_groupi_n_3688, csa_tree_add_6_33_groupi_n_3689, csa_tree_add_6_33_groupi_n_3690, csa_tree_add_6_33_groupi_n_3691;
  wire csa_tree_add_6_33_groupi_n_3692, csa_tree_add_6_33_groupi_n_3693, csa_tree_add_6_33_groupi_n_3694, csa_tree_add_6_33_groupi_n_3695, csa_tree_add_6_33_groupi_n_3696, csa_tree_add_6_33_groupi_n_3697, csa_tree_add_6_33_groupi_n_3698, csa_tree_add_6_33_groupi_n_3699;
  wire csa_tree_add_6_33_groupi_n_3700, csa_tree_add_6_33_groupi_n_3701, csa_tree_add_6_33_groupi_n_3702, csa_tree_add_6_33_groupi_n_3703, csa_tree_add_6_33_groupi_n_3704, csa_tree_add_6_33_groupi_n_3705, csa_tree_add_6_33_groupi_n_3706, csa_tree_add_6_33_groupi_n_3707;
  wire csa_tree_add_6_33_groupi_n_3708, csa_tree_add_6_33_groupi_n_3709, csa_tree_add_6_33_groupi_n_3710, csa_tree_add_6_33_groupi_n_3711, csa_tree_add_6_33_groupi_n_3712, csa_tree_add_6_33_groupi_n_3713, csa_tree_add_6_33_groupi_n_3714, csa_tree_add_6_33_groupi_n_3715;
  wire csa_tree_add_6_33_groupi_n_3716, csa_tree_add_6_33_groupi_n_3717, csa_tree_add_6_33_groupi_n_3718, csa_tree_add_6_33_groupi_n_3719, csa_tree_add_6_33_groupi_n_3720, csa_tree_add_6_33_groupi_n_3721, csa_tree_add_6_33_groupi_n_3722, csa_tree_add_6_33_groupi_n_3723;
  wire csa_tree_add_6_33_groupi_n_3724, csa_tree_add_6_33_groupi_n_3725, csa_tree_add_6_33_groupi_n_3726, csa_tree_add_6_33_groupi_n_3727, csa_tree_add_6_33_groupi_n_3728, csa_tree_add_6_33_groupi_n_3729, csa_tree_add_6_33_groupi_n_3730, csa_tree_add_6_33_groupi_n_3731;
  wire csa_tree_add_6_33_groupi_n_3732, csa_tree_add_6_33_groupi_n_3733, csa_tree_add_6_33_groupi_n_3734, csa_tree_add_6_33_groupi_n_3735, csa_tree_add_6_33_groupi_n_3736, csa_tree_add_6_33_groupi_n_3737, csa_tree_add_6_33_groupi_n_3738, csa_tree_add_6_33_groupi_n_3739;
  wire csa_tree_add_6_33_groupi_n_3740, csa_tree_add_6_33_groupi_n_3741, csa_tree_add_6_33_groupi_n_3742, csa_tree_add_6_33_groupi_n_3743, csa_tree_add_6_33_groupi_n_3744, csa_tree_add_6_33_groupi_n_3745, csa_tree_add_6_33_groupi_n_3746, csa_tree_add_6_33_groupi_n_3747;
  wire csa_tree_add_6_33_groupi_n_3748, csa_tree_add_6_33_groupi_n_3749, csa_tree_add_6_33_groupi_n_3750, csa_tree_add_6_33_groupi_n_3751, csa_tree_add_6_33_groupi_n_3752, csa_tree_add_6_33_groupi_n_3753, csa_tree_add_6_33_groupi_n_3754, csa_tree_add_6_33_groupi_n_3755;
  wire csa_tree_add_6_33_groupi_n_3756, csa_tree_add_6_33_groupi_n_3757, csa_tree_add_6_33_groupi_n_3758, csa_tree_add_6_33_groupi_n_3759, csa_tree_add_6_33_groupi_n_3760, csa_tree_add_6_33_groupi_n_3761, csa_tree_add_6_33_groupi_n_3762, csa_tree_add_6_33_groupi_n_3763;
  wire csa_tree_add_6_33_groupi_n_3764, csa_tree_add_6_33_groupi_n_3765, csa_tree_add_6_33_groupi_n_3766, csa_tree_add_6_33_groupi_n_3767, csa_tree_add_6_33_groupi_n_3768, csa_tree_add_6_33_groupi_n_3769, csa_tree_add_6_33_groupi_n_3770, csa_tree_add_6_33_groupi_n_3771;
  wire csa_tree_add_6_33_groupi_n_3772, csa_tree_add_6_33_groupi_n_3773, csa_tree_add_6_33_groupi_n_3774, csa_tree_add_6_33_groupi_n_3775, csa_tree_add_6_33_groupi_n_3776, csa_tree_add_6_33_groupi_n_3777, csa_tree_add_6_33_groupi_n_3778, csa_tree_add_6_33_groupi_n_3779;
  wire csa_tree_add_6_33_groupi_n_3780, csa_tree_add_6_33_groupi_n_3781, csa_tree_add_6_33_groupi_n_3782, csa_tree_add_6_33_groupi_n_3783, csa_tree_add_6_33_groupi_n_3784, csa_tree_add_6_33_groupi_n_3785, csa_tree_add_6_33_groupi_n_3786, csa_tree_add_6_33_groupi_n_3787;
  wire csa_tree_add_6_33_groupi_n_3788, csa_tree_add_6_33_groupi_n_3789, csa_tree_add_6_33_groupi_n_3790, csa_tree_add_6_33_groupi_n_3791, csa_tree_add_6_33_groupi_n_3792, csa_tree_add_6_33_groupi_n_3793, csa_tree_add_6_33_groupi_n_3794, csa_tree_add_6_33_groupi_n_3795;
  wire csa_tree_add_6_33_groupi_n_3796, csa_tree_add_6_33_groupi_n_3797, csa_tree_add_6_33_groupi_n_3798, csa_tree_add_6_33_groupi_n_3799, csa_tree_add_6_33_groupi_n_3800, csa_tree_add_6_33_groupi_n_3801, csa_tree_add_6_33_groupi_n_3802, csa_tree_add_6_33_groupi_n_3803;
  wire csa_tree_add_6_33_groupi_n_3804, csa_tree_add_6_33_groupi_n_3805, csa_tree_add_6_33_groupi_n_3806, csa_tree_add_6_33_groupi_n_3807, csa_tree_add_6_33_groupi_n_3808, csa_tree_add_6_33_groupi_n_3809, csa_tree_add_6_33_groupi_n_3810, csa_tree_add_6_33_groupi_n_3811;
  wire csa_tree_add_6_33_groupi_n_3812, csa_tree_add_6_33_groupi_n_3813, csa_tree_add_6_33_groupi_n_3814, csa_tree_add_6_33_groupi_n_3815, csa_tree_add_6_33_groupi_n_3816, csa_tree_add_6_33_groupi_n_3817, csa_tree_add_6_33_groupi_n_3818, csa_tree_add_6_33_groupi_n_3819;
  wire csa_tree_add_6_33_groupi_n_3820, csa_tree_add_6_33_groupi_n_3821, csa_tree_add_6_33_groupi_n_3822, csa_tree_add_6_33_groupi_n_3823, csa_tree_add_6_33_groupi_n_3824, csa_tree_add_6_33_groupi_n_3825, csa_tree_add_6_33_groupi_n_3826, csa_tree_add_6_33_groupi_n_3827;
  wire csa_tree_add_6_33_groupi_n_3828, csa_tree_add_6_33_groupi_n_3829, csa_tree_add_6_33_groupi_n_3830, csa_tree_add_6_33_groupi_n_3831, csa_tree_add_6_33_groupi_n_3832, csa_tree_add_6_33_groupi_n_3833, csa_tree_add_6_33_groupi_n_3834, csa_tree_add_6_33_groupi_n_3835;
  wire csa_tree_add_6_33_groupi_n_3836, csa_tree_add_6_33_groupi_n_3837, csa_tree_add_6_33_groupi_n_3838, csa_tree_add_6_33_groupi_n_3839, csa_tree_add_6_33_groupi_n_3840, csa_tree_add_6_33_groupi_n_3841, csa_tree_add_6_33_groupi_n_3842, csa_tree_add_6_33_groupi_n_3843;
  wire csa_tree_add_6_33_groupi_n_3844, csa_tree_add_6_33_groupi_n_3845, csa_tree_add_6_33_groupi_n_3846, csa_tree_add_6_33_groupi_n_3847, csa_tree_add_6_33_groupi_n_3848, csa_tree_add_6_33_groupi_n_3849, csa_tree_add_6_33_groupi_n_3850, csa_tree_add_6_33_groupi_n_3851;
  wire csa_tree_add_6_33_groupi_n_3852, csa_tree_add_6_33_groupi_n_3853, csa_tree_add_6_33_groupi_n_3854, csa_tree_add_6_33_groupi_n_3855, csa_tree_add_6_33_groupi_n_3856, csa_tree_add_6_33_groupi_n_3857, csa_tree_add_6_33_groupi_n_3858, csa_tree_add_6_33_groupi_n_3859;
  wire csa_tree_add_6_33_groupi_n_3860, csa_tree_add_6_33_groupi_n_3861, csa_tree_add_6_33_groupi_n_3862, csa_tree_add_6_33_groupi_n_3863, csa_tree_add_6_33_groupi_n_3864, csa_tree_add_6_33_groupi_n_3865, csa_tree_add_6_33_groupi_n_3866, csa_tree_add_6_33_groupi_n_3867;
  wire csa_tree_add_6_33_groupi_n_3868, csa_tree_add_6_33_groupi_n_3869, csa_tree_add_6_33_groupi_n_3870, csa_tree_add_6_33_groupi_n_3871, csa_tree_add_6_33_groupi_n_3872, csa_tree_add_6_33_groupi_n_3873, csa_tree_add_6_33_groupi_n_3874, csa_tree_add_6_33_groupi_n_3875;
  wire csa_tree_add_6_33_groupi_n_3876, csa_tree_add_6_33_groupi_n_3877, csa_tree_add_6_33_groupi_n_3878, csa_tree_add_6_33_groupi_n_3879, csa_tree_add_6_33_groupi_n_3880, csa_tree_add_6_33_groupi_n_3881, csa_tree_add_6_33_groupi_n_3882, csa_tree_add_6_33_groupi_n_3883;
  wire csa_tree_add_6_33_groupi_n_3884, csa_tree_add_6_33_groupi_n_3885, csa_tree_add_6_33_groupi_n_3886, csa_tree_add_6_33_groupi_n_3887, csa_tree_add_6_33_groupi_n_3888, csa_tree_add_6_33_groupi_n_3889, csa_tree_add_6_33_groupi_n_3890, csa_tree_add_6_33_groupi_n_3891;
  wire csa_tree_add_6_33_groupi_n_3892, csa_tree_add_6_33_groupi_n_3893, csa_tree_add_6_33_groupi_n_3894, csa_tree_add_6_33_groupi_n_3895, csa_tree_add_6_33_groupi_n_3896, csa_tree_add_6_33_groupi_n_3897, csa_tree_add_6_33_groupi_n_3898, csa_tree_add_6_33_groupi_n_3899;
  wire csa_tree_add_6_33_groupi_n_3900, csa_tree_add_6_33_groupi_n_3901, csa_tree_add_6_33_groupi_n_3902, csa_tree_add_6_33_groupi_n_3903, csa_tree_add_6_33_groupi_n_3904, csa_tree_add_6_33_groupi_n_3905, csa_tree_add_6_33_groupi_n_3906, csa_tree_add_6_33_groupi_n_3907;
  wire csa_tree_add_6_33_groupi_n_3908, csa_tree_add_6_33_groupi_n_3909, csa_tree_add_6_33_groupi_n_3910, csa_tree_add_6_33_groupi_n_3911, csa_tree_add_6_33_groupi_n_3912, csa_tree_add_6_33_groupi_n_3913, csa_tree_add_6_33_groupi_n_3914, csa_tree_add_6_33_groupi_n_3915;
  wire csa_tree_add_6_33_groupi_n_3916, csa_tree_add_6_33_groupi_n_3917, csa_tree_add_6_33_groupi_n_3918, csa_tree_add_6_33_groupi_n_3919, csa_tree_add_6_33_groupi_n_3920, csa_tree_add_6_33_groupi_n_3921, csa_tree_add_6_33_groupi_n_3922, csa_tree_add_6_33_groupi_n_3923;
  wire csa_tree_add_6_33_groupi_n_3924, csa_tree_add_6_33_groupi_n_3925, csa_tree_add_6_33_groupi_n_3926, csa_tree_add_6_33_groupi_n_3927, csa_tree_add_6_33_groupi_n_3928, csa_tree_add_6_33_groupi_n_3929, csa_tree_add_6_33_groupi_n_3930, csa_tree_add_6_33_groupi_n_3931;
  wire csa_tree_add_6_33_groupi_n_3932, csa_tree_add_6_33_groupi_n_3933, csa_tree_add_6_33_groupi_n_3934, csa_tree_add_6_33_groupi_n_3935, csa_tree_add_6_33_groupi_n_3936, csa_tree_add_6_33_groupi_n_3937, csa_tree_add_6_33_groupi_n_3938, csa_tree_add_6_33_groupi_n_3939;
  wire csa_tree_add_6_33_groupi_n_3940, csa_tree_add_6_33_groupi_n_3941, csa_tree_add_6_33_groupi_n_3942, csa_tree_add_6_33_groupi_n_3943, csa_tree_add_6_33_groupi_n_3944, csa_tree_add_6_33_groupi_n_3945, csa_tree_add_6_33_groupi_n_3946, csa_tree_add_6_33_groupi_n_3947;
  wire csa_tree_add_6_33_groupi_n_3948, csa_tree_add_6_33_groupi_n_3949, csa_tree_add_6_33_groupi_n_3951, csa_tree_add_6_33_groupi_n_3952, csa_tree_add_6_33_groupi_n_3953, csa_tree_add_6_33_groupi_n_3954, csa_tree_add_6_33_groupi_n_3955, csa_tree_add_6_33_groupi_n_3956;
  wire csa_tree_add_6_33_groupi_n_3957, csa_tree_add_6_33_groupi_n_3958, csa_tree_add_6_33_groupi_n_3959, csa_tree_add_6_33_groupi_n_3960, csa_tree_add_6_33_groupi_n_3961, csa_tree_add_6_33_groupi_n_3962, csa_tree_add_6_33_groupi_n_3963, csa_tree_add_6_33_groupi_n_3964;
  wire csa_tree_add_6_33_groupi_n_3965, csa_tree_add_6_33_groupi_n_3966, csa_tree_add_6_33_groupi_n_3967, csa_tree_add_6_33_groupi_n_3968, csa_tree_add_6_33_groupi_n_3969, csa_tree_add_6_33_groupi_n_3970, csa_tree_add_6_33_groupi_n_3971, csa_tree_add_6_33_groupi_n_3972;
  wire csa_tree_add_6_33_groupi_n_3973, csa_tree_add_6_33_groupi_n_3974, csa_tree_add_6_33_groupi_n_3975, csa_tree_add_6_33_groupi_n_3976, csa_tree_add_6_33_groupi_n_3977, csa_tree_add_6_33_groupi_n_3978, csa_tree_add_6_33_groupi_n_3979, csa_tree_add_6_33_groupi_n_3980;
  wire csa_tree_add_6_33_groupi_n_3981, csa_tree_add_6_33_groupi_n_3982, csa_tree_add_6_33_groupi_n_3983, csa_tree_add_6_33_groupi_n_3984, csa_tree_add_6_33_groupi_n_3985, csa_tree_add_6_33_groupi_n_3986, csa_tree_add_6_33_groupi_n_3987, csa_tree_add_6_33_groupi_n_3988;
  wire csa_tree_add_6_33_groupi_n_3989, csa_tree_add_6_33_groupi_n_3990, csa_tree_add_6_33_groupi_n_3991, csa_tree_add_6_33_groupi_n_3992, csa_tree_add_6_33_groupi_n_3993, csa_tree_add_6_33_groupi_n_3994, csa_tree_add_6_33_groupi_n_3995, csa_tree_add_6_33_groupi_n_3996;
  wire csa_tree_add_6_33_groupi_n_3997, csa_tree_add_6_33_groupi_n_3998, csa_tree_add_6_33_groupi_n_3999, csa_tree_add_6_33_groupi_n_4000, csa_tree_add_6_33_groupi_n_4001, csa_tree_add_6_33_groupi_n_4002, csa_tree_add_6_33_groupi_n_4003, csa_tree_add_6_33_groupi_n_4004;
  wire csa_tree_add_6_33_groupi_n_4005, csa_tree_add_6_33_groupi_n_4006, csa_tree_add_6_33_groupi_n_4007, csa_tree_add_6_33_groupi_n_4008, csa_tree_add_6_33_groupi_n_4009, csa_tree_add_6_33_groupi_n_4010, csa_tree_add_6_33_groupi_n_4011, csa_tree_add_6_33_groupi_n_4012;
  wire csa_tree_add_6_33_groupi_n_4013, csa_tree_add_6_33_groupi_n_4014, csa_tree_add_6_33_groupi_n_4015, csa_tree_add_6_33_groupi_n_4016, csa_tree_add_6_33_groupi_n_4017, csa_tree_add_6_33_groupi_n_4018, csa_tree_add_6_33_groupi_n_4019, csa_tree_add_6_33_groupi_n_4020;
  wire csa_tree_add_6_33_groupi_n_4021, csa_tree_add_6_33_groupi_n_4022, csa_tree_add_6_33_groupi_n_4023, csa_tree_add_6_33_groupi_n_4024, csa_tree_add_6_33_groupi_n_4025, csa_tree_add_6_33_groupi_n_4026, csa_tree_add_6_33_groupi_n_4027, csa_tree_add_6_33_groupi_n_4028;
  wire csa_tree_add_6_33_groupi_n_4029, csa_tree_add_6_33_groupi_n_4030, csa_tree_add_6_33_groupi_n_4031, csa_tree_add_6_33_groupi_n_4032, csa_tree_add_6_33_groupi_n_4033, csa_tree_add_6_33_groupi_n_4034, csa_tree_add_6_33_groupi_n_4035, csa_tree_add_6_33_groupi_n_4036;
  wire csa_tree_add_6_33_groupi_n_4037, csa_tree_add_6_33_groupi_n_4038, csa_tree_add_6_33_groupi_n_4039, csa_tree_add_6_33_groupi_n_4040, csa_tree_add_6_33_groupi_n_4041, csa_tree_add_6_33_groupi_n_4042, csa_tree_add_6_33_groupi_n_4043, csa_tree_add_6_33_groupi_n_4044;
  wire csa_tree_add_6_33_groupi_n_4045, csa_tree_add_6_33_groupi_n_4046, csa_tree_add_6_33_groupi_n_4047, csa_tree_add_6_33_groupi_n_4048, csa_tree_add_6_33_groupi_n_4049, csa_tree_add_6_33_groupi_n_4050, csa_tree_add_6_33_groupi_n_4051, csa_tree_add_6_33_groupi_n_4052;
  wire csa_tree_add_6_33_groupi_n_4053, csa_tree_add_6_33_groupi_n_4054, csa_tree_add_6_33_groupi_n_4055, csa_tree_add_6_33_groupi_n_4056, csa_tree_add_6_33_groupi_n_4057, csa_tree_add_6_33_groupi_n_4058, csa_tree_add_6_33_groupi_n_4059, csa_tree_add_6_33_groupi_n_4060;
  wire csa_tree_add_6_33_groupi_n_4061, csa_tree_add_6_33_groupi_n_4062, csa_tree_add_6_33_groupi_n_4063, csa_tree_add_6_33_groupi_n_4064, csa_tree_add_6_33_groupi_n_4065, csa_tree_add_6_33_groupi_n_4066, csa_tree_add_6_33_groupi_n_4067, csa_tree_add_6_33_groupi_n_4068;
  wire csa_tree_add_6_33_groupi_n_4069, csa_tree_add_6_33_groupi_n_4070, csa_tree_add_6_33_groupi_n_4071, csa_tree_add_6_33_groupi_n_4072, csa_tree_add_6_33_groupi_n_4073, csa_tree_add_6_33_groupi_n_4074, csa_tree_add_6_33_groupi_n_4075, csa_tree_add_6_33_groupi_n_4076;
  wire csa_tree_add_6_33_groupi_n_4077, csa_tree_add_6_33_groupi_n_4078, csa_tree_add_6_33_groupi_n_4079, csa_tree_add_6_33_groupi_n_4080, csa_tree_add_6_33_groupi_n_4081, csa_tree_add_6_33_groupi_n_4082, csa_tree_add_6_33_groupi_n_4083, csa_tree_add_6_33_groupi_n_4084;
  wire csa_tree_add_6_33_groupi_n_4085, csa_tree_add_6_33_groupi_n_4086, csa_tree_add_6_33_groupi_n_4087, csa_tree_add_6_33_groupi_n_4088, csa_tree_add_6_33_groupi_n_4089, csa_tree_add_6_33_groupi_n_4090, csa_tree_add_6_33_groupi_n_4091, csa_tree_add_6_33_groupi_n_4092;
  wire csa_tree_add_6_33_groupi_n_4093, csa_tree_add_6_33_groupi_n_4094, csa_tree_add_6_33_groupi_n_4095, csa_tree_add_6_33_groupi_n_4096, csa_tree_add_6_33_groupi_n_4097, csa_tree_add_6_33_groupi_n_4098, csa_tree_add_6_33_groupi_n_4099, csa_tree_add_6_33_groupi_n_4100;
  wire csa_tree_add_6_33_groupi_n_4101, csa_tree_add_6_33_groupi_n_4102, csa_tree_add_6_33_groupi_n_4103, csa_tree_add_6_33_groupi_n_4104, csa_tree_add_6_33_groupi_n_4105, csa_tree_add_6_33_groupi_n_4106, csa_tree_add_6_33_groupi_n_4107, csa_tree_add_6_33_groupi_n_4108;
  wire csa_tree_add_6_33_groupi_n_4109, csa_tree_add_6_33_groupi_n_4110, csa_tree_add_6_33_groupi_n_4111, csa_tree_add_6_33_groupi_n_4112, csa_tree_add_6_33_groupi_n_4113, csa_tree_add_6_33_groupi_n_4114, csa_tree_add_6_33_groupi_n_4115, csa_tree_add_6_33_groupi_n_4116;
  wire csa_tree_add_6_33_groupi_n_4117, csa_tree_add_6_33_groupi_n_4118, csa_tree_add_6_33_groupi_n_4119, csa_tree_add_6_33_groupi_n_4120, csa_tree_add_6_33_groupi_n_4121, csa_tree_add_6_33_groupi_n_4122, csa_tree_add_6_33_groupi_n_4123, csa_tree_add_6_33_groupi_n_4124;
  wire csa_tree_add_6_33_groupi_n_4125, csa_tree_add_6_33_groupi_n_4126, csa_tree_add_6_33_groupi_n_4127, csa_tree_add_6_33_groupi_n_4128, csa_tree_add_6_33_groupi_n_4129, csa_tree_add_6_33_groupi_n_4130, csa_tree_add_6_33_groupi_n_4131, csa_tree_add_6_33_groupi_n_4132;
  wire csa_tree_add_6_33_groupi_n_4133, csa_tree_add_6_33_groupi_n_4134, csa_tree_add_6_33_groupi_n_4135, csa_tree_add_6_33_groupi_n_4136, csa_tree_add_6_33_groupi_n_4137, csa_tree_add_6_33_groupi_n_4138, csa_tree_add_6_33_groupi_n_4139, csa_tree_add_6_33_groupi_n_4140;
  wire csa_tree_add_6_33_groupi_n_4141, csa_tree_add_6_33_groupi_n_4142, csa_tree_add_6_33_groupi_n_4143, csa_tree_add_6_33_groupi_n_4144, csa_tree_add_6_33_groupi_n_4145, csa_tree_add_6_33_groupi_n_4146, csa_tree_add_6_33_groupi_n_4147, csa_tree_add_6_33_groupi_n_4148;
  wire csa_tree_add_6_33_groupi_n_4149, csa_tree_add_6_33_groupi_n_4150, csa_tree_add_6_33_groupi_n_4151, csa_tree_add_6_33_groupi_n_4152, csa_tree_add_6_33_groupi_n_4153, csa_tree_add_6_33_groupi_n_4154, csa_tree_add_6_33_groupi_n_4155, csa_tree_add_6_33_groupi_n_4156;
  wire csa_tree_add_6_33_groupi_n_4157, csa_tree_add_6_33_groupi_n_4158, csa_tree_add_6_33_groupi_n_4159, csa_tree_add_6_33_groupi_n_4160, csa_tree_add_6_33_groupi_n_4161, csa_tree_add_6_33_groupi_n_4162, csa_tree_add_6_33_groupi_n_4163, csa_tree_add_6_33_groupi_n_4164;
  wire csa_tree_add_6_33_groupi_n_4165, csa_tree_add_6_33_groupi_n_4166, csa_tree_add_6_33_groupi_n_4167, csa_tree_add_6_33_groupi_n_4168, csa_tree_add_6_33_groupi_n_4169, csa_tree_add_6_33_groupi_n_4170, csa_tree_add_6_33_groupi_n_4171, csa_tree_add_6_33_groupi_n_4172;
  wire csa_tree_add_6_33_groupi_n_4173, csa_tree_add_6_33_groupi_n_4174, csa_tree_add_6_33_groupi_n_4175, csa_tree_add_6_33_groupi_n_4176, csa_tree_add_6_33_groupi_n_4177, csa_tree_add_6_33_groupi_n_4178, csa_tree_add_6_33_groupi_n_4179, csa_tree_add_6_33_groupi_n_4180;
  wire csa_tree_add_6_33_groupi_n_4181, csa_tree_add_6_33_groupi_n_4182, csa_tree_add_6_33_groupi_n_4183, csa_tree_add_6_33_groupi_n_4184, csa_tree_add_6_33_groupi_n_4185, csa_tree_add_6_33_groupi_n_4186, csa_tree_add_6_33_groupi_n_4187, csa_tree_add_6_33_groupi_n_4188;
  wire csa_tree_add_6_33_groupi_n_4189, csa_tree_add_6_33_groupi_n_4190, csa_tree_add_6_33_groupi_n_4192, csa_tree_add_6_33_groupi_n_4193, csa_tree_add_6_33_groupi_n_4194, csa_tree_add_6_33_groupi_n_4195, csa_tree_add_6_33_groupi_n_4196, csa_tree_add_6_33_groupi_n_4197;
  wire csa_tree_add_6_33_groupi_n_4198, csa_tree_add_6_33_groupi_n_4199, csa_tree_add_6_33_groupi_n_4200, csa_tree_add_6_33_groupi_n_4201, csa_tree_add_6_33_groupi_n_4202, csa_tree_add_6_33_groupi_n_4203, csa_tree_add_6_33_groupi_n_4204, csa_tree_add_6_33_groupi_n_4205;
  wire csa_tree_add_6_33_groupi_n_4206, csa_tree_add_6_33_groupi_n_4207, csa_tree_add_6_33_groupi_n_4208, csa_tree_add_6_33_groupi_n_4209, csa_tree_add_6_33_groupi_n_4210, csa_tree_add_6_33_groupi_n_4211, csa_tree_add_6_33_groupi_n_4212, csa_tree_add_6_33_groupi_n_4213;
  wire csa_tree_add_6_33_groupi_n_4214, csa_tree_add_6_33_groupi_n_4215, csa_tree_add_6_33_groupi_n_4216, csa_tree_add_6_33_groupi_n_4217, csa_tree_add_6_33_groupi_n_4218, csa_tree_add_6_33_groupi_n_4219, csa_tree_add_6_33_groupi_n_4220, csa_tree_add_6_33_groupi_n_4221;
  wire csa_tree_add_6_33_groupi_n_4222, csa_tree_add_6_33_groupi_n_4223, csa_tree_add_6_33_groupi_n_4224, csa_tree_add_6_33_groupi_n_4225, csa_tree_add_6_33_groupi_n_4226, csa_tree_add_6_33_groupi_n_4227, csa_tree_add_6_33_groupi_n_4228, csa_tree_add_6_33_groupi_n_4229;
  wire csa_tree_add_6_33_groupi_n_4230, csa_tree_add_6_33_groupi_n_4231, csa_tree_add_6_33_groupi_n_4232, csa_tree_add_6_33_groupi_n_4233, csa_tree_add_6_33_groupi_n_4234, csa_tree_add_6_33_groupi_n_4235, csa_tree_add_6_33_groupi_n_4236, csa_tree_add_6_33_groupi_n_4237;
  wire csa_tree_add_6_33_groupi_n_4238, csa_tree_add_6_33_groupi_n_4239, csa_tree_add_6_33_groupi_n_4240, csa_tree_add_6_33_groupi_n_4241, csa_tree_add_6_33_groupi_n_4242, csa_tree_add_6_33_groupi_n_4243, csa_tree_add_6_33_groupi_n_4244, csa_tree_add_6_33_groupi_n_4245;
  wire csa_tree_add_6_33_groupi_n_4246, csa_tree_add_6_33_groupi_n_4247, csa_tree_add_6_33_groupi_n_4248, csa_tree_add_6_33_groupi_n_4249, csa_tree_add_6_33_groupi_n_4250, csa_tree_add_6_33_groupi_n_4251, csa_tree_add_6_33_groupi_n_4252, csa_tree_add_6_33_groupi_n_4253;
  wire csa_tree_add_6_33_groupi_n_4254, csa_tree_add_6_33_groupi_n_4255, csa_tree_add_6_33_groupi_n_4256, csa_tree_add_6_33_groupi_n_4257, csa_tree_add_6_33_groupi_n_4258, csa_tree_add_6_33_groupi_n_4259, csa_tree_add_6_33_groupi_n_4260, csa_tree_add_6_33_groupi_n_4261;
  wire csa_tree_add_6_33_groupi_n_4262, csa_tree_add_6_33_groupi_n_4263, csa_tree_add_6_33_groupi_n_4264, csa_tree_add_6_33_groupi_n_4265, csa_tree_add_6_33_groupi_n_4266, csa_tree_add_6_33_groupi_n_4267, csa_tree_add_6_33_groupi_n_4268, csa_tree_add_6_33_groupi_n_4269;
  wire csa_tree_add_6_33_groupi_n_4270, csa_tree_add_6_33_groupi_n_4271, csa_tree_add_6_33_groupi_n_4272, csa_tree_add_6_33_groupi_n_4273, csa_tree_add_6_33_groupi_n_4274, csa_tree_add_6_33_groupi_n_4275, csa_tree_add_6_33_groupi_n_4276, csa_tree_add_6_33_groupi_n_4277;
  wire csa_tree_add_6_33_groupi_n_4278, csa_tree_add_6_33_groupi_n_4279, csa_tree_add_6_33_groupi_n_4280, csa_tree_add_6_33_groupi_n_4281, csa_tree_add_6_33_groupi_n_4282, csa_tree_add_6_33_groupi_n_4283, csa_tree_add_6_33_groupi_n_4284, csa_tree_add_6_33_groupi_n_4285;
  wire csa_tree_add_6_33_groupi_n_4286, csa_tree_add_6_33_groupi_n_4287, csa_tree_add_6_33_groupi_n_4288, csa_tree_add_6_33_groupi_n_4289, csa_tree_add_6_33_groupi_n_4290, csa_tree_add_6_33_groupi_n_4291, csa_tree_add_6_33_groupi_n_4292, csa_tree_add_6_33_groupi_n_4293;
  wire csa_tree_add_6_33_groupi_n_4294, csa_tree_add_6_33_groupi_n_4295, csa_tree_add_6_33_groupi_n_4296, csa_tree_add_6_33_groupi_n_4297, csa_tree_add_6_33_groupi_n_4298, csa_tree_add_6_33_groupi_n_4299, csa_tree_add_6_33_groupi_n_4300, csa_tree_add_6_33_groupi_n_4301;
  wire csa_tree_add_6_33_groupi_n_4302, csa_tree_add_6_33_groupi_n_4303, csa_tree_add_6_33_groupi_n_4304, csa_tree_add_6_33_groupi_n_4305, csa_tree_add_6_33_groupi_n_4306, csa_tree_add_6_33_groupi_n_4307, csa_tree_add_6_33_groupi_n_4308, csa_tree_add_6_33_groupi_n_4309;
  wire csa_tree_add_6_33_groupi_n_4310, csa_tree_add_6_33_groupi_n_4311, csa_tree_add_6_33_groupi_n_4312, csa_tree_add_6_33_groupi_n_4313, csa_tree_add_6_33_groupi_n_4314, csa_tree_add_6_33_groupi_n_4315, csa_tree_add_6_33_groupi_n_4316, csa_tree_add_6_33_groupi_n_4317;
  wire csa_tree_add_6_33_groupi_n_4318, csa_tree_add_6_33_groupi_n_4319, csa_tree_add_6_33_groupi_n_4320, csa_tree_add_6_33_groupi_n_4321, csa_tree_add_6_33_groupi_n_4322, csa_tree_add_6_33_groupi_n_4323, csa_tree_add_6_33_groupi_n_4324, csa_tree_add_6_33_groupi_n_4325;
  wire csa_tree_add_6_33_groupi_n_4326, csa_tree_add_6_33_groupi_n_4327, csa_tree_add_6_33_groupi_n_4328, csa_tree_add_6_33_groupi_n_4329, csa_tree_add_6_33_groupi_n_4330, csa_tree_add_6_33_groupi_n_4331, csa_tree_add_6_33_groupi_n_4332, csa_tree_add_6_33_groupi_n_4333;
  wire csa_tree_add_6_33_groupi_n_4334, csa_tree_add_6_33_groupi_n_4335, csa_tree_add_6_33_groupi_n_4336, csa_tree_add_6_33_groupi_n_4337, csa_tree_add_6_33_groupi_n_4338, csa_tree_add_6_33_groupi_n_4339, csa_tree_add_6_33_groupi_n_4340, csa_tree_add_6_33_groupi_n_4341;
  wire csa_tree_add_6_33_groupi_n_4342, csa_tree_add_6_33_groupi_n_4343, csa_tree_add_6_33_groupi_n_4344, csa_tree_add_6_33_groupi_n_4345, csa_tree_add_6_33_groupi_n_4346, csa_tree_add_6_33_groupi_n_4347, csa_tree_add_6_33_groupi_n_4348, csa_tree_add_6_33_groupi_n_4349;
  wire csa_tree_add_6_33_groupi_n_4350, csa_tree_add_6_33_groupi_n_4351, csa_tree_add_6_33_groupi_n_4352, csa_tree_add_6_33_groupi_n_4353, csa_tree_add_6_33_groupi_n_4354, csa_tree_add_6_33_groupi_n_4355, csa_tree_add_6_33_groupi_n_4356, csa_tree_add_6_33_groupi_n_4357;
  wire csa_tree_add_6_33_groupi_n_4358, csa_tree_add_6_33_groupi_n_4359, csa_tree_add_6_33_groupi_n_4360, csa_tree_add_6_33_groupi_n_4361, csa_tree_add_6_33_groupi_n_4362, csa_tree_add_6_33_groupi_n_4363, csa_tree_add_6_33_groupi_n_4364, csa_tree_add_6_33_groupi_n_4365;
  wire csa_tree_add_6_33_groupi_n_4366, csa_tree_add_6_33_groupi_n_4367, csa_tree_add_6_33_groupi_n_4368, csa_tree_add_6_33_groupi_n_4369, csa_tree_add_6_33_groupi_n_4370, csa_tree_add_6_33_groupi_n_4371, csa_tree_add_6_33_groupi_n_4372, csa_tree_add_6_33_groupi_n_4373;
  wire csa_tree_add_6_33_groupi_n_4374, csa_tree_add_6_33_groupi_n_4375, csa_tree_add_6_33_groupi_n_4376, csa_tree_add_6_33_groupi_n_4377, csa_tree_add_6_33_groupi_n_4378, csa_tree_add_6_33_groupi_n_4379, csa_tree_add_6_33_groupi_n_4380, csa_tree_add_6_33_groupi_n_4381;
  wire csa_tree_add_6_33_groupi_n_4382, csa_tree_add_6_33_groupi_n_4383, csa_tree_add_6_33_groupi_n_4384, csa_tree_add_6_33_groupi_n_4385, csa_tree_add_6_33_groupi_n_4386, csa_tree_add_6_33_groupi_n_4387, csa_tree_add_6_33_groupi_n_4388, csa_tree_add_6_33_groupi_n_4389;
  wire csa_tree_add_6_33_groupi_n_4390, csa_tree_add_6_33_groupi_n_4391, csa_tree_add_6_33_groupi_n_4392, csa_tree_add_6_33_groupi_n_4393, csa_tree_add_6_33_groupi_n_4394, csa_tree_add_6_33_groupi_n_4395, csa_tree_add_6_33_groupi_n_4396, csa_tree_add_6_33_groupi_n_4397;
  wire csa_tree_add_6_33_groupi_n_4398, csa_tree_add_6_33_groupi_n_4399, csa_tree_add_6_33_groupi_n_4400, csa_tree_add_6_33_groupi_n_4401, csa_tree_add_6_33_groupi_n_4402, csa_tree_add_6_33_groupi_n_4403, csa_tree_add_6_33_groupi_n_4404, csa_tree_add_6_33_groupi_n_4405;
  wire csa_tree_add_6_33_groupi_n_4406, csa_tree_add_6_33_groupi_n_4407, csa_tree_add_6_33_groupi_n_4408, csa_tree_add_6_33_groupi_n_4409, csa_tree_add_6_33_groupi_n_4411, csa_tree_add_6_33_groupi_n_4412, csa_tree_add_6_33_groupi_n_4413, csa_tree_add_6_33_groupi_n_4414;
  wire csa_tree_add_6_33_groupi_n_4415, csa_tree_add_6_33_groupi_n_4416, csa_tree_add_6_33_groupi_n_4417, csa_tree_add_6_33_groupi_n_4418, csa_tree_add_6_33_groupi_n_4419, csa_tree_add_6_33_groupi_n_4420, csa_tree_add_6_33_groupi_n_4421, csa_tree_add_6_33_groupi_n_4422;
  wire csa_tree_add_6_33_groupi_n_4423, csa_tree_add_6_33_groupi_n_4424, csa_tree_add_6_33_groupi_n_4425, csa_tree_add_6_33_groupi_n_4426, csa_tree_add_6_33_groupi_n_4427, csa_tree_add_6_33_groupi_n_4428, csa_tree_add_6_33_groupi_n_4429, csa_tree_add_6_33_groupi_n_4430;
  wire csa_tree_add_6_33_groupi_n_4431, csa_tree_add_6_33_groupi_n_4432, csa_tree_add_6_33_groupi_n_4433, csa_tree_add_6_33_groupi_n_4434, csa_tree_add_6_33_groupi_n_4435, csa_tree_add_6_33_groupi_n_4436, csa_tree_add_6_33_groupi_n_4437, csa_tree_add_6_33_groupi_n_4438;
  wire csa_tree_add_6_33_groupi_n_4439, csa_tree_add_6_33_groupi_n_4440, csa_tree_add_6_33_groupi_n_4441, csa_tree_add_6_33_groupi_n_4442, csa_tree_add_6_33_groupi_n_4443, csa_tree_add_6_33_groupi_n_4444, csa_tree_add_6_33_groupi_n_4445, csa_tree_add_6_33_groupi_n_4446;
  wire csa_tree_add_6_33_groupi_n_4447, csa_tree_add_6_33_groupi_n_4448, csa_tree_add_6_33_groupi_n_4449, csa_tree_add_6_33_groupi_n_4450, csa_tree_add_6_33_groupi_n_4451, csa_tree_add_6_33_groupi_n_4452, csa_tree_add_6_33_groupi_n_4453, csa_tree_add_6_33_groupi_n_4454;
  wire csa_tree_add_6_33_groupi_n_4455, csa_tree_add_6_33_groupi_n_4456, csa_tree_add_6_33_groupi_n_4457, csa_tree_add_6_33_groupi_n_4458, csa_tree_add_6_33_groupi_n_4459, csa_tree_add_6_33_groupi_n_4460, csa_tree_add_6_33_groupi_n_4461, csa_tree_add_6_33_groupi_n_4462;
  wire csa_tree_add_6_33_groupi_n_4463, csa_tree_add_6_33_groupi_n_4464, csa_tree_add_6_33_groupi_n_4465, csa_tree_add_6_33_groupi_n_4466, csa_tree_add_6_33_groupi_n_4467, csa_tree_add_6_33_groupi_n_4468, csa_tree_add_6_33_groupi_n_4469, csa_tree_add_6_33_groupi_n_4470;
  wire csa_tree_add_6_33_groupi_n_4471, csa_tree_add_6_33_groupi_n_4472, csa_tree_add_6_33_groupi_n_4473, csa_tree_add_6_33_groupi_n_4474, csa_tree_add_6_33_groupi_n_4475, csa_tree_add_6_33_groupi_n_4476, csa_tree_add_6_33_groupi_n_4477, csa_tree_add_6_33_groupi_n_4478;
  wire csa_tree_add_6_33_groupi_n_4479, csa_tree_add_6_33_groupi_n_4480, csa_tree_add_6_33_groupi_n_4481, csa_tree_add_6_33_groupi_n_4482, csa_tree_add_6_33_groupi_n_4483, csa_tree_add_6_33_groupi_n_4484, csa_tree_add_6_33_groupi_n_4485, csa_tree_add_6_33_groupi_n_4486;
  wire csa_tree_add_6_33_groupi_n_4487, csa_tree_add_6_33_groupi_n_4488, csa_tree_add_6_33_groupi_n_4489, csa_tree_add_6_33_groupi_n_4490, csa_tree_add_6_33_groupi_n_4491, csa_tree_add_6_33_groupi_n_4492, csa_tree_add_6_33_groupi_n_4493, csa_tree_add_6_33_groupi_n_4494;
  wire csa_tree_add_6_33_groupi_n_4495, csa_tree_add_6_33_groupi_n_4496, csa_tree_add_6_33_groupi_n_4497, csa_tree_add_6_33_groupi_n_4498, csa_tree_add_6_33_groupi_n_4499, csa_tree_add_6_33_groupi_n_4500, csa_tree_add_6_33_groupi_n_4501, csa_tree_add_6_33_groupi_n_4502;
  wire csa_tree_add_6_33_groupi_n_4503, csa_tree_add_6_33_groupi_n_4504, csa_tree_add_6_33_groupi_n_4505, csa_tree_add_6_33_groupi_n_4506, csa_tree_add_6_33_groupi_n_4507, csa_tree_add_6_33_groupi_n_4508, csa_tree_add_6_33_groupi_n_4509, csa_tree_add_6_33_groupi_n_4510;
  wire csa_tree_add_6_33_groupi_n_4511, csa_tree_add_6_33_groupi_n_4512, csa_tree_add_6_33_groupi_n_4513, csa_tree_add_6_33_groupi_n_4514, csa_tree_add_6_33_groupi_n_4515, csa_tree_add_6_33_groupi_n_4516, csa_tree_add_6_33_groupi_n_4517, csa_tree_add_6_33_groupi_n_4518;
  wire csa_tree_add_6_33_groupi_n_4519, csa_tree_add_6_33_groupi_n_4520, csa_tree_add_6_33_groupi_n_4521, csa_tree_add_6_33_groupi_n_4522, csa_tree_add_6_33_groupi_n_4523, csa_tree_add_6_33_groupi_n_4524, csa_tree_add_6_33_groupi_n_4525, csa_tree_add_6_33_groupi_n_4526;
  wire csa_tree_add_6_33_groupi_n_4527, csa_tree_add_6_33_groupi_n_4528, csa_tree_add_6_33_groupi_n_4529, csa_tree_add_6_33_groupi_n_4530, csa_tree_add_6_33_groupi_n_4531, csa_tree_add_6_33_groupi_n_4532, csa_tree_add_6_33_groupi_n_4533, csa_tree_add_6_33_groupi_n_4534;
  wire csa_tree_add_6_33_groupi_n_4535, csa_tree_add_6_33_groupi_n_4536, csa_tree_add_6_33_groupi_n_4537, csa_tree_add_6_33_groupi_n_4538, csa_tree_add_6_33_groupi_n_4539, csa_tree_add_6_33_groupi_n_4540, csa_tree_add_6_33_groupi_n_4541, csa_tree_add_6_33_groupi_n_4542;
  wire csa_tree_add_6_33_groupi_n_4543, csa_tree_add_6_33_groupi_n_4544, csa_tree_add_6_33_groupi_n_4545, csa_tree_add_6_33_groupi_n_4546, csa_tree_add_6_33_groupi_n_4547, csa_tree_add_6_33_groupi_n_4548, csa_tree_add_6_33_groupi_n_4549, csa_tree_add_6_33_groupi_n_4550;
  wire csa_tree_add_6_33_groupi_n_4551, csa_tree_add_6_33_groupi_n_4553, csa_tree_add_6_33_groupi_n_4554, csa_tree_add_6_33_groupi_n_4555, csa_tree_add_6_33_groupi_n_4556, csa_tree_add_6_33_groupi_n_4557, csa_tree_add_6_33_groupi_n_4558, csa_tree_add_6_33_groupi_n_4559;
  wire csa_tree_add_6_33_groupi_n_4560, csa_tree_add_6_33_groupi_n_4561, csa_tree_add_6_33_groupi_n_4562, csa_tree_add_6_33_groupi_n_4563, csa_tree_add_6_33_groupi_n_4564, csa_tree_add_6_33_groupi_n_4565, csa_tree_add_6_33_groupi_n_4566, csa_tree_add_6_33_groupi_n_4567;
  wire csa_tree_add_6_33_groupi_n_4568, csa_tree_add_6_33_groupi_n_4569, csa_tree_add_6_33_groupi_n_4570, csa_tree_add_6_33_groupi_n_4571, csa_tree_add_6_33_groupi_n_4572, csa_tree_add_6_33_groupi_n_4573, csa_tree_add_6_33_groupi_n_4574, csa_tree_add_6_33_groupi_n_4575;
  wire csa_tree_add_6_33_groupi_n_4576, csa_tree_add_6_33_groupi_n_4577, csa_tree_add_6_33_groupi_n_4578, csa_tree_add_6_33_groupi_n_4579, csa_tree_add_6_33_groupi_n_4580, csa_tree_add_6_33_groupi_n_4581, csa_tree_add_6_33_groupi_n_4582, csa_tree_add_6_33_groupi_n_4583;
  wire csa_tree_add_6_33_groupi_n_4584, csa_tree_add_6_33_groupi_n_4585, csa_tree_add_6_33_groupi_n_4586, csa_tree_add_6_33_groupi_n_4587, csa_tree_add_6_33_groupi_n_4588, csa_tree_add_6_33_groupi_n_4589, csa_tree_add_6_33_groupi_n_4590, csa_tree_add_6_33_groupi_n_4591;
  wire csa_tree_add_6_33_groupi_n_4592, csa_tree_add_6_33_groupi_n_4593, csa_tree_add_6_33_groupi_n_4594, csa_tree_add_6_33_groupi_n_4595, csa_tree_add_6_33_groupi_n_4596, csa_tree_add_6_33_groupi_n_4597, csa_tree_add_6_33_groupi_n_4598, csa_tree_add_6_33_groupi_n_4599;
  wire csa_tree_add_6_33_groupi_n_4600, csa_tree_add_6_33_groupi_n_4601, csa_tree_add_6_33_groupi_n_4602, csa_tree_add_6_33_groupi_n_4603, csa_tree_add_6_33_groupi_n_4604, csa_tree_add_6_33_groupi_n_4605, csa_tree_add_6_33_groupi_n_4606, csa_tree_add_6_33_groupi_n_4607;
  wire csa_tree_add_6_33_groupi_n_4608, csa_tree_add_6_33_groupi_n_4609, csa_tree_add_6_33_groupi_n_4610, csa_tree_add_6_33_groupi_n_4611, csa_tree_add_6_33_groupi_n_4612, csa_tree_add_6_33_groupi_n_4613, csa_tree_add_6_33_groupi_n_4614, csa_tree_add_6_33_groupi_n_4615;
  wire csa_tree_add_6_33_groupi_n_4616, csa_tree_add_6_33_groupi_n_4617, csa_tree_add_6_33_groupi_n_4618, csa_tree_add_6_33_groupi_n_4619, csa_tree_add_6_33_groupi_n_4620, csa_tree_add_6_33_groupi_n_4621, csa_tree_add_6_33_groupi_n_4622, csa_tree_add_6_33_groupi_n_4623;
  wire csa_tree_add_6_33_groupi_n_4624, csa_tree_add_6_33_groupi_n_4625, csa_tree_add_6_33_groupi_n_4626, csa_tree_add_6_33_groupi_n_4627, csa_tree_add_6_33_groupi_n_4628, csa_tree_add_6_33_groupi_n_4629, csa_tree_add_6_33_groupi_n_4630, csa_tree_add_6_33_groupi_n_4631;
  wire csa_tree_add_6_33_groupi_n_4632, csa_tree_add_6_33_groupi_n_4633, csa_tree_add_6_33_groupi_n_4634, csa_tree_add_6_33_groupi_n_4635, csa_tree_add_6_33_groupi_n_4636, csa_tree_add_6_33_groupi_n_4637, csa_tree_add_6_33_groupi_n_4638, csa_tree_add_6_33_groupi_n_4639;
  wire csa_tree_add_6_33_groupi_n_4640, csa_tree_add_6_33_groupi_n_4641, csa_tree_add_6_33_groupi_n_4642, csa_tree_add_6_33_groupi_n_4643, csa_tree_add_6_33_groupi_n_4644, csa_tree_add_6_33_groupi_n_4645, csa_tree_add_6_33_groupi_n_4646, csa_tree_add_6_33_groupi_n_4647;
  wire csa_tree_add_6_33_groupi_n_4648, csa_tree_add_6_33_groupi_n_4649, csa_tree_add_6_33_groupi_n_4650, csa_tree_add_6_33_groupi_n_4651, csa_tree_add_6_33_groupi_n_4652, csa_tree_add_6_33_groupi_n_4653, csa_tree_add_6_33_groupi_n_4654, csa_tree_add_6_33_groupi_n_4655;
  wire csa_tree_add_6_33_groupi_n_4656, csa_tree_add_6_33_groupi_n_4657, csa_tree_add_6_33_groupi_n_4658, csa_tree_add_6_33_groupi_n_4659, csa_tree_add_6_33_groupi_n_4660, csa_tree_add_6_33_groupi_n_4661, csa_tree_add_6_33_groupi_n_4662, csa_tree_add_6_33_groupi_n_4663;
  wire csa_tree_add_6_33_groupi_n_4664, csa_tree_add_6_33_groupi_n_4665, csa_tree_add_6_33_groupi_n_4666, csa_tree_add_6_33_groupi_n_4667, csa_tree_add_6_33_groupi_n_4668, csa_tree_add_6_33_groupi_n_4669, csa_tree_add_6_33_groupi_n_4670, csa_tree_add_6_33_groupi_n_4671;
  wire csa_tree_add_6_33_groupi_n_4672, csa_tree_add_6_33_groupi_n_4673, csa_tree_add_6_33_groupi_n_4674, csa_tree_add_6_33_groupi_n_4675, csa_tree_add_6_33_groupi_n_4676, csa_tree_add_6_33_groupi_n_4677, csa_tree_add_6_33_groupi_n_4678, csa_tree_add_6_33_groupi_n_4679;
  wire csa_tree_add_6_33_groupi_n_4680, csa_tree_add_6_33_groupi_n_4681, csa_tree_add_6_33_groupi_n_4682, csa_tree_add_6_33_groupi_n_4683, csa_tree_add_6_33_groupi_n_4684, csa_tree_add_6_33_groupi_n_4685, csa_tree_add_6_33_groupi_n_4687, csa_tree_add_6_33_groupi_n_4688;
  wire csa_tree_add_6_33_groupi_n_4689, csa_tree_add_6_33_groupi_n_4690, csa_tree_add_6_33_groupi_n_4691, csa_tree_add_6_33_groupi_n_4692, csa_tree_add_6_33_groupi_n_4693, csa_tree_add_6_33_groupi_n_4694, csa_tree_add_6_33_groupi_n_4695, csa_tree_add_6_33_groupi_n_4696;
  wire csa_tree_add_6_33_groupi_n_4697, csa_tree_add_6_33_groupi_n_4698, csa_tree_add_6_33_groupi_n_4699, csa_tree_add_6_33_groupi_n_4700, csa_tree_add_6_33_groupi_n_4701, csa_tree_add_6_33_groupi_n_4702, csa_tree_add_6_33_groupi_n_4703, csa_tree_add_6_33_groupi_n_4704;
  wire csa_tree_add_6_33_groupi_n_4705, csa_tree_add_6_33_groupi_n_4706, csa_tree_add_6_33_groupi_n_4707, csa_tree_add_6_33_groupi_n_4708, csa_tree_add_6_33_groupi_n_4709, csa_tree_add_6_33_groupi_n_4710, csa_tree_add_6_33_groupi_n_4711, csa_tree_add_6_33_groupi_n_4712;
  wire csa_tree_add_6_33_groupi_n_4713, csa_tree_add_6_33_groupi_n_4714, csa_tree_add_6_33_groupi_n_4715, csa_tree_add_6_33_groupi_n_4716, csa_tree_add_6_33_groupi_n_4717, csa_tree_add_6_33_groupi_n_4718, csa_tree_add_6_33_groupi_n_4719, csa_tree_add_6_33_groupi_n_4720;
  wire csa_tree_add_6_33_groupi_n_4721, csa_tree_add_6_33_groupi_n_4722, csa_tree_add_6_33_groupi_n_4723, csa_tree_add_6_33_groupi_n_4724, csa_tree_add_6_33_groupi_n_4725, csa_tree_add_6_33_groupi_n_4726, csa_tree_add_6_33_groupi_n_4727, csa_tree_add_6_33_groupi_n_4728;
  wire csa_tree_add_6_33_groupi_n_4729, csa_tree_add_6_33_groupi_n_4730, csa_tree_add_6_33_groupi_n_4731, csa_tree_add_6_33_groupi_n_4732, csa_tree_add_6_33_groupi_n_4733, csa_tree_add_6_33_groupi_n_4734, csa_tree_add_6_33_groupi_n_4735, csa_tree_add_6_33_groupi_n_4736;
  wire csa_tree_add_6_33_groupi_n_4737, csa_tree_add_6_33_groupi_n_4738, csa_tree_add_6_33_groupi_n_4739, csa_tree_add_6_33_groupi_n_4740, csa_tree_add_6_33_groupi_n_4741, csa_tree_add_6_33_groupi_n_4742, csa_tree_add_6_33_groupi_n_4743, csa_tree_add_6_33_groupi_n_4744;
  wire csa_tree_add_6_33_groupi_n_4745, csa_tree_add_6_33_groupi_n_4746, csa_tree_add_6_33_groupi_n_4747, csa_tree_add_6_33_groupi_n_4748, csa_tree_add_6_33_groupi_n_4749, csa_tree_add_6_33_groupi_n_4750, csa_tree_add_6_33_groupi_n_4751, csa_tree_add_6_33_groupi_n_4752;
  wire csa_tree_add_6_33_groupi_n_4753, csa_tree_add_6_33_groupi_n_4754, csa_tree_add_6_33_groupi_n_4755, csa_tree_add_6_33_groupi_n_4756, csa_tree_add_6_33_groupi_n_4757, csa_tree_add_6_33_groupi_n_4758, csa_tree_add_6_33_groupi_n_4759, csa_tree_add_6_33_groupi_n_4760;
  wire csa_tree_add_6_33_groupi_n_4761, csa_tree_add_6_33_groupi_n_4762, csa_tree_add_6_33_groupi_n_4763, csa_tree_add_6_33_groupi_n_4764, csa_tree_add_6_33_groupi_n_4766, csa_tree_add_6_33_groupi_n_4767, csa_tree_add_6_33_groupi_n_4768, csa_tree_add_6_33_groupi_n_4769;
  wire csa_tree_add_6_33_groupi_n_4770, csa_tree_add_6_33_groupi_n_4771, csa_tree_add_6_33_groupi_n_4772, csa_tree_add_6_33_groupi_n_4773, csa_tree_add_6_33_groupi_n_4774, csa_tree_add_6_33_groupi_n_4775, csa_tree_add_6_33_groupi_n_4776, csa_tree_add_6_33_groupi_n_4777;
  wire csa_tree_add_6_33_groupi_n_4778, csa_tree_add_6_33_groupi_n_4779, csa_tree_add_6_33_groupi_n_4780, csa_tree_add_6_33_groupi_n_4781, csa_tree_add_6_33_groupi_n_4782, csa_tree_add_6_33_groupi_n_4783, csa_tree_add_6_33_groupi_n_4784, csa_tree_add_6_33_groupi_n_4785;
  wire csa_tree_add_6_33_groupi_n_4786, csa_tree_add_6_33_groupi_n_4787, csa_tree_add_6_33_groupi_n_4788, csa_tree_add_6_33_groupi_n_4789, csa_tree_add_6_33_groupi_n_4790, csa_tree_add_6_33_groupi_n_4791, csa_tree_add_6_33_groupi_n_4792, csa_tree_add_6_33_groupi_n_4793;
  wire csa_tree_add_6_33_groupi_n_4794, csa_tree_add_6_33_groupi_n_4795, csa_tree_add_6_33_groupi_n_4796, csa_tree_add_6_33_groupi_n_4797, csa_tree_add_6_33_groupi_n_4798, csa_tree_add_6_33_groupi_n_4799, csa_tree_add_6_33_groupi_n_4800, csa_tree_add_6_33_groupi_n_4801;
  wire csa_tree_add_6_33_groupi_n_4802, csa_tree_add_6_33_groupi_n_4803, csa_tree_add_6_33_groupi_n_4804, csa_tree_add_6_33_groupi_n_4805, csa_tree_add_6_33_groupi_n_4806, csa_tree_add_6_33_groupi_n_4807, csa_tree_add_6_33_groupi_n_4808, csa_tree_add_6_33_groupi_n_4810;
  wire csa_tree_add_6_33_groupi_n_4811, csa_tree_add_6_33_groupi_n_4812, csa_tree_add_6_33_groupi_n_4813, csa_tree_add_6_33_groupi_n_4814, csa_tree_add_6_33_groupi_n_4815, csa_tree_add_6_33_groupi_n_4816, csa_tree_add_6_33_groupi_n_4817, csa_tree_add_6_33_groupi_n_4819;
  wire csa_tree_add_6_33_groupi_n_4820, csa_tree_add_6_33_groupi_n_4822, csa_tree_add_6_33_groupi_n_4823, csa_tree_add_6_33_groupi_n_4824, csa_tree_add_6_33_groupi_n_4826, csa_tree_add_6_33_groupi_n_4827, csa_tree_add_6_33_groupi_n_4828, csa_tree_add_6_33_groupi_n_4829;
  wire csa_tree_add_6_33_groupi_n_4830, csa_tree_add_6_33_groupi_n_4831, csa_tree_add_6_33_groupi_n_4832, csa_tree_add_6_33_groupi_n_4833, csa_tree_add_6_33_groupi_n_4834, csa_tree_add_6_33_groupi_n_4835, csa_tree_add_6_33_groupi_n_4836, csa_tree_add_6_33_groupi_n_4837;
  wire csa_tree_add_6_33_groupi_n_4839, csa_tree_add_6_33_groupi_n_4840, csa_tree_add_6_33_groupi_n_4842, csa_tree_add_6_33_groupi_n_4843, csa_tree_add_6_33_groupi_n_4844, csa_tree_add_6_33_groupi_n_4846, csa_tree_add_6_33_groupi_n_4847, csa_tree_add_6_33_groupi_n_4849;
  wire csa_tree_add_6_33_groupi_n_4850, csa_tree_add_6_33_groupi_n_4852, csa_tree_add_6_33_groupi_n_4853, csa_tree_add_6_33_groupi_n_4854, csa_tree_add_6_33_groupi_n_4855, csa_tree_add_6_33_groupi_n_4856, csa_tree_add_6_33_groupi_n_4857, csa_tree_add_6_33_groupi_n_4859;
  wire csa_tree_add_6_33_groupi_n_4860, csa_tree_add_6_33_groupi_n_4862, csa_tree_add_6_33_groupi_n_4863, csa_tree_add_6_33_groupi_n_4865, csa_tree_add_6_33_groupi_n_4866, csa_tree_add_6_33_groupi_n_4868, csa_tree_add_6_33_groupi_n_4869, csa_tree_add_6_33_groupi_n_4870;
  wire csa_tree_add_6_33_groupi_n_4871, csa_tree_add_6_33_groupi_n_4873, csa_tree_add_6_33_groupi_n_4874, csa_tree_add_6_33_groupi_n_4875, csa_tree_add_6_33_groupi_n_4877, csa_tree_add_6_33_groupi_n_4878, csa_tree_add_6_33_groupi_n_4880, csa_tree_add_6_33_groupi_n_4881;
  wire csa_tree_add_6_33_groupi_n_4883, csa_tree_add_6_33_groupi_n_4884, csa_tree_add_6_33_groupi_n_4886, csa_tree_add_6_33_groupi_n_4887, csa_tree_add_6_33_groupi_n_4889, csa_tree_add_6_33_groupi_n_4890, csa_tree_add_6_33_groupi_n_4891, csa_tree_add_6_33_groupi_n_4893;
  wire csa_tree_add_6_33_groupi_n_4894, csa_tree_add_6_33_groupi_n_4896, csa_tree_add_6_33_groupi_n_4897, csa_tree_add_6_33_groupi_n_4898, csa_tree_add_6_33_groupi_n_4899, csa_tree_add_6_33_groupi_n_4901, csa_tree_add_6_33_groupi_n_4902, csa_tree_add_6_33_groupi_n_4904;
  wire csa_tree_add_6_33_groupi_n_4905, csa_tree_add_6_33_groupi_n_4907, csa_tree_add_6_33_groupi_n_4908, csa_tree_add_6_33_groupi_n_4909, csa_tree_add_6_33_groupi_n_4911, csa_tree_add_6_33_groupi_n_4912, csa_tree_add_6_33_groupi_n_4914, csa_tree_add_6_33_groupi_n_4915;
  wire csa_tree_add_6_33_groupi_n_4916, csa_tree_add_6_33_groupi_n_4918, csa_tree_add_6_33_groupi_n_4919, csa_tree_add_6_33_groupi_n_4921, csa_tree_add_6_33_groupi_n_4922, csa_tree_add_6_33_groupi_n_4923, csa_tree_add_6_33_groupi_n_4925, csa_tree_add_6_33_groupi_n_4926;
  wire csa_tree_add_6_33_groupi_n_4928, csa_tree_add_6_33_groupi_n_4929, csa_tree_add_6_33_groupi_n_4930, csa_tree_add_6_33_groupi_n_4932, csa_tree_add_6_33_groupi_n_4933, csa_tree_add_6_33_groupi_n_4935, csa_tree_add_6_33_groupi_n_4936, csa_tree_add_6_33_groupi_n_4937;
  wire csa_tree_add_6_33_groupi_n_4939, csa_tree_add_6_33_groupi_n_4940, csa_tree_add_6_33_groupi_n_4942, csa_tree_add_6_33_groupi_n_4943, csa_tree_add_6_33_groupi_n_4944, csa_tree_add_6_33_groupi_n_4945, csa_tree_add_6_33_groupi_n_4947, csa_tree_add_6_33_groupi_n_4948;
  wire csa_tree_add_6_33_groupi_n_4949, csa_tree_add_6_33_groupi_n_4950, csa_tree_add_6_33_groupi_n_4951, csa_tree_add_6_33_groupi_n_4952, csa_tree_add_6_33_groupi_n_4953, csa_tree_add_6_33_groupi_n_4954, csa_tree_add_6_33_groupi_n_4956, csa_tree_add_6_33_groupi_n_4957;
  wire csa_tree_add_6_33_groupi_n_4958, csa_tree_add_6_33_groupi_n_4959, csa_tree_add_6_33_groupi_n_4961, csa_tree_add_6_33_groupi_n_4962, csa_tree_add_6_33_groupi_n_4963, csa_tree_add_6_33_groupi_n_4964;
  buf constbuf_n1(out1[64], 1'b0);
  or csa_tree_add_6_33_groupi_g13304__2398(out1[63] ,csa_tree_add_6_33_groupi_n_1684 ,csa_tree_add_6_33_groupi_n_4964);
  xnor csa_tree_add_6_33_groupi_g13305__5107(out1[62] ,csa_tree_add_6_33_groupi_n_4963 ,csa_tree_add_6_33_groupi_n_2177);
  nor csa_tree_add_6_33_groupi_g13306__6260(csa_tree_add_6_33_groupi_n_4964 ,csa_tree_add_6_33_groupi_n_1883 ,csa_tree_add_6_33_groupi_n_4963);
  and csa_tree_add_6_33_groupi_g13307__4319(csa_tree_add_6_33_groupi_n_4963 ,csa_tree_add_6_33_groupi_n_2838 ,csa_tree_add_6_33_groupi_n_4962);
  or csa_tree_add_6_33_groupi_g13309__8428(csa_tree_add_6_33_groupi_n_4962 ,csa_tree_add_6_33_groupi_n_2824 ,csa_tree_add_6_33_groupi_n_4961);
  and csa_tree_add_6_33_groupi_g13311__5526(csa_tree_add_6_33_groupi_n_4961 ,csa_tree_add_6_33_groupi_n_3301 ,csa_tree_add_6_33_groupi_n_4959);
  xnor csa_tree_add_6_33_groupi_g13312__6783(out1[60] ,csa_tree_add_6_33_groupi_n_4958 ,csa_tree_add_6_33_groupi_n_3395);
  or csa_tree_add_6_33_groupi_g13313__3680(csa_tree_add_6_33_groupi_n_4959 ,csa_tree_add_6_33_groupi_n_3296 ,csa_tree_add_6_33_groupi_n_4958);
  and csa_tree_add_6_33_groupi_g13314__1617(csa_tree_add_6_33_groupi_n_4958 ,csa_tree_add_6_33_groupi_n_3707 ,csa_tree_add_6_33_groupi_n_4957);
  or csa_tree_add_6_33_groupi_g13316__2802(csa_tree_add_6_33_groupi_n_4957 ,csa_tree_add_6_33_groupi_n_3736 ,csa_tree_add_6_33_groupi_n_4956);
  and csa_tree_add_6_33_groupi_g13318__1705(csa_tree_add_6_33_groupi_n_4956 ,csa_tree_add_6_33_groupi_n_3730 ,csa_tree_add_6_33_groupi_n_4954);
  xnor csa_tree_add_6_33_groupi_g13319__5122(out1[58] ,csa_tree_add_6_33_groupi_n_4953 ,csa_tree_add_6_33_groupi_n_3806);
  or csa_tree_add_6_33_groupi_g13320__8246(csa_tree_add_6_33_groupi_n_4954 ,csa_tree_add_6_33_groupi_n_3749 ,csa_tree_add_6_33_groupi_n_4953);
  and csa_tree_add_6_33_groupi_g13321__7098(csa_tree_add_6_33_groupi_n_4953 ,csa_tree_add_6_33_groupi_n_3821 ,csa_tree_add_6_33_groupi_n_4952);
  or csa_tree_add_6_33_groupi_g13323__6131(csa_tree_add_6_33_groupi_n_4952 ,csa_tree_add_6_33_groupi_n_3864 ,csa_tree_add_6_33_groupi_n_4951);
  and csa_tree_add_6_33_groupi_g13325__1881(csa_tree_add_6_33_groupi_n_4951 ,csa_tree_add_6_33_groupi_n_4121 ,csa_tree_add_6_33_groupi_n_4950);
  or csa_tree_add_6_33_groupi_g13327__5115(csa_tree_add_6_33_groupi_n_4950 ,csa_tree_add_6_33_groupi_n_4123 ,csa_tree_add_6_33_groupi_n_4949);
  and csa_tree_add_6_33_groupi_g13329__7482(csa_tree_add_6_33_groupi_n_4949 ,csa_tree_add_6_33_groupi_n_4243 ,csa_tree_add_6_33_groupi_n_4948);
  or csa_tree_add_6_33_groupi_g13331__4733(csa_tree_add_6_33_groupi_n_4948 ,csa_tree_add_6_33_groupi_n_4274 ,csa_tree_add_6_33_groupi_n_4947);
  and csa_tree_add_6_33_groupi_g13333__6161(csa_tree_add_6_33_groupi_n_4947 ,csa_tree_add_6_33_groupi_n_4372 ,csa_tree_add_6_33_groupi_n_4945);
  xnor csa_tree_add_6_33_groupi_g13334__9315(out1[54] ,csa_tree_add_6_33_groupi_n_4944 ,csa_tree_add_6_33_groupi_n_4404);
  or csa_tree_add_6_33_groupi_g13335__9945(csa_tree_add_6_33_groupi_n_4945 ,csa_tree_add_6_33_groupi_n_4351 ,csa_tree_add_6_33_groupi_n_4944);
  and csa_tree_add_6_33_groupi_g13336__2883(csa_tree_add_6_33_groupi_n_4944 ,csa_tree_add_6_33_groupi_n_4350 ,csa_tree_add_6_33_groupi_n_4943);
  or csa_tree_add_6_33_groupi_g13338__2346(csa_tree_add_6_33_groupi_n_4943 ,csa_tree_add_6_33_groupi_n_4321 ,csa_tree_add_6_33_groupi_n_4942);
  and csa_tree_add_6_33_groupi_g13340__1666(csa_tree_add_6_33_groupi_n_4942 ,csa_tree_add_6_33_groupi_n_4441 ,csa_tree_add_6_33_groupi_n_4940);
  xnor csa_tree_add_6_33_groupi_g13341__7410(out1[52] ,csa_tree_add_6_33_groupi_n_4939 ,csa_tree_add_6_33_groupi_n_4480);
  or csa_tree_add_6_33_groupi_g13342__6417(csa_tree_add_6_33_groupi_n_4940 ,csa_tree_add_6_33_groupi_n_4444 ,csa_tree_add_6_33_groupi_n_4939);
  and csa_tree_add_6_33_groupi_g13343__5477(csa_tree_add_6_33_groupi_n_4939 ,csa_tree_add_6_33_groupi_n_4446 ,csa_tree_add_6_33_groupi_n_4937);
  xnor csa_tree_add_6_33_groupi_g13344__2398(out1[51] ,csa_tree_add_6_33_groupi_n_4935 ,csa_tree_add_6_33_groupi_n_4482);
  or csa_tree_add_6_33_groupi_g13345__5107(csa_tree_add_6_33_groupi_n_4937 ,csa_tree_add_6_33_groupi_n_4451 ,csa_tree_add_6_33_groupi_n_4936);
  not csa_tree_add_6_33_groupi_g13346(csa_tree_add_6_33_groupi_n_4936 ,csa_tree_add_6_33_groupi_n_4935);
  or csa_tree_add_6_33_groupi_g13347__6260(csa_tree_add_6_33_groupi_n_4935 ,csa_tree_add_6_33_groupi_n_4933 ,csa_tree_add_6_33_groupi_n_4526);
  xnor csa_tree_add_6_33_groupi_g13348__4319(out1[50] ,csa_tree_add_6_33_groupi_n_4932 ,csa_tree_add_6_33_groupi_n_4551);
  nor csa_tree_add_6_33_groupi_g13349__8428(csa_tree_add_6_33_groupi_n_4933 ,csa_tree_add_6_33_groupi_n_4523 ,csa_tree_add_6_33_groupi_n_4932);
  and csa_tree_add_6_33_groupi_g13350__5526(csa_tree_add_6_33_groupi_n_4932 ,csa_tree_add_6_33_groupi_n_4593 ,csa_tree_add_6_33_groupi_n_4930);
  xnor csa_tree_add_6_33_groupi_g13351__6783(out1[49] ,csa_tree_add_6_33_groupi_n_4928 ,csa_tree_add_6_33_groupi_n_4621);
  or csa_tree_add_6_33_groupi_g13352__3680(csa_tree_add_6_33_groupi_n_4930 ,csa_tree_add_6_33_groupi_n_4586 ,csa_tree_add_6_33_groupi_n_4929);
  not csa_tree_add_6_33_groupi_g13353(csa_tree_add_6_33_groupi_n_4929 ,csa_tree_add_6_33_groupi_n_4928);
  or csa_tree_add_6_33_groupi_g13354__1617(csa_tree_add_6_33_groupi_n_4928 ,csa_tree_add_6_33_groupi_n_4585 ,csa_tree_add_6_33_groupi_n_4926);
  xnor csa_tree_add_6_33_groupi_g13355__2802(out1[48] ,csa_tree_add_6_33_groupi_n_4925 ,csa_tree_add_6_33_groupi_n_4626);
  nor csa_tree_add_6_33_groupi_g13356__1705(csa_tree_add_6_33_groupi_n_4926 ,csa_tree_add_6_33_groupi_n_4591 ,csa_tree_add_6_33_groupi_n_4925);
  and csa_tree_add_6_33_groupi_g13357__5122(csa_tree_add_6_33_groupi_n_4925 ,csa_tree_add_6_33_groupi_n_4642 ,csa_tree_add_6_33_groupi_n_4923);
  xnor csa_tree_add_6_33_groupi_g13358__8246(out1[47] ,csa_tree_add_6_33_groupi_n_4921 ,csa_tree_add_6_33_groupi_n_4682);
  or csa_tree_add_6_33_groupi_g13359__7098(csa_tree_add_6_33_groupi_n_4923 ,csa_tree_add_6_33_groupi_n_4922 ,csa_tree_add_6_33_groupi_n_4651);
  not csa_tree_add_6_33_groupi_g13360(csa_tree_add_6_33_groupi_n_4922 ,csa_tree_add_6_33_groupi_n_4921);
  or csa_tree_add_6_33_groupi_g13361__6131(csa_tree_add_6_33_groupi_n_4921 ,csa_tree_add_6_33_groupi_n_4640 ,csa_tree_add_6_33_groupi_n_4919);
  xnor csa_tree_add_6_33_groupi_g13362__1881(out1[46] ,csa_tree_add_6_33_groupi_n_4918 ,csa_tree_add_6_33_groupi_n_4685);
  nor csa_tree_add_6_33_groupi_g13363__5115(csa_tree_add_6_33_groupi_n_4919 ,csa_tree_add_6_33_groupi_n_4668 ,csa_tree_add_6_33_groupi_n_4918);
  and csa_tree_add_6_33_groupi_g13364__7482(csa_tree_add_6_33_groupi_n_4918 ,csa_tree_add_6_33_groupi_n_4916 ,csa_tree_add_6_33_groupi_n_4652);
  xnor csa_tree_add_6_33_groupi_g13365__4733(out1[45] ,csa_tree_add_6_33_groupi_n_4914 ,csa_tree_add_6_33_groupi_n_4680);
  or csa_tree_add_6_33_groupi_g13366__6161(csa_tree_add_6_33_groupi_n_4916 ,csa_tree_add_6_33_groupi_n_4667 ,csa_tree_add_6_33_groupi_n_4915);
  not csa_tree_add_6_33_groupi_g13367(csa_tree_add_6_33_groupi_n_4915 ,csa_tree_add_6_33_groupi_n_4914);
  or csa_tree_add_6_33_groupi_g13368__9315(csa_tree_add_6_33_groupi_n_4914 ,csa_tree_add_6_33_groupi_n_4662 ,csa_tree_add_6_33_groupi_n_4912);
  xnor csa_tree_add_6_33_groupi_g13369__9945(out1[44] ,csa_tree_add_6_33_groupi_n_4911 ,csa_tree_add_6_33_groupi_n_4679);
  nor csa_tree_add_6_33_groupi_g13370__2883(csa_tree_add_6_33_groupi_n_4912 ,csa_tree_add_6_33_groupi_n_4911 ,csa_tree_add_6_33_groupi_n_4653);
  and csa_tree_add_6_33_groupi_g13371__2346(csa_tree_add_6_33_groupi_n_4911 ,csa_tree_add_6_33_groupi_n_4909 ,csa_tree_add_6_33_groupi_n_4703);
  xnor csa_tree_add_6_33_groupi_g13372__1666(out1[43] ,csa_tree_add_6_33_groupi_n_4907 ,csa_tree_add_6_33_groupi_n_4726);
  or csa_tree_add_6_33_groupi_g13373__7410(csa_tree_add_6_33_groupi_n_4909 ,csa_tree_add_6_33_groupi_n_4705 ,csa_tree_add_6_33_groupi_n_4908);
  not csa_tree_add_6_33_groupi_g13374(csa_tree_add_6_33_groupi_n_4908 ,csa_tree_add_6_33_groupi_n_4907);
  or csa_tree_add_6_33_groupi_g13375__6417(csa_tree_add_6_33_groupi_n_4907 ,csa_tree_add_6_33_groupi_n_4905 ,csa_tree_add_6_33_groupi_n_4746);
  xnor csa_tree_add_6_33_groupi_g13376__5477(out1[42] ,csa_tree_add_6_33_groupi_n_4904 ,csa_tree_add_6_33_groupi_n_4761);
  and csa_tree_add_6_33_groupi_g13377__2398(csa_tree_add_6_33_groupi_n_4905 ,csa_tree_add_6_33_groupi_n_4904 ,csa_tree_add_6_33_groupi_n_4747);
  or csa_tree_add_6_33_groupi_g13378__5107(csa_tree_add_6_33_groupi_n_4904 ,csa_tree_add_6_33_groupi_n_4745 ,csa_tree_add_6_33_groupi_n_4902);
  xnor csa_tree_add_6_33_groupi_g13379__6260(out1[41] ,csa_tree_add_6_33_groupi_n_4901 ,csa_tree_add_6_33_groupi_n_4764);
  nor csa_tree_add_6_33_groupi_g13380__4319(csa_tree_add_6_33_groupi_n_4902 ,csa_tree_add_6_33_groupi_n_4901 ,csa_tree_add_6_33_groupi_n_4748);
  and csa_tree_add_6_33_groupi_g13381__8428(csa_tree_add_6_33_groupi_n_4901 ,csa_tree_add_6_33_groupi_n_4899 ,csa_tree_add_6_33_groupi_n_4781);
  xnor csa_tree_add_6_33_groupi_g13382__5526(out1[40] ,csa_tree_add_6_33_groupi_n_4898 ,csa_tree_add_6_33_groupi_n_4790);
  or csa_tree_add_6_33_groupi_g13383__6783(csa_tree_add_6_33_groupi_n_4899 ,csa_tree_add_6_33_groupi_n_4898 ,csa_tree_add_6_33_groupi_n_4782);
  and csa_tree_add_6_33_groupi_g13384__3680(csa_tree_add_6_33_groupi_n_4898 ,csa_tree_add_6_33_groupi_n_4777 ,csa_tree_add_6_33_groupi_n_4897);
  or csa_tree_add_6_33_groupi_g13386__1617(csa_tree_add_6_33_groupi_n_4897 ,csa_tree_add_6_33_groupi_n_4788 ,csa_tree_add_6_33_groupi_n_4896);
  and csa_tree_add_6_33_groupi_g13388__2802(csa_tree_add_6_33_groupi_n_4896 ,csa_tree_add_6_33_groupi_n_4787 ,csa_tree_add_6_33_groupi_n_4894);
  xnor csa_tree_add_6_33_groupi_g13389__1705(out1[38] ,csa_tree_add_6_33_groupi_n_4893 ,csa_tree_add_6_33_groupi_n_4795);
  or csa_tree_add_6_33_groupi_g13390__5122(csa_tree_add_6_33_groupi_n_4894 ,csa_tree_add_6_33_groupi_n_4786 ,csa_tree_add_6_33_groupi_n_4893);
  and csa_tree_add_6_33_groupi_g13391__8246(csa_tree_add_6_33_groupi_n_4893 ,csa_tree_add_6_33_groupi_n_4891 ,csa_tree_add_6_33_groupi_n_4783);
  xnor csa_tree_add_6_33_groupi_g13392__7098(out1[37] ,csa_tree_add_6_33_groupi_n_4889 ,csa_tree_add_6_33_groupi_n_4791);
  or csa_tree_add_6_33_groupi_g13393__6131(csa_tree_add_6_33_groupi_n_4891 ,csa_tree_add_6_33_groupi_n_4785 ,csa_tree_add_6_33_groupi_n_4890);
  not csa_tree_add_6_33_groupi_g13394(csa_tree_add_6_33_groupi_n_4890 ,csa_tree_add_6_33_groupi_n_4889);
  or csa_tree_add_6_33_groupi_g13395__1881(csa_tree_add_6_33_groupi_n_4889 ,csa_tree_add_6_33_groupi_n_4800 ,csa_tree_add_6_33_groupi_n_4887);
  xnor csa_tree_add_6_33_groupi_g13396__5115(out1[36] ,csa_tree_add_6_33_groupi_n_4886 ,csa_tree_add_6_33_groupi_n_4815);
  nor csa_tree_add_6_33_groupi_g13397__7482(csa_tree_add_6_33_groupi_n_4887 ,csa_tree_add_6_33_groupi_n_4886 ,csa_tree_add_6_33_groupi_n_4804);
  and csa_tree_add_6_33_groupi_g13398__4733(csa_tree_add_6_33_groupi_n_4886 ,csa_tree_add_6_33_groupi_n_4884 ,csa_tree_add_6_33_groupi_n_4805);
  xnor csa_tree_add_6_33_groupi_g13399__6161(out1[35] ,csa_tree_add_6_33_groupi_n_4883 ,csa_tree_add_6_33_groupi_n_4813);
  or csa_tree_add_6_33_groupi_g13400__9315(csa_tree_add_6_33_groupi_n_4884 ,csa_tree_add_6_33_groupi_n_4883 ,csa_tree_add_6_33_groupi_n_4806);
  and csa_tree_add_6_33_groupi_g13401__9945(csa_tree_add_6_33_groupi_n_4883 ,csa_tree_add_6_33_groupi_n_4881 ,csa_tree_add_6_33_groupi_n_4802);
  xnor csa_tree_add_6_33_groupi_g13402__2883(out1[34] ,csa_tree_add_6_33_groupi_n_4880 ,csa_tree_add_6_33_groupi_n_4814);
  or csa_tree_add_6_33_groupi_g13403__2346(csa_tree_add_6_33_groupi_n_4881 ,csa_tree_add_6_33_groupi_n_4880 ,csa_tree_add_6_33_groupi_n_4803);
  and csa_tree_add_6_33_groupi_g13404__1666(csa_tree_add_6_33_groupi_n_4880 ,csa_tree_add_6_33_groupi_n_4878 ,csa_tree_add_6_33_groupi_n_4797);
  xnor csa_tree_add_6_33_groupi_g13405__7410(out1[33] ,csa_tree_add_6_33_groupi_n_4877 ,csa_tree_add_6_33_groupi_n_4812);
  or csa_tree_add_6_33_groupi_g13406__6417(csa_tree_add_6_33_groupi_n_4878 ,csa_tree_add_6_33_groupi_n_4877 ,csa_tree_add_6_33_groupi_n_4798);
  and csa_tree_add_6_33_groupi_g13407__5477(csa_tree_add_6_33_groupi_n_4877 ,csa_tree_add_6_33_groupi_n_4807 ,csa_tree_add_6_33_groupi_n_4875);
  xnor csa_tree_add_6_33_groupi_g13408__2398(out1[32] ,csa_tree_add_6_33_groupi_n_4873 ,csa_tree_add_6_33_groupi_n_4811);
  or csa_tree_add_6_33_groupi_g13409__5107(csa_tree_add_6_33_groupi_n_4875 ,csa_tree_add_6_33_groupi_n_4801 ,csa_tree_add_6_33_groupi_n_4874);
  not csa_tree_add_6_33_groupi_g13410(csa_tree_add_6_33_groupi_n_4874 ,csa_tree_add_6_33_groupi_n_4873);
  or csa_tree_add_6_33_groupi_g13411__6260(csa_tree_add_6_33_groupi_n_4873 ,csa_tree_add_6_33_groupi_n_4780 ,csa_tree_add_6_33_groupi_n_4871);
  xnor csa_tree_add_6_33_groupi_g13412__4319(out1[31] ,csa_tree_add_6_33_groupi_n_4870 ,csa_tree_add_6_33_groupi_n_4794);
  nor csa_tree_add_6_33_groupi_g13413__8428(csa_tree_add_6_33_groupi_n_4871 ,csa_tree_add_6_33_groupi_n_4870 ,csa_tree_add_6_33_groupi_n_4784);
  and csa_tree_add_6_33_groupi_g13414__5526(csa_tree_add_6_33_groupi_n_4870 ,csa_tree_add_6_33_groupi_n_4796 ,csa_tree_add_6_33_groupi_n_4869);
  or csa_tree_add_6_33_groupi_g13416__6783(csa_tree_add_6_33_groupi_n_4869 ,csa_tree_add_6_33_groupi_n_4868 ,csa_tree_add_6_33_groupi_n_4799);
  and csa_tree_add_6_33_groupi_g13418__3680(csa_tree_add_6_33_groupi_n_4868 ,csa_tree_add_6_33_groupi_n_4779 ,csa_tree_add_6_33_groupi_n_4866);
  xnor csa_tree_add_6_33_groupi_g13419__1617(out1[29] ,csa_tree_add_6_33_groupi_n_4865 ,csa_tree_add_6_33_groupi_n_4793);
  or csa_tree_add_6_33_groupi_g13420__2802(csa_tree_add_6_33_groupi_n_4866 ,csa_tree_add_6_33_groupi_n_4778 ,csa_tree_add_6_33_groupi_n_4865);
  and csa_tree_add_6_33_groupi_g13421__1705(csa_tree_add_6_33_groupi_n_4865 ,csa_tree_add_6_33_groupi_n_4863 ,csa_tree_add_6_33_groupi_n_4749);
  xnor csa_tree_add_6_33_groupi_g13422__5122(out1[28] ,csa_tree_add_6_33_groupi_n_4862 ,csa_tree_add_6_33_groupi_n_4763);
  or csa_tree_add_6_33_groupi_g13423__8246(csa_tree_add_6_33_groupi_n_4863 ,csa_tree_add_6_33_groupi_n_4862 ,csa_tree_add_6_33_groupi_n_4750);
  and csa_tree_add_6_33_groupi_g13424__7098(csa_tree_add_6_33_groupi_n_4862 ,csa_tree_add_6_33_groupi_n_4752 ,csa_tree_add_6_33_groupi_n_4860);
  xnor csa_tree_add_6_33_groupi_g13425__6131(out1[27] ,csa_tree_add_6_33_groupi_n_4859 ,csa_tree_add_6_33_groupi_n_4762);
  or csa_tree_add_6_33_groupi_g13426__1881(csa_tree_add_6_33_groupi_n_4860 ,csa_tree_add_6_33_groupi_n_4859 ,csa_tree_add_6_33_groupi_n_4751);
  and csa_tree_add_6_33_groupi_g13427__5115(csa_tree_add_6_33_groupi_n_4859 ,csa_tree_add_6_33_groupi_n_4857 ,csa_tree_add_6_33_groupi_n_4729);
  xnor csa_tree_add_6_33_groupi_g13428__7482(out1[26] ,csa_tree_add_6_33_groupi_n_4856 ,csa_tree_add_6_33_groupi_n_4758);
  or csa_tree_add_6_33_groupi_g13429__4733(csa_tree_add_6_33_groupi_n_4857 ,csa_tree_add_6_33_groupi_n_4856 ,csa_tree_add_6_33_groupi_n_4730);
  and csa_tree_add_6_33_groupi_g13430__6161(csa_tree_add_6_33_groupi_n_4856 ,csa_tree_add_6_33_groupi_n_4855 ,csa_tree_add_6_33_groupi_n_4744);
  or csa_tree_add_6_33_groupi_g13432__9315(csa_tree_add_6_33_groupi_n_4855 ,csa_tree_add_6_33_groupi_n_4732 ,csa_tree_add_6_33_groupi_n_4854);
  and csa_tree_add_6_33_groupi_g13434__9945(csa_tree_add_6_33_groupi_n_4854 ,csa_tree_add_6_33_groupi_n_4853 ,csa_tree_add_6_33_groupi_n_4731);
  or csa_tree_add_6_33_groupi_g13436__2883(csa_tree_add_6_33_groupi_n_4853 ,csa_tree_add_6_33_groupi_n_4728 ,csa_tree_add_6_33_groupi_n_4852);
  and csa_tree_add_6_33_groupi_g13438__2346(csa_tree_add_6_33_groupi_n_4852 ,csa_tree_add_6_33_groupi_n_4638 ,csa_tree_add_6_33_groupi_n_4850);
  xnor csa_tree_add_6_33_groupi_g13439__1666(out1[23] ,csa_tree_add_6_33_groupi_n_4849 ,csa_tree_add_6_33_groupi_n_4677);
  or csa_tree_add_6_33_groupi_g13440__7410(csa_tree_add_6_33_groupi_n_4850 ,csa_tree_add_6_33_groupi_n_4849 ,csa_tree_add_6_33_groupi_n_4631);
  and csa_tree_add_6_33_groupi_g13441__6417(csa_tree_add_6_33_groupi_n_4849 ,csa_tree_add_6_33_groupi_n_4637 ,csa_tree_add_6_33_groupi_n_4847);
  xnor csa_tree_add_6_33_groupi_g13442__5477(out1[22] ,csa_tree_add_6_33_groupi_n_4846 ,csa_tree_add_6_33_groupi_n_4676);
  or csa_tree_add_6_33_groupi_g13443__2398(csa_tree_add_6_33_groupi_n_4847 ,csa_tree_add_6_33_groupi_n_4636 ,csa_tree_add_6_33_groupi_n_4846);
  and csa_tree_add_6_33_groupi_g13444__5107(csa_tree_add_6_33_groupi_n_4846 ,csa_tree_add_6_33_groupi_n_4844 ,csa_tree_add_6_33_groupi_n_4632);
  xnor csa_tree_add_6_33_groupi_g13445__6260(out1[21] ,csa_tree_add_6_33_groupi_n_4842 ,csa_tree_add_6_33_groupi_n_4675);
  or csa_tree_add_6_33_groupi_g13446__4319(csa_tree_add_6_33_groupi_n_4844 ,csa_tree_add_6_33_groupi_n_4635 ,csa_tree_add_6_33_groupi_n_4843);
  not csa_tree_add_6_33_groupi_g13447(csa_tree_add_6_33_groupi_n_4843 ,csa_tree_add_6_33_groupi_n_4842);
  or csa_tree_add_6_33_groupi_g13448__8428(csa_tree_add_6_33_groupi_n_4842 ,csa_tree_add_6_33_groupi_n_4669 ,csa_tree_add_6_33_groupi_n_4840);
  xnor csa_tree_add_6_33_groupi_g13449__5526(out1[20] ,csa_tree_add_6_33_groupi_n_4839 ,csa_tree_add_6_33_groupi_n_4674);
  nor csa_tree_add_6_33_groupi_g13450__6783(csa_tree_add_6_33_groupi_n_4840 ,csa_tree_add_6_33_groupi_n_4665 ,csa_tree_add_6_33_groupi_n_4839);
  and csa_tree_add_6_33_groupi_g13451__3680(csa_tree_add_6_33_groupi_n_4839 ,csa_tree_add_6_33_groupi_n_4603 ,csa_tree_add_6_33_groupi_n_4837);
  xnor csa_tree_add_6_33_groupi_g13452__1617(out1[19] ,csa_tree_add_6_33_groupi_n_4836 ,csa_tree_add_6_33_groupi_n_4625);
  or csa_tree_add_6_33_groupi_g13453__2802(csa_tree_add_6_33_groupi_n_4837 ,csa_tree_add_6_33_groupi_n_4836 ,csa_tree_add_6_33_groupi_n_4598);
  and csa_tree_add_6_33_groupi_g13454__1705(csa_tree_add_6_33_groupi_n_4836 ,csa_tree_add_6_33_groupi_n_4634 ,csa_tree_add_6_33_groupi_n_4835);
  or csa_tree_add_6_33_groupi_g13456__5122(csa_tree_add_6_33_groupi_n_4835 ,csa_tree_add_6_33_groupi_n_4633 ,csa_tree_add_6_33_groupi_n_4834);
  and csa_tree_add_6_33_groupi_g13458__8246(csa_tree_add_6_33_groupi_n_4834 ,csa_tree_add_6_33_groupi_n_4485 ,csa_tree_add_6_33_groupi_n_4833);
  or csa_tree_add_6_33_groupi_g13460__7098(csa_tree_add_6_33_groupi_n_4833 ,csa_tree_add_6_33_groupi_n_4489 ,csa_tree_add_6_33_groupi_n_4832);
  and csa_tree_add_6_33_groupi_g13462__6131(csa_tree_add_6_33_groupi_n_4832 ,csa_tree_add_6_33_groupi_n_4521 ,csa_tree_add_6_33_groupi_n_4831);
  or csa_tree_add_6_33_groupi_g13464__1881(csa_tree_add_6_33_groupi_n_4831 ,csa_tree_add_6_33_groupi_n_4520 ,csa_tree_add_6_33_groupi_n_4830);
  and csa_tree_add_6_33_groupi_g13466__5115(csa_tree_add_6_33_groupi_n_4830 ,csa_tree_add_6_33_groupi_n_4519 ,csa_tree_add_6_33_groupi_n_4829);
  or csa_tree_add_6_33_groupi_g13468__7482(csa_tree_add_6_33_groupi_n_4829 ,csa_tree_add_6_33_groupi_n_4518 ,csa_tree_add_6_33_groupi_n_4828);
  and csa_tree_add_6_33_groupi_g13470__4733(csa_tree_add_6_33_groupi_n_4828 ,csa_tree_add_6_33_groupi_n_4361 ,csa_tree_add_6_33_groupi_n_4827);
  or csa_tree_add_6_33_groupi_g13472__6161(csa_tree_add_6_33_groupi_n_4827 ,csa_tree_add_6_33_groupi_n_4358 ,csa_tree_add_6_33_groupi_n_4826);
  and csa_tree_add_6_33_groupi_g13474__9315(csa_tree_add_6_33_groupi_n_4826 ,csa_tree_add_6_33_groupi_n_4357 ,csa_tree_add_6_33_groupi_n_4824);
  xnor csa_tree_add_6_33_groupi_g13475__9945(out1[13] ,csa_tree_add_6_33_groupi_n_4822 ,csa_tree_add_6_33_groupi_n_4389);
  or csa_tree_add_6_33_groupi_g13476__2883(csa_tree_add_6_33_groupi_n_4824 ,csa_tree_add_6_33_groupi_n_4356 ,csa_tree_add_6_33_groupi_n_4823);
  not csa_tree_add_6_33_groupi_g13477(csa_tree_add_6_33_groupi_n_4823 ,csa_tree_add_6_33_groupi_n_4822);
  or csa_tree_add_6_33_groupi_g13478__2346(csa_tree_add_6_33_groupi_n_4822 ,csa_tree_add_6_33_groupi_n_4318 ,csa_tree_add_6_33_groupi_n_4820);
  xnor csa_tree_add_6_33_groupi_g13479__1666(out1[12] ,csa_tree_add_6_33_groupi_n_4819 ,csa_tree_add_6_33_groupi_n_4388);
  and csa_tree_add_6_33_groupi_g13480__7410(csa_tree_add_6_33_groupi_n_4820 ,csa_tree_add_6_33_groupi_n_4320 ,csa_tree_add_6_33_groupi_n_4819);
  or csa_tree_add_6_33_groupi_g13481__6417(csa_tree_add_6_33_groupi_n_4819 ,csa_tree_add_6_33_groupi_n_4055 ,csa_tree_add_6_33_groupi_n_4817);
  xnor csa_tree_add_6_33_groupi_g13482__5477(out1[11] ,csa_tree_add_6_33_groupi_n_4816 ,csa_tree_add_6_33_groupi_n_4182);
  and csa_tree_add_6_33_groupi_g13483__2398(csa_tree_add_6_33_groupi_n_4817 ,csa_tree_add_6_33_groupi_n_4054 ,csa_tree_add_6_33_groupi_n_4816);
  or csa_tree_add_6_33_groupi_g13484__5107(csa_tree_add_6_33_groupi_n_4816 ,csa_tree_add_6_33_groupi_n_4053 ,csa_tree_add_6_33_groupi_n_4808);
  xnor csa_tree_add_6_33_groupi_g13485__6260(csa_tree_add_6_33_groupi_n_4815 ,csa_tree_add_6_33_groupi_n_4766 ,csa_tree_add_6_33_groupi_n_4753);
  xnor csa_tree_add_6_33_groupi_g13486__4319(csa_tree_add_6_33_groupi_n_4814 ,csa_tree_add_6_33_groupi_n_4774 ,csa_tree_add_6_33_groupi_n_4724);
  xnor csa_tree_add_6_33_groupi_g13487__8428(csa_tree_add_6_33_groupi_n_4813 ,csa_tree_add_6_33_groupi_n_4776 ,csa_tree_add_6_33_groupi_n_4757);
  xnor csa_tree_add_6_33_groupi_g13488__5526(csa_tree_add_6_33_groupi_n_4812 ,csa_tree_add_6_33_groupi_n_4771 ,csa_tree_add_6_33_groupi_n_4739);
  xnor csa_tree_add_6_33_groupi_g13489__6783(csa_tree_add_6_33_groupi_n_4811 ,csa_tree_add_6_33_groupi_n_4755 ,csa_tree_add_6_33_groupi_n_4772);
  xnor csa_tree_add_6_33_groupi_g13490__3680(csa_tree_add_6_33_groupi_n_4810 ,csa_tree_add_6_33_groupi_n_4769 ,csa_tree_add_6_33_groupi_n_4721);
  xnor csa_tree_add_6_33_groupi_g13491__1617(out1[10] ,csa_tree_add_6_33_groupi_n_4789 ,csa_tree_add_6_33_groupi_n_4181);
  and csa_tree_add_6_33_groupi_g13492__2802(csa_tree_add_6_33_groupi_n_4808 ,csa_tree_add_6_33_groupi_n_4052 ,csa_tree_add_6_33_groupi_n_4789);
  or csa_tree_add_6_33_groupi_g13493__1705(csa_tree_add_6_33_groupi_n_4807 ,csa_tree_add_6_33_groupi_n_4772 ,csa_tree_add_6_33_groupi_n_4755);
  nor csa_tree_add_6_33_groupi_g13494__5122(csa_tree_add_6_33_groupi_n_4806 ,csa_tree_add_6_33_groupi_n_4775 ,csa_tree_add_6_33_groupi_n_4757);
  or csa_tree_add_6_33_groupi_g13495__8246(csa_tree_add_6_33_groupi_n_4805 ,csa_tree_add_6_33_groupi_n_4776 ,csa_tree_add_6_33_groupi_n_4756);
  and csa_tree_add_6_33_groupi_g13496__7098(csa_tree_add_6_33_groupi_n_4804 ,csa_tree_add_6_33_groupi_n_4767 ,csa_tree_add_6_33_groupi_n_4753);
  nor csa_tree_add_6_33_groupi_g13497__6131(csa_tree_add_6_33_groupi_n_4803 ,csa_tree_add_6_33_groupi_n_4774 ,csa_tree_add_6_33_groupi_n_4723);
  or csa_tree_add_6_33_groupi_g13498__1881(csa_tree_add_6_33_groupi_n_4802 ,csa_tree_add_6_33_groupi_n_4773 ,csa_tree_add_6_33_groupi_n_4724);
  and csa_tree_add_6_33_groupi_g13499__5115(csa_tree_add_6_33_groupi_n_4801 ,csa_tree_add_6_33_groupi_n_4772 ,csa_tree_add_6_33_groupi_n_4755);
  nor csa_tree_add_6_33_groupi_g13500__7482(csa_tree_add_6_33_groupi_n_4800 ,csa_tree_add_6_33_groupi_n_4767 ,csa_tree_add_6_33_groupi_n_4753);
  nor csa_tree_add_6_33_groupi_g13501__4733(csa_tree_add_6_33_groupi_n_4799 ,csa_tree_add_6_33_groupi_n_4769 ,csa_tree_add_6_33_groupi_n_4721);
  nor csa_tree_add_6_33_groupi_g13502__6161(csa_tree_add_6_33_groupi_n_4798 ,csa_tree_add_6_33_groupi_n_4770 ,csa_tree_add_6_33_groupi_n_4739);
  or csa_tree_add_6_33_groupi_g13503__9315(csa_tree_add_6_33_groupi_n_4797 ,csa_tree_add_6_33_groupi_n_4771 ,csa_tree_add_6_33_groupi_n_4738);
  or csa_tree_add_6_33_groupi_g13504__9945(csa_tree_add_6_33_groupi_n_4796 ,csa_tree_add_6_33_groupi_n_4768 ,csa_tree_add_6_33_groupi_n_4720);
  xnor csa_tree_add_6_33_groupi_g13505__2883(csa_tree_add_6_33_groupi_n_4795 ,csa_tree_add_6_33_groupi_n_4716 ,csa_tree_add_6_33_groupi_n_4743);
  xnor csa_tree_add_6_33_groupi_g13506__2346(csa_tree_add_6_33_groupi_n_4794 ,csa_tree_add_6_33_groupi_n_4736 ,csa_tree_add_6_33_groupi_n_4722);
  xnor csa_tree_add_6_33_groupi_g13507__1666(csa_tree_add_6_33_groupi_n_4793 ,csa_tree_add_6_33_groupi_n_4719 ,csa_tree_add_6_33_groupi_n_4735);
  xnor csa_tree_add_6_33_groupi_g13508__7410(csa_tree_add_6_33_groupi_n_4792 ,csa_tree_add_6_33_groupi_n_4734 ,csa_tree_add_6_33_groupi_n_4717);
  xnor csa_tree_add_6_33_groupi_g13509__6417(csa_tree_add_6_33_groupi_n_4791 ,csa_tree_add_6_33_groupi_n_4733 ,csa_tree_add_6_33_groupi_n_4754);
  xnor csa_tree_add_6_33_groupi_g13510__5477(csa_tree_add_6_33_groupi_n_4790 ,csa_tree_add_6_33_groupi_n_4712 ,csa_tree_add_6_33_groupi_n_4741);
  and csa_tree_add_6_33_groupi_g13511__2398(csa_tree_add_6_33_groupi_n_4788 ,csa_tree_add_6_33_groupi_n_4717 ,csa_tree_add_6_33_groupi_n_4734);
  or csa_tree_add_6_33_groupi_g13512__5107(csa_tree_add_6_33_groupi_n_4787 ,csa_tree_add_6_33_groupi_n_4716 ,csa_tree_add_6_33_groupi_n_4742);
  nor csa_tree_add_6_33_groupi_g13513__6260(csa_tree_add_6_33_groupi_n_4786 ,csa_tree_add_6_33_groupi_n_4715 ,csa_tree_add_6_33_groupi_n_4743);
  and csa_tree_add_6_33_groupi_g13514__4319(csa_tree_add_6_33_groupi_n_4785 ,csa_tree_add_6_33_groupi_n_4754 ,csa_tree_add_6_33_groupi_n_4733);
  and csa_tree_add_6_33_groupi_g13515__8428(csa_tree_add_6_33_groupi_n_4784 ,csa_tree_add_6_33_groupi_n_4737 ,csa_tree_add_6_33_groupi_n_4722);
  or csa_tree_add_6_33_groupi_g13516__5526(csa_tree_add_6_33_groupi_n_4783 ,csa_tree_add_6_33_groupi_n_4754 ,csa_tree_add_6_33_groupi_n_4733);
  nor csa_tree_add_6_33_groupi_g13517__6783(csa_tree_add_6_33_groupi_n_4782 ,csa_tree_add_6_33_groupi_n_4711 ,csa_tree_add_6_33_groupi_n_4741);
  or csa_tree_add_6_33_groupi_g13518__3680(csa_tree_add_6_33_groupi_n_4781 ,csa_tree_add_6_33_groupi_n_4712 ,csa_tree_add_6_33_groupi_n_4740);
  nor csa_tree_add_6_33_groupi_g13519__1617(csa_tree_add_6_33_groupi_n_4780 ,csa_tree_add_6_33_groupi_n_4737 ,csa_tree_add_6_33_groupi_n_4722);
  or csa_tree_add_6_33_groupi_g13520__2802(csa_tree_add_6_33_groupi_n_4779 ,csa_tree_add_6_33_groupi_n_4719 ,csa_tree_add_6_33_groupi_n_1);
  nor csa_tree_add_6_33_groupi_g13521__1705(csa_tree_add_6_33_groupi_n_4778 ,csa_tree_add_6_33_groupi_n_4718 ,csa_tree_add_6_33_groupi_n_4735);
  or csa_tree_add_6_33_groupi_g13522__5122(csa_tree_add_6_33_groupi_n_4777 ,csa_tree_add_6_33_groupi_n_4717 ,csa_tree_add_6_33_groupi_n_4734);
  or csa_tree_add_6_33_groupi_g13523__8246(csa_tree_add_6_33_groupi_n_4789 ,csa_tree_add_6_33_groupi_n_4061 ,csa_tree_add_6_33_groupi_n_4727);
  not csa_tree_add_6_33_groupi_g13524(csa_tree_add_6_33_groupi_n_4775 ,csa_tree_add_6_33_groupi_n_4776);
  not csa_tree_add_6_33_groupi_g13525(csa_tree_add_6_33_groupi_n_4773 ,csa_tree_add_6_33_groupi_n_4774);
  not csa_tree_add_6_33_groupi_g13526(csa_tree_add_6_33_groupi_n_4771 ,csa_tree_add_6_33_groupi_n_4770);
  not csa_tree_add_6_33_groupi_g13527(csa_tree_add_6_33_groupi_n_4769 ,csa_tree_add_6_33_groupi_n_4768);
  not csa_tree_add_6_33_groupi_g13528(csa_tree_add_6_33_groupi_n_4767 ,csa_tree_add_6_33_groupi_n_4766);
  xnor csa_tree_add_6_33_groupi_g13529__7098(out1[9] ,csa_tree_add_6_33_groupi_n_4725 ,csa_tree_add_6_33_groupi_n_4180);
  xnor csa_tree_add_6_33_groupi_g13530__6131(csa_tree_add_6_33_groupi_n_4764 ,csa_tree_add_6_33_groupi_n_4708 ,csa_tree_add_6_33_groupi_n_4695);
  xnor csa_tree_add_6_33_groupi_g13531__1881(csa_tree_add_6_33_groupi_n_4763 ,csa_tree_add_6_33_groupi_n_4710 ,csa_tree_add_6_33_groupi_n_4688);
  xnor csa_tree_add_6_33_groupi_g13532__5115(csa_tree_add_6_33_groupi_n_4762 ,csa_tree_add_6_33_groupi_n_4645 ,csa_tree_add_6_33_groupi_n_4694);
  xnor csa_tree_add_6_33_groupi_g13533__7482(csa_tree_add_6_33_groupi_n_4761 ,csa_tree_add_6_33_groupi_n_4672 ,csa_tree_add_6_33_groupi_n_4689);
  xnor csa_tree_add_6_33_groupi_g13534__4733(csa_tree_add_6_33_groupi_n_4760 ,csa_tree_add_6_33_groupi_n_4692 ,csa_tree_add_6_33_groupi_n_4643);
  xnor csa_tree_add_6_33_groupi_g13535__6161(csa_tree_add_6_33_groupi_n_4759 ,csa_tree_add_6_33_groupi_n_4612 ,csa_tree_add_6_33_groupi_n_4698);
  xnor csa_tree_add_6_33_groupi_g13536__9315(csa_tree_add_6_33_groupi_n_4758 ,csa_tree_add_6_33_groupi_n_4714 ,csa_tree_add_6_33_groupi_n_4691);
  xnor csa_tree_add_6_33_groupi_g13537__9945(csa_tree_add_6_33_groupi_n_4776 ,csa_tree_add_6_33_groupi_n_4617 ,csa_tree_add_6_33_groupi_n_4684);
  xnor csa_tree_add_6_33_groupi_g13538__2883(csa_tree_add_6_33_groupi_n_4774 ,csa_tree_add_6_33_groupi_n_4610 ,csa_tree_add_6_33_groupi_n_4699);
  xnor csa_tree_add_6_33_groupi_g13539__2346(csa_tree_add_6_33_groupi_n_4772 ,csa_tree_add_6_33_groupi_n_4608 ,csa_tree_add_6_33_groupi_n_4678);
  xnor csa_tree_add_6_33_groupi_g13540__1666(csa_tree_add_6_33_groupi_n_4770 ,csa_tree_add_6_33_groupi_n_4501 ,csa_tree_add_6_33_groupi_n_4681);
  xnor csa_tree_add_6_33_groupi_g13541__7410(csa_tree_add_6_33_groupi_n_4768 ,csa_tree_add_6_33_groupi_n_4494 ,csa_tree_add_6_33_groupi_n_4683);
  xnor csa_tree_add_6_33_groupi_g13542__6417(csa_tree_add_6_33_groupi_n_4766 ,csa_tree_add_6_33_groupi_n_4616 ,csa_tree_add_6_33_groupi_n_4700);
  not csa_tree_add_6_33_groupi_g13543(csa_tree_add_6_33_groupi_n_4756 ,csa_tree_add_6_33_groupi_n_4757);
  or csa_tree_add_6_33_groupi_g13544__5477(csa_tree_add_6_33_groupi_n_4752 ,csa_tree_add_6_33_groupi_n_4645 ,csa_tree_add_6_33_groupi_n_4693);
  nor csa_tree_add_6_33_groupi_g13545__2398(csa_tree_add_6_33_groupi_n_4751 ,csa_tree_add_6_33_groupi_n_4644 ,csa_tree_add_6_33_groupi_n_4694);
  nor csa_tree_add_6_33_groupi_g13546__5107(csa_tree_add_6_33_groupi_n_4750 ,csa_tree_add_6_33_groupi_n_4709 ,csa_tree_add_6_33_groupi_n_4688);
  or csa_tree_add_6_33_groupi_g13547__6260(csa_tree_add_6_33_groupi_n_4749 ,csa_tree_add_6_33_groupi_n_4710 ,csa_tree_add_6_33_groupi_n_4687);
  and csa_tree_add_6_33_groupi_g13548__4319(csa_tree_add_6_33_groupi_n_4748 ,csa_tree_add_6_33_groupi_n_4708 ,csa_tree_add_6_33_groupi_n_4696);
  or csa_tree_add_6_33_groupi_g13549__8428(csa_tree_add_6_33_groupi_n_4747 ,csa_tree_add_6_33_groupi_n_4672 ,csa_tree_add_6_33_groupi_n_4689);
  and csa_tree_add_6_33_groupi_g13550__5526(csa_tree_add_6_33_groupi_n_4746 ,csa_tree_add_6_33_groupi_n_4672 ,csa_tree_add_6_33_groupi_n_4689);
  nor csa_tree_add_6_33_groupi_g13551__6783(csa_tree_add_6_33_groupi_n_4745 ,csa_tree_add_6_33_groupi_n_4708 ,csa_tree_add_6_33_groupi_n_4696);
  or csa_tree_add_6_33_groupi_g13552__3680(csa_tree_add_6_33_groupi_n_4744 ,csa_tree_add_6_33_groupi_n_4643 ,csa_tree_add_6_33_groupi_n_4692);
  or csa_tree_add_6_33_groupi_g13553__1617(csa_tree_add_6_33_groupi_n_4757 ,csa_tree_add_6_33_groupi_n_4670 ,csa_tree_add_6_33_groupi_n_4704);
  and csa_tree_add_6_33_groupi_g13554__2802(csa_tree_add_6_33_groupi_n_4755 ,csa_tree_add_6_33_groupi_n_4650 ,csa_tree_add_6_33_groupi_n_4702);
  and csa_tree_add_6_33_groupi_g13555__1705(csa_tree_add_6_33_groupi_n_4754 ,csa_tree_add_6_33_groupi_n_4666 ,csa_tree_add_6_33_groupi_n_4707);
  and csa_tree_add_6_33_groupi_g13556__5122(csa_tree_add_6_33_groupi_n_4753 ,csa_tree_add_6_33_groupi_n_4663 ,csa_tree_add_6_33_groupi_n_4706);
  not csa_tree_add_6_33_groupi_g13557(csa_tree_add_6_33_groupi_n_4742 ,csa_tree_add_6_33_groupi_n_4743);
  not csa_tree_add_6_33_groupi_g13558(csa_tree_add_6_33_groupi_n_4740 ,csa_tree_add_6_33_groupi_n_4741);
  not csa_tree_add_6_33_groupi_g13559(csa_tree_add_6_33_groupi_n_4738 ,csa_tree_add_6_33_groupi_n_4739);
  not csa_tree_add_6_33_groupi_g13560(csa_tree_add_6_33_groupi_n_4737 ,csa_tree_add_6_33_groupi_n_4736);
  not csa_tree_add_6_33_groupi_g13561(csa_tree_add_6_33_groupi_n_4735 ,csa_tree_add_6_33_groupi_n_1);
  and csa_tree_add_6_33_groupi_g13562__8246(csa_tree_add_6_33_groupi_n_4732 ,csa_tree_add_6_33_groupi_n_4643 ,csa_tree_add_6_33_groupi_n_4692);
  or csa_tree_add_6_33_groupi_g13563__7098(csa_tree_add_6_33_groupi_n_4731 ,csa_tree_add_6_33_groupi_n_4611 ,csa_tree_add_6_33_groupi_n_4697);
  nor csa_tree_add_6_33_groupi_g13564__6131(csa_tree_add_6_33_groupi_n_4730 ,csa_tree_add_6_33_groupi_n_4713 ,csa_tree_add_6_33_groupi_n_4691);
  or csa_tree_add_6_33_groupi_g13565__1881(csa_tree_add_6_33_groupi_n_4729 ,csa_tree_add_6_33_groupi_n_4714 ,csa_tree_add_6_33_groupi_n_4690);
  nor csa_tree_add_6_33_groupi_g13566__5115(csa_tree_add_6_33_groupi_n_4728 ,csa_tree_add_6_33_groupi_n_4612 ,csa_tree_add_6_33_groupi_n_4698);
  and csa_tree_add_6_33_groupi_g13567__7482(csa_tree_add_6_33_groupi_n_4727 ,csa_tree_add_6_33_groupi_n_4062 ,csa_tree_add_6_33_groupi_n_4725);
  xnor csa_tree_add_6_33_groupi_g13568__4733(csa_tree_add_6_33_groupi_n_4726 ,csa_tree_add_6_33_groupi_n_4646 ,csa_tree_add_6_33_groupi_n_4671);
  xnor csa_tree_add_6_33_groupi_g13569__6161(csa_tree_add_6_33_groupi_n_4743 ,csa_tree_add_6_33_groupi_n_4513 ,csa_tree_add_6_33_groupi_n_4627);
  xnor csa_tree_add_6_33_groupi_g13570__9315(csa_tree_add_6_33_groupi_n_4741 ,csa_tree_add_6_33_groupi_n_4538 ,csa_tree_add_6_33_groupi_n_4619);
  or csa_tree_add_6_33_groupi_g13571__9945(csa_tree_add_6_33_groupi_n_4739 ,csa_tree_add_6_33_groupi_n_4629 ,csa_tree_add_6_33_groupi_n_4701);
  xnor csa_tree_add_6_33_groupi_g13572__2883(csa_tree_add_6_33_groupi_n_4736 ,csa_tree_add_6_33_groupi_n_4572 ,csa_tree_add_6_33_groupi_n_4620);
  xnor csa_tree_add_6_33_groupi_g13574__2346(csa_tree_add_6_33_groupi_n_4734 ,csa_tree_add_6_33_groupi_n_4540 ,csa_tree_add_6_33_groupi_n_4623);
  xnor csa_tree_add_6_33_groupi_g13575__1666(csa_tree_add_6_33_groupi_n_4733 ,csa_tree_add_6_33_groupi_n_4536 ,csa_tree_add_6_33_groupi_n_4622);
  not csa_tree_add_6_33_groupi_g13576(csa_tree_add_6_33_groupi_n_4723 ,csa_tree_add_6_33_groupi_n_4724);
  not csa_tree_add_6_33_groupi_g13577(csa_tree_add_6_33_groupi_n_4721 ,csa_tree_add_6_33_groupi_n_4720);
  not csa_tree_add_6_33_groupi_g13578(csa_tree_add_6_33_groupi_n_4718 ,csa_tree_add_6_33_groupi_n_4719);
  not csa_tree_add_6_33_groupi_g13579(csa_tree_add_6_33_groupi_n_4715 ,csa_tree_add_6_33_groupi_n_4716);
  not csa_tree_add_6_33_groupi_g13580(csa_tree_add_6_33_groupi_n_4714 ,csa_tree_add_6_33_groupi_n_4713);
  not csa_tree_add_6_33_groupi_g13581(csa_tree_add_6_33_groupi_n_4711 ,csa_tree_add_6_33_groupi_n_4712);
  not csa_tree_add_6_33_groupi_g13582(csa_tree_add_6_33_groupi_n_4709 ,csa_tree_add_6_33_groupi_n_4710);
  or csa_tree_add_6_33_groupi_g13583__7410(csa_tree_add_6_33_groupi_n_4707 ,csa_tree_add_6_33_groupi_n_4616 ,csa_tree_add_6_33_groupi_n_4664);
  or csa_tree_add_6_33_groupi_g13584__6417(csa_tree_add_6_33_groupi_n_4706 ,csa_tree_add_6_33_groupi_n_4617 ,csa_tree_add_6_33_groupi_n_4661);
  and csa_tree_add_6_33_groupi_g13585__5477(csa_tree_add_6_33_groupi_n_4705 ,csa_tree_add_6_33_groupi_n_4671 ,csa_tree_add_6_33_groupi_n_4646);
  and csa_tree_add_6_33_groupi_g13586__2398(csa_tree_add_6_33_groupi_n_4704 ,csa_tree_add_6_33_groupi_n_4656 ,csa_tree_add_6_33_groupi_n_4579);
  or csa_tree_add_6_33_groupi_g13587__5107(csa_tree_add_6_33_groupi_n_4703 ,csa_tree_add_6_33_groupi_n_4671 ,csa_tree_add_6_33_groupi_n_4646);
  or csa_tree_add_6_33_groupi_g13588__6260(csa_tree_add_6_33_groupi_n_4702 ,csa_tree_add_6_33_groupi_n_4537 ,csa_tree_add_6_33_groupi_n_4649);
  nor csa_tree_add_6_33_groupi_g13589__4319(csa_tree_add_6_33_groupi_n_4701 ,csa_tree_add_6_33_groupi_n_4628 ,csa_tree_add_6_33_groupi_n_4582);
  xnor csa_tree_add_6_33_groupi_g13590__8428(csa_tree_add_6_33_groupi_n_4700 ,csa_tree_add_6_33_groupi_n_4430 ,csa_tree_add_6_33_groupi_n_4568);
  xnor csa_tree_add_6_33_groupi_g13591__5526(csa_tree_add_6_33_groupi_n_4699 ,csa_tree_add_6_33_groupi_n_4423 ,csa_tree_add_6_33_groupi_n_4579);
  or csa_tree_add_6_33_groupi_g13592__6783(csa_tree_add_6_33_groupi_n_4725 ,csa_tree_add_6_33_groupi_n_3946 ,csa_tree_add_6_33_groupi_n_4639);
  and csa_tree_add_6_33_groupi_g13593__3680(csa_tree_add_6_33_groupi_n_4724 ,csa_tree_add_6_33_groupi_n_4602 ,csa_tree_add_6_33_groupi_n_4658);
  and csa_tree_add_6_33_groupi_g13594__1617(csa_tree_add_6_33_groupi_n_4722 ,csa_tree_add_6_33_groupi_n_4554 ,csa_tree_add_6_33_groupi_n_4648);
  and csa_tree_add_6_33_groupi_g13595__2802(csa_tree_add_6_33_groupi_n_4720 ,csa_tree_add_6_33_groupi_n_4584 ,csa_tree_add_6_33_groupi_n_4654);
  and csa_tree_add_6_33_groupi_g13596__1705(csa_tree_add_6_33_groupi_n_4719 ,csa_tree_add_6_33_groupi_n_4556 ,csa_tree_add_6_33_groupi_n_4660);
  and csa_tree_add_6_33_groupi_g13597__5122(csa_tree_add_6_33_groupi_n_4717 ,csa_tree_add_6_33_groupi_n_4600 ,csa_tree_add_6_33_groupi_n_4641);
  and csa_tree_add_6_33_groupi_g13598__8246(csa_tree_add_6_33_groupi_n_4716 ,csa_tree_add_6_33_groupi_n_4605 ,csa_tree_add_6_33_groupi_n_4657);
  or csa_tree_add_6_33_groupi_g13599__7098(csa_tree_add_6_33_groupi_n_4713 ,csa_tree_add_6_33_groupi_n_4597 ,csa_tree_add_6_33_groupi_n_4630);
  and csa_tree_add_6_33_groupi_g13600__6131(csa_tree_add_6_33_groupi_n_4712 ,csa_tree_add_6_33_groupi_n_4607 ,csa_tree_add_6_33_groupi_n_4655);
  and csa_tree_add_6_33_groupi_g13601__1881(csa_tree_add_6_33_groupi_n_4710 ,csa_tree_add_6_33_groupi_n_4595 ,csa_tree_add_6_33_groupi_n_4659);
  and csa_tree_add_6_33_groupi_g13602__5115(csa_tree_add_6_33_groupi_n_4708 ,csa_tree_add_6_33_groupi_n_4587 ,csa_tree_add_6_33_groupi_n_4647);
  not csa_tree_add_6_33_groupi_g13603(csa_tree_add_6_33_groupi_n_4698 ,csa_tree_add_6_33_groupi_n_4697);
  not csa_tree_add_6_33_groupi_g13604(csa_tree_add_6_33_groupi_n_4696 ,csa_tree_add_6_33_groupi_n_4695);
  not csa_tree_add_6_33_groupi_g13605(csa_tree_add_6_33_groupi_n_4694 ,csa_tree_add_6_33_groupi_n_4693);
  not csa_tree_add_6_33_groupi_g13606(csa_tree_add_6_33_groupi_n_4691 ,csa_tree_add_6_33_groupi_n_4690);
  not csa_tree_add_6_33_groupi_g13607(csa_tree_add_6_33_groupi_n_4688 ,csa_tree_add_6_33_groupi_n_4687);
  xnor csa_tree_add_6_33_groupi_g13608__7482(out1[8] ,csa_tree_add_6_33_groupi_n_4618 ,csa_tree_add_6_33_groupi_n_4046);
  xnor csa_tree_add_6_33_groupi_g13609__4733(csa_tree_add_6_33_groupi_n_4685 ,csa_tree_add_6_33_groupi_n_4510 ,csa_tree_add_6_33_groupi_n_4569);
  xnor csa_tree_add_6_33_groupi_g13610__6161(csa_tree_add_6_33_groupi_n_4684 ,csa_tree_add_6_33_groupi_n_4566 ,csa_tree_add_6_33_groupi_n_4382);
  xnor csa_tree_add_6_33_groupi_g13611__9315(csa_tree_add_6_33_groupi_n_4683 ,csa_tree_add_6_33_groupi_n_4329 ,csa_tree_add_6_33_groupi_n_4581);
  xnor csa_tree_add_6_33_groupi_g13612__9945(csa_tree_add_6_33_groupi_n_4682 ,csa_tree_add_6_33_groupi_n_4558 ,csa_tree_add_6_33_groupi_n_4509);
  xnor csa_tree_add_6_33_groupi_g13613__2883(csa_tree_add_6_33_groupi_n_4681 ,csa_tree_add_6_33_groupi_n_4426 ,csa_tree_add_6_33_groupi_n_4580);
  xnor csa_tree_add_6_33_groupi_g13614__2346(csa_tree_add_6_33_groupi_n_4680 ,csa_tree_add_6_33_groupi_n_4565 ,csa_tree_add_6_33_groupi_n_4535);
  xnor csa_tree_add_6_33_groupi_g13615__1666(csa_tree_add_6_33_groupi_n_4679 ,csa_tree_add_6_33_groupi_n_4615 ,csa_tree_add_6_33_groupi_n_4563);
  xnor csa_tree_add_6_33_groupi_g13616__7410(csa_tree_add_6_33_groupi_n_4678 ,csa_tree_add_6_33_groupi_n_4431 ,csa_tree_add_6_33_groupi_n_4582);
  xnor csa_tree_add_6_33_groupi_g13617__6417(csa_tree_add_6_33_groupi_n_4677 ,csa_tree_add_6_33_groupi_n_4614 ,csa_tree_add_6_33_groupi_n_4562);
  xnor csa_tree_add_6_33_groupi_g13618__5477(csa_tree_add_6_33_groupi_n_4676 ,csa_tree_add_6_33_groupi_n_4534 ,csa_tree_add_6_33_groupi_n_4560);
  xnor csa_tree_add_6_33_groupi_g13619__2398(csa_tree_add_6_33_groupi_n_4675 ,csa_tree_add_6_33_groupi_n_4512 ,csa_tree_add_6_33_groupi_n_4578);
  xnor csa_tree_add_6_33_groupi_g13620__5107(csa_tree_add_6_33_groupi_n_4674 ,csa_tree_add_6_33_groupi_n_4531 ,csa_tree_add_6_33_groupi_n_4575);
  xnor csa_tree_add_6_33_groupi_g13621__6260(csa_tree_add_6_33_groupi_n_4673 ,csa_tree_add_6_33_groupi_n_4463 ,csa_tree_add_6_33_groupi_n_4574);
  xnor csa_tree_add_6_33_groupi_g13622__4319(csa_tree_add_6_33_groupi_n_4697 ,csa_tree_add_6_33_groupi_n_4323 ,csa_tree_add_6_33_groupi_n_4550);
  xnor csa_tree_add_6_33_groupi_g13623__8428(csa_tree_add_6_33_groupi_n_4695 ,csa_tree_add_6_33_groupi_n_4473 ,csa_tree_add_6_33_groupi_n_4541);
  xnor csa_tree_add_6_33_groupi_g13624__5526(csa_tree_add_6_33_groupi_n_4693 ,csa_tree_add_6_33_groupi_n_4497 ,csa_tree_add_6_33_groupi_n_4549);
  xnor csa_tree_add_6_33_groupi_g13625__6783(csa_tree_add_6_33_groupi_n_4692 ,csa_tree_add_6_33_groupi_n_4504 ,csa_tree_add_6_33_groupi_n_4546);
  xnor csa_tree_add_6_33_groupi_g13626__3680(csa_tree_add_6_33_groupi_n_4690 ,csa_tree_add_6_33_groupi_n_4433 ,csa_tree_add_6_33_groupi_n_4548);
  xnor csa_tree_add_6_33_groupi_g13627__1617(csa_tree_add_6_33_groupi_n_4689 ,csa_tree_add_6_33_groupi_n_4479 ,csa_tree_add_6_33_groupi_n_4542);
  xnor csa_tree_add_6_33_groupi_g13628__2802(csa_tree_add_6_33_groupi_n_4687 ,csa_tree_add_6_33_groupi_n_4498 ,csa_tree_add_6_33_groupi_n_4547);
  nor csa_tree_add_6_33_groupi_g13629__1705(csa_tree_add_6_33_groupi_n_4670 ,csa_tree_add_6_33_groupi_n_4423 ,csa_tree_add_6_33_groupi_n_4610);
  nor csa_tree_add_6_33_groupi_g13630__5122(csa_tree_add_6_33_groupi_n_4669 ,csa_tree_add_6_33_groupi_n_4531 ,csa_tree_add_6_33_groupi_n_4576);
  and csa_tree_add_6_33_groupi_g13631__8246(csa_tree_add_6_33_groupi_n_4668 ,csa_tree_add_6_33_groupi_n_4510 ,csa_tree_add_6_33_groupi_n_4570);
  and csa_tree_add_6_33_groupi_g13632__7098(csa_tree_add_6_33_groupi_n_4667 ,csa_tree_add_6_33_groupi_n_4535 ,csa_tree_add_6_33_groupi_n_4565);
  or csa_tree_add_6_33_groupi_g13633__6131(csa_tree_add_6_33_groupi_n_4666 ,csa_tree_add_6_33_groupi_n_4430 ,csa_tree_add_6_33_groupi_n_4567);
  and csa_tree_add_6_33_groupi_g13634__1881(csa_tree_add_6_33_groupi_n_4665 ,csa_tree_add_6_33_groupi_n_4531 ,csa_tree_add_6_33_groupi_n_4576);
  nor csa_tree_add_6_33_groupi_g13635__5115(csa_tree_add_6_33_groupi_n_4664 ,csa_tree_add_6_33_groupi_n_4429 ,csa_tree_add_6_33_groupi_n_4568);
  or csa_tree_add_6_33_groupi_g13636__7482(csa_tree_add_6_33_groupi_n_4663 ,csa_tree_add_6_33_groupi_n_4382 ,csa_tree_add_6_33_groupi_n_4566);
  nor csa_tree_add_6_33_groupi_g13637__4733(csa_tree_add_6_33_groupi_n_4662 ,csa_tree_add_6_33_groupi_n_4615 ,csa_tree_add_6_33_groupi_n_4564);
  and csa_tree_add_6_33_groupi_g13638__6161(csa_tree_add_6_33_groupi_n_4661 ,csa_tree_add_6_33_groupi_n_4382 ,csa_tree_add_6_33_groupi_n_4566);
  or csa_tree_add_6_33_groupi_g13639__9315(csa_tree_add_6_33_groupi_n_4660 ,csa_tree_add_6_33_groupi_n_4340 ,csa_tree_add_6_33_groupi_n_4555);
  or csa_tree_add_6_33_groupi_g13640__9945(csa_tree_add_6_33_groupi_n_4659 ,csa_tree_add_6_33_groupi_n_4471 ,csa_tree_add_6_33_groupi_n_4594);
  or csa_tree_add_6_33_groupi_g13641__2883(csa_tree_add_6_33_groupi_n_4658 ,csa_tree_add_6_33_groupi_n_4553 ,csa_tree_add_6_33_groupi_n_4580);
  or csa_tree_add_6_33_groupi_g13642__2346(csa_tree_add_6_33_groupi_n_4657 ,csa_tree_add_6_33_groupi_n_4536 ,csa_tree_add_6_33_groupi_n_4604);
  or csa_tree_add_6_33_groupi_g13643__1666(csa_tree_add_6_33_groupi_n_4656 ,csa_tree_add_6_33_groupi_n_4422 ,csa_tree_add_6_33_groupi_n_4609);
  or csa_tree_add_6_33_groupi_g13644__7410(csa_tree_add_6_33_groupi_n_4655 ,csa_tree_add_6_33_groupi_n_4540 ,csa_tree_add_6_33_groupi_n_4590);
  or csa_tree_add_6_33_groupi_g13645__6417(csa_tree_add_6_33_groupi_n_4654 ,csa_tree_add_6_33_groupi_n_4539 ,csa_tree_add_6_33_groupi_n_4583);
  and csa_tree_add_6_33_groupi_g13646__5477(csa_tree_add_6_33_groupi_n_4653 ,csa_tree_add_6_33_groupi_n_4615 ,csa_tree_add_6_33_groupi_n_4564);
  or csa_tree_add_6_33_groupi_g13647__2398(csa_tree_add_6_33_groupi_n_4652 ,csa_tree_add_6_33_groupi_n_4535 ,csa_tree_add_6_33_groupi_n_4565);
  and csa_tree_add_6_33_groupi_g13648__5107(csa_tree_add_6_33_groupi_n_4651 ,csa_tree_add_6_33_groupi_n_4509 ,csa_tree_add_6_33_groupi_n_4558);
  or csa_tree_add_6_33_groupi_g13649__6260(csa_tree_add_6_33_groupi_n_4650 ,csa_tree_add_6_33_groupi_n_4468 ,csa_tree_add_6_33_groupi_n_4571);
  nor csa_tree_add_6_33_groupi_g13650__4319(csa_tree_add_6_33_groupi_n_4649 ,csa_tree_add_6_33_groupi_n_4467 ,csa_tree_add_6_33_groupi_n_4572);
  or csa_tree_add_6_33_groupi_g13651__8428(csa_tree_add_6_33_groupi_n_4648 ,csa_tree_add_6_33_groupi_n_4557 ,csa_tree_add_6_33_groupi_n_4581);
  or csa_tree_add_6_33_groupi_g13652__5526(csa_tree_add_6_33_groupi_n_4647 ,csa_tree_add_6_33_groupi_n_4538 ,csa_tree_add_6_33_groupi_n_4592);
  or csa_tree_add_6_33_groupi_g13653__6783(csa_tree_add_6_33_groupi_n_4672 ,csa_tree_add_6_33_groupi_n_4525 ,csa_tree_add_6_33_groupi_n_4589);
  and csa_tree_add_6_33_groupi_g13654__3680(csa_tree_add_6_33_groupi_n_4671 ,csa_tree_add_6_33_groupi_n_4515 ,csa_tree_add_6_33_groupi_n_4588);
  not csa_tree_add_6_33_groupi_g13655(csa_tree_add_6_33_groupi_n_4644 ,csa_tree_add_6_33_groupi_n_4645);
  or csa_tree_add_6_33_groupi_g13656__1617(csa_tree_add_6_33_groupi_n_4642 ,csa_tree_add_6_33_groupi_n_4509 ,csa_tree_add_6_33_groupi_n_4558);
  or csa_tree_add_6_33_groupi_g13657__2802(csa_tree_add_6_33_groupi_n_4641 ,csa_tree_add_6_33_groupi_n_4513 ,csa_tree_add_6_33_groupi_n_4606);
  nor csa_tree_add_6_33_groupi_g13658__1705(csa_tree_add_6_33_groupi_n_4640 ,csa_tree_add_6_33_groupi_n_4510 ,csa_tree_add_6_33_groupi_n_4570);
  and csa_tree_add_6_33_groupi_g13659__5122(csa_tree_add_6_33_groupi_n_4639 ,csa_tree_add_6_33_groupi_n_3947 ,csa_tree_add_6_33_groupi_n_4618);
  or csa_tree_add_6_33_groupi_g13660__8246(csa_tree_add_6_33_groupi_n_4638 ,csa_tree_add_6_33_groupi_n_4614 ,csa_tree_add_6_33_groupi_n_4561);
  or csa_tree_add_6_33_groupi_g13661__7098(csa_tree_add_6_33_groupi_n_4637 ,csa_tree_add_6_33_groupi_n_4534 ,csa_tree_add_6_33_groupi_n_4559);
  nor csa_tree_add_6_33_groupi_g13662__6131(csa_tree_add_6_33_groupi_n_4636 ,csa_tree_add_6_33_groupi_n_4533 ,csa_tree_add_6_33_groupi_n_4560);
  nor csa_tree_add_6_33_groupi_g13663__1881(csa_tree_add_6_33_groupi_n_4635 ,csa_tree_add_6_33_groupi_n_4512 ,csa_tree_add_6_33_groupi_n_4578);
  or csa_tree_add_6_33_groupi_g13664__5115(csa_tree_add_6_33_groupi_n_4634 ,csa_tree_add_6_33_groupi_n_4462 ,csa_tree_add_6_33_groupi_n_4573);
  nor csa_tree_add_6_33_groupi_g13665__7482(csa_tree_add_6_33_groupi_n_4633 ,csa_tree_add_6_33_groupi_n_4463 ,csa_tree_add_6_33_groupi_n_4574);
  or csa_tree_add_6_33_groupi_g13666__4733(csa_tree_add_6_33_groupi_n_4632 ,csa_tree_add_6_33_groupi_n_4511 ,csa_tree_add_6_33_groupi_n_4577);
  nor csa_tree_add_6_33_groupi_g13667__6161(csa_tree_add_6_33_groupi_n_4631 ,csa_tree_add_6_33_groupi_n_4613 ,csa_tree_add_6_33_groupi_n_4562);
  nor csa_tree_add_6_33_groupi_g13668__9315(csa_tree_add_6_33_groupi_n_4630 ,csa_tree_add_6_33_groupi_n_4477 ,csa_tree_add_6_33_groupi_n_4596);
  and csa_tree_add_6_33_groupi_g13669__9945(csa_tree_add_6_33_groupi_n_4629 ,csa_tree_add_6_33_groupi_n_4431 ,csa_tree_add_6_33_groupi_n_4608);
  nor csa_tree_add_6_33_groupi_g13670__2883(csa_tree_add_6_33_groupi_n_4628 ,csa_tree_add_6_33_groupi_n_4431 ,csa_tree_add_6_33_groupi_n_4608);
  xnor csa_tree_add_6_33_groupi_g13671__2346(csa_tree_add_6_33_groupi_n_4627 ,csa_tree_add_6_33_groupi_n_4417 ,csa_tree_add_6_33_groupi_n_4491);
  xnor csa_tree_add_6_33_groupi_g13672__1666(csa_tree_add_6_33_groupi_n_4626 ,csa_tree_add_6_33_groupi_n_4532 ,csa_tree_add_6_33_groupi_n_4505);
  xnor csa_tree_add_6_33_groupi_g13673__7410(csa_tree_add_6_33_groupi_n_4625 ,csa_tree_add_6_33_groupi_n_4460 ,csa_tree_add_6_33_groupi_n_4503);
  xnor csa_tree_add_6_33_groupi_g13674__6417(csa_tree_add_6_33_groupi_n_4624 ,csa_tree_add_6_33_groupi_n_4384 ,csa_tree_add_6_33_groupi_n_4500);
  xnor csa_tree_add_6_33_groupi_g13675__5477(csa_tree_add_6_33_groupi_n_4623 ,csa_tree_add_6_33_groupi_n_4496 ,csa_tree_add_6_33_groupi_n_4219);
  xnor csa_tree_add_6_33_groupi_g13676__2398(csa_tree_add_6_33_groupi_n_4622 ,csa_tree_add_6_33_groupi_n_4495 ,csa_tree_add_6_33_groupi_n_4411);
  xnor csa_tree_add_6_33_groupi_g13677__5107(csa_tree_add_6_33_groupi_n_4621 ,csa_tree_add_6_33_groupi_n_4492 ,csa_tree_add_6_33_groupi_n_4466);
  xnor csa_tree_add_6_33_groupi_g13678__6260(csa_tree_add_6_33_groupi_n_4620 ,csa_tree_add_6_33_groupi_n_4537 ,csa_tree_add_6_33_groupi_n_4468);
  xnor csa_tree_add_6_33_groupi_g13679__4319(csa_tree_add_6_33_groupi_n_4619 ,csa_tree_add_6_33_groupi_n_4163 ,csa_tree_add_6_33_groupi_n_4508);
  xnor csa_tree_add_6_33_groupi_g13680__8428(csa_tree_add_6_33_groupi_n_4646 ,csa_tree_add_6_33_groupi_n_4475 ,csa_tree_add_6_33_groupi_n_4481);
  and csa_tree_add_6_33_groupi_g13681__5526(csa_tree_add_6_33_groupi_n_4645 ,csa_tree_add_6_33_groupi_n_4483 ,csa_tree_add_6_33_groupi_n_4599);
  and csa_tree_add_6_33_groupi_g13682__6783(csa_tree_add_6_33_groupi_n_4643 ,csa_tree_add_6_33_groupi_n_4484 ,csa_tree_add_6_33_groupi_n_4601);
  not csa_tree_add_6_33_groupi_g13683(csa_tree_add_6_33_groupi_n_4613 ,csa_tree_add_6_33_groupi_n_4614);
  not csa_tree_add_6_33_groupi_g13684(csa_tree_add_6_33_groupi_n_4611 ,csa_tree_add_6_33_groupi_n_4612);
  not csa_tree_add_6_33_groupi_g13685(csa_tree_add_6_33_groupi_n_4609 ,csa_tree_add_6_33_groupi_n_4610);
  or csa_tree_add_6_33_groupi_g13686__3680(csa_tree_add_6_33_groupi_n_4607 ,csa_tree_add_6_33_groupi_n_4219 ,csa_tree_add_6_33_groupi_n_4496);
  nor csa_tree_add_6_33_groupi_g13687__1617(csa_tree_add_6_33_groupi_n_4606 ,csa_tree_add_6_33_groupi_n_4417 ,csa_tree_add_6_33_groupi_n_4490);
  or csa_tree_add_6_33_groupi_g13688__2802(csa_tree_add_6_33_groupi_n_4605 ,csa_tree_add_6_33_groupi_n_4411 ,csa_tree_add_6_33_groupi_n_4495);
  and csa_tree_add_6_33_groupi_g13689__1705(csa_tree_add_6_33_groupi_n_4604 ,csa_tree_add_6_33_groupi_n_4411 ,csa_tree_add_6_33_groupi_n_4495);
  or csa_tree_add_6_33_groupi_g13690__5122(csa_tree_add_6_33_groupi_n_4603 ,csa_tree_add_6_33_groupi_n_4460 ,csa_tree_add_6_33_groupi_n_4502);
  or csa_tree_add_6_33_groupi_g13691__8246(csa_tree_add_6_33_groupi_n_4602 ,csa_tree_add_6_33_groupi_n_4427 ,csa_tree_add_6_33_groupi_n_4501);
  or csa_tree_add_6_33_groupi_g13692__7098(csa_tree_add_6_33_groupi_n_4601 ,csa_tree_add_6_33_groupi_n_4108 ,csa_tree_add_6_33_groupi_n_4487);
  or csa_tree_add_6_33_groupi_g13693__6131(csa_tree_add_6_33_groupi_n_4600 ,csa_tree_add_6_33_groupi_n_4416 ,csa_tree_add_6_33_groupi_n_4491);
  or csa_tree_add_6_33_groupi_g13694__1881(csa_tree_add_6_33_groupi_n_4599 ,csa_tree_add_6_33_groupi_n_4472 ,csa_tree_add_6_33_groupi_n_4488);
  nor csa_tree_add_6_33_groupi_g13695__5115(csa_tree_add_6_33_groupi_n_4598 ,csa_tree_add_6_33_groupi_n_4459 ,csa_tree_add_6_33_groupi_n_4503);
  and csa_tree_add_6_33_groupi_g13696__7482(csa_tree_add_6_33_groupi_n_4597 ,csa_tree_add_6_33_groupi_n_3960 ,csa_tree_add_6_33_groupi_n_4504);
  nor csa_tree_add_6_33_groupi_g13697__4733(csa_tree_add_6_33_groupi_n_4596 ,csa_tree_add_6_33_groupi_n_3960 ,csa_tree_add_6_33_groupi_n_4504);
  or csa_tree_add_6_33_groupi_g13698__6161(csa_tree_add_6_33_groupi_n_4595 ,csa_tree_add_6_33_groupi_n_4202 ,csa_tree_add_6_33_groupi_n_4497);
  and csa_tree_add_6_33_groupi_g13699__9315(csa_tree_add_6_33_groupi_n_4594 ,csa_tree_add_6_33_groupi_n_4202 ,csa_tree_add_6_33_groupi_n_4497);
  or csa_tree_add_6_33_groupi_g13700__9945(csa_tree_add_6_33_groupi_n_4593 ,csa_tree_add_6_33_groupi_n_4466 ,csa_tree_add_6_33_groupi_n_4492);
  nor csa_tree_add_6_33_groupi_g13701__2883(csa_tree_add_6_33_groupi_n_4592 ,csa_tree_add_6_33_groupi_n_4162 ,csa_tree_add_6_33_groupi_n_4508);
  and csa_tree_add_6_33_groupi_g13702__2346(csa_tree_add_6_33_groupi_n_4591 ,csa_tree_add_6_33_groupi_n_4532 ,csa_tree_add_6_33_groupi_n_4506);
  and csa_tree_add_6_33_groupi_g13703__1666(csa_tree_add_6_33_groupi_n_4590 ,csa_tree_add_6_33_groupi_n_4219 ,csa_tree_add_6_33_groupi_n_4496);
  nor csa_tree_add_6_33_groupi_g13704__7410(csa_tree_add_6_33_groupi_n_4589 ,csa_tree_add_6_33_groupi_n_4473 ,csa_tree_add_6_33_groupi_n_4529);
  or csa_tree_add_6_33_groupi_g13705__6417(csa_tree_add_6_33_groupi_n_4588 ,csa_tree_add_6_33_groupi_n_4479 ,csa_tree_add_6_33_groupi_n_4527);
  or csa_tree_add_6_33_groupi_g13706__5477(csa_tree_add_6_33_groupi_n_4587 ,csa_tree_add_6_33_groupi_n_4163 ,csa_tree_add_6_33_groupi_n_4507);
  and csa_tree_add_6_33_groupi_g13707__2398(csa_tree_add_6_33_groupi_n_4586 ,csa_tree_add_6_33_groupi_n_4466 ,csa_tree_add_6_33_groupi_n_4492);
  nor csa_tree_add_6_33_groupi_g13708__5107(csa_tree_add_6_33_groupi_n_4585 ,csa_tree_add_6_33_groupi_n_4532 ,csa_tree_add_6_33_groupi_n_4506);
  or csa_tree_add_6_33_groupi_g13709__6260(csa_tree_add_6_33_groupi_n_4584 ,csa_tree_add_6_33_groupi_n_4384 ,csa_tree_add_6_33_groupi_n_4499);
  nor csa_tree_add_6_33_groupi_g13710__4319(csa_tree_add_6_33_groupi_n_4583 ,csa_tree_add_6_33_groupi_n_4383 ,csa_tree_add_6_33_groupi_n_4500);
  or csa_tree_add_6_33_groupi_g13711__8428(csa_tree_add_6_33_groupi_n_4618 ,csa_tree_add_6_33_groupi_n_3601 ,csa_tree_add_6_33_groupi_n_4486);
  and csa_tree_add_6_33_groupi_g13712__5526(csa_tree_add_6_33_groupi_n_4617 ,csa_tree_add_6_33_groupi_n_4359 ,csa_tree_add_6_33_groupi_n_4516);
  and csa_tree_add_6_33_groupi_g13713__6783(csa_tree_add_6_33_groupi_n_4616 ,csa_tree_add_6_33_groupi_n_4370 ,csa_tree_add_6_33_groupi_n_4522);
  and csa_tree_add_6_33_groupi_g13714__3680(csa_tree_add_6_33_groupi_n_4615 ,csa_tree_add_6_33_groupi_n_4448 ,csa_tree_add_6_33_groupi_n_4530);
  and csa_tree_add_6_33_groupi_g13715__1617(csa_tree_add_6_33_groupi_n_4614 ,csa_tree_add_6_33_groupi_n_4445 ,csa_tree_add_6_33_groupi_n_4528);
  or csa_tree_add_6_33_groupi_g13716__2802(csa_tree_add_6_33_groupi_n_4612 ,csa_tree_add_6_33_groupi_n_4307 ,csa_tree_add_6_33_groupi_n_4517);
  and csa_tree_add_6_33_groupi_g13717__1705(csa_tree_add_6_33_groupi_n_4610 ,csa_tree_add_6_33_groupi_n_4346 ,csa_tree_add_6_33_groupi_n_4514);
  or csa_tree_add_6_33_groupi_g13718__5122(csa_tree_add_6_33_groupi_n_4608 ,csa_tree_add_6_33_groupi_n_4352 ,csa_tree_add_6_33_groupi_n_4524);
  not csa_tree_add_6_33_groupi_g13719(csa_tree_add_6_33_groupi_n_4578 ,csa_tree_add_6_33_groupi_n_4577);
  not csa_tree_add_6_33_groupi_g13720(csa_tree_add_6_33_groupi_n_4576 ,csa_tree_add_6_33_groupi_n_4575);
  not csa_tree_add_6_33_groupi_g13721(csa_tree_add_6_33_groupi_n_4574 ,csa_tree_add_6_33_groupi_n_4573);
  not csa_tree_add_6_33_groupi_g13722(csa_tree_add_6_33_groupi_n_4572 ,csa_tree_add_6_33_groupi_n_4571);
  not csa_tree_add_6_33_groupi_g13723(csa_tree_add_6_33_groupi_n_4570 ,csa_tree_add_6_33_groupi_n_4569);
  not csa_tree_add_6_33_groupi_g13724(csa_tree_add_6_33_groupi_n_4567 ,csa_tree_add_6_33_groupi_n_4568);
  not csa_tree_add_6_33_groupi_g13725(csa_tree_add_6_33_groupi_n_4564 ,csa_tree_add_6_33_groupi_n_4563);
  not csa_tree_add_6_33_groupi_g13726(csa_tree_add_6_33_groupi_n_4562 ,csa_tree_add_6_33_groupi_n_4561);
  not csa_tree_add_6_33_groupi_g13727(csa_tree_add_6_33_groupi_n_4560 ,csa_tree_add_6_33_groupi_n_4559);
  nor csa_tree_add_6_33_groupi_g13728__8246(csa_tree_add_6_33_groupi_n_4557 ,csa_tree_add_6_33_groupi_n_4329 ,csa_tree_add_6_33_groupi_n_4494);
  or csa_tree_add_6_33_groupi_g13729__7098(csa_tree_add_6_33_groupi_n_4556 ,csa_tree_add_6_33_groupi_n_4464 ,csa_tree_add_6_33_groupi_n_4498);
  and csa_tree_add_6_33_groupi_g13730__6131(csa_tree_add_6_33_groupi_n_4555 ,csa_tree_add_6_33_groupi_n_4464 ,csa_tree_add_6_33_groupi_n_4498);
  or csa_tree_add_6_33_groupi_g13731__1881(csa_tree_add_6_33_groupi_n_4554 ,csa_tree_add_6_33_groupi_n_4328 ,csa_tree_add_6_33_groupi_n_4493);
  and csa_tree_add_6_33_groupi_g13732__5115(csa_tree_add_6_33_groupi_n_4553 ,csa_tree_add_6_33_groupi_n_4427 ,csa_tree_add_6_33_groupi_n_4501);
  xnor csa_tree_add_6_33_groupi_g13733__7482(out1[7] ,csa_tree_add_6_33_groupi_n_4476 ,csa_tree_add_6_33_groupi_n_3798);
  xnor csa_tree_add_6_33_groupi_g13734__4733(csa_tree_add_6_33_groupi_n_4551 ,csa_tree_add_6_33_groupi_n_4461 ,csa_tree_add_6_33_groupi_n_4414);
  xnor csa_tree_add_6_33_groupi_g13735__6161(csa_tree_add_6_33_groupi_n_4550 ,csa_tree_add_6_33_groupi_n_4428 ,csa_tree_add_6_33_groupi_n_4108);
  xnor csa_tree_add_6_33_groupi_g13736__9315(csa_tree_add_6_33_groupi_n_4549 ,csa_tree_add_6_33_groupi_n_4471 ,csa_tree_add_6_33_groupi_n_4202);
  xnor csa_tree_add_6_33_groupi_g13737__9945(csa_tree_add_6_33_groupi_n_4548 ,csa_tree_add_6_33_groupi_n_4226 ,csa_tree_add_6_33_groupi_n_4472);
  xnor csa_tree_add_6_33_groupi_g13738__2883(csa_tree_add_6_33_groupi_n_4547 ,csa_tree_add_6_33_groupi_n_4464 ,csa_tree_add_6_33_groupi_n_4340);
  xnor csa_tree_add_6_33_groupi_g13739__2346(csa_tree_add_6_33_groupi_n_4546 ,csa_tree_add_6_33_groupi_n_3960 ,csa_tree_add_6_33_groupi_n_4477);
  xnor csa_tree_add_6_33_groupi_g13740__1666(csa_tree_add_6_33_groupi_n_4545 ,csa_tree_add_6_33_groupi_n_4470 ,csa_tree_add_6_33_groupi_n_4421);
  xnor csa_tree_add_6_33_groupi_g13741__7410(csa_tree_add_6_33_groupi_n_4544 ,csa_tree_add_6_33_groupi_n_4424 ,csa_tree_add_6_33_groupi_n_4465);
  xnor csa_tree_add_6_33_groupi_g13742__6417(csa_tree_add_6_33_groupi_n_4543 ,csa_tree_add_6_33_groupi_n_4425 ,csa_tree_add_6_33_groupi_n_4381);
  xnor csa_tree_add_6_33_groupi_g13743__5477(csa_tree_add_6_33_groupi_n_4542 ,csa_tree_add_6_33_groupi_n_4150 ,csa_tree_add_6_33_groupi_n_4413);
  xnor csa_tree_add_6_33_groupi_g13744__2398(csa_tree_add_6_33_groupi_n_4541 ,csa_tree_add_6_33_groupi_n_4154 ,csa_tree_add_6_33_groupi_n_4418);
  xnor csa_tree_add_6_33_groupi_g13745__5107(csa_tree_add_6_33_groupi_n_4582 ,csa_tree_add_6_33_groupi_n_4332 ,csa_tree_add_6_33_groupi_n_4403);
  xnor csa_tree_add_6_33_groupi_g13746__6260(csa_tree_add_6_33_groupi_n_4581 ,csa_tree_add_6_33_groupi_n_4387 ,csa_tree_add_6_33_groupi_n_4405);
  xnor csa_tree_add_6_33_groupi_g13747__4319(csa_tree_add_6_33_groupi_n_4580 ,csa_tree_add_6_33_groupi_n_4478 ,csa_tree_add_6_33_groupi_n_4396);
  xnor csa_tree_add_6_33_groupi_g13748__8428(csa_tree_add_6_33_groupi_n_4579 ,csa_tree_add_6_33_groupi_n_4474 ,csa_tree_add_6_33_groupi_n_4407);
  xnor csa_tree_add_6_33_groupi_g13749__5526(csa_tree_add_6_33_groupi_n_4577 ,csa_tree_add_6_33_groupi_n_4165 ,csa_tree_add_6_33_groupi_n_4399);
  xnor csa_tree_add_6_33_groupi_g13750__6783(csa_tree_add_6_33_groupi_n_4575 ,csa_tree_add_6_33_groupi_n_4287 ,csa_tree_add_6_33_groupi_n_4398);
  xnor csa_tree_add_6_33_groupi_g13751__3680(csa_tree_add_6_33_groupi_n_4573 ,csa_tree_add_6_33_groupi_n_4020 ,csa_tree_add_6_33_groupi_n_4397);
  xnor csa_tree_add_6_33_groupi_g13752__1617(csa_tree_add_6_33_groupi_n_4571 ,csa_tree_add_6_33_groupi_n_4436 ,csa_tree_add_6_33_groupi_n_4402);
  xnor csa_tree_add_6_33_groupi_g13753__2802(csa_tree_add_6_33_groupi_n_4569 ,csa_tree_add_6_33_groupi_n_4289 ,csa_tree_add_6_33_groupi_n_4390);
  xnor csa_tree_add_6_33_groupi_g13754__1705(csa_tree_add_6_33_groupi_n_4568 ,csa_tree_add_6_33_groupi_n_4386 ,csa_tree_add_6_33_groupi_n_4408);
  xnor csa_tree_add_6_33_groupi_g13755__5122(csa_tree_add_6_33_groupi_n_4566 ,csa_tree_add_6_33_groupi_n_4434 ,csa_tree_add_6_33_groupi_n_4394);
  xnor csa_tree_add_6_33_groupi_g13756__8246(csa_tree_add_6_33_groupi_n_4565 ,csa_tree_add_6_33_groupi_n_4336 ,csa_tree_add_6_33_groupi_n_4395);
  xnor csa_tree_add_6_33_groupi_g13757__7098(csa_tree_add_6_33_groupi_n_4563 ,csa_tree_add_6_33_groupi_n_4385 ,csa_tree_add_6_33_groupi_n_4393);
  xnor csa_tree_add_6_33_groupi_g13758__6131(csa_tree_add_6_33_groupi_n_4561 ,csa_tree_add_6_33_groupi_n_4435 ,csa_tree_add_6_33_groupi_n_4392);
  xnor csa_tree_add_6_33_groupi_g13759__1881(csa_tree_add_6_33_groupi_n_4559 ,csa_tree_add_6_33_groupi_n_4325 ,csa_tree_add_6_33_groupi_n_4400);
  xnor csa_tree_add_6_33_groupi_g13760__5115(csa_tree_add_6_33_groupi_n_4558 ,csa_tree_add_6_33_groupi_n_4291 ,csa_tree_add_6_33_groupi_n_4406);
  not csa_tree_add_6_33_groupi_g13762(csa_tree_add_6_33_groupi_n_4534 ,csa_tree_add_6_33_groupi_n_4533);
  or csa_tree_add_6_33_groupi_g13763__7482(csa_tree_add_6_33_groupi_n_4530 ,csa_tree_add_6_33_groupi_n_4475 ,csa_tree_add_6_33_groupi_n_4458);
  and csa_tree_add_6_33_groupi_g13764__4733(csa_tree_add_6_33_groupi_n_4529 ,csa_tree_add_6_33_groupi_n_4154 ,csa_tree_add_6_33_groupi_n_4419);
  or csa_tree_add_6_33_groupi_g13765__6161(csa_tree_add_6_33_groupi_n_4528 ,csa_tree_add_6_33_groupi_n_4286 ,csa_tree_add_6_33_groupi_n_4457);
  nor csa_tree_add_6_33_groupi_g13766__9315(csa_tree_add_6_33_groupi_n_4527 ,csa_tree_add_6_33_groupi_n_4149 ,csa_tree_add_6_33_groupi_n_4413);
  nor csa_tree_add_6_33_groupi_g13767__9945(csa_tree_add_6_33_groupi_n_4526 ,csa_tree_add_6_33_groupi_n_4461 ,csa_tree_add_6_33_groupi_n_4415);
  nor csa_tree_add_6_33_groupi_g13768__2883(csa_tree_add_6_33_groupi_n_4525 ,csa_tree_add_6_33_groupi_n_4154 ,csa_tree_add_6_33_groupi_n_4419);
  nor csa_tree_add_6_33_groupi_g13769__2346(csa_tree_add_6_33_groupi_n_4524 ,csa_tree_add_6_33_groupi_n_4376 ,csa_tree_add_6_33_groupi_n_4436);
  and csa_tree_add_6_33_groupi_g13770__1666(csa_tree_add_6_33_groupi_n_4523 ,csa_tree_add_6_33_groupi_n_4461 ,csa_tree_add_6_33_groupi_n_4415);
  or csa_tree_add_6_33_groupi_g13771__7410(csa_tree_add_6_33_groupi_n_4522 ,csa_tree_add_6_33_groupi_n_4366 ,csa_tree_add_6_33_groupi_n_4434);
  or csa_tree_add_6_33_groupi_g13772__6417(csa_tree_add_6_33_groupi_n_4521 ,csa_tree_add_6_33_groupi_n_4465 ,csa_tree_add_6_33_groupi_n_4424);
  and csa_tree_add_6_33_groupi_g13773__5477(csa_tree_add_6_33_groupi_n_4520 ,csa_tree_add_6_33_groupi_n_4465 ,csa_tree_add_6_33_groupi_n_4424);
  or csa_tree_add_6_33_groupi_g13774__2398(csa_tree_add_6_33_groupi_n_4519 ,csa_tree_add_6_33_groupi_n_4381 ,csa_tree_add_6_33_groupi_n_4425);
  and csa_tree_add_6_33_groupi_g13775__5107(csa_tree_add_6_33_groupi_n_4518 ,csa_tree_add_6_33_groupi_n_4381 ,csa_tree_add_6_33_groupi_n_4425);
  nor csa_tree_add_6_33_groupi_g13776__6260(csa_tree_add_6_33_groupi_n_4517 ,csa_tree_add_6_33_groupi_n_4380 ,csa_tree_add_6_33_groupi_n_4435);
  or csa_tree_add_6_33_groupi_g13777__4319(csa_tree_add_6_33_groupi_n_4516 ,csa_tree_add_6_33_groupi_n_4355 ,csa_tree_add_6_33_groupi_n_4474);
  or csa_tree_add_6_33_groupi_g13778__8428(csa_tree_add_6_33_groupi_n_4515 ,csa_tree_add_6_33_groupi_n_4150 ,csa_tree_add_6_33_groupi_n_4412);
  or csa_tree_add_6_33_groupi_g13779__5526(csa_tree_add_6_33_groupi_n_4514 ,csa_tree_add_6_33_groupi_n_4345 ,csa_tree_add_6_33_groupi_n_4478);
  and csa_tree_add_6_33_groupi_g13780__6783(csa_tree_add_6_33_groupi_n_4540 ,csa_tree_add_6_33_groupi_n_4281 ,csa_tree_add_6_33_groupi_n_4447);
  and csa_tree_add_6_33_groupi_g13781__3680(csa_tree_add_6_33_groupi_n_4539 ,csa_tree_add_6_33_groupi_n_4242 ,csa_tree_add_6_33_groupi_n_4440);
  and csa_tree_add_6_33_groupi_g13782__1617(csa_tree_add_6_33_groupi_n_4538 ,csa_tree_add_6_33_groupi_n_4245 ,csa_tree_add_6_33_groupi_n_4438);
  and csa_tree_add_6_33_groupi_g13783__2802(csa_tree_add_6_33_groupi_n_4537 ,csa_tree_add_6_33_groupi_n_4362 ,csa_tree_add_6_33_groupi_n_4443);
  and csa_tree_add_6_33_groupi_g13784__1705(csa_tree_add_6_33_groupi_n_4536 ,csa_tree_add_6_33_groupi_n_4379 ,csa_tree_add_6_33_groupi_n_4456);
  and csa_tree_add_6_33_groupi_g13785__5122(csa_tree_add_6_33_groupi_n_4535 ,csa_tree_add_6_33_groupi_n_4374 ,csa_tree_add_6_33_groupi_n_4452);
  or csa_tree_add_6_33_groupi_g13786__8246(csa_tree_add_6_33_groupi_n_4533 ,csa_tree_add_6_33_groupi_n_4378 ,csa_tree_add_6_33_groupi_n_4455);
  and csa_tree_add_6_33_groupi_g13787__7098(csa_tree_add_6_33_groupi_n_4532 ,csa_tree_add_6_33_groupi_n_4364 ,csa_tree_add_6_33_groupi_n_4442);
  and csa_tree_add_6_33_groupi_g13788__6131(csa_tree_add_6_33_groupi_n_4531 ,csa_tree_add_6_33_groupi_n_4311 ,csa_tree_add_6_33_groupi_n_4454);
  not csa_tree_add_6_33_groupi_g13789(csa_tree_add_6_33_groupi_n_4512 ,csa_tree_add_6_33_groupi_n_4511);
  not csa_tree_add_6_33_groupi_g13790(csa_tree_add_6_33_groupi_n_4507 ,csa_tree_add_6_33_groupi_n_4508);
  not csa_tree_add_6_33_groupi_g13791(csa_tree_add_6_33_groupi_n_4506 ,csa_tree_add_6_33_groupi_n_4505);
  not csa_tree_add_6_33_groupi_g13792(csa_tree_add_6_33_groupi_n_4503 ,csa_tree_add_6_33_groupi_n_4502);
  not csa_tree_add_6_33_groupi_g13793(csa_tree_add_6_33_groupi_n_4500 ,csa_tree_add_6_33_groupi_n_4499);
  not csa_tree_add_6_33_groupi_g13794(csa_tree_add_6_33_groupi_n_4494 ,csa_tree_add_6_33_groupi_n_4493);
  not csa_tree_add_6_33_groupi_g13795(csa_tree_add_6_33_groupi_n_4490 ,csa_tree_add_6_33_groupi_n_4491);
  nor csa_tree_add_6_33_groupi_g13796__1881(csa_tree_add_6_33_groupi_n_4489 ,csa_tree_add_6_33_groupi_n_4470 ,csa_tree_add_6_33_groupi_n_4421);
  nor csa_tree_add_6_33_groupi_g13797__5115(csa_tree_add_6_33_groupi_n_4488 ,csa_tree_add_6_33_groupi_n_4226 ,csa_tree_add_6_33_groupi_n_4433);
  and csa_tree_add_6_33_groupi_g13798__7482(csa_tree_add_6_33_groupi_n_4487 ,csa_tree_add_6_33_groupi_n_4323 ,csa_tree_add_6_33_groupi_n_4428);
  and csa_tree_add_6_33_groupi_g13799__4733(csa_tree_add_6_33_groupi_n_4486 ,csa_tree_add_6_33_groupi_n_3600 ,csa_tree_add_6_33_groupi_n_4476);
  or csa_tree_add_6_33_groupi_g13800__6161(csa_tree_add_6_33_groupi_n_4485 ,csa_tree_add_6_33_groupi_n_4469 ,csa_tree_add_6_33_groupi_n_4420);
  or csa_tree_add_6_33_groupi_g13801__9315(csa_tree_add_6_33_groupi_n_4484 ,csa_tree_add_6_33_groupi_n_4323 ,csa_tree_add_6_33_groupi_n_4428);
  or csa_tree_add_6_33_groupi_g13802__9945(csa_tree_add_6_33_groupi_n_4483 ,csa_tree_add_6_33_groupi_n_4225 ,csa_tree_add_6_33_groupi_n_4432);
  xnor csa_tree_add_6_33_groupi_g13803__2883(csa_tree_add_6_33_groupi_n_4482 ,csa_tree_add_6_33_groupi_n_4330 ,csa_tree_add_6_33_groupi_n_4331);
  xnor csa_tree_add_6_33_groupi_g13804__2346(csa_tree_add_6_33_groupi_n_4481 ,csa_tree_add_6_33_groupi_n_4322 ,csa_tree_add_6_33_groupi_n_4104);
  xnor csa_tree_add_6_33_groupi_g13805__1666(csa_tree_add_6_33_groupi_n_4480 ,csa_tree_add_6_33_groupi_n_4284 ,csa_tree_add_6_33_groupi_n_4327);
  and csa_tree_add_6_33_groupi_g13806__7410(csa_tree_add_6_33_groupi_n_4513 ,csa_tree_add_6_33_groupi_n_4279 ,csa_tree_add_6_33_groupi_n_4439);
  and csa_tree_add_6_33_groupi_g13807__6417(csa_tree_add_6_33_groupi_n_4511 ,csa_tree_add_6_33_groupi_n_4306 ,csa_tree_add_6_33_groupi_n_4450);
  and csa_tree_add_6_33_groupi_g13808__5477(csa_tree_add_6_33_groupi_n_4510 ,csa_tree_add_6_33_groupi_n_4305 ,csa_tree_add_6_33_groupi_n_4449);
  and csa_tree_add_6_33_groupi_g13809__2398(csa_tree_add_6_33_groupi_n_4509 ,csa_tree_add_6_33_groupi_n_4316 ,csa_tree_add_6_33_groupi_n_4437);
  xnor csa_tree_add_6_33_groupi_g13810__5107(csa_tree_add_6_33_groupi_n_4508 ,csa_tree_add_6_33_groupi_n_4233 ,csa_tree_add_6_33_groupi_n_4299);
  xnor csa_tree_add_6_33_groupi_g13811__6260(csa_tree_add_6_33_groupi_n_4505 ,csa_tree_add_6_33_groupi_n_4290 ,csa_tree_add_6_33_groupi_n_4301);
  xnor csa_tree_add_6_33_groupi_g13812__4319(csa_tree_add_6_33_groupi_n_4504 ,csa_tree_add_6_33_groupi_n_4166 ,csa_tree_add_6_33_groupi_n_4300);
  xnor csa_tree_add_6_33_groupi_g13813__8428(csa_tree_add_6_33_groupi_n_4502 ,csa_tree_add_6_33_groupi_n_4224 ,csa_tree_add_6_33_groupi_n_4298);
  and csa_tree_add_6_33_groupi_g13814__5526(csa_tree_add_6_33_groupi_n_4501 ,csa_tree_add_6_33_groupi_n_4349 ,csa_tree_add_6_33_groupi_n_4453);
  xnor csa_tree_add_6_33_groupi_g13815__6783(csa_tree_add_6_33_groupi_n_4499 ,csa_tree_add_6_33_groupi_n_4337 ,csa_tree_add_6_33_groupi_n_4302);
  xnor csa_tree_add_6_33_groupi_g13816__3680(csa_tree_add_6_33_groupi_n_4498 ,csa_tree_add_6_33_groupi_n_4339 ,csa_tree_add_6_33_groupi_n_4295);
  xnor csa_tree_add_6_33_groupi_g13817__1617(csa_tree_add_6_33_groupi_n_4497 ,csa_tree_add_6_33_groupi_n_4169 ,csa_tree_add_6_33_groupi_n_4294);
  xnor csa_tree_add_6_33_groupi_g13818__2802(csa_tree_add_6_33_groupi_n_4496 ,csa_tree_add_6_33_groupi_n_4335 ,csa_tree_add_6_33_groupi_n_4293);
  xnor csa_tree_add_6_33_groupi_g13819__1705(csa_tree_add_6_33_groupi_n_4495 ,csa_tree_add_6_33_groupi_n_4334 ,csa_tree_add_6_33_groupi_n_4292);
  and csa_tree_add_6_33_groupi_g13820__5122(csa_tree_add_6_33_groupi_n_4493 ,csa_tree_add_6_33_groupi_n_4248 ,csa_tree_add_6_33_groupi_n_4409);
  xnor csa_tree_add_6_33_groupi_g13821__8246(csa_tree_add_6_33_groupi_n_4492 ,csa_tree_add_6_33_groupi_n_4035 ,csa_tree_add_6_33_groupi_n_4296);
  xnor csa_tree_add_6_33_groupi_g13822__7098(csa_tree_add_6_33_groupi_n_4491 ,csa_tree_add_6_33_groupi_n_4341 ,csa_tree_add_6_33_groupi_n_4297);
  not csa_tree_add_6_33_groupi_g13823(csa_tree_add_6_33_groupi_n_4470 ,csa_tree_add_6_33_groupi_n_4469);
  not csa_tree_add_6_33_groupi_g13824(csa_tree_add_6_33_groupi_n_4467 ,csa_tree_add_6_33_groupi_n_4468);
  not csa_tree_add_6_33_groupi_g13825(csa_tree_add_6_33_groupi_n_4463 ,csa_tree_add_6_33_groupi_n_4462);
  not csa_tree_add_6_33_groupi_g13826(csa_tree_add_6_33_groupi_n_4459 ,csa_tree_add_6_33_groupi_n_4460);
  and csa_tree_add_6_33_groupi_g13827__6131(csa_tree_add_6_33_groupi_n_4458 ,csa_tree_add_6_33_groupi_n_4104 ,csa_tree_add_6_33_groupi_n_4322);
  nor csa_tree_add_6_33_groupi_g13828__1881(csa_tree_add_6_33_groupi_n_4457 ,csa_tree_add_6_33_groupi_n_4085 ,csa_tree_add_6_33_groupi_n_4325);
  or csa_tree_add_6_33_groupi_g13829__5115(csa_tree_add_6_33_groupi_n_4456 ,csa_tree_add_6_33_groupi_n_4386 ,csa_tree_add_6_33_groupi_n_4373);
  and csa_tree_add_6_33_groupi_g13830__7482(csa_tree_add_6_33_groupi_n_4455 ,csa_tree_add_6_33_groupi_n_4165 ,csa_tree_add_6_33_groupi_n_4377);
  or csa_tree_add_6_33_groupi_g13831__4733(csa_tree_add_6_33_groupi_n_4454 ,csa_tree_add_6_33_groupi_n_4167 ,csa_tree_add_6_33_groupi_n_4314);
  or csa_tree_add_6_33_groupi_g13832__6161(csa_tree_add_6_33_groupi_n_4453 ,csa_tree_add_6_33_groupi_n_4333 ,csa_tree_add_6_33_groupi_n_4348);
  or csa_tree_add_6_33_groupi_g13833__9315(csa_tree_add_6_33_groupi_n_4452 ,csa_tree_add_6_33_groupi_n_4385 ,csa_tree_add_6_33_groupi_n_4360);
  and csa_tree_add_6_33_groupi_g13834__9945(csa_tree_add_6_33_groupi_n_4451 ,csa_tree_add_6_33_groupi_n_4331 ,csa_tree_add_6_33_groupi_n_4330);
  or csa_tree_add_6_33_groupi_g13835__2883(csa_tree_add_6_33_groupi_n_4450 ,csa_tree_add_6_33_groupi_n_4287 ,csa_tree_add_6_33_groupi_n_4309);
  or csa_tree_add_6_33_groupi_g13836__2346(csa_tree_add_6_33_groupi_n_4449 ,csa_tree_add_6_33_groupi_n_4336 ,csa_tree_add_6_33_groupi_n_4375);
  or csa_tree_add_6_33_groupi_g13837__1666(csa_tree_add_6_33_groupi_n_4448 ,csa_tree_add_6_33_groupi_n_4104 ,csa_tree_add_6_33_groupi_n_4322);
  or csa_tree_add_6_33_groupi_g13838__7410(csa_tree_add_6_33_groupi_n_4447 ,csa_tree_add_6_33_groupi_n_4278 ,csa_tree_add_6_33_groupi_n_4341);
  or csa_tree_add_6_33_groupi_g13839__6417(csa_tree_add_6_33_groupi_n_4446 ,csa_tree_add_6_33_groupi_n_4331 ,csa_tree_add_6_33_groupi_n_4330);
  or csa_tree_add_6_33_groupi_g13840__5477(csa_tree_add_6_33_groupi_n_4445 ,csa_tree_add_6_33_groupi_n_4084 ,csa_tree_add_6_33_groupi_n_4324);
  nor csa_tree_add_6_33_groupi_g13841__2398(csa_tree_add_6_33_groupi_n_4444 ,csa_tree_add_6_33_groupi_n_4283 ,csa_tree_add_6_33_groupi_n_4327);
  or csa_tree_add_6_33_groupi_g13842__5107(csa_tree_add_6_33_groupi_n_4443 ,csa_tree_add_6_33_groupi_n_4387 ,csa_tree_add_6_33_groupi_n_4371);
  or csa_tree_add_6_33_groupi_g13843__6260(csa_tree_add_6_33_groupi_n_4442 ,csa_tree_add_6_33_groupi_n_4291 ,csa_tree_add_6_33_groupi_n_4317);
  or csa_tree_add_6_33_groupi_g13844__4319(csa_tree_add_6_33_groupi_n_4441 ,csa_tree_add_6_33_groupi_n_4284 ,csa_tree_add_6_33_groupi_n_4326);
  or csa_tree_add_6_33_groupi_g13845__8428(csa_tree_add_6_33_groupi_n_4440 ,csa_tree_add_6_33_groupi_n_4240 ,csa_tree_add_6_33_groupi_n_4339);
  or csa_tree_add_6_33_groupi_g13846__5526(csa_tree_add_6_33_groupi_n_4439 ,csa_tree_add_6_33_groupi_n_4334 ,csa_tree_add_6_33_groupi_n_4282);
  or csa_tree_add_6_33_groupi_g13847__6783(csa_tree_add_6_33_groupi_n_4438 ,csa_tree_add_6_33_groupi_n_4238 ,csa_tree_add_6_33_groupi_n_4335);
  or csa_tree_add_6_33_groupi_g13848__3680(csa_tree_add_6_33_groupi_n_4437 ,csa_tree_add_6_33_groupi_n_4289 ,csa_tree_add_6_33_groupi_n_4310);
  and csa_tree_add_6_33_groupi_g13849__1617(csa_tree_add_6_33_groupi_n_4479 ,csa_tree_add_6_33_groupi_n_4253 ,csa_tree_add_6_33_groupi_n_4343);
  and csa_tree_add_6_33_groupi_g13850__2802(csa_tree_add_6_33_groupi_n_4478 ,csa_tree_add_6_33_groupi_n_4256 ,csa_tree_add_6_33_groupi_n_4347);
  and csa_tree_add_6_33_groupi_g13851__1705(csa_tree_add_6_33_groupi_n_4477 ,csa_tree_add_6_33_groupi_n_4192 ,csa_tree_add_6_33_groupi_n_4308);
  or csa_tree_add_6_33_groupi_g13852__5122(csa_tree_add_6_33_groupi_n_4476 ,csa_tree_add_6_33_groupi_n_3596 ,csa_tree_add_6_33_groupi_n_4304);
  and csa_tree_add_6_33_groupi_g13853__8246(csa_tree_add_6_33_groupi_n_4475 ,csa_tree_add_6_33_groupi_n_4263 ,csa_tree_add_6_33_groupi_n_4354);
  and csa_tree_add_6_33_groupi_g13854__7098(csa_tree_add_6_33_groupi_n_4474 ,csa_tree_add_6_33_groupi_n_4262 ,csa_tree_add_6_33_groupi_n_4353);
  and csa_tree_add_6_33_groupi_g13855__6131(csa_tree_add_6_33_groupi_n_4473 ,csa_tree_add_6_33_groupi_n_4246 ,csa_tree_add_6_33_groupi_n_4315);
  and csa_tree_add_6_33_groupi_g13856__1881(csa_tree_add_6_33_groupi_n_4472 ,csa_tree_add_6_33_groupi_n_4258 ,csa_tree_add_6_33_groupi_n_4313);
  and csa_tree_add_6_33_groupi_g13857__5115(csa_tree_add_6_33_groupi_n_4471 ,csa_tree_add_6_33_groupi_n_4195 ,csa_tree_add_6_33_groupi_n_4312);
  and csa_tree_add_6_33_groupi_g13858__7482(csa_tree_add_6_33_groupi_n_4469 ,csa_tree_add_6_33_groupi_n_4270 ,csa_tree_add_6_33_groupi_n_4365);
  and csa_tree_add_6_33_groupi_g13859__4733(csa_tree_add_6_33_groupi_n_4468 ,csa_tree_add_6_33_groupi_n_4197 ,csa_tree_add_6_33_groupi_n_4342);
  and csa_tree_add_6_33_groupi_g13860__6161(csa_tree_add_6_33_groupi_n_4466 ,csa_tree_add_6_33_groupi_n_4254 ,csa_tree_add_6_33_groupi_n_4344);
  and csa_tree_add_6_33_groupi_g13861__9315(csa_tree_add_6_33_groupi_n_4465 ,csa_tree_add_6_33_groupi_n_4267 ,csa_tree_add_6_33_groupi_n_4363);
  and csa_tree_add_6_33_groupi_g13862__9945(csa_tree_add_6_33_groupi_n_4464 ,csa_tree_add_6_33_groupi_n_4239 ,csa_tree_add_6_33_groupi_n_4319);
  and csa_tree_add_6_33_groupi_g13863__2883(csa_tree_add_6_33_groupi_n_4462 ,csa_tree_add_6_33_groupi_n_4272 ,csa_tree_add_6_33_groupi_n_4368);
  and csa_tree_add_6_33_groupi_g13864__2346(csa_tree_add_6_33_groupi_n_4461 ,csa_tree_add_6_33_groupi_n_4273 ,csa_tree_add_6_33_groupi_n_4367);
  and csa_tree_add_6_33_groupi_g13865__1666(csa_tree_add_6_33_groupi_n_4460 ,csa_tree_add_6_33_groupi_n_4131 ,csa_tree_add_6_33_groupi_n_4369);
  not csa_tree_add_6_33_groupi_g13866(csa_tree_add_6_33_groupi_n_4433 ,csa_tree_add_6_33_groupi_n_4432);
  not csa_tree_add_6_33_groupi_g13867(csa_tree_add_6_33_groupi_n_4429 ,csa_tree_add_6_33_groupi_n_4430);
  not csa_tree_add_6_33_groupi_g13868(csa_tree_add_6_33_groupi_n_4427 ,csa_tree_add_6_33_groupi_n_4426);
  not csa_tree_add_6_33_groupi_g13869(csa_tree_add_6_33_groupi_n_4422 ,csa_tree_add_6_33_groupi_n_4423);
  not csa_tree_add_6_33_groupi_g13870(csa_tree_add_6_33_groupi_n_4421 ,csa_tree_add_6_33_groupi_n_4420);
  not csa_tree_add_6_33_groupi_g13871(csa_tree_add_6_33_groupi_n_4419 ,csa_tree_add_6_33_groupi_n_4418);
  not csa_tree_add_6_33_groupi_g13872(csa_tree_add_6_33_groupi_n_4416 ,csa_tree_add_6_33_groupi_n_4417);
  not csa_tree_add_6_33_groupi_g13873(csa_tree_add_6_33_groupi_n_4415 ,csa_tree_add_6_33_groupi_n_4414);
  not csa_tree_add_6_33_groupi_g13874(csa_tree_add_6_33_groupi_n_4412 ,csa_tree_add_6_33_groupi_n_4413);
  xnor csa_tree_add_6_33_groupi_g13875__7410(out1[6] ,csa_tree_add_6_33_groupi_n_4288 ,csa_tree_add_6_33_groupi_n_3797);
  or csa_tree_add_6_33_groupi_g13876__6417(csa_tree_add_6_33_groupi_n_4409 ,csa_tree_add_6_33_groupi_n_4247 ,csa_tree_add_6_33_groupi_n_4338);
  xnor csa_tree_add_6_33_groupi_g13877__5477(csa_tree_add_6_33_groupi_n_4408 ,csa_tree_add_6_33_groupi_n_4147 ,csa_tree_add_6_33_groupi_n_4213);
  xnor csa_tree_add_6_33_groupi_g13878__2398(csa_tree_add_6_33_groupi_n_4407 ,csa_tree_add_6_33_groupi_n_4160 ,csa_tree_add_6_33_groupi_n_4232);
  xnor csa_tree_add_6_33_groupi_g13879__5107(csa_tree_add_6_33_groupi_n_4406 ,csa_tree_add_6_33_groupi_n_4203 ,csa_tree_add_6_33_groupi_n_3842);
  xnor csa_tree_add_6_33_groupi_g13880__6260(csa_tree_add_6_33_groupi_n_4405 ,csa_tree_add_6_33_groupi_n_4205 ,csa_tree_add_6_33_groupi_n_4013);
  xnor csa_tree_add_6_33_groupi_g13881__4319(csa_tree_add_6_33_groupi_n_4404 ,csa_tree_add_6_33_groupi_n_4153 ,csa_tree_add_6_33_groupi_n_4221);
  xnor csa_tree_add_6_33_groupi_g13882__8428(csa_tree_add_6_33_groupi_n_4403 ,csa_tree_add_6_33_groupi_n_4157 ,csa_tree_add_6_33_groupi_n_4207);
  xnor csa_tree_add_6_33_groupi_g13883__5526(csa_tree_add_6_33_groupi_n_4402 ,csa_tree_add_6_33_groupi_n_4208 ,csa_tree_add_6_33_groupi_n_4148);
  xnor csa_tree_add_6_33_groupi_g13884__6783(csa_tree_add_6_33_groupi_n_4401 ,csa_tree_add_6_33_groupi_n_4204 ,csa_tree_add_6_33_groupi_n_4285);
  xnor csa_tree_add_6_33_groupi_g13885__3680(csa_tree_add_6_33_groupi_n_4400 ,csa_tree_add_6_33_groupi_n_4085 ,csa_tree_add_6_33_groupi_n_4286);
  xnor csa_tree_add_6_33_groupi_g13886__1617(csa_tree_add_6_33_groupi_n_4399 ,csa_tree_add_6_33_groupi_n_4066 ,csa_tree_add_6_33_groupi_n_4230);
  xnor csa_tree_add_6_33_groupi_g13887__2802(csa_tree_add_6_33_groupi_n_4398 ,csa_tree_add_6_33_groupi_n_4071 ,csa_tree_add_6_33_groupi_n_4228);
  xnor csa_tree_add_6_33_groupi_g13888__1705(csa_tree_add_6_33_groupi_n_4397 ,csa_tree_add_6_33_groupi_n_4235 ,csa_tree_add_6_33_groupi_n_3965);
  xnor csa_tree_add_6_33_groupi_g13889__5122(csa_tree_add_6_33_groupi_n_4396 ,csa_tree_add_6_33_groupi_n_4211 ,csa_tree_add_6_33_groupi_n_4151);
  xnor csa_tree_add_6_33_groupi_g13890__8246(csa_tree_add_6_33_groupi_n_4395 ,csa_tree_add_6_33_groupi_n_4218 ,csa_tree_add_6_33_groupi_n_4068);
  xnor csa_tree_add_6_33_groupi_g13891__7098(csa_tree_add_6_33_groupi_n_4394 ,csa_tree_add_6_33_groupi_n_4215 ,csa_tree_add_6_33_groupi_n_4155);
  xnor csa_tree_add_6_33_groupi_g13892__6131(csa_tree_add_6_33_groupi_n_4393 ,csa_tree_add_6_33_groupi_n_4075 ,csa_tree_add_6_33_groupi_n_4223);
  xnor csa_tree_add_6_33_groupi_g13893__1881(csa_tree_add_6_33_groupi_n_4392 ,csa_tree_add_6_33_groupi_n_4201 ,csa_tree_add_6_33_groupi_n_4096);
  xnor csa_tree_add_6_33_groupi_g13894__5115(csa_tree_add_6_33_groupi_n_4391 ,csa_tree_add_6_33_groupi_n_4217 ,csa_tree_add_6_33_groupi_n_4158);
  xnor csa_tree_add_6_33_groupi_g13895__7482(csa_tree_add_6_33_groupi_n_4390 ,csa_tree_add_6_33_groupi_n_3964 ,csa_tree_add_6_33_groupi_n_4210);
  xnor csa_tree_add_6_33_groupi_g13896__4733(csa_tree_add_6_33_groupi_n_4389 ,csa_tree_add_6_33_groupi_n_4216 ,csa_tree_add_6_33_groupi_n_4161);
  xnor csa_tree_add_6_33_groupi_g13897__6161(csa_tree_add_6_33_groupi_n_4388 ,csa_tree_add_6_33_groupi_n_4028 ,csa_tree_add_6_33_groupi_n_4214);
  xnor csa_tree_add_6_33_groupi_g13898__9315(csa_tree_add_6_33_groupi_n_4436 ,csa_tree_add_6_33_groupi_n_4109 ,csa_tree_add_6_33_groupi_n_4184);
  xnor csa_tree_add_6_33_groupi_g13899__9945(csa_tree_add_6_33_groupi_n_4435 ,csa_tree_add_6_33_groupi_n_4111 ,csa_tree_add_6_33_groupi_n_4188);
  xnor csa_tree_add_6_33_groupi_g13900__2883(csa_tree_add_6_33_groupi_n_4434 ,csa_tree_add_6_33_groupi_n_4044 ,csa_tree_add_6_33_groupi_n_4173);
  xnor csa_tree_add_6_33_groupi_g13901__2346(csa_tree_add_6_33_groupi_n_4432 ,csa_tree_add_6_33_groupi_n_4093 ,csa_tree_add_6_33_groupi_n_4178);
  xnor csa_tree_add_6_33_groupi_g13902__1666(csa_tree_add_6_33_groupi_n_4431 ,csa_tree_add_6_33_groupi_n_4079 ,csa_tree_add_6_33_groupi_n_4183);
  xnor csa_tree_add_6_33_groupi_g13903__7410(csa_tree_add_6_33_groupi_n_4430 ,csa_tree_add_6_33_groupi_n_3983 ,csa_tree_add_6_33_groupi_n_4175);
  xnor csa_tree_add_6_33_groupi_g13904__6417(csa_tree_add_6_33_groupi_n_4428 ,csa_tree_add_6_33_groupi_n_4091 ,csa_tree_add_6_33_groupi_n_0);
  xnor csa_tree_add_6_33_groupi_g13905__5477(csa_tree_add_6_33_groupi_n_4426 ,csa_tree_add_6_33_groupi_n_4083 ,csa_tree_add_6_33_groupi_n_4185);
  xnor csa_tree_add_6_33_groupi_g13906__2398(csa_tree_add_6_33_groupi_n_4425 ,csa_tree_add_6_33_groupi_n_4105 ,csa_tree_add_6_33_groupi_n_4172);
  xnor csa_tree_add_6_33_groupi_g13907__5107(csa_tree_add_6_33_groupi_n_4424 ,csa_tree_add_6_33_groupi_n_4107 ,csa_tree_add_6_33_groupi_n_4186);
  xnor csa_tree_add_6_33_groupi_g13908__6260(csa_tree_add_6_33_groupi_n_4423 ,csa_tree_add_6_33_groupi_n_4110 ,csa_tree_add_6_33_groupi_n_4174);
  xnor csa_tree_add_6_33_groupi_g13909__4319(csa_tree_add_6_33_groupi_n_4420 ,csa_tree_add_6_33_groupi_n_4089 ,csa_tree_add_6_33_groupi_n_4187);
  xnor csa_tree_add_6_33_groupi_g13910__8428(csa_tree_add_6_33_groupi_n_4418 ,csa_tree_add_6_33_groupi_n_4082 ,csa_tree_add_6_33_groupi_n_4177);
  xnor csa_tree_add_6_33_groupi_g13911__5526(csa_tree_add_6_33_groupi_n_4417 ,csa_tree_add_6_33_groupi_n_3847 ,csa_tree_add_6_33_groupi_n_4189);
  xnor csa_tree_add_6_33_groupi_g13912__6783(csa_tree_add_6_33_groupi_n_4414 ,csa_tree_add_6_33_groupi_n_4164 ,csa_tree_add_6_33_groupi_n_4179);
  xnor csa_tree_add_6_33_groupi_g13913__3680(csa_tree_add_6_33_groupi_n_4413 ,csa_tree_add_6_33_groupi_n_4098 ,csa_tree_add_6_33_groupi_n_4171);
  xnor csa_tree_add_6_33_groupi_g13914__1617(csa_tree_add_6_33_groupi_n_4411 ,csa_tree_add_6_33_groupi_n_3962 ,csa_tree_add_6_33_groupi_n_4176);
  not csa_tree_add_6_33_groupi_g13915(csa_tree_add_6_33_groupi_n_4383 ,csa_tree_add_6_33_groupi_n_4384);
  and csa_tree_add_6_33_groupi_g13916__2802(csa_tree_add_6_33_groupi_n_4380 ,csa_tree_add_6_33_groupi_n_4096 ,csa_tree_add_6_33_groupi_n_4201);
  or csa_tree_add_6_33_groupi_g13917__1705(csa_tree_add_6_33_groupi_n_4379 ,csa_tree_add_6_33_groupi_n_4147 ,csa_tree_add_6_33_groupi_n_4212);
  nor csa_tree_add_6_33_groupi_g13918__5122(csa_tree_add_6_33_groupi_n_4378 ,csa_tree_add_6_33_groupi_n_4065 ,csa_tree_add_6_33_groupi_n_4230);
  or csa_tree_add_6_33_groupi_g13919__8246(csa_tree_add_6_33_groupi_n_4377 ,csa_tree_add_6_33_groupi_n_4066 ,csa_tree_add_6_33_groupi_n_4229);
  and csa_tree_add_6_33_groupi_g13920__7098(csa_tree_add_6_33_groupi_n_4376 ,csa_tree_add_6_33_groupi_n_4148 ,csa_tree_add_6_33_groupi_n_4208);
  and csa_tree_add_6_33_groupi_g13921__6131(csa_tree_add_6_33_groupi_n_4375 ,csa_tree_add_6_33_groupi_n_4068 ,csa_tree_add_6_33_groupi_n_4218);
  or csa_tree_add_6_33_groupi_g13922__1881(csa_tree_add_6_33_groupi_n_4374 ,csa_tree_add_6_33_groupi_n_4074 ,csa_tree_add_6_33_groupi_n_4223);
  nor csa_tree_add_6_33_groupi_g13923__5115(csa_tree_add_6_33_groupi_n_4373 ,csa_tree_add_6_33_groupi_n_4146 ,csa_tree_add_6_33_groupi_n_4213);
  or csa_tree_add_6_33_groupi_g13924__7482(csa_tree_add_6_33_groupi_n_4372 ,csa_tree_add_6_33_groupi_n_4153 ,csa_tree_add_6_33_groupi_n_4220);
  and csa_tree_add_6_33_groupi_g13925__4733(csa_tree_add_6_33_groupi_n_4371 ,csa_tree_add_6_33_groupi_n_4013 ,csa_tree_add_6_33_groupi_n_4205);
  or csa_tree_add_6_33_groupi_g13926__6161(csa_tree_add_6_33_groupi_n_4370 ,csa_tree_add_6_33_groupi_n_4155 ,csa_tree_add_6_33_groupi_n_4215);
  or csa_tree_add_6_33_groupi_g13927__9315(csa_tree_add_6_33_groupi_n_4369 ,csa_tree_add_6_33_groupi_n_4129 ,csa_tree_add_6_33_groupi_n_4235);
  or csa_tree_add_6_33_groupi_g13928__9945(csa_tree_add_6_33_groupi_n_4368 ,csa_tree_add_6_33_groupi_n_4030 ,csa_tree_add_6_33_groupi_n_4271);
  or csa_tree_add_6_33_groupi_g13929__2883(csa_tree_add_6_33_groupi_n_4367 ,csa_tree_add_6_33_groupi_n_4035 ,csa_tree_add_6_33_groupi_n_4257);
  and csa_tree_add_6_33_groupi_g13930__2346(csa_tree_add_6_33_groupi_n_4366 ,csa_tree_add_6_33_groupi_n_4155 ,csa_tree_add_6_33_groupi_n_4215);
  or csa_tree_add_6_33_groupi_g13931__1666(csa_tree_add_6_33_groupi_n_4365 ,csa_tree_add_6_33_groupi_n_4031 ,csa_tree_add_6_33_groupi_n_4269);
  or csa_tree_add_6_33_groupi_g13932__7410(csa_tree_add_6_33_groupi_n_4364 ,csa_tree_add_6_33_groupi_n_3842 ,csa_tree_add_6_33_groupi_n_4203);
  or csa_tree_add_6_33_groupi_g13933__6417(csa_tree_add_6_33_groupi_n_4363 ,csa_tree_add_6_33_groupi_n_4033 ,csa_tree_add_6_33_groupi_n_4266);
  or csa_tree_add_6_33_groupi_g13934__5477(csa_tree_add_6_33_groupi_n_4362 ,csa_tree_add_6_33_groupi_n_4013 ,csa_tree_add_6_33_groupi_n_4205);
  or csa_tree_add_6_33_groupi_g13935__2398(csa_tree_add_6_33_groupi_n_4361 ,csa_tree_add_6_33_groupi_n_4158 ,csa_tree_add_6_33_groupi_n_4217);
  nor csa_tree_add_6_33_groupi_g13936__5107(csa_tree_add_6_33_groupi_n_4360 ,csa_tree_add_6_33_groupi_n_4075 ,csa_tree_add_6_33_groupi_n_4222);
  or csa_tree_add_6_33_groupi_g13937__6260(csa_tree_add_6_33_groupi_n_4359 ,csa_tree_add_6_33_groupi_n_4160 ,csa_tree_add_6_33_groupi_n_4231);
  and csa_tree_add_6_33_groupi_g13938__4319(csa_tree_add_6_33_groupi_n_4358 ,csa_tree_add_6_33_groupi_n_4158 ,csa_tree_add_6_33_groupi_n_4217);
  or csa_tree_add_6_33_groupi_g13939__8428(csa_tree_add_6_33_groupi_n_4357 ,csa_tree_add_6_33_groupi_n_4161 ,csa_tree_add_6_33_groupi_n_4216);
  and csa_tree_add_6_33_groupi_g13940__5526(csa_tree_add_6_33_groupi_n_4356 ,csa_tree_add_6_33_groupi_n_4161 ,csa_tree_add_6_33_groupi_n_4216);
  nor csa_tree_add_6_33_groupi_g13941__6783(csa_tree_add_6_33_groupi_n_4355 ,csa_tree_add_6_33_groupi_n_4159 ,csa_tree_add_6_33_groupi_n_4232);
  or csa_tree_add_6_33_groupi_g13942__3680(csa_tree_add_6_33_groupi_n_4354 ,csa_tree_add_6_33_groupi_n_4036 ,csa_tree_add_6_33_groupi_n_4259);
  or csa_tree_add_6_33_groupi_g13943__1617(csa_tree_add_6_33_groupi_n_4353 ,csa_tree_add_6_33_groupi_n_4038 ,csa_tree_add_6_33_groupi_n_4261);
  nor csa_tree_add_6_33_groupi_g13944__2802(csa_tree_add_6_33_groupi_n_4352 ,csa_tree_add_6_33_groupi_n_4148 ,csa_tree_add_6_33_groupi_n_4208);
  nor csa_tree_add_6_33_groupi_g13945__1705(csa_tree_add_6_33_groupi_n_4351 ,csa_tree_add_6_33_groupi_n_4152 ,csa_tree_add_6_33_groupi_n_4221);
  or csa_tree_add_6_33_groupi_g13946__5122(csa_tree_add_6_33_groupi_n_4350 ,csa_tree_add_6_33_groupi_n_4285 ,csa_tree_add_6_33_groupi_n_4204);
  or csa_tree_add_6_33_groupi_g13947__8246(csa_tree_add_6_33_groupi_n_4349 ,csa_tree_add_6_33_groupi_n_4157 ,csa_tree_add_6_33_groupi_n_4206);
  nor csa_tree_add_6_33_groupi_g13948__7098(csa_tree_add_6_33_groupi_n_4348 ,csa_tree_add_6_33_groupi_n_4156 ,csa_tree_add_6_33_groupi_n_4207);
  or csa_tree_add_6_33_groupi_g13949__6131(csa_tree_add_6_33_groupi_n_4347 ,csa_tree_add_6_33_groupi_n_4029 ,csa_tree_add_6_33_groupi_n_4255);
  or csa_tree_add_6_33_groupi_g13950__1881(csa_tree_add_6_33_groupi_n_4346 ,csa_tree_add_6_33_groupi_n_4151 ,csa_tree_add_6_33_groupi_n_4211);
  and csa_tree_add_6_33_groupi_g13951__5115(csa_tree_add_6_33_groupi_n_4345 ,csa_tree_add_6_33_groupi_n_4151 ,csa_tree_add_6_33_groupi_n_4211);
  or csa_tree_add_6_33_groupi_g13952__7482(csa_tree_add_6_33_groupi_n_4344 ,csa_tree_add_6_33_groupi_n_4290 ,csa_tree_add_6_33_groupi_n_4250);
  or csa_tree_add_6_33_groupi_g13953__4733(csa_tree_add_6_33_groupi_n_4343 ,csa_tree_add_6_33_groupi_n_4042 ,csa_tree_add_6_33_groupi_n_4251);
  or csa_tree_add_6_33_groupi_g13954__6161(csa_tree_add_6_33_groupi_n_4342 ,csa_tree_add_6_33_groupi_n_3920 ,csa_tree_add_6_33_groupi_n_4196);
  and csa_tree_add_6_33_groupi_g13955__9315(csa_tree_add_6_33_groupi_n_4387 ,csa_tree_add_6_33_groupi_n_4112 ,csa_tree_add_6_33_groupi_n_4249);
  and csa_tree_add_6_33_groupi_g13956__9945(csa_tree_add_6_33_groupi_n_4386 ,csa_tree_add_6_33_groupi_n_4138 ,csa_tree_add_6_33_groupi_n_4275);
  and csa_tree_add_6_33_groupi_g13957__2883(csa_tree_add_6_33_groupi_n_4385 ,csa_tree_add_6_33_groupi_n_3889 ,csa_tree_add_6_33_groupi_n_4268);
  and csa_tree_add_6_33_groupi_g13958__2346(csa_tree_add_6_33_groupi_n_4384 ,csa_tree_add_6_33_groupi_n_4116 ,csa_tree_add_6_33_groupi_n_4244);
  and csa_tree_add_6_33_groupi_g13959__1666(csa_tree_add_6_33_groupi_n_4382 ,csa_tree_add_6_33_groupi_n_4128 ,csa_tree_add_6_33_groupi_n_4264);
  and csa_tree_add_6_33_groupi_g13960__7410(csa_tree_add_6_33_groupi_n_4381 ,csa_tree_add_6_33_groupi_n_4057 ,csa_tree_add_6_33_groupi_n_4265);
  not csa_tree_add_6_33_groupi_g13961(csa_tree_add_6_33_groupi_n_4338 ,csa_tree_add_6_33_groupi_n_4337);
  not csa_tree_add_6_33_groupi_g13962(csa_tree_add_6_33_groupi_n_4333 ,csa_tree_add_6_33_groupi_n_4332);
  not csa_tree_add_6_33_groupi_g13963(csa_tree_add_6_33_groupi_n_4329 ,csa_tree_add_6_33_groupi_n_4328);
  not csa_tree_add_6_33_groupi_g13964(csa_tree_add_6_33_groupi_n_4326 ,csa_tree_add_6_33_groupi_n_4327);
  not csa_tree_add_6_33_groupi_g13965(csa_tree_add_6_33_groupi_n_4324 ,csa_tree_add_6_33_groupi_n_4325);
  and csa_tree_add_6_33_groupi_g13966__6417(csa_tree_add_6_33_groupi_n_4321 ,csa_tree_add_6_33_groupi_n_4285 ,csa_tree_add_6_33_groupi_n_4204);
  or csa_tree_add_6_33_groupi_g13967__5477(csa_tree_add_6_33_groupi_n_4320 ,csa_tree_add_6_33_groupi_n_4028 ,csa_tree_add_6_33_groupi_n_4214);
  or csa_tree_add_6_33_groupi_g13968__2398(csa_tree_add_6_33_groupi_n_4319 ,csa_tree_add_6_33_groupi_n_4170 ,csa_tree_add_6_33_groupi_n_4236);
  and csa_tree_add_6_33_groupi_g13969__5107(csa_tree_add_6_33_groupi_n_4318 ,csa_tree_add_6_33_groupi_n_4028 ,csa_tree_add_6_33_groupi_n_4214);
  and csa_tree_add_6_33_groupi_g13970__6260(csa_tree_add_6_33_groupi_n_4317 ,csa_tree_add_6_33_groupi_n_3842 ,csa_tree_add_6_33_groupi_n_4203);
  or csa_tree_add_6_33_groupi_g13971__4319(csa_tree_add_6_33_groupi_n_4316 ,csa_tree_add_6_33_groupi_n_3964 ,csa_tree_add_6_33_groupi_n_4209);
  or csa_tree_add_6_33_groupi_g13972__8428(csa_tree_add_6_33_groupi_n_4315 ,csa_tree_add_6_33_groupi_n_4252 ,csa_tree_add_6_33_groupi_n_4234);
  and csa_tree_add_6_33_groupi_g13973__5526(csa_tree_add_6_33_groupi_n_4314 ,csa_tree_add_6_33_groupi_n_3913 ,csa_tree_add_6_33_groupi_n_4224);
  or csa_tree_add_6_33_groupi_g13974__6783(csa_tree_add_6_33_groupi_n_4313 ,csa_tree_add_6_33_groupi_n_4166 ,csa_tree_add_6_33_groupi_n_4260);
  or csa_tree_add_6_33_groupi_g13975__3680(csa_tree_add_6_33_groupi_n_4312 ,csa_tree_add_6_33_groupi_n_4037 ,csa_tree_add_6_33_groupi_n_4194);
  or csa_tree_add_6_33_groupi_g13976__1617(csa_tree_add_6_33_groupi_n_4311 ,csa_tree_add_6_33_groupi_n_3913 ,csa_tree_add_6_33_groupi_n_4224);
  nor csa_tree_add_6_33_groupi_g13977__2802(csa_tree_add_6_33_groupi_n_4310 ,csa_tree_add_6_33_groupi_n_3963 ,csa_tree_add_6_33_groupi_n_4210);
  nor csa_tree_add_6_33_groupi_g13978__1705(csa_tree_add_6_33_groupi_n_4309 ,csa_tree_add_6_33_groupi_n_4070 ,csa_tree_add_6_33_groupi_n_4228);
  or csa_tree_add_6_33_groupi_g13979__5122(csa_tree_add_6_33_groupi_n_4308 ,csa_tree_add_6_33_groupi_n_3848 ,csa_tree_add_6_33_groupi_n_4200);
  nor csa_tree_add_6_33_groupi_g13980__8246(csa_tree_add_6_33_groupi_n_4307 ,csa_tree_add_6_33_groupi_n_4096 ,csa_tree_add_6_33_groupi_n_4201);
  or csa_tree_add_6_33_groupi_g13981__7098(csa_tree_add_6_33_groupi_n_4306 ,csa_tree_add_6_33_groupi_n_4071 ,csa_tree_add_6_33_groupi_n_4227);
  or csa_tree_add_6_33_groupi_g13982__6131(csa_tree_add_6_33_groupi_n_4305 ,csa_tree_add_6_33_groupi_n_4068 ,csa_tree_add_6_33_groupi_n_4218);
  and csa_tree_add_6_33_groupi_g13983__1881(csa_tree_add_6_33_groupi_n_4304 ,csa_tree_add_6_33_groupi_n_3597 ,csa_tree_add_6_33_groupi_n_4288);
  xnor csa_tree_add_6_33_groupi_g13984__5115(csa_tree_add_6_33_groupi_n_4303 ,csa_tree_add_6_33_groupi_n_4067 ,csa_tree_add_6_33_groupi_n_4144);
  xnor csa_tree_add_6_33_groupi_g13985__7482(csa_tree_add_6_33_groupi_n_4302 ,csa_tree_add_6_33_groupi_n_3978 ,csa_tree_add_6_33_groupi_n_4078);
  xnor csa_tree_add_6_33_groupi_g13986__4733(csa_tree_add_6_33_groupi_n_4301 ,csa_tree_add_6_33_groupi_n_3631 ,csa_tree_add_6_33_groupi_n_4081);
  xnor csa_tree_add_6_33_groupi_g13987__6161(csa_tree_add_6_33_groupi_n_4300 ,csa_tree_add_6_33_groupi_n_4015 ,csa_tree_add_6_33_groupi_n_4087);
  xnor csa_tree_add_6_33_groupi_g13988__9315(csa_tree_add_6_33_groupi_n_4299 ,csa_tree_add_6_33_groupi_n_4076 ,csa_tree_add_6_33_groupi_n_4011);
  xnor csa_tree_add_6_33_groupi_g13989__9945(csa_tree_add_6_33_groupi_n_4298 ,csa_tree_add_6_33_groupi_n_4167 ,csa_tree_add_6_33_groupi_n_3913);
  xnor csa_tree_add_6_33_groupi_g13990__2883(csa_tree_add_6_33_groupi_n_4297 ,csa_tree_add_6_33_groupi_n_4072 ,csa_tree_add_6_33_groupi_n_3836);
  xnor csa_tree_add_6_33_groupi_g13991__2346(csa_tree_add_6_33_groupi_n_4296 ,csa_tree_add_6_33_groupi_n_4103 ,csa_tree_add_6_33_groupi_n_3536);
  xnor csa_tree_add_6_33_groupi_g13992__1666(csa_tree_add_6_33_groupi_n_4295 ,csa_tree_add_6_33_groupi_n_3976 ,csa_tree_add_6_33_groupi_n_4095);
  xnor csa_tree_add_6_33_groupi_g13993__7410(csa_tree_add_6_33_groupi_n_4294 ,csa_tree_add_6_33_groupi_n_3967 ,csa_tree_add_6_33_groupi_n_4102);
  xnor csa_tree_add_6_33_groupi_g13994__6417(csa_tree_add_6_33_groupi_n_4293 ,csa_tree_add_6_33_groupi_n_4073 ,csa_tree_add_6_33_groupi_n_4009);
  xnor csa_tree_add_6_33_groupi_g13995__5477(csa_tree_add_6_33_groupi_n_4292 ,csa_tree_add_6_33_groupi_n_4069 ,csa_tree_add_6_33_groupi_n_4145);
  and csa_tree_add_6_33_groupi_g13996__2398(csa_tree_add_6_33_groupi_n_4341 ,csa_tree_add_6_33_groupi_n_4135 ,csa_tree_add_6_33_groupi_n_4276);
  and csa_tree_add_6_33_groupi_g13997__5107(csa_tree_add_6_33_groupi_n_4340 ,csa_tree_add_6_33_groupi_n_4125 ,csa_tree_add_6_33_groupi_n_4241);
  xnor csa_tree_add_6_33_groupi_g13998__6260(csa_tree_add_6_33_groupi_n_4339 ,csa_tree_add_6_33_groupi_n_4010 ,csa_tree_add_6_33_groupi_n_4049);
  xnor csa_tree_add_6_33_groupi_g13999__4319(csa_tree_add_6_33_groupi_n_4337 ,csa_tree_add_6_33_groupi_n_4012 ,csa_tree_add_6_33_groupi_n_4051);
  and csa_tree_add_6_33_groupi_g14000__8428(csa_tree_add_6_33_groupi_n_4336 ,csa_tree_add_6_33_groupi_n_4059 ,csa_tree_add_6_33_groupi_n_4277);
  and csa_tree_add_6_33_groupi_g14001__5526(csa_tree_add_6_33_groupi_n_4335 ,csa_tree_add_6_33_groupi_n_4124 ,csa_tree_add_6_33_groupi_n_4237);
  and csa_tree_add_6_33_groupi_g14002__6783(csa_tree_add_6_33_groupi_n_4334 ,csa_tree_add_6_33_groupi_n_4063 ,csa_tree_add_6_33_groupi_n_4199);
  or csa_tree_add_6_33_groupi_g14003__3680(csa_tree_add_6_33_groupi_n_4332 ,csa_tree_add_6_33_groupi_n_4122 ,csa_tree_add_6_33_groupi_n_4198);
  and csa_tree_add_6_33_groupi_g14004__1617(csa_tree_add_6_33_groupi_n_4331 ,csa_tree_add_6_33_groupi_n_4060 ,csa_tree_add_6_33_groupi_n_4280);
  xnor csa_tree_add_6_33_groupi_g14005__2802(csa_tree_add_6_33_groupi_n_4330 ,csa_tree_add_6_33_groupi_n_3846 ,csa_tree_add_6_33_groupi_n_4048);
  xnor csa_tree_add_6_33_groupi_g14006__1705(csa_tree_add_6_33_groupi_n_4328 ,csa_tree_add_6_33_groupi_n_4100 ,csa_tree_add_6_33_groupi_n_4047);
  xnor csa_tree_add_6_33_groupi_g14007__5122(csa_tree_add_6_33_groupi_n_4327 ,csa_tree_add_6_33_groupi_n_3918 ,csa_tree_add_6_33_groupi_n_4045);
  xnor csa_tree_add_6_33_groupi_g14008__8246(csa_tree_add_6_33_groupi_n_4325 ,csa_tree_add_6_33_groupi_n_3982 ,csa_tree_add_6_33_groupi_n_4050);
  and csa_tree_add_6_33_groupi_g14009__7098(csa_tree_add_6_33_groupi_n_4323 ,csa_tree_add_6_33_groupi_n_4140 ,csa_tree_add_6_33_groupi_n_4193);
  xnor csa_tree_add_6_33_groupi_g14010__6131(csa_tree_add_6_33_groupi_n_4322 ,csa_tree_add_6_33_groupi_n_4168 ,csa_tree_add_6_33_groupi_n_3929);
  not csa_tree_add_6_33_groupi_g14011(csa_tree_add_6_33_groupi_n_4283 ,csa_tree_add_6_33_groupi_n_4284);
  and csa_tree_add_6_33_groupi_g14012__1881(csa_tree_add_6_33_groupi_n_4282 ,csa_tree_add_6_33_groupi_n_4145 ,csa_tree_add_6_33_groupi_n_4069);
  or csa_tree_add_6_33_groupi_g14013__5115(csa_tree_add_6_33_groupi_n_4281 ,csa_tree_add_6_33_groupi_n_3836 ,csa_tree_add_6_33_groupi_n_4072);
  or csa_tree_add_6_33_groupi_g14014__7482(csa_tree_add_6_33_groupi_n_4280 ,csa_tree_add_6_33_groupi_n_4164 ,csa_tree_add_6_33_groupi_n_4134);
  or csa_tree_add_6_33_groupi_g14015__4733(csa_tree_add_6_33_groupi_n_4279 ,csa_tree_add_6_33_groupi_n_4145 ,csa_tree_add_6_33_groupi_n_4069);
  and csa_tree_add_6_33_groupi_g14016__6161(csa_tree_add_6_33_groupi_n_4278 ,csa_tree_add_6_33_groupi_n_3836 ,csa_tree_add_6_33_groupi_n_4072);
  or csa_tree_add_6_33_groupi_g14017__9315(csa_tree_add_6_33_groupi_n_4277 ,csa_tree_add_6_33_groupi_n_3766 ,csa_tree_add_6_33_groupi_n_4136);
  or csa_tree_add_6_33_groupi_g14018__9945(csa_tree_add_6_33_groupi_n_4276 ,csa_tree_add_6_33_groupi_n_4034 ,csa_tree_add_6_33_groupi_n_4142);
  or csa_tree_add_6_33_groupi_g14019__2883(csa_tree_add_6_33_groupi_n_4275 ,csa_tree_add_6_33_groupi_n_4044 ,csa_tree_add_6_33_groupi_n_4133);
  and csa_tree_add_6_33_groupi_g14020__2346(csa_tree_add_6_33_groupi_n_4274 ,csa_tree_add_6_33_groupi_n_4144 ,csa_tree_add_6_33_groupi_n_4067);
  or csa_tree_add_6_33_groupi_g14021__1666(csa_tree_add_6_33_groupi_n_4273 ,csa_tree_add_6_33_groupi_n_3536 ,csa_tree_add_6_33_groupi_n_4103);
  or csa_tree_add_6_33_groupi_g14022__7410(csa_tree_add_6_33_groupi_n_4272 ,csa_tree_add_6_33_groupi_n_3955 ,csa_tree_add_6_33_groupi_n_4088);
  nor csa_tree_add_6_33_groupi_g14023__6417(csa_tree_add_6_33_groupi_n_4271 ,csa_tree_add_6_33_groupi_n_3956 ,csa_tree_add_6_33_groupi_n_4089);
  or csa_tree_add_6_33_groupi_g14024__5477(csa_tree_add_6_33_groupi_n_4270 ,csa_tree_add_6_33_groupi_n_3654 ,csa_tree_add_6_33_groupi_n_4106);
  nor csa_tree_add_6_33_groupi_g14025__2398(csa_tree_add_6_33_groupi_n_4269 ,csa_tree_add_6_33_groupi_n_3655 ,csa_tree_add_6_33_groupi_n_4107);
  or csa_tree_add_6_33_groupi_g14026__5107(csa_tree_add_6_33_groupi_n_4268 ,csa_tree_add_6_33_groupi_n_3882 ,csa_tree_add_6_33_groupi_n_4168);
  or csa_tree_add_6_33_groupi_g14027__6260(csa_tree_add_6_33_groupi_n_4267 ,csa_tree_add_6_33_groupi_n_3652 ,csa_tree_add_6_33_groupi_n_4105);
  and csa_tree_add_6_33_groupi_g14028__4319(csa_tree_add_6_33_groupi_n_4266 ,csa_tree_add_6_33_groupi_n_3652 ,csa_tree_add_6_33_groupi_n_4105);
  or csa_tree_add_6_33_groupi_g14029__8428(csa_tree_add_6_33_groupi_n_4265 ,csa_tree_add_6_33_groupi_n_3677 ,csa_tree_add_6_33_groupi_n_4056);
  or csa_tree_add_6_33_groupi_g14030__5526(csa_tree_add_6_33_groupi_n_4264 ,csa_tree_add_6_33_groupi_n_4126 ,csa_tree_add_6_33_groupi_n_4110);
  or csa_tree_add_6_33_groupi_g14031__6783(csa_tree_add_6_33_groupi_n_4263 ,csa_tree_add_6_33_groupi_n_3972 ,csa_tree_add_6_33_groupi_n_4097);
  or csa_tree_add_6_33_groupi_g14032__3680(csa_tree_add_6_33_groupi_n_4262 ,csa_tree_add_6_33_groupi_n_3657 ,csa_tree_add_6_33_groupi_n_4083);
  and csa_tree_add_6_33_groupi_g14033__1617(csa_tree_add_6_33_groupi_n_4261 ,csa_tree_add_6_33_groupi_n_3657 ,csa_tree_add_6_33_groupi_n_4083);
  nor csa_tree_add_6_33_groupi_g14034__2802(csa_tree_add_6_33_groupi_n_4260 ,csa_tree_add_6_33_groupi_n_4014 ,csa_tree_add_6_33_groupi_n_4087);
  nor csa_tree_add_6_33_groupi_g14035__1705(csa_tree_add_6_33_groupi_n_4259 ,csa_tree_add_6_33_groupi_n_3971 ,csa_tree_add_6_33_groupi_n_4098);
  or csa_tree_add_6_33_groupi_g14036__5122(csa_tree_add_6_33_groupi_n_4258 ,csa_tree_add_6_33_groupi_n_4015 ,csa_tree_add_6_33_groupi_n_4086);
  and csa_tree_add_6_33_groupi_g14037__8246(csa_tree_add_6_33_groupi_n_4257 ,csa_tree_add_6_33_groupi_n_3536 ,csa_tree_add_6_33_groupi_n_4103);
  or csa_tree_add_6_33_groupi_g14038__7098(csa_tree_add_6_33_groupi_n_4256 ,csa_tree_add_6_33_groupi_n_3606 ,csa_tree_add_6_33_groupi_n_4079);
  and csa_tree_add_6_33_groupi_g14039__6131(csa_tree_add_6_33_groupi_n_4255 ,csa_tree_add_6_33_groupi_n_3606 ,csa_tree_add_6_33_groupi_n_4079);
  or csa_tree_add_6_33_groupi_g14040__1881(csa_tree_add_6_33_groupi_n_4254 ,csa_tree_add_6_33_groupi_n_3630 ,csa_tree_add_6_33_groupi_n_4081);
  or csa_tree_add_6_33_groupi_g14041__5115(csa_tree_add_6_33_groupi_n_4253 ,csa_tree_add_6_33_groupi_n_3969 ,csa_tree_add_6_33_groupi_n_4082);
  and csa_tree_add_6_33_groupi_g14042__7482(csa_tree_add_6_33_groupi_n_4252 ,csa_tree_add_6_33_groupi_n_4011 ,csa_tree_add_6_33_groupi_n_4076);
  and csa_tree_add_6_33_groupi_g14043__4733(csa_tree_add_6_33_groupi_n_4251 ,csa_tree_add_6_33_groupi_n_3969 ,csa_tree_add_6_33_groupi_n_4082);
  nor csa_tree_add_6_33_groupi_g14044__6161(csa_tree_add_6_33_groupi_n_4250 ,csa_tree_add_6_33_groupi_n_3631 ,csa_tree_add_6_33_groupi_n_4080);
  or csa_tree_add_6_33_groupi_g14045__9315(csa_tree_add_6_33_groupi_n_4249 ,csa_tree_add_6_33_groupi_n_3919 ,csa_tree_add_6_33_groupi_n_4115);
  or csa_tree_add_6_33_groupi_g14046__9945(csa_tree_add_6_33_groupi_n_4248 ,csa_tree_add_6_33_groupi_n_3977 ,csa_tree_add_6_33_groupi_n_4078);
  nor csa_tree_add_6_33_groupi_g14047__2883(csa_tree_add_6_33_groupi_n_4247 ,csa_tree_add_6_33_groupi_n_3978 ,csa_tree_add_6_33_groupi_n_4077);
  or csa_tree_add_6_33_groupi_g14048__2346(csa_tree_add_6_33_groupi_n_4246 ,csa_tree_add_6_33_groupi_n_4011 ,csa_tree_add_6_33_groupi_n_4076);
  or csa_tree_add_6_33_groupi_g14049__1666(csa_tree_add_6_33_groupi_n_4245 ,csa_tree_add_6_33_groupi_n_4009 ,csa_tree_add_6_33_groupi_n_4073);
  or csa_tree_add_6_33_groupi_g14050__7410(csa_tree_add_6_33_groupi_n_4244 ,csa_tree_add_6_33_groupi_n_3915 ,csa_tree_add_6_33_groupi_n_4120);
  or csa_tree_add_6_33_groupi_g14051__6417(csa_tree_add_6_33_groupi_n_4243 ,csa_tree_add_6_33_groupi_n_4144 ,csa_tree_add_6_33_groupi_n_4067);
  or csa_tree_add_6_33_groupi_g14052__5477(csa_tree_add_6_33_groupi_n_4242 ,csa_tree_add_6_33_groupi_n_3975 ,csa_tree_add_6_33_groupi_n_4094);
  or csa_tree_add_6_33_groupi_g14053__2398(csa_tree_add_6_33_groupi_n_4241 ,csa_tree_add_6_33_groupi_n_3772 ,csa_tree_add_6_33_groupi_n_4130);
  nor csa_tree_add_6_33_groupi_g14054__5107(csa_tree_add_6_33_groupi_n_4240 ,csa_tree_add_6_33_groupi_n_3976 ,csa_tree_add_6_33_groupi_n_4095);
  or csa_tree_add_6_33_groupi_g14055__6260(csa_tree_add_6_33_groupi_n_4239 ,csa_tree_add_6_33_groupi_n_3967 ,csa_tree_add_6_33_groupi_n_4101);
  and csa_tree_add_6_33_groupi_g14056__4319(csa_tree_add_6_33_groupi_n_4238 ,csa_tree_add_6_33_groupi_n_4009 ,csa_tree_add_6_33_groupi_n_4073);
  or csa_tree_add_6_33_groupi_g14057__8428(csa_tree_add_6_33_groupi_n_4237 ,csa_tree_add_6_33_groupi_n_3847 ,csa_tree_add_6_33_groupi_n_4132);
  nor csa_tree_add_6_33_groupi_g14058__5526(csa_tree_add_6_33_groupi_n_4236 ,csa_tree_add_6_33_groupi_n_3966 ,csa_tree_add_6_33_groupi_n_4102);
  and csa_tree_add_6_33_groupi_g14059__6783(csa_tree_add_6_33_groupi_n_4291 ,csa_tree_add_6_33_groupi_n_3868 ,csa_tree_add_6_33_groupi_n_4118);
  and csa_tree_add_6_33_groupi_g14060__3680(csa_tree_add_6_33_groupi_n_4290 ,csa_tree_add_6_33_groupi_n_3719 ,csa_tree_add_6_33_groupi_n_4113);
  and csa_tree_add_6_33_groupi_g14061__1617(csa_tree_add_6_33_groupi_n_4289 ,csa_tree_add_6_33_groupi_n_3827 ,csa_tree_add_6_33_groupi_n_4139);
  or csa_tree_add_6_33_groupi_g14062__2802(csa_tree_add_6_33_groupi_n_4288 ,csa_tree_add_6_33_groupi_n_3493 ,csa_tree_add_6_33_groupi_n_4119);
  and csa_tree_add_6_33_groupi_g14063__1705(csa_tree_add_6_33_groupi_n_4287 ,csa_tree_add_6_33_groupi_n_3898 ,csa_tree_add_6_33_groupi_n_4137);
  and csa_tree_add_6_33_groupi_g14064__5122(csa_tree_add_6_33_groupi_n_4286 ,csa_tree_add_6_33_groupi_n_3908 ,csa_tree_add_6_33_groupi_n_4141);
  and csa_tree_add_6_33_groupi_g14065__8246(csa_tree_add_6_33_groupi_n_4285 ,csa_tree_add_6_33_groupi_n_3988 ,csa_tree_add_6_33_groupi_n_4114);
  and csa_tree_add_6_33_groupi_g14066__7098(csa_tree_add_6_33_groupi_n_4284 ,csa_tree_add_6_33_groupi_n_3990 ,csa_tree_add_6_33_groupi_n_4127);
  not csa_tree_add_6_33_groupi_g14067(csa_tree_add_6_33_groupi_n_4234 ,csa_tree_add_6_33_groupi_n_4233);
  not csa_tree_add_6_33_groupi_g14068(csa_tree_add_6_33_groupi_n_4231 ,csa_tree_add_6_33_groupi_n_4232);
  not csa_tree_add_6_33_groupi_g14069(csa_tree_add_6_33_groupi_n_4230 ,csa_tree_add_6_33_groupi_n_4229);
  not csa_tree_add_6_33_groupi_g14070(csa_tree_add_6_33_groupi_n_4228 ,csa_tree_add_6_33_groupi_n_4227);
  not csa_tree_add_6_33_groupi_g14071(csa_tree_add_6_33_groupi_n_4226 ,csa_tree_add_6_33_groupi_n_4225);
  not csa_tree_add_6_33_groupi_g14072(csa_tree_add_6_33_groupi_n_4223 ,csa_tree_add_6_33_groupi_n_4222);
  not csa_tree_add_6_33_groupi_g14073(csa_tree_add_6_33_groupi_n_4220 ,csa_tree_add_6_33_groupi_n_4221);
  not csa_tree_add_6_33_groupi_g14074(csa_tree_add_6_33_groupi_n_4212 ,csa_tree_add_6_33_groupi_n_4213);
  not csa_tree_add_6_33_groupi_g14075(csa_tree_add_6_33_groupi_n_4209 ,csa_tree_add_6_33_groupi_n_4210);
  not csa_tree_add_6_33_groupi_g14076(csa_tree_add_6_33_groupi_n_4206 ,csa_tree_add_6_33_groupi_n_4207);
  nor csa_tree_add_6_33_groupi_g14077__6131(csa_tree_add_6_33_groupi_n_4200 ,csa_tree_add_6_33_groupi_n_3979 ,csa_tree_add_6_33_groupi_n_4091);
  or csa_tree_add_6_33_groupi_g14078__1881(csa_tree_add_6_33_groupi_n_4199 ,csa_tree_add_6_33_groupi_n_3983 ,csa_tree_add_6_33_groupi_n_4143);
  and csa_tree_add_6_33_groupi_g14079__5115(csa_tree_add_6_33_groupi_n_4198 ,csa_tree_add_6_33_groupi_n_4117 ,csa_tree_add_6_33_groupi_n_4109);
  or csa_tree_add_6_33_groupi_g14080__7482(csa_tree_add_6_33_groupi_n_4197 ,csa_tree_add_6_33_groupi_n_3524 ,csa_tree_add_6_33_groupi_n_4099);
  nor csa_tree_add_6_33_groupi_g14081__4733(csa_tree_add_6_33_groupi_n_4196 ,csa_tree_add_6_33_groupi_n_3525 ,csa_tree_add_6_33_groupi_n_4100);
  or csa_tree_add_6_33_groupi_g14082__6161(csa_tree_add_6_33_groupi_n_4195 ,csa_tree_add_6_33_groupi_n_4018 ,csa_tree_add_6_33_groupi_n_4092);
  nor csa_tree_add_6_33_groupi_g14083__9315(csa_tree_add_6_33_groupi_n_4194 ,csa_tree_add_6_33_groupi_n_4019 ,csa_tree_add_6_33_groupi_n_4093);
  or csa_tree_add_6_33_groupi_g14084__9945(csa_tree_add_6_33_groupi_n_4193 ,csa_tree_add_6_33_groupi_n_4064 ,csa_tree_add_6_33_groupi_n_4111);
  or csa_tree_add_6_33_groupi_g14085__2883(csa_tree_add_6_33_groupi_n_4192 ,csa_tree_add_6_33_groupi_n_1007 ,csa_tree_add_6_33_groupi_n_4090);
  xnor csa_tree_add_6_33_groupi_g14086__2346(out1[5] ,csa_tree_add_6_33_groupi_n_4039 ,csa_tree_add_6_33_groupi_n_3579);
  xnor csa_tree_add_6_33_groupi_g14087__1666(csa_tree_add_6_33_groupi_n_4190 ,csa_tree_add_6_33_groupi_n_4017 ,csa_tree_add_6_33_groupi_n_3845);
  xnor csa_tree_add_6_33_groupi_g14088__7410(csa_tree_add_6_33_groupi_n_4189 ,csa_tree_add_6_33_groupi_n_3668 ,csa_tree_add_6_33_groupi_n_4025);
  xnor csa_tree_add_6_33_groupi_g14089__6417(csa_tree_add_6_33_groupi_n_4188 ,csa_tree_add_6_33_groupi_n_3961 ,csa_tree_add_6_33_groupi_n_3764);
  xnor csa_tree_add_6_33_groupi_g14090__5477(csa_tree_add_6_33_groupi_n_4187 ,csa_tree_add_6_33_groupi_n_3956 ,csa_tree_add_6_33_groupi_n_4030);
  xnor csa_tree_add_6_33_groupi_g14091__2398(csa_tree_add_6_33_groupi_n_4186 ,csa_tree_add_6_33_groupi_n_3655 ,csa_tree_add_6_33_groupi_n_4031);
  xor csa_tree_add_6_33_groupi_g14092__5107(csa_tree_add_6_33_groupi_n_4185 ,csa_tree_add_6_33_groupi_n_4038 ,csa_tree_add_6_33_groupi_n_3657);
  xnor csa_tree_add_6_33_groupi_g14093__6260(csa_tree_add_6_33_groupi_n_4184 ,csa_tree_add_6_33_groupi_n_3671 ,csa_tree_add_6_33_groupi_n_4023);
  xor csa_tree_add_6_33_groupi_g14094__4319(csa_tree_add_6_33_groupi_n_4183 ,csa_tree_add_6_33_groupi_n_4029 ,csa_tree_add_6_33_groupi_n_3606);
  xnor csa_tree_add_6_33_groupi_g14095__8428(csa_tree_add_6_33_groupi_n_4182 ,csa_tree_add_6_33_groupi_n_3912 ,csa_tree_add_6_33_groupi_n_3974);
  xnor csa_tree_add_6_33_groupi_g14096__5526(csa_tree_add_6_33_groupi_n_4181 ,csa_tree_add_6_33_groupi_n_3968 ,csa_tree_add_6_33_groupi_n_3973);
  xnor csa_tree_add_6_33_groupi_g14097__6783(csa_tree_add_6_33_groupi_n_4180 ,csa_tree_add_6_33_groupi_n_3911 ,csa_tree_add_6_33_groupi_n_3970);
  xnor csa_tree_add_6_33_groupi_g14098__3680(csa_tree_add_6_33_groupi_n_4179 ,csa_tree_add_6_33_groupi_n_3651 ,csa_tree_add_6_33_groupi_n_3958);
  xnor csa_tree_add_6_33_groupi_g14099__1617(csa_tree_add_6_33_groupi_n_4178 ,csa_tree_add_6_33_groupi_n_4037 ,csa_tree_add_6_33_groupi_n_4019);
  xor csa_tree_add_6_33_groupi_g14100__2802(csa_tree_add_6_33_groupi_n_4177 ,csa_tree_add_6_33_groupi_n_3969 ,csa_tree_add_6_33_groupi_n_4042);
  xnor csa_tree_add_6_33_groupi_g14102__1705(csa_tree_add_6_33_groupi_n_4176 ,csa_tree_add_6_33_groupi_n_4034 ,csa_tree_add_6_33_groupi_n_3624);
  xnor csa_tree_add_6_33_groupi_g14103__5122(csa_tree_add_6_33_groupi_n_4175 ,csa_tree_add_6_33_groupi_n_3959 ,csa_tree_add_6_33_groupi_n_3477);
  xnor csa_tree_add_6_33_groupi_g14104__8246(csa_tree_add_6_33_groupi_n_4174 ,csa_tree_add_6_33_groupi_n_4008 ,csa_tree_add_6_33_groupi_n_3761);
  xnor csa_tree_add_6_33_groupi_g14105__7098(csa_tree_add_6_33_groupi_n_4173 ,csa_tree_add_6_33_groupi_n_3980 ,csa_tree_add_6_33_groupi_n_3762);
  xnor csa_tree_add_6_33_groupi_g14106__6131(csa_tree_add_6_33_groupi_n_4172 ,csa_tree_add_6_33_groupi_n_4033 ,csa_tree_add_6_33_groupi_n_3652);
  xnor csa_tree_add_6_33_groupi_g14107__1881(csa_tree_add_6_33_groupi_n_4171 ,csa_tree_add_6_33_groupi_n_3972 ,csa_tree_add_6_33_groupi_n_4036);
  xnor csa_tree_add_6_33_groupi_g14108__5115(csa_tree_add_6_33_groupi_n_4235 ,csa_tree_add_6_33_groupi_n_3916 ,csa_tree_add_6_33_groupi_n_3931);
  xnor csa_tree_add_6_33_groupi_g14109__7482(csa_tree_add_6_33_groupi_n_4233 ,csa_tree_add_6_33_groupi_n_3566 ,csa_tree_add_6_33_groupi_n_3943);
  xnor csa_tree_add_6_33_groupi_g14110__4733(csa_tree_add_6_33_groupi_n_4232 ,csa_tree_add_6_33_groupi_n_3678 ,csa_tree_add_6_33_groupi_n_3921);
  xnor csa_tree_add_6_33_groupi_g14111__6161(csa_tree_add_6_33_groupi_n_4229 ,csa_tree_add_6_33_groupi_n_4041 ,csa_tree_add_6_33_groupi_n_3941);
  xnor csa_tree_add_6_33_groupi_g14112__9315(csa_tree_add_6_33_groupi_n_4227 ,csa_tree_add_6_33_groupi_n_3917 ,csa_tree_add_6_33_groupi_n_3940);
  xnor csa_tree_add_6_33_groupi_g14113__9945(csa_tree_add_6_33_groupi_n_4225 ,csa_tree_add_6_33_groupi_n_3680 ,csa_tree_add_6_33_groupi_n_3936);
  xnor csa_tree_add_6_33_groupi_g14114__2883(csa_tree_add_6_33_groupi_n_4224 ,csa_tree_add_6_33_groupi_n_3981 ,csa_tree_add_6_33_groupi_n_3945);
  xnor csa_tree_add_6_33_groupi_g14115__2346(csa_tree_add_6_33_groupi_n_4222 ,csa_tree_add_6_33_groupi_n_4027 ,csa_tree_add_6_33_groupi_n_3932);
  xnor csa_tree_add_6_33_groupi_g14116__1666(csa_tree_add_6_33_groupi_n_4221 ,csa_tree_add_6_33_groupi_n_3765 ,csa_tree_add_6_33_groupi_n_3933);
  xnor csa_tree_add_6_33_groupi_g14117__7410(csa_tree_add_6_33_groupi_n_4219 ,csa_tree_add_6_33_groupi_n_3636 ,csa_tree_add_6_33_groupi_n_3935);
  xnor csa_tree_add_6_33_groupi_g14118__6417(csa_tree_add_6_33_groupi_n_4218 ,csa_tree_add_6_33_groupi_n_4032 ,csa_tree_add_6_33_groupi_n_3922);
  xnor csa_tree_add_6_33_groupi_g14119__5477(csa_tree_add_6_33_groupi_n_4217 ,csa_tree_add_6_33_groupi_n_3954 ,csa_tree_add_6_33_groupi_n_3939);
  xnor csa_tree_add_6_33_groupi_g14120__2398(csa_tree_add_6_33_groupi_n_4216 ,csa_tree_add_6_33_groupi_n_3561 ,csa_tree_add_6_33_groupi_n_3938);
  xnor csa_tree_add_6_33_groupi_g14121__5107(csa_tree_add_6_33_groupi_n_4215 ,csa_tree_add_6_33_groupi_n_3679 ,csa_tree_add_6_33_groupi_n_3930);
  xnor csa_tree_add_6_33_groupi_g14122__6260(csa_tree_add_6_33_groupi_n_4214 ,csa_tree_add_6_33_groupi_n_3760 ,csa_tree_add_6_33_groupi_n_3937);
  xnor csa_tree_add_6_33_groupi_g14123__4319(csa_tree_add_6_33_groupi_n_4213 ,csa_tree_add_6_33_groupi_n_3647 ,csa_tree_add_6_33_groupi_n_3934);
  xnor csa_tree_add_6_33_groupi_g14124__8428(csa_tree_add_6_33_groupi_n_4211 ,csa_tree_add_6_33_groupi_n_3767 ,csa_tree_add_6_33_groupi_n_3928);
  xnor csa_tree_add_6_33_groupi_g14125__5526(csa_tree_add_6_33_groupi_n_4210 ,csa_tree_add_6_33_groupi_n_4040 ,csa_tree_add_6_33_groupi_n_3942);
  xnor csa_tree_add_6_33_groupi_g14126__6783(csa_tree_add_6_33_groupi_n_4208 ,csa_tree_add_6_33_groupi_n_3768 ,csa_tree_add_6_33_groupi_n_3927);
  xnor csa_tree_add_6_33_groupi_g14127__3680(csa_tree_add_6_33_groupi_n_4207 ,csa_tree_add_6_33_groupi_n_3769 ,csa_tree_add_6_33_groupi_n_3944);
  xnor csa_tree_add_6_33_groupi_g14128__1617(csa_tree_add_6_33_groupi_n_4205 ,csa_tree_add_6_33_groupi_n_3675 ,csa_tree_add_6_33_groupi_n_3925);
  xnor csa_tree_add_6_33_groupi_g14129__2802(csa_tree_add_6_33_groupi_n_4204 ,csa_tree_add_6_33_groupi_n_3914 ,csa_tree_add_6_33_groupi_n_3924);
  xnor csa_tree_add_6_33_groupi_g14130__1705(csa_tree_add_6_33_groupi_n_4203 ,csa_tree_add_6_33_groupi_n_4043 ,csa_tree_add_6_33_groupi_n_3777);
  xnor csa_tree_add_6_33_groupi_g14131__5122(csa_tree_add_6_33_groupi_n_4202 ,csa_tree_add_6_33_groupi_n_4021 ,csa_tree_add_6_33_groupi_n_3923);
  and csa_tree_add_6_33_groupi_g14132__8246(csa_tree_add_6_33_groupi_n_4201 ,csa_tree_add_6_33_groupi_n_3949 ,csa_tree_add_6_33_groupi_n_4058);
  not csa_tree_add_6_33_groupi_g14133(csa_tree_add_6_33_groupi_n_4170 ,csa_tree_add_6_33_groupi_n_4169);
  not csa_tree_add_6_33_groupi_g14134(csa_tree_add_6_33_groupi_n_4162 ,csa_tree_add_6_33_groupi_n_4163);
  not csa_tree_add_6_33_groupi_g14135(csa_tree_add_6_33_groupi_n_4159 ,csa_tree_add_6_33_groupi_n_4160);
  not csa_tree_add_6_33_groupi_g14136(csa_tree_add_6_33_groupi_n_4156 ,csa_tree_add_6_33_groupi_n_4157);
  not csa_tree_add_6_33_groupi_g14137(csa_tree_add_6_33_groupi_n_4152 ,csa_tree_add_6_33_groupi_n_4153);
  not csa_tree_add_6_33_groupi_g14138(csa_tree_add_6_33_groupi_n_4149 ,csa_tree_add_6_33_groupi_n_4150);
  not csa_tree_add_6_33_groupi_g14139(csa_tree_add_6_33_groupi_n_4146 ,csa_tree_add_6_33_groupi_n_4147);
  and csa_tree_add_6_33_groupi_g14140__7098(csa_tree_add_6_33_groupi_n_4143 ,csa_tree_add_6_33_groupi_n_3477 ,csa_tree_add_6_33_groupi_n_3959);
  and csa_tree_add_6_33_groupi_g14141__6131(csa_tree_add_6_33_groupi_n_4142 ,csa_tree_add_6_33_groupi_n_3624 ,csa_tree_add_6_33_groupi_n_3962);
  or csa_tree_add_6_33_groupi_g14142__1881(csa_tree_add_6_33_groupi_n_4141 ,csa_tree_add_6_33_groupi_n_3906 ,csa_tree_add_6_33_groupi_n_4041);
  or csa_tree_add_6_33_groupi_g14143__5115(csa_tree_add_6_33_groupi_n_4140 ,csa_tree_add_6_33_groupi_n_3764 ,csa_tree_add_6_33_groupi_n_3961);
  or csa_tree_add_6_33_groupi_g14144__7482(csa_tree_add_6_33_groupi_n_4139 ,csa_tree_add_6_33_groupi_n_3820 ,csa_tree_add_6_33_groupi_n_4032);
  or csa_tree_add_6_33_groupi_g14145__4733(csa_tree_add_6_33_groupi_n_4138 ,csa_tree_add_6_33_groupi_n_3762 ,csa_tree_add_6_33_groupi_n_3980);
  or csa_tree_add_6_33_groupi_g14146__6161(csa_tree_add_6_33_groupi_n_4137 ,csa_tree_add_6_33_groupi_n_3897 ,csa_tree_add_6_33_groupi_n_3981);
  nor csa_tree_add_6_33_groupi_g14147__9315(csa_tree_add_6_33_groupi_n_4136 ,csa_tree_add_6_33_groupi_n_3609 ,csa_tree_add_6_33_groupi_n_4027);
  or csa_tree_add_6_33_groupi_g14148__9945(csa_tree_add_6_33_groupi_n_4135 ,csa_tree_add_6_33_groupi_n_3624 ,csa_tree_add_6_33_groupi_n_3962);
  nor csa_tree_add_6_33_groupi_g14149__2883(csa_tree_add_6_33_groupi_n_4134 ,csa_tree_add_6_33_groupi_n_3651 ,csa_tree_add_6_33_groupi_n_3957);
  and csa_tree_add_6_33_groupi_g14150__2346(csa_tree_add_6_33_groupi_n_4133 ,csa_tree_add_6_33_groupi_n_3762 ,csa_tree_add_6_33_groupi_n_3980);
  nor csa_tree_add_6_33_groupi_g14151__1666(csa_tree_add_6_33_groupi_n_4132 ,csa_tree_add_6_33_groupi_n_3668 ,csa_tree_add_6_33_groupi_n_4024);
  or csa_tree_add_6_33_groupi_g14152__7410(csa_tree_add_6_33_groupi_n_4131 ,csa_tree_add_6_33_groupi_n_3965 ,csa_tree_add_6_33_groupi_n_4020);
  and csa_tree_add_6_33_groupi_g14153__6417(csa_tree_add_6_33_groupi_n_4130 ,csa_tree_add_6_33_groupi_n_3627 ,csa_tree_add_6_33_groupi_n_4021);
  and csa_tree_add_6_33_groupi_g14154__5477(csa_tree_add_6_33_groupi_n_4129 ,csa_tree_add_6_33_groupi_n_3965 ,csa_tree_add_6_33_groupi_n_4020);
  or csa_tree_add_6_33_groupi_g14155__2398(csa_tree_add_6_33_groupi_n_4128 ,csa_tree_add_6_33_groupi_n_3761 ,csa_tree_add_6_33_groupi_n_4008);
  or csa_tree_add_6_33_groupi_g14156__5107(csa_tree_add_6_33_groupi_n_4127 ,csa_tree_add_6_33_groupi_n_3846 ,csa_tree_add_6_33_groupi_n_3952);
  and csa_tree_add_6_33_groupi_g14157__6260(csa_tree_add_6_33_groupi_n_4126 ,csa_tree_add_6_33_groupi_n_3761 ,csa_tree_add_6_33_groupi_n_4008);
  or csa_tree_add_6_33_groupi_g14158__4319(csa_tree_add_6_33_groupi_n_4125 ,csa_tree_add_6_33_groupi_n_3627 ,csa_tree_add_6_33_groupi_n_4021);
  or csa_tree_add_6_33_groupi_g14159__8428(csa_tree_add_6_33_groupi_n_4124 ,csa_tree_add_6_33_groupi_n_3667 ,csa_tree_add_6_33_groupi_n_4025);
  nor csa_tree_add_6_33_groupi_g14160__5526(csa_tree_add_6_33_groupi_n_4123 ,csa_tree_add_6_33_groupi_n_4017 ,csa_tree_add_6_33_groupi_n_3845);
  nor csa_tree_add_6_33_groupi_g14161__6783(csa_tree_add_6_33_groupi_n_4122 ,csa_tree_add_6_33_groupi_n_3670 ,csa_tree_add_6_33_groupi_n_4023);
  or csa_tree_add_6_33_groupi_g14162__3680(csa_tree_add_6_33_groupi_n_4121 ,csa_tree_add_6_33_groupi_n_4016 ,csa_tree_add_6_33_groupi_n_3844);
  and csa_tree_add_6_33_groupi_g14163__1617(csa_tree_add_6_33_groupi_n_4120 ,csa_tree_add_6_33_groupi_n_3632 ,csa_tree_add_6_33_groupi_n_4010);
  and csa_tree_add_6_33_groupi_g14164__2802(csa_tree_add_6_33_groupi_n_4119 ,csa_tree_add_6_33_groupi_n_3488 ,csa_tree_add_6_33_groupi_n_4039);
  or csa_tree_add_6_33_groupi_g14165__1705(csa_tree_add_6_33_groupi_n_4118 ,csa_tree_add_6_33_groupi_n_3891 ,csa_tree_add_6_33_groupi_n_4040);
  or csa_tree_add_6_33_groupi_g14166__5122(csa_tree_add_6_33_groupi_n_4117 ,csa_tree_add_6_33_groupi_n_3671 ,csa_tree_add_6_33_groupi_n_4022);
  or csa_tree_add_6_33_groupi_g14167__8246(csa_tree_add_6_33_groupi_n_4116 ,csa_tree_add_6_33_groupi_n_3632 ,csa_tree_add_6_33_groupi_n_4010);
  and csa_tree_add_6_33_groupi_g14168__7098(csa_tree_add_6_33_groupi_n_4115 ,csa_tree_add_6_33_groupi_n_3635 ,csa_tree_add_6_33_groupi_n_4012);
  or csa_tree_add_6_33_groupi_g14169__6131(csa_tree_add_6_33_groupi_n_4114 ,csa_tree_add_6_33_groupi_n_3918 ,csa_tree_add_6_33_groupi_n_3989);
  or csa_tree_add_6_33_groupi_g14170__1881(csa_tree_add_6_33_groupi_n_4113 ,csa_tree_add_6_33_groupi_n_3710 ,csa_tree_add_6_33_groupi_n_4043);
  or csa_tree_add_6_33_groupi_g14171__5115(csa_tree_add_6_33_groupi_n_4112 ,csa_tree_add_6_33_groupi_n_3635 ,csa_tree_add_6_33_groupi_n_4012);
  or csa_tree_add_6_33_groupi_g14172__7482(csa_tree_add_6_33_groupi_n_4169 ,csa_tree_add_6_33_groupi_n_3835 ,csa_tree_add_6_33_groupi_n_3991);
  and csa_tree_add_6_33_groupi_g14173__4733(csa_tree_add_6_33_groupi_n_4168 ,csa_tree_add_6_33_groupi_n_3880 ,csa_tree_add_6_33_groupi_n_3997);
  and csa_tree_add_6_33_groupi_g14174__6161(csa_tree_add_6_33_groupi_n_4167 ,csa_tree_add_6_33_groupi_n_3893 ,csa_tree_add_6_33_groupi_n_4002);
  and csa_tree_add_6_33_groupi_g14175__9315(csa_tree_add_6_33_groupi_n_4166 ,csa_tree_add_6_33_groupi_n_3822 ,csa_tree_add_6_33_groupi_n_3999);
  or csa_tree_add_6_33_groupi_g14176__9945(csa_tree_add_6_33_groupi_n_4165 ,csa_tree_add_6_33_groupi_n_3902 ,csa_tree_add_6_33_groupi_n_4004);
  and csa_tree_add_6_33_groupi_g14177__2883(csa_tree_add_6_33_groupi_n_4164 ,csa_tree_add_6_33_groupi_n_3909 ,csa_tree_add_6_33_groupi_n_4006);
  and csa_tree_add_6_33_groupi_g14178__2346(csa_tree_add_6_33_groupi_n_4163 ,csa_tree_add_6_33_groupi_n_3852 ,csa_tree_add_6_33_groupi_n_3987);
  and csa_tree_add_6_33_groupi_g14179__1666(csa_tree_add_6_33_groupi_n_4161 ,csa_tree_add_6_33_groupi_n_3830 ,csa_tree_add_6_33_groupi_n_3992);
  and csa_tree_add_6_33_groupi_g14180__7410(csa_tree_add_6_33_groupi_n_4160 ,csa_tree_add_6_33_groupi_n_3876 ,csa_tree_add_6_33_groupi_n_3993);
  and csa_tree_add_6_33_groupi_g14181__6417(csa_tree_add_6_33_groupi_n_4158 ,csa_tree_add_6_33_groupi_n_3877 ,csa_tree_add_6_33_groupi_n_3994);
  and csa_tree_add_6_33_groupi_g14182__5477(csa_tree_add_6_33_groupi_n_4157 ,csa_tree_add_6_33_groupi_n_3901 ,csa_tree_add_6_33_groupi_n_3984);
  and csa_tree_add_6_33_groupi_g14183__2398(csa_tree_add_6_33_groupi_n_4155 ,csa_tree_add_6_33_groupi_n_3886 ,csa_tree_add_6_33_groupi_n_4000);
  and csa_tree_add_6_33_groupi_g14184__5107(csa_tree_add_6_33_groupi_n_4154 ,csa_tree_add_6_33_groupi_n_3826 ,csa_tree_add_6_33_groupi_n_3995);
  and csa_tree_add_6_33_groupi_g14185__6260(csa_tree_add_6_33_groupi_n_4153 ,csa_tree_add_6_33_groupi_n_3888 ,csa_tree_add_6_33_groupi_n_3996);
  and csa_tree_add_6_33_groupi_g14186__4319(csa_tree_add_6_33_groupi_n_4151 ,csa_tree_add_6_33_groupi_n_3858 ,csa_tree_add_6_33_groupi_n_3985);
  and csa_tree_add_6_33_groupi_g14187__8428(csa_tree_add_6_33_groupi_n_4150 ,csa_tree_add_6_33_groupi_n_3860 ,csa_tree_add_6_33_groupi_n_3986);
  and csa_tree_add_6_33_groupi_g14188__5526(csa_tree_add_6_33_groupi_n_4148 ,csa_tree_add_6_33_groupi_n_3862 ,csa_tree_add_6_33_groupi_n_4007);
  and csa_tree_add_6_33_groupi_g14189__6783(csa_tree_add_6_33_groupi_n_4147 ,csa_tree_add_6_33_groupi_n_3903 ,csa_tree_add_6_33_groupi_n_4005);
  and csa_tree_add_6_33_groupi_g14190__3680(csa_tree_add_6_33_groupi_n_4145 ,csa_tree_add_6_33_groupi_n_3816 ,csa_tree_add_6_33_groupi_n_4001);
  and csa_tree_add_6_33_groupi_g14191__1617(csa_tree_add_6_33_groupi_n_4144 ,csa_tree_add_6_33_groupi_n_3910 ,csa_tree_add_6_33_groupi_n_3998);
  not csa_tree_add_6_33_groupi_g14192(csa_tree_add_6_33_groupi_n_4107 ,csa_tree_add_6_33_groupi_n_4106);
  not csa_tree_add_6_33_groupi_g14193(csa_tree_add_6_33_groupi_n_4101 ,csa_tree_add_6_33_groupi_n_4102);
  not csa_tree_add_6_33_groupi_g14194(csa_tree_add_6_33_groupi_n_4100 ,csa_tree_add_6_33_groupi_n_4099);
  not csa_tree_add_6_33_groupi_g14195(csa_tree_add_6_33_groupi_n_4097 ,csa_tree_add_6_33_groupi_n_4098);
  not csa_tree_add_6_33_groupi_g14196(csa_tree_add_6_33_groupi_n_4095 ,csa_tree_add_6_33_groupi_n_4094);
  not csa_tree_add_6_33_groupi_g14197(csa_tree_add_6_33_groupi_n_4093 ,csa_tree_add_6_33_groupi_n_4092);
  not csa_tree_add_6_33_groupi_g14198(csa_tree_add_6_33_groupi_n_4091 ,csa_tree_add_6_33_groupi_n_4090);
  not csa_tree_add_6_33_groupi_g14199(csa_tree_add_6_33_groupi_n_4088 ,csa_tree_add_6_33_groupi_n_4089);
  not csa_tree_add_6_33_groupi_g14200(csa_tree_add_6_33_groupi_n_4086 ,csa_tree_add_6_33_groupi_n_4087);
  not csa_tree_add_6_33_groupi_g14201(csa_tree_add_6_33_groupi_n_4085 ,csa_tree_add_6_33_groupi_n_4084);
  not csa_tree_add_6_33_groupi_g14202(csa_tree_add_6_33_groupi_n_4080 ,csa_tree_add_6_33_groupi_n_4081);
  not csa_tree_add_6_33_groupi_g14203(csa_tree_add_6_33_groupi_n_4077 ,csa_tree_add_6_33_groupi_n_4078);
  not csa_tree_add_6_33_groupi_g14204(csa_tree_add_6_33_groupi_n_4074 ,csa_tree_add_6_33_groupi_n_4075);
  not csa_tree_add_6_33_groupi_g14205(csa_tree_add_6_33_groupi_n_4071 ,csa_tree_add_6_33_groupi_n_4070);
  not csa_tree_add_6_33_groupi_g14206(csa_tree_add_6_33_groupi_n_4065 ,csa_tree_add_6_33_groupi_n_4066);
  and csa_tree_add_6_33_groupi_g14207__2802(csa_tree_add_6_33_groupi_n_4064 ,csa_tree_add_6_33_groupi_n_3764 ,csa_tree_add_6_33_groupi_n_3961);
  or csa_tree_add_6_33_groupi_g14208__1705(csa_tree_add_6_33_groupi_n_4063 ,csa_tree_add_6_33_groupi_n_3477 ,csa_tree_add_6_33_groupi_n_3959);
  or csa_tree_add_6_33_groupi_g14209__5122(csa_tree_add_6_33_groupi_n_4062 ,csa_tree_add_6_33_groupi_n_3911 ,csa_tree_add_6_33_groupi_n_3970);
  and csa_tree_add_6_33_groupi_g14210__8246(csa_tree_add_6_33_groupi_n_4061 ,csa_tree_add_6_33_groupi_n_3911 ,csa_tree_add_6_33_groupi_n_3970);
  or csa_tree_add_6_33_groupi_g14211__7098(csa_tree_add_6_33_groupi_n_4060 ,csa_tree_add_6_33_groupi_n_3650 ,csa_tree_add_6_33_groupi_n_3958);
  or csa_tree_add_6_33_groupi_g14212__6131(csa_tree_add_6_33_groupi_n_4059 ,csa_tree_add_6_33_groupi_n_3610 ,csa_tree_add_6_33_groupi_n_4026);
  or csa_tree_add_6_33_groupi_g14213__1881(csa_tree_add_6_33_groupi_n_4058 ,csa_tree_add_6_33_groupi_n_3948 ,csa_tree_add_6_33_groupi_n_3982);
  or csa_tree_add_6_33_groupi_g14214__5115(csa_tree_add_6_33_groupi_n_4057 ,csa_tree_add_6_33_groupi_n_3613 ,csa_tree_add_6_33_groupi_n_3953);
  nor csa_tree_add_6_33_groupi_g14215__7482(csa_tree_add_6_33_groupi_n_4056 ,csa_tree_add_6_33_groupi_n_3614 ,csa_tree_add_6_33_groupi_n_3954);
  and csa_tree_add_6_33_groupi_g14216__4733(csa_tree_add_6_33_groupi_n_4055 ,csa_tree_add_6_33_groupi_n_3912 ,csa_tree_add_6_33_groupi_n_3974);
  or csa_tree_add_6_33_groupi_g14217__6161(csa_tree_add_6_33_groupi_n_4054 ,csa_tree_add_6_33_groupi_n_3912 ,csa_tree_add_6_33_groupi_n_3974);
  and csa_tree_add_6_33_groupi_g14218__9315(csa_tree_add_6_33_groupi_n_4053 ,csa_tree_add_6_33_groupi_n_3968 ,csa_tree_add_6_33_groupi_n_3973);
  or csa_tree_add_6_33_groupi_g14219__9945(csa_tree_add_6_33_groupi_n_4052 ,csa_tree_add_6_33_groupi_n_3968 ,csa_tree_add_6_33_groupi_n_3973);
  xor csa_tree_add_6_33_groupi_g14220__2883(csa_tree_add_6_33_groupi_n_4051 ,csa_tree_add_6_33_groupi_n_3919 ,csa_tree_add_6_33_groupi_n_3635);
  xnor csa_tree_add_6_33_groupi_g14221__2346(csa_tree_add_6_33_groupi_n_4050 ,csa_tree_add_6_33_groupi_n_3608 ,csa_tree_add_6_33_groupi_n_3840);
  xnor csa_tree_add_6_33_groupi_g14222__1666(csa_tree_add_6_33_groupi_n_4049 ,csa_tree_add_6_33_groupi_n_3632 ,csa_tree_add_6_33_groupi_n_3915);
  xnor csa_tree_add_6_33_groupi_g14223__7410(csa_tree_add_6_33_groupi_n_4048 ,csa_tree_add_6_33_groupi_n_3843 ,csa_tree_add_6_33_groupi_n_3427);
  xnor csa_tree_add_6_33_groupi_g14224__6417(csa_tree_add_6_33_groupi_n_4047 ,csa_tree_add_6_33_groupi_n_3525 ,csa_tree_add_6_33_groupi_n_3920);
  xnor csa_tree_add_6_33_groupi_g14225__5477(csa_tree_add_6_33_groupi_n_4046 ,csa_tree_add_6_33_groupi_n_3363 ,csa_tree_add_6_33_groupi_n_3841);
  xnor csa_tree_add_6_33_groupi_g14226__2398(csa_tree_add_6_33_groupi_n_4045 ,csa_tree_add_6_33_groupi_n_3369 ,csa_tree_add_6_33_groupi_n_3838);
  xnor csa_tree_add_6_33_groupi_g14227__5107(csa_tree_add_6_33_groupi_n_4111 ,csa_tree_add_6_33_groupi_n_3617 ,csa_tree_add_6_33_groupi_n_3800);
  xnor csa_tree_add_6_33_groupi_g14228__6260(csa_tree_add_6_33_groupi_n_4110 ,csa_tree_add_6_33_groupi_n_3552 ,csa_tree_add_6_33_groupi_n_3786);
  xnor csa_tree_add_6_33_groupi_g14229__4319(csa_tree_add_6_33_groupi_n_4109 ,csa_tree_add_6_33_groupi_n_3443 ,csa_tree_add_6_33_groupi_n_3799);
  and csa_tree_add_6_33_groupi_g14230__8428(csa_tree_add_6_33_groupi_n_4108 ,csa_tree_add_6_33_groupi_n_3813 ,csa_tree_add_6_33_groupi_n_4003);
  xnor csa_tree_add_6_33_groupi_g14231__5526(csa_tree_add_6_33_groupi_n_4106 ,csa_tree_add_6_33_groupi_n_3476 ,csa_tree_add_6_33_groupi_n_3788);
  xnor csa_tree_add_6_33_groupi_g14232__6783(csa_tree_add_6_33_groupi_n_4105 ,csa_tree_add_6_33_groupi_n_3416 ,csa_tree_add_6_33_groupi_n_3802);
  xnor csa_tree_add_6_33_groupi_g14233__3680(csa_tree_add_6_33_groupi_n_4104 ,csa_tree_add_6_33_groupi_n_3463 ,csa_tree_add_6_33_groupi_n_3801);
  xnor csa_tree_add_6_33_groupi_g14234__1617(csa_tree_add_6_33_groupi_n_4103 ,csa_tree_add_6_33_groupi_n_3666 ,csa_tree_add_6_33_groupi_n_3787);
  xnor csa_tree_add_6_33_groupi_g14235__2802(csa_tree_add_6_33_groupi_n_4102 ,csa_tree_add_6_33_groupi_n_3562 ,csa_tree_add_6_33_groupi_n_3805);
  xnor csa_tree_add_6_33_groupi_g14236__1705(csa_tree_add_6_33_groupi_n_4099 ,csa_tree_add_6_33_groupi_n_3468 ,csa_tree_add_6_33_groupi_n_3779);
  xnor csa_tree_add_6_33_groupi_g14237__5122(csa_tree_add_6_33_groupi_n_4098 ,csa_tree_add_6_33_groupi_n_3622 ,csa_tree_add_6_33_groupi_n_3785);
  and csa_tree_add_6_33_groupi_g14238__8246(csa_tree_add_6_33_groupi_n_4096 ,csa_tree_add_6_33_groupi_n_3811 ,csa_tree_add_6_33_groupi_n_3951);
  xnor csa_tree_add_6_33_groupi_g14239__7098(csa_tree_add_6_33_groupi_n_4094 ,csa_tree_add_6_33_groupi_n_3436 ,csa_tree_add_6_33_groupi_n_3796);
  xnor csa_tree_add_6_33_groupi_g14240__6131(csa_tree_add_6_33_groupi_n_4092 ,csa_tree_add_6_33_groupi_n_3373 ,csa_tree_add_6_33_groupi_n_3795);
  xnor csa_tree_add_6_33_groupi_g14241__1881(csa_tree_add_6_33_groupi_n_4090 ,csa_tree_add_6_33_groupi_n_3620 ,csa_tree_add_6_33_groupi_n_3794);
  xnor csa_tree_add_6_33_groupi_g14242__5115(csa_tree_add_6_33_groupi_n_4089 ,csa_tree_add_6_33_groupi_n_3553 ,csa_tree_add_6_33_groupi_n_3773);
  xnor csa_tree_add_6_33_groupi_g14243__7482(csa_tree_add_6_33_groupi_n_4087 ,csa_tree_add_6_33_groupi_n_3681 ,csa_tree_add_6_33_groupi_n_3807);
  xnor csa_tree_add_6_33_groupi_g14244__4733(csa_tree_add_6_33_groupi_n_4084 ,csa_tree_add_6_33_groupi_n_3669 ,csa_tree_add_6_33_groupi_n_3793);
  xnor csa_tree_add_6_33_groupi_g14245__6161(csa_tree_add_6_33_groupi_n_4083 ,csa_tree_add_6_33_groupi_n_3569 ,csa_tree_add_6_33_groupi_n_3784);
  xnor csa_tree_add_6_33_groupi_g14246__9315(csa_tree_add_6_33_groupi_n_4082 ,csa_tree_add_6_33_groupi_n_3642 ,csa_tree_add_6_33_groupi_n_3781);
  xnor csa_tree_add_6_33_groupi_g14247__9945(csa_tree_add_6_33_groupi_n_4081 ,csa_tree_add_6_33_groupi_n_3771 ,csa_tree_add_6_33_groupi_n_3780);
  xnor csa_tree_add_6_33_groupi_g14248__2883(csa_tree_add_6_33_groupi_n_4079 ,csa_tree_add_6_33_groupi_n_3460 ,csa_tree_add_6_33_groupi_n_3783);
  xnor csa_tree_add_6_33_groupi_g14249__2346(csa_tree_add_6_33_groupi_n_4078 ,csa_tree_add_6_33_groupi_n_3674 ,csa_tree_add_6_33_groupi_n_3776);
  xnor csa_tree_add_6_33_groupi_g14250__1666(csa_tree_add_6_33_groupi_n_4076 ,csa_tree_add_6_33_groupi_n_3558 ,csa_tree_add_6_33_groupi_n_3775);
  xnor csa_tree_add_6_33_groupi_g14251__7410(csa_tree_add_6_33_groupi_n_4075 ,csa_tree_add_6_33_groupi_n_3448 ,csa_tree_add_6_33_groupi_n_3789);
  xnor csa_tree_add_6_33_groupi_g14252__6417(csa_tree_add_6_33_groupi_n_4073 ,csa_tree_add_6_33_groupi_n_3431 ,csa_tree_add_6_33_groupi_n_3774);
  xnor csa_tree_add_6_33_groupi_g14253__5477(csa_tree_add_6_33_groupi_n_4072 ,csa_tree_add_6_33_groupi_n_3559 ,csa_tree_add_6_33_groupi_n_3778);
  xnor csa_tree_add_6_33_groupi_g14254__2398(csa_tree_add_6_33_groupi_n_4070 ,csa_tree_add_6_33_groupi_n_3407 ,csa_tree_add_6_33_groupi_n_3791);
  xnor csa_tree_add_6_33_groupi_g14255__5107(csa_tree_add_6_33_groupi_n_4069 ,csa_tree_add_6_33_groupi_n_3424 ,csa_tree_add_6_33_groupi_n_3803);
  xnor csa_tree_add_6_33_groupi_g14256__6260(csa_tree_add_6_33_groupi_n_4068 ,csa_tree_add_6_33_groupi_n_3426 ,csa_tree_add_6_33_groupi_n_3804);
  xnor csa_tree_add_6_33_groupi_g14257__4319(csa_tree_add_6_33_groupi_n_4067 ,csa_tree_add_6_33_groupi_n_3572 ,csa_tree_add_6_33_groupi_n_3790);
  xnor csa_tree_add_6_33_groupi_g14258__8428(csa_tree_add_6_33_groupi_n_4066 ,csa_tree_add_6_33_groupi_n_3465 ,csa_tree_add_6_33_groupi_n_3792);
  not csa_tree_add_6_33_groupi_g14259(csa_tree_add_6_33_groupi_n_4027 ,csa_tree_add_6_33_groupi_n_4026);
  not csa_tree_add_6_33_groupi_g14260(csa_tree_add_6_33_groupi_n_4024 ,csa_tree_add_6_33_groupi_n_4025);
  not csa_tree_add_6_33_groupi_g14261(csa_tree_add_6_33_groupi_n_4022 ,csa_tree_add_6_33_groupi_n_4023);
  not csa_tree_add_6_33_groupi_g14262(csa_tree_add_6_33_groupi_n_4019 ,csa_tree_add_6_33_groupi_n_4018);
  not csa_tree_add_6_33_groupi_g14263(csa_tree_add_6_33_groupi_n_4017 ,csa_tree_add_6_33_groupi_n_4016);
  not csa_tree_add_6_33_groupi_g14264(csa_tree_add_6_33_groupi_n_4014 ,csa_tree_add_6_33_groupi_n_4015);
  or csa_tree_add_6_33_groupi_g14265__5526(csa_tree_add_6_33_groupi_n_4007 ,csa_tree_add_6_33_groupi_n_3675 ,csa_tree_add_6_33_groupi_n_3863);
  or csa_tree_add_6_33_groupi_g14266__6783(csa_tree_add_6_33_groupi_n_4006 ,csa_tree_add_6_33_groupi_n_3549 ,csa_tree_add_6_33_groupi_n_3895);
  or csa_tree_add_6_33_groupi_g14267__3680(csa_tree_add_6_33_groupi_n_4005 ,csa_tree_add_6_33_groupi_n_3679 ,csa_tree_add_6_33_groupi_n_3900);
  and csa_tree_add_6_33_groupi_g14268__1617(csa_tree_add_6_33_groupi_n_4004 ,csa_tree_add_6_33_groupi_n_3917 ,csa_tree_add_6_33_groupi_n_3899);
  or csa_tree_add_6_33_groupi_g14269__2802(csa_tree_add_6_33_groupi_n_4003 ,csa_tree_add_6_33_groupi_n_3483 ,csa_tree_add_6_33_groupi_n_3812);
  or csa_tree_add_6_33_groupi_g14270__1705(csa_tree_add_6_33_groupi_n_4002 ,csa_tree_add_6_33_groupi_n_3916 ,csa_tree_add_6_33_groupi_n_3890);
  or csa_tree_add_6_33_groupi_g14271__5122(csa_tree_add_6_33_groupi_n_4001 ,csa_tree_add_6_33_groupi_n_3481 ,csa_tree_add_6_33_groupi_n_3815);
  or csa_tree_add_6_33_groupi_g14272__8246(csa_tree_add_6_33_groupi_n_4000 ,csa_tree_add_6_33_groupi_n_3678 ,csa_tree_add_6_33_groupi_n_3885);
  or csa_tree_add_6_33_groupi_g14273__7098(csa_tree_add_6_33_groupi_n_3999 ,csa_tree_add_6_33_groupi_n_3547 ,csa_tree_add_6_33_groupi_n_3818);
  or csa_tree_add_6_33_groupi_g14274__6131(csa_tree_add_6_33_groupi_n_3998 ,csa_tree_add_6_33_groupi_n_3765 ,csa_tree_add_6_33_groupi_n_3892);
  or csa_tree_add_6_33_groupi_g14275__1881(csa_tree_add_6_33_groupi_n_3997 ,csa_tree_add_6_33_groupi_n_3560 ,csa_tree_add_6_33_groupi_n_3875);
  or csa_tree_add_6_33_groupi_g14276__5115(csa_tree_add_6_33_groupi_n_3996 ,csa_tree_add_6_33_groupi_n_3914 ,csa_tree_add_6_33_groupi_n_3869);
  or csa_tree_add_6_33_groupi_g14277__7482(csa_tree_add_6_33_groupi_n_3995 ,csa_tree_add_6_33_groupi_n_3566 ,csa_tree_add_6_33_groupi_n_3825);
  or csa_tree_add_6_33_groupi_g14278__4733(csa_tree_add_6_33_groupi_n_3994 ,csa_tree_add_6_33_groupi_n_3561 ,csa_tree_add_6_33_groupi_n_3874);
  or csa_tree_add_6_33_groupi_g14279__6161(csa_tree_add_6_33_groupi_n_3993 ,csa_tree_add_6_33_groupi_n_3767 ,csa_tree_add_6_33_groupi_n_3870);
  or csa_tree_add_6_33_groupi_g14280__9315(csa_tree_add_6_33_groupi_n_3992 ,csa_tree_add_6_33_groupi_n_3831 ,csa_tree_add_6_33_groupi_n_3676);
  and csa_tree_add_6_33_groupi_g14281__9945(csa_tree_add_6_33_groupi_n_3991 ,csa_tree_add_6_33_groupi_n_3680 ,csa_tree_add_6_33_groupi_n_3832);
  or csa_tree_add_6_33_groupi_g14282__2883(csa_tree_add_6_33_groupi_n_3990 ,csa_tree_add_6_33_groupi_n_3427 ,csa_tree_add_6_33_groupi_n_3843);
  nor csa_tree_add_6_33_groupi_g14283__2346(csa_tree_add_6_33_groupi_n_3989 ,csa_tree_add_6_33_groupi_n_3368 ,csa_tree_add_6_33_groupi_n_3838);
  or csa_tree_add_6_33_groupi_g14284__1666(csa_tree_add_6_33_groupi_n_3988 ,csa_tree_add_6_33_groupi_n_3369 ,csa_tree_add_6_33_groupi_n_3837);
  or csa_tree_add_6_33_groupi_g14285__7410(csa_tree_add_6_33_groupi_n_3987 ,csa_tree_add_6_33_groupi_n_3770 ,csa_tree_add_6_33_groupi_n_3850);
  or csa_tree_add_6_33_groupi_g14286__6417(csa_tree_add_6_33_groupi_n_3986 ,csa_tree_add_6_33_groupi_n_3564 ,csa_tree_add_6_33_groupi_n_3904);
  or csa_tree_add_6_33_groupi_g14287__5477(csa_tree_add_6_33_groupi_n_3985 ,csa_tree_add_6_33_groupi_n_3769 ,csa_tree_add_6_33_groupi_n_3859);
  or csa_tree_add_6_33_groupi_g14288__2398(csa_tree_add_6_33_groupi_n_3984 ,csa_tree_add_6_33_groupi_n_3768 ,csa_tree_add_6_33_groupi_n_3857);
  and csa_tree_add_6_33_groupi_g14289__5107(csa_tree_add_6_33_groupi_n_4044 ,csa_tree_add_6_33_groupi_n_3748 ,csa_tree_add_6_33_groupi_n_3894);
  and csa_tree_add_6_33_groupi_g14290__6260(csa_tree_add_6_33_groupi_n_4043 ,csa_tree_add_6_33_groupi_n_3709 ,csa_tree_add_6_33_groupi_n_3851);
  and csa_tree_add_6_33_groupi_g14291__4319(csa_tree_add_6_33_groupi_n_4042 ,csa_tree_add_6_33_groupi_n_3715 ,csa_tree_add_6_33_groupi_n_3854);
  and csa_tree_add_6_33_groupi_g14292__8428(csa_tree_add_6_33_groupi_n_4041 ,csa_tree_add_6_33_groupi_n_3754 ,csa_tree_add_6_33_groupi_n_3905);
  and csa_tree_add_6_33_groupi_g14293__5526(csa_tree_add_6_33_groupi_n_4040 ,csa_tree_add_6_33_groupi_n_3691 ,csa_tree_add_6_33_groupi_n_3834);
  or csa_tree_add_6_33_groupi_g14294__6783(csa_tree_add_6_33_groupi_n_4039 ,csa_tree_add_6_33_groupi_n_3299 ,csa_tree_add_6_33_groupi_n_3861);
  and csa_tree_add_6_33_groupi_g14295__3680(csa_tree_add_6_33_groupi_n_4038 ,csa_tree_add_6_33_groupi_n_3726 ,csa_tree_add_6_33_groupi_n_3867);
  and csa_tree_add_6_33_groupi_g14296__1617(csa_tree_add_6_33_groupi_n_4037 ,csa_tree_add_6_33_groupi_n_3690 ,csa_tree_add_6_33_groupi_n_3828);
  and csa_tree_add_6_33_groupi_g14297__2802(csa_tree_add_6_33_groupi_n_4036 ,csa_tree_add_6_33_groupi_n_3729 ,csa_tree_add_6_33_groupi_n_3865);
  and csa_tree_add_6_33_groupi_g14298__1705(csa_tree_add_6_33_groupi_n_4035 ,csa_tree_add_6_33_groupi_n_3734 ,csa_tree_add_6_33_groupi_n_3873);
  and csa_tree_add_6_33_groupi_g14299__5122(csa_tree_add_6_33_groupi_n_4034 ,csa_tree_add_6_33_groupi_n_3743 ,csa_tree_add_6_33_groupi_n_3819);
  and csa_tree_add_6_33_groupi_g14300__8246(csa_tree_add_6_33_groupi_n_4033 ,csa_tree_add_6_33_groupi_n_3605 ,csa_tree_add_6_33_groupi_n_3881);
  and csa_tree_add_6_33_groupi_g14301__7098(csa_tree_add_6_33_groupi_n_4032 ,csa_tree_add_6_33_groupi_n_3751 ,csa_tree_add_6_33_groupi_n_3817);
  and csa_tree_add_6_33_groupi_g14302__6131(csa_tree_add_6_33_groupi_n_4031 ,csa_tree_add_6_33_groupi_n_3739 ,csa_tree_add_6_33_groupi_n_3883);
  and csa_tree_add_6_33_groupi_g14303__1881(csa_tree_add_6_33_groupi_n_4030 ,csa_tree_add_6_33_groupi_n_3741 ,csa_tree_add_6_33_groupi_n_3884);
  and csa_tree_add_6_33_groupi_g14304__5115(csa_tree_add_6_33_groupi_n_4029 ,csa_tree_add_6_33_groupi_n_3712 ,csa_tree_add_6_33_groupi_n_3856);
  or csa_tree_add_6_33_groupi_g14305__7482(csa_tree_add_6_33_groupi_n_4028 ,csa_tree_add_6_33_groupi_n_3503 ,csa_tree_add_6_33_groupi_n_3872);
  and csa_tree_add_6_33_groupi_g14306__4733(csa_tree_add_6_33_groupi_n_4026 ,csa_tree_add_6_33_groupi_n_3714 ,csa_tree_add_6_33_groupi_n_3907);
  and csa_tree_add_6_33_groupi_g14307__6161(csa_tree_add_6_33_groupi_n_4025 ,csa_tree_add_6_33_groupi_n_3688 ,csa_tree_add_6_33_groupi_n_3833);
  and csa_tree_add_6_33_groupi_g14308__9315(csa_tree_add_6_33_groupi_n_4023 ,csa_tree_add_6_33_groupi_n_3758 ,csa_tree_add_6_33_groupi_n_3866);
  and csa_tree_add_6_33_groupi_g14309__9945(csa_tree_add_6_33_groupi_n_4021 ,csa_tree_add_6_33_groupi_n_3687 ,csa_tree_add_6_33_groupi_n_3829);
  and csa_tree_add_6_33_groupi_g14310__2883(csa_tree_add_6_33_groupi_n_4020 ,csa_tree_add_6_33_groupi_n_3744 ,csa_tree_add_6_33_groupi_n_3887);
  and csa_tree_add_6_33_groupi_g14311__2346(csa_tree_add_6_33_groupi_n_4018 ,csa_tree_add_6_33_groupi_n_3711 ,csa_tree_add_6_33_groupi_n_3824);
  and csa_tree_add_6_33_groupi_g14312__1666(csa_tree_add_6_33_groupi_n_4016 ,csa_tree_add_6_33_groupi_n_3720 ,csa_tree_add_6_33_groupi_n_3855);
  and csa_tree_add_6_33_groupi_g14313__7410(csa_tree_add_6_33_groupi_n_4015 ,csa_tree_add_6_33_groupi_n_3732 ,csa_tree_add_6_33_groupi_n_3823);
  and csa_tree_add_6_33_groupi_g14314__6417(csa_tree_add_6_33_groupi_n_4013 ,csa_tree_add_6_33_groupi_n_3705 ,csa_tree_add_6_33_groupi_n_3849);
  and csa_tree_add_6_33_groupi_g14315__5477(csa_tree_add_6_33_groupi_n_4012 ,csa_tree_add_6_33_groupi_n_3703 ,csa_tree_add_6_33_groupi_n_3853);
  and csa_tree_add_6_33_groupi_g14316__2398(csa_tree_add_6_33_groupi_n_4011 ,csa_tree_add_6_33_groupi_n_3699 ,csa_tree_add_6_33_groupi_n_3871);
  and csa_tree_add_6_33_groupi_g14317__5107(csa_tree_add_6_33_groupi_n_4010 ,csa_tree_add_6_33_groupi_n_3697 ,csa_tree_add_6_33_groupi_n_3878);
  and csa_tree_add_6_33_groupi_g14318__6260(csa_tree_add_6_33_groupi_n_4009 ,csa_tree_add_6_33_groupi_n_3694 ,csa_tree_add_6_33_groupi_n_3896);
  and csa_tree_add_6_33_groupi_g14319__4319(csa_tree_add_6_33_groupi_n_4008 ,csa_tree_add_6_33_groupi_n_3735 ,csa_tree_add_6_33_groupi_n_3879);
  not csa_tree_add_6_33_groupi_g14321(csa_tree_add_6_33_groupi_n_3977 ,csa_tree_add_6_33_groupi_n_3978);
  not csa_tree_add_6_33_groupi_g14322(csa_tree_add_6_33_groupi_n_3975 ,csa_tree_add_6_33_groupi_n_3976);
  not csa_tree_add_6_33_groupi_g14323(csa_tree_add_6_33_groupi_n_3971 ,csa_tree_add_6_33_groupi_n_3972);
  not csa_tree_add_6_33_groupi_g14324(csa_tree_add_6_33_groupi_n_3967 ,csa_tree_add_6_33_groupi_n_3966);
  not csa_tree_add_6_33_groupi_g14325(csa_tree_add_6_33_groupi_n_3963 ,csa_tree_add_6_33_groupi_n_3964);
  not csa_tree_add_6_33_groupi_g14326(csa_tree_add_6_33_groupi_n_3957 ,csa_tree_add_6_33_groupi_n_3958);
  not csa_tree_add_6_33_groupi_g14327(csa_tree_add_6_33_groupi_n_3956 ,csa_tree_add_6_33_groupi_n_3955);
  not csa_tree_add_6_33_groupi_g14328(csa_tree_add_6_33_groupi_n_3954 ,csa_tree_add_6_33_groupi_n_3953);
  and csa_tree_add_6_33_groupi_g14329__8428(csa_tree_add_6_33_groupi_n_3952 ,csa_tree_add_6_33_groupi_n_3427 ,csa_tree_add_6_33_groupi_n_3843);
  or csa_tree_add_6_33_groupi_g14330__5526(csa_tree_add_6_33_groupi_n_3951 ,csa_tree_add_6_33_groupi_n_3487 ,csa_tree_add_6_33_groupi_n_3810);
  xnor csa_tree_add_6_33_groupi_g14331__6783(out1[4] ,csa_tree_add_6_33_groupi_n_3672 ,csa_tree_add_6_33_groupi_n_3397);
  or csa_tree_add_6_33_groupi_g14332__3680(csa_tree_add_6_33_groupi_n_3949 ,csa_tree_add_6_33_groupi_n_3608 ,csa_tree_add_6_33_groupi_n_3839);
  nor csa_tree_add_6_33_groupi_g14333__1617(csa_tree_add_6_33_groupi_n_3948 ,csa_tree_add_6_33_groupi_n_3607 ,csa_tree_add_6_33_groupi_n_3840);
  or csa_tree_add_6_33_groupi_g14334__2802(csa_tree_add_6_33_groupi_n_3947 ,csa_tree_add_6_33_groupi_n_3363 ,csa_tree_add_6_33_groupi_n_3841);
  and csa_tree_add_6_33_groupi_g14335__1705(csa_tree_add_6_33_groupi_n_3946 ,csa_tree_add_6_33_groupi_n_3363 ,csa_tree_add_6_33_groupi_n_3841);
  xnor csa_tree_add_6_33_groupi_g14336__5122(csa_tree_add_6_33_groupi_n_3945 ,csa_tree_add_6_33_groupi_n_3661 ,csa_tree_add_6_33_groupi_n_3459);
  xnor csa_tree_add_6_33_groupi_g14337__8246(csa_tree_add_6_33_groupi_n_3944 ,csa_tree_add_6_33_groupi_n_3639 ,csa_tree_add_6_33_groupi_n_3634);
  xnor csa_tree_add_6_33_groupi_g14338__7098(csa_tree_add_6_33_groupi_n_3943 ,csa_tree_add_6_33_groupi_n_3435 ,csa_tree_add_6_33_groupi_n_3645);
  xnor csa_tree_add_6_33_groupi_g14339__6131(csa_tree_add_6_33_groupi_n_3942 ,csa_tree_add_6_33_groupi_n_3531 ,csa_tree_add_6_33_groupi_n_3660);
  xnor csa_tree_add_6_33_groupi_g14340__1881(csa_tree_add_6_33_groupi_n_3941 ,csa_tree_add_6_33_groupi_n_3523 ,csa_tree_add_6_33_groupi_n_3665);
  xnor csa_tree_add_6_33_groupi_g14341__5115(csa_tree_add_6_33_groupi_n_3940 ,csa_tree_add_6_33_groupi_n_3409 ,csa_tree_add_6_33_groupi_n_3612);
  xnor csa_tree_add_6_33_groupi_g14342__7482(csa_tree_add_6_33_groupi_n_3939 ,csa_tree_add_6_33_groupi_n_3614 ,csa_tree_add_6_33_groupi_n_3677);
  xnor csa_tree_add_6_33_groupi_g14343__4733(csa_tree_add_6_33_groupi_n_3938 ,csa_tree_add_6_33_groupi_n_3663 ,csa_tree_add_6_33_groupi_n_3450);
  xnor csa_tree_add_6_33_groupi_g14344__6161(csa_tree_add_6_33_groupi_n_3937 ,csa_tree_add_6_33_groupi_n_3473 ,csa_tree_add_6_33_groupi_n_3676);
  xnor csa_tree_add_6_33_groupi_g14345__9315(csa_tree_add_6_33_groupi_n_3936 ,csa_tree_add_6_33_groupi_n_3541 ,csa_tree_add_6_33_groupi_n_3629);
  xnor csa_tree_add_6_33_groupi_g14346__9945(csa_tree_add_6_33_groupi_n_3935 ,csa_tree_add_6_33_groupi_n_3637 ,csa_tree_add_6_33_groupi_n_3770);
  xnor csa_tree_add_6_33_groupi_g14347__2883(csa_tree_add_6_33_groupi_n_3934 ,csa_tree_add_6_33_groupi_n_3619 ,csa_tree_add_6_33_groupi_n_3481);
  xnor csa_tree_add_6_33_groupi_g14348__2346(csa_tree_add_6_33_groupi_n_3933 ,csa_tree_add_6_33_groupi_n_3036 ,csa_tree_add_6_33_groupi_n_3626);
  xnor csa_tree_add_6_33_groupi_g14349__1666(csa_tree_add_6_33_groupi_n_3932 ,csa_tree_add_6_33_groupi_n_3610 ,csa_tree_add_6_33_groupi_n_3766);
  xnor csa_tree_add_6_33_groupi_g14350__7410(csa_tree_add_6_33_groupi_n_3931 ,csa_tree_add_6_33_groupi_n_3658 ,csa_tree_add_6_33_groupi_n_3533);
  xnor csa_tree_add_6_33_groupi_g14351__6417(csa_tree_add_6_33_groupi_n_3930 ,csa_tree_add_6_33_groupi_n_3662 ,csa_tree_add_6_33_groupi_n_3535);
  xnor csa_tree_add_6_33_groupi_g14352__5477(csa_tree_add_6_33_groupi_n_3929 ,csa_tree_add_6_33_groupi_n_3653 ,csa_tree_add_6_33_groupi_n_3763);
  xnor csa_tree_add_6_33_groupi_g14353__2398(csa_tree_add_6_33_groupi_n_3928 ,csa_tree_add_6_33_groupi_n_3648 ,csa_tree_add_6_33_groupi_n_3537);
  xnor csa_tree_add_6_33_groupi_g14354__5107(csa_tree_add_6_33_groupi_n_3927 ,csa_tree_add_6_33_groupi_n_3640 ,csa_tree_add_6_33_groupi_n_3444);
  xnor csa_tree_add_6_33_groupi_g14355__6260(csa_tree_add_6_33_groupi_n_3926 ,csa_tree_add_6_33_groupi_n_3649 ,csa_tree_add_6_33_groupi_n_3641);
  xnor csa_tree_add_6_33_groupi_g14356__4319(csa_tree_add_6_33_groupi_n_3925 ,csa_tree_add_6_33_groupi_n_3643 ,csa_tree_add_6_33_groupi_n_3542);
  xnor csa_tree_add_6_33_groupi_g14357__8428(csa_tree_add_6_33_groupi_n_3924 ,csa_tree_add_6_33_groupi_n_3656 ,csa_tree_add_6_33_groupi_n_3055);
  xnor csa_tree_add_6_33_groupi_g14358__5526(csa_tree_add_6_33_groupi_n_3923 ,csa_tree_add_6_33_groupi_n_3627 ,csa_tree_add_6_33_groupi_n_3772);
  xnor csa_tree_add_6_33_groupi_g14359__6783(csa_tree_add_6_33_groupi_n_3922 ,csa_tree_add_6_33_groupi_n_3623 ,csa_tree_add_6_33_groupi_n_3528);
  xnor csa_tree_add_6_33_groupi_g14360__3680(csa_tree_add_6_33_groupi_n_3921 ,csa_tree_add_6_33_groupi_n_3539 ,csa_tree_add_6_33_groupi_n_3616);
  and csa_tree_add_6_33_groupi_g14361__1617(csa_tree_add_6_33_groupi_n_3983 ,csa_tree_add_6_33_groupi_n_3603 ,csa_tree_add_6_33_groupi_n_3809);
  and csa_tree_add_6_33_groupi_g14362__2802(csa_tree_add_6_33_groupi_n_3982 ,csa_tree_add_6_33_groupi_n_3602 ,csa_tree_add_6_33_groupi_n_3808);
  xnor csa_tree_add_6_33_groupi_g14363__1705(csa_tree_add_6_33_groupi_n_3981 ,csa_tree_add_6_33_groupi_n_3551 ,csa_tree_add_6_33_groupi_n_3574);
  xnor csa_tree_add_6_33_groupi_g14364__5122(csa_tree_add_6_33_groupi_n_3980 ,csa_tree_add_6_33_groupi_n_3412 ,csa_tree_add_6_33_groupi_n_3585);
  xnor csa_tree_add_6_33_groupi_g14365__8246(csa_tree_add_6_33_groupi_n_3979 ,csa_tree_add_6_33_groupi_n_3440 ,csa_tree_add_6_33_groupi_n_3593);
  xnor csa_tree_add_6_33_groupi_g14366__7098(csa_tree_add_6_33_groupi_n_3978 ,csa_tree_add_6_33_groupi_n_3570 ,csa_tree_add_6_33_groupi_n_3584);
  xnor csa_tree_add_6_33_groupi_g14367__6131(csa_tree_add_6_33_groupi_n_3976 ,csa_tree_add_6_33_groupi_n_3382 ,csa_tree_add_6_33_groupi_n_3582);
  xnor csa_tree_add_6_33_groupi_g14368__1881(csa_tree_add_6_33_groupi_n_3974 ,csa_tree_add_6_33_groupi_n_3673 ,csa_tree_add_6_33_groupi_n_3580);
  xnor csa_tree_add_6_33_groupi_g14369__5115(csa_tree_add_6_33_groupi_n_3973 ,csa_tree_add_6_33_groupi_n_3485 ,csa_tree_add_6_33_groupi_n_3577);
  xnor csa_tree_add_6_33_groupi_g14370__7482(csa_tree_add_6_33_groupi_n_3972 ,csa_tree_add_6_33_groupi_n_3187 ,csa_tree_add_6_33_groupi_n_3586);
  xnor csa_tree_add_6_33_groupi_g14371__4733(csa_tree_add_6_33_groupi_n_3970 ,csa_tree_add_6_33_groupi_n_3471 ,csa_tree_add_6_33_groupi_n_3578);
  xnor csa_tree_add_6_33_groupi_g14372__6161(csa_tree_add_6_33_groupi_n_3969 ,csa_tree_add_6_33_groupi_n_3526 ,csa_tree_add_6_33_groupi_n_3587);
  or csa_tree_add_6_33_groupi_g14373__9315(csa_tree_add_6_33_groupi_n_3968 ,csa_tree_add_6_33_groupi_n_3727 ,csa_tree_add_6_33_groupi_n_3814);
  xnor csa_tree_add_6_33_groupi_g14374__9945(csa_tree_add_6_33_groupi_n_3966 ,csa_tree_add_6_33_groupi_n_3275 ,csa_tree_add_6_33_groupi_n_3588);
  xnor csa_tree_add_6_33_groupi_g14375__2883(csa_tree_add_6_33_groupi_n_3965 ,csa_tree_add_6_33_groupi_n_3478 ,csa_tree_add_6_33_groupi_n_3573);
  xnor csa_tree_add_6_33_groupi_g14376__2346(csa_tree_add_6_33_groupi_n_3964 ,csa_tree_add_6_33_groupi_n_3438 ,csa_tree_add_6_33_groupi_n_3589);
  xnor csa_tree_add_6_33_groupi_g14377__1666(csa_tree_add_6_33_groupi_n_3962 ,csa_tree_add_6_33_groupi_n_3550 ,csa_tree_add_6_33_groupi_n_3590);
  xnor csa_tree_add_6_33_groupi_g14378__7410(csa_tree_add_6_33_groupi_n_3961 ,csa_tree_add_6_33_groupi_n_3266 ,csa_tree_add_6_33_groupi_n_3592);
  xor csa_tree_add_6_33_groupi_g14379__6417(csa_tree_add_6_33_groupi_n_3960 ,csa_tree_add_6_33_groupi_n_3529 ,csa_tree_add_6_33_groupi_n_3581);
  xnor csa_tree_add_6_33_groupi_g14380__5477(csa_tree_add_6_33_groupi_n_3959 ,csa_tree_add_6_33_groupi_n_3417 ,csa_tree_add_6_33_groupi_n_3591);
  xnor csa_tree_add_6_33_groupi_g14381__2398(csa_tree_add_6_33_groupi_n_3958 ,csa_tree_add_6_33_groupi_n_3548 ,csa_tree_add_6_33_groupi_n_3583);
  xnor csa_tree_add_6_33_groupi_g14382__5107(csa_tree_add_6_33_groupi_n_3955 ,csa_tree_add_6_33_groupi_n_3190 ,csa_tree_add_6_33_groupi_n_3575);
  xnor csa_tree_add_6_33_groupi_g14383__6260(csa_tree_add_6_33_groupi_n_3953 ,csa_tree_add_6_33_groupi_n_3475 ,csa_tree_add_6_33_groupi_n_3576);
  or csa_tree_add_6_33_groupi_g14384__4319(csa_tree_add_6_33_groupi_n_3910 ,csa_tree_add_6_33_groupi_n_3036 ,csa_tree_add_6_33_groupi_n_3625);
  or csa_tree_add_6_33_groupi_g14385__8428(csa_tree_add_6_33_groupi_n_3909 ,csa_tree_add_6_33_groupi_n_3462 ,csa_tree_add_6_33_groupi_n_3666);
  or csa_tree_add_6_33_groupi_g14386__5526(csa_tree_add_6_33_groupi_n_3908 ,csa_tree_add_6_33_groupi_n_3522 ,csa_tree_add_6_33_groupi_n_3665);
  or csa_tree_add_6_33_groupi_g14387__6783(csa_tree_add_6_33_groupi_n_3907 ,csa_tree_add_6_33_groupi_n_3565 ,csa_tree_add_6_33_groupi_n_3753);
  nor csa_tree_add_6_33_groupi_g14388__3680(csa_tree_add_6_33_groupi_n_3906 ,csa_tree_add_6_33_groupi_n_3523 ,csa_tree_add_6_33_groupi_n_3664);
  or csa_tree_add_6_33_groupi_g14389__1617(csa_tree_add_6_33_groupi_n_3905 ,csa_tree_add_6_33_groupi_n_3546 ,csa_tree_add_6_33_groupi_n_3752);
  and csa_tree_add_6_33_groupi_g14390__2802(csa_tree_add_6_33_groupi_n_3904 ,csa_tree_add_6_33_groupi_n_3446 ,csa_tree_add_6_33_groupi_n_3642);
  or csa_tree_add_6_33_groupi_g14391__1705(csa_tree_add_6_33_groupi_n_3903 ,csa_tree_add_6_33_groupi_n_3535 ,csa_tree_add_6_33_groupi_n_3662);
  nor csa_tree_add_6_33_groupi_g14392__5122(csa_tree_add_6_33_groupi_n_3902 ,csa_tree_add_6_33_groupi_n_3408 ,csa_tree_add_6_33_groupi_n_3612);
  or csa_tree_add_6_33_groupi_g14393__8246(csa_tree_add_6_33_groupi_n_3901 ,csa_tree_add_6_33_groupi_n_3444 ,csa_tree_add_6_33_groupi_n_3640);
  and csa_tree_add_6_33_groupi_g14394__7098(csa_tree_add_6_33_groupi_n_3900 ,csa_tree_add_6_33_groupi_n_3535 ,csa_tree_add_6_33_groupi_n_3662);
  or csa_tree_add_6_33_groupi_g14395__6131(csa_tree_add_6_33_groupi_n_3899 ,csa_tree_add_6_33_groupi_n_3409 ,csa_tree_add_6_33_groupi_n_3611);
  or csa_tree_add_6_33_groupi_g14396__1881(csa_tree_add_6_33_groupi_n_3898 ,csa_tree_add_6_33_groupi_n_3459 ,csa_tree_add_6_33_groupi_n_3661);
  and csa_tree_add_6_33_groupi_g14397__5115(csa_tree_add_6_33_groupi_n_3897 ,csa_tree_add_6_33_groupi_n_3459 ,csa_tree_add_6_33_groupi_n_3661);
  or csa_tree_add_6_33_groupi_g14398__7482(csa_tree_add_6_33_groupi_n_3896 ,csa_tree_add_6_33_groupi_n_3559 ,csa_tree_add_6_33_groupi_n_3689);
  and csa_tree_add_6_33_groupi_g14399__4733(csa_tree_add_6_33_groupi_n_3895 ,csa_tree_add_6_33_groupi_n_3462 ,csa_tree_add_6_33_groupi_n_3666);
  or csa_tree_add_6_33_groupi_g14400__6161(csa_tree_add_6_33_groupi_n_3894 ,csa_tree_add_6_33_groupi_n_3552 ,csa_tree_add_6_33_groupi_n_3746);
  or csa_tree_add_6_33_groupi_g14401__9315(csa_tree_add_6_33_groupi_n_3893 ,csa_tree_add_6_33_groupi_n_3533 ,csa_tree_add_6_33_groupi_n_3658);
  nor csa_tree_add_6_33_groupi_g14402__9945(csa_tree_add_6_33_groupi_n_3892 ,csa_tree_add_6_33_groupi_n_3035 ,csa_tree_add_6_33_groupi_n_3626);
  nor csa_tree_add_6_33_groupi_g14403__2883(csa_tree_add_6_33_groupi_n_3891 ,csa_tree_add_6_33_groupi_n_3530 ,csa_tree_add_6_33_groupi_n_3660);
  and csa_tree_add_6_33_groupi_g14404__2346(csa_tree_add_6_33_groupi_n_3890 ,csa_tree_add_6_33_groupi_n_3533 ,csa_tree_add_6_33_groupi_n_3658);
  or csa_tree_add_6_33_groupi_g14405__1666(csa_tree_add_6_33_groupi_n_3889 ,csa_tree_add_6_33_groupi_n_3763 ,csa_tree_add_6_33_groupi_n_3653);
  or csa_tree_add_6_33_groupi_g14406__7410(csa_tree_add_6_33_groupi_n_3888 ,csa_tree_add_6_33_groupi_n_3055 ,csa_tree_add_6_33_groupi_n_3656);
  or csa_tree_add_6_33_groupi_g14407__6417(csa_tree_add_6_33_groupi_n_3887 ,csa_tree_add_6_33_groupi_n_3553 ,csa_tree_add_6_33_groupi_n_3742);
  or csa_tree_add_6_33_groupi_g14408__5477(csa_tree_add_6_33_groupi_n_3886 ,csa_tree_add_6_33_groupi_n_3539 ,csa_tree_add_6_33_groupi_n_3615);
  nor csa_tree_add_6_33_groupi_g14409__2398(csa_tree_add_6_33_groupi_n_3885 ,csa_tree_add_6_33_groupi_n_3538 ,csa_tree_add_6_33_groupi_n_3616);
  or csa_tree_add_6_33_groupi_g14410__5107(csa_tree_add_6_33_groupi_n_3884 ,csa_tree_add_6_33_groupi_n_3554 ,csa_tree_add_6_33_groupi_n_3740);
  or csa_tree_add_6_33_groupi_g14411__6260(csa_tree_add_6_33_groupi_n_3883 ,csa_tree_add_6_33_groupi_n_3555 ,csa_tree_add_6_33_groupi_n_3737);
  and csa_tree_add_6_33_groupi_g14412__4319(csa_tree_add_6_33_groupi_n_3882 ,csa_tree_add_6_33_groupi_n_3763 ,csa_tree_add_6_33_groupi_n_3653);
  or csa_tree_add_6_33_groupi_g14413__8428(csa_tree_add_6_33_groupi_n_3881 ,csa_tree_add_6_33_groupi_n_3380 ,csa_tree_add_6_33_groupi_n_3598);
  or csa_tree_add_6_33_groupi_g14414__5526(csa_tree_add_6_33_groupi_n_3880 ,csa_tree_add_6_33_groupi_n_3454 ,csa_tree_add_6_33_groupi_n_3621);
  or csa_tree_add_6_33_groupi_g14415__6783(csa_tree_add_6_33_groupi_n_3879 ,csa_tree_add_6_33_groupi_n_3569 ,csa_tree_add_6_33_groupi_n_3755);
  or csa_tree_add_6_33_groupi_g14416__3680(csa_tree_add_6_33_groupi_n_3878 ,csa_tree_add_6_33_groupi_n_3562 ,csa_tree_add_6_33_groupi_n_3695);
  or csa_tree_add_6_33_groupi_g14417__1617(csa_tree_add_6_33_groupi_n_3877 ,csa_tree_add_6_33_groupi_n_3450 ,csa_tree_add_6_33_groupi_n_3663);
  or csa_tree_add_6_33_groupi_g14418__2802(csa_tree_add_6_33_groupi_n_3876 ,csa_tree_add_6_33_groupi_n_3537 ,csa_tree_add_6_33_groupi_n_3648);
  nor csa_tree_add_6_33_groupi_g14419__1705(csa_tree_add_6_33_groupi_n_3875 ,csa_tree_add_6_33_groupi_n_3453 ,csa_tree_add_6_33_groupi_n_3622);
  and csa_tree_add_6_33_groupi_g14420__5122(csa_tree_add_6_33_groupi_n_3874 ,csa_tree_add_6_33_groupi_n_3450 ,csa_tree_add_6_33_groupi_n_3663);
  or csa_tree_add_6_33_groupi_g14421__8246(csa_tree_add_6_33_groupi_n_3873 ,csa_tree_add_6_33_groupi_n_3771 ,csa_tree_add_6_33_groupi_n_3718);
  and csa_tree_add_6_33_groupi_g14422__7098(csa_tree_add_6_33_groupi_n_3872 ,csa_tree_add_6_33_groupi_n_3496 ,csa_tree_add_6_33_groupi_n_3673);
  or csa_tree_add_6_33_groupi_g14423__6131(csa_tree_add_6_33_groupi_n_3871 ,csa_tree_add_6_33_groupi_n_3563 ,csa_tree_add_6_33_groupi_n_3696);
  and csa_tree_add_6_33_groupi_g14424__1881(csa_tree_add_6_33_groupi_n_3870 ,csa_tree_add_6_33_groupi_n_3537 ,csa_tree_add_6_33_groupi_n_3648);
  and csa_tree_add_6_33_groupi_g14425__5115(csa_tree_add_6_33_groupi_n_3869 ,csa_tree_add_6_33_groupi_n_3055 ,csa_tree_add_6_33_groupi_n_3656);
  or csa_tree_add_6_33_groupi_g14426__7482(csa_tree_add_6_33_groupi_n_3868 ,csa_tree_add_6_33_groupi_n_3531 ,csa_tree_add_6_33_groupi_n_3659);
  or csa_tree_add_6_33_groupi_g14427__4733(csa_tree_add_6_33_groupi_n_3867 ,csa_tree_add_6_33_groupi_n_3384 ,csa_tree_add_6_33_groupi_n_3723);
  or csa_tree_add_6_33_groupi_g14428__6161(csa_tree_add_6_33_groupi_n_3866 ,csa_tree_add_6_33_groupi_n_3486 ,csa_tree_add_6_33_groupi_n_3713);
  or csa_tree_add_6_33_groupi_g14429__9315(csa_tree_add_6_33_groupi_n_3865 ,csa_tree_add_6_33_groupi_n_3386 ,csa_tree_add_6_33_groupi_n_3721);
  and csa_tree_add_6_33_groupi_g14430__9945(csa_tree_add_6_33_groupi_n_3864 ,csa_tree_add_6_33_groupi_n_3641 ,csa_tree_add_6_33_groupi_n_3649);
  and csa_tree_add_6_33_groupi_g14431__2883(csa_tree_add_6_33_groupi_n_3863 ,csa_tree_add_6_33_groupi_n_3542 ,csa_tree_add_6_33_groupi_n_3643);
  or csa_tree_add_6_33_groupi_g14432__2346(csa_tree_add_6_33_groupi_n_3862 ,csa_tree_add_6_33_groupi_n_3542 ,csa_tree_add_6_33_groupi_n_3643);
  and csa_tree_add_6_33_groupi_g14433__1666(csa_tree_add_6_33_groupi_n_3861 ,csa_tree_add_6_33_groupi_n_3295 ,csa_tree_add_6_33_groupi_n_3672);
  or csa_tree_add_6_33_groupi_g14434__7410(csa_tree_add_6_33_groupi_n_3860 ,csa_tree_add_6_33_groupi_n_3446 ,csa_tree_add_6_33_groupi_n_3642);
  nor csa_tree_add_6_33_groupi_g14435__6417(csa_tree_add_6_33_groupi_n_3859 ,csa_tree_add_6_33_groupi_n_3639 ,csa_tree_add_6_33_groupi_n_3633);
  or csa_tree_add_6_33_groupi_g14436__5477(csa_tree_add_6_33_groupi_n_3858 ,csa_tree_add_6_33_groupi_n_3638 ,csa_tree_add_6_33_groupi_n_3634);
  and csa_tree_add_6_33_groupi_g14437__2398(csa_tree_add_6_33_groupi_n_3857 ,csa_tree_add_6_33_groupi_n_3444 ,csa_tree_add_6_33_groupi_n_3640);
  or csa_tree_add_6_33_groupi_g14438__5107(csa_tree_add_6_33_groupi_n_3856 ,csa_tree_add_6_33_groupi_n_3571 ,csa_tree_add_6_33_groupi_n_3722);
  or csa_tree_add_6_33_groupi_g14439__6260(csa_tree_add_6_33_groupi_n_3855 ,csa_tree_add_6_33_groupi_n_3572 ,csa_tree_add_6_33_groupi_n_3693);
  or csa_tree_add_6_33_groupi_g14440__4319(csa_tree_add_6_33_groupi_n_3854 ,csa_tree_add_6_33_groupi_n_3558 ,csa_tree_add_6_33_groupi_n_3716);
  or csa_tree_add_6_33_groupi_g14441__8428(csa_tree_add_6_33_groupi_n_3853 ,csa_tree_add_6_33_groupi_n_3568 ,csa_tree_add_6_33_groupi_n_3700);
  or csa_tree_add_6_33_groupi_g14442__5526(csa_tree_add_6_33_groupi_n_3852 ,csa_tree_add_6_33_groupi_n_3637 ,csa_tree_add_6_33_groupi_n_3636);
  or csa_tree_add_6_33_groupi_g14443__6783(csa_tree_add_6_33_groupi_n_3851 ,csa_tree_add_6_33_groupi_n_3387 ,csa_tree_add_6_33_groupi_n_3701);
  and csa_tree_add_6_33_groupi_g14444__3680(csa_tree_add_6_33_groupi_n_3850 ,csa_tree_add_6_33_groupi_n_3637 ,csa_tree_add_6_33_groupi_n_3636);
  or csa_tree_add_6_33_groupi_g14445__1617(csa_tree_add_6_33_groupi_n_3849 ,csa_tree_add_6_33_groupi_n_3674 ,csa_tree_add_6_33_groupi_n_3704);
  and csa_tree_add_6_33_groupi_g14446__2802(csa_tree_add_6_33_groupi_n_3920 ,csa_tree_add_6_33_groupi_n_3489 ,csa_tree_add_6_33_groupi_n_3708);
  and csa_tree_add_6_33_groupi_g14447__1705(csa_tree_add_6_33_groupi_n_3919 ,csa_tree_add_6_33_groupi_n_3492 ,csa_tree_add_6_33_groupi_n_3698);
  and csa_tree_add_6_33_groupi_g14448__5122(csa_tree_add_6_33_groupi_n_3918 ,csa_tree_add_6_33_groupi_n_3332 ,csa_tree_add_6_33_groupi_n_3702);
  or csa_tree_add_6_33_groupi_g14449__8246(csa_tree_add_6_33_groupi_n_3917 ,csa_tree_add_6_33_groupi_n_3518 ,csa_tree_add_6_33_groupi_n_3750);
  and csa_tree_add_6_33_groupi_g14450__7098(csa_tree_add_6_33_groupi_n_3916 ,csa_tree_add_6_33_groupi_n_3509 ,csa_tree_add_6_33_groupi_n_3745);
  and csa_tree_add_6_33_groupi_g14451__6131(csa_tree_add_6_33_groupi_n_3915 ,csa_tree_add_6_33_groupi_n_3500 ,csa_tree_add_6_33_groupi_n_3692);
  and csa_tree_add_6_33_groupi_g14452__1881(csa_tree_add_6_33_groupi_n_3914 ,csa_tree_add_6_33_groupi_n_3138 ,csa_tree_add_6_33_groupi_n_3731);
  and csa_tree_add_6_33_groupi_g14453__5115(csa_tree_add_6_33_groupi_n_3913 ,csa_tree_add_6_33_groupi_n_3513 ,csa_tree_add_6_33_groupi_n_3747);
  or csa_tree_add_6_33_groupi_g14454__7482(csa_tree_add_6_33_groupi_n_3912 ,csa_tree_add_6_33_groupi_n_3504 ,csa_tree_add_6_33_groupi_n_3728);
  or csa_tree_add_6_33_groupi_g14455__4733(csa_tree_add_6_33_groupi_n_3911 ,csa_tree_add_6_33_groupi_n_3116 ,csa_tree_add_6_33_groupi_n_3724);
  not csa_tree_add_6_33_groupi_g14456(csa_tree_add_6_33_groupi_n_3844 ,csa_tree_add_6_33_groupi_n_3845);
  not csa_tree_add_6_33_groupi_g14457(csa_tree_add_6_33_groupi_n_3839 ,csa_tree_add_6_33_groupi_n_3840);
  not csa_tree_add_6_33_groupi_g14458(csa_tree_add_6_33_groupi_n_3837 ,csa_tree_add_6_33_groupi_n_3838);
  nor csa_tree_add_6_33_groupi_g14459__6161(csa_tree_add_6_33_groupi_n_3835 ,csa_tree_add_6_33_groupi_n_3540 ,csa_tree_add_6_33_groupi_n_3629);
  or csa_tree_add_6_33_groupi_g14460(csa_tree_add_6_33_groupi_n_3834 ,csa_tree_add_6_33_groupi_n_3557 ,csa_tree_add_6_33_groupi_n_3685);
  or csa_tree_add_6_33_groupi_g14461(csa_tree_add_6_33_groupi_n_3833 ,csa_tree_add_6_33_groupi_n_3556 ,csa_tree_add_6_33_groupi_n_3686);
  or csa_tree_add_6_33_groupi_g14462(csa_tree_add_6_33_groupi_n_3832 ,csa_tree_add_6_33_groupi_n_3541 ,csa_tree_add_6_33_groupi_n_3628);
  nor csa_tree_add_6_33_groupi_g14463(csa_tree_add_6_33_groupi_n_3831 ,csa_tree_add_6_33_groupi_n_3473 ,csa_tree_add_6_33_groupi_n_3759);
  or csa_tree_add_6_33_groupi_g14464(csa_tree_add_6_33_groupi_n_3830 ,csa_tree_add_6_33_groupi_n_3472 ,csa_tree_add_6_33_groupi_n_3760);
  or csa_tree_add_6_33_groupi_g14465(csa_tree_add_6_33_groupi_n_3829 ,csa_tree_add_6_33_groupi_n_3373 ,csa_tree_add_6_33_groupi_n_3684);
  or csa_tree_add_6_33_groupi_g14466(csa_tree_add_6_33_groupi_n_3828 ,csa_tree_add_6_33_groupi_n_3291 ,csa_tree_add_6_33_groupi_n_3706);
  or csa_tree_add_6_33_groupi_g14467(csa_tree_add_6_33_groupi_n_3827 ,csa_tree_add_6_33_groupi_n_3528 ,csa_tree_add_6_33_groupi_n_3623);
  or csa_tree_add_6_33_groupi_g14468(csa_tree_add_6_33_groupi_n_3826 ,csa_tree_add_6_33_groupi_n_3435 ,csa_tree_add_6_33_groupi_n_3644);
  nor csa_tree_add_6_33_groupi_g14469(csa_tree_add_6_33_groupi_n_3825 ,csa_tree_add_6_33_groupi_n_3434 ,csa_tree_add_6_33_groupi_n_3645);
  or csa_tree_add_6_33_groupi_g14470(csa_tree_add_6_33_groupi_n_3824 ,csa_tree_add_6_33_groupi_n_3682 ,csa_tree_add_6_33_groupi_n_3717);
  or csa_tree_add_6_33_groupi_g14471(csa_tree_add_6_33_groupi_n_3823 ,csa_tree_add_6_33_groupi_n_3290 ,csa_tree_add_6_33_groupi_n_3738);
  or csa_tree_add_6_33_groupi_g14472(csa_tree_add_6_33_groupi_n_3822 ,csa_tree_add_6_33_groupi_n_3466 ,csa_tree_add_6_33_groupi_n_3620);
  or csa_tree_add_6_33_groupi_g14473(csa_tree_add_6_33_groupi_n_3821 ,csa_tree_add_6_33_groupi_n_3641 ,csa_tree_add_6_33_groupi_n_3649);
  and csa_tree_add_6_33_groupi_g14474(csa_tree_add_6_33_groupi_n_3820 ,csa_tree_add_6_33_groupi_n_3528 ,csa_tree_add_6_33_groupi_n_3623);
  or csa_tree_add_6_33_groupi_g14475(csa_tree_add_6_33_groupi_n_3819 ,csa_tree_add_6_33_groupi_n_3289 ,csa_tree_add_6_33_groupi_n_3594);
  and csa_tree_add_6_33_groupi_g14476(csa_tree_add_6_33_groupi_n_3818 ,csa_tree_add_6_33_groupi_n_3466 ,csa_tree_add_6_33_groupi_n_3620);
  or csa_tree_add_6_33_groupi_g14477(csa_tree_add_6_33_groupi_n_3817 ,csa_tree_add_6_33_groupi_n_3283 ,csa_tree_add_6_33_groupi_n_3604);
  or csa_tree_add_6_33_groupi_g14478(csa_tree_add_6_33_groupi_n_3816 ,csa_tree_add_6_33_groupi_n_3619 ,csa_tree_add_6_33_groupi_n_3646);
  nor csa_tree_add_6_33_groupi_g14479(csa_tree_add_6_33_groupi_n_3815 ,csa_tree_add_6_33_groupi_n_3618 ,csa_tree_add_6_33_groupi_n_3647);
  nor csa_tree_add_6_33_groupi_g14480(csa_tree_add_6_33_groupi_n_3814 ,csa_tree_add_6_33_groupi_n_3284 ,csa_tree_add_6_33_groupi_n_3725);
  or csa_tree_add_6_33_groupi_g14481(csa_tree_add_6_33_groupi_n_3813 ,csa_tree_add_6_33_groupi_n_3414 ,csa_tree_add_6_33_groupi_n_3617);
  and csa_tree_add_6_33_groupi_g14482(csa_tree_add_6_33_groupi_n_3812 ,csa_tree_add_6_33_groupi_n_3414 ,csa_tree_add_6_33_groupi_n_3617);
  or csa_tree_add_6_33_groupi_g14483(csa_tree_add_6_33_groupi_n_3811 ,csa_tree_add_6_33_groupi_n_3413 ,csa_tree_add_6_33_groupi_n_3669);
  and csa_tree_add_6_33_groupi_g14484(csa_tree_add_6_33_groupi_n_3810 ,csa_tree_add_6_33_groupi_n_3413 ,csa_tree_add_6_33_groupi_n_3669);
  or csa_tree_add_6_33_groupi_g14485(csa_tree_add_6_33_groupi_n_3809 ,csa_tree_add_6_33_groupi_n_3281 ,csa_tree_add_6_33_groupi_n_3756);
  or csa_tree_add_6_33_groupi_g14486(csa_tree_add_6_33_groupi_n_3808 ,csa_tree_add_6_33_groupi_n_3482 ,csa_tree_add_6_33_groupi_n_3757);
  xnor csa_tree_add_6_33_groupi_g14487(csa_tree_add_6_33_groupi_n_3807 ,csa_tree_add_6_33_groupi_n_3418 ,csa_tree_add_6_33_groupi_n_3419);
  xnor csa_tree_add_6_33_groupi_g14488(csa_tree_add_6_33_groupi_n_3806 ,csa_tree_add_6_33_groupi_n_3544 ,csa_tree_add_6_33_groupi_n_3433);
  xnor csa_tree_add_6_33_groupi_g14489(csa_tree_add_6_33_groupi_n_3805 ,csa_tree_add_6_33_groupi_n_3423 ,csa_tree_add_6_33_groupi_n_3430);
  xnor csa_tree_add_6_33_groupi_g14490(csa_tree_add_6_33_groupi_n_3804 ,csa_tree_add_6_33_groupi_n_3557 ,csa_tree_add_6_33_groupi_n_3189);
  xnor csa_tree_add_6_33_groupi_g14491(csa_tree_add_6_33_groupi_n_3803 ,csa_tree_add_6_33_groupi_n_3556 ,csa_tree_add_6_33_groupi_n_3425);
  xnor csa_tree_add_6_33_groupi_g14492(csa_tree_add_6_33_groupi_n_3802 ,csa_tree_add_6_33_groupi_n_3277 ,csa_tree_add_6_33_groupi_n_3555);
  xnor csa_tree_add_6_33_groupi_g14493(csa_tree_add_6_33_groupi_n_3801 ,csa_tree_add_6_33_groupi_n_3461 ,csa_tree_add_6_33_groupi_n_3565);
  xnor csa_tree_add_6_33_groupi_g14494(csa_tree_add_6_33_groupi_n_3800 ,csa_tree_add_6_33_groupi_n_3414 ,csa_tree_add_6_33_groupi_n_3483);
  xnor csa_tree_add_6_33_groupi_g14495(csa_tree_add_6_33_groupi_n_3799 ,csa_tree_add_6_33_groupi_n_3345 ,csa_tree_add_6_33_groupi_n_3571);
  xnor csa_tree_add_6_33_groupi_g14496(csa_tree_add_6_33_groupi_n_3798 ,csa_tree_add_6_33_groupi_n_3370 ,csa_tree_add_6_33_groupi_n_3469);
  xnor csa_tree_add_6_33_groupi_g14497(csa_tree_add_6_33_groupi_n_3797 ,csa_tree_add_6_33_groupi_n_3270 ,csa_tree_add_6_33_groupi_n_3470);
  xnor csa_tree_add_6_33_groupi_g14498(csa_tree_add_6_33_groupi_n_3796 ,csa_tree_add_6_33_groupi_n_3568 ,csa_tree_add_6_33_groupi_n_3467);
  xnor csa_tree_add_6_33_groupi_g14499(csa_tree_add_6_33_groupi_n_3795 ,csa_tree_add_6_33_groupi_n_3420 ,csa_tree_add_6_33_groupi_n_3278);
  xnor csa_tree_add_6_33_groupi_g14500(csa_tree_add_6_33_groupi_n_3794 ,csa_tree_add_6_33_groupi_n_3547 ,csa_tree_add_6_33_groupi_n_3466);
  xnor csa_tree_add_6_33_groupi_g14501(csa_tree_add_6_33_groupi_n_3793 ,csa_tree_add_6_33_groupi_n_3413 ,csa_tree_add_6_33_groupi_n_3487);
  xnor csa_tree_add_6_33_groupi_g14502(csa_tree_add_6_33_groupi_n_3792 ,csa_tree_add_6_33_groupi_n_3411 ,csa_tree_add_6_33_groupi_n_3482);
  xnor csa_tree_add_6_33_groupi_g14503(csa_tree_add_6_33_groupi_n_3791 ,csa_tree_add_6_33_groupi_n_3546 ,csa_tree_add_6_33_groupi_n_3352);
  xnor csa_tree_add_6_33_groupi_g14504(csa_tree_add_6_33_groupi_n_3790 ,csa_tree_add_6_33_groupi_n_3445 ,csa_tree_add_6_33_groupi_n_2682);
  xnor csa_tree_add_6_33_groupi_g14505(csa_tree_add_6_33_groupi_n_3789 ,csa_tree_add_6_33_groupi_n_3527 ,csa_tree_add_6_33_groupi_n_3283);
  xnor csa_tree_add_6_33_groupi_g14506(csa_tree_add_6_33_groupi_n_3788 ,csa_tree_add_6_33_groupi_n_3554 ,csa_tree_add_6_33_groupi_n_3365);
  xnor csa_tree_add_6_33_groupi_g14507(csa_tree_add_6_33_groupi_n_3787 ,csa_tree_add_6_33_groupi_n_3549 ,csa_tree_add_6_33_groupi_n_3462);
  xnor csa_tree_add_6_33_groupi_g14508(csa_tree_add_6_33_groupi_n_3786 ,csa_tree_add_6_33_groupi_n_3457 ,csa_tree_add_6_33_groupi_n_3458);
  xnor csa_tree_add_6_33_groupi_g14509(csa_tree_add_6_33_groupi_n_3785 ,csa_tree_add_6_33_groupi_n_3454 ,csa_tree_add_6_33_groupi_n_3560);
  xnor csa_tree_add_6_33_groupi_g14510(csa_tree_add_6_33_groupi_n_3784 ,csa_tree_add_6_33_groupi_n_3451 ,csa_tree_add_6_33_groupi_n_3452);
  xnor csa_tree_add_6_33_groupi_g14511(csa_tree_add_6_33_groupi_n_3783 ,csa_tree_add_6_33_groupi_n_3545 ,csa_tree_add_6_33_groupi_n_3384);
  xnor csa_tree_add_6_33_groupi_g14512(csa_tree_add_6_33_groupi_n_3782 ,csa_tree_add_6_33_groupi_n_3532 ,csa_tree_add_6_33_groupi_n_3048);
  xnor csa_tree_add_6_33_groupi_g14513(csa_tree_add_6_33_groupi_n_3781 ,csa_tree_add_6_33_groupi_n_3446 ,csa_tree_add_6_33_groupi_n_3564);
  xnor csa_tree_add_6_33_groupi_g14514(csa_tree_add_6_33_groupi_n_3780 ,csa_tree_add_6_33_groupi_n_3447 ,csa_tree_add_6_33_groupi_n_3269);
  xnor csa_tree_add_6_33_groupi_g14515(csa_tree_add_6_33_groupi_n_3779 ,csa_tree_add_6_33_groupi_n_3486 ,csa_tree_add_6_33_groupi_n_3186);
  xnor csa_tree_add_6_33_groupi_g14516(csa_tree_add_6_33_groupi_n_3778 ,csa_tree_add_6_33_groupi_n_3428 ,csa_tree_add_6_33_groupi_n_3364);
  xnor csa_tree_add_6_33_groupi_g14517(csa_tree_add_6_33_groupi_n_3777 ,csa_tree_add_6_33_groupi_n_3421 ,csa_tree_add_6_33_groupi_n_3534);
  xnor csa_tree_add_6_33_groupi_g14518(csa_tree_add_6_33_groupi_n_3776 ,csa_tree_add_6_33_groupi_n_3437 ,csa_tree_add_6_33_groupi_n_3367);
  xnor csa_tree_add_6_33_groupi_g14519(csa_tree_add_6_33_groupi_n_3775 ,csa_tree_add_6_33_groupi_n_3441 ,csa_tree_add_6_33_groupi_n_3371);
  xnor csa_tree_add_6_33_groupi_g14520(csa_tree_add_6_33_groupi_n_3774 ,csa_tree_add_6_33_groupi_n_3563 ,csa_tree_add_6_33_groupi_n_3366);
  xnor csa_tree_add_6_33_groupi_g14521(csa_tree_add_6_33_groupi_n_3773 ,csa_tree_add_6_33_groupi_n_3273 ,csa_tree_add_6_33_groupi_n_3456);
  and csa_tree_add_6_33_groupi_g14522(csa_tree_add_6_33_groupi_n_3848 ,csa_tree_add_6_33_groupi_n_3401 ,csa_tree_add_6_33_groupi_n_3599);
  and csa_tree_add_6_33_groupi_g14523(csa_tree_add_6_33_groupi_n_3847 ,csa_tree_add_6_33_groupi_n_3507 ,csa_tree_add_6_33_groupi_n_3683);
  and csa_tree_add_6_33_groupi_g14524(csa_tree_add_6_33_groupi_n_3846 ,csa_tree_add_6_33_groupi_n_3505 ,csa_tree_add_6_33_groupi_n_3733);
  xnor csa_tree_add_6_33_groupi_g14525(csa_tree_add_6_33_groupi_n_3845 ,csa_tree_add_6_33_groupi_n_3372 ,csa_tree_add_6_33_groupi_n_3393);
  xnor csa_tree_add_6_33_groupi_g14526(csa_tree_add_6_33_groupi_n_3843 ,csa_tree_add_6_33_groupi_n_3567 ,csa_tree_add_6_33_groupi_n_3396);
  xnor csa_tree_add_6_33_groupi_g14527(csa_tree_add_6_33_groupi_n_3842 ,csa_tree_add_6_33_groupi_n_3388 ,csa_tree_add_6_33_groupi_n_3394);
  xnor csa_tree_add_6_33_groupi_g14528(csa_tree_add_6_33_groupi_n_3841 ,csa_tree_add_6_33_groupi_n_3480 ,csa_tree_add_6_33_groupi_n_3216);
  xnor csa_tree_add_6_33_groupi_g14529(csa_tree_add_6_33_groupi_n_3840 ,csa_tree_add_6_33_groupi_n_3286 ,csa_tree_add_6_33_groupi_n_3392);
  xnor csa_tree_add_6_33_groupi_g14530(csa_tree_add_6_33_groupi_n_3838 ,csa_tree_add_6_33_groupi_n_3484 ,csa_tree_add_6_33_groupi_n_3233);
  xnor csa_tree_add_6_33_groupi_g14531(csa_tree_add_6_33_groupi_n_3836 ,csa_tree_add_6_33_groupi_n_3385 ,csa_tree_add_6_33_groupi_n_3391);
  not csa_tree_add_6_33_groupi_g14532(csa_tree_add_6_33_groupi_n_3759 ,csa_tree_add_6_33_groupi_n_3760);
  or csa_tree_add_6_33_groupi_g14533(csa_tree_add_6_33_groupi_n_3758 ,csa_tree_add_6_33_groupi_n_3186 ,csa_tree_add_6_33_groupi_n_3468);
  nor csa_tree_add_6_33_groupi_g14534(csa_tree_add_6_33_groupi_n_3757 ,csa_tree_add_6_33_groupi_n_3465 ,csa_tree_add_6_33_groupi_n_3410);
  and csa_tree_add_6_33_groupi_g14535(csa_tree_add_6_33_groupi_n_3756 ,csa_tree_add_6_33_groupi_n_3279 ,csa_tree_add_6_33_groupi_n_3412);
  and csa_tree_add_6_33_groupi_g14536(csa_tree_add_6_33_groupi_n_3755 ,csa_tree_add_6_33_groupi_n_3452 ,csa_tree_add_6_33_groupi_n_3451);
  or csa_tree_add_6_33_groupi_g14537(csa_tree_add_6_33_groupi_n_3754 ,csa_tree_add_6_33_groupi_n_3352 ,csa_tree_add_6_33_groupi_n_3406);
  and csa_tree_add_6_33_groupi_g14538(csa_tree_add_6_33_groupi_n_3753 ,csa_tree_add_6_33_groupi_n_3463 ,csa_tree_add_6_33_groupi_n_3461);
  nor csa_tree_add_6_33_groupi_g14539(csa_tree_add_6_33_groupi_n_3752 ,csa_tree_add_6_33_groupi_n_3351 ,csa_tree_add_6_33_groupi_n_3407);
  or csa_tree_add_6_33_groupi_g14540(csa_tree_add_6_33_groupi_n_3751 ,csa_tree_add_6_33_groupi_n_3527 ,csa_tree_add_6_33_groupi_n_3449);
  nor csa_tree_add_6_33_groupi_g14541(csa_tree_add_6_33_groupi_n_3750 ,csa_tree_add_6_33_groupi_n_3516 ,csa_tree_add_6_33_groupi_n_3551);
  nor csa_tree_add_6_33_groupi_g14542(csa_tree_add_6_33_groupi_n_3749 ,csa_tree_add_6_33_groupi_n_3543 ,csa_tree_add_6_33_groupi_n_3433);
  or csa_tree_add_6_33_groupi_g14543(csa_tree_add_6_33_groupi_n_3748 ,csa_tree_add_6_33_groupi_n_3458 ,csa_tree_add_6_33_groupi_n_3457);
  or csa_tree_add_6_33_groupi_g14544(csa_tree_add_6_33_groupi_n_3747 ,csa_tree_add_6_33_groupi_n_3511 ,csa_tree_add_6_33_groupi_n_3479);
  and csa_tree_add_6_33_groupi_g14545(csa_tree_add_6_33_groupi_n_3746 ,csa_tree_add_6_33_groupi_n_3458 ,csa_tree_add_6_33_groupi_n_3457);
  or csa_tree_add_6_33_groupi_g14546(csa_tree_add_6_33_groupi_n_3745 ,csa_tree_add_6_33_groupi_n_3190 ,csa_tree_add_6_33_groupi_n_3508);
  or csa_tree_add_6_33_groupi_g14547(csa_tree_add_6_33_groupi_n_3744 ,csa_tree_add_6_33_groupi_n_3272 ,csa_tree_add_6_33_groupi_n_3456);
  or csa_tree_add_6_33_groupi_g14548(csa_tree_add_6_33_groupi_n_3743 ,csa_tree_add_6_33_groupi_n_3044 ,csa_tree_add_6_33_groupi_n_3417);
  nor csa_tree_add_6_33_groupi_g14549(csa_tree_add_6_33_groupi_n_3742 ,csa_tree_add_6_33_groupi_n_3273 ,csa_tree_add_6_33_groupi_n_3455);
  or csa_tree_add_6_33_groupi_g14550(csa_tree_add_6_33_groupi_n_3741 ,csa_tree_add_6_33_groupi_n_3365 ,csa_tree_add_6_33_groupi_n_3476);
  and csa_tree_add_6_33_groupi_g14551(csa_tree_add_6_33_groupi_n_3740 ,csa_tree_add_6_33_groupi_n_3365 ,csa_tree_add_6_33_groupi_n_3476);
  or csa_tree_add_6_33_groupi_g14552(csa_tree_add_6_33_groupi_n_3739 ,csa_tree_add_6_33_groupi_n_3276 ,csa_tree_add_6_33_groupi_n_3415);
  nor csa_tree_add_6_33_groupi_g14553(csa_tree_add_6_33_groupi_n_3738 ,csa_tree_add_6_33_groupi_n_3041 ,csa_tree_add_6_33_groupi_n_3440);
  nor csa_tree_add_6_33_groupi_g14554(csa_tree_add_6_33_groupi_n_3737 ,csa_tree_add_6_33_groupi_n_3277 ,csa_tree_add_6_33_groupi_n_3416);
  and csa_tree_add_6_33_groupi_g14555(csa_tree_add_6_33_groupi_n_3736 ,csa_tree_add_6_33_groupi_n_3048 ,csa_tree_add_6_33_groupi_n_3532);
  or csa_tree_add_6_33_groupi_g14556(csa_tree_add_6_33_groupi_n_3735 ,csa_tree_add_6_33_groupi_n_3452 ,csa_tree_add_6_33_groupi_n_3451);
  or csa_tree_add_6_33_groupi_g14557(csa_tree_add_6_33_groupi_n_3734 ,csa_tree_add_6_33_groupi_n_3269 ,csa_tree_add_6_33_groupi_n_3447);
  or csa_tree_add_6_33_groupi_g14558(csa_tree_add_6_33_groupi_n_3733 ,csa_tree_add_6_33_groupi_n_3520 ,csa_tree_add_6_33_groupi_n_3548);
  or csa_tree_add_6_33_groupi_g14559(csa_tree_add_6_33_groupi_n_3732 ,csa_tree_add_6_33_groupi_n_3042 ,csa_tree_add_6_33_groupi_n_3439);
  or csa_tree_add_6_33_groupi_g14560(csa_tree_add_6_33_groupi_n_3731 ,csa_tree_add_6_33_groupi_n_3123 ,csa_tree_add_6_33_groupi_n_3484);
  or csa_tree_add_6_33_groupi_g14561(csa_tree_add_6_33_groupi_n_3730 ,csa_tree_add_6_33_groupi_n_3544 ,csa_tree_add_6_33_groupi_n_3432);
  or csa_tree_add_6_33_groupi_g14562(csa_tree_add_6_33_groupi_n_3729 ,csa_tree_add_6_33_groupi_n_3047 ,csa_tree_add_6_33_groupi_n_3526);
  and csa_tree_add_6_33_groupi_g14563(csa_tree_add_6_33_groupi_n_3728 ,csa_tree_add_6_33_groupi_n_3495 ,csa_tree_add_6_33_groupi_n_3485);
  and csa_tree_add_6_33_groupi_g14564(csa_tree_add_6_33_groupi_n_3727 ,csa_tree_add_6_33_groupi_n_2676 ,csa_tree_add_6_33_groupi_n_3471);
  or csa_tree_add_6_33_groupi_g14565(csa_tree_add_6_33_groupi_n_3726 ,csa_tree_add_6_33_groupi_n_3545 ,csa_tree_add_6_33_groupi_n_3460);
  nor csa_tree_add_6_33_groupi_g14566(csa_tree_add_6_33_groupi_n_3725 ,csa_tree_add_6_33_groupi_n_2676 ,csa_tree_add_6_33_groupi_n_3471);
  nor csa_tree_add_6_33_groupi_g14567(csa_tree_add_6_33_groupi_n_3724 ,csa_tree_add_6_33_groupi_n_2995 ,csa_tree_add_6_33_groupi_n_3480);
  and csa_tree_add_6_33_groupi_g14568(csa_tree_add_6_33_groupi_n_3723 ,csa_tree_add_6_33_groupi_n_3545 ,csa_tree_add_6_33_groupi_n_3460);
  nor csa_tree_add_6_33_groupi_g14569(csa_tree_add_6_33_groupi_n_3722 ,csa_tree_add_6_33_groupi_n_3345 ,csa_tree_add_6_33_groupi_n_3442);
  and csa_tree_add_6_33_groupi_g14570(csa_tree_add_6_33_groupi_n_3721 ,csa_tree_add_6_33_groupi_n_3047 ,csa_tree_add_6_33_groupi_n_3526);
  or csa_tree_add_6_33_groupi_g14571(csa_tree_add_6_33_groupi_n_3720 ,csa_tree_add_6_33_groupi_n_2682 ,csa_tree_add_6_33_groupi_n_3445);
  or csa_tree_add_6_33_groupi_g14572(csa_tree_add_6_33_groupi_n_3719 ,csa_tree_add_6_33_groupi_n_3534 ,csa_tree_add_6_33_groupi_n_3421);
  and csa_tree_add_6_33_groupi_g14573(csa_tree_add_6_33_groupi_n_3718 ,csa_tree_add_6_33_groupi_n_3269 ,csa_tree_add_6_33_groupi_n_3447);
  and csa_tree_add_6_33_groupi_g14574(csa_tree_add_6_33_groupi_n_3717 ,csa_tree_add_6_33_groupi_n_3419 ,csa_tree_add_6_33_groupi_n_3418);
  and csa_tree_add_6_33_groupi_g14575(csa_tree_add_6_33_groupi_n_3716 ,csa_tree_add_6_33_groupi_n_3371 ,csa_tree_add_6_33_groupi_n_3441);
  or csa_tree_add_6_33_groupi_g14576(csa_tree_add_6_33_groupi_n_3715 ,csa_tree_add_6_33_groupi_n_3371 ,csa_tree_add_6_33_groupi_n_3441);
  or csa_tree_add_6_33_groupi_g14577(csa_tree_add_6_33_groupi_n_3714 ,csa_tree_add_6_33_groupi_n_3463 ,csa_tree_add_6_33_groupi_n_3461);
  and csa_tree_add_6_33_groupi_g14578(csa_tree_add_6_33_groupi_n_3713 ,csa_tree_add_6_33_groupi_n_3186 ,csa_tree_add_6_33_groupi_n_3468);
  or csa_tree_add_6_33_groupi_g14579(csa_tree_add_6_33_groupi_n_3712 ,csa_tree_add_6_33_groupi_n_3344 ,csa_tree_add_6_33_groupi_n_3443);
  or csa_tree_add_6_33_groupi_g14580(csa_tree_add_6_33_groupi_n_3711 ,csa_tree_add_6_33_groupi_n_3419 ,csa_tree_add_6_33_groupi_n_3418);
  and csa_tree_add_6_33_groupi_g14581(csa_tree_add_6_33_groupi_n_3710 ,csa_tree_add_6_33_groupi_n_3534 ,csa_tree_add_6_33_groupi_n_3421);
  or csa_tree_add_6_33_groupi_g14582(csa_tree_add_6_33_groupi_n_3709 ,csa_tree_add_6_33_groupi_n_2659 ,csa_tree_add_6_33_groupi_n_3438);
  or csa_tree_add_6_33_groupi_g14583(csa_tree_add_6_33_groupi_n_3708 ,csa_tree_add_6_33_groupi_n_3490 ,csa_tree_add_6_33_groupi_n_3570);
  or csa_tree_add_6_33_groupi_g14584(csa_tree_add_6_33_groupi_n_3707 ,csa_tree_add_6_33_groupi_n_3048 ,csa_tree_add_6_33_groupi_n_3532);
  and csa_tree_add_6_33_groupi_g14585(csa_tree_add_6_33_groupi_n_3706 ,csa_tree_add_6_33_groupi_n_3346 ,csa_tree_add_6_33_groupi_n_3529);
  or csa_tree_add_6_33_groupi_g14586(csa_tree_add_6_33_groupi_n_3705 ,csa_tree_add_6_33_groupi_n_3367 ,csa_tree_add_6_33_groupi_n_3437);
  and csa_tree_add_6_33_groupi_g14587(csa_tree_add_6_33_groupi_n_3704 ,csa_tree_add_6_33_groupi_n_3367 ,csa_tree_add_6_33_groupi_n_3437);
  or csa_tree_add_6_33_groupi_g14588(csa_tree_add_6_33_groupi_n_3703 ,csa_tree_add_6_33_groupi_n_3467 ,csa_tree_add_6_33_groupi_n_3436);
  or csa_tree_add_6_33_groupi_g14589(csa_tree_add_6_33_groupi_n_3702 ,csa_tree_add_6_33_groupi_n_3307 ,csa_tree_add_6_33_groupi_n_3567);
  and csa_tree_add_6_33_groupi_g14590(csa_tree_add_6_33_groupi_n_3701 ,csa_tree_add_6_33_groupi_n_2659 ,csa_tree_add_6_33_groupi_n_3438);
  and csa_tree_add_6_33_groupi_g14591(csa_tree_add_6_33_groupi_n_3700 ,csa_tree_add_6_33_groupi_n_3467 ,csa_tree_add_6_33_groupi_n_3436);
  or csa_tree_add_6_33_groupi_g14592(csa_tree_add_6_33_groupi_n_3699 ,csa_tree_add_6_33_groupi_n_3366 ,csa_tree_add_6_33_groupi_n_3431);
  or csa_tree_add_6_33_groupi_g14593(csa_tree_add_6_33_groupi_n_3698 ,csa_tree_add_6_33_groupi_n_3382 ,csa_tree_add_6_33_groupi_n_3499);
  or csa_tree_add_6_33_groupi_g14594(csa_tree_add_6_33_groupi_n_3697 ,csa_tree_add_6_33_groupi_n_3422 ,csa_tree_add_6_33_groupi_n_3430);
  and csa_tree_add_6_33_groupi_g14595(csa_tree_add_6_33_groupi_n_3696 ,csa_tree_add_6_33_groupi_n_3366 ,csa_tree_add_6_33_groupi_n_3431);
  nor csa_tree_add_6_33_groupi_g14596(csa_tree_add_6_33_groupi_n_3695 ,csa_tree_add_6_33_groupi_n_3423 ,csa_tree_add_6_33_groupi_n_3429);
  or csa_tree_add_6_33_groupi_g14597(csa_tree_add_6_33_groupi_n_3694 ,csa_tree_add_6_33_groupi_n_3364 ,csa_tree_add_6_33_groupi_n_3428);
  and csa_tree_add_6_33_groupi_g14598(csa_tree_add_6_33_groupi_n_3693 ,csa_tree_add_6_33_groupi_n_2682 ,csa_tree_add_6_33_groupi_n_3445);
  or csa_tree_add_6_33_groupi_g14599(csa_tree_add_6_33_groupi_n_3692 ,csa_tree_add_6_33_groupi_n_3377 ,csa_tree_add_6_33_groupi_n_3502);
  or csa_tree_add_6_33_groupi_g14600(csa_tree_add_6_33_groupi_n_3691 ,csa_tree_add_6_33_groupi_n_3189 ,csa_tree_add_6_33_groupi_n_3426);
  or csa_tree_add_6_33_groupi_g14601(csa_tree_add_6_33_groupi_n_3690 ,csa_tree_add_6_33_groupi_n_3346 ,csa_tree_add_6_33_groupi_n_3529);
  and csa_tree_add_6_33_groupi_g14602(csa_tree_add_6_33_groupi_n_3689 ,csa_tree_add_6_33_groupi_n_3364 ,csa_tree_add_6_33_groupi_n_3428);
  or csa_tree_add_6_33_groupi_g14603(csa_tree_add_6_33_groupi_n_3688 ,csa_tree_add_6_33_groupi_n_3425 ,csa_tree_add_6_33_groupi_n_3424);
  or csa_tree_add_6_33_groupi_g14604(csa_tree_add_6_33_groupi_n_3687 ,csa_tree_add_6_33_groupi_n_3278 ,csa_tree_add_6_33_groupi_n_3420);
  and csa_tree_add_6_33_groupi_g14605(csa_tree_add_6_33_groupi_n_3686 ,csa_tree_add_6_33_groupi_n_3425 ,csa_tree_add_6_33_groupi_n_3424);
  and csa_tree_add_6_33_groupi_g14606(csa_tree_add_6_33_groupi_n_3685 ,csa_tree_add_6_33_groupi_n_3189 ,csa_tree_add_6_33_groupi_n_3426);
  and csa_tree_add_6_33_groupi_g14607(csa_tree_add_6_33_groupi_n_3684 ,csa_tree_add_6_33_groupi_n_3278 ,csa_tree_add_6_33_groupi_n_3420);
  or csa_tree_add_6_33_groupi_g14608(csa_tree_add_6_33_groupi_n_3683 ,csa_tree_add_6_33_groupi_n_3519 ,csa_tree_add_6_33_groupi_n_3550);
  and csa_tree_add_6_33_groupi_g14609(csa_tree_add_6_33_groupi_n_3772 ,csa_tree_add_6_33_groupi_n_3025 ,csa_tree_add_6_33_groupi_n_3510);
  and csa_tree_add_6_33_groupi_g14610(csa_tree_add_6_33_groupi_n_3771 ,csa_tree_add_6_33_groupi_n_3339 ,csa_tree_add_6_33_groupi_n_3494);
  and csa_tree_add_6_33_groupi_g14611(csa_tree_add_6_33_groupi_n_3770 ,csa_tree_add_6_33_groupi_n_3303 ,csa_tree_add_6_33_groupi_n_3491);
  and csa_tree_add_6_33_groupi_g14612(csa_tree_add_6_33_groupi_n_3769 ,csa_tree_add_6_33_groupi_n_3098 ,csa_tree_add_6_33_groupi_n_3515);
  and csa_tree_add_6_33_groupi_g14613(csa_tree_add_6_33_groupi_n_3768 ,csa_tree_add_6_33_groupi_n_3064 ,csa_tree_add_6_33_groupi_n_3521);
  and csa_tree_add_6_33_groupi_g14614(csa_tree_add_6_33_groupi_n_3767 ,csa_tree_add_6_33_groupi_n_2983 ,csa_tree_add_6_33_groupi_n_3497);
  and csa_tree_add_6_33_groupi_g14615(csa_tree_add_6_33_groupi_n_3766 ,csa_tree_add_6_33_groupi_n_3170 ,csa_tree_add_6_33_groupi_n_3517);
  and csa_tree_add_6_33_groupi_g14616(csa_tree_add_6_33_groupi_n_3765 ,csa_tree_add_6_33_groupi_n_3007 ,csa_tree_add_6_33_groupi_n_3402);
  and csa_tree_add_6_33_groupi_g14617(csa_tree_add_6_33_groupi_n_3764 ,csa_tree_add_6_33_groupi_n_3258 ,csa_tree_add_6_33_groupi_n_3405);
  and csa_tree_add_6_33_groupi_g14618(csa_tree_add_6_33_groupi_n_3763 ,csa_tree_add_6_33_groupi_n_3325 ,csa_tree_add_6_33_groupi_n_3506);
  and csa_tree_add_6_33_groupi_g14619(csa_tree_add_6_33_groupi_n_3762 ,csa_tree_add_6_33_groupi_n_3166 ,csa_tree_add_6_33_groupi_n_3514);
  and csa_tree_add_6_33_groupi_g14620(csa_tree_add_6_33_groupi_n_3761 ,csa_tree_add_6_33_groupi_n_3143 ,csa_tree_add_6_33_groupi_n_3501);
  and csa_tree_add_6_33_groupi_g14621(csa_tree_add_6_33_groupi_n_3760 ,csa_tree_add_6_33_groupi_n_3102 ,csa_tree_add_6_33_groupi_n_3498);
  not csa_tree_add_6_33_groupi_g14622(csa_tree_add_6_33_groupi_n_3682 ,csa_tree_add_6_33_groupi_n_3681);
  not csa_tree_add_6_33_groupi_g14623(csa_tree_add_6_33_groupi_n_3670 ,csa_tree_add_6_33_groupi_n_3671);
  not csa_tree_add_6_33_groupi_g14624(csa_tree_add_6_33_groupi_n_3667 ,csa_tree_add_6_33_groupi_n_3668);
  not csa_tree_add_6_33_groupi_g14625(csa_tree_add_6_33_groupi_n_3664 ,csa_tree_add_6_33_groupi_n_3665);
  not csa_tree_add_6_33_groupi_g14626(csa_tree_add_6_33_groupi_n_3659 ,csa_tree_add_6_33_groupi_n_3660);
  not csa_tree_add_6_33_groupi_g14627(csa_tree_add_6_33_groupi_n_3655 ,csa_tree_add_6_33_groupi_n_3654);
  not csa_tree_add_6_33_groupi_g14628(csa_tree_add_6_33_groupi_n_3650 ,csa_tree_add_6_33_groupi_n_3651);
  not csa_tree_add_6_33_groupi_g14629(csa_tree_add_6_33_groupi_n_3646 ,csa_tree_add_6_33_groupi_n_3647);
  not csa_tree_add_6_33_groupi_g14630(csa_tree_add_6_33_groupi_n_3644 ,csa_tree_add_6_33_groupi_n_3645);
  not csa_tree_add_6_33_groupi_g14631(csa_tree_add_6_33_groupi_n_3638 ,csa_tree_add_6_33_groupi_n_3639);
  not csa_tree_add_6_33_groupi_g14632(csa_tree_add_6_33_groupi_n_3633 ,csa_tree_add_6_33_groupi_n_3634);
  not csa_tree_add_6_33_groupi_g14633(csa_tree_add_6_33_groupi_n_3630 ,csa_tree_add_6_33_groupi_n_3631);
  not csa_tree_add_6_33_groupi_g14634(csa_tree_add_6_33_groupi_n_3628 ,csa_tree_add_6_33_groupi_n_3629);
  not csa_tree_add_6_33_groupi_g14635(csa_tree_add_6_33_groupi_n_3625 ,csa_tree_add_6_33_groupi_n_3626);
  not csa_tree_add_6_33_groupi_g14636(csa_tree_add_6_33_groupi_n_3621 ,csa_tree_add_6_33_groupi_n_3622);
  not csa_tree_add_6_33_groupi_g14637(csa_tree_add_6_33_groupi_n_3618 ,csa_tree_add_6_33_groupi_n_3619);
  not csa_tree_add_6_33_groupi_g14638(csa_tree_add_6_33_groupi_n_3615 ,csa_tree_add_6_33_groupi_n_3616);
  not csa_tree_add_6_33_groupi_g14639(csa_tree_add_6_33_groupi_n_3613 ,csa_tree_add_6_33_groupi_n_3614);
  not csa_tree_add_6_33_groupi_g14640(csa_tree_add_6_33_groupi_n_3612 ,csa_tree_add_6_33_groupi_n_3611);
  not csa_tree_add_6_33_groupi_g14641(csa_tree_add_6_33_groupi_n_3609 ,csa_tree_add_6_33_groupi_n_3610);
  not csa_tree_add_6_33_groupi_g14642(csa_tree_add_6_33_groupi_n_3607 ,csa_tree_add_6_33_groupi_n_3608);
  or csa_tree_add_6_33_groupi_g14643(csa_tree_add_6_33_groupi_n_3605 ,csa_tree_add_6_33_groupi_n_2902 ,csa_tree_add_6_33_groupi_n_3474);
  and csa_tree_add_6_33_groupi_g14644(csa_tree_add_6_33_groupi_n_3604 ,csa_tree_add_6_33_groupi_n_3527 ,csa_tree_add_6_33_groupi_n_3449);
  or csa_tree_add_6_33_groupi_g14645(csa_tree_add_6_33_groupi_n_3603 ,csa_tree_add_6_33_groupi_n_3279 ,csa_tree_add_6_33_groupi_n_3412);
  or csa_tree_add_6_33_groupi_g14646(csa_tree_add_6_33_groupi_n_3602 ,csa_tree_add_6_33_groupi_n_3464 ,csa_tree_add_6_33_groupi_n_3411);
  and csa_tree_add_6_33_groupi_g14647(csa_tree_add_6_33_groupi_n_3601 ,csa_tree_add_6_33_groupi_n_3370 ,csa_tree_add_6_33_groupi_n_3469);
  or csa_tree_add_6_33_groupi_g14648(csa_tree_add_6_33_groupi_n_3600 ,csa_tree_add_6_33_groupi_n_3370 ,csa_tree_add_6_33_groupi_n_3469);
  or csa_tree_add_6_33_groupi_g14649(csa_tree_add_6_33_groupi_n_3599 ,csa_tree_add_6_33_groupi_n_3285 ,csa_tree_add_6_33_groupi_n_3400);
  nor csa_tree_add_6_33_groupi_g14650(csa_tree_add_6_33_groupi_n_3598 ,csa_tree_add_6_33_groupi_n_2903 ,csa_tree_add_6_33_groupi_n_3475);
  or csa_tree_add_6_33_groupi_g14651(csa_tree_add_6_33_groupi_n_3597 ,csa_tree_add_6_33_groupi_n_3270 ,csa_tree_add_6_33_groupi_n_3470);
  and csa_tree_add_6_33_groupi_g14652(csa_tree_add_6_33_groupi_n_3596 ,csa_tree_add_6_33_groupi_n_3270 ,csa_tree_add_6_33_groupi_n_3470);
  xnor csa_tree_add_6_33_groupi_g14653(out1[3] ,csa_tree_add_6_33_groupi_n_3282 ,csa_tree_add_6_33_groupi_n_2968);
  and csa_tree_add_6_33_groupi_g14654(csa_tree_add_6_33_groupi_n_3594 ,csa_tree_add_6_33_groupi_n_3044 ,csa_tree_add_6_33_groupi_n_3417);
  xnor csa_tree_add_6_33_groupi_g14655(csa_tree_add_6_33_groupi_n_3593 ,csa_tree_add_6_33_groupi_n_3290 ,csa_tree_add_6_33_groupi_n_3042);
  xnor csa_tree_add_6_33_groupi_g14656(csa_tree_add_6_33_groupi_n_3592 ,csa_tree_add_6_33_groupi_n_3046 ,csa_tree_add_6_33_groupi_n_3285);
  xnor csa_tree_add_6_33_groupi_g14657(csa_tree_add_6_33_groupi_n_3591 ,csa_tree_add_6_33_groupi_n_3289 ,csa_tree_add_6_33_groupi_n_3044);
  xnor csa_tree_add_6_33_groupi_g14658(csa_tree_add_6_33_groupi_n_3590 ,csa_tree_add_6_33_groupi_n_3347 ,csa_tree_add_6_33_groupi_n_2621);
  xnor csa_tree_add_6_33_groupi_g14659(csa_tree_add_6_33_groupi_n_3589 ,csa_tree_add_6_33_groupi_n_3387 ,csa_tree_add_6_33_groupi_n_2659);
  xnor csa_tree_add_6_33_groupi_g14660(csa_tree_add_6_33_groupi_n_3588 ,csa_tree_add_6_33_groupi_n_3377 ,csa_tree_add_6_33_groupi_n_2632);
  xnor csa_tree_add_6_33_groupi_g14661(csa_tree_add_6_33_groupi_n_3587 ,csa_tree_add_6_33_groupi_n_3047 ,csa_tree_add_6_33_groupi_n_3386);
  xnor csa_tree_add_6_33_groupi_g14662(csa_tree_add_6_33_groupi_n_3586 ,csa_tree_add_6_33_groupi_n_3378 ,csa_tree_add_6_33_groupi_n_2609);
  xnor csa_tree_add_6_33_groupi_g14663(csa_tree_add_6_33_groupi_n_3585 ,csa_tree_add_6_33_groupi_n_3279 ,csa_tree_add_6_33_groupi_n_3281);
  xnor csa_tree_add_6_33_groupi_g14664(csa_tree_add_6_33_groupi_n_3584 ,csa_tree_add_6_33_groupi_n_3355 ,csa_tree_add_6_33_groupi_n_3268);
  xnor csa_tree_add_6_33_groupi_g14665(csa_tree_add_6_33_groupi_n_3583 ,csa_tree_add_6_33_groupi_n_3050 ,csa_tree_add_6_33_groupi_n_3348);
  xnor csa_tree_add_6_33_groupi_g14666(csa_tree_add_6_33_groupi_n_3582 ,csa_tree_add_6_33_groupi_n_3052 ,csa_tree_add_6_33_groupi_n_3350);
  xnor csa_tree_add_6_33_groupi_g14667(csa_tree_add_6_33_groupi_n_3581 ,csa_tree_add_6_33_groupi_n_3291 ,csa_tree_add_6_33_groupi_n_3346);
  xnor csa_tree_add_6_33_groupi_g14668(csa_tree_add_6_33_groupi_n_3580 ,csa_tree_add_6_33_groupi_n_3357 ,csa_tree_add_6_33_groupi_n_2890);
  xnor csa_tree_add_6_33_groupi_g14669(csa_tree_add_6_33_groupi_n_3579 ,csa_tree_add_6_33_groupi_n_3185 ,csa_tree_add_6_33_groupi_n_3271);
  xor csa_tree_add_6_33_groupi_g14670(csa_tree_add_6_33_groupi_n_3578 ,csa_tree_add_6_33_groupi_n_2676 ,csa_tree_add_6_33_groupi_n_3284);
  xnor csa_tree_add_6_33_groupi_g14671(csa_tree_add_6_33_groupi_n_3577 ,csa_tree_add_6_33_groupi_n_3359 ,csa_tree_add_6_33_groupi_n_2681);
  xnor csa_tree_add_6_33_groupi_g14672(csa_tree_add_6_33_groupi_n_3576 ,csa_tree_add_6_33_groupi_n_2903 ,csa_tree_add_6_33_groupi_n_3380);
  xnor csa_tree_add_6_33_groupi_g14673(csa_tree_add_6_33_groupi_n_3575 ,csa_tree_add_6_33_groupi_n_3362 ,csa_tree_add_6_33_groupi_n_2692);
  xnor csa_tree_add_6_33_groupi_g14674(csa_tree_add_6_33_groupi_n_3574 ,csa_tree_add_6_33_groupi_n_2897 ,csa_tree_add_6_33_groupi_n_3353);
  xnor csa_tree_add_6_33_groupi_g14675(csa_tree_add_6_33_groupi_n_3573 ,csa_tree_add_6_33_groupi_n_2614 ,csa_tree_add_6_33_groupi_n_3361);
  xnor csa_tree_add_6_33_groupi_g14676(csa_tree_add_6_33_groupi_n_3681 ,csa_tree_add_6_33_groupi_n_2724 ,csa_tree_add_6_33_groupi_n_3248);
  xnor csa_tree_add_6_33_groupi_g14677(csa_tree_add_6_33_groupi_n_3680 ,csa_tree_add_6_33_groupi_n_3375 ,csa_tree_add_6_33_groupi_n_3214);
  xnor csa_tree_add_6_33_groupi_g14678(csa_tree_add_6_33_groupi_n_3679 ,csa_tree_add_6_33_groupi_n_3057 ,csa_tree_add_6_33_groupi_n_3207);
  xnor csa_tree_add_6_33_groupi_g14679(csa_tree_add_6_33_groupi_n_3678 ,csa_tree_add_6_33_groupi_n_3376 ,csa_tree_add_6_33_groupi_n_3204);
  xnor csa_tree_add_6_33_groupi_g14680(csa_tree_add_6_33_groupi_n_3677 ,csa_tree_add_6_33_groupi_n_2685 ,csa_tree_add_6_33_groupi_n_3244);
  xnor csa_tree_add_6_33_groupi_g14681(csa_tree_add_6_33_groupi_n_3676 ,csa_tree_add_6_33_groupi_n_3192 ,csa_tree_add_6_33_groupi_n_3213);
  xnor csa_tree_add_6_33_groupi_g14682(csa_tree_add_6_33_groupi_n_3675 ,csa_tree_add_6_33_groupi_n_3381 ,csa_tree_add_6_33_groupi_n_3230);
  xnor csa_tree_add_6_33_groupi_g14683(csa_tree_add_6_33_groupi_n_3674 ,csa_tree_add_6_33_groupi_n_2684 ,csa_tree_add_6_33_groupi_n_3236);
  xnor csa_tree_add_6_33_groupi_g14684(csa_tree_add_6_33_groupi_n_3673 ,csa_tree_add_6_33_groupi_n_3287 ,csa_tree_add_6_33_groupi_n_3220);
  or csa_tree_add_6_33_groupi_g14685(csa_tree_add_6_33_groupi_n_3672 ,csa_tree_add_6_33_groupi_n_2830 ,csa_tree_add_6_33_groupi_n_3399);
  xnor csa_tree_add_6_33_groupi_g14686(csa_tree_add_6_33_groupi_n_3671 ,csa_tree_add_6_33_groupi_n_3389 ,csa_tree_add_6_33_groupi_n_3227);
  xnor csa_tree_add_6_33_groupi_g14687(csa_tree_add_6_33_groupi_n_3669 ,csa_tree_add_6_33_groupi_n_2597 ,csa_tree_add_6_33_groupi_n_3212);
  xnor csa_tree_add_6_33_groupi_g14688(csa_tree_add_6_33_groupi_n_3668 ,csa_tree_add_6_33_groupi_n_2735 ,csa_tree_add_6_33_groupi_n_3223);
  xnor csa_tree_add_6_33_groupi_g14689(csa_tree_add_6_33_groupi_n_3666 ,csa_tree_add_6_33_groupi_n_2606 ,csa_tree_add_6_33_groupi_n_3210);
  xnor csa_tree_add_6_33_groupi_g14690(csa_tree_add_6_33_groupi_n_3665 ,csa_tree_add_6_33_groupi_n_3292 ,csa_tree_add_6_33_groupi_n_3211);
  xnor csa_tree_add_6_33_groupi_g14691(csa_tree_add_6_33_groupi_n_3663 ,csa_tree_add_6_33_groupi_n_3390 ,csa_tree_add_6_33_groupi_n_3231);
  xnor csa_tree_add_6_33_groupi_g14692(csa_tree_add_6_33_groupi_n_3662 ,csa_tree_add_6_33_groupi_n_2599 ,csa_tree_add_6_33_groupi_n_3208);
  xnor csa_tree_add_6_33_groupi_g14693(csa_tree_add_6_33_groupi_n_3661 ,csa_tree_add_6_33_groupi_n_2649 ,csa_tree_add_6_33_groupi_n_3206);
  xnor csa_tree_add_6_33_groupi_g14694(csa_tree_add_6_33_groupi_n_3660 ,csa_tree_add_6_33_groupi_n_2715 ,csa_tree_add_6_33_groupi_n_3240);
  xnor csa_tree_add_6_33_groupi_g14695(csa_tree_add_6_33_groupi_n_3658 ,csa_tree_add_6_33_groupi_n_2620 ,csa_tree_add_6_33_groupi_n_3205);
  xnor csa_tree_add_6_33_groupi_g14696(csa_tree_add_6_33_groupi_n_3657 ,csa_tree_add_6_33_groupi_n_3379 ,csa_tree_add_6_33_groupi_n_3217);
  xnor csa_tree_add_6_33_groupi_g14697(csa_tree_add_6_33_groupi_n_3656 ,csa_tree_add_6_33_groupi_n_3280 ,csa_tree_add_6_33_groupi_n_3203);
  xnor csa_tree_add_6_33_groupi_g14698(csa_tree_add_6_33_groupi_n_3654 ,csa_tree_add_6_33_groupi_n_3059 ,csa_tree_add_6_33_groupi_n_3202);
  xnor csa_tree_add_6_33_groupi_g14699(csa_tree_add_6_33_groupi_n_3653 ,csa_tree_add_6_33_groupi_n_3374 ,csa_tree_add_6_33_groupi_n_3201);
  xnor csa_tree_add_6_33_groupi_g14700(csa_tree_add_6_33_groupi_n_3652 ,csa_tree_add_6_33_groupi_n_2716 ,csa_tree_add_6_33_groupi_n_3200);
  xnor csa_tree_add_6_33_groupi_g14701(csa_tree_add_6_33_groupi_n_3651 ,csa_tree_add_6_33_groupi_n_2736 ,csa_tree_add_6_33_groupi_n_3218);
  xnor csa_tree_add_6_33_groupi_g14702(csa_tree_add_6_33_groupi_n_3649 ,csa_tree_add_6_33_groupi_n_3193 ,csa_tree_add_6_33_groupi_n_3196);
  xnor csa_tree_add_6_33_groupi_g14703(csa_tree_add_6_33_groupi_n_3648 ,csa_tree_add_6_33_groupi_n_2751 ,csa_tree_add_6_33_groupi_n_3197);
  xnor csa_tree_add_6_33_groupi_g14704(csa_tree_add_6_33_groupi_n_3647 ,csa_tree_add_6_33_groupi_n_2619 ,csa_tree_add_6_33_groupi_n_3219);
  xnor csa_tree_add_6_33_groupi_g14705(csa_tree_add_6_33_groupi_n_3645 ,csa_tree_add_6_33_groupi_n_2675 ,csa_tree_add_6_33_groupi_n_3224);
  xnor csa_tree_add_6_33_groupi_g14706(csa_tree_add_6_33_groupi_n_3643 ,csa_tree_add_6_33_groupi_n_2753 ,csa_tree_add_6_33_groupi_n_3229);
  xnor csa_tree_add_6_33_groupi_g14707(csa_tree_add_6_33_groupi_n_3642 ,csa_tree_add_6_33_groupi_n_2708 ,csa_tree_add_6_33_groupi_n_3237);
  and csa_tree_add_6_33_groupi_g14708(csa_tree_add_6_33_groupi_n_3641 ,csa_tree_add_6_33_groupi_n_3264 ,csa_tree_add_6_33_groupi_n_3512);
  xnor csa_tree_add_6_33_groupi_g14709(csa_tree_add_6_33_groupi_n_3640 ,csa_tree_add_6_33_groupi_n_2744 ,csa_tree_add_6_33_groupi_n_3232);
  xnor csa_tree_add_6_33_groupi_g14710(csa_tree_add_6_33_groupi_n_3639 ,csa_tree_add_6_33_groupi_n_2749 ,csa_tree_add_6_33_groupi_n_3226);
  xnor csa_tree_add_6_33_groupi_g14711(csa_tree_add_6_33_groupi_n_3637 ,csa_tree_add_6_33_groupi_n_2742 ,csa_tree_add_6_33_groupi_n_3234);
  xnor csa_tree_add_6_33_groupi_g14712(csa_tree_add_6_33_groupi_n_3636 ,csa_tree_add_6_33_groupi_n_3195 ,csa_tree_add_6_33_groupi_n_3235);
  xnor csa_tree_add_6_33_groupi_g14713(csa_tree_add_6_33_groupi_n_3635 ,csa_tree_add_6_33_groupi_n_3194 ,csa_tree_add_6_33_groupi_n_3238);
  xnor csa_tree_add_6_33_groupi_g14714(csa_tree_add_6_33_groupi_n_3634 ,csa_tree_add_6_33_groupi_n_2740 ,csa_tree_add_6_33_groupi_n_3225);
  xnor csa_tree_add_6_33_groupi_g14715(csa_tree_add_6_33_groupi_n_3632 ,csa_tree_add_6_33_groupi_n_2755 ,csa_tree_add_6_33_groupi_n_3239);
  xnor csa_tree_add_6_33_groupi_g14716(csa_tree_add_6_33_groupi_n_3631 ,csa_tree_add_6_33_groupi_n_3191 ,csa_tree_add_6_33_groupi_n_3228);
  xnor csa_tree_add_6_33_groupi_g14717(csa_tree_add_6_33_groupi_n_3629 ,csa_tree_add_6_33_groupi_n_2733 ,csa_tree_add_6_33_groupi_n_3242);
  xnor csa_tree_add_6_33_groupi_g14718(csa_tree_add_6_33_groupi_n_3627 ,csa_tree_add_6_33_groupi_n_2647 ,csa_tree_add_6_33_groupi_n_3247);
  xnor csa_tree_add_6_33_groupi_g14719(csa_tree_add_6_33_groupi_n_3626 ,csa_tree_add_6_33_groupi_n_2658 ,csa_tree_add_6_33_groupi_n_3221);
  xnor csa_tree_add_6_33_groupi_g14720(csa_tree_add_6_33_groupi_n_3624 ,csa_tree_add_6_33_groupi_n_2629 ,csa_tree_add_6_33_groupi_n_3241);
  xnor csa_tree_add_6_33_groupi_g14721(csa_tree_add_6_33_groupi_n_3623 ,csa_tree_add_6_33_groupi_n_2639 ,csa_tree_add_6_33_groupi_n_3246);
  xnor csa_tree_add_6_33_groupi_g14722(csa_tree_add_6_33_groupi_n_3622 ,csa_tree_add_6_33_groupi_n_2913 ,csa_tree_add_6_33_groupi_n_3198);
  xnor csa_tree_add_6_33_groupi_g14723(csa_tree_add_6_33_groupi_n_3620 ,csa_tree_add_6_33_groupi_n_2617 ,csa_tree_add_6_33_groupi_n_3243);
  xnor csa_tree_add_6_33_groupi_g14724(csa_tree_add_6_33_groupi_n_3619 ,csa_tree_add_6_33_groupi_n_2623 ,csa_tree_add_6_33_groupi_n_3249);
  xnor csa_tree_add_6_33_groupi_g14725(csa_tree_add_6_33_groupi_n_3617 ,csa_tree_add_6_33_groupi_n_2607 ,csa_tree_add_6_33_groupi_n_3245);
  xnor csa_tree_add_6_33_groupi_g14726(csa_tree_add_6_33_groupi_n_3616 ,csa_tree_add_6_33_groupi_n_2644 ,csa_tree_add_6_33_groupi_n_3222);
  or csa_tree_add_6_33_groupi_g14727(csa_tree_add_6_33_groupi_n_3614 ,csa_tree_add_6_33_groupi_n_3135 ,csa_tree_add_6_33_groupi_n_3403);
  xnor csa_tree_add_6_33_groupi_g14728(csa_tree_add_6_33_groupi_n_3611 ,csa_tree_add_6_33_groupi_n_2915 ,csa_tree_add_6_33_groupi_n_3199);
  xnor csa_tree_add_6_33_groupi_g14729(csa_tree_add_6_33_groupi_n_3610 ,csa_tree_add_6_33_groupi_n_3058 ,csa_tree_add_6_33_groupi_n_3209);
  and csa_tree_add_6_33_groupi_g14730(csa_tree_add_6_33_groupi_n_3608 ,csa_tree_add_6_33_groupi_n_2990 ,csa_tree_add_6_33_groupi_n_3398);
  xnor csa_tree_add_6_33_groupi_g14731(csa_tree_add_6_33_groupi_n_3606 ,csa_tree_add_6_33_groupi_n_3383 ,csa_tree_add_6_33_groupi_n_3215);
  not csa_tree_add_6_33_groupi_g14732(csa_tree_add_6_33_groupi_n_3543 ,csa_tree_add_6_33_groupi_n_3544);
  not csa_tree_add_6_33_groupi_g14733(csa_tree_add_6_33_groupi_n_3541 ,csa_tree_add_6_33_groupi_n_3540);
  not csa_tree_add_6_33_groupi_g14734(csa_tree_add_6_33_groupi_n_3538 ,csa_tree_add_6_33_groupi_n_3539);
  not csa_tree_add_6_33_groupi_g14735(csa_tree_add_6_33_groupi_n_3530 ,csa_tree_add_6_33_groupi_n_3531);
  not csa_tree_add_6_33_groupi_g14736(csa_tree_add_6_33_groupi_n_3524 ,csa_tree_add_6_33_groupi_n_3525);
  not csa_tree_add_6_33_groupi_g14737(csa_tree_add_6_33_groupi_n_3522 ,csa_tree_add_6_33_groupi_n_3523);
  or csa_tree_add_6_33_groupi_g14738(csa_tree_add_6_33_groupi_n_3521 ,csa_tree_add_6_33_groupi_n_3008 ,csa_tree_add_6_33_groupi_n_3381);
  and csa_tree_add_6_33_groupi_g14739(csa_tree_add_6_33_groupi_n_3520 ,csa_tree_add_6_33_groupi_n_3348 ,csa_tree_add_6_33_groupi_n_3050);
  and csa_tree_add_6_33_groupi_g14740(csa_tree_add_6_33_groupi_n_3519 ,csa_tree_add_6_33_groupi_n_2621 ,csa_tree_add_6_33_groupi_n_3347);
  and csa_tree_add_6_33_groupi_g14741(csa_tree_add_6_33_groupi_n_3518 ,csa_tree_add_6_33_groupi_n_2897 ,csa_tree_add_6_33_groupi_n_3353);
  or csa_tree_add_6_33_groupi_g14742(csa_tree_add_6_33_groupi_n_3517 ,csa_tree_add_6_33_groupi_n_3168 ,csa_tree_add_6_33_groupi_n_3374);
  nor csa_tree_add_6_33_groupi_g14743(csa_tree_add_6_33_groupi_n_3516 ,csa_tree_add_6_33_groupi_n_2897 ,csa_tree_add_6_33_groupi_n_3353);
  or csa_tree_add_6_33_groupi_g14744(csa_tree_add_6_33_groupi_n_3515 ,csa_tree_add_6_33_groupi_n_3091 ,csa_tree_add_6_33_groupi_n_3389);
  or csa_tree_add_6_33_groupi_g14745(csa_tree_add_6_33_groupi_n_3514 ,csa_tree_add_6_33_groupi_n_3164 ,csa_tree_add_6_33_groupi_n_3376);
  or csa_tree_add_6_33_groupi_g14746(csa_tree_add_6_33_groupi_n_3513 ,csa_tree_add_6_33_groupi_n_2614 ,csa_tree_add_6_33_groupi_n_3360);
  or csa_tree_add_6_33_groupi_g14747(csa_tree_add_6_33_groupi_n_3512 ,csa_tree_add_6_33_groupi_n_3372 ,csa_tree_add_6_33_groupi_n_3311);
  nor csa_tree_add_6_33_groupi_g14748(csa_tree_add_6_33_groupi_n_3511 ,csa_tree_add_6_33_groupi_n_2613 ,csa_tree_add_6_33_groupi_n_3361);
  or csa_tree_add_6_33_groupi_g14749(csa_tree_add_6_33_groupi_n_3510 ,csa_tree_add_6_33_groupi_n_3024 ,csa_tree_add_6_33_groupi_n_3375);
  or csa_tree_add_6_33_groupi_g14750(csa_tree_add_6_33_groupi_n_3509 ,csa_tree_add_6_33_groupi_n_2692 ,csa_tree_add_6_33_groupi_n_3362);
  and csa_tree_add_6_33_groupi_g14751(csa_tree_add_6_33_groupi_n_3508 ,csa_tree_add_6_33_groupi_n_2692 ,csa_tree_add_6_33_groupi_n_3362);
  or csa_tree_add_6_33_groupi_g14752(csa_tree_add_6_33_groupi_n_3507 ,csa_tree_add_6_33_groupi_n_2621 ,csa_tree_add_6_33_groupi_n_3347);
  or csa_tree_add_6_33_groupi_g14753(csa_tree_add_6_33_groupi_n_3506 ,csa_tree_add_6_33_groupi_n_3320 ,csa_tree_add_6_33_groupi_n_3378);
  or csa_tree_add_6_33_groupi_g14754(csa_tree_add_6_33_groupi_n_3505 ,csa_tree_add_6_33_groupi_n_3348 ,csa_tree_add_6_33_groupi_n_3050);
  nor csa_tree_add_6_33_groupi_g14755(csa_tree_add_6_33_groupi_n_3504 ,csa_tree_add_6_33_groupi_n_2681 ,csa_tree_add_6_33_groupi_n_3359);
  nor csa_tree_add_6_33_groupi_g14756(csa_tree_add_6_33_groupi_n_3503 ,csa_tree_add_6_33_groupi_n_2890 ,csa_tree_add_6_33_groupi_n_3357);
  nor csa_tree_add_6_33_groupi_g14757(csa_tree_add_6_33_groupi_n_3502 ,csa_tree_add_6_33_groupi_n_2631 ,csa_tree_add_6_33_groupi_n_3275);
  or csa_tree_add_6_33_groupi_g14758(csa_tree_add_6_33_groupi_n_3501 ,csa_tree_add_6_33_groupi_n_3141 ,csa_tree_add_6_33_groupi_n_3379);
  or csa_tree_add_6_33_groupi_g14759(csa_tree_add_6_33_groupi_n_3500 ,csa_tree_add_6_33_groupi_n_2632 ,csa_tree_add_6_33_groupi_n_3274);
  nor csa_tree_add_6_33_groupi_g14760(csa_tree_add_6_33_groupi_n_3499 ,csa_tree_add_6_33_groupi_n_3052 ,csa_tree_add_6_33_groupi_n_3349);
  or csa_tree_add_6_33_groupi_g14761(csa_tree_add_6_33_groupi_n_3498 ,csa_tree_add_6_33_groupi_n_3125 ,csa_tree_add_6_33_groupi_n_3288);
  or csa_tree_add_6_33_groupi_g14762(csa_tree_add_6_33_groupi_n_3497 ,csa_tree_add_6_33_groupi_n_2982 ,csa_tree_add_6_33_groupi_n_3383);
  or csa_tree_add_6_33_groupi_g14763(csa_tree_add_6_33_groupi_n_3496 ,csa_tree_add_6_33_groupi_n_2889 ,csa_tree_add_6_33_groupi_n_3356);
  or csa_tree_add_6_33_groupi_g14764(csa_tree_add_6_33_groupi_n_3495 ,csa_tree_add_6_33_groupi_n_2680 ,csa_tree_add_6_33_groupi_n_3358);
  or csa_tree_add_6_33_groupi_g14765(csa_tree_add_6_33_groupi_n_3494 ,csa_tree_add_6_33_groupi_n_3388 ,csa_tree_add_6_33_groupi_n_3331);
  and csa_tree_add_6_33_groupi_g14766(csa_tree_add_6_33_groupi_n_3493 ,csa_tree_add_6_33_groupi_n_3185 ,csa_tree_add_6_33_groupi_n_3271);
  or csa_tree_add_6_33_groupi_g14767(csa_tree_add_6_33_groupi_n_3492 ,csa_tree_add_6_33_groupi_n_3051 ,csa_tree_add_6_33_groupi_n_3350);
  or csa_tree_add_6_33_groupi_g14768(csa_tree_add_6_33_groupi_n_3491 ,csa_tree_add_6_33_groupi_n_3385 ,csa_tree_add_6_33_groupi_n_3304);
  nor csa_tree_add_6_33_groupi_g14769(csa_tree_add_6_33_groupi_n_3490 ,csa_tree_add_6_33_groupi_n_3354 ,csa_tree_add_6_33_groupi_n_3268);
  or csa_tree_add_6_33_groupi_g14770(csa_tree_add_6_33_groupi_n_3489 ,csa_tree_add_6_33_groupi_n_3355 ,csa_tree_add_6_33_groupi_n_3267);
  or csa_tree_add_6_33_groupi_g14771(csa_tree_add_6_33_groupi_n_3488 ,csa_tree_add_6_33_groupi_n_3185 ,csa_tree_add_6_33_groupi_n_3271);
  and csa_tree_add_6_33_groupi_g14772(csa_tree_add_6_33_groupi_n_3572 ,csa_tree_add_6_33_groupi_n_3090 ,csa_tree_add_6_33_groupi_n_3316);
  and csa_tree_add_6_33_groupi_g14773(csa_tree_add_6_33_groupi_n_3571 ,csa_tree_add_6_33_groupi_n_3093 ,csa_tree_add_6_33_groupi_n_3297);
  and csa_tree_add_6_33_groupi_g14774(csa_tree_add_6_33_groupi_n_3570 ,csa_tree_add_6_33_groupi_n_3079 ,csa_tree_add_6_33_groupi_n_3302);
  and csa_tree_add_6_33_groupi_g14775(csa_tree_add_6_33_groupi_n_3569 ,csa_tree_add_6_33_groupi_n_3136 ,csa_tree_add_6_33_groupi_n_3313);
  and csa_tree_add_6_33_groupi_g14776(csa_tree_add_6_33_groupi_n_3568 ,csa_tree_add_6_33_groupi_n_3073 ,csa_tree_add_6_33_groupi_n_3314);
  and csa_tree_add_6_33_groupi_g14777(csa_tree_add_6_33_groupi_n_3567 ,csa_tree_add_6_33_groupi_n_3072 ,csa_tree_add_6_33_groupi_n_3315);
  and csa_tree_add_6_33_groupi_g14778(csa_tree_add_6_33_groupi_n_3566 ,csa_tree_add_6_33_groupi_n_3071 ,csa_tree_add_6_33_groupi_n_3308);
  and csa_tree_add_6_33_groupi_g14779(csa_tree_add_6_33_groupi_n_3565 ,csa_tree_add_6_33_groupi_n_3179 ,csa_tree_add_6_33_groupi_n_3338);
  and csa_tree_add_6_33_groupi_g14780(csa_tree_add_6_33_groupi_n_3564 ,csa_tree_add_6_33_groupi_n_3103 ,csa_tree_add_6_33_groupi_n_3293);
  and csa_tree_add_6_33_groupi_g14781(csa_tree_add_6_33_groupi_n_3563 ,csa_tree_add_6_33_groupi_n_3062 ,csa_tree_add_6_33_groupi_n_3319);
  and csa_tree_add_6_33_groupi_g14782(csa_tree_add_6_33_groupi_n_3562 ,csa_tree_add_6_33_groupi_n_3084 ,csa_tree_add_6_33_groupi_n_3326);
  and csa_tree_add_6_33_groupi_g14783(csa_tree_add_6_33_groupi_n_3561 ,csa_tree_add_6_33_groupi_n_2992 ,csa_tree_add_6_33_groupi_n_3310);
  and csa_tree_add_6_33_groupi_g14784(csa_tree_add_6_33_groupi_n_3560 ,csa_tree_add_6_33_groupi_n_3134 ,csa_tree_add_6_33_groupi_n_3312);
  and csa_tree_add_6_33_groupi_g14785(csa_tree_add_6_33_groupi_n_3559 ,csa_tree_add_6_33_groupi_n_3155 ,csa_tree_add_6_33_groupi_n_3329);
  and csa_tree_add_6_33_groupi_g14786(csa_tree_add_6_33_groupi_n_3558 ,csa_tree_add_6_33_groupi_n_3061 ,csa_tree_add_6_33_groupi_n_3294);
  and csa_tree_add_6_33_groupi_g14787(csa_tree_add_6_33_groupi_n_3557 ,csa_tree_add_6_33_groupi_n_3033 ,csa_tree_add_6_33_groupi_n_3335);
  and csa_tree_add_6_33_groupi_g14788(csa_tree_add_6_33_groupi_n_3556 ,csa_tree_add_6_33_groupi_n_3030 ,csa_tree_add_6_33_groupi_n_3342);
  and csa_tree_add_6_33_groupi_g14789(csa_tree_add_6_33_groupi_n_3555 ,csa_tree_add_6_33_groupi_n_3142 ,csa_tree_add_6_33_groupi_n_3317);
  and csa_tree_add_6_33_groupi_g14790(csa_tree_add_6_33_groupi_n_3554 ,csa_tree_add_6_33_groupi_n_3146 ,csa_tree_add_6_33_groupi_n_3318);
  and csa_tree_add_6_33_groupi_g14791(csa_tree_add_6_33_groupi_n_3553 ,csa_tree_add_6_33_groupi_n_3151 ,csa_tree_add_6_33_groupi_n_3324);
  and csa_tree_add_6_33_groupi_g14792(csa_tree_add_6_33_groupi_n_3552 ,csa_tree_add_6_33_groupi_n_3160 ,csa_tree_add_6_33_groupi_n_3327);
  and csa_tree_add_6_33_groupi_g14793(csa_tree_add_6_33_groupi_n_3551 ,csa_tree_add_6_33_groupi_n_3167 ,csa_tree_add_6_33_groupi_n_3333);
  and csa_tree_add_6_33_groupi_g14794(csa_tree_add_6_33_groupi_n_3550 ,csa_tree_add_6_33_groupi_n_3022 ,csa_tree_add_6_33_groupi_n_3263);
  and csa_tree_add_6_33_groupi_g14795(csa_tree_add_6_33_groupi_n_3549 ,csa_tree_add_6_33_groupi_n_3173 ,csa_tree_add_6_33_groupi_n_3330);
  and csa_tree_add_6_33_groupi_g14796(csa_tree_add_6_33_groupi_n_3548 ,csa_tree_add_6_33_groupi_n_3012 ,csa_tree_add_6_33_groupi_n_3253);
  and csa_tree_add_6_33_groupi_g14797(csa_tree_add_6_33_groupi_n_3547 ,csa_tree_add_6_33_groupi_n_3011 ,csa_tree_add_6_33_groupi_n_3259);
  and csa_tree_add_6_33_groupi_g14798(csa_tree_add_6_33_groupi_n_3546 ,csa_tree_add_6_33_groupi_n_3176 ,csa_tree_add_6_33_groupi_n_3337);
  and csa_tree_add_6_33_groupi_g14799(csa_tree_add_6_33_groupi_n_3545 ,csa_tree_add_6_33_groupi_n_3101 ,csa_tree_add_6_33_groupi_n_3306);
  and csa_tree_add_6_33_groupi_g14800(csa_tree_add_6_33_groupi_n_3544 ,csa_tree_add_6_33_groupi_n_3120 ,csa_tree_add_6_33_groupi_n_3261);
  and csa_tree_add_6_33_groupi_g14801(csa_tree_add_6_33_groupi_n_3542 ,csa_tree_add_6_33_groupi_n_3109 ,csa_tree_add_6_33_groupi_n_3298);
  and csa_tree_add_6_33_groupi_g14802(csa_tree_add_6_33_groupi_n_3540 ,csa_tree_add_6_33_groupi_n_2979 ,csa_tree_add_6_33_groupi_n_3334);
  and csa_tree_add_6_33_groupi_g14803(csa_tree_add_6_33_groupi_n_3539 ,csa_tree_add_6_33_groupi_n_3150 ,csa_tree_add_6_33_groupi_n_3323);
  and csa_tree_add_6_33_groupi_g14804(csa_tree_add_6_33_groupi_n_3537 ,csa_tree_add_6_33_groupi_n_3129 ,csa_tree_add_6_33_groupi_n_3309);
  and csa_tree_add_6_33_groupi_g14805(csa_tree_add_6_33_groupi_n_3536 ,csa_tree_add_6_33_groupi_n_3149 ,csa_tree_add_6_33_groupi_n_3322);
  and csa_tree_add_6_33_groupi_g14806(csa_tree_add_6_33_groupi_n_3535 ,csa_tree_add_6_33_groupi_n_3175 ,csa_tree_add_6_33_groupi_n_3336);
  and csa_tree_add_6_33_groupi_g14807(csa_tree_add_6_33_groupi_n_3534 ,csa_tree_add_6_33_groupi_n_3095 ,csa_tree_add_6_33_groupi_n_3340);
  and csa_tree_add_6_33_groupi_g14808(csa_tree_add_6_33_groupi_n_3533 ,csa_tree_add_6_33_groupi_n_3115 ,csa_tree_add_6_33_groupi_n_3328);
  and csa_tree_add_6_33_groupi_g14809(csa_tree_add_6_33_groupi_n_3532 ,csa_tree_add_6_33_groupi_n_3028 ,csa_tree_add_6_33_groupi_n_3262);
  and csa_tree_add_6_33_groupi_g14810(csa_tree_add_6_33_groupi_n_3531 ,csa_tree_add_6_33_groupi_n_3063 ,csa_tree_add_6_33_groupi_n_3321);
  and csa_tree_add_6_33_groupi_g14811(csa_tree_add_6_33_groupi_n_3529 ,csa_tree_add_6_33_groupi_n_3019 ,csa_tree_add_6_33_groupi_n_3257);
  and csa_tree_add_6_33_groupi_g14812(csa_tree_add_6_33_groupi_n_3528 ,csa_tree_add_6_33_groupi_n_3015 ,csa_tree_add_6_33_groupi_n_3260);
  and csa_tree_add_6_33_groupi_g14813(csa_tree_add_6_33_groupi_n_3527 ,csa_tree_add_6_33_groupi_n_3009 ,csa_tree_add_6_33_groupi_n_3256);
  and csa_tree_add_6_33_groupi_g14814(csa_tree_add_6_33_groupi_n_3526 ,csa_tree_add_6_33_groupi_n_3119 ,csa_tree_add_6_33_groupi_n_3305);
  or csa_tree_add_6_33_groupi_g14815(csa_tree_add_6_33_groupi_n_3525 ,csa_tree_add_6_33_groupi_n_3086 ,csa_tree_add_6_33_groupi_n_3300);
  or csa_tree_add_6_33_groupi_g14816(csa_tree_add_6_33_groupi_n_3523 ,csa_tree_add_6_33_groupi_n_3180 ,csa_tree_add_6_33_groupi_n_3341);
  not csa_tree_add_6_33_groupi_g14817(csa_tree_add_6_33_groupi_n_3479 ,csa_tree_add_6_33_groupi_n_3478);
  not csa_tree_add_6_33_groupi_g14818(csa_tree_add_6_33_groupi_n_3475 ,csa_tree_add_6_33_groupi_n_3474);
  not csa_tree_add_6_33_groupi_g14819(csa_tree_add_6_33_groupi_n_3473 ,csa_tree_add_6_33_groupi_n_3472);
  not csa_tree_add_6_33_groupi_g14820(csa_tree_add_6_33_groupi_n_3464 ,csa_tree_add_6_33_groupi_n_3465);
  not csa_tree_add_6_33_groupi_g14821(csa_tree_add_6_33_groupi_n_3455 ,csa_tree_add_6_33_groupi_n_3456);
  not csa_tree_add_6_33_groupi_g14822(csa_tree_add_6_33_groupi_n_3453 ,csa_tree_add_6_33_groupi_n_3454);
  not csa_tree_add_6_33_groupi_g14823(csa_tree_add_6_33_groupi_n_3449 ,csa_tree_add_6_33_groupi_n_3448);
  not csa_tree_add_6_33_groupi_g14824(csa_tree_add_6_33_groupi_n_3442 ,csa_tree_add_6_33_groupi_n_3443);
  not csa_tree_add_6_33_groupi_g14825(csa_tree_add_6_33_groupi_n_3439 ,csa_tree_add_6_33_groupi_n_3440);
  not csa_tree_add_6_33_groupi_g14826(csa_tree_add_6_33_groupi_n_3434 ,csa_tree_add_6_33_groupi_n_3435);
  not csa_tree_add_6_33_groupi_g14827(csa_tree_add_6_33_groupi_n_3432 ,csa_tree_add_6_33_groupi_n_3433);
  not csa_tree_add_6_33_groupi_g14828(csa_tree_add_6_33_groupi_n_3429 ,csa_tree_add_6_33_groupi_n_3430);
  not csa_tree_add_6_33_groupi_g14829(csa_tree_add_6_33_groupi_n_3422 ,csa_tree_add_6_33_groupi_n_3423);
  not csa_tree_add_6_33_groupi_g14830(csa_tree_add_6_33_groupi_n_3415 ,csa_tree_add_6_33_groupi_n_3416);
  not csa_tree_add_6_33_groupi_g14831(csa_tree_add_6_33_groupi_n_3410 ,csa_tree_add_6_33_groupi_n_3411);
  not csa_tree_add_6_33_groupi_g14832(csa_tree_add_6_33_groupi_n_3408 ,csa_tree_add_6_33_groupi_n_3409);
  not csa_tree_add_6_33_groupi_g14833(csa_tree_add_6_33_groupi_n_3407 ,csa_tree_add_6_33_groupi_n_3406);
  or csa_tree_add_6_33_groupi_g14834(csa_tree_add_6_33_groupi_n_3405 ,csa_tree_add_6_33_groupi_n_3286 ,csa_tree_add_6_33_groupi_n_3255);
  xnor csa_tree_add_6_33_groupi_g14835(out1[2] ,csa_tree_add_6_33_groupi_n_2912 ,csa_tree_add_6_33_groupi_n_2972);
  and csa_tree_add_6_33_groupi_g14836(csa_tree_add_6_33_groupi_n_3403 ,csa_tree_add_6_33_groupi_n_3390 ,csa_tree_add_6_33_groupi_n_3132);
  or csa_tree_add_6_33_groupi_g14837(csa_tree_add_6_33_groupi_n_3402 ,csa_tree_add_6_33_groupi_n_2994 ,csa_tree_add_6_33_groupi_n_3280);
  or csa_tree_add_6_33_groupi_g14838(csa_tree_add_6_33_groupi_n_3401 ,csa_tree_add_6_33_groupi_n_3045 ,csa_tree_add_6_33_groupi_n_3265);
  nor csa_tree_add_6_33_groupi_g14839(csa_tree_add_6_33_groupi_n_3400 ,csa_tree_add_6_33_groupi_n_3046 ,csa_tree_add_6_33_groupi_n_3266);
  nor csa_tree_add_6_33_groupi_g14840(csa_tree_add_6_33_groupi_n_3399 ,csa_tree_add_6_33_groupi_n_2882 ,csa_tree_add_6_33_groupi_n_3282);
  or csa_tree_add_6_33_groupi_g14841(csa_tree_add_6_33_groupi_n_3398 ,csa_tree_add_6_33_groupi_n_3292 ,csa_tree_add_6_33_groupi_n_2987);
  xnor csa_tree_add_6_33_groupi_g14842(csa_tree_add_6_33_groupi_n_3397 ,csa_tree_add_6_33_groupi_n_2349 ,csa_tree_add_6_33_groupi_n_3056);
  xnor csa_tree_add_6_33_groupi_g14843(csa_tree_add_6_33_groupi_n_3396 ,csa_tree_add_6_33_groupi_n_2653 ,csa_tree_add_6_33_groupi_n_3188);
  xnor csa_tree_add_6_33_groupi_g14844(csa_tree_add_6_33_groupi_n_3395 ,csa_tree_add_6_33_groupi_n_3038 ,csa_tree_add_6_33_groupi_n_2892);
  xnor csa_tree_add_6_33_groupi_g14845(csa_tree_add_6_33_groupi_n_3394 ,csa_tree_add_6_33_groupi_n_3043 ,csa_tree_add_6_33_groupi_n_2650);
  xnor csa_tree_add_6_33_groupi_g14846(csa_tree_add_6_33_groupi_n_3393 ,csa_tree_add_6_33_groupi_n_2698 ,csa_tree_add_6_33_groupi_n_3040);
  xnor csa_tree_add_6_33_groupi_g14847(csa_tree_add_6_33_groupi_n_3392 ,csa_tree_add_6_33_groupi_n_2602 ,csa_tree_add_6_33_groupi_n_3054);
  xnor csa_tree_add_6_33_groupi_g14848(csa_tree_add_6_33_groupi_n_3391 ,csa_tree_add_6_33_groupi_n_3049 ,csa_tree_add_6_33_groupi_n_2651);
  and csa_tree_add_6_33_groupi_g14849(csa_tree_add_6_33_groupi_n_3487 ,csa_tree_add_6_33_groupi_n_2993 ,csa_tree_add_6_33_groupi_n_3250);
  xnor csa_tree_add_6_33_groupi_g14850(csa_tree_add_6_33_groupi_n_3486 ,csa_tree_add_6_33_groupi_n_2505 ,csa_tree_add_6_33_groupi_n_2943);
  xnor csa_tree_add_6_33_groupi_g14851(csa_tree_add_6_33_groupi_n_3485 ,csa_tree_add_6_33_groupi_n_2746 ,csa_tree_add_6_33_groupi_n_2976);
  xnor csa_tree_add_6_33_groupi_g14852(csa_tree_add_6_33_groupi_n_3484 ,csa_tree_add_6_33_groupi_n_2527 ,csa_tree_add_6_33_groupi_n_2938);
  and csa_tree_add_6_33_groupi_g14853(csa_tree_add_6_33_groupi_n_3483 ,csa_tree_add_6_33_groupi_n_3001 ,csa_tree_add_6_33_groupi_n_3254);
  and csa_tree_add_6_33_groupi_g14854(csa_tree_add_6_33_groupi_n_3482 ,csa_tree_add_6_33_groupi_n_2986 ,csa_tree_add_6_33_groupi_n_3343);
  and csa_tree_add_6_33_groupi_g14855(csa_tree_add_6_33_groupi_n_3481 ,csa_tree_add_6_33_groupi_n_3002 ,csa_tree_add_6_33_groupi_n_3252);
  xnor csa_tree_add_6_33_groupi_g14856(csa_tree_add_6_33_groupi_n_3480 ,csa_tree_add_6_33_groupi_n_2355 ,csa_tree_add_6_33_groupi_n_2960);
  xnor csa_tree_add_6_33_groupi_g14857(csa_tree_add_6_33_groupi_n_3478 ,csa_tree_add_6_33_groupi_n_2340 ,csa_tree_add_6_33_groupi_n_2964);
  and csa_tree_add_6_33_groupi_g14858(csa_tree_add_6_33_groupi_n_3477 ,csa_tree_add_6_33_groupi_n_2996 ,csa_tree_add_6_33_groupi_n_3251);
  xnor csa_tree_add_6_33_groupi_g14859(csa_tree_add_6_33_groupi_n_3476 ,csa_tree_add_6_33_groupi_n_2348 ,csa_tree_add_6_33_groupi_n_2969);
  xnor csa_tree_add_6_33_groupi_g14860(csa_tree_add_6_33_groupi_n_3474 ,csa_tree_add_6_33_groupi_n_2365 ,csa_tree_add_6_33_groupi_n_2963);
  xnor csa_tree_add_6_33_groupi_g14861(csa_tree_add_6_33_groupi_n_3472 ,csa_tree_add_6_33_groupi_n_2419 ,csa_tree_add_6_33_groupi_n_2955);
  xnor csa_tree_add_6_33_groupi_g14862(csa_tree_add_6_33_groupi_n_3471 ,csa_tree_add_6_33_groupi_n_2395 ,csa_tree_add_6_33_groupi_n_2958);
  xnor csa_tree_add_6_33_groupi_g14863(csa_tree_add_6_33_groupi_n_3470 ,csa_tree_add_6_33_groupi_n_2745 ,csa_tree_add_6_33_groupi_n_2956);
  xnor csa_tree_add_6_33_groupi_g14864(csa_tree_add_6_33_groupi_n_3469 ,csa_tree_add_6_33_groupi_n_2739 ,csa_tree_add_6_33_groupi_n_2948);
  xnor csa_tree_add_6_33_groupi_g14865(csa_tree_add_6_33_groupi_n_3468 ,csa_tree_add_6_33_groupi_n_2545 ,csa_tree_add_6_33_groupi_n_2954);
  xnor csa_tree_add_6_33_groupi_g14866(csa_tree_add_6_33_groupi_n_3467 ,csa_tree_add_6_33_groupi_n_2472 ,csa_tree_add_6_33_groupi_n_2953);
  xnor csa_tree_add_6_33_groupi_g14867(csa_tree_add_6_33_groupi_n_3466 ,csa_tree_add_6_33_groupi_n_2463 ,csa_tree_add_6_33_groupi_n_2952);
  xnor csa_tree_add_6_33_groupi_g14868(csa_tree_add_6_33_groupi_n_3465 ,csa_tree_add_6_33_groupi_n_2378 ,csa_tree_add_6_33_groupi_n_2959);
  xnor csa_tree_add_6_33_groupi_g14869(csa_tree_add_6_33_groupi_n_3463 ,csa_tree_add_6_33_groupi_n_2515 ,csa_tree_add_6_33_groupi_n_2951);
  xnor csa_tree_add_6_33_groupi_g14870(csa_tree_add_6_33_groupi_n_3462 ,csa_tree_add_6_33_groupi_n_2452 ,csa_tree_add_6_33_groupi_n_2949);
  xnor csa_tree_add_6_33_groupi_g14871(csa_tree_add_6_33_groupi_n_3461 ,csa_tree_add_6_33_groupi_n_2604 ,csa_tree_add_6_33_groupi_n_2950);
  xnor csa_tree_add_6_33_groupi_g14872(csa_tree_add_6_33_groupi_n_3460 ,csa_tree_add_6_33_groupi_n_2455 ,csa_tree_add_6_33_groupi_n_2936);
  xnor csa_tree_add_6_33_groupi_g14873(csa_tree_add_6_33_groupi_n_3459 ,csa_tree_add_6_33_groupi_n_2568 ,csa_tree_add_6_33_groupi_n_2947);
  xnor csa_tree_add_6_33_groupi_g14874(csa_tree_add_6_33_groupi_n_3458 ,csa_tree_add_6_33_groupi_n_2422 ,csa_tree_add_6_33_groupi_n_2946);
  xnor csa_tree_add_6_33_groupi_g14875(csa_tree_add_6_33_groupi_n_3457 ,csa_tree_add_6_33_groupi_n_2536 ,csa_tree_add_6_33_groupi_n_2920);
  xnor csa_tree_add_6_33_groupi_g14876(csa_tree_add_6_33_groupi_n_3456 ,csa_tree_add_6_33_groupi_n_2611 ,csa_tree_add_6_33_groupi_n_2944);
  xnor csa_tree_add_6_33_groupi_g14877(csa_tree_add_6_33_groupi_n_3454 ,csa_tree_add_6_33_groupi_n_2582 ,csa_tree_add_6_33_groupi_n_2961);
  xnor csa_tree_add_6_33_groupi_g14878(csa_tree_add_6_33_groupi_n_3452 ,csa_tree_add_6_33_groupi_n_2539 ,csa_tree_add_6_33_groupi_n_2941);
  xnor csa_tree_add_6_33_groupi_g14879(csa_tree_add_6_33_groupi_n_3451 ,csa_tree_add_6_33_groupi_n_2596 ,csa_tree_add_6_33_groupi_n_2940);
  xnor csa_tree_add_6_33_groupi_g14880(csa_tree_add_6_33_groupi_n_3450 ,csa_tree_add_6_33_groupi_n_2453 ,csa_tree_add_6_33_groupi_n_2939);
  xnor csa_tree_add_6_33_groupi_g14881(csa_tree_add_6_33_groupi_n_3448 ,csa_tree_add_6_33_groupi_n_2665 ,csa_tree_add_6_33_groupi_n_2966);
  xnor csa_tree_add_6_33_groupi_g14882(csa_tree_add_6_33_groupi_n_3447 ,csa_tree_add_6_33_groupi_n_2622 ,csa_tree_add_6_33_groupi_n_2937);
  xnor csa_tree_add_6_33_groupi_g14883(csa_tree_add_6_33_groupi_n_3446 ,csa_tree_add_6_33_groupi_n_2513 ,csa_tree_add_6_33_groupi_n_2934);
  xnor csa_tree_add_6_33_groupi_g14884(csa_tree_add_6_33_groupi_n_3445 ,csa_tree_add_6_33_groupi_n_2508 ,csa_tree_add_6_33_groupi_n_2928);
  xnor csa_tree_add_6_33_groupi_g14885(csa_tree_add_6_33_groupi_n_3444 ,csa_tree_add_6_33_groupi_n_2544 ,csa_tree_add_6_33_groupi_n_2931);
  xnor csa_tree_add_6_33_groupi_g14886(csa_tree_add_6_33_groupi_n_3443 ,csa_tree_add_6_33_groupi_n_2503 ,csa_tree_add_6_33_groupi_n_2932);
  xnor csa_tree_add_6_33_groupi_g14887(csa_tree_add_6_33_groupi_n_3441 ,csa_tree_add_6_33_groupi_n_2662 ,csa_tree_add_6_33_groupi_n_2929);
  xnor csa_tree_add_6_33_groupi_g14888(csa_tree_add_6_33_groupi_n_3440 ,csa_tree_add_6_33_groupi_n_2727 ,csa_tree_add_6_33_groupi_n_2962);
  xnor csa_tree_add_6_33_groupi_g14889(csa_tree_add_6_33_groupi_n_3438 ,csa_tree_add_6_33_groupi_n_2530 ,csa_tree_add_6_33_groupi_n_2927);
  xnor csa_tree_add_6_33_groupi_g14890(csa_tree_add_6_33_groupi_n_3437 ,csa_tree_add_6_33_groupi_n_2547 ,csa_tree_add_6_33_groupi_n_2925);
  xnor csa_tree_add_6_33_groupi_g14891(csa_tree_add_6_33_groupi_n_3436 ,csa_tree_add_6_33_groupi_n_2738 ,csa_tree_add_6_33_groupi_n_2923);
  xnor csa_tree_add_6_33_groupi_g14892(csa_tree_add_6_33_groupi_n_3435 ,csa_tree_add_6_33_groupi_n_2529 ,csa_tree_add_6_33_groupi_n_2922);
  xnor csa_tree_add_6_33_groupi_g14893(csa_tree_add_6_33_groupi_n_3433 ,csa_tree_add_6_33_groupi_n_2718 ,csa_tree_add_6_33_groupi_n_2942);
  xnor csa_tree_add_6_33_groupi_g14894(csa_tree_add_6_33_groupi_n_3431 ,csa_tree_add_6_33_groupi_n_2497 ,csa_tree_add_6_33_groupi_n_2921);
  xnor csa_tree_add_6_33_groupi_g14895(csa_tree_add_6_33_groupi_n_3430 ,csa_tree_add_6_33_groupi_n_2429 ,csa_tree_add_6_33_groupi_n_2919);
  xnor csa_tree_add_6_33_groupi_g14896(csa_tree_add_6_33_groupi_n_3428 ,csa_tree_add_6_33_groupi_n_2556 ,csa_tree_add_6_33_groupi_n_2918);
  xnor csa_tree_add_6_33_groupi_g14897(csa_tree_add_6_33_groupi_n_3427 ,csa_tree_add_6_33_groupi_n_2741 ,csa_tree_add_6_33_groupi_n_2916);
  xnor csa_tree_add_6_33_groupi_g14898(csa_tree_add_6_33_groupi_n_3426 ,csa_tree_add_6_33_groupi_n_2393 ,csa_tree_add_6_33_groupi_n_2917);
  xnor csa_tree_add_6_33_groupi_g14899(csa_tree_add_6_33_groupi_n_3425 ,csa_tree_add_6_33_groupi_n_2440 ,csa_tree_add_6_33_groupi_n_2924);
  xnor csa_tree_add_6_33_groupi_g14900(csa_tree_add_6_33_groupi_n_3424 ,csa_tree_add_6_33_groupi_n_2481 ,csa_tree_add_6_33_groupi_n_2926);
  xnor csa_tree_add_6_33_groupi_g14901(csa_tree_add_6_33_groupi_n_3423 ,csa_tree_add_6_33_groupi_n_2581 ,csa_tree_add_6_33_groupi_n_2965);
  xnor csa_tree_add_6_33_groupi_g14902(csa_tree_add_6_33_groupi_n_3421 ,csa_tree_add_6_33_groupi_n_2747 ,csa_tree_add_6_33_groupi_n_2930);
  xnor csa_tree_add_6_33_groupi_g14903(csa_tree_add_6_33_groupi_n_3420 ,csa_tree_add_6_33_groupi_n_2441 ,csa_tree_add_6_33_groupi_n_2935);
  xnor csa_tree_add_6_33_groupi_g14904(csa_tree_add_6_33_groupi_n_3419 ,csa_tree_add_6_33_groupi_n_2448 ,csa_tree_add_6_33_groupi_n_2967);
  xnor csa_tree_add_6_33_groupi_g14905(csa_tree_add_6_33_groupi_n_3418 ,csa_tree_add_6_33_groupi_n_2730 ,csa_tree_add_6_33_groupi_n_2970);
  xnor csa_tree_add_6_33_groupi_g14906(csa_tree_add_6_33_groupi_n_3417 ,csa_tree_add_6_33_groupi_n_2451 ,csa_tree_add_6_33_groupi_n_2974);
  xnor csa_tree_add_6_33_groupi_g14907(csa_tree_add_6_33_groupi_n_3416 ,csa_tree_add_6_33_groupi_n_2555 ,csa_tree_add_6_33_groupi_n_2973);
  xnor csa_tree_add_6_33_groupi_g14908(csa_tree_add_6_33_groupi_n_3414 ,csa_tree_add_6_33_groupi_n_2460 ,csa_tree_add_6_33_groupi_n_2977);
  xnor csa_tree_add_6_33_groupi_g14909(csa_tree_add_6_33_groupi_n_3413 ,csa_tree_add_6_33_groupi_n_2430 ,csa_tree_add_6_33_groupi_n_2975);
  xnor csa_tree_add_6_33_groupi_g14910(csa_tree_add_6_33_groupi_n_3412 ,csa_tree_add_6_33_groupi_n_2474 ,csa_tree_add_6_33_groupi_n_2945);
  xnor csa_tree_add_6_33_groupi_g14911(csa_tree_add_6_33_groupi_n_3411 ,csa_tree_add_6_33_groupi_n_2593 ,csa_tree_add_6_33_groupi_n_2978);
  xnor csa_tree_add_6_33_groupi_g14912(csa_tree_add_6_33_groupi_n_3409 ,csa_tree_add_6_33_groupi_n_2569 ,csa_tree_add_6_33_groupi_n_2971);
  xnor csa_tree_add_6_33_groupi_g14913(csa_tree_add_6_33_groupi_n_3406 ,csa_tree_add_6_33_groupi_n_2688 ,csa_tree_add_6_33_groupi_n_2957);
  not csa_tree_add_6_33_groupi_g14914(csa_tree_add_6_33_groupi_n_3368 ,csa_tree_add_6_33_groupi_n_3369);
  not csa_tree_add_6_33_groupi_g14915(csa_tree_add_6_33_groupi_n_3361 ,csa_tree_add_6_33_groupi_n_3360);
  not csa_tree_add_6_33_groupi_g14916(csa_tree_add_6_33_groupi_n_3358 ,csa_tree_add_6_33_groupi_n_3359);
  not csa_tree_add_6_33_groupi_g14917(csa_tree_add_6_33_groupi_n_3356 ,csa_tree_add_6_33_groupi_n_3357);
  not csa_tree_add_6_33_groupi_g14918(csa_tree_add_6_33_groupi_n_3354 ,csa_tree_add_6_33_groupi_n_3355);
  not csa_tree_add_6_33_groupi_g14919(csa_tree_add_6_33_groupi_n_3351 ,csa_tree_add_6_33_groupi_n_3352);
  not csa_tree_add_6_33_groupi_g14920(csa_tree_add_6_33_groupi_n_3349 ,csa_tree_add_6_33_groupi_n_3350);
  not csa_tree_add_6_33_groupi_g14921(csa_tree_add_6_33_groupi_n_3344 ,csa_tree_add_6_33_groupi_n_3345);
  or csa_tree_add_6_33_groupi_g14922(csa_tree_add_6_33_groupi_n_3343 ,csa_tree_add_6_33_groupi_n_2561 ,csa_tree_add_6_33_groupi_n_3183);
  or csa_tree_add_6_33_groupi_g14923(csa_tree_add_6_33_groupi_n_3342 ,csa_tree_add_6_33_groupi_n_2731 ,csa_tree_add_6_33_groupi_n_3029);
  and csa_tree_add_6_33_groupi_g14924(csa_tree_add_6_33_groupi_n_3341 ,csa_tree_add_6_33_groupi_n_2915 ,csa_tree_add_6_33_groupi_n_3178);
  or csa_tree_add_6_33_groupi_g14925(csa_tree_add_6_33_groupi_n_3340 ,csa_tree_add_6_33_groupi_n_2543 ,csa_tree_add_6_33_groupi_n_3087);
  or csa_tree_add_6_33_groupi_g14926(csa_tree_add_6_33_groupi_n_3339 ,csa_tree_add_6_33_groupi_n_2650 ,csa_tree_add_6_33_groupi_n_3043);
  or csa_tree_add_6_33_groupi_g14927(csa_tree_add_6_33_groupi_n_3338 ,csa_tree_add_6_33_groupi_n_2914 ,csa_tree_add_6_33_groupi_n_3172);
  or csa_tree_add_6_33_groupi_g14928(csa_tree_add_6_33_groupi_n_3337 ,csa_tree_add_6_33_groupi_n_2549 ,csa_tree_add_6_33_groupi_n_3174);
  or csa_tree_add_6_33_groupi_g14929(csa_tree_add_6_33_groupi_n_3336 ,csa_tree_add_6_33_groupi_n_2752 ,csa_tree_add_6_33_groupi_n_3171);
  or csa_tree_add_6_33_groupi_g14930(csa_tree_add_6_33_groupi_n_3335 ,csa_tree_add_6_33_groupi_n_2456 ,csa_tree_add_6_33_groupi_n_3027);
  or csa_tree_add_6_33_groupi_g14931(csa_tree_add_6_33_groupi_n_3334 ,csa_tree_add_6_33_groupi_n_2725 ,csa_tree_add_6_33_groupi_n_3032);
  or csa_tree_add_6_33_groupi_g14932(csa_tree_add_6_33_groupi_n_3333 ,csa_tree_add_6_33_groupi_n_2572 ,csa_tree_add_6_33_groupi_n_3165);
  or csa_tree_add_6_33_groupi_g14933(csa_tree_add_6_33_groupi_n_3332 ,csa_tree_add_6_33_groupi_n_3188 ,csa_tree_add_6_33_groupi_n_2653);
  and csa_tree_add_6_33_groupi_g14934(csa_tree_add_6_33_groupi_n_3331 ,csa_tree_add_6_33_groupi_n_2650 ,csa_tree_add_6_33_groupi_n_3043);
  or csa_tree_add_6_33_groupi_g14935(csa_tree_add_6_33_groupi_n_3330 ,csa_tree_add_6_33_groupi_n_2541 ,csa_tree_add_6_33_groupi_n_3159);
  or csa_tree_add_6_33_groupi_g14936(csa_tree_add_6_33_groupi_n_3329 ,csa_tree_add_6_33_groupi_n_2732 ,csa_tree_add_6_33_groupi_n_3034);
  or csa_tree_add_6_33_groupi_g14937(csa_tree_add_6_33_groupi_n_3328 ,csa_tree_add_6_33_groupi_n_2580 ,csa_tree_add_6_33_groupi_n_3158);
  or csa_tree_add_6_33_groupi_g14938(csa_tree_add_6_33_groupi_n_3327 ,csa_tree_add_6_33_groupi_n_2558 ,csa_tree_add_6_33_groupi_n_3156);
  or csa_tree_add_6_33_groupi_g14939(csa_tree_add_6_33_groupi_n_3326 ,csa_tree_add_6_33_groupi_n_2733 ,csa_tree_add_6_33_groupi_n_3085);
  or csa_tree_add_6_33_groupi_g14940(csa_tree_add_6_33_groupi_n_3325 ,csa_tree_add_6_33_groupi_n_3187 ,csa_tree_add_6_33_groupi_n_2609);
  or csa_tree_add_6_33_groupi_g14941(csa_tree_add_6_33_groupi_n_3324 ,csa_tree_add_6_33_groupi_n_3059 ,csa_tree_add_6_33_groupi_n_3148);
  or csa_tree_add_6_33_groupi_g14942(csa_tree_add_6_33_groupi_n_3323 ,csa_tree_add_6_33_groupi_n_2751 ,csa_tree_add_6_33_groupi_n_3088);
  or csa_tree_add_6_33_groupi_g14943(csa_tree_add_6_33_groupi_n_3322 ,csa_tree_add_6_33_groupi_n_3191 ,csa_tree_add_6_33_groupi_n_3139);
  or csa_tree_add_6_33_groupi_g14944(csa_tree_add_6_33_groupi_n_3321 ,csa_tree_add_6_33_groupi_n_2734 ,csa_tree_add_6_33_groupi_n_3092);
  and csa_tree_add_6_33_groupi_g14945(csa_tree_add_6_33_groupi_n_3320 ,csa_tree_add_6_33_groupi_n_3187 ,csa_tree_add_6_33_groupi_n_2609);
  or csa_tree_add_6_33_groupi_g14946(csa_tree_add_6_33_groupi_n_3319 ,csa_tree_add_6_33_groupi_n_2735 ,csa_tree_add_6_33_groupi_n_3083);
  or csa_tree_add_6_33_groupi_g14947(csa_tree_add_6_33_groupi_n_3318 ,csa_tree_add_6_33_groupi_n_2750 ,csa_tree_add_6_33_groupi_n_3145);
  or csa_tree_add_6_33_groupi_g14948(csa_tree_add_6_33_groupi_n_3317 ,csa_tree_add_6_33_groupi_n_2570 ,csa_tree_add_6_33_groupi_n_3182);
  or csa_tree_add_6_33_groupi_g14949(csa_tree_add_6_33_groupi_n_3316 ,csa_tree_add_6_33_groupi_n_2723 ,csa_tree_add_6_33_groupi_n_3060);
  or csa_tree_add_6_33_groupi_g14950(csa_tree_add_6_33_groupi_n_3315 ,csa_tree_add_6_33_groupi_n_2736 ,csa_tree_add_6_33_groupi_n_3081);
  or csa_tree_add_6_33_groupi_g14951(csa_tree_add_6_33_groupi_n_3314 ,csa_tree_add_6_33_groupi_n_2737 ,csa_tree_add_6_33_groupi_n_3069);
  or csa_tree_add_6_33_groupi_g14952(csa_tree_add_6_33_groupi_n_3313 ,csa_tree_add_6_33_groupi_n_2749 ,csa_tree_add_6_33_groupi_n_3153);
  or csa_tree_add_6_33_groupi_g14953(csa_tree_add_6_33_groupi_n_3312 ,csa_tree_add_6_33_groupi_n_2743 ,csa_tree_add_6_33_groupi_n_3130);
  nor csa_tree_add_6_33_groupi_g14954(csa_tree_add_6_33_groupi_n_3311 ,csa_tree_add_6_33_groupi_n_2698 ,csa_tree_add_6_33_groupi_n_3039);
  or csa_tree_add_6_33_groupi_g14955(csa_tree_add_6_33_groupi_n_3310 ,csa_tree_add_6_33_groupi_n_3192 ,csa_tree_add_6_33_groupi_n_3127);
  or csa_tree_add_6_33_groupi_g14956(csa_tree_add_6_33_groupi_n_3309 ,csa_tree_add_6_33_groupi_n_2740 ,csa_tree_add_6_33_groupi_n_3126);
  or csa_tree_add_6_33_groupi_g14957(csa_tree_add_6_33_groupi_n_3308 ,csa_tree_add_6_33_groupi_n_3195 ,csa_tree_add_6_33_groupi_n_3070);
  and csa_tree_add_6_33_groupi_g14958(csa_tree_add_6_33_groupi_n_3307 ,csa_tree_add_6_33_groupi_n_3188 ,csa_tree_add_6_33_groupi_n_2653);
  or csa_tree_add_6_33_groupi_g14959(csa_tree_add_6_33_groupi_n_3306 ,csa_tree_add_6_33_groupi_n_2744 ,csa_tree_add_6_33_groupi_n_3117);
  or csa_tree_add_6_33_groupi_g14960(csa_tree_add_6_33_groupi_n_3305 ,csa_tree_add_6_33_groupi_n_2754 ,csa_tree_add_6_33_groupi_n_3113);
  and csa_tree_add_6_33_groupi_g14961(csa_tree_add_6_33_groupi_n_3304 ,csa_tree_add_6_33_groupi_n_2651 ,csa_tree_add_6_33_groupi_n_3049);
  or csa_tree_add_6_33_groupi_g14962(csa_tree_add_6_33_groupi_n_3303 ,csa_tree_add_6_33_groupi_n_2651 ,csa_tree_add_6_33_groupi_n_3049);
  or csa_tree_add_6_33_groupi_g14963(csa_tree_add_6_33_groupi_n_3302 ,csa_tree_add_6_33_groupi_n_2755 ,csa_tree_add_6_33_groupi_n_3078);
  or csa_tree_add_6_33_groupi_g14964(csa_tree_add_6_33_groupi_n_3301 ,csa_tree_add_6_33_groupi_n_3038 ,csa_tree_add_6_33_groupi_n_2891);
  nor csa_tree_add_6_33_groupi_g14965(csa_tree_add_6_33_groupi_n_3300 ,csa_tree_add_6_33_groupi_n_3194 ,csa_tree_add_6_33_groupi_n_3082);
  and csa_tree_add_6_33_groupi_g14966(csa_tree_add_6_33_groupi_n_3299 ,csa_tree_add_6_33_groupi_n_2349 ,csa_tree_add_6_33_groupi_n_3056);
  or csa_tree_add_6_33_groupi_g14967(csa_tree_add_6_33_groupi_n_3298 ,csa_tree_add_6_33_groupi_n_2550 ,csa_tree_add_6_33_groupi_n_3106);
  or csa_tree_add_6_33_groupi_g14968(csa_tree_add_6_33_groupi_n_3297 ,csa_tree_add_6_33_groupi_n_2753 ,csa_tree_add_6_33_groupi_n_3104);
  nor csa_tree_add_6_33_groupi_g14969(csa_tree_add_6_33_groupi_n_3296 ,csa_tree_add_6_33_groupi_n_3037 ,csa_tree_add_6_33_groupi_n_2892);
  or csa_tree_add_6_33_groupi_g14970(csa_tree_add_6_33_groupi_n_3295 ,csa_tree_add_6_33_groupi_n_2349 ,csa_tree_add_6_33_groupi_n_3056);
  or csa_tree_add_6_33_groupi_g14971(csa_tree_add_6_33_groupi_n_3294 ,csa_tree_add_6_33_groupi_n_2742 ,csa_tree_add_6_33_groupi_n_3157);
  or csa_tree_add_6_33_groupi_g14972(csa_tree_add_6_33_groupi_n_3293 ,csa_tree_add_6_33_groupi_n_2552 ,csa_tree_add_6_33_groupi_n_3089);
  or csa_tree_add_6_33_groupi_g14973(csa_tree_add_6_33_groupi_n_3390 ,csa_tree_add_6_33_groupi_n_2856 ,csa_tree_add_6_33_groupi_n_3133);
  and csa_tree_add_6_33_groupi_g14974(csa_tree_add_6_33_groupi_n_3389 ,csa_tree_add_6_33_groupi_n_2818 ,csa_tree_add_6_33_groupi_n_3097);
  and csa_tree_add_6_33_groupi_g14975(csa_tree_add_6_33_groupi_n_3388 ,csa_tree_add_6_33_groupi_n_2836 ,csa_tree_add_6_33_groupi_n_3105);
  and csa_tree_add_6_33_groupi_g14976(csa_tree_add_6_33_groupi_n_3387 ,csa_tree_add_6_33_groupi_n_2808 ,csa_tree_add_6_33_groupi_n_3077);
  and csa_tree_add_6_33_groupi_g14977(csa_tree_add_6_33_groupi_n_3386 ,csa_tree_add_6_33_groupi_n_2840 ,csa_tree_add_6_33_groupi_n_3110);
  and csa_tree_add_6_33_groupi_g14978(csa_tree_add_6_33_groupi_n_3385 ,csa_tree_add_6_33_groupi_n_2806 ,csa_tree_add_6_33_groupi_n_3074);
  and csa_tree_add_6_33_groupi_g14979(csa_tree_add_6_33_groupi_n_3384 ,csa_tree_add_6_33_groupi_n_2760 ,csa_tree_add_6_33_groupi_n_3114);
  and csa_tree_add_6_33_groupi_g14980(csa_tree_add_6_33_groupi_n_3383 ,csa_tree_add_6_33_groupi_n_2849 ,csa_tree_add_6_33_groupi_n_3065);
  and csa_tree_add_6_33_groupi_g14981(csa_tree_add_6_33_groupi_n_3382 ,csa_tree_add_6_33_groupi_n_2799 ,csa_tree_add_6_33_groupi_n_3067);
  and csa_tree_add_6_33_groupi_g14982(csa_tree_add_6_33_groupi_n_3381 ,csa_tree_add_6_33_groupi_n_2885 ,csa_tree_add_6_33_groupi_n_3100);
  and csa_tree_add_6_33_groupi_g14983(csa_tree_add_6_33_groupi_n_3380 ,csa_tree_add_6_33_groupi_n_2778 ,csa_tree_add_6_33_groupi_n_3137);
  and csa_tree_add_6_33_groupi_g14984(csa_tree_add_6_33_groupi_n_3379 ,csa_tree_add_6_33_groupi_n_2861 ,csa_tree_add_6_33_groupi_n_3140);
  and csa_tree_add_6_33_groupi_g14985(csa_tree_add_6_33_groupi_n_3378 ,csa_tree_add_6_33_groupi_n_2867 ,csa_tree_add_6_33_groupi_n_3144);
  and csa_tree_add_6_33_groupi_g14986(csa_tree_add_6_33_groupi_n_3377 ,csa_tree_add_6_33_groupi_n_2791 ,csa_tree_add_6_33_groupi_n_3128);
  and csa_tree_add_6_33_groupi_g14987(csa_tree_add_6_33_groupi_n_3376 ,csa_tree_add_6_33_groupi_n_2876 ,csa_tree_add_6_33_groupi_n_3118);
  and csa_tree_add_6_33_groupi_g14988(csa_tree_add_6_33_groupi_n_3375 ,csa_tree_add_6_33_groupi_n_2839 ,csa_tree_add_6_33_groupi_n_3031);
  and csa_tree_add_6_33_groupi_g14989(csa_tree_add_6_33_groupi_n_3374 ,csa_tree_add_6_33_groupi_n_2878 ,csa_tree_add_6_33_groupi_n_3162);
  and csa_tree_add_6_33_groupi_g14990(csa_tree_add_6_33_groupi_n_3373 ,csa_tree_add_6_33_groupi_n_2782 ,csa_tree_add_6_33_groupi_n_3026);
  and csa_tree_add_6_33_groupi_g14991(csa_tree_add_6_33_groupi_n_3372 ,csa_tree_add_6_33_groupi_n_2879 ,csa_tree_add_6_33_groupi_n_3096);
  and csa_tree_add_6_33_groupi_g14992(csa_tree_add_6_33_groupi_n_3371 ,csa_tree_add_6_33_groupi_n_2816 ,csa_tree_add_6_33_groupi_n_3094);
  or csa_tree_add_6_33_groupi_g14993(csa_tree_add_6_33_groupi_n_3370 ,csa_tree_add_6_33_groupi_n_2853 ,csa_tree_add_6_33_groupi_n_3111);
  and csa_tree_add_6_33_groupi_g14994(csa_tree_add_6_33_groupi_n_3369 ,csa_tree_add_6_33_groupi_n_2826 ,csa_tree_add_6_33_groupi_n_3163);
  and csa_tree_add_6_33_groupi_g14995(csa_tree_add_6_33_groupi_n_3367 ,csa_tree_add_6_33_groupi_n_2807 ,csa_tree_add_6_33_groupi_n_3076);
  and csa_tree_add_6_33_groupi_g14996(csa_tree_add_6_33_groupi_n_3366 ,csa_tree_add_6_33_groupi_n_2798 ,csa_tree_add_6_33_groupi_n_3066);
  and csa_tree_add_6_33_groupi_g14997(csa_tree_add_6_33_groupi_n_3365 ,csa_tree_add_6_33_groupi_n_2787 ,csa_tree_add_6_33_groupi_n_3147);
  and csa_tree_add_6_33_groupi_g14998(csa_tree_add_6_33_groupi_n_3364 ,csa_tree_add_6_33_groupi_n_2794 ,csa_tree_add_6_33_groupi_n_3107);
  or csa_tree_add_6_33_groupi_g14999(csa_tree_add_6_33_groupi_n_3363 ,csa_tree_add_6_33_groupi_n_2841 ,csa_tree_add_6_33_groupi_n_3112);
  and csa_tree_add_6_33_groupi_g15000(csa_tree_add_6_33_groupi_n_3362 ,csa_tree_add_6_33_groupi_n_2873 ,csa_tree_add_6_33_groupi_n_3154);
  and csa_tree_add_6_33_groupi_g15001(csa_tree_add_6_33_groupi_n_3360 ,csa_tree_add_6_33_groupi_n_2874 ,csa_tree_add_6_33_groupi_n_3161);
  and csa_tree_add_6_33_groupi_g15002(csa_tree_add_6_33_groupi_n_3359 ,csa_tree_add_6_33_groupi_n_2822 ,csa_tree_add_6_33_groupi_n_3121);
  and csa_tree_add_6_33_groupi_g15003(csa_tree_add_6_33_groupi_n_3357 ,csa_tree_add_6_33_groupi_n_2848 ,csa_tree_add_6_33_groupi_n_3122);
  and csa_tree_add_6_33_groupi_g15004(csa_tree_add_6_33_groupi_n_3355 ,csa_tree_add_6_33_groupi_n_2810 ,csa_tree_add_6_33_groupi_n_3080);
  or csa_tree_add_6_33_groupi_g15005(csa_tree_add_6_33_groupi_n_3353 ,csa_tree_add_6_33_groupi_n_2870 ,csa_tree_add_6_33_groupi_n_3169);
  and csa_tree_add_6_33_groupi_g15006(csa_tree_add_6_33_groupi_n_3352 ,csa_tree_add_6_33_groupi_n_2884 ,csa_tree_add_6_33_groupi_n_3177);
  and csa_tree_add_6_33_groupi_g15007(csa_tree_add_6_33_groupi_n_3350 ,csa_tree_add_6_33_groupi_n_2801 ,csa_tree_add_6_33_groupi_n_3068);
  and csa_tree_add_6_33_groupi_g15008(csa_tree_add_6_33_groupi_n_3348 ,csa_tree_add_6_33_groupi_n_2781 ,csa_tree_add_6_33_groupi_n_3020);
  and csa_tree_add_6_33_groupi_g15009(csa_tree_add_6_33_groupi_n_3347 ,csa_tree_add_6_33_groupi_n_2780 ,csa_tree_add_6_33_groupi_n_3023);
  and csa_tree_add_6_33_groupi_g15010(csa_tree_add_6_33_groupi_n_3346 ,csa_tree_add_6_33_groupi_n_2776 ,csa_tree_add_6_33_groupi_n_3021);
  or csa_tree_add_6_33_groupi_g15011(csa_tree_add_6_33_groupi_n_3345 ,csa_tree_add_6_33_groupi_n_2821 ,csa_tree_add_6_33_groupi_n_3099);
  not csa_tree_add_6_33_groupi_g15012(csa_tree_add_6_33_groupi_n_3288 ,csa_tree_add_6_33_groupi_n_3287);
  not csa_tree_add_6_33_groupi_g15013(csa_tree_add_6_33_groupi_n_3276 ,csa_tree_add_6_33_groupi_n_3277);
  not csa_tree_add_6_33_groupi_g15014(csa_tree_add_6_33_groupi_n_3274 ,csa_tree_add_6_33_groupi_n_3275);
  not csa_tree_add_6_33_groupi_g15015(csa_tree_add_6_33_groupi_n_3272 ,csa_tree_add_6_33_groupi_n_3273);
  not csa_tree_add_6_33_groupi_g15016(csa_tree_add_6_33_groupi_n_3267 ,csa_tree_add_6_33_groupi_n_3268);
  not csa_tree_add_6_33_groupi_g15017(csa_tree_add_6_33_groupi_n_3265 ,csa_tree_add_6_33_groupi_n_3266);
  or csa_tree_add_6_33_groupi_g15018(csa_tree_add_6_33_groupi_n_3264 ,csa_tree_add_6_33_groupi_n_2697 ,csa_tree_add_6_33_groupi_n_3040);
  or csa_tree_add_6_33_groupi_g15019(csa_tree_add_6_33_groupi_n_3263 ,csa_tree_add_6_33_groupi_n_2729 ,csa_tree_add_6_33_groupi_n_3018);
  or csa_tree_add_6_33_groupi_g15020(csa_tree_add_6_33_groupi_n_3262 ,csa_tree_add_6_33_groupi_n_2562 ,csa_tree_add_6_33_groupi_n_3131);
  or csa_tree_add_6_33_groupi_g15021(csa_tree_add_6_33_groupi_n_3261 ,csa_tree_add_6_33_groupi_n_3193 ,csa_tree_add_6_33_groupi_n_3152);
  or csa_tree_add_6_33_groupi_g15022(csa_tree_add_6_33_groupi_n_3260 ,csa_tree_add_6_33_groupi_n_3058 ,csa_tree_add_6_33_groupi_n_3013);
  or csa_tree_add_6_33_groupi_g15023(csa_tree_add_6_33_groupi_n_3259 ,csa_tree_add_6_33_groupi_n_2748 ,csa_tree_add_6_33_groupi_n_3010);
  or csa_tree_add_6_33_groupi_g15024(csa_tree_add_6_33_groupi_n_3258 ,csa_tree_add_6_33_groupi_n_2602 ,csa_tree_add_6_33_groupi_n_3053);
  or csa_tree_add_6_33_groupi_g15025(csa_tree_add_6_33_groupi_n_3257 ,csa_tree_add_6_33_groupi_n_2728 ,csa_tree_add_6_33_groupi_n_3017);
  or csa_tree_add_6_33_groupi_g15026(csa_tree_add_6_33_groupi_n_3256 ,csa_tree_add_6_33_groupi_n_2475 ,csa_tree_add_6_33_groupi_n_3004);
  nor csa_tree_add_6_33_groupi_g15027(csa_tree_add_6_33_groupi_n_3255 ,csa_tree_add_6_33_groupi_n_2601 ,csa_tree_add_6_33_groupi_n_3054);
  or csa_tree_add_6_33_groupi_g15028(csa_tree_add_6_33_groupi_n_3254 ,csa_tree_add_6_33_groupi_n_2726 ,csa_tree_add_6_33_groupi_n_3000);
  or csa_tree_add_6_33_groupi_g15029(csa_tree_add_6_33_groupi_n_3253 ,csa_tree_add_6_33_groupi_n_2476 ,csa_tree_add_6_33_groupi_n_2999);
  or csa_tree_add_6_33_groupi_g15030(csa_tree_add_6_33_groupi_n_3252 ,csa_tree_add_6_33_groupi_n_2482 ,csa_tree_add_6_33_groupi_n_2997);
  or csa_tree_add_6_33_groupi_g15031(csa_tree_add_6_33_groupi_n_3251 ,csa_tree_add_6_33_groupi_n_3057 ,csa_tree_add_6_33_groupi_n_3075);
  or csa_tree_add_6_33_groupi_g15032(csa_tree_add_6_33_groupi_n_3250 ,csa_tree_add_6_33_groupi_n_2546 ,csa_tree_add_6_33_groupi_n_2991);
  xnor csa_tree_add_6_33_groupi_g15033(csa_tree_add_6_33_groupi_n_3249 ,csa_tree_add_6_33_groupi_n_2731 ,csa_tree_add_6_33_groupi_n_2450);
  xnor csa_tree_add_6_33_groupi_g15034(csa_tree_add_6_33_groupi_n_3248 ,csa_tree_add_6_33_groupi_n_2626 ,csa_tree_add_6_33_groupi_n_2660);
  xnor csa_tree_add_6_33_groupi_g15035(csa_tree_add_6_33_groupi_n_3247 ,csa_tree_add_6_33_groupi_n_2737 ,csa_tree_add_6_33_groupi_n_2648);
  xnor csa_tree_add_6_33_groupi_g15036(csa_tree_add_6_33_groupi_n_3246 ,csa_tree_add_6_33_groupi_n_2734 ,csa_tree_add_6_33_groupi_n_2642);
  xnor csa_tree_add_6_33_groupi_g15037(csa_tree_add_6_33_groupi_n_3245 ,csa_tree_add_6_33_groupi_n_2605 ,csa_tree_add_6_33_groupi_n_2748);
  xnor csa_tree_add_6_33_groupi_g15038(csa_tree_add_6_33_groupi_n_3244 ,csa_tree_add_6_33_groupi_n_2712 ,csa_tree_add_6_33_groupi_n_2570);
  xnor csa_tree_add_6_33_groupi_g15039(csa_tree_add_6_33_groupi_n_3243 ,csa_tree_add_6_33_groupi_n_2616 ,csa_tree_add_6_33_groupi_n_2728);
  xnor csa_tree_add_6_33_groupi_g15040(csa_tree_add_6_33_groupi_n_3242 ,csa_tree_add_6_33_groupi_n_2634 ,csa_tree_add_6_33_groupi_n_2635);
  xnor csa_tree_add_6_33_groupi_g15041(csa_tree_add_6_33_groupi_n_3241 ,csa_tree_add_6_33_groupi_n_2732 ,csa_tree_add_6_33_groupi_n_2630);
  xnor csa_tree_add_6_33_groupi_g15042(csa_tree_add_6_33_groupi_n_3240 ,csa_tree_add_6_33_groupi_n_2668 ,csa_tree_add_6_33_groupi_n_2543);
  xnor csa_tree_add_6_33_groupi_g15043(csa_tree_add_6_33_groupi_n_3239 ,csa_tree_add_6_33_groupi_n_2654 ,csa_tree_add_6_33_groupi_n_2655);
  xnor csa_tree_add_6_33_groupi_g15044(csa_tree_add_6_33_groupi_n_3238 ,csa_tree_add_6_33_groupi_n_2661 ,csa_tree_add_6_33_groupi_n_2588);
  xnor csa_tree_add_6_33_groupi_g15045(csa_tree_add_6_33_groupi_n_3237 ,csa_tree_add_6_33_groupi_n_2704 ,csa_tree_add_6_33_groupi_n_2743);
  xnor csa_tree_add_6_33_groupi_g15046(csa_tree_add_6_33_groupi_n_3236 ,csa_tree_add_6_33_groupi_n_2683 ,csa_tree_add_6_33_groupi_n_2550);
  xnor csa_tree_add_6_33_groupi_g15047(csa_tree_add_6_33_groupi_n_3235 ,csa_tree_add_6_33_groupi_n_2657 ,csa_tree_add_6_33_groupi_n_2656);
  xnor csa_tree_add_6_33_groupi_g15048(csa_tree_add_6_33_groupi_n_3234 ,csa_tree_add_6_33_groupi_n_2666 ,csa_tree_add_6_33_groupi_n_2504);
  xnor csa_tree_add_6_33_groupi_g15049(csa_tree_add_6_33_groupi_n_3233 ,csa_tree_add_6_33_groupi_n_2696 ,csa_tree_add_6_33_groupi_n_2703);
  xnor csa_tree_add_6_33_groupi_g15050(csa_tree_add_6_33_groupi_n_3232 ,csa_tree_add_6_33_groupi_n_2689 ,csa_tree_add_6_33_groupi_n_2672);
  xnor csa_tree_add_6_33_groupi_g15051(csa_tree_add_6_33_groupi_n_3231 ,csa_tree_add_6_33_groupi_n_2710 ,csa_tree_add_6_33_groupi_n_2896);
  xnor csa_tree_add_6_33_groupi_g15052(csa_tree_add_6_33_groupi_n_3230 ,csa_tree_add_6_33_groupi_n_2713 ,csa_tree_add_6_33_groupi_n_2678);
  xnor csa_tree_add_6_33_groupi_g15053(csa_tree_add_6_33_groupi_n_3229 ,csa_tree_add_6_33_groupi_n_2645 ,csa_tree_add_6_33_groupi_n_2608);
  xnor csa_tree_add_6_33_groupi_g15054(csa_tree_add_6_33_groupi_n_3228 ,csa_tree_add_6_33_groupi_n_2899 ,csa_tree_add_6_33_groupi_n_2674);
  xnor csa_tree_add_6_33_groupi_g15055(csa_tree_add_6_33_groupi_n_3227 ,csa_tree_add_6_33_groupi_n_2671 ,csa_tree_add_6_33_groupi_n_2907);
  xnor csa_tree_add_6_33_groupi_g15056(csa_tree_add_6_33_groupi_n_3226 ,csa_tree_add_6_33_groupi_n_2520 ,csa_tree_add_6_33_groupi_n_2894);
  xnor csa_tree_add_6_33_groupi_g15057(csa_tree_add_6_33_groupi_n_3225 ,csa_tree_add_6_33_groupi_n_2699 ,csa_tree_add_6_33_groupi_n_2701);
  xor csa_tree_add_6_33_groupi_g15058(csa_tree_add_6_33_groupi_n_3224 ,csa_tree_add_6_33_groupi_n_2687 ,csa_tree_add_6_33_groupi_n_2754);
  xnor csa_tree_add_6_33_groupi_g15059(csa_tree_add_6_33_groupi_n_3223 ,csa_tree_add_6_33_groupi_n_2694 ,csa_tree_add_6_33_groupi_n_2641);
  xnor csa_tree_add_6_33_groupi_g15060(csa_tree_add_6_33_groupi_n_3222 ,csa_tree_add_6_33_groupi_n_2905 ,csa_tree_add_6_33_groupi_n_2752);
  xor csa_tree_add_6_33_groupi_g15061(csa_tree_add_6_33_groupi_n_3221 ,csa_tree_add_6_33_groupi_n_2723 ,csa_tree_add_6_33_groupi_n_2514);
  xnor csa_tree_add_6_33_groupi_g15062(csa_tree_add_6_33_groupi_n_3220 ,csa_tree_add_6_33_groupi_n_2679 ,csa_tree_add_6_33_groupi_n_2386);
  xnor csa_tree_add_6_33_groupi_g15063(csa_tree_add_6_33_groupi_n_3219 ,csa_tree_add_6_33_groupi_n_2638 ,csa_tree_add_6_33_groupi_n_2729);
  xnor csa_tree_add_6_33_groupi_g15064(csa_tree_add_6_33_groupi_n_3218 ,csa_tree_add_6_33_groupi_n_2426 ,csa_tree_add_6_33_groupi_n_2706);
  xnor csa_tree_add_6_33_groupi_g15065(csa_tree_add_6_33_groupi_n_3217 ,csa_tree_add_6_33_groupi_n_2711 ,csa_tree_add_6_33_groupi_n_2888);
  xnor csa_tree_add_6_33_groupi_g15066(csa_tree_add_6_33_groupi_n_3216 ,csa_tree_add_6_33_groupi_n_2900 ,csa_tree_add_6_33_groupi_n_2686);
  xnor csa_tree_add_6_33_groupi_g15067(csa_tree_add_6_33_groupi_n_3215 ,csa_tree_add_6_33_groupi_n_2911 ,csa_tree_add_6_33_groupi_n_2691);
  xnor csa_tree_add_6_33_groupi_g15068(csa_tree_add_6_33_groupi_n_3214 ,csa_tree_add_6_33_groupi_n_2909 ,csa_tree_add_6_33_groupi_n_2625);
  xnor csa_tree_add_6_33_groupi_g15069(csa_tree_add_6_33_groupi_n_3213 ,csa_tree_add_6_33_groupi_n_2700 ,csa_tree_add_6_33_groupi_n_2594);
  xnor csa_tree_add_6_33_groupi_g15070(csa_tree_add_6_33_groupi_n_3212 ,csa_tree_add_6_33_groupi_n_2726 ,csa_tree_add_6_33_groupi_n_2335);
  xnor csa_tree_add_6_33_groupi_g15071(csa_tree_add_6_33_groupi_n_3211 ,csa_tree_add_6_33_groupi_n_2591 ,csa_tree_add_6_33_groupi_n_2592);
  xnor csa_tree_add_6_33_groupi_g15072(csa_tree_add_6_33_groupi_n_3210 ,csa_tree_add_6_33_groupi_n_2603 ,csa_tree_add_6_33_groupi_n_2476);
  xnor csa_tree_add_6_33_groupi_g15073(csa_tree_add_6_33_groupi_n_3209 ,csa_tree_add_6_33_groupi_n_2610 ,csa_tree_add_6_33_groupi_n_2612);
  xnor csa_tree_add_6_33_groupi_g15074(csa_tree_add_6_33_groupi_n_3208 ,csa_tree_add_6_33_groupi_n_2598 ,csa_tree_add_6_33_groupi_n_2482);
  xnor csa_tree_add_6_33_groupi_g15075(csa_tree_add_6_33_groupi_n_3207 ,csa_tree_add_6_33_groupi_n_2627 ,csa_tree_add_6_33_groupi_n_2595);
  xnor csa_tree_add_6_33_groupi_g15076(csa_tree_add_6_33_groupi_n_3206 ,csa_tree_add_6_33_groupi_n_2646 ,csa_tree_add_6_33_groupi_n_2549);
  xnor csa_tree_add_6_33_groupi_g15077(csa_tree_add_6_33_groupi_n_3205 ,csa_tree_add_6_33_groupi_n_2633 ,csa_tree_add_6_33_groupi_n_2572);
  xnor csa_tree_add_6_33_groupi_g15078(csa_tree_add_6_33_groupi_n_3204 ,csa_tree_add_6_33_groupi_n_2615 ,csa_tree_add_6_33_groupi_n_2628);
  xnor csa_tree_add_6_33_groupi_g15079(csa_tree_add_6_33_groupi_n_3203 ,csa_tree_add_6_33_groupi_n_2600 ,csa_tree_add_6_33_groupi_n_2437);
  xnor csa_tree_add_6_33_groupi_g15080(csa_tree_add_6_33_groupi_n_3202 ,csa_tree_add_6_33_groupi_n_2720 ,csa_tree_add_6_33_groupi_n_2722);
  xnor csa_tree_add_6_33_groupi_g15081(csa_tree_add_6_33_groupi_n_3201 ,csa_tree_add_6_33_groupi_n_2707 ,csa_tree_add_6_33_groupi_n_2636);
  xnor csa_tree_add_6_33_groupi_g15082(csa_tree_add_6_33_groupi_n_3200 ,csa_tree_add_6_33_groupi_n_2750 ,csa_tree_add_6_33_groupi_n_2521);
  xnor csa_tree_add_6_33_groupi_g15083(csa_tree_add_6_33_groupi_n_3199 ,csa_tree_add_6_33_groupi_n_2590 ,csa_tree_add_6_33_groupi_n_2669);
  xnor csa_tree_add_6_33_groupi_g15084(csa_tree_add_6_33_groupi_n_3198 ,csa_tree_add_6_33_groupi_n_2652 ,csa_tree_add_6_33_groupi_n_2663);
  xnor csa_tree_add_6_33_groupi_g15085(csa_tree_add_6_33_groupi_n_3197 ,csa_tree_add_6_33_groupi_n_2719 ,csa_tree_add_6_33_groupi_n_2721);
  xnor csa_tree_add_6_33_groupi_g15086(csa_tree_add_6_33_groupi_n_3196 ,csa_tree_add_6_33_groupi_n_2677 ,csa_tree_add_6_33_groupi_n_2502);
  and csa_tree_add_6_33_groupi_g15087(csa_tree_add_6_33_groupi_n_3292 ,csa_tree_add_6_33_groupi_n_2852 ,csa_tree_add_6_33_groupi_n_2988);
  and csa_tree_add_6_33_groupi_g15088(csa_tree_add_6_33_groupi_n_3291 ,csa_tree_add_6_33_groupi_n_2774 ,csa_tree_add_6_33_groupi_n_3016);
  and csa_tree_add_6_33_groupi_g15089(csa_tree_add_6_33_groupi_n_3290 ,csa_tree_add_6_33_groupi_n_2770 ,csa_tree_add_6_33_groupi_n_3014);
  and csa_tree_add_6_33_groupi_g15090(csa_tree_add_6_33_groupi_n_3289 ,csa_tree_add_6_33_groupi_n_2858 ,csa_tree_add_6_33_groupi_n_3006);
  xnor csa_tree_add_6_33_groupi_g15091(csa_tree_add_6_33_groupi_n_3287 ,csa_tree_add_6_33_groupi_n_2548 ,csa_tree_add_6_33_groupi_n_2756);
  and csa_tree_add_6_33_groupi_g15092(csa_tree_add_6_33_groupi_n_3286 ,csa_tree_add_6_33_groupi_n_2766 ,csa_tree_add_6_33_groupi_n_3005);
  and csa_tree_add_6_33_groupi_g15093(csa_tree_add_6_33_groupi_n_3285 ,csa_tree_add_6_33_groupi_n_2763 ,csa_tree_add_6_33_groupi_n_3003);
  and csa_tree_add_6_33_groupi_g15094(csa_tree_add_6_33_groupi_n_3284 ,csa_tree_add_6_33_groupi_n_2844 ,csa_tree_add_6_33_groupi_n_2981);
  and csa_tree_add_6_33_groupi_g15095(csa_tree_add_6_33_groupi_n_3283 ,csa_tree_add_6_33_groupi_n_2761 ,csa_tree_add_6_33_groupi_n_2998);
  and csa_tree_add_6_33_groupi_g15096(csa_tree_add_6_33_groupi_n_3282 ,csa_tree_add_6_33_groupi_n_2829 ,csa_tree_add_6_33_groupi_n_2985);
  and csa_tree_add_6_33_groupi_g15097(csa_tree_add_6_33_groupi_n_3281 ,csa_tree_add_6_33_groupi_n_2881 ,csa_tree_add_6_33_groupi_n_3184);
  and csa_tree_add_6_33_groupi_g15098(csa_tree_add_6_33_groupi_n_3280 ,csa_tree_add_6_33_groupi_n_2851 ,csa_tree_add_6_33_groupi_n_3181);
  and csa_tree_add_6_33_groupi_g15099(csa_tree_add_6_33_groupi_n_3279 ,csa_tree_add_6_33_groupi_n_2842 ,csa_tree_add_6_33_groupi_n_2989);
  xnor csa_tree_add_6_33_groupi_g15100(csa_tree_add_6_33_groupi_n_3278 ,csa_tree_add_6_33_groupi_n_2402 ,csa_tree_add_6_33_groupi_n_2585);
  or csa_tree_add_6_33_groupi_g15101(csa_tree_add_6_33_groupi_n_3277 ,csa_tree_add_6_33_groupi_n_2866 ,csa_tree_add_6_33_groupi_n_2984);
  or csa_tree_add_6_33_groupi_g15102(csa_tree_add_6_33_groupi_n_3275 ,csa_tree_add_6_33_groupi_n_2793 ,csa_tree_add_6_33_groupi_n_2980);
  xnor csa_tree_add_6_33_groupi_g15103(csa_tree_add_6_33_groupi_n_3273 ,csa_tree_add_6_33_groupi_n_2392 ,csa_tree_add_6_33_groupi_n_2757);
  xnor csa_tree_add_6_33_groupi_g15104(csa_tree_add_6_33_groupi_n_3271 ,csa_tree_add_6_33_groupi_n_2389 ,csa_tree_add_6_33_groupi_n_2583);
  or csa_tree_add_6_33_groupi_g15105(csa_tree_add_6_33_groupi_n_3270 ,csa_tree_add_6_33_groupi_n_2835 ,csa_tree_add_6_33_groupi_n_3108);
  and csa_tree_add_6_33_groupi_g15106(csa_tree_add_6_33_groupi_n_3269 ,csa_tree_add_6_33_groupi_n_2855 ,csa_tree_add_6_33_groupi_n_3124);
  xnor csa_tree_add_6_33_groupi_g15107(csa_tree_add_6_33_groupi_n_3268 ,csa_tree_add_6_33_groupi_n_2480 ,csa_tree_add_6_33_groupi_n_2586);
  xnor csa_tree_add_6_33_groupi_g15108(csa_tree_add_6_33_groupi_n_3266 ,csa_tree_add_6_33_groupi_n_2557 ,csa_tree_add_6_33_groupi_n_2584);
  or csa_tree_add_6_33_groupi_g15109(csa_tree_add_6_33_groupi_n_3184 ,csa_tree_add_6_33_groupi_n_2575 ,csa_tree_add_6_33_groupi_n_2813);
  and csa_tree_add_6_33_groupi_g15110(csa_tree_add_6_33_groupi_n_3183 ,csa_tree_add_6_33_groupi_n_2327 ,csa_tree_add_6_33_groupi_n_2688);
  and csa_tree_add_6_33_groupi_g15111(csa_tree_add_6_33_groupi_n_3182 ,csa_tree_add_6_33_groupi_n_2685 ,csa_tree_add_6_33_groupi_n_2712);
  or csa_tree_add_6_33_groupi_g15112(csa_tree_add_6_33_groupi_n_3181 ,csa_tree_add_6_33_groupi_n_2554 ,csa_tree_add_6_33_groupi_n_2877);
  nor csa_tree_add_6_33_groupi_g15113(csa_tree_add_6_33_groupi_n_3180 ,csa_tree_add_6_33_groupi_n_877 ,csa_tree_add_6_33_groupi_n_2590);
  or csa_tree_add_6_33_groupi_g15114(csa_tree_add_6_33_groupi_n_3179 ,csa_tree_add_6_33_groupi_n_2663 ,csa_tree_add_6_33_groupi_n_2652);
  or csa_tree_add_6_33_groupi_g15115(csa_tree_add_6_33_groupi_n_3178 ,csa_tree_add_6_33_groupi_n_1006 ,csa_tree_add_6_33_groupi_n_2589);
  or csa_tree_add_6_33_groupi_g15116(csa_tree_add_6_33_groupi_n_3177 ,csa_tree_add_6_33_groupi_n_2568 ,csa_tree_add_6_33_groupi_n_2883);
  or csa_tree_add_6_33_groupi_g15117(csa_tree_add_6_33_groupi_n_3176 ,csa_tree_add_6_33_groupi_n_2649 ,csa_tree_add_6_33_groupi_n_2646);
  or csa_tree_add_6_33_groupi_g15118(csa_tree_add_6_33_groupi_n_3175 ,csa_tree_add_6_33_groupi_n_2904 ,csa_tree_add_6_33_groupi_n_2644);
  and csa_tree_add_6_33_groupi_g15119(csa_tree_add_6_33_groupi_n_3174 ,csa_tree_add_6_33_groupi_n_2649 ,csa_tree_add_6_33_groupi_n_2646);
  or csa_tree_add_6_33_groupi_g15120(csa_tree_add_6_33_groupi_n_3173 ,csa_tree_add_6_33_groupi_n_2531 ,csa_tree_add_6_33_groupi_n_2622);
  and csa_tree_add_6_33_groupi_g15121(csa_tree_add_6_33_groupi_n_3172 ,csa_tree_add_6_33_groupi_n_2663 ,csa_tree_add_6_33_groupi_n_2652);
  nor csa_tree_add_6_33_groupi_g15122(csa_tree_add_6_33_groupi_n_3171 ,csa_tree_add_6_33_groupi_n_2905 ,csa_tree_add_6_33_groupi_n_2643);
  or csa_tree_add_6_33_groupi_g15123(csa_tree_add_6_33_groupi_n_3170 ,csa_tree_add_6_33_groupi_n_2636 ,csa_tree_add_6_33_groupi_n_2707);
  nor csa_tree_add_6_33_groupi_g15124(csa_tree_add_6_33_groupi_n_3169 ,csa_tree_add_6_33_groupi_n_2542 ,csa_tree_add_6_33_groupi_n_2880);
  and csa_tree_add_6_33_groupi_g15125(csa_tree_add_6_33_groupi_n_3168 ,csa_tree_add_6_33_groupi_n_2636 ,csa_tree_add_6_33_groupi_n_2707);
  or csa_tree_add_6_33_groupi_g15126(csa_tree_add_6_33_groupi_n_3167 ,csa_tree_add_6_33_groupi_n_2633 ,csa_tree_add_6_33_groupi_n_2620);
  or csa_tree_add_6_33_groupi_g15127(csa_tree_add_6_33_groupi_n_3166 ,csa_tree_add_6_33_groupi_n_2628 ,csa_tree_add_6_33_groupi_n_2615);
  and csa_tree_add_6_33_groupi_g15128(csa_tree_add_6_33_groupi_n_3165 ,csa_tree_add_6_33_groupi_n_2633 ,csa_tree_add_6_33_groupi_n_2620);
  and csa_tree_add_6_33_groupi_g15129(csa_tree_add_6_33_groupi_n_3164 ,csa_tree_add_6_33_groupi_n_2628 ,csa_tree_add_6_33_groupi_n_2615);
  or csa_tree_add_6_33_groupi_g15130(csa_tree_add_6_33_groupi_n_3163 ,csa_tree_add_6_33_groupi_n_2825 ,csa_tree_add_6_33_groupi_n_2741);
  or csa_tree_add_6_33_groupi_g15131(csa_tree_add_6_33_groupi_n_3162 ,csa_tree_add_6_33_groupi_n_2582 ,csa_tree_add_6_33_groupi_n_2786);
  or csa_tree_add_6_33_groupi_g15132(csa_tree_add_6_33_groupi_n_3161 ,csa_tree_add_6_33_groupi_n_2363 ,csa_tree_add_6_33_groupi_n_2785);
  or csa_tree_add_6_33_groupi_g15133(csa_tree_add_6_33_groupi_n_3160 ,csa_tree_add_6_33_groupi_n_2494 ,csa_tree_add_6_33_groupi_n_2596);
  and csa_tree_add_6_33_groupi_g15134(csa_tree_add_6_33_groupi_n_3159 ,csa_tree_add_6_33_groupi_n_2531 ,csa_tree_add_6_33_groupi_n_2622);
  and csa_tree_add_6_33_groupi_g15135(csa_tree_add_6_33_groupi_n_3158 ,csa_tree_add_6_33_groupi_n_2500 ,csa_tree_add_6_33_groupi_n_2611);
  and csa_tree_add_6_33_groupi_g15136(csa_tree_add_6_33_groupi_n_3157 ,csa_tree_add_6_33_groupi_n_2504 ,csa_tree_add_6_33_groupi_n_2666);
  and csa_tree_add_6_33_groupi_g15137(csa_tree_add_6_33_groupi_n_3156 ,csa_tree_add_6_33_groupi_n_2494 ,csa_tree_add_6_33_groupi_n_2596);
  or csa_tree_add_6_33_groupi_g15138(csa_tree_add_6_33_groupi_n_3155 ,csa_tree_add_6_33_groupi_n_2630 ,csa_tree_add_6_33_groupi_n_2629);
  or csa_tree_add_6_33_groupi_g15139(csa_tree_add_6_33_groupi_n_3154 ,csa_tree_add_6_33_groupi_n_2579 ,csa_tree_add_6_33_groupi_n_2872);
  nor csa_tree_add_6_33_groupi_g15140(csa_tree_add_6_33_groupi_n_3153 ,csa_tree_add_6_33_groupi_n_2519 ,csa_tree_add_6_33_groupi_n_2894);
  and csa_tree_add_6_33_groupi_g15141(csa_tree_add_6_33_groupi_n_3152 ,csa_tree_add_6_33_groupi_n_2502 ,csa_tree_add_6_33_groupi_n_2677);
  or csa_tree_add_6_33_groupi_g15142(csa_tree_add_6_33_groupi_n_3151 ,csa_tree_add_6_33_groupi_n_2722 ,csa_tree_add_6_33_groupi_n_2720);
  or csa_tree_add_6_33_groupi_g15143(csa_tree_add_6_33_groupi_n_3150 ,csa_tree_add_6_33_groupi_n_2721 ,csa_tree_add_6_33_groupi_n_2719);
  or csa_tree_add_6_33_groupi_g15144(csa_tree_add_6_33_groupi_n_3149 ,csa_tree_add_6_33_groupi_n_2898 ,csa_tree_add_6_33_groupi_n_2674);
  and csa_tree_add_6_33_groupi_g15145(csa_tree_add_6_33_groupi_n_3148 ,csa_tree_add_6_33_groupi_n_2722 ,csa_tree_add_6_33_groupi_n_2720);
  or csa_tree_add_6_33_groupi_g15146(csa_tree_add_6_33_groupi_n_3147 ,csa_tree_add_6_33_groupi_n_2555 ,csa_tree_add_6_33_groupi_n_2868);
  or csa_tree_add_6_33_groupi_g15147(csa_tree_add_6_33_groupi_n_3146 ,csa_tree_add_6_33_groupi_n_2521 ,csa_tree_add_6_33_groupi_n_2716);
  and csa_tree_add_6_33_groupi_g15148(csa_tree_add_6_33_groupi_n_3145 ,csa_tree_add_6_33_groupi_n_2521 ,csa_tree_add_6_33_groupi_n_2716);
  or csa_tree_add_6_33_groupi_g15149(csa_tree_add_6_33_groupi_n_3144 ,csa_tree_add_6_33_groupi_n_2471 ,csa_tree_add_6_33_groupi_n_2862);
  or csa_tree_add_6_33_groupi_g15150(csa_tree_add_6_33_groupi_n_3143 ,csa_tree_add_6_33_groupi_n_2888 ,csa_tree_add_6_33_groupi_n_2711);
  or csa_tree_add_6_33_groupi_g15151(csa_tree_add_6_33_groupi_n_3142 ,csa_tree_add_6_33_groupi_n_2685 ,csa_tree_add_6_33_groupi_n_2712);
  and csa_tree_add_6_33_groupi_g15152(csa_tree_add_6_33_groupi_n_3141 ,csa_tree_add_6_33_groupi_n_2888 ,csa_tree_add_6_33_groupi_n_2711);
  or csa_tree_add_6_33_groupi_g15153(csa_tree_add_6_33_groupi_n_3140 ,csa_tree_add_6_33_groupi_n_2567 ,csa_tree_add_6_33_groupi_n_2860);
  nor csa_tree_add_6_33_groupi_g15154(csa_tree_add_6_33_groupi_n_3139 ,csa_tree_add_6_33_groupi_n_2899 ,csa_tree_add_6_33_groupi_n_2673);
  or csa_tree_add_6_33_groupi_g15155(csa_tree_add_6_33_groupi_n_3138 ,csa_tree_add_6_33_groupi_n_2695 ,csa_tree_add_6_33_groupi_n_2703);
  or csa_tree_add_6_33_groupi_g15156(csa_tree_add_6_33_groupi_n_3137 ,csa_tree_add_6_33_groupi_n_2566 ,csa_tree_add_6_33_groupi_n_2795);
  or csa_tree_add_6_33_groupi_g15157(csa_tree_add_6_33_groupi_n_3136 ,csa_tree_add_6_33_groupi_n_2520 ,csa_tree_add_6_33_groupi_n_2893);
  nor csa_tree_add_6_33_groupi_g15158(csa_tree_add_6_33_groupi_n_3135 ,csa_tree_add_6_33_groupi_n_2710 ,csa_tree_add_6_33_groupi_n_2895);
  or csa_tree_add_6_33_groupi_g15159(csa_tree_add_6_33_groupi_n_3134 ,csa_tree_add_6_33_groupi_n_2708 ,csa_tree_add_6_33_groupi_n_2704);
  nor csa_tree_add_6_33_groupi_g15160(csa_tree_add_6_33_groupi_n_3133 ,csa_tree_add_6_33_groupi_n_2565 ,csa_tree_add_6_33_groupi_n_2886);
  or csa_tree_add_6_33_groupi_g15161(csa_tree_add_6_33_groupi_n_3132 ,csa_tree_add_6_33_groupi_n_2709 ,csa_tree_add_6_33_groupi_n_2896);
  nor csa_tree_add_6_33_groupi_g15162(csa_tree_add_6_33_groupi_n_3131 ,csa_tree_add_6_33_groupi_n_1397 ,csa_tree_add_6_33_groupi_n_2718);
  and csa_tree_add_6_33_groupi_g15163(csa_tree_add_6_33_groupi_n_3130 ,csa_tree_add_6_33_groupi_n_2708 ,csa_tree_add_6_33_groupi_n_2704);
  or csa_tree_add_6_33_groupi_g15164(csa_tree_add_6_33_groupi_n_3129 ,csa_tree_add_6_33_groupi_n_2701 ,csa_tree_add_6_33_groupi_n_2699);
  or csa_tree_add_6_33_groupi_g15165(csa_tree_add_6_33_groupi_n_3128 ,csa_tree_add_6_33_groupi_n_2462 ,csa_tree_add_6_33_groupi_n_2789);
  and csa_tree_add_6_33_groupi_g15166(csa_tree_add_6_33_groupi_n_3127 ,csa_tree_add_6_33_groupi_n_2594 ,csa_tree_add_6_33_groupi_n_2700);
  and csa_tree_add_6_33_groupi_g15167(csa_tree_add_6_33_groupi_n_3126 ,csa_tree_add_6_33_groupi_n_2701 ,csa_tree_add_6_33_groupi_n_2699);
  and csa_tree_add_6_33_groupi_g15168(csa_tree_add_6_33_groupi_n_3125 ,csa_tree_add_6_33_groupi_n_2386 ,csa_tree_add_6_33_groupi_n_2679);
  or csa_tree_add_6_33_groupi_g15169(csa_tree_add_6_33_groupi_n_3124 ,csa_tree_add_6_33_groupi_n_2850 ,csa_tree_add_6_33_groupi_n_2747);
  nor csa_tree_add_6_33_groupi_g15170(csa_tree_add_6_33_groupi_n_3123 ,csa_tree_add_6_33_groupi_n_2696 ,csa_tree_add_6_33_groupi_n_2702);
  or csa_tree_add_6_33_groupi_g15171(csa_tree_add_6_33_groupi_n_3122 ,csa_tree_add_6_33_groupi_n_2746 ,csa_tree_add_6_33_groupi_n_2847);
  or csa_tree_add_6_33_groupi_g15172(csa_tree_add_6_33_groupi_n_3121 ,csa_tree_add_6_33_groupi_n_2560 ,csa_tree_add_6_33_groupi_n_2759);
  or csa_tree_add_6_33_groupi_g15173(csa_tree_add_6_33_groupi_n_3120 ,csa_tree_add_6_33_groupi_n_2502 ,csa_tree_add_6_33_groupi_n_2677);
  or csa_tree_add_6_33_groupi_g15174(csa_tree_add_6_33_groupi_n_3119 ,csa_tree_add_6_33_groupi_n_2675 ,csa_tree_add_6_33_groupi_n_2687);
  or csa_tree_add_6_33_groupi_g15175(csa_tree_add_6_33_groupi_n_3118 ,csa_tree_add_6_33_groupi_n_2539 ,csa_tree_add_6_33_groupi_n_2875);
  and csa_tree_add_6_33_groupi_g15176(csa_tree_add_6_33_groupi_n_3117 ,csa_tree_add_6_33_groupi_n_2672 ,csa_tree_add_6_33_groupi_n_2689);
  nor csa_tree_add_6_33_groupi_g15177(csa_tree_add_6_33_groupi_n_3116 ,csa_tree_add_6_33_groupi_n_2901 ,csa_tree_add_6_33_groupi_n_2686);
  or csa_tree_add_6_33_groupi_g15178(csa_tree_add_6_33_groupi_n_3115 ,csa_tree_add_6_33_groupi_n_2500 ,csa_tree_add_6_33_groupi_n_2611);
  or csa_tree_add_6_33_groupi_g15179(csa_tree_add_6_33_groupi_n_3114 ,csa_tree_add_6_33_groupi_n_2544 ,csa_tree_add_6_33_groupi_n_2845);
  and csa_tree_add_6_33_groupi_g15180(csa_tree_add_6_33_groupi_n_3113 ,csa_tree_add_6_33_groupi_n_2675 ,csa_tree_add_6_33_groupi_n_2687);
  and csa_tree_add_6_33_groupi_g15181(csa_tree_add_6_33_groupi_n_3112 ,csa_tree_add_6_33_groupi_n_2819 ,csa_tree_add_6_33_groupi_n_2739);
  nor csa_tree_add_6_33_groupi_g15182(csa_tree_add_6_33_groupi_n_3111 ,csa_tree_add_6_33_groupi_n_2837 ,csa_tree_add_6_33_groupi_n_2745);
  or csa_tree_add_6_33_groupi_g15183(csa_tree_add_6_33_groupi_n_3110 ,csa_tree_add_6_33_groupi_n_2551 ,csa_tree_add_6_33_groupi_n_2833);
  or csa_tree_add_6_33_groupi_g15184(csa_tree_add_6_33_groupi_n_3109 ,csa_tree_add_6_33_groupi_n_2684 ,csa_tree_add_6_33_groupi_n_2683);
  and csa_tree_add_6_33_groupi_g15185(csa_tree_add_6_33_groupi_n_3108 ,csa_tree_add_6_33_groupi_n_2352 ,csa_tree_add_6_33_groupi_n_2834);
  or csa_tree_add_6_33_groupi_g15186(csa_tree_add_6_33_groupi_n_3107 ,csa_tree_add_6_33_groupi_n_2465 ,csa_tree_add_6_33_groupi_n_2790);
  and csa_tree_add_6_33_groupi_g15187(csa_tree_add_6_33_groupi_n_3106 ,csa_tree_add_6_33_groupi_n_2684 ,csa_tree_add_6_33_groupi_n_2683);
  or csa_tree_add_6_33_groupi_g15188(csa_tree_add_6_33_groupi_n_3105 ,csa_tree_add_6_33_groupi_n_2553 ,csa_tree_add_6_33_groupi_n_2820);
  and csa_tree_add_6_33_groupi_g15189(csa_tree_add_6_33_groupi_n_3104 ,csa_tree_add_6_33_groupi_n_2608 ,csa_tree_add_6_33_groupi_n_2645);
  or csa_tree_add_6_33_groupi_g15190(csa_tree_add_6_33_groupi_n_3103 ,csa_tree_add_6_33_groupi_n_2518 ,csa_tree_add_6_33_groupi_n_2662);
  or csa_tree_add_6_33_groupi_g15191(csa_tree_add_6_33_groupi_n_3102 ,csa_tree_add_6_33_groupi_n_2386 ,csa_tree_add_6_33_groupi_n_2679);
  or csa_tree_add_6_33_groupi_g15192(csa_tree_add_6_33_groupi_n_3101 ,csa_tree_add_6_33_groupi_n_2672 ,csa_tree_add_6_33_groupi_n_2689);
  or csa_tree_add_6_33_groupi_g15193(csa_tree_add_6_33_groupi_n_3100 ,csa_tree_add_6_33_groupi_n_2547 ,csa_tree_add_6_33_groupi_n_2823);
  nor csa_tree_add_6_33_groupi_g15194(csa_tree_add_6_33_groupi_n_3099 ,csa_tree_add_6_33_groupi_n_2545 ,csa_tree_add_6_33_groupi_n_2815);
  or csa_tree_add_6_33_groupi_g15195(csa_tree_add_6_33_groupi_n_3098 ,csa_tree_add_6_33_groupi_n_2671 ,csa_tree_add_6_33_groupi_n_2906);
  or csa_tree_add_6_33_groupi_g15196(csa_tree_add_6_33_groupi_n_3097 ,csa_tree_add_6_33_groupi_n_2540 ,csa_tree_add_6_33_groupi_n_2814);
  or csa_tree_add_6_33_groupi_g15197(csa_tree_add_6_33_groupi_n_3096 ,csa_tree_add_6_33_groupi_n_2574 ,csa_tree_add_6_33_groupi_n_2859);
  or csa_tree_add_6_33_groupi_g15198(csa_tree_add_6_33_groupi_n_3095 ,csa_tree_add_6_33_groupi_n_2714 ,csa_tree_add_6_33_groupi_n_2668);
  or csa_tree_add_6_33_groupi_g15199(csa_tree_add_6_33_groupi_n_3094 ,csa_tree_add_6_33_groupi_n_2458 ,csa_tree_add_6_33_groupi_n_2768);
  or csa_tree_add_6_33_groupi_g15200(csa_tree_add_6_33_groupi_n_3093 ,csa_tree_add_6_33_groupi_n_2608 ,csa_tree_add_6_33_groupi_n_2645);
  and csa_tree_add_6_33_groupi_g15201(csa_tree_add_6_33_groupi_n_3092 ,csa_tree_add_6_33_groupi_n_2642 ,csa_tree_add_6_33_groupi_n_2639);
  nor csa_tree_add_6_33_groupi_g15202(csa_tree_add_6_33_groupi_n_3091 ,csa_tree_add_6_33_groupi_n_2670 ,csa_tree_add_6_33_groupi_n_2907);
  or csa_tree_add_6_33_groupi_g15203(csa_tree_add_6_33_groupi_n_3090 ,csa_tree_add_6_33_groupi_n_2514 ,csa_tree_add_6_33_groupi_n_2658);
  and csa_tree_add_6_33_groupi_g15204(csa_tree_add_6_33_groupi_n_3089 ,csa_tree_add_6_33_groupi_n_2518 ,csa_tree_add_6_33_groupi_n_2662);
  and csa_tree_add_6_33_groupi_g15205(csa_tree_add_6_33_groupi_n_3088 ,csa_tree_add_6_33_groupi_n_2721 ,csa_tree_add_6_33_groupi_n_2719);
  nor csa_tree_add_6_33_groupi_g15206(csa_tree_add_6_33_groupi_n_3087 ,csa_tree_add_6_33_groupi_n_2715 ,csa_tree_add_6_33_groupi_n_2667);
  nor csa_tree_add_6_33_groupi_g15207(csa_tree_add_6_33_groupi_n_3086 ,csa_tree_add_6_33_groupi_n_2588 ,csa_tree_add_6_33_groupi_n_2661);
  and csa_tree_add_6_33_groupi_g15208(csa_tree_add_6_33_groupi_n_3085 ,csa_tree_add_6_33_groupi_n_2635 ,csa_tree_add_6_33_groupi_n_2634);
  or csa_tree_add_6_33_groupi_g15209(csa_tree_add_6_33_groupi_n_3084 ,csa_tree_add_6_33_groupi_n_2635 ,csa_tree_add_6_33_groupi_n_2634);
  nor csa_tree_add_6_33_groupi_g15210(csa_tree_add_6_33_groupi_n_3083 ,csa_tree_add_6_33_groupi_n_2694 ,csa_tree_add_6_33_groupi_n_2640);
  and csa_tree_add_6_33_groupi_g15211(csa_tree_add_6_33_groupi_n_3082 ,csa_tree_add_6_33_groupi_n_2588 ,csa_tree_add_6_33_groupi_n_2661);
  nor csa_tree_add_6_33_groupi_g15212(csa_tree_add_6_33_groupi_n_3081 ,csa_tree_add_6_33_groupi_n_2425 ,csa_tree_add_6_33_groupi_n_2706);
  or csa_tree_add_6_33_groupi_g15213(csa_tree_add_6_33_groupi_n_3080 ,csa_tree_add_6_33_groupi_n_2472 ,csa_tree_add_6_33_groupi_n_2809);
  or csa_tree_add_6_33_groupi_g15214(csa_tree_add_6_33_groupi_n_3079 ,csa_tree_add_6_33_groupi_n_2655 ,csa_tree_add_6_33_groupi_n_2654);
  and csa_tree_add_6_33_groupi_g15215(csa_tree_add_6_33_groupi_n_3078 ,csa_tree_add_6_33_groupi_n_2655 ,csa_tree_add_6_33_groupi_n_2654);
  or csa_tree_add_6_33_groupi_g15216(csa_tree_add_6_33_groupi_n_3077 ,csa_tree_add_6_33_groupi_n_2484 ,csa_tree_add_6_33_groupi_n_2803);
  or csa_tree_add_6_33_groupi_g15217(csa_tree_add_6_33_groupi_n_3076 ,csa_tree_add_6_33_groupi_n_2738 ,csa_tree_add_6_33_groupi_n_2805);
  and csa_tree_add_6_33_groupi_g15218(csa_tree_add_6_33_groupi_n_3075 ,csa_tree_add_6_33_groupi_n_2595 ,csa_tree_add_6_33_groupi_n_2627);
  or csa_tree_add_6_33_groupi_g15219(csa_tree_add_6_33_groupi_n_3074 ,csa_tree_add_6_33_groupi_n_2481 ,csa_tree_add_6_33_groupi_n_2802);
  or csa_tree_add_6_33_groupi_g15220(csa_tree_add_6_33_groupi_n_3073 ,csa_tree_add_6_33_groupi_n_2648 ,csa_tree_add_6_33_groupi_n_2647);
  or csa_tree_add_6_33_groupi_g15221(csa_tree_add_6_33_groupi_n_3072 ,csa_tree_add_6_33_groupi_n_2426 ,csa_tree_add_6_33_groupi_n_2705);
  or csa_tree_add_6_33_groupi_g15222(csa_tree_add_6_33_groupi_n_3071 ,csa_tree_add_6_33_groupi_n_2656 ,csa_tree_add_6_33_groupi_n_2657);
  and csa_tree_add_6_33_groupi_g15223(csa_tree_add_6_33_groupi_n_3070 ,csa_tree_add_6_33_groupi_n_2656 ,csa_tree_add_6_33_groupi_n_2657);
  and csa_tree_add_6_33_groupi_g15224(csa_tree_add_6_33_groupi_n_3069 ,csa_tree_add_6_33_groupi_n_2648 ,csa_tree_add_6_33_groupi_n_2647);
  or csa_tree_add_6_33_groupi_g15225(csa_tree_add_6_33_groupi_n_3068 ,csa_tree_add_6_33_groupi_n_2477 ,csa_tree_add_6_33_groupi_n_2800);
  or csa_tree_add_6_33_groupi_g15226(csa_tree_add_6_33_groupi_n_3067 ,csa_tree_add_6_33_groupi_n_2581 ,csa_tree_add_6_33_groupi_n_2797);
  or csa_tree_add_6_33_groupi_g15227(csa_tree_add_6_33_groupi_n_3066 ,csa_tree_add_6_33_groupi_n_2556 ,csa_tree_add_6_33_groupi_n_2796);
  or csa_tree_add_6_33_groupi_g15228(csa_tree_add_6_33_groupi_n_3065 ,csa_tree_add_6_33_groupi_n_2470 ,csa_tree_add_6_33_groupi_n_2846);
  or csa_tree_add_6_33_groupi_g15229(csa_tree_add_6_33_groupi_n_3064 ,csa_tree_add_6_33_groupi_n_2678 ,csa_tree_add_6_33_groupi_n_2713);
  or csa_tree_add_6_33_groupi_g15230(csa_tree_add_6_33_groupi_n_3063 ,csa_tree_add_6_33_groupi_n_2642 ,csa_tree_add_6_33_groupi_n_2639);
  or csa_tree_add_6_33_groupi_g15231(csa_tree_add_6_33_groupi_n_3062 ,csa_tree_add_6_33_groupi_n_2693 ,csa_tree_add_6_33_groupi_n_2641);
  or csa_tree_add_6_33_groupi_g15232(csa_tree_add_6_33_groupi_n_3061 ,csa_tree_add_6_33_groupi_n_2504 ,csa_tree_add_6_33_groupi_n_2666);
  and csa_tree_add_6_33_groupi_g15233(csa_tree_add_6_33_groupi_n_3060 ,csa_tree_add_6_33_groupi_n_2514 ,csa_tree_add_6_33_groupi_n_2658);
  and csa_tree_add_6_33_groupi_g15234(csa_tree_add_6_33_groupi_n_3195 ,csa_tree_add_6_33_groupi_n_1808 ,csa_tree_add_6_33_groupi_n_2811);
  and csa_tree_add_6_33_groupi_g15235(csa_tree_add_6_33_groupi_n_3194 ,csa_tree_add_6_33_groupi_n_1810 ,csa_tree_add_6_33_groupi_n_2887);
  and csa_tree_add_6_33_groupi_g15236(csa_tree_add_6_33_groupi_n_3193 ,csa_tree_add_6_33_groupi_n_1799 ,csa_tree_add_6_33_groupi_n_2804);
  and csa_tree_add_6_33_groupi_g15237(csa_tree_add_6_33_groupi_n_3192 ,csa_tree_add_6_33_groupi_n_2371 ,csa_tree_add_6_33_groupi_n_2854);
  and csa_tree_add_6_33_groupi_g15238(csa_tree_add_6_33_groupi_n_3191 ,csa_tree_add_6_33_groupi_n_1789 ,csa_tree_add_6_33_groupi_n_2864);
  and csa_tree_add_6_33_groupi_g15239(csa_tree_add_6_33_groupi_n_3190 ,csa_tree_add_6_33_groupi_n_1685 ,csa_tree_add_6_33_groupi_n_2871);
  and csa_tree_add_6_33_groupi_g15240(csa_tree_add_6_33_groupi_n_3189 ,csa_tree_add_6_33_groupi_n_1739 ,csa_tree_add_6_33_groupi_n_2788);
  and csa_tree_add_6_33_groupi_g15241(csa_tree_add_6_33_groupi_n_3188 ,csa_tree_add_6_33_groupi_n_1848 ,csa_tree_add_6_33_groupi_n_2812);
  and csa_tree_add_6_33_groupi_g15242(csa_tree_add_6_33_groupi_n_3187 ,csa_tree_add_6_33_groupi_n_1912 ,csa_tree_add_6_33_groupi_n_2869);
  and csa_tree_add_6_33_groupi_g15243(csa_tree_add_6_33_groupi_n_3186 ,csa_tree_add_6_33_groupi_n_2486 ,csa_tree_add_6_33_groupi_n_2817);
  or csa_tree_add_6_33_groupi_g15244(csa_tree_add_6_33_groupi_n_3185 ,csa_tree_add_6_33_groupi_n_1753 ,csa_tree_add_6_33_groupi_n_2832);
  not csa_tree_add_6_33_groupi_g15245(csa_tree_add_6_33_groupi_n_3053 ,csa_tree_add_6_33_groupi_n_3054);
  not csa_tree_add_6_33_groupi_g15246(csa_tree_add_6_33_groupi_n_3051 ,csa_tree_add_6_33_groupi_n_3052);
  not csa_tree_add_6_33_groupi_g15247(csa_tree_add_6_33_groupi_n_3046 ,csa_tree_add_6_33_groupi_n_3045);
  not csa_tree_add_6_33_groupi_g15248(csa_tree_add_6_33_groupi_n_3041 ,csa_tree_add_6_33_groupi_n_3042);
  not csa_tree_add_6_33_groupi_g15249(csa_tree_add_6_33_groupi_n_3039 ,csa_tree_add_6_33_groupi_n_3040);
  not csa_tree_add_6_33_groupi_g15250(csa_tree_add_6_33_groupi_n_3037 ,csa_tree_add_6_33_groupi_n_3038);
  not csa_tree_add_6_33_groupi_g15251(csa_tree_add_6_33_groupi_n_3035 ,csa_tree_add_6_33_groupi_n_3036);
  and csa_tree_add_6_33_groupi_g15252(csa_tree_add_6_33_groupi_n_3034 ,csa_tree_add_6_33_groupi_n_2630 ,csa_tree_add_6_33_groupi_n_2629);
  or csa_tree_add_6_33_groupi_g15253(csa_tree_add_6_33_groupi_n_3033 ,csa_tree_add_6_33_groupi_n_2446 ,csa_tree_add_6_33_groupi_n_2664);
  and csa_tree_add_6_33_groupi_g15254(csa_tree_add_6_33_groupi_n_3032 ,csa_tree_add_6_33_groupi_n_2660 ,csa_tree_add_6_33_groupi_n_2626);
  or csa_tree_add_6_33_groupi_g15255(csa_tree_add_6_33_groupi_n_3031 ,csa_tree_add_6_33_groupi_n_2564 ,csa_tree_add_6_33_groupi_n_2784);
  or csa_tree_add_6_33_groupi_g15256(csa_tree_add_6_33_groupi_n_3030 ,csa_tree_add_6_33_groupi_n_2450 ,csa_tree_add_6_33_groupi_n_2623);
  and csa_tree_add_6_33_groupi_g15257(csa_tree_add_6_33_groupi_n_3029 ,csa_tree_add_6_33_groupi_n_2450 ,csa_tree_add_6_33_groupi_n_2623);
  or csa_tree_add_6_33_groupi_g15258(csa_tree_add_6_33_groupi_n_3028 ,csa_tree_add_6_33_groupi_n_1396 ,csa_tree_add_6_33_groupi_n_2717);
  nor csa_tree_add_6_33_groupi_g15259(csa_tree_add_6_33_groupi_n_3027 ,csa_tree_add_6_33_groupi_n_2445 ,csa_tree_add_6_33_groupi_n_2665);
  or csa_tree_add_6_33_groupi_g15260(csa_tree_add_6_33_groupi_n_3026 ,csa_tree_add_6_33_groupi_n_2730 ,csa_tree_add_6_33_groupi_n_2779);
  or csa_tree_add_6_33_groupi_g15261(csa_tree_add_6_33_groupi_n_3025 ,csa_tree_add_6_33_groupi_n_2908 ,csa_tree_add_6_33_groupi_n_2625);
  nor csa_tree_add_6_33_groupi_g15262(csa_tree_add_6_33_groupi_n_3024 ,csa_tree_add_6_33_groupi_n_2909 ,csa_tree_add_6_33_groupi_n_2624);
  or csa_tree_add_6_33_groupi_g15263(csa_tree_add_6_33_groupi_n_3023 ,csa_tree_add_6_33_groupi_n_2559 ,csa_tree_add_6_33_groupi_n_2777);
  or csa_tree_add_6_33_groupi_g15264(csa_tree_add_6_33_groupi_n_3022 ,csa_tree_add_6_33_groupi_n_2637 ,csa_tree_add_6_33_groupi_n_2619);
  or csa_tree_add_6_33_groupi_g15265(csa_tree_add_6_33_groupi_n_3021 ,csa_tree_add_6_33_groupi_n_2463 ,csa_tree_add_6_33_groupi_n_2775);
  or csa_tree_add_6_33_groupi_g15266(csa_tree_add_6_33_groupi_n_3020 ,csa_tree_add_6_33_groupi_n_2464 ,csa_tree_add_6_33_groupi_n_2772);
  or csa_tree_add_6_33_groupi_g15267(csa_tree_add_6_33_groupi_n_3019 ,csa_tree_add_6_33_groupi_n_2617 ,csa_tree_add_6_33_groupi_n_2616);
  nor csa_tree_add_6_33_groupi_g15268(csa_tree_add_6_33_groupi_n_3018 ,csa_tree_add_6_33_groupi_n_2638 ,csa_tree_add_6_33_groupi_n_2618);
  and csa_tree_add_6_33_groupi_g15269(csa_tree_add_6_33_groupi_n_3017 ,csa_tree_add_6_33_groupi_n_2617 ,csa_tree_add_6_33_groupi_n_2616);
  or csa_tree_add_6_33_groupi_g15270(csa_tree_add_6_33_groupi_n_3016 ,csa_tree_add_6_33_groupi_n_2727 ,csa_tree_add_6_33_groupi_n_2773);
  or csa_tree_add_6_33_groupi_g15271(csa_tree_add_6_33_groupi_n_3015 ,csa_tree_add_6_33_groupi_n_2612 ,csa_tree_add_6_33_groupi_n_2610);
  or csa_tree_add_6_33_groupi_g15272(csa_tree_add_6_33_groupi_n_3014 ,csa_tree_add_6_33_groupi_n_2460 ,csa_tree_add_6_33_groupi_n_2769);
  and csa_tree_add_6_33_groupi_g15273(csa_tree_add_6_33_groupi_n_3013 ,csa_tree_add_6_33_groupi_n_2612 ,csa_tree_add_6_33_groupi_n_2610);
  or csa_tree_add_6_33_groupi_g15274(csa_tree_add_6_33_groupi_n_3012 ,csa_tree_add_6_33_groupi_n_2606 ,csa_tree_add_6_33_groupi_n_2603);
  or csa_tree_add_6_33_groupi_g15275(csa_tree_add_6_33_groupi_n_3011 ,csa_tree_add_6_33_groupi_n_2607 ,csa_tree_add_6_33_groupi_n_2605);
  and csa_tree_add_6_33_groupi_g15276(csa_tree_add_6_33_groupi_n_3010 ,csa_tree_add_6_33_groupi_n_2607 ,csa_tree_add_6_33_groupi_n_2605);
  or csa_tree_add_6_33_groupi_g15277(csa_tree_add_6_33_groupi_n_3009 ,csa_tree_add_6_33_groupi_n_2526 ,csa_tree_add_6_33_groupi_n_2604);
  and csa_tree_add_6_33_groupi_g15278(csa_tree_add_6_33_groupi_n_3008 ,csa_tree_add_6_33_groupi_n_2678 ,csa_tree_add_6_33_groupi_n_2713);
  or csa_tree_add_6_33_groupi_g15279(csa_tree_add_6_33_groupi_n_3007 ,csa_tree_add_6_33_groupi_n_2437 ,csa_tree_add_6_33_groupi_n_2600);
  or csa_tree_add_6_33_groupi_g15280(csa_tree_add_6_33_groupi_n_3006 ,csa_tree_add_6_33_groupi_n_2474 ,csa_tree_add_6_33_groupi_n_2767);
  or csa_tree_add_6_33_groupi_g15281(csa_tree_add_6_33_groupi_n_3005 ,csa_tree_add_6_33_groupi_n_2478 ,csa_tree_add_6_33_groupi_n_2765);
  and csa_tree_add_6_33_groupi_g15282(csa_tree_add_6_33_groupi_n_3004 ,csa_tree_add_6_33_groupi_n_2526 ,csa_tree_add_6_33_groupi_n_2604);
  or csa_tree_add_6_33_groupi_g15283(csa_tree_add_6_33_groupi_n_3003 ,csa_tree_add_6_33_groupi_n_2573 ,csa_tree_add_6_33_groupi_n_2762);
  or csa_tree_add_6_33_groupi_g15284(csa_tree_add_6_33_groupi_n_3002 ,csa_tree_add_6_33_groupi_n_2599 ,csa_tree_add_6_33_groupi_n_2598);
  or csa_tree_add_6_33_groupi_g15285(csa_tree_add_6_33_groupi_n_3001 ,csa_tree_add_6_33_groupi_n_2335 ,csa_tree_add_6_33_groupi_n_2597);
  and csa_tree_add_6_33_groupi_g15286(csa_tree_add_6_33_groupi_n_3000 ,csa_tree_add_6_33_groupi_n_2335 ,csa_tree_add_6_33_groupi_n_2597);
  and csa_tree_add_6_33_groupi_g15287(csa_tree_add_6_33_groupi_n_2999 ,csa_tree_add_6_33_groupi_n_2606 ,csa_tree_add_6_33_groupi_n_2603);
  or csa_tree_add_6_33_groupi_g15288(csa_tree_add_6_33_groupi_n_2998 ,csa_tree_add_6_33_groupi_n_2479 ,csa_tree_add_6_33_groupi_n_2758);
  and csa_tree_add_6_33_groupi_g15289(csa_tree_add_6_33_groupi_n_2997 ,csa_tree_add_6_33_groupi_n_2599 ,csa_tree_add_6_33_groupi_n_2598);
  or csa_tree_add_6_33_groupi_g15290(csa_tree_add_6_33_groupi_n_2996 ,csa_tree_add_6_33_groupi_n_2595 ,csa_tree_add_6_33_groupi_n_2627);
  and csa_tree_add_6_33_groupi_g15291(csa_tree_add_6_33_groupi_n_2995 ,csa_tree_add_6_33_groupi_n_2901 ,csa_tree_add_6_33_groupi_n_2686);
  and csa_tree_add_6_33_groupi_g15292(csa_tree_add_6_33_groupi_n_2994 ,csa_tree_add_6_33_groupi_n_2437 ,csa_tree_add_6_33_groupi_n_2600);
  or csa_tree_add_6_33_groupi_g15293(csa_tree_add_6_33_groupi_n_2993 ,csa_tree_add_6_33_groupi_n_2427 ,csa_tree_add_6_33_groupi_n_2593);
  or csa_tree_add_6_33_groupi_g15294(csa_tree_add_6_33_groupi_n_2992 ,csa_tree_add_6_33_groupi_n_2594 ,csa_tree_add_6_33_groupi_n_2700);
  and csa_tree_add_6_33_groupi_g15295(csa_tree_add_6_33_groupi_n_2991 ,csa_tree_add_6_33_groupi_n_2427 ,csa_tree_add_6_33_groupi_n_2593);
  or csa_tree_add_6_33_groupi_g15296(csa_tree_add_6_33_groupi_n_2990 ,csa_tree_add_6_33_groupi_n_2592 ,csa_tree_add_6_33_groupi_n_2591);
  or csa_tree_add_6_33_groupi_g15297(csa_tree_add_6_33_groupi_n_2989 ,csa_tree_add_6_33_groupi_n_2483 ,csa_tree_add_6_33_groupi_n_2865);
  or csa_tree_add_6_33_groupi_g15298(csa_tree_add_6_33_groupi_n_2988 ,csa_tree_add_6_33_groupi_n_2569 ,csa_tree_add_6_33_groupi_n_2857);
  and csa_tree_add_6_33_groupi_g15299(csa_tree_add_6_33_groupi_n_2987 ,csa_tree_add_6_33_groupi_n_2592 ,csa_tree_add_6_33_groupi_n_2591);
  or csa_tree_add_6_33_groupi_g15300(csa_tree_add_6_33_groupi_n_2986 ,csa_tree_add_6_33_groupi_n_2327 ,csa_tree_add_6_33_groupi_n_2688);
  or csa_tree_add_6_33_groupi_g15301(csa_tree_add_6_33_groupi_n_2985 ,csa_tree_add_6_33_groupi_n_2912 ,csa_tree_add_6_33_groupi_n_2827);
  and csa_tree_add_6_33_groupi_g15302(csa_tree_add_6_33_groupi_n_2984 ,csa_tree_add_6_33_groupi_n_2365 ,csa_tree_add_6_33_groupi_n_2863);
  or csa_tree_add_6_33_groupi_g15303(csa_tree_add_6_33_groupi_n_2983 ,csa_tree_add_6_33_groupi_n_2910 ,csa_tree_add_6_33_groupi_n_2690);
  nor csa_tree_add_6_33_groupi_g15304(csa_tree_add_6_33_groupi_n_2982 ,csa_tree_add_6_33_groupi_n_2911 ,csa_tree_add_6_33_groupi_n_2691);
  or csa_tree_add_6_33_groupi_g15305(csa_tree_add_6_33_groupi_n_2981 ,csa_tree_add_6_33_groupi_n_2356 ,csa_tree_add_6_33_groupi_n_2843);
  nor csa_tree_add_6_33_groupi_g15306(csa_tree_add_6_33_groupi_n_2980 ,csa_tree_add_6_33_groupi_n_2366 ,csa_tree_add_6_33_groupi_n_2792);
  or csa_tree_add_6_33_groupi_g15307(csa_tree_add_6_33_groupi_n_2979 ,csa_tree_add_6_33_groupi_n_2660 ,csa_tree_add_6_33_groupi_n_2626);
  xnor csa_tree_add_6_33_groupi_g15308(csa_tree_add_6_33_groupi_n_2978 ,csa_tree_add_6_33_groupi_n_2546 ,csa_tree_add_6_33_groupi_n_2427);
  xnor csa_tree_add_6_33_groupi_g15309(csa_tree_add_6_33_groupi_n_2977 ,csa_tree_add_6_33_groupi_n_2379 ,csa_tree_add_6_33_groupi_n_2423);
  xnor csa_tree_add_6_33_groupi_g15310(csa_tree_add_6_33_groupi_n_2976 ,csa_tree_add_6_33_groupi_n_2535 ,csa_tree_add_6_33_groupi_n_2413);
  xnor csa_tree_add_6_33_groupi_g15311(csa_tree_add_6_33_groupi_n_2975 ,csa_tree_add_6_33_groupi_n_2573 ,csa_tree_add_6_33_groupi_n_2431);
  xnor csa_tree_add_6_33_groupi_g15312(csa_tree_add_6_33_groupi_n_2974 ,csa_tree_add_6_33_groupi_n_2454 ,csa_tree_add_6_33_groupi_n_2559);
  xnor csa_tree_add_6_33_groupi_g15313(csa_tree_add_6_33_groupi_n_2973 ,csa_tree_add_6_33_groupi_n_2342 ,csa_tree_add_6_33_groupi_n_2383);
  xnor csa_tree_add_6_33_groupi_g15314(csa_tree_add_6_33_groupi_n_2972 ,csa_tree_add_6_33_groupi_n_1138 ,csa_tree_add_6_33_groupi_n_2406);
  xnor csa_tree_add_6_33_groupi_g15315(csa_tree_add_6_33_groupi_n_2971 ,csa_tree_add_6_33_groupi_n_1134 ,csa_tree_add_6_33_groupi_n_2398);
  xnor csa_tree_add_6_33_groupi_g15316(csa_tree_add_6_33_groupi_n_2970 ,csa_tree_add_6_33_groupi_n_2380 ,csa_tree_add_6_33_groupi_n_2496);
  xnor csa_tree_add_6_33_groupi_g15317(csa_tree_add_6_33_groupi_n_2969 ,csa_tree_add_6_33_groupi_n_2579 ,csa_tree_add_6_33_groupi_n_2418);
  xnor csa_tree_add_6_33_groupi_g15318(csa_tree_add_6_33_groupi_n_2968 ,csa_tree_add_6_33_groupi_n_2330 ,csa_tree_add_6_33_groupi_n_2387);
  xnor csa_tree_add_6_33_groupi_g15319(csa_tree_add_6_33_groupi_n_2967 ,csa_tree_add_6_33_groupi_n_2564 ,csa_tree_add_6_33_groupi_n_2533);
  xnor csa_tree_add_6_33_groupi_g15320(csa_tree_add_6_33_groupi_n_2966 ,csa_tree_add_6_33_groupi_n_2456 ,csa_tree_add_6_33_groupi_n_2446);
  xnor csa_tree_add_6_33_groupi_g15321(csa_tree_add_6_33_groupi_n_2965 ,csa_tree_add_6_33_groupi_n_2333 ,csa_tree_add_6_33_groupi_n_2434);
  xnor csa_tree_add_6_33_groupi_g15322(csa_tree_add_6_33_groupi_n_2964 ,csa_tree_add_6_33_groupi_n_2542 ,csa_tree_add_6_33_groupi_n_2420);
  xnor csa_tree_add_6_33_groupi_g15323(csa_tree_add_6_33_groupi_n_2963 ,csa_tree_add_6_33_groupi_n_1376 ,csa_tree_add_6_33_groupi_n_2415);
  xnor csa_tree_add_6_33_groupi_g15324(csa_tree_add_6_33_groupi_n_2962 ,csa_tree_add_6_33_groupi_n_2443 ,csa_tree_add_6_33_groupi_n_2401);
  xnor csa_tree_add_6_33_groupi_g15325(csa_tree_add_6_33_groupi_n_2961 ,csa_tree_add_6_33_groupi_n_2524 ,csa_tree_add_6_33_groupi_n_2528);
  xnor csa_tree_add_6_33_groupi_g15326(csa_tree_add_6_33_groupi_n_2960 ,csa_tree_add_6_33_groupi_n_1414 ,csa_tree_add_6_33_groupi_n_2411);
  xnor csa_tree_add_6_33_groupi_g15327(csa_tree_add_6_33_groupi_n_2959 ,csa_tree_add_6_33_groupi_n_2344 ,csa_tree_add_6_33_groupi_n_2478);
  xnor csa_tree_add_6_33_groupi_g15328(csa_tree_add_6_33_groupi_n_2958 ,csa_tree_add_6_33_groupi_n_2346 ,csa_tree_add_6_33_groupi_n_2560);
  xnor csa_tree_add_6_33_groupi_g15329(csa_tree_add_6_33_groupi_n_2957 ,csa_tree_add_6_33_groupi_n_2561 ,csa_tree_add_6_33_groupi_n_2327);
  xnor csa_tree_add_6_33_groupi_g15330(csa_tree_add_6_33_groupi_n_2956 ,csa_tree_add_6_33_groupi_n_2337 ,csa_tree_add_6_33_groupi_n_2408);
  xnor csa_tree_add_6_33_groupi_g15331(csa_tree_add_6_33_groupi_n_2955 ,csa_tree_add_6_33_groupi_n_2338 ,csa_tree_add_6_33_groupi_n_2565);
  xnor csa_tree_add_6_33_groupi_g15332(csa_tree_add_6_33_groupi_n_2954 ,csa_tree_add_6_33_groupi_n_2339 ,csa_tree_add_6_33_groupi_n_2416);
  xnor csa_tree_add_6_33_groupi_g15333(csa_tree_add_6_33_groupi_n_2953 ,csa_tree_add_6_33_groupi_n_2495 ,csa_tree_add_6_33_groupi_n_2334);
  xnor csa_tree_add_6_33_groupi_g15334(csa_tree_add_6_33_groupi_n_2952 ,csa_tree_add_6_33_groupi_n_2447 ,csa_tree_add_6_33_groupi_n_2336);
  xnor csa_tree_add_6_33_groupi_g15335(csa_tree_add_6_33_groupi_n_2951 ,csa_tree_add_6_33_groupi_n_1145 ,csa_tree_add_6_33_groupi_n_2479);
  xnor csa_tree_add_6_33_groupi_g15336(csa_tree_add_6_33_groupi_n_2950 ,csa_tree_add_6_33_groupi_n_2526 ,csa_tree_add_6_33_groupi_n_2475);
  xnor csa_tree_add_6_33_groupi_g15337(csa_tree_add_6_33_groupi_n_2949 ,csa_tree_add_6_33_groupi_n_1150 ,csa_tree_add_6_33_groupi_n_2464);
  xnor csa_tree_add_6_33_groupi_g15338(csa_tree_add_6_33_groupi_n_2948 ,csa_tree_add_6_33_groupi_n_2391 ,csa_tree_add_6_33_groupi_n_2499);
  xnor csa_tree_add_6_33_groupi_g15339(csa_tree_add_6_33_groupi_n_2947 ,csa_tree_add_6_33_groupi_n_2396 ,csa_tree_add_6_33_groupi_n_2510);
  xnor csa_tree_add_6_33_groupi_g15340(csa_tree_add_6_33_groupi_n_2946 ,csa_tree_add_6_33_groupi_n_1157 ,csa_tree_add_6_33_groupi_n_2575);
  xnor csa_tree_add_6_33_groupi_g15341(csa_tree_add_6_33_groupi_n_2945 ,csa_tree_add_6_33_groupi_n_2438 ,csa_tree_add_6_33_groupi_n_2439);
  xnor csa_tree_add_6_33_groupi_g15342(csa_tree_add_6_33_groupi_n_2944 ,csa_tree_add_6_33_groupi_n_2500 ,csa_tree_add_6_33_groupi_n_2580);
  xnor csa_tree_add_6_33_groupi_g15343(csa_tree_add_6_33_groupi_n_2943 ,csa_tree_add_6_33_groupi_n_2512 ,csa_tree_add_6_33_groupi_n_2540);
  xor csa_tree_add_6_33_groupi_g15344(csa_tree_add_6_33_groupi_n_2942 ,csa_tree_add_6_33_groupi_n_1397 ,csa_tree_add_6_33_groupi_n_2562);
  xnor csa_tree_add_6_33_groupi_g15345(csa_tree_add_6_33_groupi_n_2941 ,csa_tree_add_6_33_groupi_n_2517 ,csa_tree_add_6_33_groupi_n_2509);
  xnor csa_tree_add_6_33_groupi_g15346(csa_tree_add_6_33_groupi_n_2940 ,csa_tree_add_6_33_groupi_n_2494 ,csa_tree_add_6_33_groupi_n_2558);
  xnor csa_tree_add_6_33_groupi_g15347(csa_tree_add_6_33_groupi_n_2939 ,csa_tree_add_6_33_groupi_n_2381 ,csa_tree_add_6_33_groupi_n_2566);
  xnor csa_tree_add_6_33_groupi_g15348(csa_tree_add_6_33_groupi_n_2938 ,csa_tree_add_6_33_groupi_n_1417 ,csa_tree_add_6_33_groupi_n_2554);
  xnor csa_tree_add_6_33_groupi_g15349(csa_tree_add_6_33_groupi_n_2937 ,csa_tree_add_6_33_groupi_n_2541 ,csa_tree_add_6_33_groupi_n_2531);
  xnor csa_tree_add_6_33_groupi_g15350(csa_tree_add_6_33_groupi_n_2936 ,csa_tree_add_6_33_groupi_n_2567 ,csa_tree_add_6_33_groupi_n_2532);
  xnor csa_tree_add_6_33_groupi_g15351(csa_tree_add_6_33_groupi_n_2935 ,csa_tree_add_6_33_groupi_n_2444 ,csa_tree_add_6_33_groupi_n_2462);
  xnor csa_tree_add_6_33_groupi_g15352(csa_tree_add_6_33_groupi_n_2934 ,csa_tree_add_6_33_groupi_n_2523 ,csa_tree_add_6_33_groupi_n_2471);
  xnor csa_tree_add_6_33_groupi_g15353(csa_tree_add_6_33_groupi_n_2933 ,csa_tree_add_6_33_groupi_n_1370 ,csa_tree_add_6_33_groupi_n_2435);
  xnor csa_tree_add_6_33_groupi_g15354(csa_tree_add_6_33_groupi_n_2932 ,csa_tree_add_6_33_groupi_n_2470 ,csa_tree_add_6_33_groupi_n_2506);
  xnor csa_tree_add_6_33_groupi_g15355(csa_tree_add_6_33_groupi_n_2931 ,csa_tree_add_6_33_groupi_n_2385 ,csa_tree_add_6_33_groupi_n_2428);
  xnor csa_tree_add_6_33_groupi_g15356(csa_tree_add_6_33_groupi_n_2930 ,csa_tree_add_6_33_groupi_n_2511 ,csa_tree_add_6_33_groupi_n_2516);
  xnor csa_tree_add_6_33_groupi_g15357(csa_tree_add_6_33_groupi_n_2929 ,csa_tree_add_6_33_groupi_n_2552 ,csa_tree_add_6_33_groupi_n_2518);
  xnor csa_tree_add_6_33_groupi_g15358(csa_tree_add_6_33_groupi_n_2928 ,csa_tree_add_6_33_groupi_n_1072 ,csa_tree_add_6_33_groupi_n_2574);
  xnor csa_tree_add_6_33_groupi_g15359(csa_tree_add_6_33_groupi_n_2927 ,csa_tree_add_6_33_groupi_n_1206 ,csa_tree_add_6_33_groupi_n_2553);
  xnor csa_tree_add_6_33_groupi_g15360(csa_tree_add_6_33_groupi_n_2926 ,csa_tree_add_6_33_groupi_n_2407 ,csa_tree_add_6_33_groupi_n_2404);
  xnor csa_tree_add_6_33_groupi_g15361(csa_tree_add_6_33_groupi_n_2925 ,csa_tree_add_6_33_groupi_n_2449 ,csa_tree_add_6_33_groupi_n_2525);
  xnor csa_tree_add_6_33_groupi_g15362(csa_tree_add_6_33_groupi_n_2924 ,csa_tree_add_6_33_groupi_n_1481 ,csa_tree_add_6_33_groupi_n_2465);
  xnor csa_tree_add_6_33_groupi_g15363(csa_tree_add_6_33_groupi_n_2923 ,csa_tree_add_6_33_groupi_n_2403 ,csa_tree_add_6_33_groupi_n_2399);
  xnor csa_tree_add_6_33_groupi_g15364(csa_tree_add_6_33_groupi_n_2922 ,csa_tree_add_6_33_groupi_n_1404 ,csa_tree_add_6_33_groupi_n_2551);
  xnor csa_tree_add_6_33_groupi_g15365(csa_tree_add_6_33_groupi_n_2921 ,csa_tree_add_6_33_groupi_n_2458 ,csa_tree_add_6_33_groupi_n_2507);
  xnor csa_tree_add_6_33_groupi_g15366(csa_tree_add_6_33_groupi_n_2920 ,csa_tree_add_6_33_groupi_n_2483 ,csa_tree_add_6_33_groupi_n_2424);
  xnor csa_tree_add_6_33_groupi_g15367(csa_tree_add_6_33_groupi_n_2919 ,csa_tree_add_6_33_groupi_n_2384 ,csa_tree_add_6_33_groupi_n_2477);
  xnor csa_tree_add_6_33_groupi_g15368(csa_tree_add_6_33_groupi_n_2918 ,csa_tree_add_6_33_groupi_n_2436 ,csa_tree_add_6_33_groupi_n_2432);
  xnor csa_tree_add_6_33_groupi_g15369(csa_tree_add_6_33_groupi_n_2917 ,csa_tree_add_6_33_groupi_n_2484 ,csa_tree_add_6_33_groupi_n_2376);
  xnor csa_tree_add_6_33_groupi_g15370(csa_tree_add_6_33_groupi_n_2916 ,csa_tree_add_6_33_groupi_n_2522 ,csa_tree_add_6_33_groupi_n_2501);
  xnor csa_tree_add_6_33_groupi_g15371(csa_tree_add_6_33_groupi_n_3059 ,csa_tree_add_6_33_groupi_n_2577 ,csa_tree_add_6_33_groupi_n_2139);
  xnor csa_tree_add_6_33_groupi_g15372(csa_tree_add_6_33_groupi_n_3058 ,csa_tree_add_6_33_groupi_n_2461 ,csa_tree_add_6_33_groupi_n_2037);
  xnor csa_tree_add_6_33_groupi_g15373(csa_tree_add_6_33_groupi_n_3057 ,csa_tree_add_6_33_groupi_n_2563 ,csa_tree_add_6_33_groupi_n_2060);
  xnor csa_tree_add_6_33_groupi_g15374(csa_tree_add_6_33_groupi_n_3056 ,csa_tree_add_6_33_groupi_n_2457 ,csa_tree_add_6_33_groupi_n_2179);
  xnor csa_tree_add_6_33_groupi_g15375(csa_tree_add_6_33_groupi_n_3055 ,csa_tree_add_6_33_groupi_n_2459 ,csa_tree_add_6_33_groupi_n_2035);
  xnor csa_tree_add_6_33_groupi_g15376(csa_tree_add_6_33_groupi_n_3054 ,csa_tree_add_6_33_groupi_n_2468 ,csa_tree_add_6_33_groupi_n_2030);
  xnor csa_tree_add_6_33_groupi_g15377(csa_tree_add_6_33_groupi_n_3052 ,csa_tree_add_6_33_groupi_n_2466 ,csa_tree_add_6_33_groupi_n_2063);
  xnor csa_tree_add_6_33_groupi_g15378(csa_tree_add_6_33_groupi_n_3050 ,csa_tree_add_6_33_groupi_n_2537 ,csa_tree_add_6_33_groupi_n_2038);
  xnor csa_tree_add_6_33_groupi_g15379(csa_tree_add_6_33_groupi_n_3049 ,csa_tree_add_6_33_groupi_n_2538 ,csa_tree_add_6_33_groupi_n_2070);
  xnor csa_tree_add_6_33_groupi_g15380(csa_tree_add_6_33_groupi_n_3048 ,csa_tree_add_6_33_groupi_n_2578 ,csa_tree_add_6_33_groupi_n_2059);
  xnor csa_tree_add_6_33_groupi_g15381(csa_tree_add_6_33_groupi_n_3047 ,csa_tree_add_6_33_groupi_n_2576 ,csa_tree_add_6_33_groupi_n_2043);
  and csa_tree_add_6_33_groupi_g15382(csa_tree_add_6_33_groupi_n_3045 ,csa_tree_add_6_33_groupi_n_1920 ,csa_tree_add_6_33_groupi_n_2764);
  and csa_tree_add_6_33_groupi_g15383(csa_tree_add_6_33_groupi_n_3044 ,csa_tree_add_6_33_groupi_n_1850 ,csa_tree_add_6_33_groupi_n_2831);
  xnor csa_tree_add_6_33_groupi_g15384(csa_tree_add_6_33_groupi_n_3043 ,csa_tree_add_6_33_groupi_n_2571 ,csa_tree_add_6_33_groupi_n_2110);
  and csa_tree_add_6_33_groupi_g15385(csa_tree_add_6_33_groupi_n_3042 ,csa_tree_add_6_33_groupi_n_2372 ,csa_tree_add_6_33_groupi_n_2771);
  xnor csa_tree_add_6_33_groupi_g15386(csa_tree_add_6_33_groupi_n_3040 ,csa_tree_add_6_33_groupi_n_2473 ,csa_tree_add_6_33_groupi_n_2162);
  and csa_tree_add_6_33_groupi_g15387(csa_tree_add_6_33_groupi_n_3038 ,csa_tree_add_6_33_groupi_n_1759 ,csa_tree_add_6_33_groupi_n_2828);
  and csa_tree_add_6_33_groupi_g15388(csa_tree_add_6_33_groupi_n_3036 ,csa_tree_add_6_33_groupi_n_1717 ,csa_tree_add_6_33_groupi_n_2783);
  not csa_tree_add_6_33_groupi_g15389(csa_tree_add_6_33_groupi_n_2914 ,csa_tree_add_6_33_groupi_n_2913);
  not csa_tree_add_6_33_groupi_g15390(csa_tree_add_6_33_groupi_n_2911 ,csa_tree_add_6_33_groupi_n_2910);
  not csa_tree_add_6_33_groupi_g15391(csa_tree_add_6_33_groupi_n_2909 ,csa_tree_add_6_33_groupi_n_2908);
  not csa_tree_add_6_33_groupi_g15392(csa_tree_add_6_33_groupi_n_2906 ,csa_tree_add_6_33_groupi_n_2907);
  not csa_tree_add_6_33_groupi_g15393(csa_tree_add_6_33_groupi_n_2904 ,csa_tree_add_6_33_groupi_n_2905);
  not csa_tree_add_6_33_groupi_g15394(csa_tree_add_6_33_groupi_n_2903 ,csa_tree_add_6_33_groupi_n_2902);
  not csa_tree_add_6_33_groupi_g15395(csa_tree_add_6_33_groupi_n_2901 ,csa_tree_add_6_33_groupi_n_2900);
  not csa_tree_add_6_33_groupi_g15396(csa_tree_add_6_33_groupi_n_2898 ,csa_tree_add_6_33_groupi_n_2899);
  not csa_tree_add_6_33_groupi_g15397(csa_tree_add_6_33_groupi_n_2895 ,csa_tree_add_6_33_groupi_n_2896);
  not csa_tree_add_6_33_groupi_g15398(csa_tree_add_6_33_groupi_n_2893 ,csa_tree_add_6_33_groupi_n_2894);
  not csa_tree_add_6_33_groupi_g15399(csa_tree_add_6_33_groupi_n_2891 ,csa_tree_add_6_33_groupi_n_2892);
  not csa_tree_add_6_33_groupi_g15400(csa_tree_add_6_33_groupi_n_2890 ,csa_tree_add_6_33_groupi_n_2889);
  or csa_tree_add_6_33_groupi_g15401(csa_tree_add_6_33_groupi_n_2887 ,csa_tree_add_6_33_groupi_n_1681 ,csa_tree_add_6_33_groupi_n_2467);
  nor csa_tree_add_6_33_groupi_g15402(csa_tree_add_6_33_groupi_n_2886 ,csa_tree_add_6_33_groupi_n_2338 ,csa_tree_add_6_33_groupi_n_2419);
  or csa_tree_add_6_33_groupi_g15403(csa_tree_add_6_33_groupi_n_2885 ,csa_tree_add_6_33_groupi_n_2525 ,csa_tree_add_6_33_groupi_n_2449);
  or csa_tree_add_6_33_groupi_g15404(csa_tree_add_6_33_groupi_n_2884 ,csa_tree_add_6_33_groupi_n_2510 ,csa_tree_add_6_33_groupi_n_2396);
  and csa_tree_add_6_33_groupi_g15405(csa_tree_add_6_33_groupi_n_2883 ,csa_tree_add_6_33_groupi_n_2510 ,csa_tree_add_6_33_groupi_n_2396);
  and csa_tree_add_6_33_groupi_g15406(csa_tree_add_6_33_groupi_n_2882 ,csa_tree_add_6_33_groupi_n_2331 ,csa_tree_add_6_33_groupi_n_2387);
  or csa_tree_add_6_33_groupi_g15407(csa_tree_add_6_33_groupi_n_2881 ,csa_tree_add_6_33_groupi_n_1157 ,csa_tree_add_6_33_groupi_n_2422);
  and csa_tree_add_6_33_groupi_g15408(csa_tree_add_6_33_groupi_n_2880 ,csa_tree_add_6_33_groupi_n_2340 ,csa_tree_add_6_33_groupi_n_2421);
  or csa_tree_add_6_33_groupi_g15409(csa_tree_add_6_33_groupi_n_2879 ,csa_tree_add_6_33_groupi_n_1072 ,csa_tree_add_6_33_groupi_n_2508);
  or csa_tree_add_6_33_groupi_g15410(csa_tree_add_6_33_groupi_n_2878 ,csa_tree_add_6_33_groupi_n_2528 ,csa_tree_add_6_33_groupi_n_2524);
  and csa_tree_add_6_33_groupi_g15411(csa_tree_add_6_33_groupi_n_2877 ,csa_tree_add_6_33_groupi_n_1417 ,csa_tree_add_6_33_groupi_n_2527);
  or csa_tree_add_6_33_groupi_g15412(csa_tree_add_6_33_groupi_n_2876 ,csa_tree_add_6_33_groupi_n_2509 ,csa_tree_add_6_33_groupi_n_2517);
  and csa_tree_add_6_33_groupi_g15413(csa_tree_add_6_33_groupi_n_2875 ,csa_tree_add_6_33_groupi_n_2509 ,csa_tree_add_6_33_groupi_n_2517);
  or csa_tree_add_6_33_groupi_g15414(csa_tree_add_6_33_groupi_n_2874 ,csa_tree_add_6_33_groupi_n_1408 ,csa_tree_add_6_33_groupi_n_2392);
  or csa_tree_add_6_33_groupi_g15415(csa_tree_add_6_33_groupi_n_2873 ,csa_tree_add_6_33_groupi_n_2347 ,csa_tree_add_6_33_groupi_n_2417);
  nor csa_tree_add_6_33_groupi_g15416(csa_tree_add_6_33_groupi_n_2872 ,csa_tree_add_6_33_groupi_n_2348 ,csa_tree_add_6_33_groupi_n_2418);
  or csa_tree_add_6_33_groupi_g15417(csa_tree_add_6_33_groupi_n_2871 ,csa_tree_add_6_33_groupi_n_1654 ,csa_tree_add_6_33_groupi_n_2577);
  nor csa_tree_add_6_33_groupi_g15418(csa_tree_add_6_33_groupi_n_2870 ,csa_tree_add_6_33_groupi_n_2340 ,csa_tree_add_6_33_groupi_n_2421);
  or csa_tree_add_6_33_groupi_g15419(csa_tree_add_6_33_groupi_n_2869 ,csa_tree_add_6_33_groupi_n_1803 ,csa_tree_add_6_33_groupi_n_2576);
  nor csa_tree_add_6_33_groupi_g15420(csa_tree_add_6_33_groupi_n_2868 ,csa_tree_add_6_33_groupi_n_2342 ,csa_tree_add_6_33_groupi_n_2382);
  or csa_tree_add_6_33_groupi_g15421(csa_tree_add_6_33_groupi_n_2867 ,csa_tree_add_6_33_groupi_n_2523 ,csa_tree_add_6_33_groupi_n_2513);
  nor csa_tree_add_6_33_groupi_g15422(csa_tree_add_6_33_groupi_n_2866 ,csa_tree_add_6_33_groupi_n_1376 ,csa_tree_add_6_33_groupi_n_2414);
  and csa_tree_add_6_33_groupi_g15423(csa_tree_add_6_33_groupi_n_2865 ,csa_tree_add_6_33_groupi_n_2424 ,csa_tree_add_6_33_groupi_n_2536);
  or csa_tree_add_6_33_groupi_g15424(csa_tree_add_6_33_groupi_n_2864 ,csa_tree_add_6_33_groupi_n_1888 ,csa_tree_add_6_33_groupi_n_2571);
  or csa_tree_add_6_33_groupi_g15425(csa_tree_add_6_33_groupi_n_2863 ,csa_tree_add_6_33_groupi_n_1375 ,csa_tree_add_6_33_groupi_n_2415);
  and csa_tree_add_6_33_groupi_g15426(csa_tree_add_6_33_groupi_n_2862 ,csa_tree_add_6_33_groupi_n_2523 ,csa_tree_add_6_33_groupi_n_2513);
  or csa_tree_add_6_33_groupi_g15427(csa_tree_add_6_33_groupi_n_2861 ,csa_tree_add_6_33_groupi_n_2532 ,csa_tree_add_6_33_groupi_n_2455);
  and csa_tree_add_6_33_groupi_g15428(csa_tree_add_6_33_groupi_n_2860 ,csa_tree_add_6_33_groupi_n_2532 ,csa_tree_add_6_33_groupi_n_2455);
  and csa_tree_add_6_33_groupi_g15429(csa_tree_add_6_33_groupi_n_2859 ,csa_tree_add_6_33_groupi_n_1072 ,csa_tree_add_6_33_groupi_n_2508);
  or csa_tree_add_6_33_groupi_g15430(csa_tree_add_6_33_groupi_n_2858 ,csa_tree_add_6_33_groupi_n_2439 ,csa_tree_add_6_33_groupi_n_2438);
  nor csa_tree_add_6_33_groupi_g15431(csa_tree_add_6_33_groupi_n_2857 ,csa_tree_add_6_33_groupi_n_1133 ,csa_tree_add_6_33_groupi_n_2398);
  and csa_tree_add_6_33_groupi_g15432(csa_tree_add_6_33_groupi_n_2856 ,csa_tree_add_6_33_groupi_n_2338 ,csa_tree_add_6_33_groupi_n_2419);
  or csa_tree_add_6_33_groupi_g15433(csa_tree_add_6_33_groupi_n_2855 ,csa_tree_add_6_33_groupi_n_2516 ,csa_tree_add_6_33_groupi_n_2511);
  or csa_tree_add_6_33_groupi_g15434(csa_tree_add_6_33_groupi_n_2854 ,csa_tree_add_6_33_groupi_n_2490 ,csa_tree_add_6_33_groupi_n_2548);
  nor csa_tree_add_6_33_groupi_g15435(csa_tree_add_6_33_groupi_n_2853 ,csa_tree_add_6_33_groupi_n_2337 ,csa_tree_add_6_33_groupi_n_2409);
  or csa_tree_add_6_33_groupi_g15436(csa_tree_add_6_33_groupi_n_2852 ,csa_tree_add_6_33_groupi_n_1134 ,csa_tree_add_6_33_groupi_n_2397);
  or csa_tree_add_6_33_groupi_g15437(csa_tree_add_6_33_groupi_n_2851 ,csa_tree_add_6_33_groupi_n_1417 ,csa_tree_add_6_33_groupi_n_2527);
  and csa_tree_add_6_33_groupi_g15438(csa_tree_add_6_33_groupi_n_2850 ,csa_tree_add_6_33_groupi_n_2516 ,csa_tree_add_6_33_groupi_n_2511);
  or csa_tree_add_6_33_groupi_g15439(csa_tree_add_6_33_groupi_n_2849 ,csa_tree_add_6_33_groupi_n_2506 ,csa_tree_add_6_33_groupi_n_2503);
  or csa_tree_add_6_33_groupi_g15440(csa_tree_add_6_33_groupi_n_2848 ,csa_tree_add_6_33_groupi_n_2535 ,csa_tree_add_6_33_groupi_n_2412);
  nor csa_tree_add_6_33_groupi_g15441(csa_tree_add_6_33_groupi_n_2847 ,csa_tree_add_6_33_groupi_n_2534 ,csa_tree_add_6_33_groupi_n_2413);
  and csa_tree_add_6_33_groupi_g15442(csa_tree_add_6_33_groupi_n_2846 ,csa_tree_add_6_33_groupi_n_2506 ,csa_tree_add_6_33_groupi_n_2503);
  and csa_tree_add_6_33_groupi_g15443(csa_tree_add_6_33_groupi_n_2845 ,csa_tree_add_6_33_groupi_n_2428 ,csa_tree_add_6_33_groupi_n_2385);
  or csa_tree_add_6_33_groupi_g15444(csa_tree_add_6_33_groupi_n_2844 ,csa_tree_add_6_33_groupi_n_1414 ,csa_tree_add_6_33_groupi_n_2410);
  nor csa_tree_add_6_33_groupi_g15445(csa_tree_add_6_33_groupi_n_2843 ,csa_tree_add_6_33_groupi_n_1413 ,csa_tree_add_6_33_groupi_n_2411);
  or csa_tree_add_6_33_groupi_g15446(csa_tree_add_6_33_groupi_n_2842 ,csa_tree_add_6_33_groupi_n_2424 ,csa_tree_add_6_33_groupi_n_2536);
  nor csa_tree_add_6_33_groupi_g15447(csa_tree_add_6_33_groupi_n_2841 ,csa_tree_add_6_33_groupi_n_2499 ,csa_tree_add_6_33_groupi_n_2391);
  or csa_tree_add_6_33_groupi_g15448(csa_tree_add_6_33_groupi_n_2840 ,csa_tree_add_6_33_groupi_n_1404 ,csa_tree_add_6_33_groupi_n_2529);
  or csa_tree_add_6_33_groupi_g15449(csa_tree_add_6_33_groupi_n_2839 ,csa_tree_add_6_33_groupi_n_2533 ,csa_tree_add_6_33_groupi_n_2448);
  or csa_tree_add_6_33_groupi_g15450(csa_tree_add_6_33_groupi_n_2838 ,csa_tree_add_6_33_groupi_n_1370 ,csa_tree_add_6_33_groupi_n_2435);
  and csa_tree_add_6_33_groupi_g15451(csa_tree_add_6_33_groupi_n_2837 ,csa_tree_add_6_33_groupi_n_2337 ,csa_tree_add_6_33_groupi_n_2409);
  or csa_tree_add_6_33_groupi_g15452(csa_tree_add_6_33_groupi_n_2836 ,csa_tree_add_6_33_groupi_n_1206 ,csa_tree_add_6_33_groupi_n_2530);
  nor csa_tree_add_6_33_groupi_g15453(csa_tree_add_6_33_groupi_n_2835 ,csa_tree_add_6_33_groupi_n_1519 ,csa_tree_add_6_33_groupi_n_2389);
  or csa_tree_add_6_33_groupi_g15454(csa_tree_add_6_33_groupi_n_2834 ,csa_tree_add_6_33_groupi_n_1518 ,csa_tree_add_6_33_groupi_n_2388);
  and csa_tree_add_6_33_groupi_g15455(csa_tree_add_6_33_groupi_n_2833 ,csa_tree_add_6_33_groupi_n_1404 ,csa_tree_add_6_33_groupi_n_2529);
  and csa_tree_add_6_33_groupi_g15456(csa_tree_add_6_33_groupi_n_2832 ,csa_tree_add_6_33_groupi_n_1743 ,csa_tree_add_6_33_groupi_n_2457);
  or csa_tree_add_6_33_groupi_g15457(csa_tree_add_6_33_groupi_n_2831 ,csa_tree_add_6_33_groupi_n_1919 ,csa_tree_add_6_33_groupi_n_2563);
  nor csa_tree_add_6_33_groupi_g15458(csa_tree_add_6_33_groupi_n_2830 ,csa_tree_add_6_33_groupi_n_2331 ,csa_tree_add_6_33_groupi_n_2387);
  or csa_tree_add_6_33_groupi_g15459(csa_tree_add_6_33_groupi_n_2829 ,csa_tree_add_6_33_groupi_n_1138 ,csa_tree_add_6_33_groupi_n_2405);
  or csa_tree_add_6_33_groupi_g15460(csa_tree_add_6_33_groupi_n_2828 ,csa_tree_add_6_33_groupi_n_1784 ,csa_tree_add_6_33_groupi_n_2578);
  nor csa_tree_add_6_33_groupi_g15461(csa_tree_add_6_33_groupi_n_2827 ,csa_tree_add_6_33_groupi_n_1137 ,csa_tree_add_6_33_groupi_n_2406);
  or csa_tree_add_6_33_groupi_g15462(csa_tree_add_6_33_groupi_n_2826 ,csa_tree_add_6_33_groupi_n_2501 ,csa_tree_add_6_33_groupi_n_2522);
  and csa_tree_add_6_33_groupi_g15463(csa_tree_add_6_33_groupi_n_2825 ,csa_tree_add_6_33_groupi_n_2501 ,csa_tree_add_6_33_groupi_n_2522);
  and csa_tree_add_6_33_groupi_g15464(csa_tree_add_6_33_groupi_n_2824 ,csa_tree_add_6_33_groupi_n_1370 ,csa_tree_add_6_33_groupi_n_2435);
  and csa_tree_add_6_33_groupi_g15465(csa_tree_add_6_33_groupi_n_2823 ,csa_tree_add_6_33_groupi_n_2525 ,csa_tree_add_6_33_groupi_n_2449);
  or csa_tree_add_6_33_groupi_g15466(csa_tree_add_6_33_groupi_n_2822 ,csa_tree_add_6_33_groupi_n_2345 ,csa_tree_add_6_33_groupi_n_2395);
  and csa_tree_add_6_33_groupi_g15467(csa_tree_add_6_33_groupi_n_2821 ,csa_tree_add_6_33_groupi_n_2339 ,csa_tree_add_6_33_groupi_n_2416);
  and csa_tree_add_6_33_groupi_g15468(csa_tree_add_6_33_groupi_n_2820 ,csa_tree_add_6_33_groupi_n_1206 ,csa_tree_add_6_33_groupi_n_2530);
  or csa_tree_add_6_33_groupi_g15469(csa_tree_add_6_33_groupi_n_2819 ,csa_tree_add_6_33_groupi_n_2498 ,csa_tree_add_6_33_groupi_n_2390);
  or csa_tree_add_6_33_groupi_g15470(csa_tree_add_6_33_groupi_n_2818 ,csa_tree_add_6_33_groupi_n_2512 ,csa_tree_add_6_33_groupi_n_2505);
  or csa_tree_add_6_33_groupi_g15471(csa_tree_add_6_33_groupi_n_2817 ,csa_tree_add_6_33_groupi_n_2487 ,csa_tree_add_6_33_groupi_n_2480);
  or csa_tree_add_6_33_groupi_g15472(csa_tree_add_6_33_groupi_n_2816 ,csa_tree_add_6_33_groupi_n_2507 ,csa_tree_add_6_33_groupi_n_2497);
  nor csa_tree_add_6_33_groupi_g15473(csa_tree_add_6_33_groupi_n_2815 ,csa_tree_add_6_33_groupi_n_2339 ,csa_tree_add_6_33_groupi_n_2416);
  and csa_tree_add_6_33_groupi_g15474(csa_tree_add_6_33_groupi_n_2814 ,csa_tree_add_6_33_groupi_n_2512 ,csa_tree_add_6_33_groupi_n_2505);
  and csa_tree_add_6_33_groupi_g15475(csa_tree_add_6_33_groupi_n_2813 ,csa_tree_add_6_33_groupi_n_1157 ,csa_tree_add_6_33_groupi_n_2422);
  or csa_tree_add_6_33_groupi_g15476(csa_tree_add_6_33_groupi_n_2812 ,csa_tree_add_6_33_groupi_n_1807 ,csa_tree_add_6_33_groupi_n_2537);
  or csa_tree_add_6_33_groupi_g15477(csa_tree_add_6_33_groupi_n_2811 ,csa_tree_add_6_33_groupi_n_1882 ,csa_tree_add_6_33_groupi_n_2538);
  or csa_tree_add_6_33_groupi_g15478(csa_tree_add_6_33_groupi_n_2810 ,csa_tree_add_6_33_groupi_n_2334 ,csa_tree_add_6_33_groupi_n_2495);
  and csa_tree_add_6_33_groupi_g15479(csa_tree_add_6_33_groupi_n_2809 ,csa_tree_add_6_33_groupi_n_2334 ,csa_tree_add_6_33_groupi_n_2495);
  or csa_tree_add_6_33_groupi_g15480(csa_tree_add_6_33_groupi_n_2808 ,csa_tree_add_6_33_groupi_n_2376 ,csa_tree_add_6_33_groupi_n_2393);
  or csa_tree_add_6_33_groupi_g15481(csa_tree_add_6_33_groupi_n_2807 ,csa_tree_add_6_33_groupi_n_2399 ,csa_tree_add_6_33_groupi_n_2403);
  or csa_tree_add_6_33_groupi_g15482(csa_tree_add_6_33_groupi_n_2806 ,csa_tree_add_6_33_groupi_n_2404 ,csa_tree_add_6_33_groupi_n_2407);
  and csa_tree_add_6_33_groupi_g15483(csa_tree_add_6_33_groupi_n_2805 ,csa_tree_add_6_33_groupi_n_2399 ,csa_tree_add_6_33_groupi_n_2403);
  or csa_tree_add_6_33_groupi_g15484(csa_tree_add_6_33_groupi_n_2804 ,csa_tree_add_6_33_groupi_n_1773 ,csa_tree_add_6_33_groupi_n_2473);
  and csa_tree_add_6_33_groupi_g15485(csa_tree_add_6_33_groupi_n_2803 ,csa_tree_add_6_33_groupi_n_2376 ,csa_tree_add_6_33_groupi_n_2393);
  and csa_tree_add_6_33_groupi_g15486(csa_tree_add_6_33_groupi_n_2802 ,csa_tree_add_6_33_groupi_n_2404 ,csa_tree_add_6_33_groupi_n_2407);
  or csa_tree_add_6_33_groupi_g15487(csa_tree_add_6_33_groupi_n_2801 ,csa_tree_add_6_33_groupi_n_2429 ,csa_tree_add_6_33_groupi_n_2384);
  and csa_tree_add_6_33_groupi_g15488(csa_tree_add_6_33_groupi_n_2800 ,csa_tree_add_6_33_groupi_n_2429 ,csa_tree_add_6_33_groupi_n_2384);
  or csa_tree_add_6_33_groupi_g15489(csa_tree_add_6_33_groupi_n_2799 ,csa_tree_add_6_33_groupi_n_2332 ,csa_tree_add_6_33_groupi_n_2434);
  or csa_tree_add_6_33_groupi_g15490(csa_tree_add_6_33_groupi_n_2798 ,csa_tree_add_6_33_groupi_n_2432 ,csa_tree_add_6_33_groupi_n_2436);
  nor csa_tree_add_6_33_groupi_g15491(csa_tree_add_6_33_groupi_n_2797 ,csa_tree_add_6_33_groupi_n_2333 ,csa_tree_add_6_33_groupi_n_2433);
  and csa_tree_add_6_33_groupi_g15492(csa_tree_add_6_33_groupi_n_2796 ,csa_tree_add_6_33_groupi_n_2432 ,csa_tree_add_6_33_groupi_n_2436);
  and csa_tree_add_6_33_groupi_g15493(csa_tree_add_6_33_groupi_n_2795 ,csa_tree_add_6_33_groupi_n_2453 ,csa_tree_add_6_33_groupi_n_2381);
  or csa_tree_add_6_33_groupi_g15494(csa_tree_add_6_33_groupi_n_2794 ,csa_tree_add_6_33_groupi_n_1481 ,csa_tree_add_6_33_groupi_n_2440);
  and csa_tree_add_6_33_groupi_g15495(csa_tree_add_6_33_groupi_n_2793 ,csa_tree_add_6_33_groupi_n_1091 ,csa_tree_add_6_33_groupi_n_2402);
  nor csa_tree_add_6_33_groupi_g15496(csa_tree_add_6_33_groupi_n_2792 ,csa_tree_add_6_33_groupi_n_1091 ,csa_tree_add_6_33_groupi_n_2402);
  or csa_tree_add_6_33_groupi_g15497(csa_tree_add_6_33_groupi_n_2791 ,csa_tree_add_6_33_groupi_n_2441 ,csa_tree_add_6_33_groupi_n_2444);
  and csa_tree_add_6_33_groupi_g15498(csa_tree_add_6_33_groupi_n_2790 ,csa_tree_add_6_33_groupi_n_1481 ,csa_tree_add_6_33_groupi_n_2440);
  and csa_tree_add_6_33_groupi_g15499(csa_tree_add_6_33_groupi_n_2789 ,csa_tree_add_6_33_groupi_n_2441 ,csa_tree_add_6_33_groupi_n_2444);
  or csa_tree_add_6_33_groupi_g15500(csa_tree_add_6_33_groupi_n_2788 ,csa_tree_add_6_33_groupi_n_1736 ,csa_tree_add_6_33_groupi_n_2461);
  or csa_tree_add_6_33_groupi_g15501(csa_tree_add_6_33_groupi_n_2787 ,csa_tree_add_6_33_groupi_n_2341 ,csa_tree_add_6_33_groupi_n_2383);
  and csa_tree_add_6_33_groupi_g15502(csa_tree_add_6_33_groupi_n_2786 ,csa_tree_add_6_33_groupi_n_2528 ,csa_tree_add_6_33_groupi_n_2524);
  and csa_tree_add_6_33_groupi_g15503(csa_tree_add_6_33_groupi_n_2785 ,csa_tree_add_6_33_groupi_n_1408 ,csa_tree_add_6_33_groupi_n_2392);
  and csa_tree_add_6_33_groupi_g15504(csa_tree_add_6_33_groupi_n_2784 ,csa_tree_add_6_33_groupi_n_2533 ,csa_tree_add_6_33_groupi_n_2448);
  or csa_tree_add_6_33_groupi_g15505(csa_tree_add_6_33_groupi_n_2783 ,csa_tree_add_6_33_groupi_n_1660 ,csa_tree_add_6_33_groupi_n_2459);
  or csa_tree_add_6_33_groupi_g15506(csa_tree_add_6_33_groupi_n_2782 ,csa_tree_add_6_33_groupi_n_2496 ,csa_tree_add_6_33_groupi_n_2380);
  or csa_tree_add_6_33_groupi_g15507(csa_tree_add_6_33_groupi_n_2781 ,csa_tree_add_6_33_groupi_n_1150 ,csa_tree_add_6_33_groupi_n_2452);
  or csa_tree_add_6_33_groupi_g15508(csa_tree_add_6_33_groupi_n_2780 ,csa_tree_add_6_33_groupi_n_2454 ,csa_tree_add_6_33_groupi_n_2451);
  and csa_tree_add_6_33_groupi_g15509(csa_tree_add_6_33_groupi_n_2779 ,csa_tree_add_6_33_groupi_n_2496 ,csa_tree_add_6_33_groupi_n_2380);
  or csa_tree_add_6_33_groupi_g15510(csa_tree_add_6_33_groupi_n_2778 ,csa_tree_add_6_33_groupi_n_2453 ,csa_tree_add_6_33_groupi_n_2381);
  and csa_tree_add_6_33_groupi_g15511(csa_tree_add_6_33_groupi_n_2777 ,csa_tree_add_6_33_groupi_n_2454 ,csa_tree_add_6_33_groupi_n_2451);
  or csa_tree_add_6_33_groupi_g15512(csa_tree_add_6_33_groupi_n_2776 ,csa_tree_add_6_33_groupi_n_2336 ,csa_tree_add_6_33_groupi_n_2447);
  and csa_tree_add_6_33_groupi_g15513(csa_tree_add_6_33_groupi_n_2775 ,csa_tree_add_6_33_groupi_n_2336 ,csa_tree_add_6_33_groupi_n_2447);
  or csa_tree_add_6_33_groupi_g15514(csa_tree_add_6_33_groupi_n_2774 ,csa_tree_add_6_33_groupi_n_2443 ,csa_tree_add_6_33_groupi_n_2400);
  nor csa_tree_add_6_33_groupi_g15515(csa_tree_add_6_33_groupi_n_2773 ,csa_tree_add_6_33_groupi_n_2442 ,csa_tree_add_6_33_groupi_n_2401);
  and csa_tree_add_6_33_groupi_g15516(csa_tree_add_6_33_groupi_n_2772 ,csa_tree_add_6_33_groupi_n_1150 ,csa_tree_add_6_33_groupi_n_2452);
  or csa_tree_add_6_33_groupi_g15517(csa_tree_add_6_33_groupi_n_2771 ,csa_tree_add_6_33_groupi_n_2373 ,csa_tree_add_6_33_groupi_n_2557);
  or csa_tree_add_6_33_groupi_g15518(csa_tree_add_6_33_groupi_n_2770 ,csa_tree_add_6_33_groupi_n_2423 ,csa_tree_add_6_33_groupi_n_2379);
  and csa_tree_add_6_33_groupi_g15519(csa_tree_add_6_33_groupi_n_2769 ,csa_tree_add_6_33_groupi_n_2423 ,csa_tree_add_6_33_groupi_n_2379);
  and csa_tree_add_6_33_groupi_g15520(csa_tree_add_6_33_groupi_n_2768 ,csa_tree_add_6_33_groupi_n_2507 ,csa_tree_add_6_33_groupi_n_2497);
  and csa_tree_add_6_33_groupi_g15521(csa_tree_add_6_33_groupi_n_2767 ,csa_tree_add_6_33_groupi_n_2439 ,csa_tree_add_6_33_groupi_n_2438);
  or csa_tree_add_6_33_groupi_g15522(csa_tree_add_6_33_groupi_n_2766 ,csa_tree_add_6_33_groupi_n_2343 ,csa_tree_add_6_33_groupi_n_2378);
  nor csa_tree_add_6_33_groupi_g15523(csa_tree_add_6_33_groupi_n_2765 ,csa_tree_add_6_33_groupi_n_2344 ,csa_tree_add_6_33_groupi_n_2377);
  or csa_tree_add_6_33_groupi_g15524(csa_tree_add_6_33_groupi_n_2764 ,csa_tree_add_6_33_groupi_n_1924 ,csa_tree_add_6_33_groupi_n_2469);
  or csa_tree_add_6_33_groupi_g15525(csa_tree_add_6_33_groupi_n_2763 ,csa_tree_add_6_33_groupi_n_2431 ,csa_tree_add_6_33_groupi_n_2430);
  and csa_tree_add_6_33_groupi_g15526(csa_tree_add_6_33_groupi_n_2762 ,csa_tree_add_6_33_groupi_n_2431 ,csa_tree_add_6_33_groupi_n_2430);
  or csa_tree_add_6_33_groupi_g15527(csa_tree_add_6_33_groupi_n_2761 ,csa_tree_add_6_33_groupi_n_1145 ,csa_tree_add_6_33_groupi_n_2515);
  or csa_tree_add_6_33_groupi_g15528(csa_tree_add_6_33_groupi_n_2760 ,csa_tree_add_6_33_groupi_n_2428 ,csa_tree_add_6_33_groupi_n_2385);
  nor csa_tree_add_6_33_groupi_g15529(csa_tree_add_6_33_groupi_n_2759 ,csa_tree_add_6_33_groupi_n_2346 ,csa_tree_add_6_33_groupi_n_2394);
  and csa_tree_add_6_33_groupi_g15530(csa_tree_add_6_33_groupi_n_2758 ,csa_tree_add_6_33_groupi_n_1145 ,csa_tree_add_6_33_groupi_n_2515);
  xor csa_tree_add_6_33_groupi_g15531(csa_tree_add_6_33_groupi_n_2757 ,csa_tree_add_6_33_groupi_n_1408 ,csa_tree_add_6_33_groupi_n_2363);
  xnor csa_tree_add_6_33_groupi_g15532(csa_tree_add_6_33_groupi_n_2756 ,csa_tree_add_6_33_groupi_n_1143 ,csa_tree_add_6_33_groupi_n_2326);
  or csa_tree_add_6_33_groupi_g15533(csa_tree_add_6_33_groupi_n_2915 ,csa_tree_add_6_33_groupi_n_1885 ,csa_tree_add_6_33_groupi_n_2374);
  xnor csa_tree_add_6_33_groupi_g15534(csa_tree_add_6_33_groupi_n_2913 ,csa_tree_add_6_33_groupi_n_1365 ,csa_tree_add_6_33_groupi_n_2171);
  and csa_tree_add_6_33_groupi_g15535(csa_tree_add_6_33_groupi_n_2912 ,csa_tree_add_6_33_groupi_n_1347 ,csa_tree_add_6_33_groupi_n_2493);
  and csa_tree_add_6_33_groupi_g15536(csa_tree_add_6_33_groupi_n_2910 ,csa_tree_add_6_33_groupi_n_1855 ,csa_tree_add_6_33_groupi_n_2489);
  and csa_tree_add_6_33_groupi_g15537(csa_tree_add_6_33_groupi_n_2908 ,csa_tree_add_6_33_groupi_n_1902 ,csa_tree_add_6_33_groupi_n_2370);
  xnor csa_tree_add_6_33_groupi_g15538(csa_tree_add_6_33_groupi_n_2907 ,csa_tree_add_6_33_groupi_n_2353 ,csa_tree_add_6_33_groupi_n_2117);
  xnor csa_tree_add_6_33_groupi_g15539(csa_tree_add_6_33_groupi_n_2905 ,csa_tree_add_6_33_groupi_n_1440 ,csa_tree_add_6_33_groupi_n_2096);
  and csa_tree_add_6_33_groupi_g15540(csa_tree_add_6_33_groupi_n_2902 ,csa_tree_add_6_33_groupi_n_1749 ,csa_tree_add_6_33_groupi_n_2491);
  or csa_tree_add_6_33_groupi_g15541(csa_tree_add_6_33_groupi_n_2900 ,csa_tree_add_6_33_groupi_n_1704 ,csa_tree_add_6_33_groupi_n_2488);
  xnor csa_tree_add_6_33_groupi_g15542(csa_tree_add_6_33_groupi_n_2899 ,csa_tree_add_6_33_groupi_n_1388 ,csa_tree_add_6_33_groupi_n_2168);
  xnor csa_tree_add_6_33_groupi_g15543(csa_tree_add_6_33_groupi_n_2897 ,csa_tree_add_6_33_groupi_n_2367 ,csa_tree_add_6_33_groupi_n_2155);
  xnor csa_tree_add_6_33_groupi_g15544(csa_tree_add_6_33_groupi_n_2896 ,csa_tree_add_6_33_groupi_n_2360 ,csa_tree_add_6_33_groupi_n_2129);
  xnor csa_tree_add_6_33_groupi_g15545(csa_tree_add_6_33_groupi_n_2894 ,csa_tree_add_6_33_groupi_n_1494 ,csa_tree_add_6_33_groupi_n_2169);
  xnor csa_tree_add_6_33_groupi_g15546(csa_tree_add_6_33_groupi_n_2892 ,csa_tree_add_6_33_groupi_n_1407 ,csa_tree_add_6_33_groupi_n_2174);
  or csa_tree_add_6_33_groupi_g15547(csa_tree_add_6_33_groupi_n_2889 ,csa_tree_add_6_33_groupi_n_1953 ,csa_tree_add_6_33_groupi_n_2485);
  and csa_tree_add_6_33_groupi_g15548(csa_tree_add_6_33_groupi_n_2888 ,csa_tree_add_6_33_groupi_n_1838 ,csa_tree_add_6_33_groupi_n_2492);
  not csa_tree_add_6_33_groupi_g15549(csa_tree_add_6_33_groupi_n_2725 ,csa_tree_add_6_33_groupi_n_2724);
  not csa_tree_add_6_33_groupi_g15550(csa_tree_add_6_33_groupi_n_2717 ,csa_tree_add_6_33_groupi_n_2718);
  not csa_tree_add_6_33_groupi_g15551(csa_tree_add_6_33_groupi_n_2714 ,csa_tree_add_6_33_groupi_n_2715);
  not csa_tree_add_6_33_groupi_g15552(csa_tree_add_6_33_groupi_n_2709 ,csa_tree_add_6_33_groupi_n_2710);
  not csa_tree_add_6_33_groupi_g15553(csa_tree_add_6_33_groupi_n_2705 ,csa_tree_add_6_33_groupi_n_2706);
  not csa_tree_add_6_33_groupi_g15554(csa_tree_add_6_33_groupi_n_2702 ,csa_tree_add_6_33_groupi_n_2703);
  not csa_tree_add_6_33_groupi_g15555(csa_tree_add_6_33_groupi_n_2697 ,csa_tree_add_6_33_groupi_n_2698);
  not csa_tree_add_6_33_groupi_g15556(csa_tree_add_6_33_groupi_n_2695 ,csa_tree_add_6_33_groupi_n_2696);
  not csa_tree_add_6_33_groupi_g15557(csa_tree_add_6_33_groupi_n_2693 ,csa_tree_add_6_33_groupi_n_2694);
  not csa_tree_add_6_33_groupi_g15558(csa_tree_add_6_33_groupi_n_2691 ,csa_tree_add_6_33_groupi_n_2690);
  not csa_tree_add_6_33_groupi_g15559(csa_tree_add_6_33_groupi_n_2681 ,csa_tree_add_6_33_groupi_n_2680);
  not csa_tree_add_6_33_groupi_g15560(csa_tree_add_6_33_groupi_n_2673 ,csa_tree_add_6_33_groupi_n_2674);
  not csa_tree_add_6_33_groupi_g15561(csa_tree_add_6_33_groupi_n_2670 ,csa_tree_add_6_33_groupi_n_2671);
  not csa_tree_add_6_33_groupi_g15563(csa_tree_add_6_33_groupi_n_2667 ,csa_tree_add_6_33_groupi_n_2668);
  not csa_tree_add_6_33_groupi_g15564(csa_tree_add_6_33_groupi_n_2664 ,csa_tree_add_6_33_groupi_n_2665);
  not csa_tree_add_6_33_groupi_g15565(csa_tree_add_6_33_groupi_n_2643 ,csa_tree_add_6_33_groupi_n_2644);
  not csa_tree_add_6_33_groupi_g15566(csa_tree_add_6_33_groupi_n_2640 ,csa_tree_add_6_33_groupi_n_2641);
  not csa_tree_add_6_33_groupi_g15567(csa_tree_add_6_33_groupi_n_2637 ,csa_tree_add_6_33_groupi_n_2638);
  not csa_tree_add_6_33_groupi_g15568(csa_tree_add_6_33_groupi_n_2631 ,csa_tree_add_6_33_groupi_n_2632);
  not csa_tree_add_6_33_groupi_g15569(csa_tree_add_6_33_groupi_n_2624 ,csa_tree_add_6_33_groupi_n_2625);
  not csa_tree_add_6_33_groupi_g15570(csa_tree_add_6_33_groupi_n_2618 ,csa_tree_add_6_33_groupi_n_2619);
  not csa_tree_add_6_33_groupi_g15571(csa_tree_add_6_33_groupi_n_2613 ,csa_tree_add_6_33_groupi_n_2614);
  not csa_tree_add_6_33_groupi_g15572(csa_tree_add_6_33_groupi_n_2601 ,csa_tree_add_6_33_groupi_n_2602);
  not csa_tree_add_6_33_groupi_g15573(csa_tree_add_6_33_groupi_n_2589 ,csa_tree_add_6_33_groupi_n_2590);
  xnor csa_tree_add_6_33_groupi_g15574(out1[1] ,csa_tree_add_6_33_groupi_n_2358 ,csa_tree_add_6_33_groupi_n_1625);
  xnor csa_tree_add_6_33_groupi_g15575(csa_tree_add_6_33_groupi_n_2586 ,csa_tree_add_6_33_groupi_n_1484 ,csa_tree_add_6_33_groupi_n_2351);
  xnor csa_tree_add_6_33_groupi_g15576(csa_tree_add_6_33_groupi_n_2585 ,csa_tree_add_6_33_groupi_n_1091 ,csa_tree_add_6_33_groupi_n_2366);
  xnor csa_tree_add_6_33_groupi_g15577(csa_tree_add_6_33_groupi_n_2584 ,csa_tree_add_6_33_groupi_n_1410 ,csa_tree_add_6_33_groupi_n_2329);
  xnor csa_tree_add_6_33_groupi_g15578(csa_tree_add_6_33_groupi_n_2583 ,csa_tree_add_6_33_groupi_n_1519 ,csa_tree_add_6_33_groupi_n_2352);
  xnor csa_tree_add_6_33_groupi_g15579(csa_tree_add_6_33_groupi_n_2755 ,csa_tree_add_6_33_groupi_n_1227 ,csa_tree_add_6_33_groupi_n_2062);
  xor csa_tree_add_6_33_groupi_g15580(csa_tree_add_6_33_groupi_n_2754 ,csa_tree_add_6_33_groupi_n_1524 ,csa_tree_add_6_33_groupi_n_2165);
  xnor csa_tree_add_6_33_groupi_g15581(csa_tree_add_6_33_groupi_n_2753 ,csa_tree_add_6_33_groupi_n_1123 ,csa_tree_add_6_33_groupi_n_2101);
  xnor csa_tree_add_6_33_groupi_g15582(csa_tree_add_6_33_groupi_n_2752 ,csa_tree_add_6_33_groupi_n_1386 ,csa_tree_add_6_33_groupi_n_2114);
  xnor csa_tree_add_6_33_groupi_g15583(csa_tree_add_6_33_groupi_n_2751 ,csa_tree_add_6_33_groupi_n_1374 ,csa_tree_add_6_33_groupi_n_2143);
  xnor csa_tree_add_6_33_groupi_g15584(csa_tree_add_6_33_groupi_n_2750 ,csa_tree_add_6_33_groupi_n_1540 ,csa_tree_add_6_33_groupi_n_2154);
  xnor csa_tree_add_6_33_groupi_g15585(csa_tree_add_6_33_groupi_n_2749 ,csa_tree_add_6_33_groupi_n_1096 ,csa_tree_add_6_33_groupi_n_2160);
  xnor csa_tree_add_6_33_groupi_g15586(csa_tree_add_6_33_groupi_n_2748 ,csa_tree_add_6_33_groupi_n_1297 ,csa_tree_add_6_33_groupi_n_2124);
  xnor csa_tree_add_6_33_groupi_g15587(csa_tree_add_6_33_groupi_n_2747 ,csa_tree_add_6_33_groupi_n_1144 ,csa_tree_add_6_33_groupi_n_2111);
  xnor csa_tree_add_6_33_groupi_g15588(csa_tree_add_6_33_groupi_n_2746 ,csa_tree_add_6_33_groupi_n_1579 ,csa_tree_add_6_33_groupi_n_2103);
  xnor csa_tree_add_6_33_groupi_g15589(csa_tree_add_6_33_groupi_n_2745 ,csa_tree_add_6_33_groupi_n_1232 ,csa_tree_add_6_33_groupi_n_2150);
  xnor csa_tree_add_6_33_groupi_g15590(csa_tree_add_6_33_groupi_n_2744 ,csa_tree_add_6_33_groupi_n_1149 ,csa_tree_add_6_33_groupi_n_2106);
  xnor csa_tree_add_6_33_groupi_g15591(csa_tree_add_6_33_groupi_n_2743 ,csa_tree_add_6_33_groupi_n_1505 ,csa_tree_add_6_33_groupi_n_2016);
  xnor csa_tree_add_6_33_groupi_g15592(csa_tree_add_6_33_groupi_n_2742 ,csa_tree_add_6_33_groupi_n_1463 ,csa_tree_add_6_33_groupi_n_2133);
  xnor csa_tree_add_6_33_groupi_g15593(csa_tree_add_6_33_groupi_n_2741 ,csa_tree_add_6_33_groupi_n_1170 ,csa_tree_add_6_33_groupi_n_2086);
  xnor csa_tree_add_6_33_groupi_g15594(csa_tree_add_6_33_groupi_n_2740 ,csa_tree_add_6_33_groupi_n_1169 ,csa_tree_add_6_33_groupi_n_2122);
  xnor csa_tree_add_6_33_groupi_g15595(csa_tree_add_6_33_groupi_n_2739 ,csa_tree_add_6_33_groupi_n_2364 ,csa_tree_add_6_33_groupi_n_2108);
  xnor csa_tree_add_6_33_groupi_g15596(csa_tree_add_6_33_groupi_n_2738 ,csa_tree_add_6_33_groupi_n_1438 ,csa_tree_add_6_33_groupi_n_2090);
  xnor csa_tree_add_6_33_groupi_g15597(csa_tree_add_6_33_groupi_n_2737 ,csa_tree_add_6_33_groupi_n_1105 ,csa_tree_add_6_33_groupi_n_2120);
  xnor csa_tree_add_6_33_groupi_g15598(csa_tree_add_6_33_groupi_n_2736 ,csa_tree_add_6_33_groupi_n_1368 ,csa_tree_add_6_33_groupi_n_2057);
  xnor csa_tree_add_6_33_groupi_g15599(csa_tree_add_6_33_groupi_n_2735 ,csa_tree_add_6_33_groupi_n_1378 ,csa_tree_add_6_33_groupi_n_2082);
  xnor csa_tree_add_6_33_groupi_g15600(csa_tree_add_6_33_groupi_n_2734 ,csa_tree_add_6_33_groupi_n_1070 ,csa_tree_add_6_33_groupi_n_2054);
  xnor csa_tree_add_6_33_groupi_g15601(csa_tree_add_6_33_groupi_n_2733 ,csa_tree_add_6_33_groupi_n_1155 ,csa_tree_add_6_33_groupi_n_2051);
  xnor csa_tree_add_6_33_groupi_g15602(csa_tree_add_6_33_groupi_n_2732 ,csa_tree_add_6_33_groupi_n_1500 ,csa_tree_add_6_33_groupi_n_2094);
  xnor csa_tree_add_6_33_groupi_g15603(csa_tree_add_6_33_groupi_n_2731 ,csa_tree_add_6_33_groupi_n_1373 ,csa_tree_add_6_33_groupi_n_2142);
  xnor csa_tree_add_6_33_groupi_g15604(csa_tree_add_6_33_groupi_n_2730 ,csa_tree_add_6_33_groupi_n_1468 ,csa_tree_add_6_33_groupi_n_2022);
  xnor csa_tree_add_6_33_groupi_g15605(csa_tree_add_6_33_groupi_n_2729 ,csa_tree_add_6_33_groupi_n_1475 ,csa_tree_add_6_33_groupi_n_2027);
  xnor csa_tree_add_6_33_groupi_g15606(csa_tree_add_6_33_groupi_n_2728 ,csa_tree_add_6_33_groupi_n_1081 ,csa_tree_add_6_33_groupi_n_2042);
  xnor csa_tree_add_6_33_groupi_g15607(csa_tree_add_6_33_groupi_n_2727 ,csa_tree_add_6_33_groupi_n_1447 ,csa_tree_add_6_33_groupi_n_2041);
  xnor csa_tree_add_6_33_groupi_g15608(csa_tree_add_6_33_groupi_n_2726 ,csa_tree_add_6_33_groupi_n_1544 ,csa_tree_add_6_33_groupi_n_2147);
  xnor csa_tree_add_6_33_groupi_g15609(csa_tree_add_6_33_groupi_n_2724 ,csa_tree_add_6_33_groupi_n_2368 ,csa_tree_add_6_33_groupi_n_2045);
  xor csa_tree_add_6_33_groupi_g15610(csa_tree_add_6_33_groupi_n_2723 ,csa_tree_add_6_33_groupi_n_1152 ,csa_tree_add_6_33_groupi_n_2170);
  xnor csa_tree_add_6_33_groupi_g15611(csa_tree_add_6_33_groupi_n_2722 ,csa_tree_add_6_33_groupi_n_1307 ,csa_tree_add_6_33_groupi_n_2089);
  xnor csa_tree_add_6_33_groupi_g15612(csa_tree_add_6_33_groupi_n_2721 ,csa_tree_add_6_33_groupi_n_1082 ,csa_tree_add_6_33_groupi_n_2034);
  xnor csa_tree_add_6_33_groupi_g15613(csa_tree_add_6_33_groupi_n_2720 ,csa_tree_add_6_33_groupi_n_1270 ,csa_tree_add_6_33_groupi_n_2163);
  xnor csa_tree_add_6_33_groupi_g15614(csa_tree_add_6_33_groupi_n_2719 ,csa_tree_add_6_33_groupi_n_1398 ,csa_tree_add_6_33_groupi_n_2138);
  xnor csa_tree_add_6_33_groupi_g15615(csa_tree_add_6_33_groupi_n_2718 ,csa_tree_add_6_33_groupi_n_1125 ,csa_tree_add_6_33_groupi_n_2014);
  xnor csa_tree_add_6_33_groupi_g15616(csa_tree_add_6_33_groupi_n_2716 ,csa_tree_add_6_33_groupi_n_1257 ,csa_tree_add_6_33_groupi_n_2099);
  xnor csa_tree_add_6_33_groupi_g15617(csa_tree_add_6_33_groupi_n_2715 ,csa_tree_add_6_33_groupi_n_1496 ,csa_tree_add_6_33_groupi_n_2172);
  xnor csa_tree_add_6_33_groupi_g15618(csa_tree_add_6_33_groupi_n_2713 ,csa_tree_add_6_33_groupi_n_1211 ,csa_tree_add_6_33_groupi_n_2048);
  xnor csa_tree_add_6_33_groupi_g15619(csa_tree_add_6_33_groupi_n_2712 ,csa_tree_add_6_33_groupi_n_1576 ,csa_tree_add_6_33_groupi_n_2119);
  xnor csa_tree_add_6_33_groupi_g15620(csa_tree_add_6_33_groupi_n_2711 ,csa_tree_add_6_33_groupi_n_1419 ,csa_tree_add_6_33_groupi_n_2098);
  xnor csa_tree_add_6_33_groupi_g15621(csa_tree_add_6_33_groupi_n_2710 ,csa_tree_add_6_33_groupi_n_1585 ,csa_tree_add_6_33_groupi_n_2130);
  xnor csa_tree_add_6_33_groupi_g15622(csa_tree_add_6_33_groupi_n_2708 ,csa_tree_add_6_33_groupi_n_1165 ,csa_tree_add_6_33_groupi_n_2127);
  xnor csa_tree_add_6_33_groupi_g15623(csa_tree_add_6_33_groupi_n_2707 ,csa_tree_add_6_33_groupi_n_1101 ,csa_tree_add_6_33_groupi_n_2140);
  xnor csa_tree_add_6_33_groupi_g15624(csa_tree_add_6_33_groupi_n_2706 ,csa_tree_add_6_33_groupi_n_1391 ,csa_tree_add_6_33_groupi_n_2178);
  xnor csa_tree_add_6_33_groupi_g15625(csa_tree_add_6_33_groupi_n_2704 ,csa_tree_add_6_33_groupi_n_1119 ,csa_tree_add_6_33_groupi_n_2126);
  xnor csa_tree_add_6_33_groupi_g15626(csa_tree_add_6_33_groupi_n_2703 ,csa_tree_add_6_33_groupi_n_1228 ,csa_tree_add_6_33_groupi_n_2020);
  xnor csa_tree_add_6_33_groupi_g15627(csa_tree_add_6_33_groupi_n_2701 ,csa_tree_add_6_33_groupi_n_1212 ,csa_tree_add_6_33_groupi_n_2040);
  xnor csa_tree_add_6_33_groupi_g15628(csa_tree_add_6_33_groupi_n_2700 ,csa_tree_add_6_33_groupi_n_1282 ,csa_tree_add_6_33_groupi_n_2039);
  xnor csa_tree_add_6_33_groupi_g15629(csa_tree_add_6_33_groupi_n_2699 ,csa_tree_add_6_33_groupi_n_1504 ,csa_tree_add_6_33_groupi_n_2123);
  xnor csa_tree_add_6_33_groupi_g15630(csa_tree_add_6_33_groupi_n_2698 ,csa_tree_add_6_33_groupi_n_1225 ,csa_tree_add_6_33_groupi_n_2167);
  xnor csa_tree_add_6_33_groupi_g15631(csa_tree_add_6_33_groupi_n_2696 ,csa_tree_add_6_33_groupi_n_1098 ,csa_tree_add_6_33_groupi_n_2176);
  xnor csa_tree_add_6_33_groupi_g15632(csa_tree_add_6_33_groupi_n_2694 ,csa_tree_add_6_33_groupi_n_1136 ,csa_tree_add_6_33_groupi_n_2173);
  xnor csa_tree_add_6_33_groupi_g15633(csa_tree_add_6_33_groupi_n_2692 ,csa_tree_add_6_33_groupi_n_1551 ,csa_tree_add_6_33_groupi_n_2121);
  xnor csa_tree_add_6_33_groupi_g15634(csa_tree_add_6_33_groupi_n_2690 ,csa_tree_add_6_33_groupi_n_2357 ,csa_tree_add_6_33_groupi_n_2097);
  xnor csa_tree_add_6_33_groupi_g15635(csa_tree_add_6_33_groupi_n_2689 ,csa_tree_add_6_33_groupi_n_1427 ,csa_tree_add_6_33_groupi_n_2113);
  xnor csa_tree_add_6_33_groupi_g15636(csa_tree_add_6_33_groupi_n_2688 ,csa_tree_add_6_33_groupi_n_1562 ,csa_tree_add_6_33_groupi_n_2164);
  xnor csa_tree_add_6_33_groupi_g15637(csa_tree_add_6_33_groupi_n_2687 ,csa_tree_add_6_33_groupi_n_1079 ,csa_tree_add_6_33_groupi_n_2112);
  xnor csa_tree_add_6_33_groupi_g15638(csa_tree_add_6_33_groupi_n_2686 ,csa_tree_add_6_33_groupi_n_1236 ,csa_tree_add_6_33_groupi_n_2093);
  xnor csa_tree_add_6_33_groupi_g15639(csa_tree_add_6_33_groupi_n_2685 ,csa_tree_add_6_33_groupi_n_1617 ,csa_tree_add_6_33_groupi_n_2132);
  xnor csa_tree_add_6_33_groupi_g15640(csa_tree_add_6_33_groupi_n_2684 ,csa_tree_add_6_33_groupi_n_1405 ,csa_tree_add_6_33_groupi_n_2066);
  xnor csa_tree_add_6_33_groupi_g15641(csa_tree_add_6_33_groupi_n_2683 ,csa_tree_add_6_33_groupi_n_1390 ,csa_tree_add_6_33_groupi_n_2104);
  xnor csa_tree_add_6_33_groupi_g15642(csa_tree_add_6_33_groupi_n_2682 ,csa_tree_add_6_33_groupi_n_1364 ,csa_tree_add_6_33_groupi_n_2092);
  xnor csa_tree_add_6_33_groupi_g15643(csa_tree_add_6_33_groupi_n_2680 ,csa_tree_add_6_33_groupi_n_2362 ,csa_tree_add_6_33_groupi_n_2141);
  xnor csa_tree_add_6_33_groupi_g15644(csa_tree_add_6_33_groupi_n_2679 ,csa_tree_add_6_33_groupi_n_1605 ,csa_tree_add_6_33_groupi_n_2102);
  xnor csa_tree_add_6_33_groupi_g15645(csa_tree_add_6_33_groupi_n_2678 ,csa_tree_add_6_33_groupi_n_1444 ,csa_tree_add_6_33_groupi_n_2032);
  xnor csa_tree_add_6_33_groupi_g15646(csa_tree_add_6_33_groupi_n_2677 ,csa_tree_add_6_33_groupi_n_1162 ,csa_tree_add_6_33_groupi_n_2087);
  xor csa_tree_add_6_33_groupi_g15647(csa_tree_add_6_33_groupi_n_2676 ,csa_tree_add_6_33_groupi_n_1537 ,csa_tree_add_6_33_groupi_n_2083);
  xnor csa_tree_add_6_33_groupi_g15648(csa_tree_add_6_33_groupi_n_2675 ,csa_tree_add_6_33_groupi_n_1531 ,csa_tree_add_6_33_groupi_n_2137);
  xnor csa_tree_add_6_33_groupi_g15649(csa_tree_add_6_33_groupi_n_2674 ,csa_tree_add_6_33_groupi_n_1369 ,csa_tree_add_6_33_groupi_n_2134);
  xnor csa_tree_add_6_33_groupi_g15650(csa_tree_add_6_33_groupi_n_2672 ,csa_tree_add_6_33_groupi_n_1382 ,csa_tree_add_6_33_groupi_n_2125);
  xnor csa_tree_add_6_33_groupi_g15651(csa_tree_add_6_33_groupi_n_2671 ,csa_tree_add_6_33_groupi_n_1071 ,csa_tree_add_6_33_groupi_n_2100);
  xnor csa_tree_add_6_33_groupi_g15652(csa_tree_add_6_33_groupi_n_2669 ,csa_tree_add_6_33_groupi_n_1596 ,csa_tree_add_6_33_groupi_n_2128);
  xnor csa_tree_add_6_33_groupi_g15653(csa_tree_add_6_33_groupi_n_2668 ,csa_tree_add_6_33_groupi_n_1076 ,csa_tree_add_6_33_groupi_n_2085);
  xnor csa_tree_add_6_33_groupi_g15654(csa_tree_add_6_33_groupi_n_2666 ,csa_tree_add_6_33_groupi_n_1415 ,csa_tree_add_6_33_groupi_n_2088);
  xnor csa_tree_add_6_33_groupi_g15655(csa_tree_add_6_33_groupi_n_2665 ,csa_tree_add_6_33_groupi_n_1177 ,csa_tree_add_6_33_groupi_n_2175);
  xnor csa_tree_add_6_33_groupi_g15656(csa_tree_add_6_33_groupi_n_2663 ,csa_tree_add_6_33_groupi_n_1516 ,csa_tree_add_6_33_groupi_n_2161);
  xnor csa_tree_add_6_33_groupi_g15657(csa_tree_add_6_33_groupi_n_2662 ,csa_tree_add_6_33_groupi_n_1197 ,csa_tree_add_6_33_groupi_n_2091);
  xnor csa_tree_add_6_33_groupi_g15658(csa_tree_add_6_33_groupi_n_2661 ,csa_tree_add_6_33_groupi_n_1377 ,csa_tree_add_6_33_groupi_n_2076);
  xnor csa_tree_add_6_33_groupi_g15659(csa_tree_add_6_33_groupi_n_2660 ,csa_tree_add_6_33_groupi_n_1471 ,csa_tree_add_6_33_groupi_n_2078);
  xnor csa_tree_add_6_33_groupi_g15660(csa_tree_add_6_33_groupi_n_2659 ,csa_tree_add_6_33_groupi_n_1190 ,csa_tree_add_6_33_groupi_n_2075);
  xnor csa_tree_add_6_33_groupi_g15661(csa_tree_add_6_33_groupi_n_2658 ,csa_tree_add_6_33_groupi_n_1115 ,csa_tree_add_6_33_groupi_n_2069);
  xnor csa_tree_add_6_33_groupi_g15662(csa_tree_add_6_33_groupi_n_2657 ,csa_tree_add_6_33_groupi_n_1480 ,csa_tree_add_6_33_groupi_n_2074);
  xnor csa_tree_add_6_33_groupi_g15663(csa_tree_add_6_33_groupi_n_2656 ,csa_tree_add_6_33_groupi_n_1194 ,csa_tree_add_6_33_groupi_n_2073);
  xnor csa_tree_add_6_33_groupi_g15664(csa_tree_add_6_33_groupi_n_2655 ,csa_tree_add_6_33_groupi_n_1528 ,csa_tree_add_6_33_groupi_n_2052);
  xnor csa_tree_add_6_33_groupi_g15665(csa_tree_add_6_33_groupi_n_2654 ,csa_tree_add_6_33_groupi_n_1502 ,csa_tree_add_6_33_groupi_n_2072);
  xnor csa_tree_add_6_33_groupi_g15666(csa_tree_add_6_33_groupi_n_2653 ,csa_tree_add_6_33_groupi_n_1501 ,csa_tree_add_6_33_groupi_n_2068);
  xnor csa_tree_add_6_33_groupi_g15667(csa_tree_add_6_33_groupi_n_2652 ,csa_tree_add_6_33_groupi_n_1487 ,csa_tree_add_6_33_groupi_n_2067);
  xnor csa_tree_add_6_33_groupi_g15668(csa_tree_add_6_33_groupi_n_2651 ,csa_tree_add_6_33_groupi_n_1180 ,csa_tree_add_6_33_groupi_n_2071);
  xnor csa_tree_add_6_33_groupi_g15669(csa_tree_add_6_33_groupi_n_2650 ,csa_tree_add_6_33_groupi_n_1478 ,csa_tree_add_6_33_groupi_n_2047);
  xnor csa_tree_add_6_33_groupi_g15670(csa_tree_add_6_33_groupi_n_2649 ,csa_tree_add_6_33_groupi_n_1550 ,csa_tree_add_6_33_groupi_n_2081);
  xnor csa_tree_add_6_33_groupi_g15671(csa_tree_add_6_33_groupi_n_2648 ,csa_tree_add_6_33_groupi_n_1112 ,csa_tree_add_6_33_groupi_n_2065);
  xnor csa_tree_add_6_33_groupi_g15672(csa_tree_add_6_33_groupi_n_2647 ,csa_tree_add_6_33_groupi_n_1184 ,csa_tree_add_6_33_groupi_n_2064);
  xnor csa_tree_add_6_33_groupi_g15673(csa_tree_add_6_33_groupi_n_2646 ,csa_tree_add_6_33_groupi_n_1538 ,csa_tree_add_6_33_groupi_n_2080);
  xnor csa_tree_add_6_33_groupi_g15674(csa_tree_add_6_33_groupi_n_2645 ,csa_tree_add_6_33_groupi_n_1428 ,csa_tree_add_6_33_groupi_n_2061);
  xnor csa_tree_add_6_33_groupi_g15675(csa_tree_add_6_33_groupi_n_2644 ,csa_tree_add_6_33_groupi_n_1418 ,csa_tree_add_6_33_groupi_n_2107);
  xnor csa_tree_add_6_33_groupi_g15676(csa_tree_add_6_33_groupi_n_2642 ,csa_tree_add_6_33_groupi_n_1485 ,csa_tree_add_6_33_groupi_n_2058);
  xnor csa_tree_add_6_33_groupi_g15677(csa_tree_add_6_33_groupi_n_2641 ,csa_tree_add_6_33_groupi_n_1433 ,csa_tree_add_6_33_groupi_n_2056);
  xnor csa_tree_add_6_33_groupi_g15678(csa_tree_add_6_33_groupi_n_2639 ,csa_tree_add_6_33_groupi_n_1156 ,csa_tree_add_6_33_groupi_n_2055);
  xnor csa_tree_add_6_33_groupi_g15679(csa_tree_add_6_33_groupi_n_2638 ,csa_tree_add_6_33_groupi_n_1131 ,csa_tree_add_6_33_groupi_n_2166);
  xnor csa_tree_add_6_33_groupi_g15680(csa_tree_add_6_33_groupi_n_2636 ,csa_tree_add_6_33_groupi_n_1449 ,csa_tree_add_6_33_groupi_n_2148);
  xnor csa_tree_add_6_33_groupi_g15681(csa_tree_add_6_33_groupi_n_2635 ,csa_tree_add_6_33_groupi_n_1103 ,csa_tree_add_6_33_groupi_n_2021);
  xnor csa_tree_add_6_33_groupi_g15682(csa_tree_add_6_33_groupi_n_2634 ,csa_tree_add_6_33_groupi_n_1244 ,csa_tree_add_6_33_groupi_n_2019);
  xnor csa_tree_add_6_33_groupi_g15683(csa_tree_add_6_33_groupi_n_2633 ,csa_tree_add_6_33_groupi_n_1283 ,csa_tree_add_6_33_groupi_n_2149);
  xnor csa_tree_add_6_33_groupi_g15684(csa_tree_add_6_33_groupi_n_2632 ,csa_tree_add_6_33_groupi_n_1186 ,csa_tree_add_6_33_groupi_n_2036);
  xnor csa_tree_add_6_33_groupi_g15685(csa_tree_add_6_33_groupi_n_2630 ,csa_tree_add_6_33_groupi_n_1090 ,csa_tree_add_6_33_groupi_n_2050);
  xnor csa_tree_add_6_33_groupi_g15686(csa_tree_add_6_33_groupi_n_2629 ,csa_tree_add_6_33_groupi_n_1246 ,csa_tree_add_6_33_groupi_n_2118);
  xnor csa_tree_add_6_33_groupi_g15687(csa_tree_add_6_33_groupi_n_2628 ,csa_tree_add_6_33_groupi_n_1511 ,csa_tree_add_6_33_groupi_n_2157);
  xnor csa_tree_add_6_33_groupi_g15688(csa_tree_add_6_33_groupi_n_2627 ,csa_tree_add_6_33_groupi_n_1395 ,csa_tree_add_6_33_groupi_n_2049);
  xnor csa_tree_add_6_33_groupi_g15689(csa_tree_add_6_33_groupi_n_2626 ,csa_tree_add_6_33_groupi_n_1077 ,csa_tree_add_6_33_groupi_n_2144);
  xnor csa_tree_add_6_33_groupi_g15690(csa_tree_add_6_33_groupi_n_2625 ,csa_tree_add_6_33_groupi_n_1215 ,csa_tree_add_6_33_groupi_n_2044);
  xnor csa_tree_add_6_33_groupi_g15691(csa_tree_add_6_33_groupi_n_2623 ,csa_tree_add_6_33_groupi_n_1385 ,csa_tree_add_6_33_groupi_n_2135);
  xnor csa_tree_add_6_33_groupi_g15692(csa_tree_add_6_33_groupi_n_2622 ,csa_tree_add_6_33_groupi_n_1514 ,csa_tree_add_6_33_groupi_n_2152);
  xnor csa_tree_add_6_33_groupi_g15693(csa_tree_add_6_33_groupi_n_2621 ,csa_tree_add_6_33_groupi_n_1219 ,csa_tree_add_6_33_groupi_n_2158);
  xnor csa_tree_add_6_33_groupi_g15694(csa_tree_add_6_33_groupi_n_2620 ,csa_tree_add_6_33_groupi_n_1327 ,csa_tree_add_6_33_groupi_n_2153);
  xnor csa_tree_add_6_33_groupi_g15695(csa_tree_add_6_33_groupi_n_2619 ,csa_tree_add_6_33_groupi_n_1522 ,csa_tree_add_6_33_groupi_n_2018);
  xnor csa_tree_add_6_33_groupi_g15696(csa_tree_add_6_33_groupi_n_2617 ,csa_tree_add_6_33_groupi_n_1240 ,csa_tree_add_6_33_groupi_n_2015);
  xnor csa_tree_add_6_33_groupi_g15697(csa_tree_add_6_33_groupi_n_2616 ,csa_tree_add_6_33_groupi_n_1456 ,csa_tree_add_6_33_groupi_n_2024);
  xnor csa_tree_add_6_33_groupi_g15698(csa_tree_add_6_33_groupi_n_2615 ,csa_tree_add_6_33_groupi_n_1379 ,csa_tree_add_6_33_groupi_n_2151);
  xnor csa_tree_add_6_33_groupi_g15699(csa_tree_add_6_33_groupi_n_2614 ,csa_tree_add_6_33_groupi_n_1582 ,csa_tree_add_6_33_groupi_n_2028);
  xnor csa_tree_add_6_33_groupi_g15700(csa_tree_add_6_33_groupi_n_2612 ,csa_tree_add_6_33_groupi_n_1389 ,csa_tree_add_6_33_groupi_n_2029);
  xnor csa_tree_add_6_33_groupi_g15701(csa_tree_add_6_33_groupi_n_2611 ,csa_tree_add_6_33_groupi_n_1572 ,csa_tree_add_6_33_groupi_n_2084);
  xnor csa_tree_add_6_33_groupi_g15702(csa_tree_add_6_33_groupi_n_2610 ,csa_tree_add_6_33_groupi_n_1231 ,csa_tree_add_6_33_groupi_n_2046);
  xnor csa_tree_add_6_33_groupi_g15703(csa_tree_add_6_33_groupi_n_2609 ,csa_tree_add_6_33_groupi_n_1392 ,csa_tree_add_6_33_groupi_n_2136);
  xnor csa_tree_add_6_33_groupi_g15704(csa_tree_add_6_33_groupi_n_2608 ,csa_tree_add_6_33_groupi_n_1201 ,csa_tree_add_6_33_groupi_n_2079);
  xnor csa_tree_add_6_33_groupi_g15705(csa_tree_add_6_33_groupi_n_2607 ,csa_tree_add_6_33_groupi_n_1571 ,csa_tree_add_6_33_groupi_n_2115);
  xnor csa_tree_add_6_33_groupi_g15706(csa_tree_add_6_33_groupi_n_2606 ,csa_tree_add_6_33_groupi_n_1111 ,csa_tree_add_6_33_groupi_n_2033);
  xnor csa_tree_add_6_33_groupi_g15707(csa_tree_add_6_33_groupi_n_2605 ,csa_tree_add_6_33_groupi_n_1291 ,csa_tree_add_6_33_groupi_n_2116);
  xnor csa_tree_add_6_33_groupi_g15708(csa_tree_add_6_33_groupi_n_2604 ,csa_tree_add_6_33_groupi_n_1188 ,csa_tree_add_6_33_groupi_n_2031);
  xnor csa_tree_add_6_33_groupi_g15709(csa_tree_add_6_33_groupi_n_2603 ,csa_tree_add_6_33_groupi_n_1182 ,csa_tree_add_6_33_groupi_n_2156);
  xnor csa_tree_add_6_33_groupi_g15710(csa_tree_add_6_33_groupi_n_2602 ,csa_tree_add_6_33_groupi_n_1549 ,csa_tree_add_6_33_groupi_n_2145);
  xnor csa_tree_add_6_33_groupi_g15711(csa_tree_add_6_33_groupi_n_2600 ,csa_tree_add_6_33_groupi_n_1435 ,csa_tree_add_6_33_groupi_n_2017);
  xnor csa_tree_add_6_33_groupi_g15712(csa_tree_add_6_33_groupi_n_2599 ,csa_tree_add_6_33_groupi_n_1118 ,csa_tree_add_6_33_groupi_n_2026);
  xnor csa_tree_add_6_33_groupi_g15713(csa_tree_add_6_33_groupi_n_2598 ,csa_tree_add_6_33_groupi_n_1383 ,csa_tree_add_6_33_groupi_n_2146);
  xnor csa_tree_add_6_33_groupi_g15714(csa_tree_add_6_33_groupi_n_2597 ,csa_tree_add_6_33_groupi_n_1536 ,csa_tree_add_6_33_groupi_n_2131);
  xnor csa_tree_add_6_33_groupi_g15715(csa_tree_add_6_33_groupi_n_2596 ,csa_tree_add_6_33_groupi_n_1474 ,csa_tree_add_6_33_groupi_n_2105);
  xnor csa_tree_add_6_33_groupi_g15716(csa_tree_add_6_33_groupi_n_2595 ,csa_tree_add_6_33_groupi_n_1445 ,csa_tree_add_6_33_groupi_n_2025);
  xnor csa_tree_add_6_33_groupi_g15717(csa_tree_add_6_33_groupi_n_2594 ,csa_tree_add_6_33_groupi_n_1609 ,csa_tree_add_6_33_groupi_n_2159);
  xnor csa_tree_add_6_33_groupi_g15718(csa_tree_add_6_33_groupi_n_2593 ,csa_tree_add_6_33_groupi_n_1559 ,csa_tree_add_6_33_groupi_n_2109);
  xnor csa_tree_add_6_33_groupi_g15719(csa_tree_add_6_33_groupi_n_2592 ,csa_tree_add_6_33_groupi_n_1564 ,csa_tree_add_6_33_groupi_n_2023);
  xnor csa_tree_add_6_33_groupi_g15720(csa_tree_add_6_33_groupi_n_2591 ,csa_tree_add_6_33_groupi_n_1256 ,csa_tree_add_6_33_groupi_n_2053);
  xnor csa_tree_add_6_33_groupi_g15721(csa_tree_add_6_33_groupi_n_2590 ,csa_tree_add_6_33_groupi_n_1555 ,csa_tree_add_6_33_groupi_n_2095);
  xnor csa_tree_add_6_33_groupi_g15722(csa_tree_add_6_33_groupi_n_2588 ,csa_tree_add_6_33_groupi_n_1220 ,csa_tree_add_6_33_groupi_n_2077);
  not csa_tree_add_6_33_groupi_g15723(csa_tree_add_6_33_groupi_n_2534 ,csa_tree_add_6_33_groupi_n_2535);
  not csa_tree_add_6_33_groupi_g15724(csa_tree_add_6_33_groupi_n_2519 ,csa_tree_add_6_33_groupi_n_2520);
  not csa_tree_add_6_33_groupi_g15725(csa_tree_add_6_33_groupi_n_2498 ,csa_tree_add_6_33_groupi_n_2499);
  or csa_tree_add_6_33_groupi_g15726(csa_tree_add_6_33_groupi_n_2493 ,csa_tree_add_6_33_groupi_n_1042 ,csa_tree_add_6_33_groupi_n_2359);
  or csa_tree_add_6_33_groupi_g15727(csa_tree_add_6_33_groupi_n_2492 ,csa_tree_add_6_33_groupi_n_1892 ,csa_tree_add_6_33_groupi_n_2357);
  or csa_tree_add_6_33_groupi_g15728(csa_tree_add_6_33_groupi_n_2491 ,csa_tree_add_6_33_groupi_n_1998 ,csa_tree_add_6_33_groupi_n_2361);
  nor csa_tree_add_6_33_groupi_g15729(csa_tree_add_6_33_groupi_n_2490 ,csa_tree_add_6_33_groupi_n_1142 ,csa_tree_add_6_33_groupi_n_2326);
  or csa_tree_add_6_33_groupi_g15730(csa_tree_add_6_33_groupi_n_2489 ,csa_tree_add_6_33_groupi_n_1899 ,csa_tree_add_6_33_groupi_n_2354);
  and csa_tree_add_6_33_groupi_g15731(csa_tree_add_6_33_groupi_n_2488 ,csa_tree_add_6_33_groupi_n_1815 ,csa_tree_add_6_33_groupi_n_2364);
  nor csa_tree_add_6_33_groupi_g15732(csa_tree_add_6_33_groupi_n_2487 ,csa_tree_add_6_33_groupi_n_1483 ,csa_tree_add_6_33_groupi_n_2351);
  or csa_tree_add_6_33_groupi_g15733(csa_tree_add_6_33_groupi_n_2486 ,csa_tree_add_6_33_groupi_n_1484 ,csa_tree_add_6_33_groupi_n_2350);
  and csa_tree_add_6_33_groupi_g15734(csa_tree_add_6_33_groupi_n_2485 ,csa_tree_add_6_33_groupi_n_1698 ,csa_tree_add_6_33_groupi_n_2362);
  and csa_tree_add_6_33_groupi_g15735(csa_tree_add_6_33_groupi_n_2582 ,csa_tree_add_6_33_groupi_n_1886 ,csa_tree_add_6_33_groupi_n_2264);
  and csa_tree_add_6_33_groupi_g15736(csa_tree_add_6_33_groupi_n_2581 ,csa_tree_add_6_33_groupi_n_1959 ,csa_tree_add_6_33_groupi_n_2304);
  and csa_tree_add_6_33_groupi_g15737(csa_tree_add_6_33_groupi_n_2580 ,csa_tree_add_6_33_groupi_n_1830 ,csa_tree_add_6_33_groupi_n_2268);
  and csa_tree_add_6_33_groupi_g15738(csa_tree_add_6_33_groupi_n_2579 ,csa_tree_add_6_33_groupi_n_1939 ,csa_tree_add_6_33_groupi_n_2296);
  and csa_tree_add_6_33_groupi_g15739(csa_tree_add_6_33_groupi_n_2578 ,csa_tree_add_6_33_groupi_n_2000 ,csa_tree_add_6_33_groupi_n_2320);
  and csa_tree_add_6_33_groupi_g15740(csa_tree_add_6_33_groupi_n_2577 ,csa_tree_add_6_33_groupi_n_1758 ,csa_tree_add_6_33_groupi_n_2216);
  and csa_tree_add_6_33_groupi_g15741(csa_tree_add_6_33_groupi_n_2576 ,csa_tree_add_6_33_groupi_n_1757 ,csa_tree_add_6_33_groupi_n_2231);
  and csa_tree_add_6_33_groupi_g15742(csa_tree_add_6_33_groupi_n_2575 ,csa_tree_add_6_33_groupi_n_1997 ,csa_tree_add_6_33_groupi_n_2322);
  and csa_tree_add_6_33_groupi_g15743(csa_tree_add_6_33_groupi_n_2574 ,csa_tree_add_6_33_groupi_n_1914 ,csa_tree_add_6_33_groupi_n_2275);
  and csa_tree_add_6_33_groupi_g15744(csa_tree_add_6_33_groupi_n_2573 ,csa_tree_add_6_33_groupi_n_1891 ,csa_tree_add_6_33_groupi_n_2305);
  and csa_tree_add_6_33_groupi_g15745(csa_tree_add_6_33_groupi_n_2572 ,csa_tree_add_6_33_groupi_n_1893 ,csa_tree_add_6_33_groupi_n_2309);
  and csa_tree_add_6_33_groupi_g15746(csa_tree_add_6_33_groupi_n_2571 ,csa_tree_add_6_33_groupi_n_1904 ,csa_tree_add_6_33_groupi_n_2281);
  and csa_tree_add_6_33_groupi_g15747(csa_tree_add_6_33_groupi_n_2570 ,csa_tree_add_6_33_groupi_n_1819 ,csa_tree_add_6_33_groupi_n_2233);
  and csa_tree_add_6_33_groupi_g15748(csa_tree_add_6_33_groupi_n_2569 ,csa_tree_add_6_33_groupi_n_1905 ,csa_tree_add_6_33_groupi_n_2180);
  and csa_tree_add_6_33_groupi_g15749(csa_tree_add_6_33_groupi_n_2568 ,csa_tree_add_6_33_groupi_n_1816 ,csa_tree_add_6_33_groupi_n_2317);
  and csa_tree_add_6_33_groupi_g15750(csa_tree_add_6_33_groupi_n_2567 ,csa_tree_add_6_33_groupi_n_1734 ,csa_tree_add_6_33_groupi_n_2280);
  and csa_tree_add_6_33_groupi_g15751(csa_tree_add_6_33_groupi_n_2566 ,csa_tree_add_6_33_groupi_n_1710 ,csa_tree_add_6_33_groupi_n_2207);
  and csa_tree_add_6_33_groupi_g15752(csa_tree_add_6_33_groupi_n_2565 ,csa_tree_add_6_33_groupi_n_1776 ,csa_tree_add_6_33_groupi_n_2278);
  and csa_tree_add_6_33_groupi_g15753(csa_tree_add_6_33_groupi_n_2564 ,csa_tree_add_6_33_groupi_n_1714 ,csa_tree_add_6_33_groupi_n_2188);
  and csa_tree_add_6_33_groupi_g15754(csa_tree_add_6_33_groupi_n_2563 ,csa_tree_add_6_33_groupi_n_1877 ,csa_tree_add_6_33_groupi_n_2263);
  and csa_tree_add_6_33_groupi_g15755(csa_tree_add_6_33_groupi_n_2562 ,csa_tree_add_6_33_groupi_n_1712 ,csa_tree_add_6_33_groupi_n_2307);
  and csa_tree_add_6_33_groupi_g15756(csa_tree_add_6_33_groupi_n_2561 ,csa_tree_add_6_33_groupi_n_1994 ,csa_tree_add_6_33_groupi_n_2323);
  and csa_tree_add_6_33_groupi_g15757(csa_tree_add_6_33_groupi_n_2560 ,csa_tree_add_6_33_groupi_n_1725 ,csa_tree_add_6_33_groupi_n_2183);
  and csa_tree_add_6_33_groupi_g15758(csa_tree_add_6_33_groupi_n_2559 ,csa_tree_add_6_33_groupi_n_1961 ,csa_tree_add_6_33_groupi_n_2215);
  and csa_tree_add_6_33_groupi_g15759(csa_tree_add_6_33_groupi_n_2558 ,csa_tree_add_6_33_groupi_n_1897 ,csa_tree_add_6_33_groupi_n_2282);
  and csa_tree_add_6_33_groupi_g15760(csa_tree_add_6_33_groupi_n_2557 ,csa_tree_add_6_33_groupi_n_1942 ,csa_tree_add_6_33_groupi_n_2254);
  and csa_tree_add_6_33_groupi_g15761(csa_tree_add_6_33_groupi_n_2556 ,csa_tree_add_6_33_groupi_n_1979 ,csa_tree_add_6_33_groupi_n_2211);
  and csa_tree_add_6_33_groupi_g15762(csa_tree_add_6_33_groupi_n_2555 ,csa_tree_add_6_33_groupi_n_1653 ,csa_tree_add_6_33_groupi_n_2291);
  and csa_tree_add_6_33_groupi_g15763(csa_tree_add_6_33_groupi_n_2554 ,csa_tree_add_6_33_groupi_n_1867 ,csa_tree_add_6_33_groupi_n_2311);
  and csa_tree_add_6_33_groupi_g15764(csa_tree_add_6_33_groupi_n_2553 ,csa_tree_add_6_33_groupi_n_1984 ,csa_tree_add_6_33_groupi_n_2298);
  and csa_tree_add_6_33_groupi_g15765(csa_tree_add_6_33_groupi_n_2552 ,csa_tree_add_6_33_groupi_n_1847 ,csa_tree_add_6_33_groupi_n_2277);
  and csa_tree_add_6_33_groupi_g15766(csa_tree_add_6_33_groupi_n_2551 ,csa_tree_add_6_33_groupi_n_1820 ,csa_tree_add_6_33_groupi_n_2259);
  and csa_tree_add_6_33_groupi_g15767(csa_tree_add_6_33_groupi_n_2550 ,csa_tree_add_6_33_groupi_n_1996 ,csa_tree_add_6_33_groupi_n_2255);
  and csa_tree_add_6_33_groupi_g15768(csa_tree_add_6_33_groupi_n_2549 ,csa_tree_add_6_33_groupi_n_1835 ,csa_tree_add_6_33_groupi_n_2314);
  and csa_tree_add_6_33_groupi_g15769(csa_tree_add_6_33_groupi_n_2548 ,csa_tree_add_6_33_groupi_n_1752 ,csa_tree_add_6_33_groupi_n_2226);
  and csa_tree_add_6_33_groupi_g15770(csa_tree_add_6_33_groupi_n_2547 ,csa_tree_add_6_33_groupi_n_1839 ,csa_tree_add_6_33_groupi_n_2252);
  and csa_tree_add_6_33_groupi_g15771(csa_tree_add_6_33_groupi_n_2546 ,csa_tree_add_6_33_groupi_n_1976 ,csa_tree_add_6_33_groupi_n_2181);
  and csa_tree_add_6_33_groupi_g15772(csa_tree_add_6_33_groupi_n_2545 ,csa_tree_add_6_33_groupi_n_1863 ,csa_tree_add_6_33_groupi_n_2240);
  and csa_tree_add_6_33_groupi_g15773(csa_tree_add_6_33_groupi_n_2544 ,csa_tree_add_6_33_groupi_n_1846 ,csa_tree_add_6_33_groupi_n_2256);
  and csa_tree_add_6_33_groupi_g15774(csa_tree_add_6_33_groupi_n_2543 ,csa_tree_add_6_33_groupi_n_1844 ,csa_tree_add_6_33_groupi_n_2234);
  and csa_tree_add_6_33_groupi_g15775(csa_tree_add_6_33_groupi_n_2542 ,csa_tree_add_6_33_groupi_n_1958 ,csa_tree_add_6_33_groupi_n_2312);
  and csa_tree_add_6_33_groupi_g15776(csa_tree_add_6_33_groupi_n_2541 ,csa_tree_add_6_33_groupi_n_1990 ,csa_tree_add_6_33_groupi_n_2247);
  and csa_tree_add_6_33_groupi_g15777(csa_tree_add_6_33_groupi_n_2540 ,csa_tree_add_6_33_groupi_n_1729 ,csa_tree_add_6_33_groupi_n_2243);
  and csa_tree_add_6_33_groupi_g15778(csa_tree_add_6_33_groupi_n_2539 ,csa_tree_add_6_33_groupi_n_1925 ,csa_tree_add_6_33_groupi_n_2184);
  and csa_tree_add_6_33_groupi_g15779(csa_tree_add_6_33_groupi_n_2538 ,csa_tree_add_6_33_groupi_n_1806 ,csa_tree_add_6_33_groupi_n_2230);
  and csa_tree_add_6_33_groupi_g15780(csa_tree_add_6_33_groupi_n_2537 ,csa_tree_add_6_33_groupi_n_1802 ,csa_tree_add_6_33_groupi_n_2227);
  and csa_tree_add_6_33_groupi_g15781(csa_tree_add_6_33_groupi_n_2536 ,csa_tree_add_6_33_groupi_n_1874 ,csa_tree_add_6_33_groupi_n_2272);
  and csa_tree_add_6_33_groupi_g15782(csa_tree_add_6_33_groupi_n_2535 ,csa_tree_add_6_33_groupi_n_1779 ,csa_tree_add_6_33_groupi_n_2271);
  and csa_tree_add_6_33_groupi_g15783(csa_tree_add_6_33_groupi_n_2533 ,csa_tree_add_6_33_groupi_n_1706 ,csa_tree_add_6_33_groupi_n_2191);
  and csa_tree_add_6_33_groupi_g15784(csa_tree_add_6_33_groupi_n_2532 ,csa_tree_add_6_33_groupi_n_1668 ,csa_tree_add_6_33_groupi_n_2290);
  and csa_tree_add_6_33_groupi_g15785(csa_tree_add_6_33_groupi_n_2531 ,csa_tree_add_6_33_groupi_n_1879 ,csa_tree_add_6_33_groupi_n_2313);
  and csa_tree_add_6_33_groupi_g15786(csa_tree_add_6_33_groupi_n_2530 ,csa_tree_add_6_33_groupi_n_1722 ,csa_tree_add_6_33_groupi_n_2212);
  and csa_tree_add_6_33_groupi_g15787(csa_tree_add_6_33_groupi_n_2529 ,csa_tree_add_6_33_groupi_n_1745 ,csa_tree_add_6_33_groupi_n_2262);
  and csa_tree_add_6_33_groupi_g15788(csa_tree_add_6_33_groupi_n_2528 ,csa_tree_add_6_33_groupi_n_1671 ,csa_tree_add_6_33_groupi_n_2266);
  and csa_tree_add_6_33_groupi_g15789(csa_tree_add_6_33_groupi_n_2527 ,csa_tree_add_6_33_groupi_n_1765 ,csa_tree_add_6_33_groupi_n_2316);
  and csa_tree_add_6_33_groupi_g15790(csa_tree_add_6_33_groupi_n_2526 ,csa_tree_add_6_33_groupi_n_1657 ,csa_tree_add_6_33_groupi_n_2287);
  and csa_tree_add_6_33_groupi_g15791(csa_tree_add_6_33_groupi_n_2525 ,csa_tree_add_6_33_groupi_n_1724 ,csa_tree_add_6_33_groupi_n_2193);
  and csa_tree_add_6_33_groupi_g15792(csa_tree_add_6_33_groupi_n_2524 ,csa_tree_add_6_33_groupi_n_1965 ,csa_tree_add_6_33_groupi_n_2306);
  and csa_tree_add_6_33_groupi_g15793(csa_tree_add_6_33_groupi_n_2523 ,csa_tree_add_6_33_groupi_n_1917 ,csa_tree_add_6_33_groupi_n_2269);
  and csa_tree_add_6_33_groupi_g15794(csa_tree_add_6_33_groupi_n_2522 ,csa_tree_add_6_33_groupi_n_1822 ,csa_tree_add_6_33_groupi_n_2253);
  and csa_tree_add_6_33_groupi_g15795(csa_tree_add_6_33_groupi_n_2521 ,csa_tree_add_6_33_groupi_n_1995 ,csa_tree_add_6_33_groupi_n_2289);
  and csa_tree_add_6_33_groupi_g15796(csa_tree_add_6_33_groupi_n_2520 ,csa_tree_add_6_33_groupi_n_1968 ,csa_tree_add_6_33_groupi_n_2270);
  and csa_tree_add_6_33_groupi_g15797(csa_tree_add_6_33_groupi_n_2518 ,csa_tree_add_6_33_groupi_n_1894 ,csa_tree_add_6_33_groupi_n_2285);
  and csa_tree_add_6_33_groupi_g15798(csa_tree_add_6_33_groupi_n_2517 ,csa_tree_add_6_33_groupi_n_1922 ,csa_tree_add_6_33_groupi_n_2199);
  and csa_tree_add_6_33_groupi_g15799(csa_tree_add_6_33_groupi_n_2516 ,csa_tree_add_6_33_groupi_n_1661 ,csa_tree_add_6_33_groupi_n_2208);
  and csa_tree_add_6_33_groupi_g15800(csa_tree_add_6_33_groupi_n_2515 ,csa_tree_add_6_33_groupi_n_1687 ,csa_tree_add_6_33_groupi_n_2189);
  and csa_tree_add_6_33_groupi_g15801(csa_tree_add_6_33_groupi_n_2514 ,csa_tree_add_6_33_groupi_n_1973 ,csa_tree_add_6_33_groupi_n_2232);
  and csa_tree_add_6_33_groupi_g15802(csa_tree_add_6_33_groupi_n_2513 ,csa_tree_add_6_33_groupi_n_1872 ,csa_tree_add_6_33_groupi_n_2288);
  and csa_tree_add_6_33_groupi_g15803(csa_tree_add_6_33_groupi_n_2512 ,csa_tree_add_6_33_groupi_n_1826 ,csa_tree_add_6_33_groupi_n_2242);
  and csa_tree_add_6_33_groupi_g15804(csa_tree_add_6_33_groupi_n_2511 ,csa_tree_add_6_33_groupi_n_1828 ,csa_tree_add_6_33_groupi_n_2274);
  and csa_tree_add_6_33_groupi_g15805(csa_tree_add_6_33_groupi_n_2510 ,csa_tree_add_6_33_groupi_n_1682 ,csa_tree_add_6_33_groupi_n_2318);
  and csa_tree_add_6_33_groupi_g15806(csa_tree_add_6_33_groupi_n_2509 ,csa_tree_add_6_33_groupi_n_1967 ,csa_tree_add_6_33_groupi_n_2238);
  and csa_tree_add_6_33_groupi_g15807(csa_tree_add_6_33_groupi_n_2508 ,csa_tree_add_6_33_groupi_n_1873 ,csa_tree_add_6_33_groupi_n_2300);
  and csa_tree_add_6_33_groupi_g15808(csa_tree_add_6_33_groupi_n_2507 ,csa_tree_add_6_33_groupi_n_1980 ,csa_tree_add_6_33_groupi_n_2245);
  and csa_tree_add_6_33_groupi_g15809(csa_tree_add_6_33_groupi_n_2506 ,csa_tree_add_6_33_groupi_n_1699 ,csa_tree_add_6_33_groupi_n_2246);
  and csa_tree_add_6_33_groupi_g15810(csa_tree_add_6_33_groupi_n_2505 ,csa_tree_add_6_33_groupi_n_1992 ,csa_tree_add_6_33_groupi_n_2210);
  and csa_tree_add_6_33_groupi_g15811(csa_tree_add_6_33_groupi_n_2504 ,csa_tree_add_6_33_groupi_n_1907 ,csa_tree_add_6_33_groupi_n_2236);
  and csa_tree_add_6_33_groupi_g15812(csa_tree_add_6_33_groupi_n_2503 ,csa_tree_add_6_33_groupi_n_1829 ,csa_tree_add_6_33_groupi_n_2257);
  and csa_tree_add_6_33_groupi_g15813(csa_tree_add_6_33_groupi_n_2502 ,csa_tree_add_6_33_groupi_n_1703 ,csa_tree_add_6_33_groupi_n_2220);
  and csa_tree_add_6_33_groupi_g15814(csa_tree_add_6_33_groupi_n_2501 ,csa_tree_add_6_33_groupi_n_1842 ,csa_tree_add_6_33_groupi_n_2284);
  and csa_tree_add_6_33_groupi_g15815(csa_tree_add_6_33_groupi_n_2500 ,csa_tree_add_6_33_groupi_n_1809 ,csa_tree_add_6_33_groupi_n_2301);
  and csa_tree_add_6_33_groupi_g15816(csa_tree_add_6_33_groupi_n_2499 ,csa_tree_add_6_33_groupi_n_1705 ,csa_tree_add_6_33_groupi_n_2265);
  and csa_tree_add_6_33_groupi_g15817(csa_tree_add_6_33_groupi_n_2497 ,csa_tree_add_6_33_groupi_n_1730 ,csa_tree_add_6_33_groupi_n_2308);
  and csa_tree_add_6_33_groupi_g15818(csa_tree_add_6_33_groupi_n_2496 ,csa_tree_add_6_33_groupi_n_1852 ,csa_tree_add_6_33_groupi_n_2194);
  and csa_tree_add_6_33_groupi_g15819(csa_tree_add_6_33_groupi_n_2495 ,csa_tree_add_6_33_groupi_n_1754 ,csa_tree_add_6_33_groupi_n_2229);
  and csa_tree_add_6_33_groupi_g15820(csa_tree_add_6_33_groupi_n_2494 ,csa_tree_add_6_33_groupi_n_1697 ,csa_tree_add_6_33_groupi_n_2249);
  not csa_tree_add_6_33_groupi_g15821(csa_tree_add_6_33_groupi_n_2469 ,csa_tree_add_6_33_groupi_n_2468);
  not csa_tree_add_6_33_groupi_g15822(csa_tree_add_6_33_groupi_n_2467 ,csa_tree_add_6_33_groupi_n_2466);
  not csa_tree_add_6_33_groupi_g15823(csa_tree_add_6_33_groupi_n_2445 ,csa_tree_add_6_33_groupi_n_2446);
  not csa_tree_add_6_33_groupi_g15824(csa_tree_add_6_33_groupi_n_2442 ,csa_tree_add_6_33_groupi_n_2443);
  not csa_tree_add_6_33_groupi_g15825(csa_tree_add_6_33_groupi_n_2433 ,csa_tree_add_6_33_groupi_n_2434);
  not csa_tree_add_6_33_groupi_g15826(csa_tree_add_6_33_groupi_n_2425 ,csa_tree_add_6_33_groupi_n_2426);
  not csa_tree_add_6_33_groupi_g15827(csa_tree_add_6_33_groupi_n_2421 ,csa_tree_add_6_33_groupi_n_2420);
  not csa_tree_add_6_33_groupi_g15828(csa_tree_add_6_33_groupi_n_2417 ,csa_tree_add_6_33_groupi_n_2418);
  not csa_tree_add_6_33_groupi_g15829(csa_tree_add_6_33_groupi_n_2414 ,csa_tree_add_6_33_groupi_n_2415);
  not csa_tree_add_6_33_groupi_g15830(csa_tree_add_6_33_groupi_n_2412 ,csa_tree_add_6_33_groupi_n_2413);
  not csa_tree_add_6_33_groupi_g15831(csa_tree_add_6_33_groupi_n_2410 ,csa_tree_add_6_33_groupi_n_2411);
  not csa_tree_add_6_33_groupi_g15832(csa_tree_add_6_33_groupi_n_2409 ,csa_tree_add_6_33_groupi_n_2408);
  not csa_tree_add_6_33_groupi_g15833(csa_tree_add_6_33_groupi_n_2405 ,csa_tree_add_6_33_groupi_n_2406);
  not csa_tree_add_6_33_groupi_g15834(csa_tree_add_6_33_groupi_n_2400 ,csa_tree_add_6_33_groupi_n_2401);
  not csa_tree_add_6_33_groupi_g15835(csa_tree_add_6_33_groupi_n_2397 ,csa_tree_add_6_33_groupi_n_2398);
  not csa_tree_add_6_33_groupi_g15836(csa_tree_add_6_33_groupi_n_2394 ,csa_tree_add_6_33_groupi_n_2395);
  not csa_tree_add_6_33_groupi_g15837(csa_tree_add_6_33_groupi_n_2390 ,csa_tree_add_6_33_groupi_n_2391);
  not csa_tree_add_6_33_groupi_g15838(csa_tree_add_6_33_groupi_n_2388 ,csa_tree_add_6_33_groupi_n_2389);
  not csa_tree_add_6_33_groupi_g15839(csa_tree_add_6_33_groupi_n_2382 ,csa_tree_add_6_33_groupi_n_2383);
  not csa_tree_add_6_33_groupi_g15840(csa_tree_add_6_33_groupi_n_2377 ,csa_tree_add_6_33_groupi_n_2378);
  xnor csa_tree_add_6_33_groupi_g15841(out1[0] ,csa_tree_add_6_33_groupi_n_1649 ,in3[0]);
  and csa_tree_add_6_33_groupi_g15842(csa_tree_add_6_33_groupi_n_2374 ,csa_tree_add_6_33_groupi_n_1790 ,csa_tree_add_6_33_groupi_n_2367);
  nor csa_tree_add_6_33_groupi_g15843(csa_tree_add_6_33_groupi_n_2373 ,csa_tree_add_6_33_groupi_n_1409 ,csa_tree_add_6_33_groupi_n_2329);
  or csa_tree_add_6_33_groupi_g15844(csa_tree_add_6_33_groupi_n_2372 ,csa_tree_add_6_33_groupi_n_1410 ,csa_tree_add_6_33_groupi_n_2328);
  or csa_tree_add_6_33_groupi_g15845(csa_tree_add_6_33_groupi_n_2371 ,csa_tree_add_6_33_groupi_n_1143 ,csa_tree_add_6_33_groupi_n_2325);
  or csa_tree_add_6_33_groupi_g15846(csa_tree_add_6_33_groupi_n_2370 ,csa_tree_add_6_33_groupi_n_1728 ,csa_tree_add_6_33_groupi_n_2369);
  and csa_tree_add_6_33_groupi_g15847(csa_tree_add_6_33_groupi_n_2484 ,csa_tree_add_6_33_groupi_n_1688 ,csa_tree_add_6_33_groupi_n_2222);
  and csa_tree_add_6_33_groupi_g15848(csa_tree_add_6_33_groupi_n_2483 ,csa_tree_add_6_33_groupi_n_1916 ,csa_tree_add_6_33_groupi_n_2295);
  and csa_tree_add_6_33_groupi_g15849(csa_tree_add_6_33_groupi_n_2482 ,csa_tree_add_6_33_groupi_n_1774 ,csa_tree_add_6_33_groupi_n_2319);
  and csa_tree_add_6_33_groupi_g15850(csa_tree_add_6_33_groupi_n_2481 ,csa_tree_add_6_33_groupi_n_1787 ,csa_tree_add_6_33_groupi_n_2261);
  xnor csa_tree_add_6_33_groupi_g15851(csa_tree_add_6_33_groupi_n_2480 ,csa_tree_add_6_33_groupi_n_1593 ,csa_tree_add_6_33_groupi_n_1639);
  and csa_tree_add_6_33_groupi_g15852(csa_tree_add_6_33_groupi_n_2479 ,csa_tree_add_6_33_groupi_n_1677 ,csa_tree_add_6_33_groupi_n_2321);
  and csa_tree_add_6_33_groupi_g15853(csa_tree_add_6_33_groupi_n_2478 ,csa_tree_add_6_33_groupi_n_1937 ,csa_tree_add_6_33_groupi_n_2294);
  and csa_tree_add_6_33_groupi_g15854(csa_tree_add_6_33_groupi_n_2477 ,csa_tree_add_6_33_groupi_n_1986 ,csa_tree_add_6_33_groupi_n_2217);
  and csa_tree_add_6_33_groupi_g15855(csa_tree_add_6_33_groupi_n_2476 ,csa_tree_add_6_33_groupi_n_1972 ,csa_tree_add_6_33_groupi_n_2303);
  and csa_tree_add_6_33_groupi_g15856(csa_tree_add_6_33_groupi_n_2475 ,csa_tree_add_6_33_groupi_n_1890 ,csa_tree_add_6_33_groupi_n_2293);
  and csa_tree_add_6_33_groupi_g15857(csa_tree_add_6_33_groupi_n_2474 ,csa_tree_add_6_33_groupi_n_1966 ,csa_tree_add_6_33_groupi_n_2292);
  and csa_tree_add_6_33_groupi_g15858(csa_tree_add_6_33_groupi_n_2473 ,csa_tree_add_6_33_groupi_n_1900 ,csa_tree_add_6_33_groupi_n_2195);
  and csa_tree_add_6_33_groupi_g15859(csa_tree_add_6_33_groupi_n_2472 ,csa_tree_add_6_33_groupi_n_1719 ,csa_tree_add_6_33_groupi_n_2228);
  and csa_tree_add_6_33_groupi_g15860(csa_tree_add_6_33_groupi_n_2471 ,csa_tree_add_6_33_groupi_n_1853 ,csa_tree_add_6_33_groupi_n_2286);
  and csa_tree_add_6_33_groupi_g15861(csa_tree_add_6_33_groupi_n_2470 ,csa_tree_add_6_33_groupi_n_1834 ,csa_tree_add_6_33_groupi_n_2235);
  xnor csa_tree_add_6_33_groupi_g15862(csa_tree_add_6_33_groupi_n_2468 ,csa_tree_add_6_33_groupi_n_1646 ,in1[11]);
  xnor csa_tree_add_6_33_groupi_g15863(csa_tree_add_6_33_groupi_n_2466 ,csa_tree_add_6_33_groupi_n_1634 ,in1[14]);
  and csa_tree_add_6_33_groupi_g15864(csa_tree_add_6_33_groupi_n_2465 ,csa_tree_add_6_33_groupi_n_1732 ,csa_tree_add_6_33_groupi_n_2203);
  and csa_tree_add_6_33_groupi_g15865(csa_tree_add_6_33_groupi_n_2464 ,csa_tree_add_6_33_groupi_n_1726 ,csa_tree_add_6_33_groupi_n_2315);
  and csa_tree_add_6_33_groupi_g15866(csa_tree_add_6_33_groupi_n_2463 ,csa_tree_add_6_33_groupi_n_1859 ,csa_tree_add_6_33_groupi_n_2273);
  and csa_tree_add_6_33_groupi_g15867(csa_tree_add_6_33_groupi_n_2462 ,csa_tree_add_6_33_groupi_n_1709 ,csa_tree_add_6_33_groupi_n_2201);
  and csa_tree_add_6_33_groupi_g15868(csa_tree_add_6_33_groupi_n_2461 ,csa_tree_add_6_33_groupi_n_1662 ,csa_tree_add_6_33_groupi_n_2196);
  and csa_tree_add_6_33_groupi_g15869(csa_tree_add_6_33_groupi_n_2460 ,csa_tree_add_6_33_groupi_n_1783 ,csa_tree_add_6_33_groupi_n_2258);
  and csa_tree_add_6_33_groupi_g15870(csa_tree_add_6_33_groupi_n_2459 ,csa_tree_add_6_33_groupi_n_1906 ,csa_tree_add_6_33_groupi_n_2250);
  and csa_tree_add_6_33_groupi_g15871(csa_tree_add_6_33_groupi_n_2458 ,csa_tree_add_6_33_groupi_n_1731 ,csa_tree_add_6_33_groupi_n_2237);
  xnor csa_tree_add_6_33_groupi_g15872(csa_tree_add_6_33_groupi_n_2457 ,csa_tree_add_6_33_groupi_n_1638 ,in1[2]);
  and csa_tree_add_6_33_groupi_g15873(csa_tree_add_6_33_groupi_n_2456 ,csa_tree_add_6_33_groupi_n_1928 ,csa_tree_add_6_33_groupi_n_2185);
  and csa_tree_add_6_33_groupi_g15874(csa_tree_add_6_33_groupi_n_2455 ,csa_tree_add_6_33_groupi_n_1936 ,csa_tree_add_6_33_groupi_n_2279);
  and csa_tree_add_6_33_groupi_g15875(csa_tree_add_6_33_groupi_n_2454 ,csa_tree_add_6_33_groupi_n_1702 ,csa_tree_add_6_33_groupi_n_2186);
  and csa_tree_add_6_33_groupi_g15876(csa_tree_add_6_33_groupi_n_2453 ,csa_tree_add_6_33_groupi_n_1938 ,csa_tree_add_6_33_groupi_n_2198);
  and csa_tree_add_6_33_groupi_g15877(csa_tree_add_6_33_groupi_n_2452 ,csa_tree_add_6_33_groupi_n_1796 ,csa_tree_add_6_33_groupi_n_2244);
  and csa_tree_add_6_33_groupi_g15878(csa_tree_add_6_33_groupi_n_2451 ,csa_tree_add_6_33_groupi_n_1870 ,csa_tree_add_6_33_groupi_n_2204);
  and csa_tree_add_6_33_groupi_g15879(csa_tree_add_6_33_groupi_n_2450 ,csa_tree_add_6_33_groupi_n_1908 ,csa_tree_add_6_33_groupi_n_2187);
  and csa_tree_add_6_33_groupi_g15880(csa_tree_add_6_33_groupi_n_2449 ,csa_tree_add_6_33_groupi_n_1824 ,csa_tree_add_6_33_groupi_n_2283);
  and csa_tree_add_6_33_groupi_g15881(csa_tree_add_6_33_groupi_n_2448 ,csa_tree_add_6_33_groupi_n_1673 ,csa_tree_add_6_33_groupi_n_2190);
  and csa_tree_add_6_33_groupi_g15882(csa_tree_add_6_33_groupi_n_2447 ,csa_tree_add_6_33_groupi_n_1670 ,csa_tree_add_6_33_groupi_n_2248);
  and csa_tree_add_6_33_groupi_g15883(csa_tree_add_6_33_groupi_n_2446 ,csa_tree_add_6_33_groupi_n_1849 ,csa_tree_add_6_33_groupi_n_2192);
  and csa_tree_add_6_33_groupi_g15884(csa_tree_add_6_33_groupi_n_2444 ,csa_tree_add_6_33_groupi_n_1742 ,csa_tree_add_6_33_groupi_n_2202);
  and csa_tree_add_6_33_groupi_g15885(csa_tree_add_6_33_groupi_n_2443 ,csa_tree_add_6_33_groupi_n_1683 ,csa_tree_add_6_33_groupi_n_2251);
  and csa_tree_add_6_33_groupi_g15886(csa_tree_add_6_33_groupi_n_2441 ,csa_tree_add_6_33_groupi_n_1744 ,csa_tree_add_6_33_groupi_n_2197);
  and csa_tree_add_6_33_groupi_g15887(csa_tree_add_6_33_groupi_n_2440 ,csa_tree_add_6_33_groupi_n_1656 ,csa_tree_add_6_33_groupi_n_2205);
  and csa_tree_add_6_33_groupi_g15888(csa_tree_add_6_33_groupi_n_2439 ,csa_tree_add_6_33_groupi_n_1993 ,csa_tree_add_6_33_groupi_n_2267);
  and csa_tree_add_6_33_groupi_g15889(csa_tree_add_6_33_groupi_n_2438 ,csa_tree_add_6_33_groupi_n_1930 ,csa_tree_add_6_33_groupi_n_2302);
  and csa_tree_add_6_33_groupi_g15890(csa_tree_add_6_33_groupi_n_2437 ,csa_tree_add_6_33_groupi_n_1767 ,csa_tree_add_6_33_groupi_n_2297);
  and csa_tree_add_6_33_groupi_g15891(csa_tree_add_6_33_groupi_n_2436 ,csa_tree_add_6_33_groupi_n_1768 ,csa_tree_add_6_33_groupi_n_2310);
  and csa_tree_add_6_33_groupi_g15892(csa_tree_add_6_33_groupi_n_2435 ,csa_tree_add_6_33_groupi_n_1686 ,csa_tree_add_6_33_groupi_n_2276);
  and csa_tree_add_6_33_groupi_g15893(csa_tree_add_6_33_groupi_n_2434 ,csa_tree_add_6_33_groupi_n_1956 ,csa_tree_add_6_33_groupi_n_2213);
  and csa_tree_add_6_33_groupi_g15894(csa_tree_add_6_33_groupi_n_2432 ,csa_tree_add_6_33_groupi_n_1770 ,csa_tree_add_6_33_groupi_n_2214);
  and csa_tree_add_6_33_groupi_g15895(csa_tree_add_6_33_groupi_n_2431 ,csa_tree_add_6_33_groupi_n_1962 ,csa_tree_add_6_33_groupi_n_2299);
  and csa_tree_add_6_33_groupi_g15896(csa_tree_add_6_33_groupi_n_2430 ,csa_tree_add_6_33_groupi_n_1761 ,csa_tree_add_6_33_groupi_n_2239);
  and csa_tree_add_6_33_groupi_g15897(csa_tree_add_6_33_groupi_n_2429 ,csa_tree_add_6_33_groupi_n_1896 ,csa_tree_add_6_33_groupi_n_2218);
  and csa_tree_add_6_33_groupi_g15898(csa_tree_add_6_33_groupi_n_2428 ,csa_tree_add_6_33_groupi_n_1694 ,csa_tree_add_6_33_groupi_n_2200);
  and csa_tree_add_6_33_groupi_g15899(csa_tree_add_6_33_groupi_n_2427 ,csa_tree_add_6_33_groupi_n_1667 ,csa_tree_add_6_33_groupi_n_2182);
  and csa_tree_add_6_33_groupi_g15900(csa_tree_add_6_33_groupi_n_2426 ,csa_tree_add_6_33_groupi_n_1887 ,csa_tree_add_6_33_groupi_n_2219);
  and csa_tree_add_6_33_groupi_g15901(csa_tree_add_6_33_groupi_n_2424 ,csa_tree_add_6_33_groupi_n_1695 ,csa_tree_add_6_33_groupi_n_2260);
  and csa_tree_add_6_33_groupi_g15902(csa_tree_add_6_33_groupi_n_2423 ,csa_tree_add_6_33_groupi_n_1733 ,csa_tree_add_6_33_groupi_n_2206);
  and csa_tree_add_6_33_groupi_g15903(csa_tree_add_6_33_groupi_n_2422 ,csa_tree_add_6_33_groupi_n_1785 ,csa_tree_add_6_33_groupi_n_2324);
  xnor csa_tree_add_6_33_groupi_g15904(csa_tree_add_6_33_groupi_n_2420 ,csa_tree_add_6_33_groupi_n_1641 ,in1[9]);
  xnor csa_tree_add_6_33_groupi_g15905(csa_tree_add_6_33_groupi_n_2419 ,csa_tree_add_6_33_groupi_n_1645 ,in1[6]);
  xnor csa_tree_add_6_33_groupi_g15906(csa_tree_add_6_33_groupi_n_2418 ,csa_tree_add_6_33_groupi_n_1640 ,in1[8]);
  xnor csa_tree_add_6_33_groupi_g15907(csa_tree_add_6_33_groupi_n_2416 ,csa_tree_add_6_33_groupi_n_1624 ,in1[15]);
  xnor csa_tree_add_6_33_groupi_g15908(csa_tree_add_6_33_groupi_n_2415 ,csa_tree_add_6_33_groupi_n_1636 ,in1[7]);
  xnor csa_tree_add_6_33_groupi_g15909(csa_tree_add_6_33_groupi_n_2413 ,csa_tree_add_6_33_groupi_n_1648 ,in1[5]);
  xnor csa_tree_add_6_33_groupi_g15910(csa_tree_add_6_33_groupi_n_2411 ,csa_tree_add_6_33_groupi_n_1644 ,in1[4]);
  xnor csa_tree_add_6_33_groupi_g15911(csa_tree_add_6_33_groupi_n_2408 ,csa_tree_add_6_33_groupi_n_1635 ,in1[3]);
  and csa_tree_add_6_33_groupi_g15912(csa_tree_add_6_33_groupi_n_2407 ,csa_tree_add_6_33_groupi_n_1781 ,csa_tree_add_6_33_groupi_n_2221);
  xnor csa_tree_add_6_33_groupi_g15913(csa_tree_add_6_33_groupi_n_2406 ,csa_tree_add_6_33_groupi_n_1650 ,in2[2]);
  and csa_tree_add_6_33_groupi_g15914(csa_tree_add_6_33_groupi_n_2404 ,csa_tree_add_6_33_groupi_n_1792 ,csa_tree_add_6_33_groupi_n_2241);
  and csa_tree_add_6_33_groupi_g15915(csa_tree_add_6_33_groupi_n_2403 ,csa_tree_add_6_33_groupi_n_1860 ,csa_tree_add_6_33_groupi_n_2224);
  xnor csa_tree_add_6_33_groupi_g15916(csa_tree_add_6_33_groupi_n_2402 ,csa_tree_add_6_33_groupi_n_1627 ,in1[13]);
  xnor csa_tree_add_6_33_groupi_g15917(csa_tree_add_6_33_groupi_n_2401 ,csa_tree_add_6_33_groupi_n_1626 ,in1[12]);
  and csa_tree_add_6_33_groupi_g15918(csa_tree_add_6_33_groupi_n_2399 ,csa_tree_add_6_33_groupi_n_1793 ,csa_tree_add_6_33_groupi_n_2225);
  xnor csa_tree_add_6_33_groupi_g15919(csa_tree_add_6_33_groupi_n_2398 ,csa_tree_add_6_33_groupi_n_1628 ,in1[10]);
  xnor csa_tree_add_6_33_groupi_g15920(csa_tree_add_6_33_groupi_n_2396 ,csa_tree_add_6_33_groupi_n_1581 ,csa_tree_add_6_33_groupi_n_1629);
  xnor csa_tree_add_6_33_groupi_g15921(csa_tree_add_6_33_groupi_n_2395 ,csa_tree_add_6_33_groupi_n_1570 ,csa_tree_add_6_33_groupi_n_1642);
  and csa_tree_add_6_33_groupi_g15922(csa_tree_add_6_33_groupi_n_2393 ,csa_tree_add_6_33_groupi_n_1794 ,csa_tree_add_6_33_groupi_n_2223);
  xnor csa_tree_add_6_33_groupi_g15923(csa_tree_add_6_33_groupi_n_2392 ,csa_tree_add_6_33_groupi_n_1316 ,csa_tree_add_6_33_groupi_n_1631);
  xnor csa_tree_add_6_33_groupi_g15924(csa_tree_add_6_33_groupi_n_2391 ,csa_tree_add_6_33_groupi_n_1600 ,csa_tree_add_6_33_groupi_n_1633);
  xnor csa_tree_add_6_33_groupi_g15925(csa_tree_add_6_33_groupi_n_2389 ,csa_tree_add_6_33_groupi_n_1569 ,csa_tree_add_6_33_groupi_n_1620);
  xnor csa_tree_add_6_33_groupi_g15926(csa_tree_add_6_33_groupi_n_2387 ,csa_tree_add_6_33_groupi_n_1251 ,csa_tree_add_6_33_groupi_n_1622);
  xnor csa_tree_add_6_33_groupi_g15927(csa_tree_add_6_33_groupi_n_2386 ,csa_tree_add_6_33_groupi_n_1563 ,csa_tree_add_6_33_groupi_n_1643);
  xnor csa_tree_add_6_33_groupi_g15928(csa_tree_add_6_33_groupi_n_2385 ,csa_tree_add_6_33_groupi_n_1295 ,csa_tree_add_6_33_groupi_n_1621);
  xnor csa_tree_add_6_33_groupi_g15929(csa_tree_add_6_33_groupi_n_2384 ,csa_tree_add_6_33_groupi_n_1558 ,csa_tree_add_6_33_groupi_n_1647);
  xnor csa_tree_add_6_33_groupi_g15930(csa_tree_add_6_33_groupi_n_2383 ,csa_tree_add_6_33_groupi_n_1543 ,csa_tree_add_6_33_groupi_n_1637);
  xnor csa_tree_add_6_33_groupi_g15931(csa_tree_add_6_33_groupi_n_2381 ,csa_tree_add_6_33_groupi_n_1281 ,csa_tree_add_6_33_groupi_n_1619);
  xnor csa_tree_add_6_33_groupi_g15932(csa_tree_add_6_33_groupi_n_2380 ,csa_tree_add_6_33_groupi_n_1561 ,csa_tree_add_6_33_groupi_n_1632);
  xnor csa_tree_add_6_33_groupi_g15933(csa_tree_add_6_33_groupi_n_2379 ,csa_tree_add_6_33_groupi_n_1262 ,csa_tree_add_6_33_groupi_n_1630);
  xnor csa_tree_add_6_33_groupi_g15934(csa_tree_add_6_33_groupi_n_2378 ,csa_tree_add_6_33_groupi_n_1566 ,csa_tree_add_6_33_groupi_n_1623);
  and csa_tree_add_6_33_groupi_g15935(csa_tree_add_6_33_groupi_n_2376 ,csa_tree_add_6_33_groupi_n_1927 ,csa_tree_add_6_33_groupi_n_2209);
  not csa_tree_add_6_33_groupi_g15936(csa_tree_add_6_33_groupi_n_2369 ,csa_tree_add_6_33_groupi_n_2368);
  not csa_tree_add_6_33_groupi_g15937(csa_tree_add_6_33_groupi_n_2361 ,csa_tree_add_6_33_groupi_n_2360);
  not csa_tree_add_6_33_groupi_g15938(csa_tree_add_6_33_groupi_n_2359 ,csa_tree_add_6_33_groupi_n_2358);
  not csa_tree_add_6_33_groupi_g15939(csa_tree_add_6_33_groupi_n_2356 ,csa_tree_add_6_33_groupi_n_2355);
  not csa_tree_add_6_33_groupi_g15940(csa_tree_add_6_33_groupi_n_2354 ,csa_tree_add_6_33_groupi_n_2353);
  not csa_tree_add_6_33_groupi_g15941(csa_tree_add_6_33_groupi_n_2350 ,csa_tree_add_6_33_groupi_n_2351);
  not csa_tree_add_6_33_groupi_g15942(csa_tree_add_6_33_groupi_n_2347 ,csa_tree_add_6_33_groupi_n_2348);
  not csa_tree_add_6_33_groupi_g15943(csa_tree_add_6_33_groupi_n_2345 ,csa_tree_add_6_33_groupi_n_2346);
  not csa_tree_add_6_33_groupi_g15944(csa_tree_add_6_33_groupi_n_2343 ,csa_tree_add_6_33_groupi_n_2344);
  not csa_tree_add_6_33_groupi_g15945(csa_tree_add_6_33_groupi_n_2341 ,csa_tree_add_6_33_groupi_n_2342);
  not csa_tree_add_6_33_groupi_g15946(csa_tree_add_6_33_groupi_n_2332 ,csa_tree_add_6_33_groupi_n_2333);
  not csa_tree_add_6_33_groupi_g15947(csa_tree_add_6_33_groupi_n_2331 ,csa_tree_add_6_33_groupi_n_2330);
  not csa_tree_add_6_33_groupi_g15948(csa_tree_add_6_33_groupi_n_2328 ,csa_tree_add_6_33_groupi_n_2329);
  not csa_tree_add_6_33_groupi_g15949(csa_tree_add_6_33_groupi_n_2325 ,csa_tree_add_6_33_groupi_n_2326);
  or csa_tree_add_6_33_groupi_g15950(csa_tree_add_6_33_groupi_n_2324 ,csa_tree_add_6_33_groupi_n_1298 ,csa_tree_add_6_33_groupi_n_1999);
  or csa_tree_add_6_33_groupi_g15951(csa_tree_add_6_33_groupi_n_2323 ,csa_tree_add_6_33_groupi_n_1550 ,csa_tree_add_6_33_groupi_n_1880);
  or csa_tree_add_6_33_groupi_g15952(csa_tree_add_6_33_groupi_n_2322 ,csa_tree_add_6_33_groupi_n_1264 ,csa_tree_add_6_33_groupi_n_1678);
  or csa_tree_add_6_33_groupi_g15953(csa_tree_add_6_33_groupi_n_2321 ,csa_tree_add_6_33_groupi_n_1574 ,csa_tree_add_6_33_groupi_n_1663);
  or csa_tree_add_6_33_groupi_g15955(csa_tree_add_6_33_groupi_n_2319 ,csa_tree_add_6_33_groupi_n_1578 ,csa_tree_add_6_33_groupi_n_1862);
  or csa_tree_add_6_33_groupi_g15956(csa_tree_add_6_33_groupi_n_2318 ,csa_tree_add_6_33_groupi_n_1327 ,csa_tree_add_6_33_groupi_n_1988);
  or csa_tree_add_6_33_groupi_g15957(csa_tree_add_6_33_groupi_n_2317 ,csa_tree_add_6_33_groupi_n_1283 ,csa_tree_add_6_33_groupi_n_1665);
  or csa_tree_add_6_33_groupi_g15958(csa_tree_add_6_33_groupi_n_2316 ,csa_tree_add_6_33_groupi_n_1280 ,csa_tree_add_6_33_groupi_n_1987);
  or csa_tree_add_6_33_groupi_g15959(csa_tree_add_6_33_groupi_n_2315 ,csa_tree_add_6_33_groupi_n_1310 ,csa_tree_add_6_33_groupi_n_1921);
  or csa_tree_add_6_33_groupi_g15960(csa_tree_add_6_33_groupi_n_2314 ,csa_tree_add_6_33_groupi_n_1582 ,csa_tree_add_6_33_groupi_n_1832);
  or csa_tree_add_6_33_groupi_g15961(csa_tree_add_6_33_groupi_n_2313 ,csa_tree_add_6_33_groupi_n_1255 ,csa_tree_add_6_33_groupi_n_1845);
  or csa_tree_add_6_33_groupi_g15962(csa_tree_add_6_33_groupi_n_2312 ,csa_tree_add_6_33_groupi_n_1572 ,csa_tree_add_6_33_groupi_n_1878);
  or csa_tree_add_6_33_groupi_g15963(csa_tree_add_6_33_groupi_n_2311 ,csa_tree_add_6_33_groupi_n_1587 ,csa_tree_add_6_33_groupi_n_1971);
  or csa_tree_add_6_33_groupi_g15964(csa_tree_add_6_33_groupi_n_2310 ,csa_tree_add_6_33_groupi_n_1302 ,csa_tree_add_6_33_groupi_n_1827);
  or csa_tree_add_6_33_groupi_g15965(csa_tree_add_6_33_groupi_n_2309 ,csa_tree_add_6_33_groupi_n_1551 ,csa_tree_add_6_33_groupi_n_1929);
  or csa_tree_add_6_33_groupi_g15966(csa_tree_add_6_33_groupi_n_2308 ,csa_tree_add_6_33_groupi_n_1268 ,csa_tree_add_6_33_groupi_n_1664);
  or csa_tree_add_6_33_groupi_g15967(csa_tree_add_6_33_groupi_n_2307 ,csa_tree_add_6_33_groupi_n_1553 ,csa_tree_add_6_33_groupi_n_1945);
  or csa_tree_add_6_33_groupi_g15968(csa_tree_add_6_33_groupi_n_2306 ,csa_tree_add_6_33_groupi_n_1321 ,csa_tree_add_6_33_groupi_n_1659);
  or csa_tree_add_6_33_groupi_g15969(csa_tree_add_6_33_groupi_n_2305 ,csa_tree_add_6_33_groupi_n_1564 ,csa_tree_add_6_33_groupi_n_1737);
  or csa_tree_add_6_33_groupi_g15970(csa_tree_add_6_33_groupi_n_2304 ,csa_tree_add_6_33_groupi_n_1253 ,csa_tree_add_6_33_groupi_n_1978);
  or csa_tree_add_6_33_groupi_g15971(csa_tree_add_6_33_groupi_n_2303 ,csa_tree_add_6_33_groupi_n_1278 ,csa_tree_add_6_33_groupi_n_1947);
  or csa_tree_add_6_33_groupi_g15972(csa_tree_add_6_33_groupi_n_2302 ,csa_tree_add_6_33_groupi_n_1604 ,csa_tree_add_6_33_groupi_n_1954);
  or csa_tree_add_6_33_groupi_g15973(csa_tree_add_6_33_groupi_n_2301 ,csa_tree_add_6_33_groupi_n_1270 ,csa_tree_add_6_33_groupi_n_1823);
  or csa_tree_add_6_33_groupi_g15974(csa_tree_add_6_33_groupi_n_2300 ,csa_tree_add_6_33_groupi_n_1567 ,csa_tree_add_6_33_groupi_n_1910);
  or csa_tree_add_6_33_groupi_g15975(csa_tree_add_6_33_groupi_n_2299 ,csa_tree_add_6_33_groupi_n_1559 ,csa_tree_add_6_33_groupi_n_1669);
  or csa_tree_add_6_33_groupi_g15976(csa_tree_add_6_33_groupi_n_2298 ,csa_tree_add_6_33_groupi_n_1575 ,csa_tree_add_6_33_groupi_n_1840);
  or csa_tree_add_6_33_groupi_g15978(csa_tree_add_6_33_groupi_n_2296 ,csa_tree_add_6_33_groupi_n_1540 ,csa_tree_add_6_33_groupi_n_1943);
  or csa_tree_add_6_33_groupi_g15979(csa_tree_add_6_33_groupi_n_2295 ,csa_tree_add_6_33_groupi_n_1304 ,csa_tree_add_6_33_groupi_n_1944);
  or csa_tree_add_6_33_groupi_g15980(csa_tree_add_6_33_groupi_n_2294 ,csa_tree_add_6_33_groupi_n_1562 ,csa_tree_add_6_33_groupi_n_1674);
  or csa_tree_add_6_33_groupi_g15981(csa_tree_add_6_33_groupi_n_2293 ,csa_tree_add_6_33_groupi_n_1580 ,csa_tree_add_6_33_groupi_n_1833);
  or csa_tree_add_6_33_groupi_g15982(csa_tree_add_6_33_groupi_n_2292 ,csa_tree_add_6_33_groupi_n_1315 ,csa_tree_add_6_33_groupi_n_1975);
  or csa_tree_add_6_33_groupi_g15983(csa_tree_add_6_33_groupi_n_2291 ,csa_tree_add_6_33_groupi_n_1576 ,csa_tree_add_6_33_groupi_n_1812);
  or csa_tree_add_6_33_groupi_g15984(csa_tree_add_6_33_groupi_n_2290 ,csa_tree_add_6_33_groupi_n_1275 ,csa_tree_add_6_33_groupi_n_1740);
  or csa_tree_add_6_33_groupi_g15985(csa_tree_add_6_33_groupi_n_2289 ,csa_tree_add_6_33_groupi_n_1617 ,csa_tree_add_6_33_groupi_n_1843);
  or csa_tree_add_6_33_groupi_g15986(csa_tree_add_6_33_groupi_n_2288 ,csa_tree_add_6_33_groupi_n_1556 ,csa_tree_add_6_33_groupi_n_1983);
  or csa_tree_add_6_33_groupi_g15987(csa_tree_add_6_33_groupi_n_2287 ,csa_tree_add_6_33_groupi_n_1301 ,csa_tree_add_6_33_groupi_n_1931);
  or csa_tree_add_6_33_groupi_g15988(csa_tree_add_6_33_groupi_n_2286 ,csa_tree_add_6_33_groupi_n_1261 ,csa_tree_add_6_33_groupi_n_1778);
  or csa_tree_add_6_33_groupi_g15989(csa_tree_add_6_33_groupi_n_2285 ,csa_tree_add_6_33_groupi_n_1294 ,csa_tree_add_6_33_groupi_n_1869);
  or csa_tree_add_6_33_groupi_g15991(csa_tree_add_6_33_groupi_n_2283 ,csa_tree_add_6_33_groupi_n_1274 ,csa_tree_add_6_33_groupi_n_1989);
  or csa_tree_add_6_33_groupi_g15992(csa_tree_add_6_33_groupi_n_2282 ,csa_tree_add_6_33_groupi_n_1595 ,csa_tree_add_6_33_groupi_n_1949);
  or csa_tree_add_6_33_groupi_g15993(csa_tree_add_6_33_groupi_n_2281 ,csa_tree_add_6_33_groupi_n_1560 ,csa_tree_add_6_33_groupi_n_1696);
  or csa_tree_add_6_33_groupi_g15994(csa_tree_add_6_33_groupi_n_2280 ,csa_tree_add_6_33_groupi_n_1286 ,csa_tree_add_6_33_groupi_n_1716);
  or csa_tree_add_6_33_groupi_g15995(csa_tree_add_6_33_groupi_n_2279 ,csa_tree_add_6_33_groupi_n_1597 ,csa_tree_add_6_33_groupi_n_1690);
  or csa_tree_add_6_33_groupi_g15996(csa_tree_add_6_33_groupi_n_2278 ,csa_tree_add_6_33_groupi_n_1605 ,csa_tree_add_6_33_groupi_n_1738);
  or csa_tree_add_6_33_groupi_g15997(csa_tree_add_6_33_groupi_n_2277 ,csa_tree_add_6_33_groupi_n_1601 ,csa_tree_add_6_33_groupi_n_1763);
  or csa_tree_add_6_33_groupi_g15998(csa_tree_add_6_33_groupi_n_2276 ,csa_tree_add_6_33_groupi_n_1263 ,csa_tree_add_6_33_groupi_n_2013);
  or csa_tree_add_6_33_groupi_g16000(csa_tree_add_6_33_groupi_n_2274 ,csa_tree_add_6_33_groupi_n_1326 ,csa_tree_add_6_33_groupi_n_1746);
  or csa_tree_add_6_33_groupi_g16001(csa_tree_add_6_33_groupi_n_2273 ,csa_tree_add_6_33_groupi_n_1297 ,csa_tree_add_6_33_groupi_n_1689);
  or csa_tree_add_6_33_groupi_g16002(csa_tree_add_6_33_groupi_n_2272 ,csa_tree_add_6_33_groupi_n_1584 ,csa_tree_add_6_33_groupi_n_1655);
  or csa_tree_add_6_33_groupi_g16003(csa_tree_add_6_33_groupi_n_2271 ,csa_tree_add_6_33_groupi_n_1537 ,csa_tree_add_6_33_groupi_n_1948);
  or csa_tree_add_6_33_groupi_g16004(csa_tree_add_6_33_groupi_n_2270 ,csa_tree_add_6_33_groupi_n_1541 ,csa_tree_add_6_33_groupi_n_1951);
  or csa_tree_add_6_33_groupi_g16005(csa_tree_add_6_33_groupi_n_2269 ,csa_tree_add_6_33_groupi_n_1252 ,csa_tree_add_6_33_groupi_n_1901);
  or csa_tree_add_6_33_groupi_g16006(csa_tree_add_6_33_groupi_n_2268 ,csa_tree_add_6_33_groupi_n_1307 ,csa_tree_add_6_33_groupi_n_1932);
  or csa_tree_add_6_33_groupi_g16007(csa_tree_add_6_33_groupi_n_2267 ,csa_tree_add_6_33_groupi_n_1266 ,csa_tree_add_6_33_groupi_n_1960);
  or csa_tree_add_6_33_groupi_g16008(csa_tree_add_6_33_groupi_n_2266 ,csa_tree_add_6_33_groupi_n_1613 ,csa_tree_add_6_33_groupi_n_1851);
  or csa_tree_add_6_33_groupi_g16009(csa_tree_add_6_33_groupi_n_2265 ,csa_tree_add_6_33_groupi_n_1288 ,csa_tree_add_6_33_groupi_n_1861);
  or csa_tree_add_6_33_groupi_g16010(csa_tree_add_6_33_groupi_n_2264 ,csa_tree_add_6_33_groupi_n_1290 ,csa_tree_add_6_33_groupi_n_1718);
  or csa_tree_add_6_33_groupi_g16011(csa_tree_add_6_33_groupi_n_2263 ,csa_tree_add_6_33_groupi_n_1292 ,csa_tree_add_6_33_groupi_n_1881);
  or csa_tree_add_6_33_groupi_g16012(csa_tree_add_6_33_groupi_n_2262 ,csa_tree_add_6_33_groupi_n_1300 ,csa_tree_add_6_33_groupi_n_1857);
  or csa_tree_add_6_33_groupi_g16013(csa_tree_add_6_33_groupi_n_2261 ,csa_tree_add_6_33_groupi_n_1273 ,csa_tree_add_6_33_groupi_n_1801);
  or csa_tree_add_6_33_groupi_g16014(csa_tree_add_6_33_groupi_n_2260 ,csa_tree_add_6_33_groupi_n_1308 ,csa_tree_add_6_33_groupi_n_1875);
  or csa_tree_add_6_33_groupi_g16015(csa_tree_add_6_33_groupi_n_2259 ,csa_tree_add_6_33_groupi_n_1258 ,csa_tree_add_6_33_groupi_n_1858);
  or csa_tree_add_6_33_groupi_g16016(csa_tree_add_6_33_groupi_n_2258 ,csa_tree_add_6_33_groupi_n_1544 ,csa_tree_add_6_33_groupi_n_1970);
  or csa_tree_add_6_33_groupi_g16017(csa_tree_add_6_33_groupi_n_2257 ,csa_tree_add_6_33_groupi_n_1607 ,csa_tree_add_6_33_groupi_n_1772);
  or csa_tree_add_6_33_groupi_g16018(csa_tree_add_6_33_groupi_n_2256 ,csa_tree_add_6_33_groupi_n_1586 ,csa_tree_add_6_33_groupi_n_1854);
  or csa_tree_add_6_33_groupi_g16019(csa_tree_add_6_33_groupi_n_2255 ,csa_tree_add_6_33_groupi_n_1324 ,csa_tree_add_6_33_groupi_n_1760);
  or csa_tree_add_6_33_groupi_g16020(csa_tree_add_6_33_groupi_n_2254 ,csa_tree_add_6_33_groupi_n_1536 ,csa_tree_add_6_33_groupi_n_1766);
  or csa_tree_add_6_33_groupi_g16021(csa_tree_add_6_33_groupi_n_2253 ,csa_tree_add_6_33_groupi_n_1616 ,csa_tree_add_6_33_groupi_n_1797);
  or csa_tree_add_6_33_groupi_g16022(csa_tree_add_6_33_groupi_n_2252 ,csa_tree_add_6_33_groupi_n_1309 ,csa_tree_add_6_33_groupi_n_1841);
  or csa_tree_add_6_33_groupi_g16023(csa_tree_add_6_33_groupi_n_2251 ,csa_tree_add_6_33_groupi_n_1291 ,csa_tree_add_6_33_groupi_n_1727);
  or csa_tree_add_6_33_groupi_g16024(csa_tree_add_6_33_groupi_n_2250 ,csa_tree_add_6_33_groupi_n_1554 ,csa_tree_add_6_33_groupi_n_1676);
  or csa_tree_add_6_33_groupi_g16025(csa_tree_add_6_33_groupi_n_2249 ,csa_tree_add_6_33_groupi_n_1592 ,csa_tree_add_6_33_groupi_n_1969);
  or csa_tree_add_6_33_groupi_g16026(csa_tree_add_6_33_groupi_n_2248 ,csa_tree_add_6_33_groupi_n_1571 ,csa_tree_add_6_33_groupi_n_1692);
  or csa_tree_add_6_33_groupi_g16027(csa_tree_add_6_33_groupi_n_2247 ,csa_tree_add_6_33_groupi_n_1317 ,csa_tree_add_6_33_groupi_n_1751);
  or csa_tree_add_6_33_groupi_g16028(csa_tree_add_6_33_groupi_n_2246 ,csa_tree_add_6_33_groupi_n_1612 ,csa_tree_add_6_33_groupi_n_1821);
  or csa_tree_add_6_33_groupi_g16030(csa_tree_add_6_33_groupi_n_2244 ,csa_tree_add_6_33_groupi_n_1319 ,csa_tree_add_6_33_groupi_n_1691);
  or csa_tree_add_6_33_groupi_g16031(csa_tree_add_6_33_groupi_n_2243 ,csa_tree_add_6_33_groupi_n_1311 ,csa_tree_add_6_33_groupi_n_1786);
  or csa_tree_add_6_33_groupi_g16032(csa_tree_add_6_33_groupi_n_2242 ,csa_tree_add_6_33_groupi_n_1557 ,csa_tree_add_6_33_groupi_n_1775);
  or csa_tree_add_6_33_groupi_g16033(csa_tree_add_6_33_groupi_n_2241 ,csa_tree_add_6_33_groupi_n_1615 ,csa_tree_add_6_33_groupi_n_1836);
  or csa_tree_add_6_33_groupi_g16034(csa_tree_add_6_33_groupi_n_2240 ,csa_tree_add_6_33_groupi_n_1314 ,csa_tree_add_6_33_groupi_n_1876);
  or csa_tree_add_6_33_groupi_g16035(csa_tree_add_6_33_groupi_n_2239 ,csa_tree_add_6_33_groupi_n_1256 ,csa_tree_add_6_33_groupi_n_1791);
  or csa_tree_add_6_33_groupi_g16037(csa_tree_add_6_33_groupi_n_2237 ,csa_tree_add_6_33_groupi_n_1565 ,csa_tree_add_6_33_groupi_n_1818);
  or csa_tree_add_6_33_groupi_g16038(csa_tree_add_6_33_groupi_n_2236 ,csa_tree_add_6_33_groupi_n_1269 ,csa_tree_add_6_33_groupi_n_1898);
  or csa_tree_add_6_33_groupi_g16039(csa_tree_add_6_33_groupi_n_2235 ,csa_tree_add_6_33_groupi_n_1602 ,csa_tree_add_6_33_groupi_n_1813);
  or csa_tree_add_6_33_groupi_g16040(csa_tree_add_6_33_groupi_n_2234 ,csa_tree_add_6_33_groupi_n_1608 ,csa_tree_add_6_33_groupi_n_1913);
  or csa_tree_add_6_33_groupi_g16041(csa_tree_add_6_33_groupi_n_2233 ,csa_tree_add_6_33_groupi_n_1585 ,csa_tree_add_6_33_groupi_n_1831);
  or csa_tree_add_6_33_groupi_g16042(csa_tree_add_6_33_groupi_n_2232 ,csa_tree_add_6_33_groupi_n_1260 ,csa_tree_add_6_33_groupi_n_1805);
  or csa_tree_add_6_33_groupi_g16043(csa_tree_add_6_33_groupi_n_2231 ,csa_tree_add_6_33_groupi_n_1603 ,csa_tree_add_6_33_groupi_n_1981);
  or csa_tree_add_6_33_groupi_g16044(csa_tree_add_6_33_groupi_n_2230 ,csa_tree_add_6_33_groupi_n_1594 ,csa_tree_add_6_33_groupi_n_1713);
  or csa_tree_add_6_33_groupi_g16045(csa_tree_add_6_33_groupi_n_2229 ,csa_tree_add_6_33_groupi_n_1589 ,csa_tree_add_6_33_groupi_n_1804);
  or csa_tree_add_6_33_groupi_g16046(csa_tree_add_6_33_groupi_n_2228 ,csa_tree_add_6_33_groupi_n_1259 ,csa_tree_add_6_33_groupi_n_1764);
  or csa_tree_add_6_33_groupi_g16047(csa_tree_add_6_33_groupi_n_2227 ,csa_tree_add_6_33_groupi_n_1614 ,csa_tree_add_6_33_groupi_n_1777);
  or csa_tree_add_6_33_groupi_g16048(csa_tree_add_6_33_groupi_n_2226 ,csa_tree_add_6_33_groupi_n_1579 ,csa_tree_add_6_33_groupi_n_1814);
  or csa_tree_add_6_33_groupi_g16049(csa_tree_add_6_33_groupi_n_2225 ,csa_tree_add_6_33_groupi_n_1323 ,csa_tree_add_6_33_groupi_n_1720);
  or csa_tree_add_6_33_groupi_g16050(csa_tree_add_6_33_groupi_n_2224 ,csa_tree_add_6_33_groupi_n_1299 ,csa_tree_add_6_33_groupi_n_1811);
  or csa_tree_add_6_33_groupi_g16051(csa_tree_add_6_33_groupi_n_2223 ,csa_tree_add_6_33_groupi_n_1287 ,csa_tree_add_6_33_groupi_n_1825);
  or csa_tree_add_6_33_groupi_g16052(csa_tree_add_6_33_groupi_n_2222 ,csa_tree_add_6_33_groupi_n_1303 ,csa_tree_add_6_33_groupi_n_1782);
  or csa_tree_add_6_33_groupi_g16053(csa_tree_add_6_33_groupi_n_2221 ,csa_tree_add_6_33_groupi_n_1606 ,csa_tree_add_6_33_groupi_n_1788);
  or csa_tree_add_6_33_groupi_g16055(csa_tree_add_6_33_groupi_n_2219 ,csa_tree_add_6_33_groupi_n_1254 ,csa_tree_add_6_33_groupi_n_1771);
  or csa_tree_add_6_33_groupi_g16056(csa_tree_add_6_33_groupi_n_2218 ,csa_tree_add_6_33_groupi_n_1312 ,csa_tree_add_6_33_groupi_n_1903);
  or csa_tree_add_6_33_groupi_g16057(csa_tree_add_6_33_groupi_n_2217 ,csa_tree_add_6_33_groupi_n_1573 ,csa_tree_add_6_33_groupi_n_1934);
  or csa_tree_add_6_33_groupi_g16058(csa_tree_add_6_33_groupi_n_2216 ,csa_tree_add_6_33_groupi_n_1257 ,csa_tree_add_6_33_groupi_n_1941);
  or csa_tree_add_6_33_groupi_g16059(csa_tree_add_6_33_groupi_n_2215 ,csa_tree_add_6_33_groupi_n_1289 ,csa_tree_add_6_33_groupi_n_1723);
  or csa_tree_add_6_33_groupi_g16060(csa_tree_add_6_33_groupi_n_2214 ,csa_tree_add_6_33_groupi_n_1618 ,csa_tree_add_6_33_groupi_n_1769);
  or csa_tree_add_6_33_groupi_g16061(csa_tree_add_6_33_groupi_n_2213 ,csa_tree_add_6_33_groupi_n_1271 ,csa_tree_add_6_33_groupi_n_1952);
  or csa_tree_add_6_33_groupi_g16062(csa_tree_add_6_33_groupi_n_2212 ,csa_tree_add_6_33_groupi_n_1591 ,csa_tree_add_6_33_groupi_n_1911);
  or csa_tree_add_6_33_groupi_g16063(csa_tree_add_6_33_groupi_n_2211 ,csa_tree_add_6_33_groupi_n_1599 ,csa_tree_add_6_33_groupi_n_1935);
  or csa_tree_add_6_33_groupi_g16064(csa_tree_add_6_33_groupi_n_2210 ,csa_tree_add_6_33_groupi_n_1610 ,csa_tree_add_6_33_groupi_n_1982);
  or csa_tree_add_6_33_groupi_g16067(csa_tree_add_6_33_groupi_n_2207 ,csa_tree_add_6_33_groupi_n_1282 ,csa_tree_add_6_33_groupi_n_1762);
  or csa_tree_add_6_33_groupi_g16068(csa_tree_add_6_33_groupi_n_2206 ,csa_tree_add_6_33_groupi_n_1549 ,csa_tree_add_6_33_groupi_n_1680);
  or csa_tree_add_6_33_groupi_g16069(csa_tree_add_6_33_groupi_n_2205 ,csa_tree_add_6_33_groupi_n_1276 ,csa_tree_add_6_33_groupi_n_1748);
  or csa_tree_add_6_33_groupi_g16070(csa_tree_add_6_33_groupi_n_2204 ,csa_tree_add_6_33_groupi_n_1542 ,csa_tree_add_6_33_groupi_n_1856);
  or csa_tree_add_6_33_groupi_g16071(csa_tree_add_6_33_groupi_n_2203 ,csa_tree_add_6_33_groupi_n_1318 ,csa_tree_add_6_33_groupi_n_1741);
  or csa_tree_add_6_33_groupi_g16072(csa_tree_add_6_33_groupi_n_2202 ,csa_tree_add_6_33_groupi_n_1611 ,csa_tree_add_6_33_groupi_n_1711);
  or csa_tree_add_6_33_groupi_g16073(csa_tree_add_6_33_groupi_n_2201 ,csa_tree_add_6_33_groupi_n_1277 ,csa_tree_add_6_33_groupi_n_1800);
  or csa_tree_add_6_33_groupi_g16074(csa_tree_add_6_33_groupi_n_2200 ,csa_tree_add_6_33_groupi_n_1545 ,csa_tree_add_6_33_groupi_n_1666);
  or csa_tree_add_6_33_groupi_g16075(csa_tree_add_6_33_groupi_n_2199 ,csa_tree_add_6_33_groupi_n_1577 ,csa_tree_add_6_33_groupi_n_1866);
  or csa_tree_add_6_33_groupi_g16076(csa_tree_add_6_33_groupi_n_2198 ,csa_tree_add_6_33_groupi_n_1609 ,csa_tree_add_6_33_groupi_n_1679);
  or csa_tree_add_6_33_groupi_g16077(csa_tree_add_6_33_groupi_n_2197 ,csa_tree_add_6_33_groupi_n_1588 ,csa_tree_add_6_33_groupi_n_1701);
  or csa_tree_add_6_33_groupi_g16078(csa_tree_add_6_33_groupi_n_2196 ,csa_tree_add_6_33_groupi_n_1267 ,csa_tree_add_6_33_groupi_n_1864);
  or csa_tree_add_6_33_groupi_g16079(csa_tree_add_6_33_groupi_n_2195 ,csa_tree_add_6_33_groupi_n_1548 ,csa_tree_add_6_33_groupi_n_1795);
  or csa_tree_add_6_33_groupi_g16080(csa_tree_add_6_33_groupi_n_2194 ,csa_tree_add_6_33_groupi_n_1305 ,csa_tree_add_6_33_groupi_n_1985);
  or csa_tree_add_6_33_groupi_g16081(csa_tree_add_6_33_groupi_n_2193 ,csa_tree_add_6_33_groupi_n_1552 ,csa_tree_add_6_33_groupi_n_1780);
  or csa_tree_add_6_33_groupi_g16082(csa_tree_add_6_33_groupi_n_2192 ,csa_tree_add_6_33_groupi_n_1306 ,csa_tree_add_6_33_groupi_n_1871);
  or csa_tree_add_6_33_groupi_g16083(csa_tree_add_6_33_groupi_n_2191 ,csa_tree_add_6_33_groupi_n_1590 ,csa_tree_add_6_33_groupi_n_1658);
  or csa_tree_add_6_33_groupi_g16084(csa_tree_add_6_33_groupi_n_2190 ,csa_tree_add_6_33_groupi_n_1325 ,csa_tree_add_6_33_groupi_n_1909);
  or csa_tree_add_6_33_groupi_g16085(csa_tree_add_6_33_groupi_n_2189 ,csa_tree_add_6_33_groupi_n_1583 ,csa_tree_add_6_33_groupi_n_1750);
  or csa_tree_add_6_33_groupi_g16086(csa_tree_add_6_33_groupi_n_2188 ,csa_tree_add_6_33_groupi_n_1284 ,csa_tree_add_6_33_groupi_n_1923);
  or csa_tree_add_6_33_groupi_g16087(csa_tree_add_6_33_groupi_n_2187 ,csa_tree_add_6_33_groupi_n_1296 ,csa_tree_add_6_33_groupi_n_1817);
  or csa_tree_add_6_33_groupi_g16088(csa_tree_add_6_33_groupi_n_2186 ,csa_tree_add_6_33_groupi_n_1546 ,csa_tree_add_6_33_groupi_n_1721);
  or csa_tree_add_6_33_groupi_g16089(csa_tree_add_6_33_groupi_n_2185 ,csa_tree_add_6_33_groupi_n_1272 ,csa_tree_add_6_33_groupi_n_1837);
  or csa_tree_add_6_33_groupi_g16090(csa_tree_add_6_33_groupi_n_2368 ,csa_tree_add_6_33_groupi_n_1063 ,csa_tree_add_6_33_groupi_n_2009);
  or csa_tree_add_6_33_groupi_g16091(csa_tree_add_6_33_groupi_n_2367 ,csa_tree_add_6_33_groupi_n_1049 ,csa_tree_add_6_33_groupi_n_1915);
  and csa_tree_add_6_33_groupi_g16092(csa_tree_add_6_33_groupi_n_2366 ,csa_tree_add_6_33_groupi_n_1067 ,csa_tree_add_6_33_groupi_n_1747);
  or csa_tree_add_6_33_groupi_g16093(csa_tree_add_6_33_groupi_n_2365 ,csa_tree_add_6_33_groupi_n_1342 ,csa_tree_add_6_33_groupi_n_1798);
  or csa_tree_add_6_33_groupi_g16094(csa_tree_add_6_33_groupi_n_2364 ,csa_tree_add_6_33_groupi_n_1058 ,csa_tree_add_6_33_groupi_n_1756);
  and csa_tree_add_6_33_groupi_g16095(csa_tree_add_6_33_groupi_n_2363 ,csa_tree_add_6_33_groupi_n_1044 ,csa_tree_add_6_33_groupi_n_2004);
  or csa_tree_add_6_33_groupi_g16096(csa_tree_add_6_33_groupi_n_2362 ,csa_tree_add_6_33_groupi_n_1338 ,csa_tree_add_6_33_groupi_n_1889);
  or csa_tree_add_6_33_groupi_g16097(csa_tree_add_6_33_groupi_n_2360 ,csa_tree_add_6_33_groupi_n_1052 ,csa_tree_add_6_33_groupi_n_2012);
  or csa_tree_add_6_33_groupi_g16098(csa_tree_add_6_33_groupi_n_2358 ,csa_tree_add_6_33_groupi_n_1341 ,csa_tree_add_6_33_groupi_n_1675);
  and csa_tree_add_6_33_groupi_g16099(csa_tree_add_6_33_groupi_n_2357 ,csa_tree_add_6_33_groupi_n_1352 ,csa_tree_add_6_33_groupi_n_1946);
  or csa_tree_add_6_33_groupi_g16100(csa_tree_add_6_33_groupi_n_2355 ,csa_tree_add_6_33_groupi_n_1353 ,csa_tree_add_6_33_groupi_n_1652);
  or csa_tree_add_6_33_groupi_g16101(csa_tree_add_6_33_groupi_n_2353 ,csa_tree_add_6_33_groupi_n_1053 ,csa_tree_add_6_33_groupi_n_2001);
  or csa_tree_add_6_33_groupi_g16102(csa_tree_add_6_33_groupi_n_2352 ,csa_tree_add_6_33_groupi_n_1358 ,csa_tree_add_6_33_groupi_n_2011);
  or csa_tree_add_6_33_groupi_g16103(csa_tree_add_6_33_groupi_n_2351 ,csa_tree_add_6_33_groupi_n_1048 ,csa_tree_add_6_33_groupi_n_2005);
  or csa_tree_add_6_33_groupi_g16104(csa_tree_add_6_33_groupi_n_2349 ,csa_tree_add_6_33_groupi_n_1359 ,csa_tree_add_6_33_groupi_n_1926);
  or csa_tree_add_6_33_groupi_g16105(csa_tree_add_6_33_groupi_n_2348 ,csa_tree_add_6_33_groupi_n_1330 ,csa_tree_add_6_33_groupi_n_1950);
  or csa_tree_add_6_33_groupi_g16106(csa_tree_add_6_33_groupi_n_2346 ,csa_tree_add_6_33_groupi_n_1047 ,csa_tree_add_6_33_groupi_n_1918);
  or csa_tree_add_6_33_groupi_g16107(csa_tree_add_6_33_groupi_n_2344 ,csa_tree_add_6_33_groupi_n_1050 ,csa_tree_add_6_33_groupi_n_2002);
  or csa_tree_add_6_33_groupi_g16108(csa_tree_add_6_33_groupi_n_2342 ,csa_tree_add_6_33_groupi_n_1344 ,csa_tree_add_6_33_groupi_n_2006);
  and csa_tree_add_6_33_groupi_g16109(csa_tree_add_6_33_groupi_n_2340 ,csa_tree_add_6_33_groupi_n_1062 ,csa_tree_add_6_33_groupi_n_1933);
  or csa_tree_add_6_33_groupi_g16110(csa_tree_add_6_33_groupi_n_2339 ,csa_tree_add_6_33_groupi_n_1363 ,csa_tree_add_6_33_groupi_n_1963);
  or csa_tree_add_6_33_groupi_g16111(csa_tree_add_6_33_groupi_n_2338 ,csa_tree_add_6_33_groupi_n_1329 ,csa_tree_add_6_33_groupi_n_1955);
  and csa_tree_add_6_33_groupi_g16112(csa_tree_add_6_33_groupi_n_2337 ,csa_tree_add_6_33_groupi_n_1046 ,csa_tree_add_6_33_groupi_n_1735);
  and csa_tree_add_6_33_groupi_g16113(csa_tree_add_6_33_groupi_n_2336 ,csa_tree_add_6_33_groupi_n_1336 ,csa_tree_add_6_33_groupi_n_1884);
  and csa_tree_add_6_33_groupi_g16114(csa_tree_add_6_33_groupi_n_2335 ,csa_tree_add_6_33_groupi_n_1066 ,csa_tree_add_6_33_groupi_n_1868);
  and csa_tree_add_6_33_groupi_g16115(csa_tree_add_6_33_groupi_n_2334 ,csa_tree_add_6_33_groupi_n_1069 ,csa_tree_add_6_33_groupi_n_1707);
  or csa_tree_add_6_33_groupi_g16116(csa_tree_add_6_33_groupi_n_2333 ,csa_tree_add_6_33_groupi_n_1045 ,csa_tree_add_6_33_groupi_n_2008);
  or csa_tree_add_6_33_groupi_g16117(csa_tree_add_6_33_groupi_n_2330 ,csa_tree_add_6_33_groupi_n_1068 ,csa_tree_add_6_33_groupi_n_2010);
  or csa_tree_add_6_33_groupi_g16118(csa_tree_add_6_33_groupi_n_2329 ,csa_tree_add_6_33_groupi_n_1360 ,csa_tree_add_6_33_groupi_n_2003);
  and csa_tree_add_6_33_groupi_g16119(csa_tree_add_6_33_groupi_n_2327 ,csa_tree_add_6_33_groupi_n_1054 ,csa_tree_add_6_33_groupi_n_1715);
  or csa_tree_add_6_33_groupi_g16120(csa_tree_add_6_33_groupi_n_2326 ,csa_tree_add_6_33_groupi_n_1051 ,csa_tree_add_6_33_groupi_n_2007);
  or csa_tree_add_6_33_groupi_g16121(csa_tree_add_6_33_groupi_n_2184 ,csa_tree_add_6_33_groupi_n_1322 ,csa_tree_add_6_33_groupi_n_1700);
  or csa_tree_add_6_33_groupi_g16122(csa_tree_add_6_33_groupi_n_2183 ,csa_tree_add_6_33_groupi_n_1293 ,csa_tree_add_6_33_groupi_n_1651);
  or csa_tree_add_6_33_groupi_g16123(csa_tree_add_6_33_groupi_n_2182 ,csa_tree_add_6_33_groupi_n_1596 ,csa_tree_add_6_33_groupi_n_1693);
  or csa_tree_add_6_33_groupi_g16124(csa_tree_add_6_33_groupi_n_2181 ,csa_tree_add_6_33_groupi_n_1555 ,csa_tree_add_6_33_groupi_n_1964);
  or csa_tree_add_6_33_groupi_g16125(csa_tree_add_6_33_groupi_n_2180 ,csa_tree_add_6_33_groupi_n_1538 ,csa_tree_add_6_33_groupi_n_1755);
  xnor csa_tree_add_6_33_groupi_g16126(csa_tree_add_6_33_groupi_n_2179 ,csa_tree_add_6_33_groupi_n_1509 ,csa_tree_add_6_33_groupi_n_1210);
  xnor csa_tree_add_6_33_groupi_g16127(csa_tree_add_6_33_groupi_n_2178 ,csa_tree_add_6_33_groupi_n_1285 ,in1[25]);
  xnor csa_tree_add_6_33_groupi_g16128(csa_tree_add_6_33_groupi_n_2177 ,csa_tree_add_6_33_groupi_n_1245 ,in1[31]);
  xnor csa_tree_add_6_33_groupi_g16129(csa_tree_add_6_33_groupi_n_2176 ,csa_tree_add_6_33_groupi_n_1547 ,in1[26]);
  xnor csa_tree_add_6_33_groupi_g16130(csa_tree_add_6_33_groupi_n_2175 ,csa_tree_add_6_33_groupi_n_1313 ,in1[22]);
  xnor csa_tree_add_6_33_groupi_g16131(csa_tree_add_6_33_groupi_n_2174 ,csa_tree_add_6_33_groupi_n_1263 ,in1[30]);
  xnor csa_tree_add_6_33_groupi_g16132(csa_tree_add_6_33_groupi_n_2173 ,csa_tree_add_6_33_groupi_n_1279 ,in1[19]);
  xnor csa_tree_add_6_33_groupi_g16133(csa_tree_add_6_33_groupi_n_2172 ,csa_tree_add_6_33_groupi_n_1598 ,in1[23]);
  xnor csa_tree_add_6_33_groupi_g16134(csa_tree_add_6_33_groupi_n_2171 ,csa_tree_add_6_33_groupi_n_1574 ,in1[21]);
  xnor csa_tree_add_6_33_groupi_g16135(csa_tree_add_6_33_groupi_n_2170 ,csa_tree_add_6_33_groupi_n_1265 ,in1[27]);
  xnor csa_tree_add_6_33_groupi_g16136(csa_tree_add_6_33_groupi_n_2169 ,csa_tree_add_6_33_groupi_n_1568 ,in1[16]);
  xnor csa_tree_add_6_33_groupi_g16137(csa_tree_add_6_33_groupi_n_2168 ,csa_tree_add_6_33_groupi_n_1310 ,in1[24]);
  xnor csa_tree_add_6_33_groupi_g16138(csa_tree_add_6_33_groupi_n_2167 ,csa_tree_add_6_33_groupi_n_1539 ,in1[28]);
  xnor csa_tree_add_6_33_groupi_g16139(csa_tree_add_6_33_groupi_n_2166 ,csa_tree_add_6_33_groupi_n_1615 ,in1[18]);
  xnor csa_tree_add_6_33_groupi_g16140(csa_tree_add_6_33_groupi_n_2165 ,csa_tree_add_6_33_groupi_n_1261 ,in1[20]);
  xnor csa_tree_add_6_33_groupi_g16141(csa_tree_add_6_33_groupi_n_2164 ,csa_tree_add_6_33_groupi_n_1089 ,csa_tree_add_6_33_groupi_n_1117);
  xnor csa_tree_add_6_33_groupi_g16142(csa_tree_add_6_33_groupi_n_2163 ,csa_tree_add_6_33_groupi_n_1146 ,csa_tree_add_6_33_groupi_n_1491);
  xnor csa_tree_add_6_33_groupi_g16143(csa_tree_add_6_33_groupi_n_2162 ,csa_tree_add_6_33_groupi_n_1372 ,csa_tree_add_6_33_groupi_n_1380);
  xnor csa_tree_add_6_33_groupi_g16144(csa_tree_add_6_33_groupi_n_2161 ,csa_tree_add_6_33_groupi_n_1078 ,csa_tree_add_6_33_groupi_n_1583);
  xnor csa_tree_add_6_33_groupi_g16145(csa_tree_add_6_33_groupi_n_2160 ,csa_tree_add_6_33_groupi_n_1217 ,csa_tree_add_6_33_groupi_n_1592);
  xnor csa_tree_add_6_33_groupi_g16146(csa_tree_add_6_33_groupi_n_2159 ,csa_tree_add_6_33_groupi_n_1087 ,csa_tree_add_6_33_groupi_n_1151);
  xnor csa_tree_add_6_33_groupi_g16147(csa_tree_add_6_33_groupi_n_2158 ,csa_tree_add_6_33_groupi_n_1473 ,csa_tree_add_6_33_groupi_n_1594);
  xnor csa_tree_add_6_33_groupi_g16148(csa_tree_add_6_33_groupi_n_2157 ,csa_tree_add_6_33_groupi_n_1520 ,csa_tree_add_6_33_groupi_n_1604);
  xnor csa_tree_add_6_33_groupi_g16149(csa_tree_add_6_33_groupi_n_2156 ,csa_tree_add_6_33_groupi_n_1254 ,csa_tree_add_6_33_groupi_n_1172);
  xnor csa_tree_add_6_33_groupi_g16150(csa_tree_add_6_33_groupi_n_2155 ,csa_tree_add_6_33_groupi_n_1425 ,csa_tree_add_6_33_groupi_n_1535);
  xnor csa_tree_add_6_33_groupi_g16151(csa_tree_add_6_33_groupi_n_2154 ,csa_tree_add_6_33_groupi_n_1455 ,csa_tree_add_6_33_groupi_n_1167);
  xnor csa_tree_add_6_33_groupi_g16152(csa_tree_add_6_33_groupi_n_2153 ,csa_tree_add_6_33_groupi_n_1432 ,csa_tree_add_6_33_groupi_n_1148);
  xnor csa_tree_add_6_33_groupi_g16153(csa_tree_add_6_33_groupi_n_2152 ,csa_tree_add_6_33_groupi_n_1526 ,csa_tree_add_6_33_groupi_n_1278);
  xnor csa_tree_add_6_33_groupi_g16154(csa_tree_add_6_33_groupi_n_2151 ,csa_tree_add_6_33_groupi_n_1499 ,csa_tree_add_6_33_groupi_n_1266);
  xnor csa_tree_add_6_33_groupi_g16155(csa_tree_add_6_33_groupi_n_2150 ,csa_tree_add_6_33_groupi_n_1288 ,csa_tree_add_6_33_groupi_n_1216);
  xnor csa_tree_add_6_33_groupi_g16156(csa_tree_add_6_33_groupi_n_2149 ,csa_tree_add_6_33_groupi_n_1113 ,csa_tree_add_6_33_groupi_n_1384);
  xnor csa_tree_add_6_33_groupi_g16157(csa_tree_add_6_33_groupi_n_2148 ,csa_tree_add_6_33_groupi_n_1371 ,csa_tree_add_6_33_groupi_n_1267);
  xnor csa_tree_add_6_33_groupi_g16158(csa_tree_add_6_33_groupi_n_2147 ,csa_tree_add_6_33_groupi_n_1493 ,csa_tree_add_6_33_groupi_n_1158);
  xnor csa_tree_add_6_33_groupi_g16159(csa_tree_add_6_33_groupi_n_2146 ,csa_tree_add_6_33_groupi_n_1213 ,csa_tree_add_6_33_groupi_n_1546);
  xnor csa_tree_add_6_33_groupi_g16160(csa_tree_add_6_33_groupi_n_2145 ,csa_tree_add_6_33_groupi_n_1460 ,csa_tree_add_6_33_groupi_n_1420);
  xnor csa_tree_add_6_33_groupi_g16161(csa_tree_add_6_33_groupi_n_2144 ,csa_tree_add_6_33_groupi_n_1442 ,csa_tree_add_6_33_groupi_n_1611);
  xnor csa_tree_add_6_33_groupi_g16162(csa_tree_add_6_33_groupi_n_2143 ,csa_tree_add_6_33_groupi_n_1304 ,csa_tree_add_6_33_groupi_n_1530);
  xnor csa_tree_add_6_33_groupi_g16163(csa_tree_add_6_33_groupi_n_2142 ,csa_tree_add_6_33_groupi_n_1147 ,csa_tree_add_6_33_groupi_n_1273);
  xnor csa_tree_add_6_33_groupi_g16164(csa_tree_add_6_33_groupi_n_2141 ,csa_tree_add_6_33_groupi_n_1161 ,csa_tree_add_6_33_groupi_n_1477);
  xnor csa_tree_add_6_33_groupi_g16165(csa_tree_add_6_33_groupi_n_2140 ,csa_tree_add_6_33_groupi_n_1208 ,csa_tree_add_6_33_groupi_n_1306);
  xnor csa_tree_add_6_33_groupi_g16166(csa_tree_add_6_33_groupi_n_2139 ,csa_tree_add_6_33_groupi_n_1192 ,csa_tree_add_6_33_groupi_n_1174);
  xnor csa_tree_add_6_33_groupi_g16167(csa_tree_add_6_33_groupi_n_2138 ,csa_tree_add_6_33_groupi_n_1429 ,csa_tree_add_6_33_groupi_n_1584);
  xnor csa_tree_add_6_33_groupi_g16168(csa_tree_add_6_33_groupi_n_2137 ,csa_tree_add_6_33_groupi_n_1489 ,csa_tree_add_6_33_groupi_n_1252);
  xnor csa_tree_add_6_33_groupi_g16169(csa_tree_add_6_33_groupi_n_2136 ,csa_tree_add_6_33_groupi_n_1459 ,csa_tree_add_6_33_groupi_n_1580);
  xnor csa_tree_add_6_33_groupi_g16170(csa_tree_add_6_33_groupi_n_2135 ,csa_tree_add_6_33_groupi_n_1196 ,csa_tree_add_6_33_groupi_n_1606);
  xnor csa_tree_add_6_33_groupi_g16171(csa_tree_add_6_33_groupi_n_2134 ,csa_tree_add_6_33_groupi_n_1234 ,csa_tree_add_6_33_groupi_n_1319);
  xnor csa_tree_add_6_33_groupi_g16172(csa_tree_add_6_33_groupi_n_2133 ,csa_tree_add_6_33_groupi_n_1181 ,csa_tree_add_6_33_groupi_n_1300);
  xnor csa_tree_add_6_33_groupi_g16173(csa_tree_add_6_33_groupi_n_2132 ,csa_tree_add_6_33_groupi_n_1233 ,csa_tree_add_6_33_groupi_n_1452);
  xnor csa_tree_add_6_33_groupi_g16174(csa_tree_add_6_33_groupi_n_2131 ,csa_tree_add_6_33_groupi_n_1486 ,csa_tree_add_6_33_groupi_n_1205);
  xnor csa_tree_add_6_33_groupi_g16175(csa_tree_add_6_33_groupi_n_2130 ,csa_tree_add_6_33_groupi_n_1073 ,csa_tree_add_6_33_groupi_n_1110);
  xnor csa_tree_add_6_33_groupi_g16176(csa_tree_add_6_33_groupi_n_2129 ,csa_tree_add_6_33_groupi_n_1099 ,csa_tree_add_6_33_groupi_n_1189);
  xnor csa_tree_add_6_33_groupi_g16177(csa_tree_add_6_33_groupi_n_2128 ,csa_tree_add_6_33_groupi_n_1497 ,csa_tree_add_6_33_groupi_n_1187);
  xnor csa_tree_add_6_33_groupi_g16178(csa_tree_add_6_33_groupi_n_2127 ,csa_tree_add_6_33_groupi_n_1492 ,csa_tree_add_6_33_groupi_n_1613);
  xnor csa_tree_add_6_33_groupi_g16179(csa_tree_add_6_33_groupi_n_2126 ,csa_tree_add_6_33_groupi_n_1226 ,csa_tree_add_6_33_groupi_n_1321);
  xnor csa_tree_add_6_33_groupi_g16180(csa_tree_add_6_33_groupi_n_2125 ,csa_tree_add_6_33_groupi_n_1275 ,csa_tree_add_6_33_groupi_n_1109);
  xnor csa_tree_add_6_33_groupi_g16181(csa_tree_add_6_33_groupi_n_2124 ,csa_tree_add_6_33_groupi_n_1202 ,csa_tree_add_6_33_groupi_n_1367);
  xnor csa_tree_add_6_33_groupi_g16182(csa_tree_add_6_33_groupi_n_2123 ,csa_tree_add_6_33_groupi_n_1595 ,csa_tree_add_6_33_groupi_n_1436);
  xnor csa_tree_add_6_33_groupi_g16183(csa_tree_add_6_33_groupi_n_2122 ,csa_tree_add_6_33_groupi_n_1482 ,csa_tree_add_6_33_groupi_n_1577);
  xnor csa_tree_add_6_33_groupi_g16184(csa_tree_add_6_33_groupi_n_2121 ,csa_tree_add_6_33_groupi_n_1529 ,csa_tree_add_6_33_groupi_n_1204);
  xnor csa_tree_add_6_33_groupi_g16185(csa_tree_add_6_33_groupi_n_2120 ,csa_tree_add_6_33_groupi_n_1085 ,csa_tree_add_6_33_groupi_n_1299);
  xnor csa_tree_add_6_33_groupi_g16186(csa_tree_add_6_33_groupi_n_2119 ,csa_tree_add_6_33_groupi_n_1506 ,csa_tree_add_6_33_groupi_n_1080);
  xnor csa_tree_add_6_33_groupi_g16187(csa_tree_add_6_33_groupi_n_2118 ,csa_tree_add_6_33_groupi_n_1527 ,csa_tree_add_6_33_groupi_n_1618);
  xnor csa_tree_add_6_33_groupi_g16188(csa_tree_add_6_33_groupi_n_2117 ,csa_tree_add_6_33_groupi_n_1168 ,csa_tree_add_6_33_groupi_n_1242);
  xnor csa_tree_add_6_33_groupi_g16189(csa_tree_add_6_33_groupi_n_2116 ,csa_tree_add_6_33_groupi_n_1507 ,csa_tree_add_6_33_groupi_n_1431);
  xnor csa_tree_add_6_33_groupi_g16190(csa_tree_add_6_33_groupi_n_2115 ,csa_tree_add_6_33_groupi_n_1175 ,csa_tree_add_6_33_groupi_n_1224);
  xnor csa_tree_add_6_33_groupi_g16191(csa_tree_add_6_33_groupi_n_2114 ,csa_tree_add_6_33_groupi_n_1292 ,csa_tree_add_6_33_groupi_n_1222);
  xnor csa_tree_add_6_33_groupi_g16192(csa_tree_add_6_33_groupi_n_2113 ,csa_tree_add_6_33_groupi_n_1597 ,csa_tree_add_6_33_groupi_n_1127);
  xnor csa_tree_add_6_33_groupi_g16193(csa_tree_add_6_33_groupi_n_2112 ,csa_tree_add_6_33_groupi_n_1092 ,csa_tree_add_6_33_groupi_n_1556);
  xnor csa_tree_add_6_33_groupi_g16194(csa_tree_add_6_33_groupi_n_2111 ,csa_tree_add_6_33_groupi_n_1465 ,csa_tree_add_6_33_groupi_n_1255);
  xnor csa_tree_add_6_33_groupi_g16195(csa_tree_add_6_33_groupi_n_2110 ,csa_tree_add_6_33_groupi_n_1139 ,csa_tree_add_6_33_groupi_n_1439);
  xnor csa_tree_add_6_33_groupi_g16196(csa_tree_add_6_33_groupi_n_2109 ,csa_tree_add_6_33_groupi_n_1203 ,csa_tree_add_6_33_groupi_n_1141);
  xnor csa_tree_add_6_33_groupi_g16197(csa_tree_add_6_33_groupi_n_2108 ,csa_tree_add_6_33_groupi_n_1400 ,csa_tree_add_6_33_groupi_n_1107);
  xnor csa_tree_add_6_33_groupi_g16198(csa_tree_add_6_33_groupi_n_2107 ,csa_tree_add_6_33_groupi_n_1191 ,csa_tree_add_6_33_groupi_n_1315);
  xnor csa_tree_add_6_33_groupi_g16199(csa_tree_add_6_33_groupi_n_2106 ,csa_tree_add_6_33_groupi_n_1394 ,csa_tree_add_6_33_groupi_n_1541);
  xnor csa_tree_add_6_33_groupi_g16200(csa_tree_add_6_33_groupi_n_2105 ,csa_tree_add_6_33_groupi_n_1121 ,csa_tree_add_6_33_groupi_n_1298);
  xnor csa_tree_add_6_33_groupi_g16201(csa_tree_add_6_33_groupi_n_2104 ,csa_tree_add_6_33_groupi_n_1610 ,csa_tree_add_6_33_groupi_n_1130);
  xnor csa_tree_add_6_33_groupi_g16202(csa_tree_add_6_33_groupi_n_2103 ,csa_tree_add_6_33_groupi_n_1159 ,csa_tree_add_6_33_groupi_n_1532);
  xnor csa_tree_add_6_33_groupi_g16203(csa_tree_add_6_33_groupi_n_2102 ,csa_tree_add_6_33_groupi_n_1223 ,csa_tree_add_6_33_groupi_n_1128);
  xnor csa_tree_add_6_33_groupi_g16204(csa_tree_add_6_33_groupi_n_2101 ,csa_tree_add_6_33_groupi_n_1176 ,csa_tree_add_6_33_groupi_n_1612);
  xnor csa_tree_add_6_33_groupi_g16205(csa_tree_add_6_33_groupi_n_2100 ,csa_tree_add_6_33_groupi_n_1235 ,csa_tree_add_6_33_groupi_n_1286);
  xnor csa_tree_add_6_33_groupi_g16206(csa_tree_add_6_33_groupi_n_2099 ,csa_tree_add_6_33_groupi_n_1104 ,csa_tree_add_6_33_groupi_n_1097);
  xnor csa_tree_add_6_33_groupi_g16207(csa_tree_add_6_33_groupi_n_2098 ,csa_tree_add_6_33_groupi_n_1416 ,csa_tree_add_6_33_groupi_n_1308);
  xnor csa_tree_add_6_33_groupi_g16208(csa_tree_add_6_33_groupi_n_2097 ,csa_tree_add_6_33_groupi_n_1450 ,csa_tree_add_6_33_groupi_n_1178);
  xnor csa_tree_add_6_33_groupi_g16209(csa_tree_add_6_33_groupi_n_2096 ,csa_tree_add_6_33_groupi_n_1578 ,in1[17]);
  xnor csa_tree_add_6_33_groupi_g16210(csa_tree_add_6_33_groupi_n_2095 ,csa_tree_add_6_33_groupi_n_1513 ,csa_tree_add_6_33_groupi_n_1166);
  xnor csa_tree_add_6_33_groupi_g16211(csa_tree_add_6_33_groupi_n_2094 ,csa_tree_add_6_33_groupi_n_1495 ,csa_tree_add_6_33_groupi_n_1302);
  xnor csa_tree_add_6_33_groupi_g16212(csa_tree_add_6_33_groupi_n_2093 ,csa_tree_add_6_33_groupi_n_1293 ,csa_tree_add_6_33_groupi_n_1464);
  xnor csa_tree_add_6_33_groupi_g16213(csa_tree_add_6_33_groupi_n_2092 ,csa_tree_add_6_33_groupi_n_1479 ,csa_tree_add_6_33_groupi_n_1548);
  xnor csa_tree_add_6_33_groupi_g16214(csa_tree_add_6_33_groupi_n_2091 ,csa_tree_add_6_33_groupi_n_1472 ,csa_tree_add_6_33_groupi_n_1603);
  xnor csa_tree_add_6_33_groupi_g16215(csa_tree_add_6_33_groupi_n_2090 ,csa_tree_add_6_33_groupi_n_1083 ,csa_tree_add_6_33_groupi_n_1324);
  xnor csa_tree_add_6_33_groupi_g16216(csa_tree_add_6_33_groupi_n_2089 ,csa_tree_add_6_33_groupi_n_1458 ,csa_tree_add_6_33_groupi_n_1075);
  xnor csa_tree_add_6_33_groupi_g16217(csa_tree_add_6_33_groupi_n_2088 ,csa_tree_add_6_33_groupi_n_1467 ,csa_tree_add_6_33_groupi_n_1258);
  xnor csa_tree_add_6_33_groupi_g16218(csa_tree_add_6_33_groupi_n_2087 ,csa_tree_add_6_33_groupi_n_1488 ,csa_tree_add_6_33_groupi_n_1553);
  xnor csa_tree_add_6_33_groupi_g16219(csa_tree_add_6_33_groupi_n_2086 ,csa_tree_add_6_33_groupi_n_1074 ,csa_tree_add_6_33_groupi_n_1587);
  xnor csa_tree_add_6_33_groupi_g16220(csa_tree_add_6_33_groupi_n_2085 ,csa_tree_add_6_33_groupi_n_1560 ,csa_tree_add_6_33_groupi_n_1401);
  xnor csa_tree_add_6_33_groupi_g16221(csa_tree_add_6_33_groupi_n_2084 ,csa_tree_add_6_33_groupi_n_1183 ,csa_tree_add_6_33_groupi_n_1094);
  xnor csa_tree_add_6_33_groupi_g16222(csa_tree_add_6_33_groupi_n_2083 ,csa_tree_add_6_33_groupi_n_1243 ,csa_tree_add_6_33_groupi_n_1237);
  xnor csa_tree_add_6_33_groupi_g16223(csa_tree_add_6_33_groupi_n_2082 ,csa_tree_add_6_33_groupi_n_1140 ,csa_tree_add_6_33_groupi_n_1268);
  xnor csa_tree_add_6_33_groupi_g16224(csa_tree_add_6_33_groupi_n_2081 ,csa_tree_add_6_33_groupi_n_1114 ,csa_tree_add_6_33_groupi_n_1393);
  xnor csa_tree_add_6_33_groupi_g16225(csa_tree_add_6_33_groupi_n_2080 ,csa_tree_add_6_33_groupi_n_1173 ,csa_tree_add_6_33_groupi_n_1116);
  xnor csa_tree_add_6_33_groupi_g16226(csa_tree_add_6_33_groupi_n_2079 ,csa_tree_add_6_33_groupi_n_1247 ,csa_tree_add_6_33_groupi_n_1607);
  xnor csa_tree_add_6_33_groupi_g16227(csa_tree_add_6_33_groupi_n_2078 ,csa_tree_add_6_33_groupi_n_1448 ,csa_tree_add_6_33_groupi_n_1277);
  xnor csa_tree_add_6_33_groupi_g16228(csa_tree_add_6_33_groupi_n_2077 ,csa_tree_add_6_33_groupi_n_1193 ,csa_tree_add_6_33_groupi_n_1311);
  xnor csa_tree_add_6_33_groupi_g16229(csa_tree_add_6_33_groupi_n_2076 ,csa_tree_add_6_33_groupi_n_1387 ,csa_tree_add_6_33_groupi_n_1314);
  xnor csa_tree_add_6_33_groupi_g16230(csa_tree_add_6_33_groupi_n_2075 ,csa_tree_add_6_33_groupi_n_1403 ,csa_tree_add_6_33_groupi_n_1326);
  xnor csa_tree_add_6_33_groupi_g16231(csa_tree_add_6_33_groupi_n_2074 ,csa_tree_add_6_33_groupi_n_1443 ,csa_tree_add_6_33_groupi_n_1601);
  xnor csa_tree_add_6_33_groupi_g16232(csa_tree_add_6_33_groupi_n_2073 ,csa_tree_add_6_33_groupi_n_1457 ,csa_tree_add_6_33_groupi_n_1294);
  xnor csa_tree_add_6_33_groupi_g16233(csa_tree_add_6_33_groupi_n_2072 ,csa_tree_add_6_33_groupi_n_1552 ,csa_tree_add_6_33_groupi_n_1129);
  xnor csa_tree_add_6_33_groupi_g16234(csa_tree_add_6_33_groupi_n_2071 ,csa_tree_add_6_33_groupi_n_1406 ,csa_tree_add_6_33_groupi_n_1565);
  xnor csa_tree_add_6_33_groupi_g16235(csa_tree_add_6_33_groupi_n_2070 ,csa_tree_add_6_33_groupi_n_1153 ,csa_tree_add_6_33_groupi_n_1241);
  xnor csa_tree_add_6_33_groupi_g16236(csa_tree_add_6_33_groupi_n_2069 ,csa_tree_add_6_33_groupi_n_1567 ,csa_tree_add_6_33_groupi_n_1238);
  xnor csa_tree_add_6_33_groupi_g16237(csa_tree_add_6_33_groupi_n_2068 ,csa_tree_add_6_33_groupi_n_1280 ,csa_tree_add_6_33_groupi_n_1095);
  xnor csa_tree_add_6_33_groupi_g16238(csa_tree_add_6_33_groupi_n_2067 ,csa_tree_add_6_33_groupi_n_1411 ,csa_tree_add_6_33_groupi_n_1301);
  xnor csa_tree_add_6_33_groupi_g16239(csa_tree_add_6_33_groupi_n_2066 ,csa_tree_add_6_33_groupi_n_1512 ,csa_tree_add_6_33_groupi_n_1557);
  xnor csa_tree_add_6_33_groupi_g16240(csa_tree_add_6_33_groupi_n_2065 ,csa_tree_add_6_33_groupi_n_1250 ,csa_tree_add_6_33_groupi_n_1589);
  xnor csa_tree_add_6_33_groupi_g16241(csa_tree_add_6_33_groupi_n_2064 ,csa_tree_add_6_33_groupi_n_1086 ,csa_tree_add_6_33_groupi_n_1259);
  xnor csa_tree_add_6_33_groupi_g16242(csa_tree_add_6_33_groupi_n_2063 ,csa_tree_add_6_33_groupi_n_1423 ,csa_tree_add_6_33_groupi_n_1102);
  xnor csa_tree_add_6_33_groupi_g16243(csa_tree_add_6_33_groupi_n_2062 ,csa_tree_add_6_33_groupi_n_1274 ,csa_tree_add_6_33_groupi_n_1171);
  xnor csa_tree_add_6_33_groupi_g16244(csa_tree_add_6_33_groupi_n_2061 ,csa_tree_add_6_33_groupi_n_1545 ,csa_tree_add_6_33_groupi_n_1221);
  xnor csa_tree_add_6_33_groupi_g16245(csa_tree_add_6_33_groupi_n_2060 ,csa_tree_add_6_33_groupi_n_1515 ,csa_tree_add_6_33_groupi_n_1525);
  xnor csa_tree_add_6_33_groupi_g16246(csa_tree_add_6_33_groupi_n_2059 ,csa_tree_add_6_33_groupi_n_1466 ,csa_tree_add_6_33_groupi_n_1437);
  xnor csa_tree_add_6_33_groupi_g16247(csa_tree_add_6_33_groupi_n_2058 ,csa_tree_add_6_33_groupi_n_1230 ,csa_tree_add_6_33_groupi_n_1575);
  xnor csa_tree_add_6_33_groupi_g16248(csa_tree_add_6_33_groupi_n_2057 ,csa_tree_add_6_33_groupi_n_1616 ,csa_tree_add_6_33_groupi_n_1100);
  xnor csa_tree_add_6_33_groupi_g16249(csa_tree_add_6_33_groupi_n_2056 ,csa_tree_add_6_33_groupi_n_1412 ,csa_tree_add_6_33_groupi_n_1269);
  xnor csa_tree_add_6_33_groupi_g16250(csa_tree_add_6_33_groupi_n_2055 ,csa_tree_add_6_33_groupi_n_1462 ,csa_tree_add_6_33_groupi_n_1591);
  xnor csa_tree_add_6_33_groupi_g16251(csa_tree_add_6_33_groupi_n_2054 ,csa_tree_add_6_33_groupi_n_1366 ,csa_tree_add_6_33_groupi_n_1608);
  xnor csa_tree_add_6_33_groupi_g16252(csa_tree_add_6_33_groupi_n_2053 ,csa_tree_add_6_33_groupi_n_1154 ,csa_tree_add_6_33_groupi_n_1093);
  xnor csa_tree_add_6_33_groupi_g16253(csa_tree_add_6_33_groupi_n_2052 ,csa_tree_add_6_33_groupi_n_1185 ,csa_tree_add_6_33_groupi_n_1309);
  xnor csa_tree_add_6_33_groupi_g16254(csa_tree_add_6_33_groupi_n_2051 ,csa_tree_add_6_33_groupi_n_1253 ,csa_tree_add_6_33_groupi_n_1135);
  xnor csa_tree_add_6_33_groupi_g16255(csa_tree_add_6_33_groupi_n_2050 ,csa_tree_add_6_33_groupi_n_1088 ,csa_tree_add_6_33_groupi_n_1599);
  xnor csa_tree_add_6_33_groupi_g16256(csa_tree_add_6_33_groupi_n_2049 ,csa_tree_add_6_33_groupi_n_1218 ,csa_tree_add_6_33_groupi_n_1296);
  xnor csa_tree_add_6_33_groupi_g16257(csa_tree_add_6_33_groupi_n_2048 ,csa_tree_add_6_33_groupi_n_1122 ,csa_tree_add_6_33_groupi_n_1602);
  xnor csa_tree_add_6_33_groupi_g16258(csa_tree_add_6_33_groupi_n_2047 ,csa_tree_add_6_33_groupi_n_1317 ,csa_tree_add_6_33_groupi_n_1521);
  xnor csa_tree_add_6_33_groupi_g16259(csa_tree_add_6_33_groupi_n_2046 ,csa_tree_add_6_33_groupi_n_1120 ,csa_tree_add_6_33_groupi_n_1287);
  xnor csa_tree_add_6_33_groupi_g16260(csa_tree_add_6_33_groupi_n_2045 ,csa_tree_add_6_33_groupi_n_1199 ,csa_tree_add_6_33_groupi_n_1430);
  xnor csa_tree_add_6_33_groupi_g16261(csa_tree_add_6_33_groupi_n_2044 ,csa_tree_add_6_33_groupi_n_1271 ,csa_tree_add_6_33_groupi_n_1179);
  xnor csa_tree_add_6_33_groupi_g16262(csa_tree_add_6_33_groupi_n_2043 ,csa_tree_add_6_33_groupi_n_1124 ,csa_tree_add_6_33_groupi_n_1214);
  xnor csa_tree_add_6_33_groupi_g16263(csa_tree_add_6_33_groupi_n_2042 ,csa_tree_add_6_33_groupi_n_1195 ,csa_tree_add_6_33_groupi_n_1590);
  xnor csa_tree_add_6_33_groupi_g16264(csa_tree_add_6_33_groupi_n_2041 ,csa_tree_add_6_33_groupi_n_1305 ,csa_tree_add_6_33_groupi_n_1198);
  xnor csa_tree_add_6_33_groupi_g16265(csa_tree_add_6_33_groupi_n_2040 ,csa_tree_add_6_33_groupi_n_1322 ,csa_tree_add_6_33_groupi_n_1422);
  xnor csa_tree_add_6_33_groupi_g16266(csa_tree_add_6_33_groupi_n_2039 ,csa_tree_add_6_33_groupi_n_1108 ,csa_tree_add_6_33_groupi_n_1426);
  xnor csa_tree_add_6_33_groupi_g16267(csa_tree_add_6_33_groupi_n_2038 ,csa_tree_add_6_33_groupi_n_1239 ,csa_tree_add_6_33_groupi_n_1084);
  xnor csa_tree_add_6_33_groupi_g16268(csa_tree_add_6_33_groupi_n_2037 ,csa_tree_add_6_33_groupi_n_1229 ,csa_tree_add_6_33_groupi_n_1446);
  xnor csa_tree_add_6_33_groupi_g16269(csa_tree_add_6_33_groupi_n_2036 ,csa_tree_add_6_33_groupi_n_1503 ,csa_tree_add_6_33_groupi_n_1323);
  xnor csa_tree_add_6_33_groupi_g16270(csa_tree_add_6_33_groupi_n_2035 ,csa_tree_add_6_33_groupi_n_1164 ,csa_tree_add_6_33_groupi_n_1441);
  xnor csa_tree_add_6_33_groupi_g16271(csa_tree_add_6_33_groupi_n_2034 ,csa_tree_add_6_33_groupi_n_1498 ,csa_tree_add_6_33_groupi_n_1264);
  xnor csa_tree_add_6_33_groupi_g16272(csa_tree_add_6_33_groupi_n_2033 ,csa_tree_add_6_33_groupi_n_1490 ,csa_tree_add_6_33_groupi_n_1614);
  xnor csa_tree_add_6_33_groupi_g16273(csa_tree_add_6_33_groupi_n_2032 ,csa_tree_add_6_33_groupi_n_1248 ,csa_tree_add_6_33_groupi_n_1586);
  xnor csa_tree_add_6_33_groupi_g16274(csa_tree_add_6_33_groupi_n_2031 ,csa_tree_add_6_33_groupi_n_1272 ,csa_tree_add_6_33_groupi_n_1402);
  xnor csa_tree_add_6_33_groupi_g16275(csa_tree_add_6_33_groupi_n_2030 ,csa_tree_add_6_33_groupi_n_1510 ,csa_tree_add_6_33_groupi_n_1249);
  xnor csa_tree_add_6_33_groupi_g16276(csa_tree_add_6_33_groupi_n_2029 ,csa_tree_add_6_33_groupi_n_1469 ,csa_tree_add_6_33_groupi_n_1303);
  xnor csa_tree_add_6_33_groupi_g16277(csa_tree_add_6_33_groupi_n_2028 ,csa_tree_add_6_33_groupi_n_1207 ,csa_tree_add_6_33_groupi_n_1454);
  xnor csa_tree_add_6_33_groupi_g16278(csa_tree_add_6_33_groupi_n_2027 ,csa_tree_add_6_33_groupi_n_1461 ,csa_tree_add_6_33_groupi_n_1276);
  xnor csa_tree_add_6_33_groupi_g16279(csa_tree_add_6_33_groupi_n_2026 ,csa_tree_add_6_33_groupi_n_1381 ,csa_tree_add_6_33_groupi_n_1289);
  xnor csa_tree_add_6_33_groupi_g16280(csa_tree_add_6_33_groupi_n_2025 ,csa_tree_add_6_33_groupi_n_1200 ,csa_tree_add_6_33_groupi_n_1542);
  xnor csa_tree_add_6_33_groupi_g16281(csa_tree_add_6_33_groupi_n_2024 ,csa_tree_add_6_33_groupi_n_1284 ,csa_tree_add_6_33_groupi_n_1451);
  xnor csa_tree_add_6_33_groupi_g16282(csa_tree_add_6_33_groupi_n_2023 ,csa_tree_add_6_33_groupi_n_1470 ,csa_tree_add_6_33_groupi_n_1132);
  xnor csa_tree_add_6_33_groupi_g16283(csa_tree_add_6_33_groupi_n_2022 ,csa_tree_add_6_33_groupi_n_1453 ,csa_tree_add_6_33_groupi_n_1588);
  xnor csa_tree_add_6_33_groupi_g16284(csa_tree_add_6_33_groupi_n_2021 ,csa_tree_add_6_33_groupi_n_1312 ,csa_tree_add_6_33_groupi_n_1533);
  xnor csa_tree_add_6_33_groupi_g16285(csa_tree_add_6_33_groupi_n_2020 ,csa_tree_add_6_33_groupi_n_1554 ,csa_tree_add_6_33_groupi_n_1523);
  xnor csa_tree_add_6_33_groupi_g16286(csa_tree_add_6_33_groupi_n_2019 ,csa_tree_add_6_33_groupi_n_1573 ,csa_tree_add_6_33_groupi_n_1517);
  xnor csa_tree_add_6_33_groupi_g16287(csa_tree_add_6_33_groupi_n_2018 ,csa_tree_add_6_33_groupi_n_1421 ,csa_tree_add_6_33_groupi_n_1318);
  xnor csa_tree_add_6_33_groupi_g16288(csa_tree_add_6_33_groupi_n_2017 ,csa_tree_add_6_33_groupi_n_1434 ,csa_tree_add_6_33_groupi_n_1260);
  xnor csa_tree_add_6_33_groupi_g16289(csa_tree_add_6_33_groupi_n_2016 ,csa_tree_add_6_33_groupi_n_1163 ,csa_tree_add_6_33_groupi_n_1290);
  xnor csa_tree_add_6_33_groupi_g16290(csa_tree_add_6_33_groupi_n_2015 ,csa_tree_add_6_33_groupi_n_1126 ,csa_tree_add_6_33_groupi_n_1325);
  xnor csa_tree_add_6_33_groupi_g16291(csa_tree_add_6_33_groupi_n_2014 ,csa_tree_add_6_33_groupi_n_1320 ,in1[29]);
  and csa_tree_add_6_33_groupi_g16293(csa_tree_add_6_33_groupi_n_2012 ,in2[12] ,csa_tree_add_6_33_groupi_n_1335);
  and csa_tree_add_6_33_groupi_g16294(csa_tree_add_6_33_groupi_n_2011 ,in3[4] ,csa_tree_add_6_33_groupi_n_1064);
  and csa_tree_add_6_33_groupi_g16295(csa_tree_add_6_33_groupi_n_2010 ,in2[2] ,csa_tree_add_6_33_groupi_n_1361);
  and csa_tree_add_6_33_groupi_g16296(csa_tree_add_6_33_groupi_n_2009 ,in2[24] ,csa_tree_add_6_33_groupi_n_1060);
  and csa_tree_add_6_33_groupi_g16297(csa_tree_add_6_33_groupi_n_2008 ,in2[26] ,csa_tree_add_6_33_groupi_n_1355);
  and csa_tree_add_6_33_groupi_g16298(csa_tree_add_6_33_groupi_n_2007 ,in2[10] ,csa_tree_add_6_33_groupi_n_1343);
  and csa_tree_add_6_33_groupi_g16299(csa_tree_add_6_33_groupi_n_2006 ,in2[14] ,csa_tree_add_6_33_groupi_n_1340);
  and csa_tree_add_6_33_groupi_g16300(csa_tree_add_6_33_groupi_n_2005 ,in2[28] ,csa_tree_add_6_33_groupi_n_1339);
  or csa_tree_add_6_33_groupi_g16301(csa_tree_add_6_33_groupi_n_2004 ,csa_tree_add_6_33_groupi_n_1022 ,csa_tree_add_6_33_groupi_n_1328);
  and csa_tree_add_6_33_groupi_g16302(csa_tree_add_6_33_groupi_n_2003 ,in2[22] ,csa_tree_add_6_33_groupi_n_1337);
  and csa_tree_add_6_33_groupi_g16303(csa_tree_add_6_33_groupi_n_2002 ,in2[20] ,csa_tree_add_6_33_groupi_n_1331);
  and csa_tree_add_6_33_groupi_g16304(csa_tree_add_6_33_groupi_n_2001 ,in2[30] ,csa_tree_add_6_33_groupi_n_1349);
  or csa_tree_add_6_33_groupi_g16305(csa_tree_add_6_33_groupi_n_2000 ,csa_tree_add_6_33_groupi_n_304 ,csa_tree_add_6_33_groupi_n_1125);
  and csa_tree_add_6_33_groupi_g16306(csa_tree_add_6_33_groupi_n_1999 ,csa_tree_add_6_33_groupi_n_1474 ,csa_tree_add_6_33_groupi_n_1121);
  and csa_tree_add_6_33_groupi_g16307(csa_tree_add_6_33_groupi_n_1998 ,csa_tree_add_6_33_groupi_n_1099 ,csa_tree_add_6_33_groupi_n_1189);
  or csa_tree_add_6_33_groupi_g16308(csa_tree_add_6_33_groupi_n_1997 ,csa_tree_add_6_33_groupi_n_1498 ,csa_tree_add_6_33_groupi_n_1082);
  or csa_tree_add_6_33_groupi_g16309(csa_tree_add_6_33_groupi_n_1996 ,csa_tree_add_6_33_groupi_n_1438 ,csa_tree_add_6_33_groupi_n_1083);
  or csa_tree_add_6_33_groupi_g16310(csa_tree_add_6_33_groupi_n_1995 ,csa_tree_add_6_33_groupi_n_1233 ,csa_tree_add_6_33_groupi_n_1452);
  or csa_tree_add_6_33_groupi_g16311(csa_tree_add_6_33_groupi_n_1994 ,csa_tree_add_6_33_groupi_n_1114 ,csa_tree_add_6_33_groupi_n_1393);
  or csa_tree_add_6_33_groupi_g16312(csa_tree_add_6_33_groupi_n_1993 ,csa_tree_add_6_33_groupi_n_1499 ,csa_tree_add_6_33_groupi_n_1379);
  or csa_tree_add_6_33_groupi_g16313(csa_tree_add_6_33_groupi_n_1992 ,csa_tree_add_6_33_groupi_n_1130 ,csa_tree_add_6_33_groupi_n_1390);
  or csa_tree_add_6_33_groupi_g16315(csa_tree_add_6_33_groupi_n_1990 ,csa_tree_add_6_33_groupi_n_1478 ,csa_tree_add_6_33_groupi_n_1521);
  and csa_tree_add_6_33_groupi_g16316(csa_tree_add_6_33_groupi_n_1989 ,csa_tree_add_6_33_groupi_n_1227 ,csa_tree_add_6_33_groupi_n_1171);
  and csa_tree_add_6_33_groupi_g16317(csa_tree_add_6_33_groupi_n_1988 ,csa_tree_add_6_33_groupi_n_1432 ,csa_tree_add_6_33_groupi_n_1148);
  and csa_tree_add_6_33_groupi_g16318(csa_tree_add_6_33_groupi_n_1987 ,csa_tree_add_6_33_groupi_n_1095 ,csa_tree_add_6_33_groupi_n_1501);
  or csa_tree_add_6_33_groupi_g16319(csa_tree_add_6_33_groupi_n_1986 ,csa_tree_add_6_33_groupi_n_1517 ,csa_tree_add_6_33_groupi_n_1244);
  and csa_tree_add_6_33_groupi_g16320(csa_tree_add_6_33_groupi_n_1985 ,csa_tree_add_6_33_groupi_n_1198 ,csa_tree_add_6_33_groupi_n_1447);
  or csa_tree_add_6_33_groupi_g16321(csa_tree_add_6_33_groupi_n_1984 ,csa_tree_add_6_33_groupi_n_1230 ,csa_tree_add_6_33_groupi_n_1485);
  and csa_tree_add_6_33_groupi_g16322(csa_tree_add_6_33_groupi_n_1983 ,csa_tree_add_6_33_groupi_n_1079 ,csa_tree_add_6_33_groupi_n_1092);
  and csa_tree_add_6_33_groupi_g16323(csa_tree_add_6_33_groupi_n_1982 ,csa_tree_add_6_33_groupi_n_1130 ,csa_tree_add_6_33_groupi_n_1390);
  and csa_tree_add_6_33_groupi_g16324(csa_tree_add_6_33_groupi_n_1981 ,csa_tree_add_6_33_groupi_n_1472 ,csa_tree_add_6_33_groupi_n_1197);
  or csa_tree_add_6_33_groupi_g16325(csa_tree_add_6_33_groupi_n_1980 ,csa_tree_add_6_33_groupi_n_427 ,csa_tree_add_6_33_groupi_n_1136);
  or csa_tree_add_6_33_groupi_g16326(csa_tree_add_6_33_groupi_n_1979 ,csa_tree_add_6_33_groupi_n_1088 ,csa_tree_add_6_33_groupi_n_1090);
  and csa_tree_add_6_33_groupi_g16327(csa_tree_add_6_33_groupi_n_1978 ,csa_tree_add_6_33_groupi_n_1135 ,csa_tree_add_6_33_groupi_n_1155);
  or csa_tree_add_6_33_groupi_g16329(csa_tree_add_6_33_groupi_n_1976 ,csa_tree_add_6_33_groupi_n_1513 ,csa_tree_add_6_33_groupi_n_1166);
  and csa_tree_add_6_33_groupi_g16330(csa_tree_add_6_33_groupi_n_1975 ,csa_tree_add_6_33_groupi_n_1191 ,csa_tree_add_6_33_groupi_n_1418);
  or csa_tree_add_6_33_groupi_g16332(csa_tree_add_6_33_groupi_n_1973 ,csa_tree_add_6_33_groupi_n_1434 ,csa_tree_add_6_33_groupi_n_1435);
  or csa_tree_add_6_33_groupi_g16333(csa_tree_add_6_33_groupi_n_1972 ,csa_tree_add_6_33_groupi_n_1526 ,csa_tree_add_6_33_groupi_n_1514);
  and csa_tree_add_6_33_groupi_g16334(csa_tree_add_6_33_groupi_n_1971 ,csa_tree_add_6_33_groupi_n_1074 ,csa_tree_add_6_33_groupi_n_1170);
  and csa_tree_add_6_33_groupi_g16335(csa_tree_add_6_33_groupi_n_1970 ,csa_tree_add_6_33_groupi_n_1493 ,csa_tree_add_6_33_groupi_n_1158);
  and csa_tree_add_6_33_groupi_g16336(csa_tree_add_6_33_groupi_n_1969 ,csa_tree_add_6_33_groupi_n_1096 ,csa_tree_add_6_33_groupi_n_1217);
  or csa_tree_add_6_33_groupi_g16337(csa_tree_add_6_33_groupi_n_1968 ,csa_tree_add_6_33_groupi_n_1149 ,csa_tree_add_6_33_groupi_n_1394);
  or csa_tree_add_6_33_groupi_g16338(csa_tree_add_6_33_groupi_n_1967 ,csa_tree_add_6_33_groupi_n_478 ,csa_tree_add_6_33_groupi_n_1494);
  or csa_tree_add_6_33_groupi_g16339(csa_tree_add_6_33_groupi_n_1966 ,csa_tree_add_6_33_groupi_n_1191 ,csa_tree_add_6_33_groupi_n_1418);
  or csa_tree_add_6_33_groupi_g16340(csa_tree_add_6_33_groupi_n_1965 ,csa_tree_add_6_33_groupi_n_1119 ,csa_tree_add_6_33_groupi_n_1226);
  and csa_tree_add_6_33_groupi_g16341(csa_tree_add_6_33_groupi_n_1964 ,csa_tree_add_6_33_groupi_n_1513 ,csa_tree_add_6_33_groupi_n_1166);
  nor csa_tree_add_6_33_groupi_g16342(csa_tree_add_6_33_groupi_n_1963 ,csa_tree_add_6_33_groupi_n_1593 ,csa_tree_add_6_33_groupi_n_1061);
  or csa_tree_add_6_33_groupi_g16343(csa_tree_add_6_33_groupi_n_1962 ,csa_tree_add_6_33_groupi_n_1203 ,csa_tree_add_6_33_groupi_n_1141);
  or csa_tree_add_6_33_groupi_g16344(csa_tree_add_6_33_groupi_n_1961 ,csa_tree_add_6_33_groupi_n_1381 ,csa_tree_add_6_33_groupi_n_1118);
  and csa_tree_add_6_33_groupi_g16345(csa_tree_add_6_33_groupi_n_1960 ,csa_tree_add_6_33_groupi_n_1499 ,csa_tree_add_6_33_groupi_n_1379);
  or csa_tree_add_6_33_groupi_g16346(csa_tree_add_6_33_groupi_n_1959 ,csa_tree_add_6_33_groupi_n_1135 ,csa_tree_add_6_33_groupi_n_1155);
  or csa_tree_add_6_33_groupi_g16347(csa_tree_add_6_33_groupi_n_1958 ,csa_tree_add_6_33_groupi_n_1183 ,csa_tree_add_6_33_groupi_n_1094);
  or csa_tree_add_6_33_groupi_g16349(csa_tree_add_6_33_groupi_n_1956 ,csa_tree_add_6_33_groupi_n_1215 ,csa_tree_add_6_33_groupi_n_1179);
  nor csa_tree_add_6_33_groupi_g16350(csa_tree_add_6_33_groupi_n_1955 ,csa_tree_add_6_33_groupi_n_1563 ,csa_tree_add_6_33_groupi_n_1345);
  and csa_tree_add_6_33_groupi_g16351(csa_tree_add_6_33_groupi_n_1954 ,csa_tree_add_6_33_groupi_n_1520 ,csa_tree_add_6_33_groupi_n_1511);
  nor csa_tree_add_6_33_groupi_g16352(csa_tree_add_6_33_groupi_n_1953 ,csa_tree_add_6_33_groupi_n_1161 ,csa_tree_add_6_33_groupi_n_1477);
  and csa_tree_add_6_33_groupi_g16353(csa_tree_add_6_33_groupi_n_1952 ,csa_tree_add_6_33_groupi_n_1215 ,csa_tree_add_6_33_groupi_n_1179);
  and csa_tree_add_6_33_groupi_g16354(csa_tree_add_6_33_groupi_n_1951 ,csa_tree_add_6_33_groupi_n_1149 ,csa_tree_add_6_33_groupi_n_1394);
  nor csa_tree_add_6_33_groupi_g16355(csa_tree_add_6_33_groupi_n_1950 ,csa_tree_add_6_33_groupi_n_1543 ,csa_tree_add_6_33_groupi_n_1332);
  and csa_tree_add_6_33_groupi_g16356(csa_tree_add_6_33_groupi_n_1949 ,csa_tree_add_6_33_groupi_n_1504 ,csa_tree_add_6_33_groupi_n_1436);
  and csa_tree_add_6_33_groupi_g16357(csa_tree_add_6_33_groupi_n_1948 ,csa_tree_add_6_33_groupi_n_1243 ,csa_tree_add_6_33_groupi_n_1237);
  and csa_tree_add_6_33_groupi_g16358(csa_tree_add_6_33_groupi_n_1947 ,csa_tree_add_6_33_groupi_n_1526 ,csa_tree_add_6_33_groupi_n_1514);
  or csa_tree_add_6_33_groupi_g16359(csa_tree_add_6_33_groupi_n_1946 ,csa_tree_add_6_33_groupi_n_1295 ,csa_tree_add_6_33_groupi_n_1351);
  and csa_tree_add_6_33_groupi_g16360(csa_tree_add_6_33_groupi_n_1945 ,csa_tree_add_6_33_groupi_n_1488 ,csa_tree_add_6_33_groupi_n_1162);
  and csa_tree_add_6_33_groupi_g16361(csa_tree_add_6_33_groupi_n_1944 ,csa_tree_add_6_33_groupi_n_1530 ,csa_tree_add_6_33_groupi_n_1374);
  and csa_tree_add_6_33_groupi_g16362(csa_tree_add_6_33_groupi_n_1943 ,csa_tree_add_6_33_groupi_n_1455 ,csa_tree_add_6_33_groupi_n_1167);
  or csa_tree_add_6_33_groupi_g16363(csa_tree_add_6_33_groupi_n_1942 ,csa_tree_add_6_33_groupi_n_1486 ,csa_tree_add_6_33_groupi_n_1205);
  and csa_tree_add_6_33_groupi_g16364(csa_tree_add_6_33_groupi_n_1941 ,csa_tree_add_6_33_groupi_n_1104 ,csa_tree_add_6_33_groupi_n_1097);
  or csa_tree_add_6_33_groupi_g16366(csa_tree_add_6_33_groupi_n_1939 ,csa_tree_add_6_33_groupi_n_1455 ,csa_tree_add_6_33_groupi_n_1167);
  or csa_tree_add_6_33_groupi_g16367(csa_tree_add_6_33_groupi_n_1938 ,csa_tree_add_6_33_groupi_n_1087 ,csa_tree_add_6_33_groupi_n_1151);
  or csa_tree_add_6_33_groupi_g16368(csa_tree_add_6_33_groupi_n_1937 ,csa_tree_add_6_33_groupi_n_1089 ,csa_tree_add_6_33_groupi_n_1117);
  or csa_tree_add_6_33_groupi_g16369(csa_tree_add_6_33_groupi_n_1936 ,csa_tree_add_6_33_groupi_n_1427 ,csa_tree_add_6_33_groupi_n_1127);
  and csa_tree_add_6_33_groupi_g16370(csa_tree_add_6_33_groupi_n_1935 ,csa_tree_add_6_33_groupi_n_1088 ,csa_tree_add_6_33_groupi_n_1090);
  and csa_tree_add_6_33_groupi_g16371(csa_tree_add_6_33_groupi_n_1934 ,csa_tree_add_6_33_groupi_n_1517 ,csa_tree_add_6_33_groupi_n_1244);
  or csa_tree_add_6_33_groupi_g16372(csa_tree_add_6_33_groupi_n_1933 ,csa_tree_add_6_33_groupi_n_1316 ,csa_tree_add_6_33_groupi_n_1043);
  and csa_tree_add_6_33_groupi_g16373(csa_tree_add_6_33_groupi_n_1932 ,csa_tree_add_6_33_groupi_n_1458 ,csa_tree_add_6_33_groupi_n_1075);
  and csa_tree_add_6_33_groupi_g16374(csa_tree_add_6_33_groupi_n_1931 ,csa_tree_add_6_33_groupi_n_1487 ,csa_tree_add_6_33_groupi_n_1411);
  or csa_tree_add_6_33_groupi_g16375(csa_tree_add_6_33_groupi_n_1930 ,csa_tree_add_6_33_groupi_n_1520 ,csa_tree_add_6_33_groupi_n_1511);
  and csa_tree_add_6_33_groupi_g16376(csa_tree_add_6_33_groupi_n_1929 ,csa_tree_add_6_33_groupi_n_1529 ,csa_tree_add_6_33_groupi_n_1204);
  or csa_tree_add_6_33_groupi_g16377(csa_tree_add_6_33_groupi_n_1928 ,csa_tree_add_6_33_groupi_n_1188 ,csa_tree_add_6_33_groupi_n_1402);
  or csa_tree_add_6_33_groupi_g16378(csa_tree_add_6_33_groupi_n_1927 ,csa_tree_add_6_33_groupi_n_782 ,csa_tree_add_6_33_groupi_n_1177);
  nor csa_tree_add_6_33_groupi_g16379(csa_tree_add_6_33_groupi_n_1926 ,csa_tree_add_6_33_groupi_n_1251 ,csa_tree_add_6_33_groupi_n_1346);
  or csa_tree_add_6_33_groupi_g16380(csa_tree_add_6_33_groupi_n_1925 ,csa_tree_add_6_33_groupi_n_1422 ,csa_tree_add_6_33_groupi_n_1212);
  and csa_tree_add_6_33_groupi_g16381(csa_tree_add_6_33_groupi_n_1924 ,csa_tree_add_6_33_groupi_n_1510 ,csa_tree_add_6_33_groupi_n_1249);
  and csa_tree_add_6_33_groupi_g16382(csa_tree_add_6_33_groupi_n_1923 ,csa_tree_add_6_33_groupi_n_1456 ,csa_tree_add_6_33_groupi_n_1451);
  or csa_tree_add_6_33_groupi_g16383(csa_tree_add_6_33_groupi_n_1922 ,csa_tree_add_6_33_groupi_n_1482 ,csa_tree_add_6_33_groupi_n_1169);
  or csa_tree_add_6_33_groupi_g16385(csa_tree_add_6_33_groupi_n_1920 ,csa_tree_add_6_33_groupi_n_1510 ,csa_tree_add_6_33_groupi_n_1249);
  and csa_tree_add_6_33_groupi_g16386(csa_tree_add_6_33_groupi_n_1919 ,csa_tree_add_6_33_groupi_n_1515 ,csa_tree_add_6_33_groupi_n_1525);
  nor csa_tree_add_6_33_groupi_g16387(csa_tree_add_6_33_groupi_n_1918 ,csa_tree_add_6_33_groupi_n_128 ,csa_tree_add_6_33_groupi_n_1348);
  or csa_tree_add_6_33_groupi_g16388(csa_tree_add_6_33_groupi_n_1917 ,csa_tree_add_6_33_groupi_n_1531 ,csa_tree_add_6_33_groupi_n_1489);
  or csa_tree_add_6_33_groupi_g16389(csa_tree_add_6_33_groupi_n_1916 ,csa_tree_add_6_33_groupi_n_1530 ,csa_tree_add_6_33_groupi_n_1374);
  and csa_tree_add_6_33_groupi_g16390(csa_tree_add_6_33_groupi_n_1915 ,in2[18] ,csa_tree_add_6_33_groupi_n_1055);
  or csa_tree_add_6_33_groupi_g16391(csa_tree_add_6_33_groupi_n_1914 ,csa_tree_add_6_33_groupi_n_271 ,csa_tree_add_6_33_groupi_n_1152);
  and csa_tree_add_6_33_groupi_g16392(csa_tree_add_6_33_groupi_n_1913 ,csa_tree_add_6_33_groupi_n_1366 ,csa_tree_add_6_33_groupi_n_1070);
  or csa_tree_add_6_33_groupi_g16393(csa_tree_add_6_33_groupi_n_1912 ,csa_tree_add_6_33_groupi_n_1124 ,csa_tree_add_6_33_groupi_n_1214);
  and csa_tree_add_6_33_groupi_g16394(csa_tree_add_6_33_groupi_n_1911 ,csa_tree_add_6_33_groupi_n_1156 ,csa_tree_add_6_33_groupi_n_1462);
  and csa_tree_add_6_33_groupi_g16395(csa_tree_add_6_33_groupi_n_1910 ,csa_tree_add_6_33_groupi_n_1238 ,csa_tree_add_6_33_groupi_n_1115);
  and csa_tree_add_6_33_groupi_g16396(csa_tree_add_6_33_groupi_n_1909 ,csa_tree_add_6_33_groupi_n_1126 ,csa_tree_add_6_33_groupi_n_1240);
  or csa_tree_add_6_33_groupi_g16397(csa_tree_add_6_33_groupi_n_1908 ,csa_tree_add_6_33_groupi_n_1218 ,csa_tree_add_6_33_groupi_n_1395);
  or csa_tree_add_6_33_groupi_g16398(csa_tree_add_6_33_groupi_n_1907 ,csa_tree_add_6_33_groupi_n_1433 ,csa_tree_add_6_33_groupi_n_1412);
  or csa_tree_add_6_33_groupi_g16399(csa_tree_add_6_33_groupi_n_1906 ,csa_tree_add_6_33_groupi_n_1523 ,csa_tree_add_6_33_groupi_n_1228);
  or csa_tree_add_6_33_groupi_g16400(csa_tree_add_6_33_groupi_n_1905 ,csa_tree_add_6_33_groupi_n_1173 ,csa_tree_add_6_33_groupi_n_1116);
  or csa_tree_add_6_33_groupi_g16401(csa_tree_add_6_33_groupi_n_1904 ,csa_tree_add_6_33_groupi_n_1076 ,csa_tree_add_6_33_groupi_n_1401);
  and csa_tree_add_6_33_groupi_g16402(csa_tree_add_6_33_groupi_n_1903 ,csa_tree_add_6_33_groupi_n_1533 ,csa_tree_add_6_33_groupi_n_1103);
  or csa_tree_add_6_33_groupi_g16403(csa_tree_add_6_33_groupi_n_1902 ,csa_tree_add_6_33_groupi_n_1199 ,csa_tree_add_6_33_groupi_n_1430);
  and csa_tree_add_6_33_groupi_g16404(csa_tree_add_6_33_groupi_n_1901 ,csa_tree_add_6_33_groupi_n_1531 ,csa_tree_add_6_33_groupi_n_1489);
  or csa_tree_add_6_33_groupi_g16405(csa_tree_add_6_33_groupi_n_1900 ,csa_tree_add_6_33_groupi_n_1479 ,csa_tree_add_6_33_groupi_n_1364);
  and csa_tree_add_6_33_groupi_g16406(csa_tree_add_6_33_groupi_n_1899 ,csa_tree_add_6_33_groupi_n_1168 ,csa_tree_add_6_33_groupi_n_1242);
  and csa_tree_add_6_33_groupi_g16407(csa_tree_add_6_33_groupi_n_1898 ,csa_tree_add_6_33_groupi_n_1433 ,csa_tree_add_6_33_groupi_n_1412);
  or csa_tree_add_6_33_groupi_g16408(csa_tree_add_6_33_groupi_n_1897 ,csa_tree_add_6_33_groupi_n_1504 ,csa_tree_add_6_33_groupi_n_1436);
  or csa_tree_add_6_33_groupi_g16409(csa_tree_add_6_33_groupi_n_1896 ,csa_tree_add_6_33_groupi_n_1533 ,csa_tree_add_6_33_groupi_n_1103);
  or csa_tree_add_6_33_groupi_g16411(csa_tree_add_6_33_groupi_n_1894 ,csa_tree_add_6_33_groupi_n_1457 ,csa_tree_add_6_33_groupi_n_1194);
  or csa_tree_add_6_33_groupi_g16412(csa_tree_add_6_33_groupi_n_1893 ,csa_tree_add_6_33_groupi_n_1529 ,csa_tree_add_6_33_groupi_n_1204);
  and csa_tree_add_6_33_groupi_g16413(csa_tree_add_6_33_groupi_n_1892 ,csa_tree_add_6_33_groupi_n_1450 ,csa_tree_add_6_33_groupi_n_1178);
  or csa_tree_add_6_33_groupi_g16414(csa_tree_add_6_33_groupi_n_1891 ,csa_tree_add_6_33_groupi_n_1470 ,csa_tree_add_6_33_groupi_n_1132);
  or csa_tree_add_6_33_groupi_g16415(csa_tree_add_6_33_groupi_n_1890 ,csa_tree_add_6_33_groupi_n_1459 ,csa_tree_add_6_33_groupi_n_1392);
  nor csa_tree_add_6_33_groupi_g16416(csa_tree_add_6_33_groupi_n_1889 ,csa_tree_add_6_33_groupi_n_1570 ,csa_tree_add_6_33_groupi_n_1333);
  and csa_tree_add_6_33_groupi_g16417(csa_tree_add_6_33_groupi_n_1888 ,csa_tree_add_6_33_groupi_n_1139 ,csa_tree_add_6_33_groupi_n_1439);
  or csa_tree_add_6_33_groupi_g16418(csa_tree_add_6_33_groupi_n_1887 ,csa_tree_add_6_33_groupi_n_1172 ,csa_tree_add_6_33_groupi_n_1182);
  or csa_tree_add_6_33_groupi_g16419(csa_tree_add_6_33_groupi_n_1886 ,csa_tree_add_6_33_groupi_n_1505 ,csa_tree_add_6_33_groupi_n_1163);
  nor csa_tree_add_6_33_groupi_g16420(csa_tree_add_6_33_groupi_n_1885 ,csa_tree_add_6_33_groupi_n_1425 ,csa_tree_add_6_33_groupi_n_1535);
  or csa_tree_add_6_33_groupi_g16421(csa_tree_add_6_33_groupi_n_1884 ,csa_tree_add_6_33_groupi_n_1262 ,csa_tree_add_6_33_groupi_n_1334);
  and csa_tree_add_6_33_groupi_g16422(csa_tree_add_6_33_groupi_n_1883 ,csa_tree_add_6_33_groupi_n_770 ,csa_tree_add_6_33_groupi_n_1245);
  and csa_tree_add_6_33_groupi_g16423(csa_tree_add_6_33_groupi_n_1882 ,csa_tree_add_6_33_groupi_n_1153 ,csa_tree_add_6_33_groupi_n_1241);
  and csa_tree_add_6_33_groupi_g16424(csa_tree_add_6_33_groupi_n_1881 ,csa_tree_add_6_33_groupi_n_1222 ,csa_tree_add_6_33_groupi_n_1386);
  and csa_tree_add_6_33_groupi_g16425(csa_tree_add_6_33_groupi_n_1880 ,csa_tree_add_6_33_groupi_n_1114 ,csa_tree_add_6_33_groupi_n_1393);
  or csa_tree_add_6_33_groupi_g16426(csa_tree_add_6_33_groupi_n_1879 ,csa_tree_add_6_33_groupi_n_1465 ,csa_tree_add_6_33_groupi_n_1144);
  and csa_tree_add_6_33_groupi_g16427(csa_tree_add_6_33_groupi_n_1878 ,csa_tree_add_6_33_groupi_n_1183 ,csa_tree_add_6_33_groupi_n_1094);
  or csa_tree_add_6_33_groupi_g16428(csa_tree_add_6_33_groupi_n_1877 ,csa_tree_add_6_33_groupi_n_1222 ,csa_tree_add_6_33_groupi_n_1386);
  and csa_tree_add_6_33_groupi_g16429(csa_tree_add_6_33_groupi_n_1876 ,csa_tree_add_6_33_groupi_n_1387 ,csa_tree_add_6_33_groupi_n_1377);
  and csa_tree_add_6_33_groupi_g16430(csa_tree_add_6_33_groupi_n_1875 ,csa_tree_add_6_33_groupi_n_1419 ,csa_tree_add_6_33_groupi_n_1416);
  or csa_tree_add_6_33_groupi_g16431(csa_tree_add_6_33_groupi_n_1874 ,csa_tree_add_6_33_groupi_n_1429 ,csa_tree_add_6_33_groupi_n_1398);
  or csa_tree_add_6_33_groupi_g16432(csa_tree_add_6_33_groupi_n_1873 ,csa_tree_add_6_33_groupi_n_1238 ,csa_tree_add_6_33_groupi_n_1115);
  or csa_tree_add_6_33_groupi_g16433(csa_tree_add_6_33_groupi_n_1872 ,csa_tree_add_6_33_groupi_n_1079 ,csa_tree_add_6_33_groupi_n_1092);
  and csa_tree_add_6_33_groupi_g16434(csa_tree_add_6_33_groupi_n_1871 ,csa_tree_add_6_33_groupi_n_1101 ,csa_tree_add_6_33_groupi_n_1208);
  or csa_tree_add_6_33_groupi_g16435(csa_tree_add_6_33_groupi_n_1870 ,csa_tree_add_6_33_groupi_n_1445 ,csa_tree_add_6_33_groupi_n_1200);
  and csa_tree_add_6_33_groupi_g16436(csa_tree_add_6_33_groupi_n_1869 ,csa_tree_add_6_33_groupi_n_1457 ,csa_tree_add_6_33_groupi_n_1194);
  or csa_tree_add_6_33_groupi_g16437(csa_tree_add_6_33_groupi_n_1868 ,csa_tree_add_6_33_groupi_n_1566 ,csa_tree_add_6_33_groupi_n_1057);
  or csa_tree_add_6_33_groupi_g16438(csa_tree_add_6_33_groupi_n_1867 ,csa_tree_add_6_33_groupi_n_1074 ,csa_tree_add_6_33_groupi_n_1170);
  and csa_tree_add_6_33_groupi_g16439(csa_tree_add_6_33_groupi_n_1866 ,csa_tree_add_6_33_groupi_n_1482 ,csa_tree_add_6_33_groupi_n_1169);
  and csa_tree_add_6_33_groupi_g16441(csa_tree_add_6_33_groupi_n_1864 ,csa_tree_add_6_33_groupi_n_1371 ,csa_tree_add_6_33_groupi_n_1449);
  or csa_tree_add_6_33_groupi_g16442(csa_tree_add_6_33_groupi_n_1863 ,csa_tree_add_6_33_groupi_n_1387 ,csa_tree_add_6_33_groupi_n_1377);
  and csa_tree_add_6_33_groupi_g16443(csa_tree_add_6_33_groupi_n_1862 ,csa_tree_add_6_33_groupi_n_334 ,csa_tree_add_6_33_groupi_n_1440);
  and csa_tree_add_6_33_groupi_g16444(csa_tree_add_6_33_groupi_n_1861 ,csa_tree_add_6_33_groupi_n_1232 ,csa_tree_add_6_33_groupi_n_1216);
  or csa_tree_add_6_33_groupi_g16445(csa_tree_add_6_33_groupi_n_1860 ,csa_tree_add_6_33_groupi_n_1085 ,csa_tree_add_6_33_groupi_n_1105);
  or csa_tree_add_6_33_groupi_g16446(csa_tree_add_6_33_groupi_n_1859 ,csa_tree_add_6_33_groupi_n_1202 ,csa_tree_add_6_33_groupi_n_1367);
  and csa_tree_add_6_33_groupi_g16447(csa_tree_add_6_33_groupi_n_1858 ,csa_tree_add_6_33_groupi_n_1415 ,csa_tree_add_6_33_groupi_n_1467);
  and csa_tree_add_6_33_groupi_g16448(csa_tree_add_6_33_groupi_n_1857 ,csa_tree_add_6_33_groupi_n_1181 ,csa_tree_add_6_33_groupi_n_1463);
  and csa_tree_add_6_33_groupi_g16449(csa_tree_add_6_33_groupi_n_1856 ,csa_tree_add_6_33_groupi_n_1445 ,csa_tree_add_6_33_groupi_n_1200);
  or csa_tree_add_6_33_groupi_g16450(csa_tree_add_6_33_groupi_n_1855 ,csa_tree_add_6_33_groupi_n_1168 ,csa_tree_add_6_33_groupi_n_1242);
  and csa_tree_add_6_33_groupi_g16451(csa_tree_add_6_33_groupi_n_1854 ,csa_tree_add_6_33_groupi_n_1248 ,csa_tree_add_6_33_groupi_n_1444);
  or csa_tree_add_6_33_groupi_g16452(csa_tree_add_6_33_groupi_n_1853 ,csa_tree_add_6_33_groupi_n_598 ,csa_tree_add_6_33_groupi_n_1524);
  or csa_tree_add_6_33_groupi_g16453(csa_tree_add_6_33_groupi_n_1852 ,csa_tree_add_6_33_groupi_n_1198 ,csa_tree_add_6_33_groupi_n_1447);
  and csa_tree_add_6_33_groupi_g16454(csa_tree_add_6_33_groupi_n_1851 ,csa_tree_add_6_33_groupi_n_1492 ,csa_tree_add_6_33_groupi_n_1165);
  or csa_tree_add_6_33_groupi_g16455(csa_tree_add_6_33_groupi_n_1850 ,csa_tree_add_6_33_groupi_n_1515 ,csa_tree_add_6_33_groupi_n_1525);
  or csa_tree_add_6_33_groupi_g16456(csa_tree_add_6_33_groupi_n_1849 ,csa_tree_add_6_33_groupi_n_1101 ,csa_tree_add_6_33_groupi_n_1208);
  or csa_tree_add_6_33_groupi_g16457(csa_tree_add_6_33_groupi_n_1848 ,csa_tree_add_6_33_groupi_n_1239 ,csa_tree_add_6_33_groupi_n_1084);
  or csa_tree_add_6_33_groupi_g16458(csa_tree_add_6_33_groupi_n_1847 ,csa_tree_add_6_33_groupi_n_1480 ,csa_tree_add_6_33_groupi_n_1443);
  or csa_tree_add_6_33_groupi_g16459(csa_tree_add_6_33_groupi_n_1846 ,csa_tree_add_6_33_groupi_n_1248 ,csa_tree_add_6_33_groupi_n_1444);
  and csa_tree_add_6_33_groupi_g16460(csa_tree_add_6_33_groupi_n_1845 ,csa_tree_add_6_33_groupi_n_1465 ,csa_tree_add_6_33_groupi_n_1144);
  or csa_tree_add_6_33_groupi_g16461(csa_tree_add_6_33_groupi_n_1844 ,csa_tree_add_6_33_groupi_n_1366 ,csa_tree_add_6_33_groupi_n_1070);
  and csa_tree_add_6_33_groupi_g16462(csa_tree_add_6_33_groupi_n_1843 ,csa_tree_add_6_33_groupi_n_1233 ,csa_tree_add_6_33_groupi_n_1452);
  or csa_tree_add_6_33_groupi_g16463(csa_tree_add_6_33_groupi_n_1842 ,csa_tree_add_6_33_groupi_n_794 ,csa_tree_add_6_33_groupi_n_1391);
  and csa_tree_add_6_33_groupi_g16464(csa_tree_add_6_33_groupi_n_1841 ,csa_tree_add_6_33_groupi_n_1528 ,csa_tree_add_6_33_groupi_n_1185);
  and csa_tree_add_6_33_groupi_g16465(csa_tree_add_6_33_groupi_n_1840 ,csa_tree_add_6_33_groupi_n_1230 ,csa_tree_add_6_33_groupi_n_1485);
  or csa_tree_add_6_33_groupi_g16466(csa_tree_add_6_33_groupi_n_1839 ,csa_tree_add_6_33_groupi_n_1528 ,csa_tree_add_6_33_groupi_n_1185);
  or csa_tree_add_6_33_groupi_g16467(csa_tree_add_6_33_groupi_n_1838 ,csa_tree_add_6_33_groupi_n_1450 ,csa_tree_add_6_33_groupi_n_1178);
  and csa_tree_add_6_33_groupi_g16468(csa_tree_add_6_33_groupi_n_1837 ,csa_tree_add_6_33_groupi_n_1188 ,csa_tree_add_6_33_groupi_n_1402);
  and csa_tree_add_6_33_groupi_g16469(csa_tree_add_6_33_groupi_n_1836 ,csa_tree_add_6_33_groupi_n_736 ,csa_tree_add_6_33_groupi_n_1131);
  or csa_tree_add_6_33_groupi_g16470(csa_tree_add_6_33_groupi_n_1835 ,csa_tree_add_6_33_groupi_n_1207 ,csa_tree_add_6_33_groupi_n_1454);
  or csa_tree_add_6_33_groupi_g16471(csa_tree_add_6_33_groupi_n_1834 ,csa_tree_add_6_33_groupi_n_1122 ,csa_tree_add_6_33_groupi_n_1211);
  and csa_tree_add_6_33_groupi_g16472(csa_tree_add_6_33_groupi_n_1833 ,csa_tree_add_6_33_groupi_n_1459 ,csa_tree_add_6_33_groupi_n_1392);
  and csa_tree_add_6_33_groupi_g16473(csa_tree_add_6_33_groupi_n_1832 ,csa_tree_add_6_33_groupi_n_1207 ,csa_tree_add_6_33_groupi_n_1454);
  and csa_tree_add_6_33_groupi_g16474(csa_tree_add_6_33_groupi_n_1831 ,csa_tree_add_6_33_groupi_n_1073 ,csa_tree_add_6_33_groupi_n_1110);
  or csa_tree_add_6_33_groupi_g16475(csa_tree_add_6_33_groupi_n_1830 ,csa_tree_add_6_33_groupi_n_1458 ,csa_tree_add_6_33_groupi_n_1075);
  or csa_tree_add_6_33_groupi_g16476(csa_tree_add_6_33_groupi_n_1829 ,csa_tree_add_6_33_groupi_n_1247 ,csa_tree_add_6_33_groupi_n_1201);
  or csa_tree_add_6_33_groupi_g16477(csa_tree_add_6_33_groupi_n_1828 ,csa_tree_add_6_33_groupi_n_1190 ,csa_tree_add_6_33_groupi_n_1403);
  and csa_tree_add_6_33_groupi_g16478(csa_tree_add_6_33_groupi_n_1827 ,csa_tree_add_6_33_groupi_n_1495 ,csa_tree_add_6_33_groupi_n_1500);
  or csa_tree_add_6_33_groupi_g16479(csa_tree_add_6_33_groupi_n_1826 ,csa_tree_add_6_33_groupi_n_1512 ,csa_tree_add_6_33_groupi_n_1405);
  and csa_tree_add_6_33_groupi_g16480(csa_tree_add_6_33_groupi_n_1825 ,csa_tree_add_6_33_groupi_n_1231 ,csa_tree_add_6_33_groupi_n_1120);
  or csa_tree_add_6_33_groupi_g16481(csa_tree_add_6_33_groupi_n_1824 ,csa_tree_add_6_33_groupi_n_1227 ,csa_tree_add_6_33_groupi_n_1171);
  and csa_tree_add_6_33_groupi_g16482(csa_tree_add_6_33_groupi_n_1823 ,csa_tree_add_6_33_groupi_n_1146 ,csa_tree_add_6_33_groupi_n_1491);
  or csa_tree_add_6_33_groupi_g16483(csa_tree_add_6_33_groupi_n_1822 ,csa_tree_add_6_33_groupi_n_1368 ,csa_tree_add_6_33_groupi_n_1100);
  and csa_tree_add_6_33_groupi_g16484(csa_tree_add_6_33_groupi_n_1821 ,csa_tree_add_6_33_groupi_n_1176 ,csa_tree_add_6_33_groupi_n_1123);
  or csa_tree_add_6_33_groupi_g16485(csa_tree_add_6_33_groupi_n_1820 ,csa_tree_add_6_33_groupi_n_1415 ,csa_tree_add_6_33_groupi_n_1467);
  or csa_tree_add_6_33_groupi_g16486(csa_tree_add_6_33_groupi_n_1819 ,csa_tree_add_6_33_groupi_n_1073 ,csa_tree_add_6_33_groupi_n_1110);
  and csa_tree_add_6_33_groupi_g16487(csa_tree_add_6_33_groupi_n_1818 ,csa_tree_add_6_33_groupi_n_1406 ,csa_tree_add_6_33_groupi_n_1180);
  and csa_tree_add_6_33_groupi_g16488(csa_tree_add_6_33_groupi_n_1817 ,csa_tree_add_6_33_groupi_n_1218 ,csa_tree_add_6_33_groupi_n_1395);
  or csa_tree_add_6_33_groupi_g16489(csa_tree_add_6_33_groupi_n_1816 ,csa_tree_add_6_33_groupi_n_1113 ,csa_tree_add_6_33_groupi_n_1384);
  or csa_tree_add_6_33_groupi_g16490(csa_tree_add_6_33_groupi_n_1815 ,csa_tree_add_6_33_groupi_n_1399 ,csa_tree_add_6_33_groupi_n_1106);
  and csa_tree_add_6_33_groupi_g16491(csa_tree_add_6_33_groupi_n_1814 ,csa_tree_add_6_33_groupi_n_1159 ,csa_tree_add_6_33_groupi_n_1532);
  and csa_tree_add_6_33_groupi_g16492(csa_tree_add_6_33_groupi_n_1813 ,csa_tree_add_6_33_groupi_n_1122 ,csa_tree_add_6_33_groupi_n_1211);
  and csa_tree_add_6_33_groupi_g16493(csa_tree_add_6_33_groupi_n_1812 ,csa_tree_add_6_33_groupi_n_1506 ,csa_tree_add_6_33_groupi_n_1080);
  and csa_tree_add_6_33_groupi_g16494(csa_tree_add_6_33_groupi_n_1811 ,csa_tree_add_6_33_groupi_n_1085 ,csa_tree_add_6_33_groupi_n_1105);
  or csa_tree_add_6_33_groupi_g16495(csa_tree_add_6_33_groupi_n_1810 ,csa_tree_add_6_33_groupi_n_1423 ,csa_tree_add_6_33_groupi_n_1102);
  or csa_tree_add_6_33_groupi_g16496(csa_tree_add_6_33_groupi_n_1809 ,csa_tree_add_6_33_groupi_n_1146 ,csa_tree_add_6_33_groupi_n_1491);
  or csa_tree_add_6_33_groupi_g16497(csa_tree_add_6_33_groupi_n_1808 ,csa_tree_add_6_33_groupi_n_1153 ,csa_tree_add_6_33_groupi_n_1241);
  and csa_tree_add_6_33_groupi_g16498(csa_tree_add_6_33_groupi_n_1807 ,csa_tree_add_6_33_groupi_n_1239 ,csa_tree_add_6_33_groupi_n_1084);
  or csa_tree_add_6_33_groupi_g16499(csa_tree_add_6_33_groupi_n_1806 ,csa_tree_add_6_33_groupi_n_1219 ,csa_tree_add_6_33_groupi_n_1473);
  and csa_tree_add_6_33_groupi_g16500(csa_tree_add_6_33_groupi_n_1805 ,csa_tree_add_6_33_groupi_n_1434 ,csa_tree_add_6_33_groupi_n_1435);
  and csa_tree_add_6_33_groupi_g16501(csa_tree_add_6_33_groupi_n_1804 ,csa_tree_add_6_33_groupi_n_1112 ,csa_tree_add_6_33_groupi_n_1250);
  and csa_tree_add_6_33_groupi_g16502(csa_tree_add_6_33_groupi_n_1803 ,csa_tree_add_6_33_groupi_n_1124 ,csa_tree_add_6_33_groupi_n_1214);
  or csa_tree_add_6_33_groupi_g16503(csa_tree_add_6_33_groupi_n_1802 ,csa_tree_add_6_33_groupi_n_1490 ,csa_tree_add_6_33_groupi_n_1111);
  and csa_tree_add_6_33_groupi_g16504(csa_tree_add_6_33_groupi_n_1801 ,csa_tree_add_6_33_groupi_n_1373 ,csa_tree_add_6_33_groupi_n_1147);
  and csa_tree_add_6_33_groupi_g16505(csa_tree_add_6_33_groupi_n_1800 ,csa_tree_add_6_33_groupi_n_1471 ,csa_tree_add_6_33_groupi_n_1448);
  or csa_tree_add_6_33_groupi_g16506(csa_tree_add_6_33_groupi_n_1799 ,csa_tree_add_6_33_groupi_n_1372 ,csa_tree_add_6_33_groupi_n_1380);
  nor csa_tree_add_6_33_groupi_g16507(csa_tree_add_6_33_groupi_n_1798 ,csa_tree_add_6_33_groupi_n_1281 ,csa_tree_add_6_33_groupi_n_1065);
  and csa_tree_add_6_33_groupi_g16508(csa_tree_add_6_33_groupi_n_1797 ,csa_tree_add_6_33_groupi_n_1368 ,csa_tree_add_6_33_groupi_n_1100);
  or csa_tree_add_6_33_groupi_g16509(csa_tree_add_6_33_groupi_n_1796 ,csa_tree_add_6_33_groupi_n_1369 ,csa_tree_add_6_33_groupi_n_1234);
  and csa_tree_add_6_33_groupi_g16510(csa_tree_add_6_33_groupi_n_1795 ,csa_tree_add_6_33_groupi_n_1479 ,csa_tree_add_6_33_groupi_n_1364);
  or csa_tree_add_6_33_groupi_g16511(csa_tree_add_6_33_groupi_n_1794 ,csa_tree_add_6_33_groupi_n_1231 ,csa_tree_add_6_33_groupi_n_1120);
  or csa_tree_add_6_33_groupi_g16512(csa_tree_add_6_33_groupi_n_1793 ,csa_tree_add_6_33_groupi_n_1503 ,csa_tree_add_6_33_groupi_n_1186);
  or csa_tree_add_6_33_groupi_g16513(csa_tree_add_6_33_groupi_n_1792 ,csa_tree_add_6_33_groupi_n_785 ,csa_tree_add_6_33_groupi_n_1131);
  and csa_tree_add_6_33_groupi_g16514(csa_tree_add_6_33_groupi_n_1791 ,csa_tree_add_6_33_groupi_n_1154 ,csa_tree_add_6_33_groupi_n_1093);
  or csa_tree_add_6_33_groupi_g16515(csa_tree_add_6_33_groupi_n_1790 ,csa_tree_add_6_33_groupi_n_1424 ,csa_tree_add_6_33_groupi_n_1534);
  or csa_tree_add_6_33_groupi_g16516(csa_tree_add_6_33_groupi_n_1789 ,csa_tree_add_6_33_groupi_n_1139 ,csa_tree_add_6_33_groupi_n_1439);
  and csa_tree_add_6_33_groupi_g16517(csa_tree_add_6_33_groupi_n_1788 ,csa_tree_add_6_33_groupi_n_1196 ,csa_tree_add_6_33_groupi_n_1385);
  or csa_tree_add_6_33_groupi_g16518(csa_tree_add_6_33_groupi_n_1787 ,csa_tree_add_6_33_groupi_n_1373 ,csa_tree_add_6_33_groupi_n_1147);
  and csa_tree_add_6_33_groupi_g16519(csa_tree_add_6_33_groupi_n_1786 ,csa_tree_add_6_33_groupi_n_1193 ,csa_tree_add_6_33_groupi_n_1220);
  or csa_tree_add_6_33_groupi_g16520(csa_tree_add_6_33_groupi_n_1785 ,csa_tree_add_6_33_groupi_n_1474 ,csa_tree_add_6_33_groupi_n_1121);
  and csa_tree_add_6_33_groupi_g16521(csa_tree_add_6_33_groupi_n_1784 ,csa_tree_add_6_33_groupi_n_1466 ,csa_tree_add_6_33_groupi_n_1437);
  or csa_tree_add_6_33_groupi_g16522(csa_tree_add_6_33_groupi_n_1783 ,csa_tree_add_6_33_groupi_n_1493 ,csa_tree_add_6_33_groupi_n_1158);
  and csa_tree_add_6_33_groupi_g16523(csa_tree_add_6_33_groupi_n_1782 ,csa_tree_add_6_33_groupi_n_1389 ,csa_tree_add_6_33_groupi_n_1469);
  or csa_tree_add_6_33_groupi_g16524(csa_tree_add_6_33_groupi_n_1781 ,csa_tree_add_6_33_groupi_n_1196 ,csa_tree_add_6_33_groupi_n_1385);
  and csa_tree_add_6_33_groupi_g16525(csa_tree_add_6_33_groupi_n_1780 ,csa_tree_add_6_33_groupi_n_1502 ,csa_tree_add_6_33_groupi_n_1129);
  or csa_tree_add_6_33_groupi_g16526(csa_tree_add_6_33_groupi_n_1779 ,csa_tree_add_6_33_groupi_n_1243 ,csa_tree_add_6_33_groupi_n_1237);
  and csa_tree_add_6_33_groupi_g16527(csa_tree_add_6_33_groupi_n_1778 ,csa_tree_add_6_33_groupi_n_800 ,csa_tree_add_6_33_groupi_n_1524);
  and csa_tree_add_6_33_groupi_g16528(csa_tree_add_6_33_groupi_n_1777 ,csa_tree_add_6_33_groupi_n_1490 ,csa_tree_add_6_33_groupi_n_1111);
  or csa_tree_add_6_33_groupi_g16529(csa_tree_add_6_33_groupi_n_1776 ,csa_tree_add_6_33_groupi_n_1223 ,csa_tree_add_6_33_groupi_n_1128);
  and csa_tree_add_6_33_groupi_g16530(csa_tree_add_6_33_groupi_n_1775 ,csa_tree_add_6_33_groupi_n_1512 ,csa_tree_add_6_33_groupi_n_1405);
  or csa_tree_add_6_33_groupi_g16531(csa_tree_add_6_33_groupi_n_1774 ,csa_tree_add_6_33_groupi_n_806 ,csa_tree_add_6_33_groupi_n_1440);
  and csa_tree_add_6_33_groupi_g16532(csa_tree_add_6_33_groupi_n_1773 ,csa_tree_add_6_33_groupi_n_1372 ,csa_tree_add_6_33_groupi_n_1380);
  and csa_tree_add_6_33_groupi_g16533(csa_tree_add_6_33_groupi_n_1772 ,csa_tree_add_6_33_groupi_n_1247 ,csa_tree_add_6_33_groupi_n_1201);
  and csa_tree_add_6_33_groupi_g16534(csa_tree_add_6_33_groupi_n_1771 ,csa_tree_add_6_33_groupi_n_1172 ,csa_tree_add_6_33_groupi_n_1182);
  or csa_tree_add_6_33_groupi_g16535(csa_tree_add_6_33_groupi_n_1770 ,csa_tree_add_6_33_groupi_n_1246 ,csa_tree_add_6_33_groupi_n_1527);
  and csa_tree_add_6_33_groupi_g16536(csa_tree_add_6_33_groupi_n_1769 ,csa_tree_add_6_33_groupi_n_1246 ,csa_tree_add_6_33_groupi_n_1527);
  or csa_tree_add_6_33_groupi_g16537(csa_tree_add_6_33_groupi_n_1768 ,csa_tree_add_6_33_groupi_n_1495 ,csa_tree_add_6_33_groupi_n_1500);
  or csa_tree_add_6_33_groupi_g16538(csa_tree_add_6_33_groupi_n_1767 ,csa_tree_add_6_33_groupi_n_773 ,csa_tree_add_6_33_groupi_n_1098);
  and csa_tree_add_6_33_groupi_g16539(csa_tree_add_6_33_groupi_n_1766 ,csa_tree_add_6_33_groupi_n_1486 ,csa_tree_add_6_33_groupi_n_1205);
  or csa_tree_add_6_33_groupi_g16540(csa_tree_add_6_33_groupi_n_1765 ,csa_tree_add_6_33_groupi_n_1095 ,csa_tree_add_6_33_groupi_n_1501);
  and csa_tree_add_6_33_groupi_g16541(csa_tree_add_6_33_groupi_n_1764 ,csa_tree_add_6_33_groupi_n_1184 ,csa_tree_add_6_33_groupi_n_1086);
  and csa_tree_add_6_33_groupi_g16542(csa_tree_add_6_33_groupi_n_1763 ,csa_tree_add_6_33_groupi_n_1480 ,csa_tree_add_6_33_groupi_n_1443);
  and csa_tree_add_6_33_groupi_g16543(csa_tree_add_6_33_groupi_n_1762 ,csa_tree_add_6_33_groupi_n_1108 ,csa_tree_add_6_33_groupi_n_1426);
  or csa_tree_add_6_33_groupi_g16544(csa_tree_add_6_33_groupi_n_1761 ,csa_tree_add_6_33_groupi_n_1154 ,csa_tree_add_6_33_groupi_n_1093);
  and csa_tree_add_6_33_groupi_g16545(csa_tree_add_6_33_groupi_n_1760 ,csa_tree_add_6_33_groupi_n_1438 ,csa_tree_add_6_33_groupi_n_1083);
  or csa_tree_add_6_33_groupi_g16546(csa_tree_add_6_33_groupi_n_1759 ,csa_tree_add_6_33_groupi_n_1466 ,csa_tree_add_6_33_groupi_n_1437);
  or csa_tree_add_6_33_groupi_g16547(csa_tree_add_6_33_groupi_n_1758 ,csa_tree_add_6_33_groupi_n_1104 ,csa_tree_add_6_33_groupi_n_1097);
  or csa_tree_add_6_33_groupi_g16548(csa_tree_add_6_33_groupi_n_1757 ,csa_tree_add_6_33_groupi_n_1472 ,csa_tree_add_6_33_groupi_n_1197);
  nor csa_tree_add_6_33_groupi_g16549(csa_tree_add_6_33_groupi_n_1756 ,csa_tree_add_6_33_groupi_n_125 ,csa_tree_add_6_33_groupi_n_1056);
  and csa_tree_add_6_33_groupi_g16550(csa_tree_add_6_33_groupi_n_1755 ,csa_tree_add_6_33_groupi_n_1173 ,csa_tree_add_6_33_groupi_n_1116);
  or csa_tree_add_6_33_groupi_g16551(csa_tree_add_6_33_groupi_n_1754 ,csa_tree_add_6_33_groupi_n_1112 ,csa_tree_add_6_33_groupi_n_1250);
  nor csa_tree_add_6_33_groupi_g16552(csa_tree_add_6_33_groupi_n_1753 ,csa_tree_add_6_33_groupi_n_1509 ,csa_tree_add_6_33_groupi_n_1210);
  or csa_tree_add_6_33_groupi_g16553(csa_tree_add_6_33_groupi_n_1752 ,csa_tree_add_6_33_groupi_n_1159 ,csa_tree_add_6_33_groupi_n_1532);
  and csa_tree_add_6_33_groupi_g16554(csa_tree_add_6_33_groupi_n_1751 ,csa_tree_add_6_33_groupi_n_1478 ,csa_tree_add_6_33_groupi_n_1521);
  and csa_tree_add_6_33_groupi_g16555(csa_tree_add_6_33_groupi_n_1750 ,csa_tree_add_6_33_groupi_n_1516 ,csa_tree_add_6_33_groupi_n_1078);
  or csa_tree_add_6_33_groupi_g16556(csa_tree_add_6_33_groupi_n_1749 ,csa_tree_add_6_33_groupi_n_1099 ,csa_tree_add_6_33_groupi_n_1189);
  and csa_tree_add_6_33_groupi_g16557(csa_tree_add_6_33_groupi_n_1748 ,csa_tree_add_6_33_groupi_n_1461 ,csa_tree_add_6_33_groupi_n_1475);
  or csa_tree_add_6_33_groupi_g16558(csa_tree_add_6_33_groupi_n_1747 ,csa_tree_add_6_33_groupi_n_1561 ,csa_tree_add_6_33_groupi_n_1059);
  and csa_tree_add_6_33_groupi_g16559(csa_tree_add_6_33_groupi_n_1746 ,csa_tree_add_6_33_groupi_n_1190 ,csa_tree_add_6_33_groupi_n_1403);
  or csa_tree_add_6_33_groupi_g16560(csa_tree_add_6_33_groupi_n_1745 ,csa_tree_add_6_33_groupi_n_1181 ,csa_tree_add_6_33_groupi_n_1463);
  or csa_tree_add_6_33_groupi_g16561(csa_tree_add_6_33_groupi_n_1744 ,csa_tree_add_6_33_groupi_n_1468 ,csa_tree_add_6_33_groupi_n_1453);
  or csa_tree_add_6_33_groupi_g16562(csa_tree_add_6_33_groupi_n_1743 ,csa_tree_add_6_33_groupi_n_1508 ,csa_tree_add_6_33_groupi_n_1209);
  or csa_tree_add_6_33_groupi_g16563(csa_tree_add_6_33_groupi_n_1742 ,csa_tree_add_6_33_groupi_n_1442 ,csa_tree_add_6_33_groupi_n_1077);
  and csa_tree_add_6_33_groupi_g16564(csa_tree_add_6_33_groupi_n_1741 ,csa_tree_add_6_33_groupi_n_1522 ,csa_tree_add_6_33_groupi_n_1421);
  and csa_tree_add_6_33_groupi_g16565(csa_tree_add_6_33_groupi_n_1740 ,csa_tree_add_6_33_groupi_n_1109 ,csa_tree_add_6_33_groupi_n_1382);
  or csa_tree_add_6_33_groupi_g16566(csa_tree_add_6_33_groupi_n_1739 ,csa_tree_add_6_33_groupi_n_1229 ,csa_tree_add_6_33_groupi_n_1446);
  and csa_tree_add_6_33_groupi_g16567(csa_tree_add_6_33_groupi_n_1738 ,csa_tree_add_6_33_groupi_n_1223 ,csa_tree_add_6_33_groupi_n_1128);
  and csa_tree_add_6_33_groupi_g16568(csa_tree_add_6_33_groupi_n_1737 ,csa_tree_add_6_33_groupi_n_1470 ,csa_tree_add_6_33_groupi_n_1132);
  and csa_tree_add_6_33_groupi_g16569(csa_tree_add_6_33_groupi_n_1736 ,csa_tree_add_6_33_groupi_n_1229 ,csa_tree_add_6_33_groupi_n_1446);
  or csa_tree_add_6_33_groupi_g16570(csa_tree_add_6_33_groupi_n_1735 ,csa_tree_add_6_33_groupi_n_1569 ,csa_tree_add_6_33_groupi_n_1357);
  or csa_tree_add_6_33_groupi_g16571(csa_tree_add_6_33_groupi_n_1734 ,csa_tree_add_6_33_groupi_n_1235 ,csa_tree_add_6_33_groupi_n_1071);
  or csa_tree_add_6_33_groupi_g16572(csa_tree_add_6_33_groupi_n_1733 ,csa_tree_add_6_33_groupi_n_1460 ,csa_tree_add_6_33_groupi_n_1420);
  or csa_tree_add_6_33_groupi_g16573(csa_tree_add_6_33_groupi_n_1732 ,csa_tree_add_6_33_groupi_n_1522 ,csa_tree_add_6_33_groupi_n_1421);
  or csa_tree_add_6_33_groupi_g16574(csa_tree_add_6_33_groupi_n_1731 ,csa_tree_add_6_33_groupi_n_1406 ,csa_tree_add_6_33_groupi_n_1180);
  or csa_tree_add_6_33_groupi_g16575(csa_tree_add_6_33_groupi_n_1730 ,csa_tree_add_6_33_groupi_n_1378 ,csa_tree_add_6_33_groupi_n_1140);
  or csa_tree_add_6_33_groupi_g16576(csa_tree_add_6_33_groupi_n_1729 ,csa_tree_add_6_33_groupi_n_1193 ,csa_tree_add_6_33_groupi_n_1220);
  and csa_tree_add_6_33_groupi_g16577(csa_tree_add_6_33_groupi_n_1728 ,csa_tree_add_6_33_groupi_n_1199 ,csa_tree_add_6_33_groupi_n_1430);
  and csa_tree_add_6_33_groupi_g16578(csa_tree_add_6_33_groupi_n_1727 ,csa_tree_add_6_33_groupi_n_1507 ,csa_tree_add_6_33_groupi_n_1431);
  or csa_tree_add_6_33_groupi_g16579(csa_tree_add_6_33_groupi_n_1726 ,csa_tree_add_6_33_groupi_n_809 ,csa_tree_add_6_33_groupi_n_1388);
  or csa_tree_add_6_33_groupi_g16580(csa_tree_add_6_33_groupi_n_1725 ,csa_tree_add_6_33_groupi_n_1236 ,csa_tree_add_6_33_groupi_n_1464);
  or csa_tree_add_6_33_groupi_g16581(csa_tree_add_6_33_groupi_n_1724 ,csa_tree_add_6_33_groupi_n_1502 ,csa_tree_add_6_33_groupi_n_1129);
  and csa_tree_add_6_33_groupi_g16582(csa_tree_add_6_33_groupi_n_1723 ,csa_tree_add_6_33_groupi_n_1381 ,csa_tree_add_6_33_groupi_n_1118);
  or csa_tree_add_6_33_groupi_g16583(csa_tree_add_6_33_groupi_n_1722 ,csa_tree_add_6_33_groupi_n_1156 ,csa_tree_add_6_33_groupi_n_1462);
  and csa_tree_add_6_33_groupi_g16584(csa_tree_add_6_33_groupi_n_1721 ,csa_tree_add_6_33_groupi_n_1383 ,csa_tree_add_6_33_groupi_n_1213);
  and csa_tree_add_6_33_groupi_g16585(csa_tree_add_6_33_groupi_n_1720 ,csa_tree_add_6_33_groupi_n_1503 ,csa_tree_add_6_33_groupi_n_1186);
  or csa_tree_add_6_33_groupi_g16586(csa_tree_add_6_33_groupi_n_1719 ,csa_tree_add_6_33_groupi_n_1184 ,csa_tree_add_6_33_groupi_n_1086);
  and csa_tree_add_6_33_groupi_g16587(csa_tree_add_6_33_groupi_n_1718 ,csa_tree_add_6_33_groupi_n_1505 ,csa_tree_add_6_33_groupi_n_1163);
  or csa_tree_add_6_33_groupi_g16588(csa_tree_add_6_33_groupi_n_1717 ,csa_tree_add_6_33_groupi_n_1164 ,csa_tree_add_6_33_groupi_n_1441);
  and csa_tree_add_6_33_groupi_g16589(csa_tree_add_6_33_groupi_n_1716 ,csa_tree_add_6_33_groupi_n_1235 ,csa_tree_add_6_33_groupi_n_1071);
  or csa_tree_add_6_33_groupi_g16590(csa_tree_add_6_33_groupi_n_1715 ,csa_tree_add_6_33_groupi_n_1581 ,csa_tree_add_6_33_groupi_n_1354);
  or csa_tree_add_6_33_groupi_g16591(csa_tree_add_6_33_groupi_n_1714 ,csa_tree_add_6_33_groupi_n_1456 ,csa_tree_add_6_33_groupi_n_1451);
  and csa_tree_add_6_33_groupi_g16592(csa_tree_add_6_33_groupi_n_1713 ,csa_tree_add_6_33_groupi_n_1219 ,csa_tree_add_6_33_groupi_n_1473);
  or csa_tree_add_6_33_groupi_g16593(csa_tree_add_6_33_groupi_n_1712 ,csa_tree_add_6_33_groupi_n_1488 ,csa_tree_add_6_33_groupi_n_1162);
  and csa_tree_add_6_33_groupi_g16594(csa_tree_add_6_33_groupi_n_1711 ,csa_tree_add_6_33_groupi_n_1442 ,csa_tree_add_6_33_groupi_n_1077);
  or csa_tree_add_6_33_groupi_g16595(csa_tree_add_6_33_groupi_n_1710 ,csa_tree_add_6_33_groupi_n_1108 ,csa_tree_add_6_33_groupi_n_1426);
  or csa_tree_add_6_33_groupi_g16596(csa_tree_add_6_33_groupi_n_1709 ,csa_tree_add_6_33_groupi_n_1471 ,csa_tree_add_6_33_groupi_n_1448);
  or csa_tree_add_6_33_groupi_g16598(csa_tree_add_6_33_groupi_n_1707 ,csa_tree_add_6_33_groupi_n_1558 ,csa_tree_add_6_33_groupi_n_1350);
  or csa_tree_add_6_33_groupi_g16599(csa_tree_add_6_33_groupi_n_1706 ,csa_tree_add_6_33_groupi_n_1195 ,csa_tree_add_6_33_groupi_n_1081);
  or csa_tree_add_6_33_groupi_g16600(csa_tree_add_6_33_groupi_n_1705 ,csa_tree_add_6_33_groupi_n_1232 ,csa_tree_add_6_33_groupi_n_1216);
  nor csa_tree_add_6_33_groupi_g16601(csa_tree_add_6_33_groupi_n_1704 ,csa_tree_add_6_33_groupi_n_1400 ,csa_tree_add_6_33_groupi_n_1107);
  or csa_tree_add_6_33_groupi_g16602(csa_tree_add_6_33_groupi_n_1703 ,csa_tree_add_6_33_groupi_n_776 ,csa_tree_add_6_33_groupi_n_1225);
  or csa_tree_add_6_33_groupi_g16603(csa_tree_add_6_33_groupi_n_1702 ,csa_tree_add_6_33_groupi_n_1383 ,csa_tree_add_6_33_groupi_n_1213);
  and csa_tree_add_6_33_groupi_g16604(csa_tree_add_6_33_groupi_n_1701 ,csa_tree_add_6_33_groupi_n_1468 ,csa_tree_add_6_33_groupi_n_1453);
  and csa_tree_add_6_33_groupi_g16605(csa_tree_add_6_33_groupi_n_1700 ,csa_tree_add_6_33_groupi_n_1422 ,csa_tree_add_6_33_groupi_n_1212);
  or csa_tree_add_6_33_groupi_g16606(csa_tree_add_6_33_groupi_n_1699 ,csa_tree_add_6_33_groupi_n_1176 ,csa_tree_add_6_33_groupi_n_1123);
  or csa_tree_add_6_33_groupi_g16607(csa_tree_add_6_33_groupi_n_1698 ,csa_tree_add_6_33_groupi_n_1160 ,csa_tree_add_6_33_groupi_n_1476);
  or csa_tree_add_6_33_groupi_g16608(csa_tree_add_6_33_groupi_n_1697 ,csa_tree_add_6_33_groupi_n_1096 ,csa_tree_add_6_33_groupi_n_1217);
  and csa_tree_add_6_33_groupi_g16609(csa_tree_add_6_33_groupi_n_1696 ,csa_tree_add_6_33_groupi_n_1076 ,csa_tree_add_6_33_groupi_n_1401);
  or csa_tree_add_6_33_groupi_g16610(csa_tree_add_6_33_groupi_n_1695 ,csa_tree_add_6_33_groupi_n_1419 ,csa_tree_add_6_33_groupi_n_1416);
  or csa_tree_add_6_33_groupi_g16611(csa_tree_add_6_33_groupi_n_1694 ,csa_tree_add_6_33_groupi_n_1428 ,csa_tree_add_6_33_groupi_n_1221);
  and csa_tree_add_6_33_groupi_g16612(csa_tree_add_6_33_groupi_n_1693 ,csa_tree_add_6_33_groupi_n_1497 ,csa_tree_add_6_33_groupi_n_1187);
  and csa_tree_add_6_33_groupi_g16613(csa_tree_add_6_33_groupi_n_1692 ,csa_tree_add_6_33_groupi_n_1175 ,csa_tree_add_6_33_groupi_n_1224);
  and csa_tree_add_6_33_groupi_g16614(csa_tree_add_6_33_groupi_n_1691 ,csa_tree_add_6_33_groupi_n_1369 ,csa_tree_add_6_33_groupi_n_1234);
  and csa_tree_add_6_33_groupi_g16615(csa_tree_add_6_33_groupi_n_1690 ,csa_tree_add_6_33_groupi_n_1427 ,csa_tree_add_6_33_groupi_n_1127);
  and csa_tree_add_6_33_groupi_g16616(csa_tree_add_6_33_groupi_n_1689 ,csa_tree_add_6_33_groupi_n_1202 ,csa_tree_add_6_33_groupi_n_1367);
  or csa_tree_add_6_33_groupi_g16617(csa_tree_add_6_33_groupi_n_1688 ,csa_tree_add_6_33_groupi_n_1389 ,csa_tree_add_6_33_groupi_n_1469);
  or csa_tree_add_6_33_groupi_g16618(csa_tree_add_6_33_groupi_n_1687 ,csa_tree_add_6_33_groupi_n_1516 ,csa_tree_add_6_33_groupi_n_1078);
  or csa_tree_add_6_33_groupi_g16619(csa_tree_add_6_33_groupi_n_1686 ,csa_tree_add_6_33_groupi_n_346 ,csa_tree_add_6_33_groupi_n_1407);
  or csa_tree_add_6_33_groupi_g16620(csa_tree_add_6_33_groupi_n_1685 ,csa_tree_add_6_33_groupi_n_1192 ,csa_tree_add_6_33_groupi_n_1174);
  nor csa_tree_add_6_33_groupi_g16621(csa_tree_add_6_33_groupi_n_1684 ,csa_tree_add_6_33_groupi_n_770 ,csa_tree_add_6_33_groupi_n_1245);
  or csa_tree_add_6_33_groupi_g16622(csa_tree_add_6_33_groupi_n_1683 ,csa_tree_add_6_33_groupi_n_1507 ,csa_tree_add_6_33_groupi_n_1431);
  or csa_tree_add_6_33_groupi_g16623(csa_tree_add_6_33_groupi_n_1682 ,csa_tree_add_6_33_groupi_n_1432 ,csa_tree_add_6_33_groupi_n_1148);
  and csa_tree_add_6_33_groupi_g16624(csa_tree_add_6_33_groupi_n_1681 ,csa_tree_add_6_33_groupi_n_1423 ,csa_tree_add_6_33_groupi_n_1102);
  and csa_tree_add_6_33_groupi_g16625(csa_tree_add_6_33_groupi_n_1680 ,csa_tree_add_6_33_groupi_n_1460 ,csa_tree_add_6_33_groupi_n_1420);
  and csa_tree_add_6_33_groupi_g16626(csa_tree_add_6_33_groupi_n_1679 ,csa_tree_add_6_33_groupi_n_1087 ,csa_tree_add_6_33_groupi_n_1151);
  and csa_tree_add_6_33_groupi_g16627(csa_tree_add_6_33_groupi_n_1678 ,csa_tree_add_6_33_groupi_n_1498 ,csa_tree_add_6_33_groupi_n_1082);
  or csa_tree_add_6_33_groupi_g16628(csa_tree_add_6_33_groupi_n_1677 ,csa_tree_add_6_33_groupi_n_676 ,csa_tree_add_6_33_groupi_n_1365);
  and csa_tree_add_6_33_groupi_g16629(csa_tree_add_6_33_groupi_n_1676 ,csa_tree_add_6_33_groupi_n_1523 ,csa_tree_add_6_33_groupi_n_1228);
  nor csa_tree_add_6_33_groupi_g16630(csa_tree_add_6_33_groupi_n_1675 ,csa_tree_add_6_33_groupi_n_122 ,csa_tree_add_6_33_groupi_n_1362);
  and csa_tree_add_6_33_groupi_g16631(csa_tree_add_6_33_groupi_n_1674 ,csa_tree_add_6_33_groupi_n_1089 ,csa_tree_add_6_33_groupi_n_1117);
  or csa_tree_add_6_33_groupi_g16632(csa_tree_add_6_33_groupi_n_1673 ,csa_tree_add_6_33_groupi_n_1126 ,csa_tree_add_6_33_groupi_n_1240);
  or csa_tree_add_6_33_groupi_g16634(csa_tree_add_6_33_groupi_n_1671 ,csa_tree_add_6_33_groupi_n_1492 ,csa_tree_add_6_33_groupi_n_1165);
  or csa_tree_add_6_33_groupi_g16635(csa_tree_add_6_33_groupi_n_1670 ,csa_tree_add_6_33_groupi_n_1175 ,csa_tree_add_6_33_groupi_n_1224);
  and csa_tree_add_6_33_groupi_g16636(csa_tree_add_6_33_groupi_n_1669 ,csa_tree_add_6_33_groupi_n_1203 ,csa_tree_add_6_33_groupi_n_1141);
  or csa_tree_add_6_33_groupi_g16637(csa_tree_add_6_33_groupi_n_1668 ,csa_tree_add_6_33_groupi_n_1109 ,csa_tree_add_6_33_groupi_n_1382);
  or csa_tree_add_6_33_groupi_g16638(csa_tree_add_6_33_groupi_n_1667 ,csa_tree_add_6_33_groupi_n_1497 ,csa_tree_add_6_33_groupi_n_1187);
  and csa_tree_add_6_33_groupi_g16639(csa_tree_add_6_33_groupi_n_1666 ,csa_tree_add_6_33_groupi_n_1428 ,csa_tree_add_6_33_groupi_n_1221);
  and csa_tree_add_6_33_groupi_g16640(csa_tree_add_6_33_groupi_n_1665 ,csa_tree_add_6_33_groupi_n_1113 ,csa_tree_add_6_33_groupi_n_1384);
  and csa_tree_add_6_33_groupi_g16641(csa_tree_add_6_33_groupi_n_1664 ,csa_tree_add_6_33_groupi_n_1378 ,csa_tree_add_6_33_groupi_n_1140);
  and csa_tree_add_6_33_groupi_g16642(csa_tree_add_6_33_groupi_n_1663 ,csa_tree_add_6_33_groupi_n_803 ,csa_tree_add_6_33_groupi_n_1365);
  or csa_tree_add_6_33_groupi_g16643(csa_tree_add_6_33_groupi_n_1662 ,csa_tree_add_6_33_groupi_n_1371 ,csa_tree_add_6_33_groupi_n_1449);
  or csa_tree_add_6_33_groupi_g16644(csa_tree_add_6_33_groupi_n_1661 ,csa_tree_add_6_33_groupi_n_791 ,csa_tree_add_6_33_groupi_n_1496);
  and csa_tree_add_6_33_groupi_g16645(csa_tree_add_6_33_groupi_n_1660 ,csa_tree_add_6_33_groupi_n_1164 ,csa_tree_add_6_33_groupi_n_1441);
  and csa_tree_add_6_33_groupi_g16646(csa_tree_add_6_33_groupi_n_1659 ,csa_tree_add_6_33_groupi_n_1119 ,csa_tree_add_6_33_groupi_n_1226);
  and csa_tree_add_6_33_groupi_g16647(csa_tree_add_6_33_groupi_n_1658 ,csa_tree_add_6_33_groupi_n_1195 ,csa_tree_add_6_33_groupi_n_1081);
  or csa_tree_add_6_33_groupi_g16648(csa_tree_add_6_33_groupi_n_1657 ,csa_tree_add_6_33_groupi_n_1487 ,csa_tree_add_6_33_groupi_n_1411);
  or csa_tree_add_6_33_groupi_g16649(csa_tree_add_6_33_groupi_n_1656 ,csa_tree_add_6_33_groupi_n_1461 ,csa_tree_add_6_33_groupi_n_1475);
  and csa_tree_add_6_33_groupi_g16650(csa_tree_add_6_33_groupi_n_1655 ,csa_tree_add_6_33_groupi_n_1429 ,csa_tree_add_6_33_groupi_n_1398);
  and csa_tree_add_6_33_groupi_g16651(csa_tree_add_6_33_groupi_n_1654 ,csa_tree_add_6_33_groupi_n_1192 ,csa_tree_add_6_33_groupi_n_1174);
  or csa_tree_add_6_33_groupi_g16652(csa_tree_add_6_33_groupi_n_1653 ,csa_tree_add_6_33_groupi_n_1506 ,csa_tree_add_6_33_groupi_n_1080);
  nor csa_tree_add_6_33_groupi_g16653(csa_tree_add_6_33_groupi_n_1652 ,csa_tree_add_6_33_groupi_n_1600 ,csa_tree_add_6_33_groupi_n_1356);
  and csa_tree_add_6_33_groupi_g16654(csa_tree_add_6_33_groupi_n_1651 ,csa_tree_add_6_33_groupi_n_1236 ,csa_tree_add_6_33_groupi_n_1464);
  xnor csa_tree_add_6_33_groupi_g16655(csa_tree_add_6_33_groupi_n_1650 ,in1[1] ,in3[2]);
  xnor csa_tree_add_6_33_groupi_g16656(csa_tree_add_6_33_groupi_n_1649 ,in1[0] ,in2[0]);
  xnor csa_tree_add_6_33_groupi_g16657(csa_tree_add_6_33_groupi_n_1648 ,in3[10] ,in2[10]);
  xnor csa_tree_add_6_33_groupi_g16658(csa_tree_add_6_33_groupi_n_1647 ,in3[27] ,in2[27]);
  xnor csa_tree_add_6_33_groupi_g16659(csa_tree_add_6_33_groupi_n_1646 ,in3[22] ,in2[22]);
  xnor csa_tree_add_6_33_groupi_g16660(csa_tree_add_6_33_groupi_n_1645 ,in3[12] ,in2[12]);
  xnor csa_tree_add_6_33_groupi_g16661(csa_tree_add_6_33_groupi_n_1644 ,in3[8] ,in2[8]);
  xnor csa_tree_add_6_33_groupi_g16662(csa_tree_add_6_33_groupi_n_1643 ,in3[11] ,in2[11]);
  xnor csa_tree_add_6_33_groupi_g16663(csa_tree_add_6_33_groupi_n_1642 ,in3[9] ,in2[9]);
  xnor csa_tree_add_6_33_groupi_g16664(csa_tree_add_6_33_groupi_n_1641 ,in3[18] ,in2[18]);
  xnor csa_tree_add_6_33_groupi_g16665(csa_tree_add_6_33_groupi_n_1640 ,in3[16] ,in2[16]);
  xnor csa_tree_add_6_33_groupi_g16666(csa_tree_add_6_33_groupi_n_1639 ,in3[29] ,in2[29]);
  xnor csa_tree_add_6_33_groupi_g16667(csa_tree_add_6_33_groupi_n_1638 ,in3[4] ,in2[4]);
  xnor csa_tree_add_6_33_groupi_g16668(csa_tree_add_6_33_groupi_n_1637 ,in3[15] ,in2[15]);
  xnor csa_tree_add_6_33_groupi_g16669(csa_tree_add_6_33_groupi_n_1636 ,in3[14] ,in2[14]);
  xnor csa_tree_add_6_33_groupi_g16670(csa_tree_add_6_33_groupi_n_1635 ,in3[6] ,in2[6]);
  xnor csa_tree_add_6_33_groupi_g16671(csa_tree_add_6_33_groupi_n_1634 ,in3[28] ,in2[28]);
  xnor csa_tree_add_6_33_groupi_g16672(csa_tree_add_6_33_groupi_n_1633 ,in3[7] ,in2[7]);
  xnor csa_tree_add_6_33_groupi_g16673(csa_tree_add_6_33_groupi_n_1632 ,in3[25] ,in2[25]);
  xnor csa_tree_add_6_33_groupi_g16674(csa_tree_add_6_33_groupi_n_1631 ,in3[17] ,in2[17]);
  xnor csa_tree_add_6_33_groupi_g16675(csa_tree_add_6_33_groupi_n_1630 ,in3[23] ,in2[23]);
  xnor csa_tree_add_6_33_groupi_g16676(csa_tree_add_6_33_groupi_n_1629 ,in3[19] ,in2[19]);
  xnor csa_tree_add_6_33_groupi_g16677(csa_tree_add_6_33_groupi_n_1628 ,in3[20] ,in2[20]);
  xnor csa_tree_add_6_33_groupi_g16678(csa_tree_add_6_33_groupi_n_1627 ,in3[26] ,in2[26]);
  xnor csa_tree_add_6_33_groupi_g16679(csa_tree_add_6_33_groupi_n_1626 ,in3[24] ,in2[24]);
  xnor csa_tree_add_6_33_groupi_g16680(csa_tree_add_6_33_groupi_n_1625 ,in3[1] ,in2[1]);
  xnor csa_tree_add_6_33_groupi_g16681(csa_tree_add_6_33_groupi_n_1624 ,in3[30] ,in2[30]);
  xnor csa_tree_add_6_33_groupi_g16682(csa_tree_add_6_33_groupi_n_1623 ,in3[21] ,in2[21]);
  xnor csa_tree_add_6_33_groupi_g16683(csa_tree_add_6_33_groupi_n_1622 ,in3[3] ,in2[3]);
  xnor csa_tree_add_6_33_groupi_g16684(csa_tree_add_6_33_groupi_n_1621 ,in3[31] ,in2[31]);
  xnor csa_tree_add_6_33_groupi_g16685(csa_tree_add_6_33_groupi_n_1620 ,in3[5] ,in2[5]);
  xnor csa_tree_add_6_33_groupi_g16686(csa_tree_add_6_33_groupi_n_1619 ,in3[13] ,in2[13]);
  not csa_tree_add_6_33_groupi_g16687(csa_tree_add_6_33_groupi_n_1534 ,csa_tree_add_6_33_groupi_n_1535);
  not csa_tree_add_6_33_groupi_g16688(csa_tree_add_6_33_groupi_n_1518 ,csa_tree_add_6_33_groupi_n_1519);
  not csa_tree_add_6_33_groupi_g16689(csa_tree_add_6_33_groupi_n_1508 ,csa_tree_add_6_33_groupi_n_1509);
  not csa_tree_add_6_33_groupi_g16690(csa_tree_add_6_33_groupi_n_1483 ,csa_tree_add_6_33_groupi_n_1484);
  not csa_tree_add_6_33_groupi_g16691(csa_tree_add_6_33_groupi_n_1476 ,csa_tree_add_6_33_groupi_n_1477);
  not csa_tree_add_6_33_groupi_g16692(csa_tree_add_6_33_groupi_n_1424 ,csa_tree_add_6_33_groupi_n_1425);
  not csa_tree_add_6_33_groupi_g16693(csa_tree_add_6_33_groupi_n_1414 ,csa_tree_add_6_33_groupi_n_1413);
  not csa_tree_add_6_33_groupi_g16694(csa_tree_add_6_33_groupi_n_1409 ,csa_tree_add_6_33_groupi_n_1410);
  not csa_tree_add_6_33_groupi_g16695(csa_tree_add_6_33_groupi_n_1399 ,csa_tree_add_6_33_groupi_n_1400);
  not csa_tree_add_6_33_groupi_g16696(csa_tree_add_6_33_groupi_n_1396 ,csa_tree_add_6_33_groupi_n_1397);
  not csa_tree_add_6_33_groupi_g16697(csa_tree_add_6_33_groupi_n_1375 ,csa_tree_add_6_33_groupi_n_1376);
  and csa_tree_add_6_33_groupi_g16698(csa_tree_add_6_33_groupi_n_1363 ,in3[29] ,in2[29]);
  nor csa_tree_add_6_33_groupi_g16699(csa_tree_add_6_33_groupi_n_1362 ,in3[0] ,in2[0]);
  or csa_tree_add_6_33_groupi_g16700(csa_tree_add_6_33_groupi_n_1361 ,in1[1] ,in3[2]);
  and csa_tree_add_6_33_groupi_g16701(csa_tree_add_6_33_groupi_n_1360 ,in1[11] ,in3[22]);
  and csa_tree_add_6_33_groupi_g16702(csa_tree_add_6_33_groupi_n_1359 ,in3[3] ,in2[3]);
  and csa_tree_add_6_33_groupi_g16703(csa_tree_add_6_33_groupi_n_1358 ,in1[2] ,in2[4]);
  nor csa_tree_add_6_33_groupi_g16704(csa_tree_add_6_33_groupi_n_1357 ,in3[5] ,in2[5]);
  nor csa_tree_add_6_33_groupi_g16705(csa_tree_add_6_33_groupi_n_1356 ,in3[7] ,in2[7]);
  or csa_tree_add_6_33_groupi_g16706(csa_tree_add_6_33_groupi_n_1355 ,in1[13] ,in3[26]);
  nor csa_tree_add_6_33_groupi_g16707(csa_tree_add_6_33_groupi_n_1354 ,in3[19] ,in2[19]);
  and csa_tree_add_6_33_groupi_g16708(csa_tree_add_6_33_groupi_n_1353 ,in3[7] ,in2[7]);
  nand csa_tree_add_6_33_groupi_g16709(csa_tree_add_6_33_groupi_n_1352 ,in3[31] ,in2[31]);
  nor csa_tree_add_6_33_groupi_g16710(csa_tree_add_6_33_groupi_n_1351 ,in3[31] ,in2[31]);
  nor csa_tree_add_6_33_groupi_g16711(csa_tree_add_6_33_groupi_n_1350 ,in3[27] ,in2[27]);
  or csa_tree_add_6_33_groupi_g16712(csa_tree_add_6_33_groupi_n_1349 ,in1[15] ,in3[30]);
  nor csa_tree_add_6_33_groupi_g16713(csa_tree_add_6_33_groupi_n_1348 ,in3[8] ,in2[8]);
  nand csa_tree_add_6_33_groupi_g16714(csa_tree_add_6_33_groupi_n_1347 ,in3[1] ,in2[1]);
  nor csa_tree_add_6_33_groupi_g16715(csa_tree_add_6_33_groupi_n_1346 ,in3[3] ,in2[3]);
  nor csa_tree_add_6_33_groupi_g16716(csa_tree_add_6_33_groupi_n_1345 ,in3[11] ,in2[11]);
  and csa_tree_add_6_33_groupi_g16717(csa_tree_add_6_33_groupi_n_1344 ,in1[7] ,in3[14]);
  or csa_tree_add_6_33_groupi_g16718(csa_tree_add_6_33_groupi_n_1343 ,in1[5] ,in3[10]);
  and csa_tree_add_6_33_groupi_g16719(csa_tree_add_6_33_groupi_n_1342 ,in3[13] ,in2[13]);
  and csa_tree_add_6_33_groupi_g16720(csa_tree_add_6_33_groupi_n_1341 ,in3[0] ,in2[0]);
  or csa_tree_add_6_33_groupi_g16721(csa_tree_add_6_33_groupi_n_1340 ,in1[7] ,in3[14]);
  or csa_tree_add_6_33_groupi_g16722(csa_tree_add_6_33_groupi_n_1339 ,in1[14] ,in3[28]);
  and csa_tree_add_6_33_groupi_g16723(csa_tree_add_6_33_groupi_n_1338 ,in3[9] ,in2[9]);
  or csa_tree_add_6_33_groupi_g16724(csa_tree_add_6_33_groupi_n_1337 ,in1[11] ,in3[22]);
  nand csa_tree_add_6_33_groupi_g16725(csa_tree_add_6_33_groupi_n_1336 ,in3[23] ,in2[23]);
  or csa_tree_add_6_33_groupi_g16726(csa_tree_add_6_33_groupi_n_1335 ,in1[6] ,in3[12]);
  nor csa_tree_add_6_33_groupi_g16727(csa_tree_add_6_33_groupi_n_1334 ,in3[23] ,in2[23]);
  nor csa_tree_add_6_33_groupi_g16728(csa_tree_add_6_33_groupi_n_1333 ,in3[9] ,in2[9]);
  nor csa_tree_add_6_33_groupi_g16729(csa_tree_add_6_33_groupi_n_1332 ,in3[15] ,in2[15]);
  or csa_tree_add_6_33_groupi_g16730(csa_tree_add_6_33_groupi_n_1331 ,in1[10] ,in3[20]);
  and csa_tree_add_6_33_groupi_g16731(csa_tree_add_6_33_groupi_n_1330 ,in3[15] ,in2[15]);
  and csa_tree_add_6_33_groupi_g16732(csa_tree_add_6_33_groupi_n_1329 ,in3[11] ,in2[11]);
  nor csa_tree_add_6_33_groupi_g16733(csa_tree_add_6_33_groupi_n_1328 ,in1[8] ,in3[16]);
  or csa_tree_add_6_33_groupi_g16734(csa_tree_add_6_33_groupi_n_1618 ,csa_tree_add_6_33_groupi_n_532 ,csa_tree_add_6_33_groupi_n_469);
  or csa_tree_add_6_33_groupi_g16735(csa_tree_add_6_33_groupi_n_1617 ,csa_tree_add_6_33_groupi_n_580 ,csa_tree_add_6_33_groupi_n_310);
  or csa_tree_add_6_33_groupi_g16736(csa_tree_add_6_33_groupi_n_1616 ,csa_tree_add_6_33_groupi_n_202 ,csa_tree_add_6_33_groupi_n_247);
  or csa_tree_add_6_33_groupi_g16737(csa_tree_add_6_33_groupi_n_1615 ,csa_tree_add_6_33_groupi_n_406 ,csa_tree_add_6_33_groupi_n_316);
  or csa_tree_add_6_33_groupi_g16738(csa_tree_add_6_33_groupi_n_1614 ,csa_tree_add_6_33_groupi_n_484 ,csa_tree_add_6_33_groupi_n_604);
  or csa_tree_add_6_33_groupi_g16739(csa_tree_add_6_33_groupi_n_1613 ,csa_tree_add_6_33_groupi_n_592 ,csa_tree_add_6_33_groupi_n_388);
  or csa_tree_add_6_33_groupi_g16740(csa_tree_add_6_33_groupi_n_1612 ,csa_tree_add_6_33_groupi_n_616 ,csa_tree_add_6_33_groupi_n_382);
  or csa_tree_add_6_33_groupi_g16741(csa_tree_add_6_33_groupi_n_1611 ,csa_tree_add_6_33_groupi_n_157 ,csa_tree_add_6_33_groupi_n_520);
  or csa_tree_add_6_33_groupi_g16742(csa_tree_add_6_33_groupi_n_1610 ,csa_tree_add_6_33_groupi_n_640 ,csa_tree_add_6_33_groupi_n_586);
  or csa_tree_add_6_33_groupi_g16743(csa_tree_add_6_33_groupi_n_1609 ,csa_tree_add_6_33_groupi_n_562 ,csa_tree_add_6_33_groupi_n_394);
  or csa_tree_add_6_33_groupi_g16744(csa_tree_add_6_33_groupi_n_1608 ,csa_tree_add_6_33_groupi_n_184 ,csa_tree_add_6_33_groupi_n_655);
  or csa_tree_add_6_33_groupi_g16745(csa_tree_add_6_33_groupi_n_1607 ,csa_tree_add_6_33_groupi_n_544 ,csa_tree_add_6_33_groupi_n_646);
  or csa_tree_add_6_33_groupi_g16746(csa_tree_add_6_33_groupi_n_1606 ,csa_tree_add_6_33_groupi_n_328 ,csa_tree_add_6_33_groupi_n_445);
  or csa_tree_add_6_33_groupi_g16747(csa_tree_add_6_33_groupi_n_1605 ,csa_tree_add_6_33_groupi_n_722 ,csa_tree_add_6_33_groupi_n_142);
  or csa_tree_add_6_33_groupi_g16748(csa_tree_add_6_33_groupi_n_1604 ,csa_tree_add_6_33_groupi_n_538 ,csa_tree_add_6_33_groupi_n_220);
  or csa_tree_add_6_33_groupi_g16749(csa_tree_add_6_33_groupi_n_1603 ,csa_tree_add_6_33_groupi_n_322 ,csa_tree_add_6_33_groupi_n_583);
  or csa_tree_add_6_33_groupi_g16750(csa_tree_add_6_33_groupi_n_1602 ,csa_tree_add_6_33_groupi_n_238 ,csa_tree_add_6_33_groupi_n_377);
  or csa_tree_add_6_33_groupi_g16751(csa_tree_add_6_33_groupi_n_1601 ,csa_tree_add_6_33_groupi_n_688 ,csa_tree_add_6_33_groupi_n_760);
  or csa_tree_add_6_33_groupi_g16752(csa_tree_add_6_33_groupi_n_1600 ,csa_tree_add_6_33_groupi_n_464 ,csa_tree_add_6_33_groupi_n_206);
  or csa_tree_add_6_33_groupi_g16753(csa_tree_add_6_33_groupi_n_1599 ,csa_tree_add_6_33_groupi_n_574 ,csa_tree_add_6_33_groupi_n_670);
  or csa_tree_add_6_33_groupi_g16754(csa_tree_add_6_33_groupi_n_1598 ,csa_tree_add_6_33_groupi_n_448 ,csa_tree_add_6_33_groupi_n_607);
  or csa_tree_add_6_33_groupi_g16755(csa_tree_add_6_33_groupi_n_1597 ,csa_tree_add_6_33_groupi_n_160 ,csa_tree_add_6_33_groupi_n_496);
  or csa_tree_add_6_33_groupi_g16756(csa_tree_add_6_33_groupi_n_1596 ,csa_tree_add_6_33_groupi_n_280 ,csa_tree_add_6_33_groupi_n_514);
  or csa_tree_add_6_33_groupi_g16757(csa_tree_add_6_33_groupi_n_1595 ,csa_tree_add_6_33_groupi_n_250 ,csa_tree_add_6_33_groupi_n_754);
  or csa_tree_add_6_33_groupi_g16758(csa_tree_add_6_33_groupi_n_1594 ,csa_tree_add_6_33_groupi_n_424 ,csa_tree_add_6_33_groupi_n_577);
  or csa_tree_add_6_33_groupi_g16759(csa_tree_add_6_33_groupi_n_1593 ,csa_tree_add_6_33_groupi_n_475 ,csa_tree_add_6_33_groupi_n_256);
  or csa_tree_add_6_33_groupi_g16760(csa_tree_add_6_33_groupi_n_1592 ,csa_tree_add_6_33_groupi_n_226 ,csa_tree_add_6_33_groupi_n_167);
  or csa_tree_add_6_33_groupi_g16761(csa_tree_add_6_33_groupi_n_1591 ,csa_tree_add_6_33_groupi_n_682 ,csa_tree_add_6_33_groupi_n_746);
  or csa_tree_add_6_33_groupi_g16762(csa_tree_add_6_33_groupi_n_1590 ,csa_tree_add_6_33_groupi_n_139 ,csa_tree_add_6_33_groupi_n_674);
  or csa_tree_add_6_33_groupi_g16763(csa_tree_add_6_33_groupi_n_1589 ,csa_tree_add_6_33_groupi_n_550 ,csa_tree_add_6_33_groupi_n_763);
  or csa_tree_add_6_33_groupi_g16764(csa_tree_add_6_33_groupi_n_1588 ,csa_tree_add_6_33_groupi_n_451 ,csa_tree_add_6_33_groupi_n_622);
  or csa_tree_add_6_33_groupi_g16765(csa_tree_add_6_33_groupi_n_1587 ,csa_tree_add_6_33_groupi_n_283 ,csa_tree_add_6_33_groupi_n_163);
  or csa_tree_add_6_33_groupi_g16766(csa_tree_add_6_33_groupi_n_1586 ,csa_tree_add_6_33_groupi_n_259 ,csa_tree_add_6_33_groupi_n_559);
  or csa_tree_add_6_33_groupi_g16767(csa_tree_add_6_33_groupi_n_1585 ,csa_tree_add_6_33_groupi_n_460 ,csa_tree_add_6_33_groupi_n_353);
  or csa_tree_add_6_33_groupi_g16768(csa_tree_add_6_33_groupi_n_1584 ,csa_tree_add_6_33_groupi_n_343 ,csa_tree_add_6_33_groupi_n_752);
  or csa_tree_add_6_33_groupi_g16769(csa_tree_add_6_33_groupi_n_1583 ,csa_tree_add_6_33_groupi_n_217 ,csa_tree_add_6_33_groupi_n_292);
  or csa_tree_add_6_33_groupi_g16770(csa_tree_add_6_33_groupi_n_1582 ,csa_tree_add_6_33_groupi_n_53 ,csa_tree_add_6_33_groupi_n_358);
  or csa_tree_add_6_33_groupi_g16771(csa_tree_add_6_33_groupi_n_1581 ,csa_tree_add_6_33_groupi_n_370 ,csa_tree_add_6_33_groupi_n_700);
  or csa_tree_add_6_33_groupi_g16772(csa_tree_add_6_33_groupi_n_1580 ,csa_tree_add_6_33_groupi_n_523 ,csa_tree_add_6_33_groupi_n_230);
  or csa_tree_add_6_33_groupi_g16773(csa_tree_add_6_33_groupi_n_1579 ,csa_tree_add_6_33_groupi_n_170 ,csa_tree_add_6_33_groupi_n_658);
  or csa_tree_add_6_33_groupi_g16774(csa_tree_add_6_33_groupi_n_1578 ,csa_tree_add_6_33_groupi_n_331 ,csa_tree_add_6_33_groupi_n_667);
  or csa_tree_add_6_33_groupi_g16775(csa_tree_add_6_33_groupi_n_1577 ,csa_tree_add_6_33_groupi_n_337 ,csa_tree_add_6_33_groupi_n_698);
  or csa_tree_add_6_33_groupi_g16776(csa_tree_add_6_33_groupi_n_1576 ,csa_tree_add_6_33_groupi_n_728 ,csa_tree_add_6_33_groupi_n_662);
  or csa_tree_add_6_33_groupi_g16777(csa_tree_add_6_33_groupi_n_1575 ,csa_tree_add_6_33_groupi_n_436 ,csa_tree_add_6_33_groupi_n_595);
  or csa_tree_add_6_33_groupi_g16778(csa_tree_add_6_33_groupi_n_1574 ,csa_tree_add_6_33_groupi_n_706 ,csa_tree_add_6_33_groupi_n_571);
  or csa_tree_add_6_33_groupi_g16779(csa_tree_add_6_33_groupi_n_1573 ,csa_tree_add_6_33_groupi_n_694 ,csa_tree_add_6_33_groupi_n_587);
  or csa_tree_add_6_33_groupi_g16780(csa_tree_add_6_33_groupi_n_1572 ,csa_tree_add_6_33_groupi_n_275 ,csa_tree_add_6_33_groupi_n_236);
  or csa_tree_add_6_33_groupi_g16781(csa_tree_add_6_33_groupi_n_1571 ,csa_tree_add_6_33_groupi_n_490 ,csa_tree_add_6_33_groupi_n_196);
  or csa_tree_add_6_33_groupi_g16782(csa_tree_add_6_33_groupi_n_1570 ,csa_tree_add_6_33_groupi_n_130 ,csa_tree_add_6_33_groupi_n_391);
  or csa_tree_add_6_33_groupi_g16783(csa_tree_add_6_33_groupi_n_1569 ,csa_tree_add_6_33_groupi_n_307 ,csa_tree_add_6_33_groupi_n_710);
  or csa_tree_add_6_33_groupi_g16784(csa_tree_add_6_33_groupi_n_1568 ,csa_tree_add_6_33_groupi_n_796 ,csa_tree_add_6_33_groupi_n_418);
  or csa_tree_add_6_33_groupi_g16785(csa_tree_add_6_33_groupi_n_1567 ,csa_tree_add_6_33_groupi_n_199 ,csa_tree_add_6_33_groupi_n_241);
  or csa_tree_add_6_33_groupi_g16786(csa_tree_add_6_33_groupi_n_1566 ,csa_tree_add_6_33_groupi_n_704 ,csa_tree_add_6_33_groupi_n_397);
  or csa_tree_add_6_33_groupi_g16787(csa_tree_add_6_33_groupi_n_1565 ,csa_tree_add_6_33_groupi_n_508 ,csa_tree_add_6_33_groupi_n_379);
  or csa_tree_add_6_33_groupi_g16788(csa_tree_add_6_33_groupi_n_1564 ,csa_tree_add_6_33_groupi_n_364 ,csa_tree_add_6_33_groupi_n_581);
  or csa_tree_add_6_33_groupi_g16789(csa_tree_add_6_33_groupi_n_1563 ,csa_tree_add_6_33_groupi_n_466 ,csa_tree_add_6_33_groupi_n_455);
  or csa_tree_add_6_33_groupi_g16790(csa_tree_add_6_33_groupi_n_1562 ,csa_tree_add_6_33_groupi_n_748 ,csa_tree_add_6_33_groupi_n_692);
  or csa_tree_add_6_33_groupi_g16791(csa_tree_add_6_33_groupi_n_1561 ,csa_tree_add_6_33_groupi_n_401 ,csa_tree_add_6_33_groupi_n_686);
  or csa_tree_add_6_33_groupi_g16792(csa_tree_add_6_33_groupi_n_1560 ,csa_tree_add_6_33_groupi_n_190 ,csa_tree_add_6_33_groupi_n_253);
  or csa_tree_add_6_33_groupi_g16793(csa_tree_add_6_33_groupi_n_1559 ,csa_tree_add_6_33_groupi_n_149 ,csa_tree_add_6_33_groupi_n_649);
  or csa_tree_add_6_33_groupi_g16794(csa_tree_add_6_33_groupi_n_1558 ,csa_tree_add_6_33_groupi_n_715 ,csa_tree_add_6_33_groupi_n_208);
  or csa_tree_add_6_33_groupi_g16795(csa_tree_add_6_33_groupi_n_1557 ,csa_tree_add_6_33_groupi_n_403 ,csa_tree_add_6_33_groupi_n_263);
  or csa_tree_add_6_33_groupi_g16796(csa_tree_add_6_33_groupi_n_1556 ,csa_tree_add_6_33_groupi_n_430 ,csa_tree_add_6_33_groupi_n_742);
  or csa_tree_add_6_33_groupi_g16797(csa_tree_add_6_33_groupi_n_1555 ,csa_tree_add_6_33_groupi_n_412 ,csa_tree_add_6_33_groupi_n_127);
  or csa_tree_add_6_33_groupi_g16798(csa_tree_add_6_33_groupi_n_1554 ,csa_tree_add_6_33_groupi_n_277 ,csa_tree_add_6_33_groupi_n_151);
  or csa_tree_add_6_33_groupi_g16799(csa_tree_add_6_33_groupi_n_1553 ,csa_tree_add_6_33_groupi_n_325 ,csa_tree_add_6_33_groupi_n_472);
  or csa_tree_add_6_33_groupi_g16800(csa_tree_add_6_33_groupi_n_1552 ,csa_tree_add_6_33_groupi_n_634 ,csa_tree_add_6_33_groupi_n_355);
  or csa_tree_add_6_33_groupi_g16801(csa_tree_add_6_33_groupi_n_1551 ,csa_tree_add_6_33_groupi_n_758 ,csa_tree_add_6_33_groupi_n_664);
  or csa_tree_add_6_33_groupi_g16802(csa_tree_add_6_33_groupi_n_1550 ,csa_tree_add_6_33_groupi_n_266 ,csa_tree_add_6_33_groupi_n_107);
  or csa_tree_add_6_33_groupi_g16803(csa_tree_add_6_33_groupi_n_1549 ,csa_tree_add_6_33_groupi_n_361 ,csa_tree_add_6_33_groupi_n_229);
  or csa_tree_add_6_33_groupi_g16804(csa_tree_add_6_33_groupi_n_1548 ,csa_tree_add_6_33_groupi_n_565 ,csa_tree_add_6_33_groupi_n_553);
  or csa_tree_add_6_33_groupi_g16805(csa_tree_add_6_33_groupi_n_1547 ,csa_tree_add_6_33_groupi_n_766 ,csa_tree_add_6_33_groupi_n_541);
  or csa_tree_add_6_33_groupi_g16806(csa_tree_add_6_33_groupi_n_1546 ,csa_tree_add_6_33_groupi_n_499 ,csa_tree_add_6_33_groupi_n_349);
  or csa_tree_add_6_33_groupi_g16807(csa_tree_add_6_33_groupi_n_1545 ,csa_tree_add_6_33_groupi_n_145 ,csa_tree_add_6_33_groupi_n_65);
  or csa_tree_add_6_33_groupi_g16808(csa_tree_add_6_33_groupi_n_1544 ,csa_tree_add_6_33_groupi_n_479 ,csa_tree_add_6_33_groupi_n_463);
  or csa_tree_add_6_33_groupi_g16809(csa_tree_add_6_33_groupi_n_1543 ,csa_tree_add_6_33_groupi_n_563 ,csa_tree_add_6_33_groupi_n_113);
  or csa_tree_add_6_33_groupi_g16810(csa_tree_add_6_33_groupi_n_1542 ,csa_tree_add_6_33_groupi_n_175 ,csa_tree_add_6_33_groupi_n_116);
  or csa_tree_add_6_33_groupi_g16811(csa_tree_add_6_33_groupi_n_1541 ,csa_tree_add_6_33_groupi_n_481 ,csa_tree_add_6_33_groupi_n_110);
  or csa_tree_add_6_33_groupi_g16812(csa_tree_add_6_33_groupi_n_1540 ,csa_tree_add_6_33_groupi_n_232 ,csa_tree_add_6_33_groupi_n_517);
  or csa_tree_add_6_33_groupi_g16813(csa_tree_add_6_33_groupi_n_1539 ,csa_tree_add_6_33_groupi_n_775 ,csa_tree_add_6_33_groupi_n_433);
  or csa_tree_add_6_33_groupi_g16814(csa_tree_add_6_33_groupi_n_1538 ,csa_tree_add_6_33_groupi_n_98 ,csa_tree_add_6_33_groupi_n_221);
  or csa_tree_add_6_33_groupi_g16815(csa_tree_add_6_33_groupi_n_1537 ,csa_tree_add_6_33_groupi_n_383 ,csa_tree_add_6_33_groupi_n_77);
  or csa_tree_add_6_33_groupi_g16816(csa_tree_add_6_33_groupi_n_1536 ,csa_tree_add_6_33_groupi_n_385 ,csa_tree_add_6_33_groupi_n_629);
  or csa_tree_add_6_33_groupi_g16817(csa_tree_add_6_33_groupi_n_1535 ,csa_tree_add_6_33_groupi_n_421 ,csa_tree_add_6_33_groupi_n_302);
  or csa_tree_add_6_33_groupi_g16818(csa_tree_add_6_33_groupi_n_1533 ,csa_tree_add_6_33_groupi_n_547 ,csa_tree_add_6_33_groupi_n_50);
  or csa_tree_add_6_33_groupi_g16819(csa_tree_add_6_33_groupi_n_1532 ,csa_tree_add_6_33_groupi_n_722 ,csa_tree_add_6_33_groupi_n_740);
  or csa_tree_add_6_33_groupi_g16820(csa_tree_add_6_33_groupi_n_1531 ,csa_tree_add_6_33_groupi_n_193 ,csa_tree_add_6_33_groupi_n_656);
  or csa_tree_add_6_33_groupi_g16821(csa_tree_add_6_33_groupi_n_1530 ,csa_tree_add_6_33_groupi_n_134 ,csa_tree_add_6_33_groupi_n_311);
  or csa_tree_add_6_33_groupi_g16822(csa_tree_add_6_33_groupi_n_1529 ,csa_tree_add_6_33_groupi_n_493 ,csa_tree_add_6_33_groupi_n_511);
  or csa_tree_add_6_33_groupi_g16823(csa_tree_add_6_33_groupi_n_1528 ,csa_tree_add_6_33_groupi_n_671 ,csa_tree_add_6_33_groupi_n_367);
  or csa_tree_add_6_33_groupi_g16824(csa_tree_add_6_33_groupi_n_1527 ,csa_tree_add_6_33_groupi_n_203 ,csa_tree_add_6_33_groupi_n_359);
  or csa_tree_add_6_33_groupi_g16825(csa_tree_add_6_33_groupi_n_1526 ,csa_tree_add_6_33_groupi_n_535 ,csa_tree_add_6_33_groupi_n_601);
  or csa_tree_add_6_33_groupi_g16826(csa_tree_add_6_33_groupi_n_1525 ,csa_tree_add_6_33_groupi_n_181 ,csa_tree_add_6_33_groupi_n_619);
  or csa_tree_add_6_33_groupi_g16827(csa_tree_add_6_33_groupi_n_1524 ,csa_tree_add_6_33_groupi_n_589 ,csa_tree_add_6_33_groupi_n_313);
  or csa_tree_add_6_33_groupi_g16828(csa_tree_add_6_33_groupi_n_1523 ,csa_tree_add_6_33_groupi_n_529 ,csa_tree_add_6_33_groupi_n_781);
  or csa_tree_add_6_33_groupi_g16829(csa_tree_add_6_33_groupi_n_1522 ,csa_tree_add_6_33_groupi_n_439 ,csa_tree_add_6_33_groupi_n_161);
  or csa_tree_add_6_33_groupi_g16830(csa_tree_add_6_33_groupi_n_1521 ,csa_tree_add_6_33_groupi_n_136 ,csa_tree_add_6_33_groupi_n_173);
  or csa_tree_add_6_33_groupi_g16831(csa_tree_add_6_33_groupi_n_1520 ,csa_tree_add_6_33_groupi_n_799 ,csa_tree_add_6_33_groupi_n_734);
  or csa_tree_add_6_33_groupi_g16832(csa_tree_add_6_33_groupi_n_1519 ,csa_tree_add_6_33_groupi_n_124 ,csa_tree_add_6_33_groupi_n_211);
  or csa_tree_add_6_33_groupi_g16833(csa_tree_add_6_33_groupi_n_1517 ,csa_tree_add_6_33_groupi_n_611 ,csa_tree_add_6_33_groupi_n_80);
  or csa_tree_add_6_33_groupi_g16834(csa_tree_add_6_33_groupi_n_1516 ,csa_tree_add_6_33_groupi_n_295 ,csa_tree_add_6_33_groupi_n_268);
  or csa_tree_add_6_33_groupi_g16835(csa_tree_add_6_33_groupi_n_1515 ,csa_tree_add_6_33_groupi_n_442 ,csa_tree_add_6_33_groupi_n_719);
  or csa_tree_add_6_33_groupi_g16836(csa_tree_add_6_33_groupi_n_1514 ,csa_tree_add_6_33_groupi_n_505 ,csa_tree_add_6_33_groupi_n_784);
  or csa_tree_add_6_33_groupi_g16837(csa_tree_add_6_33_groupi_n_1513 ,csa_tree_add_6_33_groupi_n_487 ,csa_tree_add_6_33_groupi_n_569);
  or csa_tree_add_6_33_groupi_g16838(csa_tree_add_6_33_groupi_n_1512 ,csa_tree_add_6_33_groupi_n_730 ,csa_tree_add_6_33_groupi_n_289);
  or csa_tree_add_6_33_groupi_g16839(csa_tree_add_6_33_groupi_n_1511 ,csa_tree_add_6_33_groupi_n_457 ,csa_tree_add_6_33_groupi_n_712);
  or csa_tree_add_6_33_groupi_g16840(csa_tree_add_6_33_groupi_n_1510 ,csa_tree_add_6_33_groupi_n_68 ,csa_tree_add_6_33_groupi_n_95);
  or csa_tree_add_6_33_groupi_g16841(csa_tree_add_6_33_groupi_n_1509 ,csa_tree_add_6_33_groupi_n_86 ,csa_tree_add_6_33_groupi_n_205);
  or csa_tree_add_6_33_groupi_g16842(csa_tree_add_6_33_groupi_n_1507 ,csa_tree_add_6_33_groupi_n_415 ,csa_tree_add_6_33_groupi_n_461);
  or csa_tree_add_6_33_groupi_g16843(csa_tree_add_6_33_groupi_n_1506 ,csa_tree_add_6_33_groupi_n_373 ,csa_tree_add_6_33_groupi_n_395);
  or csa_tree_add_6_33_groupi_g16844(csa_tree_add_6_33_groupi_n_1505 ,csa_tree_add_6_33_groupi_n_793 ,csa_tree_add_6_33_groupi_n_409);
  or csa_tree_add_6_33_groupi_g16845(csa_tree_add_6_33_groupi_n_1504 ,csa_tree_add_6_33_groupi_n_599 ,csa_tree_add_6_33_groupi_n_74);
  or csa_tree_add_6_33_groupi_g16846(csa_tree_add_6_33_groupi_n_1503 ,csa_tree_add_6_33_groupi_n_805 ,csa_tree_add_6_33_groupi_n_584);
  or csa_tree_add_6_33_groupi_g16847(csa_tree_add_6_33_groupi_n_1502 ,csa_tree_add_6_33_groupi_n_62 ,csa_tree_add_6_33_groupi_n_274);
  or csa_tree_add_6_33_groupi_g16848(csa_tree_add_6_33_groupi_n_1501 ,csa_tree_add_6_33_groupi_n_724 ,csa_tree_add_6_33_groupi_n_637);
  or csa_tree_add_6_33_groupi_g16849(csa_tree_add_6_33_groupi_n_1500 ,csa_tree_add_6_33_groupi_n_527 ,csa_tree_add_6_33_groupi_n_446);
  or csa_tree_add_6_33_groupi_g16850(csa_tree_add_6_33_groupi_n_1499 ,csa_tree_add_6_33_groupi_n_244 ,csa_tree_add_6_33_groupi_n_761);
  or csa_tree_add_6_33_groupi_g16851(csa_tree_add_6_33_groupi_n_1498 ,csa_tree_add_6_33_groupi_n_335 ,csa_tree_add_6_33_groupi_n_716);
  or csa_tree_add_6_33_groupi_g16852(csa_tree_add_6_33_groupi_n_1497 ,csa_tree_add_6_33_groupi_n_365 ,csa_tree_add_6_33_groupi_n_197);
  or csa_tree_add_6_33_groupi_g16853(csa_tree_add_6_33_groupi_n_1496 ,csa_tree_add_6_33_groupi_n_557 ,csa_tree_add_6_33_groupi_n_575);
  or csa_tree_add_6_33_groupi_g16854(csa_tree_add_6_33_groupi_n_1495 ,csa_tree_add_6_33_groupi_n_187 ,csa_tree_add_6_33_groupi_n_119);
  or csa_tree_add_6_33_groupi_g16855(csa_tree_add_6_33_groupi_n_1494 ,csa_tree_add_6_33_groupi_n_737 ,csa_tree_add_6_33_groupi_n_83);
  or csa_tree_add_6_33_groupi_g16856(csa_tree_add_6_33_groupi_n_1493 ,csa_tree_add_6_33_groupi_n_419 ,csa_tree_add_6_33_groupi_n_104);
  or csa_tree_add_6_33_groupi_g16857(csa_tree_add_6_33_groupi_n_1492 ,csa_tree_add_6_33_groupi_n_613 ,csa_tree_add_6_33_groupi_n_631);
  or csa_tree_add_6_33_groupi_g16858(csa_tree_add_6_33_groupi_n_1491 ,csa_tree_add_6_33_groupi_n_413 ,csa_tree_add_6_33_groupi_n_121);
  or csa_tree_add_6_33_groupi_g16859(csa_tree_add_6_33_groupi_n_1490 ,csa_tree_add_6_33_groupi_n_545 ,csa_tree_add_6_33_groupi_n_643);
  or csa_tree_add_6_33_groupi_g16860(csa_tree_add_6_33_groupi_n_1489 ,csa_tree_add_6_33_groupi_n_772 ,csa_tree_add_6_33_groupi_n_59);
  or csa_tree_add_6_33_groupi_g16861(csa_tree_add_6_33_groupi_n_1488 ,csa_tree_add_6_33_groupi_n_787 ,csa_tree_add_6_33_groupi_n_223);
  or csa_tree_add_6_33_groupi_g16862(csa_tree_add_6_33_groupi_n_1487 ,csa_tree_add_6_33_groupi_n_605 ,csa_tree_add_6_33_groupi_n_778);
  or csa_tree_add_6_33_groupi_g16863(csa_tree_add_6_33_groupi_n_1486 ,csa_tree_add_6_33_groupi_n_71 ,csa_tree_add_6_33_groupi_n_578);
  or csa_tree_add_6_33_groupi_g16864(csa_tree_add_6_33_groupi_n_1485 ,csa_tree_add_6_33_groupi_n_503 ,csa_tree_add_6_33_groupi_n_407);
  or csa_tree_add_6_33_groupi_g16865(csa_tree_add_6_33_groupi_n_1484 ,csa_tree_add_6_33_groupi_n_287 ,csa_tree_add_6_33_groupi_n_101);
  or csa_tree_add_6_33_groupi_g16866(csa_tree_add_6_33_groupi_n_1482 ,csa_tree_add_6_33_groupi_n_593 ,csa_tree_add_6_33_groupi_n_560);
  or csa_tree_add_6_33_groupi_g16867(csa_tree_add_6_33_groupi_n_1481 ,csa_tree_add_6_33_groupi_n_539 ,csa_tree_add_6_33_groupi_n_371);
  or csa_tree_add_6_33_groupi_g16868(csa_tree_add_6_33_groupi_n_1480 ,csa_tree_add_6_33_groupi_n_808 ,csa_tree_add_6_33_groupi_n_755);
  or csa_tree_add_6_33_groupi_g16869(csa_tree_add_6_33_groupi_n_1479 ,csa_tree_add_6_33_groupi_n_185 ,csa_tree_add_6_33_groupi_n_485);
  or csa_tree_add_6_33_groupi_g16870(csa_tree_add_6_33_groupi_n_1478 ,csa_tree_add_6_33_groupi_n_473 ,csa_tree_add_6_33_groupi_n_551);
  or csa_tree_add_6_33_groupi_g16871(csa_tree_add_6_33_groupi_n_1477 ,csa_tree_add_6_33_groupi_n_470 ,csa_tree_add_6_33_groupi_n_521);
  or csa_tree_add_6_33_groupi_g16872(csa_tree_add_6_33_groupi_n_1475 ,csa_tree_add_6_33_groupi_n_305 ,csa_tree_add_6_33_groupi_n_764);
  or csa_tree_add_6_33_groupi_g16873(csa_tree_add_6_33_groupi_n_1474 ,csa_tree_add_6_33_groupi_n_802 ,csa_tree_add_6_33_groupi_n_209);
  or csa_tree_add_6_33_groupi_g16874(csa_tree_add_6_33_groupi_n_1473 ,csa_tree_add_6_33_groupi_n_767 ,csa_tree_add_6_33_groupi_n_686);
  or csa_tree_add_6_33_groupi_g16875(csa_tree_add_6_33_groupi_n_1472 ,csa_tree_add_6_33_groupi_n_299 ,csa_tree_add_6_33_groupi_n_173);
  or csa_tree_add_6_33_groupi_g16876(csa_tree_add_6_33_groupi_n_1471 ,csa_tree_add_6_33_groupi_n_731 ,csa_tree_add_6_33_groupi_n_52);
  or csa_tree_add_6_33_groupi_g16877(csa_tree_add_6_33_groupi_n_1470 ,csa_tree_add_6_33_groupi_n_389 ,csa_tree_add_6_33_groupi_n_515);
  or csa_tree_add_6_33_groupi_g16878(csa_tree_add_6_33_groupi_n_1469 ,csa_tree_add_6_33_groupi_n_689 ,csa_tree_add_6_33_groupi_n_416);
  or csa_tree_add_6_33_groupi_g16879(csa_tree_add_6_33_groupi_n_1468 ,csa_tree_add_6_33_groupi_n_56 ,csa_tree_add_6_33_groupi_n_758);
  or csa_tree_add_6_33_groupi_g16880(csa_tree_add_6_33_groupi_n_1467 ,csa_tree_add_6_33_groupi_n_533 ,csa_tree_add_6_33_groupi_n_586);
  or csa_tree_add_6_33_groupi_g16881(csa_tree_add_6_33_groupi_n_1466 ,csa_tree_add_6_33_groupi_n_319 ,csa_tree_add_6_33_groupi_n_218);
  or csa_tree_add_6_33_groupi_g16882(csa_tree_add_6_33_groupi_n_1465 ,csa_tree_add_6_33_groupi_n_437 ,csa_tree_add_6_33_groupi_n_158);
  or csa_tree_add_6_33_groupi_g16883(csa_tree_add_6_33_groupi_n_1464 ,csa_tree_add_6_33_groupi_n_701 ,csa_tree_add_6_33_groupi_n_89);
  or csa_tree_add_6_33_groupi_g16884(csa_tree_add_6_33_groupi_n_1463 ,csa_tree_add_6_33_groupi_n_500 ,csa_tree_add_6_33_groupi_n_179);
  or csa_tree_add_6_33_groupi_g16885(csa_tree_add_6_33_groupi_n_1462 ,csa_tree_add_6_33_groupi_n_347 ,csa_tree_add_6_33_groupi_n_497);
  or csa_tree_add_6_33_groupi_g16886(csa_tree_add_6_33_groupi_n_1461 ,csa_tree_add_6_33_groupi_n_608 ,csa_tree_add_6_33_groupi_n_293);
  or csa_tree_add_6_33_groupi_g16887(csa_tree_add_6_33_groupi_n_1460 ,csa_tree_add_6_33_groupi_n_746 ,csa_tree_add_6_33_groupi_n_398);
  or csa_tree_add_6_33_groupi_g16888(csa_tree_add_6_33_groupi_n_1459 ,csa_tree_add_6_33_groupi_n_242 ,csa_tree_add_6_33_groupi_n_476);
  or csa_tree_add_6_33_groupi_g16889(csa_tree_add_6_33_groupi_n_1458 ,csa_tree_add_6_33_groupi_n_380 ,csa_tree_add_6_33_groupi_n_728);
  or csa_tree_add_6_33_groupi_g16890(csa_tree_add_6_33_groupi_n_1457 ,csa_tree_add_6_33_groupi_n_260 ,csa_tree_add_6_33_groupi_n_140);
  or csa_tree_add_6_33_groupi_g16891(csa_tree_add_6_33_groupi_n_1456 ,csa_tree_add_6_33_groupi_n_317 ,csa_tree_add_6_33_groupi_n_377);
  or csa_tree_add_6_33_groupi_g16892(csa_tree_add_6_33_groupi_n_1455 ,csa_tree_add_6_33_groupi_n_356 ,csa_tree_add_6_33_groupi_n_170);
  or csa_tree_add_6_33_groupi_g16893(csa_tree_add_6_33_groupi_n_1454 ,csa_tree_add_6_33_groupi_n_410 ,csa_tree_add_6_33_groupi_n_752);
  or csa_tree_add_6_33_groupi_g16894(csa_tree_add_6_33_groupi_n_1453 ,csa_tree_add_6_33_groupi_n_596 ,csa_tree_add_6_33_groupi_n_647);
  or csa_tree_add_6_33_groupi_g16895(csa_tree_add_6_33_groupi_n_1452 ,csa_tree_add_6_33_groupi_n_257 ,csa_tree_add_6_33_groupi_n_92);
  or csa_tree_add_6_33_groupi_g16896(csa_tree_add_6_33_groupi_n_1451 ,csa_tree_add_6_33_groupi_n_790 ,csa_tree_add_6_33_groupi_n_680);
  or csa_tree_add_6_33_groupi_g16897(csa_tree_add_6_33_groupi_n_1450 ,csa_tree_add_6_33_groupi_n_200 ,csa_tree_add_6_33_groupi_n_626);
  or csa_tree_add_6_33_groupi_g16898(csa_tree_add_6_33_groupi_n_1449 ,csa_tree_add_6_33_groupi_n_554 ,csa_tree_add_6_33_groupi_n_281);
  or csa_tree_add_6_33_groupi_g16899(csa_tree_add_6_33_groupi_n_1448 ,csa_tree_add_6_33_groupi_n_749 ,csa_tree_add_6_33_groupi_n_662);
  or csa_tree_add_6_33_groupi_g16900(csa_tree_add_6_33_groupi_n_1447 ,csa_tree_add_6_33_groupi_n_602 ,csa_tree_add_6_33_groupi_n_215);
  or csa_tree_add_6_33_groupi_g16901(csa_tree_add_6_33_groupi_n_1446 ,csa_tree_add_6_33_groupi_n_272 ,csa_tree_add_6_33_groupi_n_668);
  or csa_tree_add_6_33_groupi_g16902(csa_tree_add_6_33_groupi_n_1445 ,csa_tree_add_6_33_groupi_n_572 ,csa_tree_add_6_33_groupi_n_491);
  or csa_tree_add_6_33_groupi_g16903(csa_tree_add_6_33_groupi_n_1444 ,csa_tree_add_6_33_groupi_n_176 ,csa_tree_add_6_33_groupi_n_143);
  or csa_tree_add_6_33_groupi_g16904(csa_tree_add_6_33_groupi_n_1443 ,csa_tree_add_6_33_groupi_n_425 ,csa_tree_add_6_33_groupi_n_362);
  or csa_tree_add_6_33_groupi_g16905(csa_tree_add_6_33_groupi_n_1442 ,csa_tree_add_6_33_groupi_n_695 ,csa_tree_add_6_33_groupi_n_350);
  or csa_tree_add_6_33_groupi_g16906(csa_tree_add_6_33_groupi_n_1441 ,csa_tree_add_6_33_groupi_n_811 ,csa_tree_add_6_33_groupi_n_677);
  or csa_tree_add_6_33_groupi_g16907(csa_tree_add_6_33_groupi_n_1440 ,csa_tree_add_6_33_groupi_n_428 ,csa_tree_add_6_33_groupi_n_401);
  or csa_tree_add_6_33_groupi_g16908(csa_tree_add_6_33_groupi_n_1439 ,csa_tree_add_6_33_groupi_n_341 ,csa_tree_add_6_33_groupi_n_26);
  or csa_tree_add_6_33_groupi_g16909(csa_tree_add_6_33_groupi_n_1438 ,csa_tree_add_6_33_groupi_n_251 ,csa_tree_add_6_33_groupi_n_263);
  or csa_tree_add_6_33_groupi_g16910(csa_tree_add_6_33_groupi_n_1437 ,csa_tree_add_6_33_groupi_n_769 ,csa_tree_add_6_33_groupi_n_227);
  or csa_tree_add_6_33_groupi_g16911(csa_tree_add_6_33_groupi_n_1436 ,csa_tree_add_6_33_groupi_n_542 ,csa_tree_add_6_33_groupi_n_131);
  or csa_tree_add_6_33_groupi_g16912(csa_tree_add_6_33_groupi_n_1435 ,csa_tree_add_6_33_groupi_n_329 ,csa_tree_add_6_33_groupi_n_590);
  or csa_tree_add_6_33_groupi_g16913(csa_tree_add_6_33_groupi_n_1434 ,csa_tree_add_6_33_groupi_n_284 ,csa_tree_add_6_33_groupi_n_536);
  or csa_tree_add_6_33_groupi_g16914(csa_tree_add_6_33_groupi_n_1433 ,csa_tree_add_6_33_groupi_n_548 ,csa_tree_add_6_33_groupi_n_332);
  or csa_tree_add_6_33_groupi_g16915(csa_tree_add_6_33_groupi_n_1432 ,csa_tree_add_6_33_groupi_n_149 ,csa_tree_add_6_33_groupi_n_167);
  or csa_tree_add_6_33_groupi_g16916(csa_tree_add_6_33_groupi_n_1431 ,csa_tree_add_6_33_groupi_n_248 ,csa_tree_add_6_33_groupi_n_698);
  or csa_tree_add_6_33_groupi_g16917(csa_tree_add_6_33_groupi_n_1430 ,csa_tree_add_6_33_groupi_n_191 ,csa_tree_add_6_33_groupi_n_47);
  or csa_tree_add_6_33_groupi_g16918(csa_tree_add_6_33_groupi_n_1429 ,csa_tree_add_6_33_groupi_n_155 ,csa_tree_add_6_33_groupi_n_580);
  or csa_tree_add_6_33_groupi_g16919(csa_tree_add_6_33_groupi_n_1428 ,csa_tree_add_6_33_groupi_n_278 ,csa_tree_add_6_33_groupi_n_392);
  or csa_tree_add_6_33_groupi_g16920(csa_tree_add_6_33_groupi_n_1427 ,csa_tree_add_6_33_groupi_n_641 ,csa_tree_add_6_33_groupi_n_368);
  or csa_tree_add_6_33_groupi_g16921(csa_tree_add_6_33_groupi_n_1426 ,csa_tree_add_6_33_groupi_n_374 ,csa_tree_add_6_33_groupi_n_653);
  or csa_tree_add_6_33_groupi_g16922(csa_tree_add_6_33_groupi_n_1425 ,csa_tree_add_6_33_groupi_n_734 ,csa_tree_add_6_33_groupi_n_674);
  or csa_tree_add_6_33_groupi_g16923(csa_tree_add_6_33_groupi_n_1423 ,csa_tree_add_6_33_groupi_n_152 ,csa_tree_add_6_33_groupi_n_623);
  or csa_tree_add_6_33_groupi_g16924(csa_tree_add_6_33_groupi_n_1422 ,csa_tree_add_6_33_groupi_n_239 ,csa_tree_add_6_33_groupi_n_220);
  or csa_tree_add_6_33_groupi_g16925(csa_tree_add_6_33_groupi_n_1421 ,csa_tree_add_6_33_groupi_n_482 ,csa_tree_add_6_33_groupi_n_562);
  or csa_tree_add_6_33_groupi_g16926(csa_tree_add_6_33_groupi_n_1420 ,csa_tree_add_6_33_groupi_n_635 ,csa_tree_add_6_33_groupi_n_518);
  or csa_tree_add_6_33_groupi_g16927(csa_tree_add_6_33_groupi_n_1419 ,csa_tree_add_6_33_groupi_n_146 ,csa_tree_add_6_33_groupi_n_290);
  or csa_tree_add_6_33_groupi_g16928(csa_tree_add_6_33_groupi_n_1418 ,csa_tree_add_6_33_groupi_n_434 ,csa_tree_add_6_33_groupi_n_106);
  or csa_tree_add_6_33_groupi_g16929(csa_tree_add_6_33_groupi_n_1417 ,csa_tree_add_6_33_groupi_n_683 ,csa_tree_add_6_33_groupi_n_24);
  or csa_tree_add_6_33_groupi_g16930(csa_tree_add_6_33_groupi_n_1416 ,csa_tree_add_6_33_groupi_n_458 ,csa_tree_add_6_33_groupi_n_131);
  or csa_tree_add_6_33_groupi_g16931(csa_tree_add_6_33_groupi_n_1415 ,csa_tree_add_6_33_groupi_n_36 ,csa_tree_add_6_33_groupi_n_478);
  and csa_tree_add_6_33_groupi_g16932(csa_tree_add_6_33_groupi_n_1413 ,in1[4] ,in1[3]);
  or csa_tree_add_6_33_groupi_g16933(csa_tree_add_6_33_groupi_n_1412 ,csa_tree_add_6_33_groupi_n_224 ,csa_tree_add_6_33_groupi_n_743);
  or csa_tree_add_6_33_groupi_g16934(csa_tree_add_6_33_groupi_n_1411 ,csa_tree_add_6_33_groupi_n_509 ,csa_tree_add_6_33_groupi_n_704);
  or csa_tree_add_6_33_groupi_g16935(csa_tree_add_6_33_groupi_n_1410 ,csa_tree_add_6_33_groupi_n_655 ,csa_tree_add_6_33_groupi_n_103);
  or csa_tree_add_6_33_groupi_g16936(csa_tree_add_6_33_groupi_n_1408 ,csa_tree_add_6_33_groupi_n_82 ,csa_tree_add_6_33_groupi_n_659);
  or csa_tree_add_6_33_groupi_g16937(csa_tree_add_6_33_groupi_n_1407 ,csa_tree_add_6_33_groupi_n_524 ,csa_tree_add_6_33_groupi_n_40);
  or csa_tree_add_6_33_groupi_g16938(csa_tree_add_6_33_groupi_n_1406 ,csa_tree_add_6_33_groupi_n_449 ,csa_tree_add_6_33_groupi_n_422);
  or csa_tree_add_6_33_groupi_g16939(csa_tree_add_6_33_groupi_n_1405 ,csa_tree_add_6_33_groupi_n_296 ,csa_tree_add_6_33_groupi_n_235);
  or csa_tree_add_6_33_groupi_g16940(csa_tree_add_6_33_groupi_n_1404 ,csa_tree_add_6_33_groupi_n_28 ,csa_tree_add_6_33_groupi_n_494);
  or csa_tree_add_6_33_groupi_g16941(csa_tree_add_6_33_groupi_n_1403 ,csa_tree_add_6_33_groupi_n_431 ,csa_tree_add_6_33_groupi_n_670);
  or csa_tree_add_6_33_groupi_g16942(csa_tree_add_6_33_groupi_n_1402 ,csa_tree_add_6_33_groupi_n_182 ,csa_tree_add_6_33_groupi_n_73);
  or csa_tree_add_6_33_groupi_g16943(csa_tree_add_6_33_groupi_n_1401 ,csa_tree_add_6_33_groupi_n_137 ,csa_tree_add_6_33_groupi_n_488);
  or csa_tree_add_6_33_groupi_g16944(csa_tree_add_6_33_groupi_n_1400 ,csa_tree_add_6_33_groupi_n_308 ,csa_tree_add_6_33_groupi_n_512);
  or csa_tree_add_6_33_groupi_g16945(csa_tree_add_6_33_groupi_n_1398 ,csa_tree_add_6_33_groupi_n_725 ,csa_tree_add_6_33_groupi_n_692);
  and csa_tree_add_6_33_groupi_g16946(csa_tree_add_6_33_groupi_n_1397 ,in1[30] ,in1[27]);
  or csa_tree_add_6_33_groupi_g16947(csa_tree_add_6_33_groupi_n_1395 ,csa_tree_add_6_33_groupi_n_323 ,csa_tree_add_6_33_groupi_n_127);
  or csa_tree_add_6_33_groupi_g16948(csa_tree_add_6_33_groupi_n_1394 ,csa_tree_add_6_33_groupi_n_556 ,csa_tree_add_6_33_groupi_n_353);
  or csa_tree_add_6_33_groupi_g16949(csa_tree_add_6_33_groupi_n_1393 ,csa_tree_add_6_33_groupi_n_160 ,csa_tree_add_6_33_groupi_n_85);
  or csa_tree_add_6_33_groupi_g16950(csa_tree_add_6_33_groupi_n_1392 ,csa_tree_add_6_33_groupi_n_42 ,csa_tree_add_6_33_groupi_n_61);
  or csa_tree_add_6_33_groupi_g16951(csa_tree_add_6_33_groupi_n_1391 ,csa_tree_add_6_33_groupi_n_286 ,csa_tree_add_6_33_groupi_n_610);
  or csa_tree_add_6_33_groupi_g16952(csa_tree_add_6_33_groupi_n_1390 ,csa_tree_add_6_33_groupi_n_502 ,csa_tree_add_6_33_groupi_n_394);
  or csa_tree_add_6_33_groupi_g16953(csa_tree_add_6_33_groupi_n_1389 ,csa_tree_add_6_33_groupi_n_544 ,csa_tree_add_6_33_groupi_n_404);
  or csa_tree_add_6_33_groupi_g16954(csa_tree_add_6_33_groupi_n_1388 ,csa_tree_add_6_33_groupi_n_484 ,csa_tree_add_6_33_groupi_n_617);
  or csa_tree_add_6_33_groupi_g16955(csa_tree_add_6_33_groupi_n_1387 ,csa_tree_add_6_33_groupi_n_598 ,csa_tree_add_6_33_groupi_n_382);
  or csa_tree_add_6_33_groupi_g16956(csa_tree_add_6_33_groupi_n_1386 ,csa_tree_add_6_33_groupi_n_566 ,csa_tree_add_6_33_groupi_n_109);
  or csa_tree_add_6_33_groupi_g16957(csa_tree_add_6_33_groupi_n_1385 ,csa_tree_add_6_33_groupi_n_526 ,csa_tree_add_6_33_groupi_n_301);
  or csa_tree_add_6_33_groupi_g16958(csa_tree_add_6_33_groupi_n_1384 ,csa_tree_add_6_33_groupi_n_475 ,csa_tree_add_6_33_groupi_n_212);
  or csa_tree_add_6_33_groupi_g16959(csa_tree_add_6_33_groupi_n_1383 ,csa_tree_add_6_33_groupi_n_604 ,csa_tree_add_6_33_groupi_n_266);
  or csa_tree_add_6_33_groupi_g16960(csa_tree_add_6_33_groupi_n_1382 ,csa_tree_add_6_33_groupi_n_164 ,csa_tree_add_6_33_groupi_n_467);
  or csa_tree_add_6_33_groupi_g16961(csa_tree_add_6_33_groupi_n_1381 ,csa_tree_add_6_33_groupi_n_386 ,csa_tree_add_6_33_groupi_n_667);
  or csa_tree_add_6_33_groupi_g16962(csa_tree_add_6_33_groupi_n_1380 ,csa_tree_add_6_33_groupi_n_812 ,csa_tree_add_6_33_groupi_n_443);
  or csa_tree_add_6_33_groupi_g16963(csa_tree_add_6_33_groupi_n_1379 ,csa_tree_add_6_33_groupi_n_188 ,csa_tree_add_6_33_groupi_n_721);
  or csa_tree_add_6_33_groupi_g16964(csa_tree_add_6_33_groupi_n_1378 ,csa_tree_add_6_33_groupi_n_592 ,csa_tree_add_6_33_groupi_n_715);
  or csa_tree_add_6_33_groupi_g16965(csa_tree_add_6_33_groupi_n_1377 ,csa_tree_add_6_33_groupi_n_452 ,csa_tree_add_6_33_groupi_n_650);
  or csa_tree_add_6_33_groupi_g16966(csa_tree_add_6_33_groupi_n_1376 ,csa_tree_add_6_33_groupi_n_230 ,csa_tree_add_6_33_groupi_n_455);
  or csa_tree_add_6_33_groupi_g16967(csa_tree_add_6_33_groupi_n_1374 ,csa_tree_add_6_33_groupi_n_530 ,csa_tree_add_6_33_groupi_n_628);
  or csa_tree_add_6_33_groupi_g16968(csa_tree_add_6_33_groupi_n_1373 ,csa_tree_add_6_33_groupi_n_707 ,csa_tree_add_6_33_groupi_n_67);
  or csa_tree_add_6_33_groupi_g16969(csa_tree_add_6_33_groupi_n_1372 ,csa_tree_add_6_33_groupi_n_506 ,csa_tree_add_6_33_groupi_n_472);
  or csa_tree_add_6_33_groupi_g16970(csa_tree_add_6_33_groupi_n_1371 ,csa_tree_add_6_33_groupi_n_157 ,csa_tree_add_6_33_groupi_n_574);
  or csa_tree_add_6_33_groupi_g16971(csa_tree_add_6_33_groupi_n_1370 ,csa_tree_add_6_33_groupi_n_769 ,csa_tree_add_6_33_groupi_n_32);
  or csa_tree_add_6_33_groupi_g16972(csa_tree_add_6_33_groupi_n_1369 ,csa_tree_add_6_33_groupi_n_271 ,csa_tree_add_6_33_groupi_n_550);
  or csa_tree_add_6_33_groupi_g16973(csa_tree_add_6_33_groupi_n_1368 ,csa_tree_add_6_33_groupi_n_766 ,csa_tree_add_6_33_groupi_n_194);
  or csa_tree_add_6_33_groupi_g16974(csa_tree_add_6_33_groupi_n_1367 ,csa_tree_add_6_33_groupi_n_259 ,csa_tree_add_6_33_groupi_n_520);
  or csa_tree_add_6_33_groupi_g16975(csa_tree_add_6_33_groupi_n_1366 ,csa_tree_add_6_33_groupi_n_538 ,csa_tree_add_6_33_groupi_n_440);
  or csa_tree_add_6_33_groupi_g16976(csa_tree_add_6_33_groupi_n_1365 ,csa_tree_add_6_33_groupi_n_245 ,csa_tree_add_6_33_groupi_n_34);
  or csa_tree_add_6_33_groupi_g16977(csa_tree_add_6_33_groupi_n_1364 ,csa_tree_add_6_33_groupi_n_682 ,csa_tree_add_6_33_groupi_n_644);
  not csa_tree_add_6_33_groupi_g16978(csa_tree_add_6_33_groupi_n_1210 ,csa_tree_add_6_33_groupi_n_1209);
  not csa_tree_add_6_33_groupi_g16979(csa_tree_add_6_33_groupi_n_1161 ,csa_tree_add_6_33_groupi_n_1160);
  not csa_tree_add_6_33_groupi_g16980(csa_tree_add_6_33_groupi_n_1143 ,csa_tree_add_6_33_groupi_n_1142);
  not csa_tree_add_6_33_groupi_g16981(csa_tree_add_6_33_groupi_n_1138 ,csa_tree_add_6_33_groupi_n_1137);
  not csa_tree_add_6_33_groupi_g16982(csa_tree_add_6_33_groupi_n_1134 ,csa_tree_add_6_33_groupi_n_1133);
  not csa_tree_add_6_33_groupi_g16983(csa_tree_add_6_33_groupi_n_1107 ,csa_tree_add_6_33_groupi_n_1106);
  nand csa_tree_add_6_33_groupi_g16984(csa_tree_add_6_33_groupi_n_1069 ,in3[27] ,in2[27]);
  and csa_tree_add_6_33_groupi_g16985(csa_tree_add_6_33_groupi_n_1068 ,in1[1] ,in3[2]);
  nand csa_tree_add_6_33_groupi_g16986(csa_tree_add_6_33_groupi_n_1067 ,in3[25] ,in2[25]);
  nand csa_tree_add_6_33_groupi_g16987(csa_tree_add_6_33_groupi_n_1066 ,in3[21] ,in2[21]);
  nor csa_tree_add_6_33_groupi_g16988(csa_tree_add_6_33_groupi_n_1065 ,in3[13] ,in2[13]);
  or csa_tree_add_6_33_groupi_g16989(csa_tree_add_6_33_groupi_n_1064 ,in1[2] ,in2[4]);
  and csa_tree_add_6_33_groupi_g16990(csa_tree_add_6_33_groupi_n_1063 ,in1[12] ,in3[24]);
  nand csa_tree_add_6_33_groupi_g16991(csa_tree_add_6_33_groupi_n_1062 ,in3[17] ,in2[17]);
  nor csa_tree_add_6_33_groupi_g16992(csa_tree_add_6_33_groupi_n_1061 ,in3[29] ,in2[29]);
  or csa_tree_add_6_33_groupi_g16993(csa_tree_add_6_33_groupi_n_1060 ,in1[12] ,in3[24]);
  nor csa_tree_add_6_33_groupi_g16994(csa_tree_add_6_33_groupi_n_1059 ,in3[25] ,in2[25]);
  and csa_tree_add_6_33_groupi_g16995(csa_tree_add_6_33_groupi_n_1058 ,in3[6] ,in2[6]);
  nor csa_tree_add_6_33_groupi_g16996(csa_tree_add_6_33_groupi_n_1057 ,in3[21] ,in2[21]);
  nor csa_tree_add_6_33_groupi_g16997(csa_tree_add_6_33_groupi_n_1056 ,in3[6] ,in2[6]);
  or csa_tree_add_6_33_groupi_g16998(csa_tree_add_6_33_groupi_n_1055 ,in1[9] ,in3[18]);
  nand csa_tree_add_6_33_groupi_g16999(csa_tree_add_6_33_groupi_n_1054 ,in3[19] ,in2[19]);
  and csa_tree_add_6_33_groupi_g17000(csa_tree_add_6_33_groupi_n_1053 ,in1[15] ,in3[30]);
  and csa_tree_add_6_33_groupi_g17001(csa_tree_add_6_33_groupi_n_1052 ,in1[6] ,in3[12]);
  and csa_tree_add_6_33_groupi_g17002(csa_tree_add_6_33_groupi_n_1051 ,in1[5] ,in3[10]);
  and csa_tree_add_6_33_groupi_g17003(csa_tree_add_6_33_groupi_n_1050 ,in1[10] ,in3[20]);
  and csa_tree_add_6_33_groupi_g17004(csa_tree_add_6_33_groupi_n_1049 ,in1[9] ,in3[18]);
  and csa_tree_add_6_33_groupi_g17005(csa_tree_add_6_33_groupi_n_1048 ,in1[14] ,in3[28]);
  and csa_tree_add_6_33_groupi_g17006(csa_tree_add_6_33_groupi_n_1047 ,in3[8] ,in2[8]);
  nand csa_tree_add_6_33_groupi_g17007(csa_tree_add_6_33_groupi_n_1046 ,in3[5] ,in2[5]);
  and csa_tree_add_6_33_groupi_g17008(csa_tree_add_6_33_groupi_n_1045 ,in1[13] ,in3[26]);
  or csa_tree_add_6_33_groupi_g17009(csa_tree_add_6_33_groupi_n_1044 ,csa_tree_add_6_33_groupi_n_358 ,csa_tree_add_6_33_groupi_n_1041);
  nor csa_tree_add_6_33_groupi_g17010(csa_tree_add_6_33_groupi_n_1043 ,in3[17] ,in2[17]);
  nor csa_tree_add_6_33_groupi_g17011(csa_tree_add_6_33_groupi_n_1042 ,in3[1] ,in2[1]);
  or csa_tree_add_6_33_groupi_g17012(csa_tree_add_6_33_groupi_n_1327 ,csa_tree_add_6_33_groupi_n_754 ,csa_tree_add_6_33_groupi_n_620);
  or csa_tree_add_6_33_groupi_g17013(csa_tree_add_6_33_groupi_n_1326 ,csa_tree_add_6_33_groupi_n_344 ,csa_tree_add_6_33_groupi_n_418);
  or csa_tree_add_6_33_groupi_g17014(csa_tree_add_6_33_groupi_n_1325 ,csa_tree_add_6_33_groupi_n_595 ,csa_tree_add_6_33_groupi_n_124);
  or csa_tree_add_6_33_groupi_g17015(csa_tree_add_6_33_groupi_n_1324 ,csa_tree_add_6_33_groupi_n_30 ,csa_tree_add_6_33_groupi_n_310);
  or csa_tree_add_6_33_groupi_g17016(csa_tree_add_6_33_groupi_n_1323 ,csa_tree_add_6_33_groupi_n_154 ,csa_tree_add_6_33_groupi_n_79);
  or csa_tree_add_6_33_groupi_g17017(csa_tree_add_6_33_groupi_n_1322 ,csa_tree_add_6_33_groupi_n_638 ,csa_tree_add_6_33_groupi_n_233);
  or csa_tree_add_6_33_groupi_g17018(csa_tree_add_6_33_groupi_n_1321 ,csa_tree_add_6_33_groupi_n_523 ,csa_tree_add_6_33_groupi_n_583);
  or csa_tree_add_6_33_groupi_g17019(csa_tree_add_6_33_groupi_n_1320 ,csa_tree_add_6_33_groupi_n_304 ,csa_tree_add_6_33_groupi_n_133);
  or csa_tree_add_6_33_groupi_g17020(csa_tree_add_6_33_groupi_n_1319 ,csa_tree_add_6_33_groupi_n_181 ,csa_tree_add_6_33_groupi_n_694);
  or csa_tree_add_6_33_groupi_g17021(csa_tree_add_6_33_groupi_n_1318 ,csa_tree_add_6_33_groupi_n_424 ,csa_tree_add_6_33_groupi_n_196);
  or csa_tree_add_6_33_groupi_g17022(csa_tree_add_6_33_groupi_n_1317 ,csa_tree_add_6_33_groupi_n_202 ,csa_tree_add_6_33_groupi_n_736);
  or csa_tree_add_6_33_groupi_g17023(csa_tree_add_6_33_groupi_n_1316 ,csa_tree_add_6_33_groupi_n_64 ,csa_tree_add_6_33_groupi_n_763);
  or csa_tree_add_6_33_groupi_g17024(csa_tree_add_6_33_groupi_n_1315 ,csa_tree_add_6_33_groupi_n_254 ,csa_tree_add_6_33_groupi_n_275);
  or csa_tree_add_6_33_groupi_g17025(csa_tree_add_6_33_groupi_n_1314 ,csa_tree_add_6_33_groupi_n_184 ,csa_tree_add_6_33_groupi_n_710);
  or csa_tree_add_6_33_groupi_g17026(csa_tree_add_6_33_groupi_n_1313 ,csa_tree_add_6_33_groupi_n_607 ,csa_tree_add_6_33_groupi_n_614);
  or csa_tree_add_6_33_groupi_g17027(csa_tree_add_6_33_groupi_n_1312 ,csa_tree_add_6_33_groupi_n_412 ,csa_tree_add_6_33_groupi_n_97);
  or csa_tree_add_6_33_groupi_g17028(csa_tree_add_6_33_groupi_n_1311 ,csa_tree_add_6_33_groupi_n_601 ,csa_tree_add_6_33_groupi_n_376);
  or csa_tree_add_6_33_groupi_g17029(csa_tree_add_6_33_groupi_n_1310 ,csa_tree_add_6_33_groupi_n_18 ,csa_tree_add_6_33_groupi_n_238);
  or csa_tree_add_6_33_groupi_g17030(csa_tree_add_6_33_groupi_n_1309 ,csa_tree_add_6_33_groupi_n_22 ,csa_tree_add_6_33_groupi_n_169);
  or csa_tree_add_6_33_groupi_g17031(csa_tree_add_6_33_groupi_n_1308 ,csa_tree_add_6_33_groupi_n_226 ,csa_tree_add_6_33_groupi_n_665);
  or csa_tree_add_6_33_groupi_g17032(csa_tree_add_6_33_groupi_n_1307 ,csa_tree_add_6_33_groupi_n_496 ,csa_tree_add_6_33_groupi_n_206);
  or csa_tree_add_6_33_groupi_g17033(csa_tree_add_6_33_groupi_n_1306 ,csa_tree_add_6_33_groupi_n_338 ,csa_tree_add_6_33_groupi_n_118);
  or csa_tree_add_6_33_groupi_g17034(csa_tree_add_6_33_groupi_n_1305 ,csa_tree_add_6_33_groupi_n_70 ,csa_tree_add_6_33_groupi_n_364);
  or csa_tree_add_6_33_groupi_g17035(csa_tree_add_6_33_groupi_n_1304 ,csa_tree_add_6_33_groupi_n_589 ,csa_tree_add_6_33_groupi_n_718);
  or csa_tree_add_6_33_groupi_g17036(csa_tree_add_6_33_groupi_n_1303 ,csa_tree_add_6_33_groupi_n_532 ,csa_tree_add_6_33_groupi_n_490);
  or csa_tree_add_6_33_groupi_g17037(csa_tree_add_6_33_groupi_n_1302 ,csa_tree_add_6_33_groupi_n_326 ,csa_tree_add_6_33_groupi_n_661);
  or csa_tree_add_6_33_groupi_g17038(csa_tree_add_6_33_groupi_n_1301 ,csa_tree_add_6_33_groupi_n_320 ,csa_tree_add_6_33_groupi_n_370);
  or csa_tree_add_6_33_groupi_g17039(csa_tree_add_6_33_groupi_n_1300 ,csa_tree_add_6_33_groupi_n_136 ,csa_tree_add_6_33_groupi_n_713);
  or csa_tree_add_6_33_groupi_g17040(csa_tree_add_6_33_groupi_n_1299 ,csa_tree_add_6_33_groupi_n_241 ,csa_tree_add_6_33_groupi_n_100);
  or csa_tree_add_6_33_groupi_g17041(csa_tree_add_6_33_groupi_n_1298 ,csa_tree_add_6_33_groupi_n_553 ,csa_tree_add_6_33_groupi_n_94);
  or csa_tree_add_6_33_groupi_g17042(csa_tree_add_6_33_groupi_n_1297 ,csa_tree_add_6_33_groupi_n_178 ,csa_tree_add_6_33_groupi_n_760);
  or csa_tree_add_6_33_groupi_g17043(csa_tree_add_6_33_groupi_n_1296 ,csa_tree_add_6_33_groupi_n_508 ,csa_tree_add_6_33_groupi_n_464);
  or csa_tree_add_6_33_groupi_g17044(csa_tree_add_6_33_groupi_n_1295 ,csa_tree_add_6_33_groupi_n_314 ,csa_tree_add_6_33_groupi_n_290);
  or csa_tree_add_6_33_groupi_g17045(csa_tree_add_6_33_groupi_n_1294 ,csa_tree_add_6_33_groupi_n_676 ,csa_tree_add_6_33_groupi_n_269);
  or csa_tree_add_6_33_groupi_g17046(csa_tree_add_6_33_groupi_n_1293 ,csa_tree_add_6_33_groupi_n_112 ,csa_tree_add_6_33_groupi_n_514);
  or csa_tree_add_6_33_groupi_g17047(csa_tree_add_6_33_groupi_n_1292 ,csa_tree_add_6_33_groupi_n_781 ,csa_tree_add_6_33_groupi_n_208);
  or csa_tree_add_6_33_groupi_g17048(csa_tree_add_6_33_groupi_n_1291 ,csa_tree_add_6_33_groupi_n_611 ,csa_tree_add_6_33_groupi_n_76);
  or csa_tree_add_6_33_groupi_g17049(csa_tree_add_6_33_groupi_n_1290 ,csa_tree_add_6_33_groupi_n_430 ,csa_tree_add_6_33_groupi_n_757);
  or csa_tree_add_6_33_groupi_g17050(csa_tree_add_6_33_groupi_n_1289 ,csa_tree_add_6_33_groupi_n_632 ,csa_tree_add_6_33_groupi_n_172);
  or csa_tree_add_6_33_groupi_g17051(csa_tree_add_6_33_groupi_n_1288 ,csa_tree_add_6_33_groupi_n_625 ,csa_tree_add_6_33_groupi_n_751);
  or csa_tree_add_6_33_groupi_g17052(csa_tree_add_6_33_groupi_n_1287 ,csa_tree_add_6_33_groupi_n_724 ,csa_tree_add_6_33_groupi_n_256);
  or csa_tree_add_6_33_groupi_g17053(csa_tree_add_6_33_groupi_n_1286 ,csa_tree_add_6_33_groupi_n_565 ,csa_tree_add_6_33_groupi_n_91);
  or csa_tree_add_6_33_groupi_g17054(csa_tree_add_6_33_groupi_n_1285 ,csa_tree_add_6_33_groupi_n_541 ,csa_tree_add_6_33_groupi_n_298);
  or csa_tree_add_6_33_groupi_g17055(csa_tree_add_6_33_groupi_n_1284 ,csa_tree_add_6_33_groupi_n_796 ,csa_tree_add_6_33_groupi_n_460);
  or csa_tree_add_6_33_groupi_g17056(csa_tree_add_6_33_groupi_n_1283 ,csa_tree_add_6_33_groupi_n_703 ,csa_tree_add_6_33_groupi_n_49);
  or csa_tree_add_6_33_groupi_g17057(csa_tree_add_6_33_groupi_n_1282 ,csa_tree_add_6_33_groupi_n_685 ,csa_tree_add_6_33_groupi_n_214);
  or csa_tree_add_6_33_groupi_g17058(csa_tree_add_6_33_groupi_n_1281 ,csa_tree_add_6_33_groupi_n_397 ,csa_tree_add_6_33_groupi_n_646);
  or csa_tree_add_6_33_groupi_g17059(csa_tree_add_6_33_groupi_n_1280 ,csa_tree_add_6_33_groupi_n_688 ,csa_tree_add_6_33_groupi_n_605);
  or csa_tree_add_6_33_groupi_g17060(csa_tree_add_6_33_groupi_n_1279 ,csa_tree_add_6_33_groupi_n_38 ,csa_tree_add_6_33_groupi_n_406);
  or csa_tree_add_6_33_groupi_g17061(csa_tree_add_6_33_groupi_n_1278 ,csa_tree_add_6_33_groupi_n_217 ,csa_tree_add_6_33_groupi_n_427);
  or csa_tree_add_6_33_groupi_g17062(csa_tree_add_6_33_groupi_n_1277 ,csa_tree_add_6_33_groupi_n_640 ,csa_tree_add_6_33_groupi_n_568);
  or csa_tree_add_6_33_groupi_g17063(csa_tree_add_6_33_groupi_n_1276 ,csa_tree_add_6_33_groupi_n_199 ,csa_tree_add_6_33_groupi_n_469);
  or csa_tree_add_6_33_groupi_g17064(csa_tree_add_6_33_groupi_n_1275 ,csa_tree_add_6_33_groupi_n_388 ,csa_tree_add_6_33_groupi_n_265);
  or csa_tree_add_6_33_groupi_g17065(csa_tree_add_6_33_groupi_n_1274 ,csa_tree_add_6_33_groupi_n_139 ,csa_tree_add_6_33_groupi_n_577);
  or csa_tree_add_6_33_groupi_g17066(csa_tree_add_6_33_groupi_n_1273 ,csa_tree_add_6_33_groupi_n_535 ,csa_tree_add_6_33_groupi_n_262);
  or csa_tree_add_6_33_groupi_g17067(csa_tree_add_6_33_groupi_n_1272 ,csa_tree_add_6_33_groupi_n_436 ,csa_tree_add_6_33_groupi_n_748);
  or csa_tree_add_6_33_groupi_g17068(csa_tree_add_6_33_groupi_n_1271 ,csa_tree_add_6_33_groupi_n_20 ,csa_tree_add_6_33_groupi_n_379);
  or csa_tree_add_6_33_groupi_g17069(csa_tree_add_6_33_groupi_n_1270 ,csa_tree_add_6_33_groupi_n_55 ,csa_tree_add_6_33_groupi_n_391);
  or csa_tree_add_6_33_groupi_g17070(csa_tree_add_6_33_groupi_n_1269 ,csa_tree_add_6_33_groupi_n_175 ,csa_tree_add_6_33_groupi_n_559);
  or csa_tree_add_6_33_groupi_g17071(csa_tree_add_6_33_groupi_n_1268 ,csa_tree_add_6_33_groupi_n_499 ,csa_tree_add_6_33_groupi_n_361);
  or csa_tree_add_6_33_groupi_g17072(csa_tree_add_6_33_groupi_n_1267 ,csa_tree_add_6_33_groupi_n_448 ,csa_tree_add_6_33_groupi_n_634);
  or csa_tree_add_6_33_groupi_g17073(csa_tree_add_6_33_groupi_n_1266 ,csa_tree_add_6_33_groupi_n_527 ,csa_tree_add_6_33_groupi_n_517);
  or csa_tree_add_6_33_groupi_g17074(csa_tree_add_6_33_groupi_n_1265 ,csa_tree_add_6_33_groupi_n_283 ,csa_tree_add_6_33_groupi_n_481);
  or csa_tree_add_6_33_groupi_g17075(csa_tree_add_6_33_groupi_n_1264 ,csa_tree_add_6_33_groupi_n_403 ,csa_tree_add_6_33_groupi_n_400);
  or csa_tree_add_6_33_groupi_g17076(csa_tree_add_6_33_groupi_n_1263 ,csa_tree_add_6_33_groupi_n_346 ,csa_tree_add_6_33_groupi_n_529);
  or csa_tree_add_6_33_groupi_g17077(csa_tree_add_6_33_groupi_n_1262 ,csa_tree_add_6_33_groupi_n_292 ,csa_tree_add_6_33_groupi_n_53);
  or csa_tree_add_6_33_groupi_g17078(csa_tree_add_6_33_groupi_n_1261 ,csa_tree_add_6_33_groupi_n_571 ,csa_tree_add_6_33_groupi_n_145);
  or csa_tree_add_6_33_groupi_g17079(csa_tree_add_6_33_groupi_n_1260 ,csa_tree_add_6_33_groupi_n_775 ,csa_tree_add_6_33_groupi_n_190);
  or csa_tree_add_6_33_groupi_g17080(csa_tree_add_6_33_groupi_n_1259 ,csa_tree_add_6_33_groupi_n_593 ,csa_tree_add_6_33_groupi_n_166);
  or csa_tree_add_6_33_groupi_g17081(csa_tree_add_6_33_groupi_n_1258 ,csa_tree_add_6_33_groupi_n_340 ,csa_tree_add_6_33_groupi_n_355);
  or csa_tree_add_6_33_groupi_g17082(csa_tree_add_6_33_groupi_n_1257 ,csa_tree_add_6_33_groupi_n_742 ,csa_tree_add_6_33_groupi_n_236);
  or csa_tree_add_6_33_groupi_g17083(csa_tree_add_6_33_groupi_n_1256 ,csa_tree_add_6_33_groupi_n_730 ,csa_tree_add_6_33_groupi_n_445);
  or csa_tree_add_6_33_groupi_g17084(csa_tree_add_6_33_groupi_n_1255 ,csa_tree_add_6_33_groupi_n_793 ,csa_tree_add_6_33_groupi_n_247);
  or csa_tree_add_6_33_groupi_g17085(csa_tree_add_6_33_groupi_n_1254 ,csa_tree_add_6_33_groupi_n_277 ,csa_tree_add_6_33_groupi_n_616);
  or csa_tree_add_6_33_groupi_g17086(csa_tree_add_6_33_groupi_n_1253 ,csa_tree_add_6_33_groupi_n_421 ,csa_tree_add_6_33_groupi_n_367);
  or csa_tree_add_6_33_groupi_g17087(csa_tree_add_6_33_groupi_n_1252 ,csa_tree_add_6_33_groupi_n_433 ,csa_tree_add_6_33_groupi_n_232);
  or csa_tree_add_6_33_groupi_g17088(csa_tree_add_6_33_groupi_n_1251 ,csa_tree_add_6_33_groupi_n_511 ,csa_tree_add_6_33_groupi_n_740);
  or csa_tree_add_6_33_groupi_g17089(csa_tree_add_6_33_groupi_n_1250 ,csa_tree_add_6_33_groupi_n_439 ,csa_tree_add_6_33_groupi_n_700);
  or csa_tree_add_6_33_groupi_g17090(csa_tree_add_6_33_groupi_n_1249 ,csa_tree_add_6_33_groupi_n_547 ,csa_tree_add_6_33_groupi_n_142);
  or csa_tree_add_6_33_groupi_g17091(csa_tree_add_6_33_groupi_n_1248 ,csa_tree_add_6_33_groupi_n_415 ,csa_tree_add_6_33_groupi_n_493);
  or csa_tree_add_6_33_groupi_g17092(csa_tree_add_6_33_groupi_n_1247 ,csa_tree_add_6_33_groupi_n_385 ,csa_tree_add_6_33_groupi_n_373);
  or csa_tree_add_6_33_groupi_g17093(csa_tree_add_6_33_groupi_n_1246 ,csa_tree_add_6_33_groupi_n_451 ,csa_tree_add_6_33_groupi_n_409);
  or csa_tree_add_6_33_groupi_g17094(csa_tree_add_6_33_groupi_n_1245 ,csa_tree_add_6_33_groupi_n_811 ,csa_tree_add_6_33_groupi_n_328);
  or csa_tree_add_6_33_groupi_g17095(csa_tree_add_6_33_groupi_n_1244 ,csa_tree_add_6_33_groupi_n_163 ,csa_tree_add_6_33_groupi_n_86);
  or csa_tree_add_6_33_groupi_g17096(csa_tree_add_6_33_groupi_n_1243 ,csa_tree_add_6_33_groupi_n_673 ,csa_tree_add_6_33_groupi_n_622);
  or csa_tree_add_6_33_groupi_g17097(csa_tree_add_6_33_groupi_n_1242 ,csa_tree_add_6_33_groupi_n_134 ,csa_tree_add_6_33_groupi_n_395);
  or csa_tree_add_6_33_groupi_g17098(csa_tree_add_6_33_groupi_n_1241 ,csa_tree_add_6_33_groupi_n_137 ,csa_tree_add_6_33_groupi_n_130);
  or csa_tree_add_6_33_groupi_g17099(csa_tree_add_6_33_groupi_n_1240 ,csa_tree_add_6_33_groupi_n_706 ,csa_tree_add_6_33_groupi_n_521);
  or csa_tree_add_6_33_groupi_g17100(csa_tree_add_6_33_groupi_n_1239 ,csa_tree_add_6_33_groupi_n_505 ,csa_tree_add_6_33_groupi_n_799);
  or csa_tree_add_6_33_groupi_g17101(csa_tree_add_6_33_groupi_n_1238 ,csa_tree_add_6_33_groupi_n_322 ,csa_tree_add_6_33_groupi_n_193);
  or csa_tree_add_6_33_groupi_g17102(csa_tree_add_6_33_groupi_n_1237 ,csa_tree_add_6_33_groupi_n_727 ,csa_tree_add_6_33_groupi_n_697);
  or csa_tree_add_6_33_groupi_g17103(csa_tree_add_6_33_groupi_n_1236 ,csa_tree_add_6_33_groupi_n_107 ,csa_tree_add_6_33_groupi_n_691);
  or csa_tree_add_6_33_groupi_g17104(csa_tree_add_6_33_groupi_n_1235 ,csa_tree_add_6_33_groupi_n_253 ,csa_tree_add_6_33_groupi_n_587);
  or csa_tree_add_6_33_groupi_g17105(csa_tree_add_6_33_groupi_n_1234 ,csa_tree_add_6_33_groupi_n_343 ,csa_tree_add_6_33_groupi_n_334);
  or csa_tree_add_6_33_groupi_g17106(csa_tree_add_6_33_groupi_n_1233 ,csa_tree_add_6_33_groupi_n_349 ,csa_tree_add_6_33_groupi_n_352);
  or csa_tree_add_6_33_groupi_g17107(csa_tree_add_6_33_groupi_n_1232 ,csa_tree_add_6_33_groupi_n_307 ,csa_tree_add_6_33_groupi_n_211);
  or csa_tree_add_6_33_groupi_g17108(csa_tree_add_6_33_groupi_n_1231 ,csa_tree_add_6_33_groupi_n_244 ,csa_tree_add_6_33_groupi_n_599);
  or csa_tree_add_6_33_groupi_g17109(csa_tree_add_6_33_groupi_n_1230 ,csa_tree_add_6_33_groupi_n_643 ,csa_tree_add_6_33_groupi_n_613);
  or csa_tree_add_6_33_groupi_g17110(csa_tree_add_6_33_groupi_n_1229 ,csa_tree_add_6_33_groupi_n_457 ,csa_tree_add_6_33_groupi_n_316);
  or csa_tree_add_6_33_groupi_g17111(csa_tree_add_6_33_groupi_n_1228 ,csa_tree_add_6_33_groupi_n_337 ,csa_tree_add_6_33_groupi_n_802);
  or csa_tree_add_6_33_groupi_g17112(csa_tree_add_6_33_groupi_n_1227 ,csa_tree_add_6_33_groupi_n_487 ,csa_tree_add_6_33_groupi_n_745);
  or csa_tree_add_6_33_groupi_g17113(csa_tree_add_6_33_groupi_n_1226 ,csa_tree_add_6_33_groupi_n_325 ,csa_tree_add_6_33_groupi_n_229);
  or csa_tree_add_6_33_groupi_g17114(csa_tree_add_6_33_groupi_n_1225 ,csa_tree_add_6_33_groupi_n_319 ,csa_tree_add_6_33_groupi_n_557);
  or csa_tree_add_6_33_groupi_g17115(csa_tree_add_6_33_groupi_n_1224 ,csa_tree_add_6_33_groupi_n_784 ,csa_tree_add_6_33_groupi_n_647);
  or csa_tree_add_6_33_groupi_g17116(csa_tree_add_6_33_groupi_n_1223 ,csa_tree_add_6_33_groupi_n_116 ,csa_tree_add_6_33_groupi_n_110);
  or csa_tree_add_6_33_groupi_g17117(csa_tree_add_6_33_groupi_n_1222 ,csa_tree_add_6_33_groupi_n_203 ,csa_tree_add_6_33_groupi_n_664);
  or csa_tree_add_6_33_groupi_g17118(csa_tree_add_6_33_groupi_n_1221 ,csa_tree_add_6_33_groupi_n_787 ,csa_tree_add_6_33_groupi_n_121);
  or csa_tree_add_6_33_groupi_g17119(csa_tree_add_6_33_groupi_n_1220 ,csa_tree_add_6_33_groupi_n_790 ,csa_tree_add_6_33_groupi_n_463);
  or csa_tree_add_6_33_groupi_g17120(csa_tree_add_6_33_groupi_n_1219 ,csa_tree_add_6_33_groupi_n_155 ,csa_tree_add_6_33_groupi_n_148);
  or csa_tree_add_6_33_groupi_g17121(csa_tree_add_6_33_groupi_n_1218 ,csa_tree_add_6_33_groupi_n_239 ,csa_tree_add_6_33_groupi_n_74);
  or csa_tree_add_6_33_groupi_g17122(csa_tree_add_6_33_groupi_n_1217 ,csa_tree_add_6_33_groupi_n_772 ,csa_tree_add_6_33_groupi_n_113);
  or csa_tree_add_6_33_groupi_g17123(csa_tree_add_6_33_groupi_n_1216 ,csa_tree_add_6_33_groupi_n_50 ,csa_tree_add_6_33_groupi_n_88);
  or csa_tree_add_6_33_groupi_g17124(csa_tree_add_6_33_groupi_n_1215 ,csa_tree_add_6_33_groupi_n_151 ,csa_tree_add_6_33_groupi_n_205);
  or csa_tree_add_6_33_groupi_g17125(csa_tree_add_6_33_groupi_n_1214 ,csa_tree_add_6_33_groupi_n_223 ,csa_tree_add_6_33_groupi_n_733);
  or csa_tree_add_6_33_groupi_g17126(csa_tree_add_6_33_groupi_n_1213 ,csa_tree_add_6_33_groupi_n_545 ,csa_tree_add_6_33_groupi_n_581);
  or csa_tree_add_6_33_groupi_g17127(csa_tree_add_6_33_groupi_n_1212 ,csa_tree_add_6_33_groupi_n_295 ,csa_tree_add_6_33_groupi_n_466);
  or csa_tree_add_6_33_groupi_g17128(csa_tree_add_6_33_groupi_n_1211 ,csa_tree_add_6_33_groupi_n_442 ,csa_tree_add_6_33_groupi_n_569);
  and csa_tree_add_6_33_groupi_g17129(csa_tree_add_6_33_groupi_n_1209 ,in1[3] ,in1[0]);
  or csa_tree_add_6_33_groupi_g17130(csa_tree_add_6_33_groupi_n_1208 ,csa_tree_add_6_33_groupi_n_305 ,csa_tree_add_6_33_groupi_n_289);
  or csa_tree_add_6_33_groupi_g17131(csa_tree_add_6_33_groupi_n_1207 ,csa_tree_add_6_33_groupi_n_65 ,csa_tree_add_6_33_groupi_n_649);
  or csa_tree_add_6_33_groupi_g17132(csa_tree_add_6_33_groupi_n_1206 ,csa_tree_add_6_33_groupi_n_185 ,csa_tree_add_6_33_groupi_n_280);
  or csa_tree_add_6_33_groupi_g17133(csa_tree_add_6_33_groupi_n_1205 ,csa_tree_add_6_33_groupi_n_250 ,csa_tree_add_6_33_groupi_n_302);
  or csa_tree_add_6_33_groupi_g17134(csa_tree_add_6_33_groupi_n_1204 ,csa_tree_add_6_33_groupi_n_62 ,csa_tree_add_6_33_groupi_n_101);
  or csa_tree_add_6_33_groupi_g17135(csa_tree_add_6_33_groupi_n_1203 ,csa_tree_add_6_33_groupi_n_479 ,csa_tree_add_6_33_groupi_n_311);
  or csa_tree_add_6_33_groupi_g17136(csa_tree_add_6_33_groupi_n_1202 ,csa_tree_add_6_33_groupi_n_637 ,csa_tree_add_6_33_groupi_n_658);
  or csa_tree_add_6_33_groupi_g17137(csa_tree_add_6_33_groupi_n_1201 ,csa_tree_add_6_33_groupi_n_503 ,csa_tree_add_6_33_groupi_n_454);
  or csa_tree_add_6_33_groupi_g17138(csa_tree_add_6_33_groupi_n_1200 ,csa_tree_add_6_33_groupi_n_287 ,csa_tree_add_6_33_groupi_n_712);
  or csa_tree_add_6_33_groupi_g17139(csa_tree_add_6_33_groupi_n_1199 ,csa_tree_add_6_33_groupi_n_331 ,csa_tree_add_6_33_groupi_n_95);
  or csa_tree_add_6_33_groupi_g17140(csa_tree_add_6_33_groupi_n_1198 ,csa_tree_add_6_33_groupi_n_716 ,csa_tree_add_6_33_groupi_n_221);
  or csa_tree_add_6_33_groupi_g17141(csa_tree_add_6_33_groupi_n_1197 ,csa_tree_add_6_33_groupi_n_683 ,csa_tree_add_6_33_groupi_n_383);
  or csa_tree_add_6_33_groupi_g17142(csa_tree_add_6_33_groupi_n_1196 ,csa_tree_add_6_33_groupi_n_449 ,csa_tree_add_6_33_groupi_n_274);
  or csa_tree_add_6_33_groupi_g17143(csa_tree_add_6_33_groupi_n_1195 ,csa_tree_add_6_33_groupi_n_83 ,csa_tree_add_6_33_groupi_n_98);
  or csa_tree_add_6_33_groupi_g17144(csa_tree_add_6_33_groupi_n_1194 ,csa_tree_add_6_33_groupi_n_164 ,csa_tree_add_6_33_groupi_n_419);
  or csa_tree_add_6_33_groupi_g17145(csa_tree_add_6_33_groupi_n_1193 ,csa_tree_add_6_33_groupi_n_313 ,csa_tree_add_6_33_groupi_n_365);
  or csa_tree_add_6_33_groupi_g17146(csa_tree_add_6_33_groupi_n_1192 ,csa_tree_add_6_33_groupi_n_719 ,csa_tree_add_6_33_groupi_n_446);
  or csa_tree_add_6_33_groupi_g17147(csa_tree_add_6_33_groupi_n_1191 ,csa_tree_add_6_33_groupi_n_737 ,csa_tree_add_6_33_groupi_n_413);
  or csa_tree_add_6_33_groupi_g17148(csa_tree_add_6_33_groupi_n_1190 ,csa_tree_add_6_33_groupi_n_485 ,csa_tree_add_6_33_groupi_n_631);
  or csa_tree_add_6_33_groupi_g17149(csa_tree_add_6_33_groupi_n_1189 ,csa_tree_add_6_33_groupi_n_371 ,csa_tree_add_6_33_groupi_n_92);
  or csa_tree_add_6_33_groupi_g17150(csa_tree_add_6_33_groupi_n_1188 ,csa_tree_add_6_33_groupi_n_272 ,csa_tree_add_6_33_groupi_n_172);
  or csa_tree_add_6_33_groupi_g17151(csa_tree_add_6_33_groupi_n_1187 ,csa_tree_add_6_33_groupi_n_656 ,csa_tree_add_6_33_groupi_n_629);
  or csa_tree_add_6_33_groupi_g17152(csa_tree_add_6_33_groupi_n_1186 ,csa_tree_add_6_33_groupi_n_187 ,csa_tree_add_6_33_groupi_n_515);
  or csa_tree_add_6_33_groupi_g17153(csa_tree_add_6_33_groupi_n_1185 ,csa_tree_add_6_33_groupi_n_575 ,csa_tree_add_6_33_groupi_n_461);
  or csa_tree_add_6_33_groupi_g17154(csa_tree_add_6_33_groupi_n_1184 ,csa_tree_add_6_33_groupi_n_68 ,csa_tree_add_6_33_groupi_n_119);
  or csa_tree_add_6_33_groupi_g17155(csa_tree_add_6_33_groupi_n_1183 ,csa_tree_add_6_33_groupi_n_563 ,csa_tree_add_6_33_groupi_n_470);
  or csa_tree_add_6_33_groupi_g17156(csa_tree_add_6_33_groupi_n_1182 ,csa_tree_add_6_33_groupi_n_347 ,csa_tree_add_6_33_groupi_n_407);
  or csa_tree_add_6_33_groupi_g17157(csa_tree_add_6_33_groupi_n_1181 ,csa_tree_add_6_33_groupi_n_539 ,csa_tree_add_6_33_groupi_n_59);
  or csa_tree_add_6_33_groupi_g17158(csa_tree_add_6_33_groupi_n_1180 ,csa_tree_add_6_33_groupi_n_341 ,csa_tree_add_6_33_groupi_n_701);
  or csa_tree_add_6_33_groupi_g17159(csa_tree_add_6_33_groupi_n_1179 ,csa_tree_add_6_33_groupi_n_242 ,csa_tree_add_6_33_groupi_n_679);
  or csa_tree_add_6_33_groupi_g17160(csa_tree_add_6_33_groupi_n_1178 ,csa_tree_add_6_33_groupi_n_533 ,csa_tree_add_6_33_groupi_n_751);
  or csa_tree_add_6_33_groupi_g17161(csa_tree_add_6_33_groupi_n_1177 ,csa_tree_add_6_33_groupi_n_808 ,csa_tree_add_6_33_groupi_n_778);
  or csa_tree_add_6_33_groupi_g17162(csa_tree_add_6_33_groupi_n_1176 ,csa_tree_add_6_33_groupi_n_671 ,csa_tree_add_6_33_groupi_n_56);
  or csa_tree_add_6_33_groupi_g17163(csa_tree_add_6_33_groupi_n_1175 ,csa_tree_add_6_33_groupi_n_268 ,csa_tree_add_6_33_groupi_n_673);
  or csa_tree_add_6_33_groupi_g17164(csa_tree_add_6_33_groupi_n_1174 ,csa_tree_add_6_33_groupi_n_209 ,csa_tree_add_6_33_groupi_n_166);
  or csa_tree_add_6_33_groupi_g17165(csa_tree_add_6_33_groupi_n_1173 ,csa_tree_add_6_33_groupi_n_805 ,csa_tree_add_6_33_groupi_n_215);
  or csa_tree_add_6_33_groupi_g17166(csa_tree_add_6_33_groupi_n_1172 ,csa_tree_add_6_33_groupi_n_509 ,csa_tree_add_6_33_groupi_n_428);
  or csa_tree_add_6_33_groupi_g17167(csa_tree_add_6_33_groupi_n_1171 ,csa_tree_add_6_33_groupi_n_425 ,csa_tree_add_6_33_groupi_n_46);
  or csa_tree_add_6_33_groupi_g17168(csa_tree_add_6_33_groupi_n_1170 ,csa_tree_add_6_33_groupi_n_431 ,csa_tree_add_6_33_groupi_n_677);
  or csa_tree_add_6_33_groupi_g17169(csa_tree_add_6_33_groupi_n_1169 ,csa_tree_add_6_33_groupi_n_524 ,csa_tree_add_6_33_groupi_n_652);
  or csa_tree_add_6_33_groupi_g17170(csa_tree_add_6_33_groupi_n_1168 ,csa_tree_add_6_33_groupi_n_227 ,csa_tree_add_6_33_groupi_n_619);
  or csa_tree_add_6_33_groupi_g17171(csa_tree_add_6_33_groupi_n_1167 ,csa_tree_add_6_33_groupi_n_757 ,csa_tree_add_6_33_groupi_n_659);
  or csa_tree_add_6_33_groupi_g17172(csa_tree_add_6_33_groupi_n_1166 ,csa_tree_add_6_33_groupi_n_641 ,csa_tree_add_6_33_groupi_n_709);
  or csa_tree_add_6_33_groupi_g17173(csa_tree_add_6_33_groupi_n_1165 ,csa_tree_add_6_33_groupi_n_299 ,csa_tree_add_6_33_groupi_n_161);
  or csa_tree_add_6_33_groupi_g17174(csa_tree_add_6_33_groupi_n_1164 ,csa_tree_add_6_33_groupi_n_566 ,csa_tree_add_6_33_groupi_n_194);
  or csa_tree_add_6_33_groupi_g17175(csa_tree_add_6_33_groupi_n_1163 ,csa_tree_add_6_33_groupi_n_689 ,csa_tree_add_6_33_groupi_n_71);
  or csa_tree_add_6_33_groupi_g17176(csa_tree_add_6_33_groupi_n_1162 ,csa_tree_add_6_33_groupi_n_182 ,csa_tree_add_6_33_groupi_n_554);
  and csa_tree_add_6_33_groupi_g17177(csa_tree_add_6_33_groupi_n_1160 ,in1[5] ,in1[4]);
  or csa_tree_add_6_33_groupi_g17178(csa_tree_add_6_33_groupi_n_1159 ,csa_tree_add_6_33_groupi_n_359 ,csa_tree_add_6_33_groupi_n_143);
  or csa_tree_add_6_33_groupi_g17179(csa_tree_add_6_33_groupi_n_1158 ,csa_tree_add_6_33_groupi_n_248 ,csa_tree_add_6_33_groupi_n_77);
  or csa_tree_add_6_33_groupi_g17180(csa_tree_add_6_33_groupi_n_1157 ,csa_tree_add_6_33_groupi_n_329 ,csa_tree_add_6_33_groupi_n_80);
  or csa_tree_add_6_33_groupi_g17181(csa_tree_add_6_33_groupi_n_1156 ,csa_tree_add_6_33_groupi_n_284 ,csa_tree_add_6_33_groupi_n_335);
  or csa_tree_add_6_33_groupi_g17182(csa_tree_add_6_33_groupi_n_1155 ,csa_tree_add_6_33_groupi_n_635 ,csa_tree_add_6_33_groupi_n_104);
  or csa_tree_add_6_33_groupi_g17183(csa_tree_add_6_33_groupi_n_1154 ,csa_tree_add_6_33_groupi_n_755 ,csa_tree_add_6_33_groupi_n_764);
  or csa_tree_add_6_33_groupi_g17184(csa_tree_add_6_33_groupi_n_1153 ,csa_tree_add_6_33_groupi_n_437 ,csa_tree_add_6_33_groupi_n_293);
  or csa_tree_add_6_33_groupi_g17185(csa_tree_add_6_33_groupi_n_1152 ,csa_tree_add_6_33_groupi_n_530 ,csa_tree_add_6_33_groupi_n_191);
  or csa_tree_add_6_33_groupi_g17186(csa_tree_add_6_33_groupi_n_1151 ,csa_tree_add_6_33_groupi_n_197 ,csa_tree_add_6_33_groupi_n_626);
  or csa_tree_add_6_33_groupi_g17187(csa_tree_add_6_33_groupi_n_1150 ,csa_tree_add_6_33_groupi_n_725 ,csa_tree_add_6_33_groupi_n_317);
  or csa_tree_add_6_33_groupi_g17188(csa_tree_add_6_33_groupi_n_1149 ,csa_tree_add_6_33_groupi_n_551 ,csa_tree_add_6_33_groupi_n_761);
  or csa_tree_add_6_33_groupi_g17189(csa_tree_add_6_33_groupi_n_1148 ,csa_tree_add_6_33_groupi_n_281 ,csa_tree_add_6_33_groupi_n_739);
  or csa_tree_add_6_33_groupi_g17190(csa_tree_add_6_33_groupi_n_1147 ,csa_tree_add_6_33_groupi_n_152 ,csa_tree_add_6_33_groupi_n_362);
  or csa_tree_add_6_33_groupi_g17191(csa_tree_add_6_33_groupi_n_1146 ,csa_tree_add_6_33_groupi_n_179 ,csa_tree_add_6_33_groupi_n_623);
  or csa_tree_add_6_33_groupi_g17192(csa_tree_add_6_33_groupi_n_1145 ,csa_tree_add_6_33_groupi_n_218 ,csa_tree_add_6_33_groupi_n_497);
  or csa_tree_add_6_33_groupi_g17193(csa_tree_add_6_33_groupi_n_1144 ,csa_tree_add_6_33_groupi_n_278 ,csa_tree_add_6_33_groupi_n_146);
  and csa_tree_add_6_33_groupi_g17194(csa_tree_add_6_33_groupi_n_1142 ,in1[10] ,in1[0]);
  or csa_tree_add_6_33_groupi_g17195(csa_tree_add_6_33_groupi_n_1141 ,csa_tree_add_6_33_groupi_n_251 ,csa_tree_add_6_33_groupi_n_454);
  or csa_tree_add_6_33_groupi_g17196(csa_tree_add_6_33_groupi_n_1140 ,csa_tree_add_6_33_groupi_n_542 ,csa_tree_add_6_33_groupi_n_257);
  or csa_tree_add_6_33_groupi_g17197(csa_tree_add_6_33_groupi_n_1139 ,csa_tree_add_6_33_groupi_n_506 ,csa_tree_add_6_33_groupi_n_332);
  and csa_tree_add_6_33_groupi_g17198(csa_tree_add_6_33_groupi_n_1137 ,in1[1] ,in1[0]);
  or csa_tree_add_6_33_groupi_g17199(csa_tree_add_6_33_groupi_n_1136 ,csa_tree_add_6_33_groupi_n_617 ,csa_tree_add_6_33_groupi_n_476);
  or csa_tree_add_6_33_groupi_g17200(csa_tree_add_6_33_groupi_n_1135 ,csa_tree_add_6_33_groupi_n_389 ,csa_tree_add_6_33_groupi_n_727);
  and csa_tree_add_6_33_groupi_g17201(csa_tree_add_6_33_groupi_n_1133 ,in1[13] ,in1[6]);
  or csa_tree_add_6_33_groupi_g17202(csa_tree_add_6_33_groupi_n_1132 ,csa_tree_add_6_33_groupi_n_440 ,csa_tree_add_6_33_groupi_n_697);
  or csa_tree_add_6_33_groupi_g17203(csa_tree_add_6_33_groupi_n_1131 ,csa_tree_add_6_33_groupi_n_260 ,csa_tree_add_6_33_groupi_n_731);
  or csa_tree_add_6_33_groupi_g17204(csa_tree_add_6_33_groupi_n_1130 ,csa_tree_add_6_33_groupi_n_536 ,csa_tree_add_6_33_groupi_n_628);
  or csa_tree_add_6_33_groupi_g17205(csa_tree_add_6_33_groupi_n_1129 ,csa_tree_add_6_33_groupi_n_473 ,csa_tree_add_6_33_groupi_n_691);
  or csa_tree_add_6_33_groupi_g17206(csa_tree_add_6_33_groupi_n_1128 ,csa_tree_add_6_33_groupi_n_398 ,csa_tree_add_6_33_groupi_n_392);
  or csa_tree_add_6_33_groupi_g17207(csa_tree_add_6_33_groupi_n_1127 ,csa_tree_add_6_33_groupi_n_296 ,csa_tree_add_6_33_groupi_n_376);
  or csa_tree_add_6_33_groupi_g17208(csa_tree_add_6_33_groupi_n_1126 ,csa_tree_add_6_33_groupi_n_491 ,csa_tree_add_6_33_groupi_n_721);
  or csa_tree_add_6_33_groupi_g17209(csa_tree_add_6_33_groupi_n_1125 ,csa_tree_add_6_33_groupi_n_526 ,csa_tree_add_6_33_groupi_n_767);
  or csa_tree_add_6_33_groupi_g17210(csa_tree_add_6_33_groupi_n_1124 ,csa_tree_add_6_33_groupi_n_500 ,csa_tree_add_6_33_groupi_n_400);
  or csa_tree_add_6_33_groupi_g17211(csa_tree_add_6_33_groupi_n_1123 ,csa_tree_add_6_33_groupi_n_158 ,csa_tree_add_6_33_groupi_n_467);
  or csa_tree_add_6_33_groupi_g17212(csa_tree_add_6_33_groupi_n_1122 ,csa_tree_add_6_33_groupi_n_314 ,csa_tree_add_6_33_groupi_n_703);
  or csa_tree_add_6_33_groupi_g17213(csa_tree_add_6_33_groupi_n_1121 ,csa_tree_add_6_33_groupi_n_443 ,csa_tree_add_6_33_groupi_n_380);
  or csa_tree_add_6_33_groupi_g17214(csa_tree_add_6_33_groupi_n_1120 ,csa_tree_add_6_33_groupi_n_323 ,csa_tree_add_6_33_groupi_n_745);
  or csa_tree_add_6_33_groupi_g17215(csa_tree_add_6_33_groupi_n_1119 ,csa_tree_add_6_33_groupi_n_245 ,csa_tree_add_6_33_groupi_n_269);
  or csa_tree_add_6_33_groupi_g17216(csa_tree_add_6_33_groupi_n_1118 ,csa_tree_add_6_33_groupi_n_452 ,csa_tree_add_6_33_groupi_n_148);
  or csa_tree_add_6_33_groupi_g17217(csa_tree_add_6_33_groupi_n_1117 ,csa_tree_add_6_33_groupi_n_265 ,csa_tree_add_6_33_groupi_n_650);
  or csa_tree_add_6_33_groupi_g17218(csa_tree_add_6_33_groupi_n_1116 ,csa_tree_add_6_33_groupi_n_140 ,csa_tree_add_6_33_groupi_n_653);
  or csa_tree_add_6_33_groupi_g17219(csa_tree_add_6_33_groupi_n_1115 ,csa_tree_add_6_33_groupi_n_44 ,csa_tree_add_6_33_groupi_n_608);
  or csa_tree_add_6_33_groupi_g17220(csa_tree_add_6_33_groupi_n_1114 ,csa_tree_add_6_33_groupi_n_416 ,csa_tree_add_6_33_groupi_n_620);
  or csa_tree_add_6_33_groupi_g17221(csa_tree_add_6_33_groupi_n_1113 ,csa_tree_add_6_33_groupi_n_368 ,csa_tree_add_6_33_groupi_n_169);
  or csa_tree_add_6_33_groupi_g17222(csa_tree_add_6_33_groupi_n_1112 ,csa_tree_add_6_33_groupi_n_668 ,csa_tree_add_6_33_groupi_n_685);
  or csa_tree_add_6_33_groupi_g17223(csa_tree_add_6_33_groupi_n_1111 ,csa_tree_add_6_33_groupi_n_200 ,csa_tree_add_6_33_groupi_n_596);
  or csa_tree_add_6_33_groupi_g17224(csa_tree_add_6_33_groupi_n_1110 ,csa_tree_add_6_33_groupi_n_233 ,csa_tree_add_6_33_groupi_n_89);
  or csa_tree_add_6_33_groupi_g17225(csa_tree_add_6_33_groupi_n_1109 ,csa_tree_add_6_33_groupi_n_602 ,csa_tree_add_6_33_groupi_n_356);
  or csa_tree_add_6_33_groupi_g17226(csa_tree_add_6_33_groupi_n_1108 ,csa_tree_add_6_33_groupi_n_661 ,csa_tree_add_6_33_groupi_n_352);
  and csa_tree_add_6_33_groupi_g17227(csa_tree_add_6_33_groupi_n_1106 ,in1[6] ,in1[0]);
  or csa_tree_add_6_33_groupi_g17228(csa_tree_add_6_33_groupi_n_1105 ,csa_tree_add_6_33_groupi_n_482 ,csa_tree_add_6_33_groupi_n_679);
  or csa_tree_add_6_33_groupi_g17229(csa_tree_add_6_33_groupi_n_1104 ,csa_tree_add_6_33_groupi_n_733 ,csa_tree_add_6_33_groupi_n_212);
  or csa_tree_add_6_33_groupi_g17230(csa_tree_add_6_33_groupi_n_1103 ,csa_tree_add_6_33_groupi_n_707 ,csa_tree_add_6_33_groupi_n_235);
  or csa_tree_add_6_33_groupi_g17231(csa_tree_add_6_33_groupi_n_1102 ,csa_tree_add_6_33_groupi_n_28 ,csa_tree_add_6_33_groupi_n_518);
  or csa_tree_add_6_33_groupi_g17232(csa_tree_add_6_33_groupi_n_1101 ,csa_tree_add_6_33_groupi_n_458 ,csa_tree_add_6_33_groupi_n_695);
  or csa_tree_add_6_33_groupi_g17233(csa_tree_add_6_33_groupi_n_1100 ,csa_tree_add_6_33_groupi_n_44 ,csa_tree_add_6_33_groupi_n_749);
  or csa_tree_add_6_33_groupi_g17234(csa_tree_add_6_33_groupi_n_1099 ,csa_tree_add_6_33_groupi_n_262 ,csa_tree_add_6_33_groupi_n_512);
  or csa_tree_add_6_33_groupi_g17235(csa_tree_add_6_33_groupi_n_1098 ,csa_tree_add_6_33_groupi_n_176 ,csa_tree_add_6_33_groupi_n_644);
  or csa_tree_add_6_33_groupi_g17236(csa_tree_add_6_33_groupi_n_1097 ,csa_tree_add_6_33_groupi_n_422 ,csa_tree_add_6_33_groupi_n_47);
  or csa_tree_add_6_33_groupi_g17237(csa_tree_add_6_33_groupi_n_1096 ,csa_tree_add_6_33_groupi_n_254 ,csa_tree_add_6_33_groupi_n_743);
  or csa_tree_add_6_33_groupi_g17238(csa_tree_add_6_33_groupi_n_1095 ,csa_tree_add_6_33_groupi_n_344 ,csa_tree_add_6_33_groupi_n_572);
  or csa_tree_add_6_33_groupi_g17239(csa_tree_add_6_33_groupi_n_1094 ,csa_tree_add_6_33_groupi_n_26 ,csa_tree_add_6_33_groupi_n_709);
  or csa_tree_add_6_33_groupi_g17240(csa_tree_add_6_33_groupi_n_1093 ,csa_tree_add_6_33_groupi_n_548 ,csa_tree_add_6_33_groupi_n_680);
  or csa_tree_add_6_33_groupi_g17241(csa_tree_add_6_33_groupi_n_1092 ,csa_tree_add_6_33_groupi_n_40 ,csa_tree_add_6_33_groupi_n_374);
  and csa_tree_add_6_33_groupi_g17242(csa_tree_add_6_33_groupi_n_1091 ,in1[13] ,in1[12]);
  or csa_tree_add_6_33_groupi_g17243(csa_tree_add_6_33_groupi_n_1090 ,csa_tree_add_6_33_groupi_n_590 ,csa_tree_add_6_33_groupi_n_494);
  or csa_tree_add_6_33_groupi_g17244(csa_tree_add_6_33_groupi_n_1089 ,csa_tree_add_6_33_groupi_n_718 ,csa_tree_add_6_33_groupi_n_584);
  or csa_tree_add_6_33_groupi_g17245(csa_tree_add_6_33_groupi_n_1088 ,csa_tree_add_6_33_groupi_n_638 ,csa_tree_add_6_33_groupi_n_20);
  or csa_tree_add_6_33_groupi_g17246(csa_tree_add_6_33_groupi_n_1087 ,csa_tree_add_6_33_groupi_n_713 ,csa_tree_add_6_33_groupi_n_308);
  or csa_tree_add_6_33_groupi_g17247(csa_tree_add_6_33_groupi_n_1086 ,csa_tree_add_6_33_groupi_n_614 ,csa_tree_add_6_33_groupi_n_665);
  or csa_tree_add_6_33_groupi_g17248(csa_tree_add_6_33_groupi_n_1085 ,csa_tree_add_6_33_groupi_n_404 ,csa_tree_add_6_33_groupi_n_350);
  or csa_tree_add_6_33_groupi_g17249(csa_tree_add_6_33_groupi_n_1084 ,csa_tree_add_6_33_groupi_n_338 ,csa_tree_add_6_33_groupi_n_632);
  or csa_tree_add_6_33_groupi_g17250(csa_tree_add_6_33_groupi_n_1083 ,csa_tree_add_6_33_groupi_n_36 ,csa_tree_add_6_33_groupi_n_568);
  or csa_tree_add_6_33_groupi_g17251(csa_tree_add_6_33_groupi_n_1082 ,csa_tree_add_6_33_groupi_n_24 ,csa_tree_add_6_33_groupi_n_178);
  or csa_tree_add_6_33_groupi_g17252(csa_tree_add_6_33_groupi_n_1081 ,csa_tree_add_6_33_groupi_n_38 ,csa_tree_add_6_33_groupi_n_301);
  or csa_tree_add_6_33_groupi_g17253(csa_tree_add_6_33_groupi_n_1080 ,csa_tree_add_6_33_groupi_n_58 ,csa_tree_add_6_33_groupi_n_739);
  or csa_tree_add_6_33_groupi_g17254(csa_tree_add_6_33_groupi_n_1079 ,csa_tree_add_6_33_groupi_n_22 ,csa_tree_add_6_33_groupi_n_386);
  or csa_tree_add_6_33_groupi_g17255(csa_tree_add_6_33_groupi_n_1078 ,csa_tree_add_6_33_groupi_n_434 ,csa_tree_add_6_33_groupi_n_488);
  or csa_tree_add_6_33_groupi_g17256(csa_tree_add_6_33_groupi_n_1077 ,csa_tree_add_6_33_groupi_n_30 ,csa_tree_add_6_33_groupi_n_214);
  or csa_tree_add_6_33_groupi_g17257(csa_tree_add_6_33_groupi_n_1076 ,csa_tree_add_6_33_groupi_n_224 ,csa_tree_add_6_33_groupi_n_34);
  or csa_tree_add_6_33_groupi_g17258(csa_tree_add_6_33_groupi_n_1075 ,csa_tree_add_6_33_groupi_n_578 ,csa_tree_add_6_33_groupi_n_115);
  or csa_tree_add_6_33_groupi_g17259(csa_tree_add_6_33_groupi_n_1074 ,csa_tree_add_6_33_groupi_n_42 ,csa_tree_add_6_33_groupi_n_188);
  or csa_tree_add_6_33_groupi_g17260(csa_tree_add_6_33_groupi_n_1073 ,csa_tree_add_6_33_groupi_n_560 ,csa_tree_add_6_33_groupi_n_625);
  or csa_tree_add_6_33_groupi_g17261(csa_tree_add_6_33_groupi_n_1072 ,csa_tree_add_6_33_groupi_n_326 ,csa_tree_add_6_33_groupi_n_18);
  or csa_tree_add_6_33_groupi_g17262(csa_tree_add_6_33_groupi_n_1071 ,csa_tree_add_6_33_groupi_n_320 ,csa_tree_add_6_33_groupi_n_652);
  or csa_tree_add_6_33_groupi_g17263(csa_tree_add_6_33_groupi_n_1070 ,csa_tree_add_6_33_groupi_n_32 ,csa_tree_add_6_33_groupi_n_410);
  not csa_tree_add_6_33_groupi_g17264(csa_tree_add_6_33_groupi_n_1041 ,in3[16]);
  not csa_tree_add_6_33_groupi_g17265(csa_tree_add_6_33_groupi_n_1040 ,in1[0]);
  not csa_tree_add_6_33_groupi_g17266(csa_tree_add_6_33_groupi_n_1039 ,in1[3]);
  not csa_tree_add_6_33_groupi_g17267(csa_tree_add_6_33_groupi_n_1038 ,in1[2]);
  not csa_tree_add_6_33_groupi_g17268(csa_tree_add_6_33_groupi_n_1037 ,in1[9]);
  not csa_tree_add_6_33_groupi_g17269(csa_tree_add_6_33_groupi_n_1036 ,in1[6]);
  not csa_tree_add_6_33_groupi_g17270(csa_tree_add_6_33_groupi_n_1035 ,in1[11]);
  not csa_tree_add_6_33_groupi_g17271(csa_tree_add_6_33_groupi_n_1034 ,in1[18]);
  not csa_tree_add_6_33_groupi_g17272(csa_tree_add_6_33_groupi_n_1033 ,in1[26]);
  not csa_tree_add_6_33_groupi_g17273(csa_tree_add_6_33_groupi_n_1032 ,in1[10]);
  not csa_tree_add_6_33_groupi_g17274(csa_tree_add_6_33_groupi_n_1031 ,in1[15]);
  not csa_tree_add_6_33_groupi_g17275(csa_tree_add_6_33_groupi_n_1030 ,in1[5]);
  not csa_tree_add_6_33_groupi_g17276(csa_tree_add_6_33_groupi_n_1029 ,in1[30]);
  not csa_tree_add_6_33_groupi_g17277(csa_tree_add_6_33_groupi_n_1028 ,in1[27]);
  not csa_tree_add_6_33_groupi_g17278(csa_tree_add_6_33_groupi_n_1027 ,in1[21]);
  not csa_tree_add_6_33_groupi_g17279(csa_tree_add_6_33_groupi_n_1026 ,in1[29]);
  not csa_tree_add_6_33_groupi_g17280(csa_tree_add_6_33_groupi_n_1025 ,in1[24]);
  not csa_tree_add_6_33_groupi_g17281(csa_tree_add_6_33_groupi_n_1024 ,in1[12]);
  not csa_tree_add_6_33_groupi_g17282(csa_tree_add_6_33_groupi_n_1023 ,in1[1]);
  not csa_tree_add_6_33_groupi_g17283(csa_tree_add_6_33_groupi_n_1022 ,in2[16]);
  not csa_tree_add_6_33_groupi_g17284(csa_tree_add_6_33_groupi_n_1021 ,in1[4]);
  not csa_tree_add_6_33_groupi_g17285(csa_tree_add_6_33_groupi_n_1020 ,in1[16]);
  not csa_tree_add_6_33_groupi_g17286(csa_tree_add_6_33_groupi_n_1019 ,in1[20]);
  not csa_tree_add_6_33_groupi_g17287(csa_tree_add_6_33_groupi_n_1018 ,in1[23]);
  not csa_tree_add_6_33_groupi_g17288(csa_tree_add_6_33_groupi_n_1017 ,in1[17]);
  not csa_tree_add_6_33_groupi_g17289(csa_tree_add_6_33_groupi_n_1016 ,in1[7]);
  not csa_tree_add_6_33_groupi_g17290(csa_tree_add_6_33_groupi_n_1015 ,in1[14]);
  not csa_tree_add_6_33_groupi_g17291(csa_tree_add_6_33_groupi_n_1014 ,in1[13]);
  not csa_tree_add_6_33_groupi_g17292(csa_tree_add_6_33_groupi_n_1013 ,in1[25]);
  not csa_tree_add_6_33_groupi_g17293(csa_tree_add_6_33_groupi_n_1012 ,in1[31]);
  not csa_tree_add_6_33_groupi_g17294(csa_tree_add_6_33_groupi_n_1011 ,in1[22]);
  not csa_tree_add_6_33_groupi_g17295(csa_tree_add_6_33_groupi_n_1010 ,in1[19]);
  not csa_tree_add_6_33_groupi_g17296(csa_tree_add_6_33_groupi_n_1009 ,in1[28]);
  not csa_tree_add_6_33_groupi_g17297(csa_tree_add_6_33_groupi_n_1008 ,in1[8]);
  not csa_tree_add_6_33_groupi_drc_bufs(csa_tree_add_6_33_groupi_n_1005 ,csa_tree_add_6_33_groupi_n_853);
  not csa_tree_add_6_33_groupi_drc_bufs17298(csa_tree_add_6_33_groupi_n_1004 ,csa_tree_add_6_33_groupi_n_854);
  not csa_tree_add_6_33_groupi_drc_bufs17299(csa_tree_add_6_33_groupi_n_1003 ,csa_tree_add_6_33_groupi_n_853);
  not csa_tree_add_6_33_groupi_drc_bufs17300(csa_tree_add_6_33_groupi_n_1002 ,csa_tree_add_6_33_groupi_n_854);
  not csa_tree_add_6_33_groupi_drc_bufs17305(csa_tree_add_6_33_groupi_n_1001 ,csa_tree_add_6_33_groupi_n_857);
  not csa_tree_add_6_33_groupi_drc_bufs17306(csa_tree_add_6_33_groupi_n_1000 ,csa_tree_add_6_33_groupi_n_858);
  not csa_tree_add_6_33_groupi_drc_bufs17307(csa_tree_add_6_33_groupi_n_999 ,csa_tree_add_6_33_groupi_n_857);
  not csa_tree_add_6_33_groupi_drc_bufs17308(csa_tree_add_6_33_groupi_n_998 ,csa_tree_add_6_33_groupi_n_858);
  not csa_tree_add_6_33_groupi_drc_bufs17313(csa_tree_add_6_33_groupi_n_997 ,csa_tree_add_6_33_groupi_n_871);
  not csa_tree_add_6_33_groupi_drc_bufs17314(csa_tree_add_6_33_groupi_n_996 ,csa_tree_add_6_33_groupi_n_872);
  not csa_tree_add_6_33_groupi_drc_bufs17315(csa_tree_add_6_33_groupi_n_995 ,csa_tree_add_6_33_groupi_n_871);
  not csa_tree_add_6_33_groupi_drc_bufs17316(csa_tree_add_6_33_groupi_n_994 ,csa_tree_add_6_33_groupi_n_872);
  not csa_tree_add_6_33_groupi_drc_bufs17321(csa_tree_add_6_33_groupi_n_993 ,csa_tree_add_6_33_groupi_n_825);
  not csa_tree_add_6_33_groupi_drc_bufs17322(csa_tree_add_6_33_groupi_n_992 ,csa_tree_add_6_33_groupi_n_826);
  not csa_tree_add_6_33_groupi_drc_bufs17323(csa_tree_add_6_33_groupi_n_991 ,csa_tree_add_6_33_groupi_n_825);
  not csa_tree_add_6_33_groupi_drc_bufs17324(csa_tree_add_6_33_groupi_n_990 ,csa_tree_add_6_33_groupi_n_826);
  not csa_tree_add_6_33_groupi_drc_bufs17329(csa_tree_add_6_33_groupi_n_989 ,csa_tree_add_6_33_groupi_n_847);
  not csa_tree_add_6_33_groupi_drc_bufs17330(csa_tree_add_6_33_groupi_n_988 ,csa_tree_add_6_33_groupi_n_848);
  not csa_tree_add_6_33_groupi_drc_bufs17331(csa_tree_add_6_33_groupi_n_987 ,csa_tree_add_6_33_groupi_n_847);
  not csa_tree_add_6_33_groupi_drc_bufs17332(csa_tree_add_6_33_groupi_n_986 ,csa_tree_add_6_33_groupi_n_848);
  not csa_tree_add_6_33_groupi_drc_bufs17337(csa_tree_add_6_33_groupi_n_985 ,csa_tree_add_6_33_groupi_n_833);
  not csa_tree_add_6_33_groupi_drc_bufs17338(csa_tree_add_6_33_groupi_n_984 ,csa_tree_add_6_33_groupi_n_834);
  not csa_tree_add_6_33_groupi_drc_bufs17339(csa_tree_add_6_33_groupi_n_983 ,csa_tree_add_6_33_groupi_n_833);
  not csa_tree_add_6_33_groupi_drc_bufs17340(csa_tree_add_6_33_groupi_n_982 ,csa_tree_add_6_33_groupi_n_834);
  not csa_tree_add_6_33_groupi_drc_bufs17345(csa_tree_add_6_33_groupi_n_981 ,csa_tree_add_6_33_groupi_n_835);
  not csa_tree_add_6_33_groupi_drc_bufs17346(csa_tree_add_6_33_groupi_n_980 ,csa_tree_add_6_33_groupi_n_836);
  not csa_tree_add_6_33_groupi_drc_bufs17347(csa_tree_add_6_33_groupi_n_979 ,csa_tree_add_6_33_groupi_n_835);
  not csa_tree_add_6_33_groupi_drc_bufs17348(csa_tree_add_6_33_groupi_n_978 ,csa_tree_add_6_33_groupi_n_836);
  not csa_tree_add_6_33_groupi_drc_bufs17353(csa_tree_add_6_33_groupi_n_977 ,csa_tree_add_6_33_groupi_n_861);
  not csa_tree_add_6_33_groupi_drc_bufs17354(csa_tree_add_6_33_groupi_n_976 ,csa_tree_add_6_33_groupi_n_862);
  not csa_tree_add_6_33_groupi_drc_bufs17355(csa_tree_add_6_33_groupi_n_975 ,csa_tree_add_6_33_groupi_n_861);
  not csa_tree_add_6_33_groupi_drc_bufs17356(csa_tree_add_6_33_groupi_n_974 ,csa_tree_add_6_33_groupi_n_862);
  not csa_tree_add_6_33_groupi_drc_bufs17361(csa_tree_add_6_33_groupi_n_973 ,csa_tree_add_6_33_groupi_n_829);
  not csa_tree_add_6_33_groupi_drc_bufs17362(csa_tree_add_6_33_groupi_n_972 ,csa_tree_add_6_33_groupi_n_830);
  not csa_tree_add_6_33_groupi_drc_bufs17363(csa_tree_add_6_33_groupi_n_971 ,csa_tree_add_6_33_groupi_n_829);
  not csa_tree_add_6_33_groupi_drc_bufs17364(csa_tree_add_6_33_groupi_n_970 ,csa_tree_add_6_33_groupi_n_830);
  not csa_tree_add_6_33_groupi_drc_bufs17369(csa_tree_add_6_33_groupi_n_969 ,csa_tree_add_6_33_groupi_n_831);
  not csa_tree_add_6_33_groupi_drc_bufs17370(csa_tree_add_6_33_groupi_n_968 ,csa_tree_add_6_33_groupi_n_832);
  not csa_tree_add_6_33_groupi_drc_bufs17371(csa_tree_add_6_33_groupi_n_967 ,csa_tree_add_6_33_groupi_n_831);
  not csa_tree_add_6_33_groupi_drc_bufs17372(csa_tree_add_6_33_groupi_n_966 ,csa_tree_add_6_33_groupi_n_832);
  not csa_tree_add_6_33_groupi_drc_bufs17377(csa_tree_add_6_33_groupi_n_965 ,csa_tree_add_6_33_groupi_n_819);
  not csa_tree_add_6_33_groupi_drc_bufs17378(csa_tree_add_6_33_groupi_n_964 ,csa_tree_add_6_33_groupi_n_820);
  not csa_tree_add_6_33_groupi_drc_bufs17379(csa_tree_add_6_33_groupi_n_963 ,csa_tree_add_6_33_groupi_n_819);
  not csa_tree_add_6_33_groupi_drc_bufs17380(csa_tree_add_6_33_groupi_n_962 ,csa_tree_add_6_33_groupi_n_820);
  not csa_tree_add_6_33_groupi_drc_bufs17385(csa_tree_add_6_33_groupi_n_961 ,csa_tree_add_6_33_groupi_n_863);
  not csa_tree_add_6_33_groupi_drc_bufs17386(csa_tree_add_6_33_groupi_n_960 ,csa_tree_add_6_33_groupi_n_864);
  not csa_tree_add_6_33_groupi_drc_bufs17387(csa_tree_add_6_33_groupi_n_959 ,csa_tree_add_6_33_groupi_n_863);
  not csa_tree_add_6_33_groupi_drc_bufs17388(csa_tree_add_6_33_groupi_n_958 ,csa_tree_add_6_33_groupi_n_864);
  not csa_tree_add_6_33_groupi_drc_bufs17393(csa_tree_add_6_33_groupi_n_957 ,csa_tree_add_6_33_groupi_n_873);
  not csa_tree_add_6_33_groupi_drc_bufs17394(csa_tree_add_6_33_groupi_n_956 ,csa_tree_add_6_33_groupi_n_874);
  not csa_tree_add_6_33_groupi_drc_bufs17395(csa_tree_add_6_33_groupi_n_955 ,csa_tree_add_6_33_groupi_n_873);
  not csa_tree_add_6_33_groupi_drc_bufs17396(csa_tree_add_6_33_groupi_n_954 ,csa_tree_add_6_33_groupi_n_874);
  not csa_tree_add_6_33_groupi_drc_bufs17401(csa_tree_add_6_33_groupi_n_953 ,csa_tree_add_6_33_groupi_n_875);
  not csa_tree_add_6_33_groupi_drc_bufs17402(csa_tree_add_6_33_groupi_n_952 ,csa_tree_add_6_33_groupi_n_876);
  not csa_tree_add_6_33_groupi_drc_bufs17403(csa_tree_add_6_33_groupi_n_951 ,csa_tree_add_6_33_groupi_n_875);
  not csa_tree_add_6_33_groupi_drc_bufs17404(csa_tree_add_6_33_groupi_n_950 ,csa_tree_add_6_33_groupi_n_876);
  not csa_tree_add_6_33_groupi_drc_bufs17409(csa_tree_add_6_33_groupi_n_949 ,csa_tree_add_6_33_groupi_n_845);
  not csa_tree_add_6_33_groupi_drc_bufs17410(csa_tree_add_6_33_groupi_n_948 ,csa_tree_add_6_33_groupi_n_846);
  not csa_tree_add_6_33_groupi_drc_bufs17411(csa_tree_add_6_33_groupi_n_947 ,csa_tree_add_6_33_groupi_n_845);
  not csa_tree_add_6_33_groupi_drc_bufs17412(csa_tree_add_6_33_groupi_n_946 ,csa_tree_add_6_33_groupi_n_846);
  not csa_tree_add_6_33_groupi_drc_bufs17417(csa_tree_add_6_33_groupi_n_945 ,csa_tree_add_6_33_groupi_n_843);
  not csa_tree_add_6_33_groupi_drc_bufs17418(csa_tree_add_6_33_groupi_n_944 ,csa_tree_add_6_33_groupi_n_844);
  not csa_tree_add_6_33_groupi_drc_bufs17419(csa_tree_add_6_33_groupi_n_943 ,csa_tree_add_6_33_groupi_n_843);
  not csa_tree_add_6_33_groupi_drc_bufs17420(csa_tree_add_6_33_groupi_n_942 ,csa_tree_add_6_33_groupi_n_844);
  not csa_tree_add_6_33_groupi_drc_bufs17425(csa_tree_add_6_33_groupi_n_941 ,csa_tree_add_6_33_groupi_n_859);
  not csa_tree_add_6_33_groupi_drc_bufs17426(csa_tree_add_6_33_groupi_n_940 ,csa_tree_add_6_33_groupi_n_860);
  not csa_tree_add_6_33_groupi_drc_bufs17427(csa_tree_add_6_33_groupi_n_939 ,csa_tree_add_6_33_groupi_n_859);
  not csa_tree_add_6_33_groupi_drc_bufs17428(csa_tree_add_6_33_groupi_n_938 ,csa_tree_add_6_33_groupi_n_860);
  not csa_tree_add_6_33_groupi_drc_bufs17433(csa_tree_add_6_33_groupi_n_937 ,csa_tree_add_6_33_groupi_n_869);
  not csa_tree_add_6_33_groupi_drc_bufs17434(csa_tree_add_6_33_groupi_n_936 ,csa_tree_add_6_33_groupi_n_870);
  not csa_tree_add_6_33_groupi_drc_bufs17435(csa_tree_add_6_33_groupi_n_935 ,csa_tree_add_6_33_groupi_n_869);
  not csa_tree_add_6_33_groupi_drc_bufs17436(csa_tree_add_6_33_groupi_n_934 ,csa_tree_add_6_33_groupi_n_870);
  not csa_tree_add_6_33_groupi_drc_bufs17441(csa_tree_add_6_33_groupi_n_933 ,csa_tree_add_6_33_groupi_n_817);
  not csa_tree_add_6_33_groupi_drc_bufs17442(csa_tree_add_6_33_groupi_n_932 ,csa_tree_add_6_33_groupi_n_818);
  not csa_tree_add_6_33_groupi_drc_bufs17443(csa_tree_add_6_33_groupi_n_931 ,csa_tree_add_6_33_groupi_n_817);
  not csa_tree_add_6_33_groupi_drc_bufs17444(csa_tree_add_6_33_groupi_n_930 ,csa_tree_add_6_33_groupi_n_818);
  not csa_tree_add_6_33_groupi_drc_bufs17449(csa_tree_add_6_33_groupi_n_929 ,csa_tree_add_6_33_groupi_n_851);
  not csa_tree_add_6_33_groupi_drc_bufs17450(csa_tree_add_6_33_groupi_n_928 ,csa_tree_add_6_33_groupi_n_852);
  not csa_tree_add_6_33_groupi_drc_bufs17451(csa_tree_add_6_33_groupi_n_927 ,csa_tree_add_6_33_groupi_n_851);
  not csa_tree_add_6_33_groupi_drc_bufs17452(csa_tree_add_6_33_groupi_n_926 ,csa_tree_add_6_33_groupi_n_852);
  not csa_tree_add_6_33_groupi_drc_bufs17457(csa_tree_add_6_33_groupi_n_925 ,csa_tree_add_6_33_groupi_n_827);
  not csa_tree_add_6_33_groupi_drc_bufs17458(csa_tree_add_6_33_groupi_n_924 ,csa_tree_add_6_33_groupi_n_828);
  not csa_tree_add_6_33_groupi_drc_bufs17459(csa_tree_add_6_33_groupi_n_923 ,csa_tree_add_6_33_groupi_n_827);
  not csa_tree_add_6_33_groupi_drc_bufs17460(csa_tree_add_6_33_groupi_n_922 ,csa_tree_add_6_33_groupi_n_828);
  not csa_tree_add_6_33_groupi_drc_bufs17465(csa_tree_add_6_33_groupi_n_921 ,csa_tree_add_6_33_groupi_n_855);
  not csa_tree_add_6_33_groupi_drc_bufs17466(csa_tree_add_6_33_groupi_n_920 ,csa_tree_add_6_33_groupi_n_856);
  not csa_tree_add_6_33_groupi_drc_bufs17467(csa_tree_add_6_33_groupi_n_919 ,csa_tree_add_6_33_groupi_n_855);
  not csa_tree_add_6_33_groupi_drc_bufs17468(csa_tree_add_6_33_groupi_n_918 ,csa_tree_add_6_33_groupi_n_856);
  not csa_tree_add_6_33_groupi_drc_bufs17473(csa_tree_add_6_33_groupi_n_917 ,csa_tree_add_6_33_groupi_n_823);
  not csa_tree_add_6_33_groupi_drc_bufs17474(csa_tree_add_6_33_groupi_n_916 ,csa_tree_add_6_33_groupi_n_824);
  not csa_tree_add_6_33_groupi_drc_bufs17475(csa_tree_add_6_33_groupi_n_915 ,csa_tree_add_6_33_groupi_n_823);
  not csa_tree_add_6_33_groupi_drc_bufs17476(csa_tree_add_6_33_groupi_n_914 ,csa_tree_add_6_33_groupi_n_824);
  not csa_tree_add_6_33_groupi_drc_bufs17481(csa_tree_add_6_33_groupi_n_913 ,csa_tree_add_6_33_groupi_n_821);
  not csa_tree_add_6_33_groupi_drc_bufs17482(csa_tree_add_6_33_groupi_n_912 ,csa_tree_add_6_33_groupi_n_822);
  not csa_tree_add_6_33_groupi_drc_bufs17483(csa_tree_add_6_33_groupi_n_911 ,csa_tree_add_6_33_groupi_n_821);
  not csa_tree_add_6_33_groupi_drc_bufs17484(csa_tree_add_6_33_groupi_n_910 ,csa_tree_add_6_33_groupi_n_822);
  not csa_tree_add_6_33_groupi_drc_bufs17489(csa_tree_add_6_33_groupi_n_909 ,csa_tree_add_6_33_groupi_n_815);
  not csa_tree_add_6_33_groupi_drc_bufs17490(csa_tree_add_6_33_groupi_n_908 ,csa_tree_add_6_33_groupi_n_816);
  not csa_tree_add_6_33_groupi_drc_bufs17491(csa_tree_add_6_33_groupi_n_907 ,csa_tree_add_6_33_groupi_n_815);
  not csa_tree_add_6_33_groupi_drc_bufs17492(csa_tree_add_6_33_groupi_n_906 ,csa_tree_add_6_33_groupi_n_816);
  not csa_tree_add_6_33_groupi_drc_bufs17497(csa_tree_add_6_33_groupi_n_905 ,csa_tree_add_6_33_groupi_n_865);
  not csa_tree_add_6_33_groupi_drc_bufs17498(csa_tree_add_6_33_groupi_n_904 ,csa_tree_add_6_33_groupi_n_866);
  not csa_tree_add_6_33_groupi_drc_bufs17499(csa_tree_add_6_33_groupi_n_903 ,csa_tree_add_6_33_groupi_n_865);
  not csa_tree_add_6_33_groupi_drc_bufs17500(csa_tree_add_6_33_groupi_n_902 ,csa_tree_add_6_33_groupi_n_866);
  not csa_tree_add_6_33_groupi_drc_bufs17505(csa_tree_add_6_33_groupi_n_901 ,csa_tree_add_6_33_groupi_n_867);
  not csa_tree_add_6_33_groupi_drc_bufs17506(csa_tree_add_6_33_groupi_n_900 ,csa_tree_add_6_33_groupi_n_868);
  not csa_tree_add_6_33_groupi_drc_bufs17507(csa_tree_add_6_33_groupi_n_899 ,csa_tree_add_6_33_groupi_n_867);
  not csa_tree_add_6_33_groupi_drc_bufs17508(csa_tree_add_6_33_groupi_n_898 ,csa_tree_add_6_33_groupi_n_868);
  not csa_tree_add_6_33_groupi_drc_bufs17513(csa_tree_add_6_33_groupi_n_897 ,csa_tree_add_6_33_groupi_n_849);
  not csa_tree_add_6_33_groupi_drc_bufs17514(csa_tree_add_6_33_groupi_n_896 ,csa_tree_add_6_33_groupi_n_850);
  not csa_tree_add_6_33_groupi_drc_bufs17515(csa_tree_add_6_33_groupi_n_895 ,csa_tree_add_6_33_groupi_n_849);
  not csa_tree_add_6_33_groupi_drc_bufs17516(csa_tree_add_6_33_groupi_n_894 ,csa_tree_add_6_33_groupi_n_850);
  not csa_tree_add_6_33_groupi_drc_bufs17521(csa_tree_add_6_33_groupi_n_893 ,csa_tree_add_6_33_groupi_n_837);
  not csa_tree_add_6_33_groupi_drc_bufs17522(csa_tree_add_6_33_groupi_n_892 ,csa_tree_add_6_33_groupi_n_838);
  not csa_tree_add_6_33_groupi_drc_bufs17523(csa_tree_add_6_33_groupi_n_891 ,csa_tree_add_6_33_groupi_n_837);
  not csa_tree_add_6_33_groupi_drc_bufs17524(csa_tree_add_6_33_groupi_n_890 ,csa_tree_add_6_33_groupi_n_838);
  not csa_tree_add_6_33_groupi_drc_bufs17529(csa_tree_add_6_33_groupi_n_889 ,csa_tree_add_6_33_groupi_n_839);
  not csa_tree_add_6_33_groupi_drc_bufs17530(csa_tree_add_6_33_groupi_n_888 ,csa_tree_add_6_33_groupi_n_840);
  not csa_tree_add_6_33_groupi_drc_bufs17531(csa_tree_add_6_33_groupi_n_887 ,csa_tree_add_6_33_groupi_n_839);
  not csa_tree_add_6_33_groupi_drc_bufs17532(csa_tree_add_6_33_groupi_n_886 ,csa_tree_add_6_33_groupi_n_840);
  not csa_tree_add_6_33_groupi_drc_bufs17537(csa_tree_add_6_33_groupi_n_885 ,csa_tree_add_6_33_groupi_n_813);
  not csa_tree_add_6_33_groupi_drc_bufs17538(csa_tree_add_6_33_groupi_n_884 ,csa_tree_add_6_33_groupi_n_814);
  not csa_tree_add_6_33_groupi_drc_bufs17539(csa_tree_add_6_33_groupi_n_883 ,csa_tree_add_6_33_groupi_n_813);
  not csa_tree_add_6_33_groupi_drc_bufs17540(csa_tree_add_6_33_groupi_n_882 ,csa_tree_add_6_33_groupi_n_814);
  not csa_tree_add_6_33_groupi_drc_bufs17545(csa_tree_add_6_33_groupi_n_881 ,csa_tree_add_6_33_groupi_n_841);
  not csa_tree_add_6_33_groupi_drc_bufs17546(csa_tree_add_6_33_groupi_n_880 ,csa_tree_add_6_33_groupi_n_842);
  not csa_tree_add_6_33_groupi_drc_bufs17547(csa_tree_add_6_33_groupi_n_879 ,csa_tree_add_6_33_groupi_n_841);
  not csa_tree_add_6_33_groupi_drc_bufs17548(csa_tree_add_6_33_groupi_n_878 ,csa_tree_add_6_33_groupi_n_842);
  not csa_tree_add_6_33_groupi_drc_bufs17563(csa_tree_add_6_33_groupi_n_877 ,csa_tree_add_6_33_groupi_n_1006);
  not csa_tree_add_6_33_groupi_drc_bufs17564(csa_tree_add_6_33_groupi_n_1006 ,csa_tree_add_6_33_groupi_n_2669);
  not csa_tree_add_6_33_groupi_drc_bufs17568(csa_tree_add_6_33_groupi_n_1007 ,csa_tree_add_6_33_groupi_n_3979);
  not csa_tree_add_6_33_groupi_drc_bufs18182(csa_tree_add_6_33_groupi_n_876 ,csa_tree_add_6_33_groupi_n_1009);
  not csa_tree_add_6_33_groupi_drc_bufs18183(csa_tree_add_6_33_groupi_n_875 ,csa_tree_add_6_33_groupi_n_1009);
  not csa_tree_add_6_33_groupi_drc_bufs18186(csa_tree_add_6_33_groupi_n_874 ,csa_tree_add_6_33_groupi_n_1010);
  not csa_tree_add_6_33_groupi_drc_bufs18187(csa_tree_add_6_33_groupi_n_873 ,csa_tree_add_6_33_groupi_n_1010);
  not csa_tree_add_6_33_groupi_drc_bufs18190(csa_tree_add_6_33_groupi_n_872 ,csa_tree_add_6_33_groupi_n_1026);
  not csa_tree_add_6_33_groupi_drc_bufs18191(csa_tree_add_6_33_groupi_n_871 ,csa_tree_add_6_33_groupi_n_1026);
  not csa_tree_add_6_33_groupi_drc_bufs18194(csa_tree_add_6_33_groupi_n_870 ,csa_tree_add_6_33_groupi_n_1031);
  not csa_tree_add_6_33_groupi_drc_bufs18195(csa_tree_add_6_33_groupi_n_869 ,csa_tree_add_6_33_groupi_n_1031);
  not csa_tree_add_6_33_groupi_drc_bufs18198(csa_tree_add_6_33_groupi_n_868 ,csa_tree_add_6_33_groupi_n_1024);
  not csa_tree_add_6_33_groupi_drc_bufs18199(csa_tree_add_6_33_groupi_n_867 ,csa_tree_add_6_33_groupi_n_1024);
  not csa_tree_add_6_33_groupi_drc_bufs18202(csa_tree_add_6_33_groupi_n_866 ,csa_tree_add_6_33_groupi_n_1030);
  not csa_tree_add_6_33_groupi_drc_bufs18203(csa_tree_add_6_33_groupi_n_865 ,csa_tree_add_6_33_groupi_n_1030);
  not csa_tree_add_6_33_groupi_drc_bufs18206(csa_tree_add_6_33_groupi_n_864 ,csa_tree_add_6_33_groupi_n_1011);
  not csa_tree_add_6_33_groupi_drc_bufs18207(csa_tree_add_6_33_groupi_n_863 ,csa_tree_add_6_33_groupi_n_1011);
  not csa_tree_add_6_33_groupi_drc_bufs18210(csa_tree_add_6_33_groupi_n_862 ,csa_tree_add_6_33_groupi_n_1017);
  not csa_tree_add_6_33_groupi_drc_bufs18211(csa_tree_add_6_33_groupi_n_861 ,csa_tree_add_6_33_groupi_n_1017);
  not csa_tree_add_6_33_groupi_drc_bufs18214(csa_tree_add_6_33_groupi_n_860 ,csa_tree_add_6_33_groupi_n_1008);
  not csa_tree_add_6_33_groupi_drc_bufs18215(csa_tree_add_6_33_groupi_n_859 ,csa_tree_add_6_33_groupi_n_1008);
  not csa_tree_add_6_33_groupi_drc_bufs18218(csa_tree_add_6_33_groupi_n_858 ,csa_tree_add_6_33_groupi_n_1027);
  not csa_tree_add_6_33_groupi_drc_bufs18219(csa_tree_add_6_33_groupi_n_857 ,csa_tree_add_6_33_groupi_n_1027);
  not csa_tree_add_6_33_groupi_drc_bufs18222(csa_tree_add_6_33_groupi_n_856 ,csa_tree_add_6_33_groupi_n_1035);
  not csa_tree_add_6_33_groupi_drc_bufs18223(csa_tree_add_6_33_groupi_n_855 ,csa_tree_add_6_33_groupi_n_1035);
  not csa_tree_add_6_33_groupi_drc_bufs18226(csa_tree_add_6_33_groupi_n_854 ,csa_tree_add_6_33_groupi_n_1012);
  not csa_tree_add_6_33_groupi_drc_bufs18227(csa_tree_add_6_33_groupi_n_853 ,csa_tree_add_6_33_groupi_n_1012);
  not csa_tree_add_6_33_groupi_drc_bufs18230(csa_tree_add_6_33_groupi_n_852 ,csa_tree_add_6_33_groupi_n_1015);
  not csa_tree_add_6_33_groupi_drc_bufs18231(csa_tree_add_6_33_groupi_n_851 ,csa_tree_add_6_33_groupi_n_1015);
  not csa_tree_add_6_33_groupi_drc_bufs18234(csa_tree_add_6_33_groupi_n_850 ,csa_tree_add_6_33_groupi_n_1023);
  not csa_tree_add_6_33_groupi_drc_bufs18235(csa_tree_add_6_33_groupi_n_849 ,csa_tree_add_6_33_groupi_n_1023);
  not csa_tree_add_6_33_groupi_drc_bufs18238(csa_tree_add_6_33_groupi_n_848 ,csa_tree_add_6_33_groupi_n_1020);
  not csa_tree_add_6_33_groupi_drc_bufs18239(csa_tree_add_6_33_groupi_n_847 ,csa_tree_add_6_33_groupi_n_1020);
  not csa_tree_add_6_33_groupi_drc_bufs18242(csa_tree_add_6_33_groupi_n_846 ,csa_tree_add_6_33_groupi_n_1028);
  not csa_tree_add_6_33_groupi_drc_bufs18243(csa_tree_add_6_33_groupi_n_845 ,csa_tree_add_6_33_groupi_n_1028);
  not csa_tree_add_6_33_groupi_drc_bufs18246(csa_tree_add_6_33_groupi_n_844 ,csa_tree_add_6_33_groupi_n_1029);
  not csa_tree_add_6_33_groupi_drc_bufs18247(csa_tree_add_6_33_groupi_n_843 ,csa_tree_add_6_33_groupi_n_1029);
  not csa_tree_add_6_33_groupi_drc_bufs18250(csa_tree_add_6_33_groupi_n_842 ,csa_tree_add_6_33_groupi_n_1040);
  not csa_tree_add_6_33_groupi_drc_bufs18251(csa_tree_add_6_33_groupi_n_841 ,csa_tree_add_6_33_groupi_n_1040);
  not csa_tree_add_6_33_groupi_drc_bufs18254(csa_tree_add_6_33_groupi_n_840 ,csa_tree_add_6_33_groupi_n_1036);
  not csa_tree_add_6_33_groupi_drc_bufs18255(csa_tree_add_6_33_groupi_n_839 ,csa_tree_add_6_33_groupi_n_1036);
  not csa_tree_add_6_33_groupi_drc_bufs18258(csa_tree_add_6_33_groupi_n_838 ,csa_tree_add_6_33_groupi_n_1032);
  not csa_tree_add_6_33_groupi_drc_bufs18259(csa_tree_add_6_33_groupi_n_837 ,csa_tree_add_6_33_groupi_n_1032);
  not csa_tree_add_6_33_groupi_drc_bufs18262(csa_tree_add_6_33_groupi_n_836 ,csa_tree_add_6_33_groupi_n_1018);
  not csa_tree_add_6_33_groupi_drc_bufs18263(csa_tree_add_6_33_groupi_n_835 ,csa_tree_add_6_33_groupi_n_1018);
  not csa_tree_add_6_33_groupi_drc_bufs18266(csa_tree_add_6_33_groupi_n_834 ,csa_tree_add_6_33_groupi_n_1019);
  not csa_tree_add_6_33_groupi_drc_bufs18267(csa_tree_add_6_33_groupi_n_833 ,csa_tree_add_6_33_groupi_n_1019);
  not csa_tree_add_6_33_groupi_drc_bufs18270(csa_tree_add_6_33_groupi_n_832 ,csa_tree_add_6_33_groupi_n_1033);
  not csa_tree_add_6_33_groupi_drc_bufs18271(csa_tree_add_6_33_groupi_n_831 ,csa_tree_add_6_33_groupi_n_1033);
  not csa_tree_add_6_33_groupi_drc_bufs18274(csa_tree_add_6_33_groupi_n_830 ,csa_tree_add_6_33_groupi_n_1034);
  not csa_tree_add_6_33_groupi_drc_bufs18275(csa_tree_add_6_33_groupi_n_829 ,csa_tree_add_6_33_groupi_n_1034);
  not csa_tree_add_6_33_groupi_drc_bufs18278(csa_tree_add_6_33_groupi_n_828 ,csa_tree_add_6_33_groupi_n_1038);
  not csa_tree_add_6_33_groupi_drc_bufs18279(csa_tree_add_6_33_groupi_n_827 ,csa_tree_add_6_33_groupi_n_1038);
  not csa_tree_add_6_33_groupi_drc_bufs18282(csa_tree_add_6_33_groupi_n_826 ,csa_tree_add_6_33_groupi_n_1025);
  not csa_tree_add_6_33_groupi_drc_bufs18283(csa_tree_add_6_33_groupi_n_825 ,csa_tree_add_6_33_groupi_n_1025);
  not csa_tree_add_6_33_groupi_drc_bufs18286(csa_tree_add_6_33_groupi_n_824 ,csa_tree_add_6_33_groupi_n_1037);
  not csa_tree_add_6_33_groupi_drc_bufs18287(csa_tree_add_6_33_groupi_n_823 ,csa_tree_add_6_33_groupi_n_1037);
  not csa_tree_add_6_33_groupi_drc_bufs18290(csa_tree_add_6_33_groupi_n_822 ,csa_tree_add_6_33_groupi_n_1021);
  not csa_tree_add_6_33_groupi_drc_bufs18291(csa_tree_add_6_33_groupi_n_821 ,csa_tree_add_6_33_groupi_n_1021);
  not csa_tree_add_6_33_groupi_drc_bufs18294(csa_tree_add_6_33_groupi_n_820 ,csa_tree_add_6_33_groupi_n_1013);
  not csa_tree_add_6_33_groupi_drc_bufs18295(csa_tree_add_6_33_groupi_n_819 ,csa_tree_add_6_33_groupi_n_1013);
  not csa_tree_add_6_33_groupi_drc_bufs18298(csa_tree_add_6_33_groupi_n_818 ,csa_tree_add_6_33_groupi_n_1016);
  not csa_tree_add_6_33_groupi_drc_bufs18299(csa_tree_add_6_33_groupi_n_817 ,csa_tree_add_6_33_groupi_n_1016);
  not csa_tree_add_6_33_groupi_drc_bufs18302(csa_tree_add_6_33_groupi_n_816 ,csa_tree_add_6_33_groupi_n_1039);
  not csa_tree_add_6_33_groupi_drc_bufs18303(csa_tree_add_6_33_groupi_n_815 ,csa_tree_add_6_33_groupi_n_1039);
  not csa_tree_add_6_33_groupi_drc_bufs18306(csa_tree_add_6_33_groupi_n_814 ,csa_tree_add_6_33_groupi_n_1014);
  not csa_tree_add_6_33_groupi_drc_bufs18307(csa_tree_add_6_33_groupi_n_813 ,csa_tree_add_6_33_groupi_n_1014);
  not csa_tree_add_6_33_groupi_drc_bufs18310(csa_tree_add_6_33_groupi_n_812 ,csa_tree_add_6_33_groupi_n_810);
  not csa_tree_add_6_33_groupi_drc_bufs18311(csa_tree_add_6_33_groupi_n_811 ,csa_tree_add_6_33_groupi_n_810);
  not csa_tree_add_6_33_groupi_drc_bufs18312(csa_tree_add_6_33_groupi_n_810 ,csa_tree_add_6_33_groupi_n_1004);
  not csa_tree_add_6_33_groupi_drc_bufs18314(csa_tree_add_6_33_groupi_n_809 ,csa_tree_add_6_33_groupi_n_807);
  not csa_tree_add_6_33_groupi_drc_bufs18315(csa_tree_add_6_33_groupi_n_808 ,csa_tree_add_6_33_groupi_n_807);
  not csa_tree_add_6_33_groupi_drc_bufs18316(csa_tree_add_6_33_groupi_n_807 ,csa_tree_add_6_33_groupi_n_993);
  not csa_tree_add_6_33_groupi_drc_bufs18318(csa_tree_add_6_33_groupi_n_806 ,csa_tree_add_6_33_groupi_n_804);
  not csa_tree_add_6_33_groupi_drc_bufs18319(csa_tree_add_6_33_groupi_n_805 ,csa_tree_add_6_33_groupi_n_804);
  not csa_tree_add_6_33_groupi_drc_bufs18320(csa_tree_add_6_33_groupi_n_804 ,csa_tree_add_6_33_groupi_n_977);
  not csa_tree_add_6_33_groupi_drc_bufs18322(csa_tree_add_6_33_groupi_n_803 ,csa_tree_add_6_33_groupi_n_801);
  not csa_tree_add_6_33_groupi_drc_bufs18323(csa_tree_add_6_33_groupi_n_802 ,csa_tree_add_6_33_groupi_n_801);
  not csa_tree_add_6_33_groupi_drc_bufs18324(csa_tree_add_6_33_groupi_n_801 ,csa_tree_add_6_33_groupi_n_1001);
  not csa_tree_add_6_33_groupi_drc_bufs18326(csa_tree_add_6_33_groupi_n_800 ,csa_tree_add_6_33_groupi_n_798);
  not csa_tree_add_6_33_groupi_drc_bufs18327(csa_tree_add_6_33_groupi_n_799 ,csa_tree_add_6_33_groupi_n_798);
  not csa_tree_add_6_33_groupi_drc_bufs18328(csa_tree_add_6_33_groupi_n_798 ,csa_tree_add_6_33_groupi_n_985);
  not csa_tree_add_6_33_groupi_drc_bufs18330(csa_tree_add_6_33_groupi_n_797 ,csa_tree_add_6_33_groupi_n_795);
  not csa_tree_add_6_33_groupi_drc_bufs18331(csa_tree_add_6_33_groupi_n_796 ,csa_tree_add_6_33_groupi_n_795);
  not csa_tree_add_6_33_groupi_drc_bufs18332(csa_tree_add_6_33_groupi_n_795 ,csa_tree_add_6_33_groupi_n_989);
  not csa_tree_add_6_33_groupi_drc_bufs18334(csa_tree_add_6_33_groupi_n_794 ,csa_tree_add_6_33_groupi_n_792);
  not csa_tree_add_6_33_groupi_drc_bufs18335(csa_tree_add_6_33_groupi_n_793 ,csa_tree_add_6_33_groupi_n_792);
  not csa_tree_add_6_33_groupi_drc_bufs18336(csa_tree_add_6_33_groupi_n_792 ,csa_tree_add_6_33_groupi_n_965);
  not csa_tree_add_6_33_groupi_drc_bufs18338(csa_tree_add_6_33_groupi_n_791 ,csa_tree_add_6_33_groupi_n_789);
  not csa_tree_add_6_33_groupi_drc_bufs18339(csa_tree_add_6_33_groupi_n_790 ,csa_tree_add_6_33_groupi_n_789);
  not csa_tree_add_6_33_groupi_drc_bufs18340(csa_tree_add_6_33_groupi_n_789 ,csa_tree_add_6_33_groupi_n_981);
  not csa_tree_add_6_33_groupi_drc_bufs18342(csa_tree_add_6_33_groupi_n_788 ,csa_tree_add_6_33_groupi_n_786);
  not csa_tree_add_6_33_groupi_drc_bufs18343(csa_tree_add_6_33_groupi_n_787 ,csa_tree_add_6_33_groupi_n_786);
  not csa_tree_add_6_33_groupi_drc_bufs18344(csa_tree_add_6_33_groupi_n_786 ,csa_tree_add_6_33_groupi_n_997);
  not csa_tree_add_6_33_groupi_drc_bufs18346(csa_tree_add_6_33_groupi_n_785 ,csa_tree_add_6_33_groupi_n_783);
  not csa_tree_add_6_33_groupi_drc_bufs18347(csa_tree_add_6_33_groupi_n_784 ,csa_tree_add_6_33_groupi_n_783);
  not csa_tree_add_6_33_groupi_drc_bufs18348(csa_tree_add_6_33_groupi_n_783 ,csa_tree_add_6_33_groupi_n_973);
  not csa_tree_add_6_33_groupi_drc_bufs18350(csa_tree_add_6_33_groupi_n_782 ,csa_tree_add_6_33_groupi_n_780);
  not csa_tree_add_6_33_groupi_drc_bufs18351(csa_tree_add_6_33_groupi_n_781 ,csa_tree_add_6_33_groupi_n_780);
  not csa_tree_add_6_33_groupi_drc_bufs18352(csa_tree_add_6_33_groupi_n_780 ,csa_tree_add_6_33_groupi_n_961);
  not csa_tree_add_6_33_groupi_drc_bufs18354(csa_tree_add_6_33_groupi_n_779 ,csa_tree_add_6_33_groupi_n_777);
  not csa_tree_add_6_33_groupi_drc_bufs18355(csa_tree_add_6_33_groupi_n_778 ,csa_tree_add_6_33_groupi_n_777);
  not csa_tree_add_6_33_groupi_drc_bufs18356(csa_tree_add_6_33_groupi_n_777 ,csa_tree_add_6_33_groupi_n_957);
  not csa_tree_add_6_33_groupi_drc_bufs18358(csa_tree_add_6_33_groupi_n_776 ,csa_tree_add_6_33_groupi_n_774);
  not csa_tree_add_6_33_groupi_drc_bufs18359(csa_tree_add_6_33_groupi_n_775 ,csa_tree_add_6_33_groupi_n_774);
  not csa_tree_add_6_33_groupi_drc_bufs18360(csa_tree_add_6_33_groupi_n_774 ,csa_tree_add_6_33_groupi_n_953);
  not csa_tree_add_6_33_groupi_drc_bufs18362(csa_tree_add_6_33_groupi_n_773 ,csa_tree_add_6_33_groupi_n_771);
  not csa_tree_add_6_33_groupi_drc_bufs18363(csa_tree_add_6_33_groupi_n_772 ,csa_tree_add_6_33_groupi_n_771);
  not csa_tree_add_6_33_groupi_drc_bufs18364(csa_tree_add_6_33_groupi_n_771 ,csa_tree_add_6_33_groupi_n_969);
  not csa_tree_add_6_33_groupi_drc_bufs18366(csa_tree_add_6_33_groupi_n_770 ,csa_tree_add_6_33_groupi_n_768);
  not csa_tree_add_6_33_groupi_drc_bufs18367(csa_tree_add_6_33_groupi_n_769 ,csa_tree_add_6_33_groupi_n_768);
  not csa_tree_add_6_33_groupi_drc_bufs18368(csa_tree_add_6_33_groupi_n_768 ,csa_tree_add_6_33_groupi_n_1005);
  not csa_tree_add_6_33_groupi_drc_bufs18370(csa_tree_add_6_33_groupi_n_767 ,csa_tree_add_6_33_groupi_n_765);
  not csa_tree_add_6_33_groupi_drc_bufs18371(csa_tree_add_6_33_groupi_n_766 ,csa_tree_add_6_33_groupi_n_765);
  not csa_tree_add_6_33_groupi_drc_bufs18372(csa_tree_add_6_33_groupi_n_765 ,csa_tree_add_6_33_groupi_n_969);
  not csa_tree_add_6_33_groupi_drc_bufs18374(csa_tree_add_6_33_groupi_n_764 ,csa_tree_add_6_33_groupi_n_762);
  not csa_tree_add_6_33_groupi_drc_bufs18375(csa_tree_add_6_33_groupi_n_763 ,csa_tree_add_6_33_groupi_n_762);
  not csa_tree_add_6_33_groupi_drc_bufs18376(csa_tree_add_6_33_groupi_n_762 ,csa_tree_add_6_33_groupi_n_889);
  not csa_tree_add_6_33_groupi_drc_bufs18378(csa_tree_add_6_33_groupi_n_761 ,csa_tree_add_6_33_groupi_n_759);
  not csa_tree_add_6_33_groupi_drc_bufs18379(csa_tree_add_6_33_groupi_n_760 ,csa_tree_add_6_33_groupi_n_759);
  not csa_tree_add_6_33_groupi_drc_bufs18380(csa_tree_add_6_33_groupi_n_759 ,csa_tree_add_6_33_groupi_n_893);
  not csa_tree_add_6_33_groupi_drc_bufs18382(csa_tree_add_6_33_groupi_n_758 ,csa_tree_add_6_33_groupi_n_756);
  not csa_tree_add_6_33_groupi_drc_bufs18383(csa_tree_add_6_33_groupi_n_757 ,csa_tree_add_6_33_groupi_n_756);
  not csa_tree_add_6_33_groupi_drc_bufs18384(csa_tree_add_6_33_groupi_n_756 ,csa_tree_add_6_33_groupi_n_918);
  not csa_tree_add_6_33_groupi_drc_bufs18386(csa_tree_add_6_33_groupi_n_755 ,csa_tree_add_6_33_groupi_n_753);
  not csa_tree_add_6_33_groupi_drc_bufs18387(csa_tree_add_6_33_groupi_n_754 ,csa_tree_add_6_33_groupi_n_753);
  not csa_tree_add_6_33_groupi_drc_bufs18388(csa_tree_add_6_33_groupi_n_753 ,csa_tree_add_6_33_groupi_n_927);
  not csa_tree_add_6_33_groupi_drc_bufs18390(csa_tree_add_6_33_groupi_n_752 ,csa_tree_add_6_33_groupi_n_750);
  not csa_tree_add_6_33_groupi_drc_bufs18391(csa_tree_add_6_33_groupi_n_751 ,csa_tree_add_6_33_groupi_n_750);
  not csa_tree_add_6_33_groupi_drc_bufs18392(csa_tree_add_6_33_groupi_n_750 ,csa_tree_add_6_33_groupi_n_922);
  not csa_tree_add_6_33_groupi_drc_bufs18394(csa_tree_add_6_33_groupi_n_749 ,csa_tree_add_6_33_groupi_n_747);
  not csa_tree_add_6_33_groupi_drc_bufs18395(csa_tree_add_6_33_groupi_n_748 ,csa_tree_add_6_33_groupi_n_747);
  not csa_tree_add_6_33_groupi_drc_bufs18396(csa_tree_add_6_33_groupi_n_747 ,csa_tree_add_6_33_groupi_n_970);
  not csa_tree_add_6_33_groupi_drc_bufs18398(csa_tree_add_6_33_groupi_n_746 ,csa_tree_add_6_33_groupi_n_744);
  not csa_tree_add_6_33_groupi_drc_bufs18399(csa_tree_add_6_33_groupi_n_745 ,csa_tree_add_6_33_groupi_n_744);
  not csa_tree_add_6_33_groupi_drc_bufs18400(csa_tree_add_6_33_groupi_n_744 ,csa_tree_add_6_33_groupi_n_882);
  not csa_tree_add_6_33_groupi_drc_bufs18402(csa_tree_add_6_33_groupi_n_743 ,csa_tree_add_6_33_groupi_n_741);
  not csa_tree_add_6_33_groupi_drc_bufs18403(csa_tree_add_6_33_groupi_n_742 ,csa_tree_add_6_33_groupi_n_741);
  not csa_tree_add_6_33_groupi_drc_bufs18404(csa_tree_add_6_33_groupi_n_741 ,csa_tree_add_6_33_groupi_n_892);
  not csa_tree_add_6_33_groupi_drc_bufs18406(csa_tree_add_6_33_groupi_n_740 ,csa_tree_add_6_33_groupi_n_738);
  not csa_tree_add_6_33_groupi_drc_bufs18407(csa_tree_add_6_33_groupi_n_739 ,csa_tree_add_6_33_groupi_n_738);
  not csa_tree_add_6_33_groupi_drc_bufs18408(csa_tree_add_6_33_groupi_n_738 ,csa_tree_add_6_33_groupi_n_880);
  not csa_tree_add_6_33_groupi_drc_bufs18410(csa_tree_add_6_33_groupi_n_737 ,csa_tree_add_6_33_groupi_n_735);
  not csa_tree_add_6_33_groupi_drc_bufs18411(csa_tree_add_6_33_groupi_n_736 ,csa_tree_add_6_33_groupi_n_735);
  not csa_tree_add_6_33_groupi_drc_bufs18412(csa_tree_add_6_33_groupi_n_735 ,csa_tree_add_6_33_groupi_n_970);
  not csa_tree_add_6_33_groupi_drc_bufs18414(csa_tree_add_6_33_groupi_n_734 ,csa_tree_add_6_33_groupi_n_732);
  not csa_tree_add_6_33_groupi_drc_bufs18415(csa_tree_add_6_33_groupi_n_733 ,csa_tree_add_6_33_groupi_n_732);
  not csa_tree_add_6_33_groupi_drc_bufs18416(csa_tree_add_6_33_groupi_n_732 ,csa_tree_add_6_33_groupi_n_884);
  not csa_tree_add_6_33_groupi_drc_bufs18418(csa_tree_add_6_33_groupi_n_731 ,csa_tree_add_6_33_groupi_n_729);
  not csa_tree_add_6_33_groupi_drc_bufs18419(csa_tree_add_6_33_groupi_n_730 ,csa_tree_add_6_33_groupi_n_729);
  not csa_tree_add_6_33_groupi_drc_bufs18420(csa_tree_add_6_33_groupi_n_729 ,csa_tree_add_6_33_groupi_n_935);
  not csa_tree_add_6_33_groupi_drc_bufs18422(csa_tree_add_6_33_groupi_n_728 ,csa_tree_add_6_33_groupi_n_726);
  not csa_tree_add_6_33_groupi_drc_bufs18423(csa_tree_add_6_33_groupi_n_727 ,csa_tree_add_6_33_groupi_n_726);
  not csa_tree_add_6_33_groupi_drc_bufs18424(csa_tree_add_6_33_groupi_n_726 ,csa_tree_add_6_33_groupi_n_930);
  not csa_tree_add_6_33_groupi_drc_bufs18426(csa_tree_add_6_33_groupi_n_725 ,csa_tree_add_6_33_groupi_n_723);
  not csa_tree_add_6_33_groupi_drc_bufs18427(csa_tree_add_6_33_groupi_n_724 ,csa_tree_add_6_33_groupi_n_723);
  not csa_tree_add_6_33_groupi_drc_bufs18428(csa_tree_add_6_33_groupi_n_723 ,csa_tree_add_6_33_groupi_n_1002);
  not csa_tree_add_6_33_groupi_drc_bufs18430(csa_tree_add_6_33_groupi_n_722 ,csa_tree_add_6_33_groupi_n_720);
  not csa_tree_add_6_33_groupi_drc_bufs18431(csa_tree_add_6_33_groupi_n_721 ,csa_tree_add_6_33_groupi_n_720);
  not csa_tree_add_6_33_groupi_drc_bufs18432(csa_tree_add_6_33_groupi_n_720 ,csa_tree_add_6_33_groupi_n_914);
  not csa_tree_add_6_33_groupi_drc_bufs18434(csa_tree_add_6_33_groupi_n_719 ,csa_tree_add_6_33_groupi_n_717);
  not csa_tree_add_6_33_groupi_drc_bufs18435(csa_tree_add_6_33_groupi_n_718 ,csa_tree_add_6_33_groupi_n_717);
  not csa_tree_add_6_33_groupi_drc_bufs18436(csa_tree_add_6_33_groupi_n_717 ,csa_tree_add_6_33_groupi_n_892);
  not csa_tree_add_6_33_groupi_drc_bufs18438(csa_tree_add_6_33_groupi_n_716 ,csa_tree_add_6_33_groupi_n_714);
  not csa_tree_add_6_33_groupi_drc_bufs18439(csa_tree_add_6_33_groupi_n_715 ,csa_tree_add_6_33_groupi_n_714);
  not csa_tree_add_6_33_groupi_drc_bufs18440(csa_tree_add_6_33_groupi_n_714 ,csa_tree_add_6_33_groupi_n_935);
  not csa_tree_add_6_33_groupi_drc_bufs18442(csa_tree_add_6_33_groupi_n_713 ,csa_tree_add_6_33_groupi_n_711);
  not csa_tree_add_6_33_groupi_drc_bufs18443(csa_tree_add_6_33_groupi_n_712 ,csa_tree_add_6_33_groupi_n_711);
  not csa_tree_add_6_33_groupi_drc_bufs18444(csa_tree_add_6_33_groupi_n_711 ,csa_tree_add_6_33_groupi_n_933);
  not csa_tree_add_6_33_groupi_drc_bufs18446(csa_tree_add_6_33_groupi_n_710 ,csa_tree_add_6_33_groupi_n_708);
  not csa_tree_add_6_33_groupi_drc_bufs18447(csa_tree_add_6_33_groupi_n_709 ,csa_tree_add_6_33_groupi_n_708);
  not csa_tree_add_6_33_groupi_drc_bufs18448(csa_tree_add_6_33_groupi_n_708 ,csa_tree_add_6_33_groupi_n_878);
  not csa_tree_add_6_33_groupi_drc_bufs18450(csa_tree_add_6_33_groupi_n_707 ,csa_tree_add_6_33_groupi_n_705);
  not csa_tree_add_6_33_groupi_drc_bufs18451(csa_tree_add_6_33_groupi_n_706 ,csa_tree_add_6_33_groupi_n_705);
  not csa_tree_add_6_33_groupi_drc_bufs18452(csa_tree_add_6_33_groupi_n_705 ,csa_tree_add_6_33_groupi_n_998);
  not csa_tree_add_6_33_groupi_drc_bufs18454(csa_tree_add_6_33_groupi_n_704 ,csa_tree_add_6_33_groupi_n_702);
  not csa_tree_add_6_33_groupi_drc_bufs18455(csa_tree_add_6_33_groupi_n_703 ,csa_tree_add_6_33_groupi_n_702);
  not csa_tree_add_6_33_groupi_drc_bufs18456(csa_tree_add_6_33_groupi_n_702 ,csa_tree_add_6_33_groupi_n_898);
  not csa_tree_add_6_33_groupi_drc_bufs18458(csa_tree_add_6_33_groupi_n_701 ,csa_tree_add_6_33_groupi_n_699);
  not csa_tree_add_6_33_groupi_drc_bufs18459(csa_tree_add_6_33_groupi_n_700 ,csa_tree_add_6_33_groupi_n_699);
  not csa_tree_add_6_33_groupi_drc_bufs18460(csa_tree_add_6_33_groupi_n_699 ,csa_tree_add_6_33_groupi_n_933);
  not csa_tree_add_6_33_groupi_drc_bufs18462(csa_tree_add_6_33_groupi_n_698 ,csa_tree_add_6_33_groupi_n_696);
  not csa_tree_add_6_33_groupi_drc_bufs18463(csa_tree_add_6_33_groupi_n_697 ,csa_tree_add_6_33_groupi_n_696);
  not csa_tree_add_6_33_groupi_drc_bufs18464(csa_tree_add_6_33_groupi_n_696 ,csa_tree_add_6_33_groupi_n_894);
  not csa_tree_add_6_33_groupi_drc_bufs18466(csa_tree_add_6_33_groupi_n_695 ,csa_tree_add_6_33_groupi_n_693);
  not csa_tree_add_6_33_groupi_drc_bufs18467(csa_tree_add_6_33_groupi_n_694 ,csa_tree_add_6_33_groupi_n_693);
  not csa_tree_add_6_33_groupi_drc_bufs18468(csa_tree_add_6_33_groupi_n_693 ,csa_tree_add_6_33_groupi_n_988);
  not csa_tree_add_6_33_groupi_drc_bufs18470(csa_tree_add_6_33_groupi_n_692 ,csa_tree_add_6_33_groupi_n_690);
  not csa_tree_add_6_33_groupi_drc_bufs18471(csa_tree_add_6_33_groupi_n_691 ,csa_tree_add_6_33_groupi_n_690);
  not csa_tree_add_6_33_groupi_drc_bufs18472(csa_tree_add_6_33_groupi_n_690 ,csa_tree_add_6_33_groupi_n_895);
  not csa_tree_add_6_33_groupi_drc_bufs18474(csa_tree_add_6_33_groupi_n_689 ,csa_tree_add_6_33_groupi_n_687);
  not csa_tree_add_6_33_groupi_drc_bufs18475(csa_tree_add_6_33_groupi_n_688 ,csa_tree_add_6_33_groupi_n_687);
  not csa_tree_add_6_33_groupi_drc_bufs18476(csa_tree_add_6_33_groupi_n_687 ,csa_tree_add_6_33_groupi_n_953);
  not csa_tree_add_6_33_groupi_drc_bufs18478(csa_tree_add_6_33_groupi_n_686 ,csa_tree_add_6_33_groupi_n_684);
  not csa_tree_add_6_33_groupi_drc_bufs18479(csa_tree_add_6_33_groupi_n_685 ,csa_tree_add_6_33_groupi_n_684);
  not csa_tree_add_6_33_groupi_drc_bufs18480(csa_tree_add_6_33_groupi_n_684 ,csa_tree_add_6_33_groupi_n_890);
  not csa_tree_add_6_33_groupi_drc_bufs18482(csa_tree_add_6_33_groupi_n_683 ,csa_tree_add_6_33_groupi_n_681);
  not csa_tree_add_6_33_groupi_drc_bufs18483(csa_tree_add_6_33_groupi_n_682 ,csa_tree_add_6_33_groupi_n_681);
  not csa_tree_add_6_33_groupi_drc_bufs18484(csa_tree_add_6_33_groupi_n_681 ,csa_tree_add_6_33_groupi_n_1002);
  not csa_tree_add_6_33_groupi_drc_bufs18486(csa_tree_add_6_33_groupi_n_680 ,csa_tree_add_6_33_groupi_n_678);
  not csa_tree_add_6_33_groupi_drc_bufs18487(csa_tree_add_6_33_groupi_n_679 ,csa_tree_add_6_33_groupi_n_678);
  not csa_tree_add_6_33_groupi_drc_bufs18488(csa_tree_add_6_33_groupi_n_678 ,csa_tree_add_6_33_groupi_n_879);
  not csa_tree_add_6_33_groupi_drc_bufs18490(csa_tree_add_6_33_groupi_n_677 ,csa_tree_add_6_33_groupi_n_675);
  not csa_tree_add_6_33_groupi_drc_bufs18491(csa_tree_add_6_33_groupi_n_676 ,csa_tree_add_6_33_groupi_n_675);
  not csa_tree_add_6_33_groupi_drc_bufs18492(csa_tree_add_6_33_groupi_n_675 ,csa_tree_add_6_33_groupi_n_998);
  not csa_tree_add_6_33_groupi_drc_bufs18494(csa_tree_add_6_33_groupi_n_674 ,csa_tree_add_6_33_groupi_n_672);
  not csa_tree_add_6_33_groupi_drc_bufs18495(csa_tree_add_6_33_groupi_n_673 ,csa_tree_add_6_33_groupi_n_672);
  not csa_tree_add_6_33_groupi_drc_bufs18496(csa_tree_add_6_33_groupi_n_672 ,csa_tree_add_6_33_groupi_n_902);
  not csa_tree_add_6_33_groupi_drc_bufs18498(csa_tree_add_6_33_groupi_n_671 ,csa_tree_add_6_33_groupi_n_669);
  not csa_tree_add_6_33_groupi_drc_bufs18499(csa_tree_add_6_33_groupi_n_670 ,csa_tree_add_6_33_groupi_n_669);
  not csa_tree_add_6_33_groupi_drc_bufs18500(csa_tree_add_6_33_groupi_n_669 ,csa_tree_add_6_33_groupi_n_988);
  not csa_tree_add_6_33_groupi_drc_bufs18502(csa_tree_add_6_33_groupi_n_668 ,csa_tree_add_6_33_groupi_n_666);
  not csa_tree_add_6_33_groupi_drc_bufs18503(csa_tree_add_6_33_groupi_n_667 ,csa_tree_add_6_33_groupi_n_666);
  not csa_tree_add_6_33_groupi_drc_bufs18504(csa_tree_add_6_33_groupi_n_666 ,csa_tree_add_6_33_groupi_n_987);
  not csa_tree_add_6_33_groupi_drc_bufs18506(csa_tree_add_6_33_groupi_n_665 ,csa_tree_add_6_33_groupi_n_663);
  not csa_tree_add_6_33_groupi_drc_bufs18507(csa_tree_add_6_33_groupi_n_664 ,csa_tree_add_6_33_groupi_n_663);
  not csa_tree_add_6_33_groupi_drc_bufs18508(csa_tree_add_6_33_groupi_n_663 ,csa_tree_add_6_33_groupi_n_904);
  not csa_tree_add_6_33_groupi_drc_bufs18510(csa_tree_add_6_33_groupi_n_662 ,csa_tree_add_6_33_groupi_n_660);
  not csa_tree_add_6_33_groupi_drc_bufs18511(csa_tree_add_6_33_groupi_n_661 ,csa_tree_add_6_33_groupi_n_660);
  not csa_tree_add_6_33_groupi_drc_bufs18512(csa_tree_add_6_33_groupi_n_660 ,csa_tree_add_6_33_groupi_n_888);
  not csa_tree_add_6_33_groupi_drc_bufs18514(csa_tree_add_6_33_groupi_n_659 ,csa_tree_add_6_33_groupi_n_657);
  not csa_tree_add_6_33_groupi_drc_bufs18515(csa_tree_add_6_33_groupi_n_658 ,csa_tree_add_6_33_groupi_n_657);
  not csa_tree_add_6_33_groupi_drc_bufs18516(csa_tree_add_6_33_groupi_n_657 ,csa_tree_add_6_33_groupi_n_909);
  not csa_tree_add_6_33_groupi_drc_bufs18518(csa_tree_add_6_33_groupi_n_656 ,csa_tree_add_6_33_groupi_n_654);
  not csa_tree_add_6_33_groupi_drc_bufs18519(csa_tree_add_6_33_groupi_n_655 ,csa_tree_add_6_33_groupi_n_654);
  not csa_tree_add_6_33_groupi_drc_bufs18520(csa_tree_add_6_33_groupi_n_654 ,csa_tree_add_6_33_groupi_n_987);
  not csa_tree_add_6_33_groupi_drc_bufs18522(csa_tree_add_6_33_groupi_n_653 ,csa_tree_add_6_33_groupi_n_651);
  not csa_tree_add_6_33_groupi_drc_bufs18523(csa_tree_add_6_33_groupi_n_652 ,csa_tree_add_6_33_groupi_n_651);
  not csa_tree_add_6_33_groupi_drc_bufs18524(csa_tree_add_6_33_groupi_n_651 ,csa_tree_add_6_33_groupi_n_881);
  not csa_tree_add_6_33_groupi_drc_bufs18526(csa_tree_add_6_33_groupi_n_650 ,csa_tree_add_6_33_groupi_n_648);
  not csa_tree_add_6_33_groupi_drc_bufs18527(csa_tree_add_6_33_groupi_n_649 ,csa_tree_add_6_33_groupi_n_648);
  not csa_tree_add_6_33_groupi_drc_bufs18528(csa_tree_add_6_33_groupi_n_648 ,csa_tree_add_6_33_groupi_n_932);
  not csa_tree_add_6_33_groupi_drc_bufs18530(csa_tree_add_6_33_groupi_n_647 ,csa_tree_add_6_33_groupi_n_645);
  not csa_tree_add_6_33_groupi_drc_bufs18531(csa_tree_add_6_33_groupi_n_646 ,csa_tree_add_6_33_groupi_n_645);
  not csa_tree_add_6_33_groupi_drc_bufs18532(csa_tree_add_6_33_groupi_n_645 ,csa_tree_add_6_33_groupi_n_913);
  not csa_tree_add_6_33_groupi_drc_bufs18534(csa_tree_add_6_33_groupi_n_644 ,csa_tree_add_6_33_groupi_n_642);
  not csa_tree_add_6_33_groupi_drc_bufs18535(csa_tree_add_6_33_groupi_n_643 ,csa_tree_add_6_33_groupi_n_642);
  not csa_tree_add_6_33_groupi_drc_bufs18536(csa_tree_add_6_33_groupi_n_642 ,csa_tree_add_6_33_groupi_n_980);
  not csa_tree_add_6_33_groupi_drc_bufs18538(csa_tree_add_6_33_groupi_n_641 ,csa_tree_add_6_33_groupi_n_639);
  not csa_tree_add_6_33_groupi_drc_bufs18539(csa_tree_add_6_33_groupi_n_640 ,csa_tree_add_6_33_groupi_n_639);
  not csa_tree_add_6_33_groupi_drc_bufs18540(csa_tree_add_6_33_groupi_n_639 ,csa_tree_add_6_33_groupi_n_955);
  not csa_tree_add_6_33_groupi_drc_bufs18542(csa_tree_add_6_33_groupi_n_638 ,csa_tree_add_6_33_groupi_n_636);
  not csa_tree_add_6_33_groupi_drc_bufs18543(csa_tree_add_6_33_groupi_n_637 ,csa_tree_add_6_33_groupi_n_636);
  not csa_tree_add_6_33_groupi_drc_bufs18544(csa_tree_add_6_33_groupi_n_636 ,csa_tree_add_6_33_groupi_n_955);
  not csa_tree_add_6_33_groupi_drc_bufs18546(csa_tree_add_6_33_groupi_n_635 ,csa_tree_add_6_33_groupi_n_633);
  not csa_tree_add_6_33_groupi_drc_bufs18547(csa_tree_add_6_33_groupi_n_634 ,csa_tree_add_6_33_groupi_n_633);
  not csa_tree_add_6_33_groupi_drc_bufs18548(csa_tree_add_6_33_groupi_n_633 ,csa_tree_add_6_33_groupi_n_956);
  not csa_tree_add_6_33_groupi_drc_bufs18550(csa_tree_add_6_33_groupi_n_632 ,csa_tree_add_6_33_groupi_n_630);
  not csa_tree_add_6_33_groupi_drc_bufs18551(csa_tree_add_6_33_groupi_n_631 ,csa_tree_add_6_33_groupi_n_630);
  not csa_tree_add_6_33_groupi_drc_bufs18552(csa_tree_add_6_33_groupi_n_630 ,csa_tree_add_6_33_groupi_n_956);
  not csa_tree_add_6_33_groupi_drc_bufs18554(csa_tree_add_6_33_groupi_n_629 ,csa_tree_add_6_33_groupi_n_627);
  not csa_tree_add_6_33_groupi_drc_bufs18555(csa_tree_add_6_33_groupi_n_628 ,csa_tree_add_6_33_groupi_n_627);
  not csa_tree_add_6_33_groupi_drc_bufs18556(csa_tree_add_6_33_groupi_n_627 ,csa_tree_add_6_33_groupi_n_907);
  not csa_tree_add_6_33_groupi_drc_bufs18558(csa_tree_add_6_33_groupi_n_626 ,csa_tree_add_6_33_groupi_n_624);
  not csa_tree_add_6_33_groupi_drc_bufs18559(csa_tree_add_6_33_groupi_n_625 ,csa_tree_add_6_33_groupi_n_624);
  not csa_tree_add_6_33_groupi_drc_bufs18560(csa_tree_add_6_33_groupi_n_624 ,csa_tree_add_6_33_groupi_n_907);
  not csa_tree_add_6_33_groupi_drc_bufs18562(csa_tree_add_6_33_groupi_n_623 ,csa_tree_add_6_33_groupi_n_621);
  not csa_tree_add_6_33_groupi_drc_bufs18563(csa_tree_add_6_33_groupi_n_622 ,csa_tree_add_6_33_groupi_n_621);
  not csa_tree_add_6_33_groupi_drc_bufs18564(csa_tree_add_6_33_groupi_n_621 ,csa_tree_add_6_33_groupi_n_908);
  not csa_tree_add_6_33_groupi_drc_bufs18566(csa_tree_add_6_33_groupi_n_620 ,csa_tree_add_6_33_groupi_n_618);
  not csa_tree_add_6_33_groupi_drc_bufs18567(csa_tree_add_6_33_groupi_n_619 ,csa_tree_add_6_33_groupi_n_618);
  not csa_tree_add_6_33_groupi_drc_bufs18568(csa_tree_add_6_33_groupi_n_618 ,csa_tree_add_6_33_groupi_n_908);
  not csa_tree_add_6_33_groupi_drc_bufs18570(csa_tree_add_6_33_groupi_n_617 ,csa_tree_add_6_33_groupi_n_615);
  not csa_tree_add_6_33_groupi_drc_bufs18571(csa_tree_add_6_33_groupi_n_616 ,csa_tree_add_6_33_groupi_n_615);
  not csa_tree_add_6_33_groupi_drc_bufs18572(csa_tree_add_6_33_groupi_n_615 ,csa_tree_add_6_33_groupi_n_1000);
  not csa_tree_add_6_33_groupi_drc_bufs18574(csa_tree_add_6_33_groupi_n_614 ,csa_tree_add_6_33_groupi_n_612);
  not csa_tree_add_6_33_groupi_drc_bufs18575(csa_tree_add_6_33_groupi_n_613 ,csa_tree_add_6_33_groupi_n_612);
  not csa_tree_add_6_33_groupi_drc_bufs18576(csa_tree_add_6_33_groupi_n_612 ,csa_tree_add_6_33_groupi_n_1000);
  not csa_tree_add_6_33_groupi_drc_bufs18578(csa_tree_add_6_33_groupi_n_611 ,csa_tree_add_6_33_groupi_n_609);
  not csa_tree_add_6_33_groupi_drc_bufs18579(csa_tree_add_6_33_groupi_n_610 ,csa_tree_add_6_33_groupi_n_609);
  not csa_tree_add_6_33_groupi_drc_bufs18580(csa_tree_add_6_33_groupi_n_609 ,csa_tree_add_6_33_groupi_n_958);
  not csa_tree_add_6_33_groupi_drc_bufs18582(csa_tree_add_6_33_groupi_n_608 ,csa_tree_add_6_33_groupi_n_606);
  not csa_tree_add_6_33_groupi_drc_bufs18583(csa_tree_add_6_33_groupi_n_607 ,csa_tree_add_6_33_groupi_n_606);
  not csa_tree_add_6_33_groupi_drc_bufs18584(csa_tree_add_6_33_groupi_n_606 ,csa_tree_add_6_33_groupi_n_958);
  not csa_tree_add_6_33_groupi_drc_bufs18586(csa_tree_add_6_33_groupi_n_605 ,csa_tree_add_6_33_groupi_n_603);
  not csa_tree_add_6_33_groupi_drc_bufs18587(csa_tree_add_6_33_groupi_n_604 ,csa_tree_add_6_33_groupi_n_603);
  not csa_tree_add_6_33_groupi_drc_bufs18588(csa_tree_add_6_33_groupi_n_603 ,csa_tree_add_6_33_groupi_n_959);
  not csa_tree_add_6_33_groupi_drc_bufs18590(csa_tree_add_6_33_groupi_n_602 ,csa_tree_add_6_33_groupi_n_600);
  not csa_tree_add_6_33_groupi_drc_bufs18591(csa_tree_add_6_33_groupi_n_601 ,csa_tree_add_6_33_groupi_n_600);
  not csa_tree_add_6_33_groupi_drc_bufs18592(csa_tree_add_6_33_groupi_n_600 ,csa_tree_add_6_33_groupi_n_959);
  not csa_tree_add_6_33_groupi_drc_bufs18594(csa_tree_add_6_33_groupi_n_599 ,csa_tree_add_6_33_groupi_n_597);
  not csa_tree_add_6_33_groupi_drc_bufs18595(csa_tree_add_6_33_groupi_n_598 ,csa_tree_add_6_33_groupi_n_597);
  not csa_tree_add_6_33_groupi_drc_bufs18596(csa_tree_add_6_33_groupi_n_597 ,csa_tree_add_6_33_groupi_n_982);
  not csa_tree_add_6_33_groupi_drc_bufs18598(csa_tree_add_6_33_groupi_n_596 ,csa_tree_add_6_33_groupi_n_594);
  not csa_tree_add_6_33_groupi_drc_bufs18599(csa_tree_add_6_33_groupi_n_595 ,csa_tree_add_6_33_groupi_n_594);
  not csa_tree_add_6_33_groupi_drc_bufs18600(csa_tree_add_6_33_groupi_n_594 ,csa_tree_add_6_33_groupi_n_982);
  not csa_tree_add_6_33_groupi_drc_bufs18602(csa_tree_add_6_33_groupi_n_593 ,csa_tree_add_6_33_groupi_n_591);
  not csa_tree_add_6_33_groupi_drc_bufs18603(csa_tree_add_6_33_groupi_n_592 ,csa_tree_add_6_33_groupi_n_591);
  not csa_tree_add_6_33_groupi_drc_bufs18604(csa_tree_add_6_33_groupi_n_591 ,csa_tree_add_6_33_groupi_n_960);
  not csa_tree_add_6_33_groupi_drc_bufs18606(csa_tree_add_6_33_groupi_n_590 ,csa_tree_add_6_33_groupi_n_588);
  not csa_tree_add_6_33_groupi_drc_bufs18607(csa_tree_add_6_33_groupi_n_589 ,csa_tree_add_6_33_groupi_n_588);
  not csa_tree_add_6_33_groupi_drc_bufs18608(csa_tree_add_6_33_groupi_n_588 ,csa_tree_add_6_33_groupi_n_960);
  not csa_tree_add_6_33_groupi_drc_bufs18610(csa_tree_add_6_33_groupi_n_587 ,csa_tree_add_6_33_groupi_n_585);
  not csa_tree_add_6_33_groupi_drc_bufs18611(csa_tree_add_6_33_groupi_n_586 ,csa_tree_add_6_33_groupi_n_585);
  not csa_tree_add_6_33_groupi_drc_bufs18612(csa_tree_add_6_33_groupi_n_585 ,csa_tree_add_6_33_groupi_n_915);
  not csa_tree_add_6_33_groupi_drc_bufs18614(csa_tree_add_6_33_groupi_n_584 ,csa_tree_add_6_33_groupi_n_582);
  not csa_tree_add_6_33_groupi_drc_bufs18615(csa_tree_add_6_33_groupi_n_583 ,csa_tree_add_6_33_groupi_n_582);
  not csa_tree_add_6_33_groupi_drc_bufs18616(csa_tree_add_6_33_groupi_n_582 ,csa_tree_add_6_33_groupi_n_915);
  not csa_tree_add_6_33_groupi_drc_bufs18618(csa_tree_add_6_33_groupi_n_581 ,csa_tree_add_6_33_groupi_n_579);
  not csa_tree_add_6_33_groupi_drc_bufs18619(csa_tree_add_6_33_groupi_n_580 ,csa_tree_add_6_33_groupi_n_579);
  not csa_tree_add_6_33_groupi_drc_bufs18620(csa_tree_add_6_33_groupi_n_579 ,csa_tree_add_6_33_groupi_n_916);
  not csa_tree_add_6_33_groupi_drc_bufs18622(csa_tree_add_6_33_groupi_n_578 ,csa_tree_add_6_33_groupi_n_576);
  not csa_tree_add_6_33_groupi_drc_bufs18623(csa_tree_add_6_33_groupi_n_577 ,csa_tree_add_6_33_groupi_n_576);
  not csa_tree_add_6_33_groupi_drc_bufs18624(csa_tree_add_6_33_groupi_n_576 ,csa_tree_add_6_33_groupi_n_916);
  not csa_tree_add_6_33_groupi_drc_bufs18626(csa_tree_add_6_33_groupi_n_575 ,csa_tree_add_6_33_groupi_n_573);
  not csa_tree_add_6_33_groupi_drc_bufs18627(csa_tree_add_6_33_groupi_n_574 ,csa_tree_add_6_33_groupi_n_573);
  not csa_tree_add_6_33_groupi_drc_bufs18628(csa_tree_add_6_33_groupi_n_573 ,csa_tree_add_6_33_groupi_n_983);
  not csa_tree_add_6_33_groupi_drc_bufs18630(csa_tree_add_6_33_groupi_n_572 ,csa_tree_add_6_33_groupi_n_570);
  not csa_tree_add_6_33_groupi_drc_bufs18631(csa_tree_add_6_33_groupi_n_571 ,csa_tree_add_6_33_groupi_n_570);
  not csa_tree_add_6_33_groupi_drc_bufs18632(csa_tree_add_6_33_groupi_n_570 ,csa_tree_add_6_33_groupi_n_983);
  not csa_tree_add_6_33_groupi_drc_bufs18634(csa_tree_add_6_33_groupi_n_569 ,csa_tree_add_6_33_groupi_n_567);
  not csa_tree_add_6_33_groupi_drc_bufs18635(csa_tree_add_6_33_groupi_n_568 ,csa_tree_add_6_33_groupi_n_567);
  not csa_tree_add_6_33_groupi_drc_bufs18636(csa_tree_add_6_33_groupi_n_567 ,csa_tree_add_6_33_groupi_n_904);
  not csa_tree_add_6_33_groupi_drc_bufs18638(csa_tree_add_6_33_groupi_n_566 ,csa_tree_add_6_33_groupi_n_564);
  not csa_tree_add_6_33_groupi_drc_bufs18639(csa_tree_add_6_33_groupi_n_565 ,csa_tree_add_6_33_groupi_n_564);
  not csa_tree_add_6_33_groupi_drc_bufs18640(csa_tree_add_6_33_groupi_n_564 ,csa_tree_add_6_33_groupi_n_994);
  not csa_tree_add_6_33_groupi_drc_bufs18642(csa_tree_add_6_33_groupi_n_563 ,csa_tree_add_6_33_groupi_n_561);
  not csa_tree_add_6_33_groupi_drc_bufs18643(csa_tree_add_6_33_groupi_n_562 ,csa_tree_add_6_33_groupi_n_561);
  not csa_tree_add_6_33_groupi_drc_bufs18644(csa_tree_add_6_33_groupi_n_561 ,csa_tree_add_6_33_groupi_n_917);
  not csa_tree_add_6_33_groupi_drc_bufs18646(csa_tree_add_6_33_groupi_n_560 ,csa_tree_add_6_33_groupi_n_558);
  not csa_tree_add_6_33_groupi_drc_bufs18647(csa_tree_add_6_33_groupi_n_559 ,csa_tree_add_6_33_groupi_n_558);
  not csa_tree_add_6_33_groupi_drc_bufs18648(csa_tree_add_6_33_groupi_n_558 ,csa_tree_add_6_33_groupi_n_917);
  not csa_tree_add_6_33_groupi_drc_bufs18650(csa_tree_add_6_33_groupi_n_557 ,csa_tree_add_6_33_groupi_n_555);
  not csa_tree_add_6_33_groupi_drc_bufs18651(csa_tree_add_6_33_groupi_n_556 ,csa_tree_add_6_33_groupi_n_555);
  not csa_tree_add_6_33_groupi_drc_bufs18652(csa_tree_add_6_33_groupi_n_555 ,csa_tree_add_6_33_groupi_n_962);
  not csa_tree_add_6_33_groupi_drc_bufs18654(csa_tree_add_6_33_groupi_n_554 ,csa_tree_add_6_33_groupi_n_552);
  not csa_tree_add_6_33_groupi_drc_bufs18655(csa_tree_add_6_33_groupi_n_553 ,csa_tree_add_6_33_groupi_n_552);
  not csa_tree_add_6_33_groupi_drc_bufs18656(csa_tree_add_6_33_groupi_n_552 ,csa_tree_add_6_33_groupi_n_962);
  not csa_tree_add_6_33_groupi_drc_bufs18658(csa_tree_add_6_33_groupi_n_551 ,csa_tree_add_6_33_groupi_n_549);
  not csa_tree_add_6_33_groupi_drc_bufs18659(csa_tree_add_6_33_groupi_n_550 ,csa_tree_add_6_33_groupi_n_549);
  not csa_tree_add_6_33_groupi_drc_bufs18660(csa_tree_add_6_33_groupi_n_549 ,csa_tree_add_6_33_groupi_n_984);
  not csa_tree_add_6_33_groupi_drc_bufs18662(csa_tree_add_6_33_groupi_n_548 ,csa_tree_add_6_33_groupi_n_546);
  not csa_tree_add_6_33_groupi_drc_bufs18663(csa_tree_add_6_33_groupi_n_547 ,csa_tree_add_6_33_groupi_n_546);
  not csa_tree_add_6_33_groupi_drc_bufs18664(csa_tree_add_6_33_groupi_n_546 ,csa_tree_add_6_33_groupi_n_984);
  not csa_tree_add_6_33_groupi_drc_bufs18666(csa_tree_add_6_33_groupi_n_545 ,csa_tree_add_6_33_groupi_n_543);
  not csa_tree_add_6_33_groupi_drc_bufs18667(csa_tree_add_6_33_groupi_n_544 ,csa_tree_add_6_33_groupi_n_543);
  not csa_tree_add_6_33_groupi_drc_bufs18668(csa_tree_add_6_33_groupi_n_543 ,csa_tree_add_6_33_groupi_n_963);
  not csa_tree_add_6_33_groupi_drc_bufs18670(csa_tree_add_6_33_groupi_n_542 ,csa_tree_add_6_33_groupi_n_540);
  not csa_tree_add_6_33_groupi_drc_bufs18671(csa_tree_add_6_33_groupi_n_541 ,csa_tree_add_6_33_groupi_n_540);
  not csa_tree_add_6_33_groupi_drc_bufs18672(csa_tree_add_6_33_groupi_n_540 ,csa_tree_add_6_33_groupi_n_963);
  not csa_tree_add_6_33_groupi_drc_bufs18674(csa_tree_add_6_33_groupi_n_539 ,csa_tree_add_6_33_groupi_n_537);
  not csa_tree_add_6_33_groupi_drc_bufs18675(csa_tree_add_6_33_groupi_n_538 ,csa_tree_add_6_33_groupi_n_537);
  not csa_tree_add_6_33_groupi_drc_bufs18676(csa_tree_add_6_33_groupi_n_537 ,csa_tree_add_6_33_groupi_n_964);
  not csa_tree_add_6_33_groupi_drc_bufs18678(csa_tree_add_6_33_groupi_n_536 ,csa_tree_add_6_33_groupi_n_534);
  not csa_tree_add_6_33_groupi_drc_bufs18679(csa_tree_add_6_33_groupi_n_535 ,csa_tree_add_6_33_groupi_n_534);
  not csa_tree_add_6_33_groupi_drc_bufs18680(csa_tree_add_6_33_groupi_n_534 ,csa_tree_add_6_33_groupi_n_964);
  not csa_tree_add_6_33_groupi_drc_bufs18682(csa_tree_add_6_33_groupi_n_533 ,csa_tree_add_6_33_groupi_n_531);
  not csa_tree_add_6_33_groupi_drc_bufs18683(csa_tree_add_6_33_groupi_n_532 ,csa_tree_add_6_33_groupi_n_531);
  not csa_tree_add_6_33_groupi_drc_bufs18684(csa_tree_add_6_33_groupi_n_531 ,csa_tree_add_6_33_groupi_n_995);
  not csa_tree_add_6_33_groupi_drc_bufs18686(csa_tree_add_6_33_groupi_n_530 ,csa_tree_add_6_33_groupi_n_528);
  not csa_tree_add_6_33_groupi_drc_bufs18687(csa_tree_add_6_33_groupi_n_529 ,csa_tree_add_6_33_groupi_n_528);
  not csa_tree_add_6_33_groupi_drc_bufs18688(csa_tree_add_6_33_groupi_n_528 ,csa_tree_add_6_33_groupi_n_995);
  not csa_tree_add_6_33_groupi_drc_bufs18690(csa_tree_add_6_33_groupi_n_527 ,csa_tree_add_6_33_groupi_n_525);
  not csa_tree_add_6_33_groupi_drc_bufs18691(csa_tree_add_6_33_groupi_n_526 ,csa_tree_add_6_33_groupi_n_525);
  not csa_tree_add_6_33_groupi_drc_bufs18692(csa_tree_add_6_33_groupi_n_525 ,csa_tree_add_6_33_groupi_n_1003);
  not csa_tree_add_6_33_groupi_drc_bufs18694(csa_tree_add_6_33_groupi_n_524 ,csa_tree_add_6_33_groupi_n_522);
  not csa_tree_add_6_33_groupi_drc_bufs18695(csa_tree_add_6_33_groupi_n_523 ,csa_tree_add_6_33_groupi_n_522);
  not csa_tree_add_6_33_groupi_drc_bufs18696(csa_tree_add_6_33_groupi_n_522 ,csa_tree_add_6_33_groupi_n_1003);
  not csa_tree_add_6_33_groupi_drc_bufs18698(csa_tree_add_6_33_groupi_n_521 ,csa_tree_add_6_33_groupi_n_519);
  not csa_tree_add_6_33_groupi_drc_bufs18699(csa_tree_add_6_33_groupi_n_520 ,csa_tree_add_6_33_groupi_n_519);
  not csa_tree_add_6_33_groupi_drc_bufs18700(csa_tree_add_6_33_groupi_n_519 ,csa_tree_add_6_33_groupi_n_924);
  not csa_tree_add_6_33_groupi_drc_bufs18702(csa_tree_add_6_33_groupi_n_518 ,csa_tree_add_6_33_groupi_n_516);
  not csa_tree_add_6_33_groupi_drc_bufs18703(csa_tree_add_6_33_groupi_n_517 ,csa_tree_add_6_33_groupi_n_516);
  not csa_tree_add_6_33_groupi_drc_bufs18704(csa_tree_add_6_33_groupi_n_516 ,csa_tree_add_6_33_groupi_n_924);
  not csa_tree_add_6_33_groupi_drc_bufs18706(csa_tree_add_6_33_groupi_n_515 ,csa_tree_add_6_33_groupi_n_513);
  not csa_tree_add_6_33_groupi_drc_bufs18707(csa_tree_add_6_33_groupi_n_514 ,csa_tree_add_6_33_groupi_n_513);
  not csa_tree_add_6_33_groupi_drc_bufs18708(csa_tree_add_6_33_groupi_n_513 ,csa_tree_add_6_33_groupi_n_925);
  not csa_tree_add_6_33_groupi_drc_bufs18710(csa_tree_add_6_33_groupi_n_512 ,csa_tree_add_6_33_groupi_n_510);
  not csa_tree_add_6_33_groupi_drc_bufs18711(csa_tree_add_6_33_groupi_n_511 ,csa_tree_add_6_33_groupi_n_510);
  not csa_tree_add_6_33_groupi_drc_bufs18712(csa_tree_add_6_33_groupi_n_510 ,csa_tree_add_6_33_groupi_n_925);
  not csa_tree_add_6_33_groupi_drc_bufs18714(csa_tree_add_6_33_groupi_n_509 ,csa_tree_add_6_33_groupi_n_507);
  not csa_tree_add_6_33_groupi_drc_bufs18715(csa_tree_add_6_33_groupi_n_508 ,csa_tree_add_6_33_groupi_n_507);
  not csa_tree_add_6_33_groupi_drc_bufs18716(csa_tree_add_6_33_groupi_n_507 ,csa_tree_add_6_33_groupi_n_996);
  not csa_tree_add_6_33_groupi_drc_bufs18718(csa_tree_add_6_33_groupi_n_506 ,csa_tree_add_6_33_groupi_n_504);
  not csa_tree_add_6_33_groupi_drc_bufs18719(csa_tree_add_6_33_groupi_n_505 ,csa_tree_add_6_33_groupi_n_504);
  not csa_tree_add_6_33_groupi_drc_bufs18720(csa_tree_add_6_33_groupi_n_504 ,csa_tree_add_6_33_groupi_n_996);
  not csa_tree_add_6_33_groupi_drc_bufs18722(csa_tree_add_6_33_groupi_n_503 ,csa_tree_add_6_33_groupi_n_501);
  not csa_tree_add_6_33_groupi_drc_bufs18723(csa_tree_add_6_33_groupi_n_502 ,csa_tree_add_6_33_groupi_n_501);
  not csa_tree_add_6_33_groupi_drc_bufs18724(csa_tree_add_6_33_groupi_n_501 ,csa_tree_add_6_33_groupi_n_966);
  not csa_tree_add_6_33_groupi_drc_bufs18726(csa_tree_add_6_33_groupi_n_500 ,csa_tree_add_6_33_groupi_n_498);
  not csa_tree_add_6_33_groupi_drc_bufs18727(csa_tree_add_6_33_groupi_n_499 ,csa_tree_add_6_33_groupi_n_498);
  not csa_tree_add_6_33_groupi_drc_bufs18728(csa_tree_add_6_33_groupi_n_498 ,csa_tree_add_6_33_groupi_n_966);
  not csa_tree_add_6_33_groupi_drc_bufs18730(csa_tree_add_6_33_groupi_n_497 ,csa_tree_add_6_33_groupi_n_495);
  not csa_tree_add_6_33_groupi_drc_bufs18731(csa_tree_add_6_33_groupi_n_496 ,csa_tree_add_6_33_groupi_n_495);
  not csa_tree_add_6_33_groupi_drc_bufs18732(csa_tree_add_6_33_groupi_n_495 ,csa_tree_add_6_33_groupi_n_928);
  not csa_tree_add_6_33_groupi_drc_bufs18734(csa_tree_add_6_33_groupi_n_494 ,csa_tree_add_6_33_groupi_n_492);
  not csa_tree_add_6_33_groupi_drc_bufs18735(csa_tree_add_6_33_groupi_n_493 ,csa_tree_add_6_33_groupi_n_492);
  not csa_tree_add_6_33_groupi_drc_bufs18736(csa_tree_add_6_33_groupi_n_492 ,csa_tree_add_6_33_groupi_n_928);
  not csa_tree_add_6_33_groupi_drc_bufs18738(csa_tree_add_6_33_groupi_n_491 ,csa_tree_add_6_33_groupi_n_489);
  not csa_tree_add_6_33_groupi_drc_bufs18739(csa_tree_add_6_33_groupi_n_490 ,csa_tree_add_6_33_groupi_n_489);
  not csa_tree_add_6_33_groupi_drc_bufs18740(csa_tree_add_6_33_groupi_n_489 ,csa_tree_add_6_33_groupi_n_929);
  not csa_tree_add_6_33_groupi_drc_bufs18742(csa_tree_add_6_33_groupi_n_488 ,csa_tree_add_6_33_groupi_n_486);
  not csa_tree_add_6_33_groupi_drc_bufs18743(csa_tree_add_6_33_groupi_n_487 ,csa_tree_add_6_33_groupi_n_486);
  not csa_tree_add_6_33_groupi_drc_bufs18744(csa_tree_add_6_33_groupi_n_486 ,csa_tree_add_6_33_groupi_n_929);
  not csa_tree_add_6_33_groupi_drc_bufs18746(csa_tree_add_6_33_groupi_n_485 ,csa_tree_add_6_33_groupi_n_483);
  not csa_tree_add_6_33_groupi_drc_bufs18747(csa_tree_add_6_33_groupi_n_484 ,csa_tree_add_6_33_groupi_n_483);
  not csa_tree_add_6_33_groupi_drc_bufs18748(csa_tree_add_6_33_groupi_n_483 ,csa_tree_add_6_33_groupi_n_967);
  not csa_tree_add_6_33_groupi_drc_bufs18750(csa_tree_add_6_33_groupi_n_482 ,csa_tree_add_6_33_groupi_n_480);
  not csa_tree_add_6_33_groupi_drc_bufs18751(csa_tree_add_6_33_groupi_n_481 ,csa_tree_add_6_33_groupi_n_480);
  not csa_tree_add_6_33_groupi_drc_bufs18752(csa_tree_add_6_33_groupi_n_480 ,csa_tree_add_6_33_groupi_n_967);
  not csa_tree_add_6_33_groupi_drc_bufs18754(csa_tree_add_6_33_groupi_n_479 ,csa_tree_add_6_33_groupi_n_477);
  not csa_tree_add_6_33_groupi_drc_bufs18755(csa_tree_add_6_33_groupi_n_478 ,csa_tree_add_6_33_groupi_n_477);
  not csa_tree_add_6_33_groupi_drc_bufs18756(csa_tree_add_6_33_groupi_n_477 ,csa_tree_add_6_33_groupi_n_986);
  not csa_tree_add_6_33_groupi_drc_bufs18758(csa_tree_add_6_33_groupi_n_476 ,csa_tree_add_6_33_groupi_n_474);
  not csa_tree_add_6_33_groupi_drc_bufs18759(csa_tree_add_6_33_groupi_n_475 ,csa_tree_add_6_33_groupi_n_474);
  not csa_tree_add_6_33_groupi_drc_bufs18760(csa_tree_add_6_33_groupi_n_474 ,csa_tree_add_6_33_groupi_n_986);
  not csa_tree_add_6_33_groupi_drc_bufs18762(csa_tree_add_6_33_groupi_n_473 ,csa_tree_add_6_33_groupi_n_471);
  not csa_tree_add_6_33_groupi_drc_bufs18763(csa_tree_add_6_33_groupi_n_472 ,csa_tree_add_6_33_groupi_n_471);
  not csa_tree_add_6_33_groupi_drc_bufs18764(csa_tree_add_6_33_groupi_n_471 ,csa_tree_add_6_33_groupi_n_968);
  not csa_tree_add_6_33_groupi_drc_bufs18766(csa_tree_add_6_33_groupi_n_470 ,csa_tree_add_6_33_groupi_n_468);
  not csa_tree_add_6_33_groupi_drc_bufs18767(csa_tree_add_6_33_groupi_n_469 ,csa_tree_add_6_33_groupi_n_468);
  not csa_tree_add_6_33_groupi_drc_bufs18768(csa_tree_add_6_33_groupi_n_468 ,csa_tree_add_6_33_groupi_n_932);
  not csa_tree_add_6_33_groupi_drc_bufs18770(csa_tree_add_6_33_groupi_n_467 ,csa_tree_add_6_33_groupi_n_465);
  not csa_tree_add_6_33_groupi_drc_bufs18771(csa_tree_add_6_33_groupi_n_466 ,csa_tree_add_6_33_groupi_n_465);
  not csa_tree_add_6_33_groupi_drc_bufs18772(csa_tree_add_6_33_groupi_n_465 ,csa_tree_add_6_33_groupi_n_931);
  not csa_tree_add_6_33_groupi_drc_bufs18774(csa_tree_add_6_33_groupi_n_464 ,csa_tree_add_6_33_groupi_n_462);
  not csa_tree_add_6_33_groupi_drc_bufs18775(csa_tree_add_6_33_groupi_n_463 ,csa_tree_add_6_33_groupi_n_462);
  not csa_tree_add_6_33_groupi_drc_bufs18776(csa_tree_add_6_33_groupi_n_462 ,csa_tree_add_6_33_groupi_n_905);
  not csa_tree_add_6_33_groupi_drc_bufs18778(csa_tree_add_6_33_groupi_n_461 ,csa_tree_add_6_33_groupi_n_459);
  not csa_tree_add_6_33_groupi_drc_bufs18779(csa_tree_add_6_33_groupi_n_460 ,csa_tree_add_6_33_groupi_n_459);
  not csa_tree_add_6_33_groupi_drc_bufs18780(csa_tree_add_6_33_groupi_n_459 ,csa_tree_add_6_33_groupi_n_931);
  not csa_tree_add_6_33_groupi_drc_bufs18782(csa_tree_add_6_33_groupi_n_458 ,csa_tree_add_6_33_groupi_n_456);
  not csa_tree_add_6_33_groupi_drc_bufs18783(csa_tree_add_6_33_groupi_n_457 ,csa_tree_add_6_33_groupi_n_456);
  not csa_tree_add_6_33_groupi_drc_bufs18784(csa_tree_add_6_33_groupi_n_456 ,csa_tree_add_6_33_groupi_n_968);
  not csa_tree_add_6_33_groupi_drc_bufs18786(csa_tree_add_6_33_groupi_n_455 ,csa_tree_add_6_33_groupi_n_453);
  not csa_tree_add_6_33_groupi_drc_bufs18787(csa_tree_add_6_33_groupi_n_454 ,csa_tree_add_6_33_groupi_n_453);
  not csa_tree_add_6_33_groupi_drc_bufs18788(csa_tree_add_6_33_groupi_n_453 ,csa_tree_add_6_33_groupi_n_906);
  not csa_tree_add_6_33_groupi_drc_bufs18790(csa_tree_add_6_33_groupi_n_452 ,csa_tree_add_6_33_groupi_n_450);
  not csa_tree_add_6_33_groupi_drc_bufs18791(csa_tree_add_6_33_groupi_n_451 ,csa_tree_add_6_33_groupi_n_450);
  not csa_tree_add_6_33_groupi_drc_bufs18792(csa_tree_add_6_33_groupi_n_450 ,csa_tree_add_6_33_groupi_n_1001);
  not csa_tree_add_6_33_groupi_drc_bufs18794(csa_tree_add_6_33_groupi_n_449 ,csa_tree_add_6_33_groupi_n_447);
  not csa_tree_add_6_33_groupi_drc_bufs18795(csa_tree_add_6_33_groupi_n_448 ,csa_tree_add_6_33_groupi_n_447);
  not csa_tree_add_6_33_groupi_drc_bufs18796(csa_tree_add_6_33_groupi_n_447 ,csa_tree_add_6_33_groupi_n_980);
  not csa_tree_add_6_33_groupi_drc_bufs18798(csa_tree_add_6_33_groupi_n_446 ,csa_tree_add_6_33_groupi_n_444);
  not csa_tree_add_6_33_groupi_drc_bufs18799(csa_tree_add_6_33_groupi_n_445 ,csa_tree_add_6_33_groupi_n_444);
  not csa_tree_add_6_33_groupi_drc_bufs18800(csa_tree_add_6_33_groupi_n_444 ,csa_tree_add_6_33_groupi_n_905);
  not csa_tree_add_6_33_groupi_drc_bufs18802(csa_tree_add_6_33_groupi_n_443 ,csa_tree_add_6_33_groupi_n_441);
  not csa_tree_add_6_33_groupi_drc_bufs18803(csa_tree_add_6_33_groupi_n_442 ,csa_tree_add_6_33_groupi_n_441);
  not csa_tree_add_6_33_groupi_drc_bufs18804(csa_tree_add_6_33_groupi_n_441 ,csa_tree_add_6_33_groupi_n_991);
  not csa_tree_add_6_33_groupi_drc_bufs18806(csa_tree_add_6_33_groupi_n_440 ,csa_tree_add_6_33_groupi_n_438);
  not csa_tree_add_6_33_groupi_drc_bufs18807(csa_tree_add_6_33_groupi_n_439 ,csa_tree_add_6_33_groupi_n_438);
  not csa_tree_add_6_33_groupi_drc_bufs18808(csa_tree_add_6_33_groupi_n_438 ,csa_tree_add_6_33_groupi_n_954);
  not csa_tree_add_6_33_groupi_drc_bufs18810(csa_tree_add_6_33_groupi_n_437 ,csa_tree_add_6_33_groupi_n_435);
  not csa_tree_add_6_33_groupi_drc_bufs18811(csa_tree_add_6_33_groupi_n_436 ,csa_tree_add_6_33_groupi_n_435);
  not csa_tree_add_6_33_groupi_drc_bufs18812(csa_tree_add_6_33_groupi_n_435 ,csa_tree_add_6_33_groupi_n_991);
  not csa_tree_add_6_33_groupi_drc_bufs18814(csa_tree_add_6_33_groupi_n_434 ,csa_tree_add_6_33_groupi_n_432);
  not csa_tree_add_6_33_groupi_drc_bufs18815(csa_tree_add_6_33_groupi_n_433 ,csa_tree_add_6_33_groupi_n_432);
  not csa_tree_add_6_33_groupi_drc_bufs18816(csa_tree_add_6_33_groupi_n_432 ,csa_tree_add_6_33_groupi_n_948);
  not csa_tree_add_6_33_groupi_drc_bufs18818(csa_tree_add_6_33_groupi_n_431 ,csa_tree_add_6_33_groupi_n_429);
  not csa_tree_add_6_33_groupi_drc_bufs18819(csa_tree_add_6_33_groupi_n_430 ,csa_tree_add_6_33_groupi_n_429);
  not csa_tree_add_6_33_groupi_drc_bufs18820(csa_tree_add_6_33_groupi_n_429 ,csa_tree_add_6_33_groupi_n_997);
  not csa_tree_add_6_33_groupi_drc_bufs18822(csa_tree_add_6_33_groupi_n_428 ,csa_tree_add_6_33_groupi_n_426);
  not csa_tree_add_6_33_groupi_drc_bufs18823(csa_tree_add_6_33_groupi_n_427 ,csa_tree_add_6_33_groupi_n_426);
  not csa_tree_add_6_33_groupi_drc_bufs18824(csa_tree_add_6_33_groupi_n_426 ,csa_tree_add_6_33_groupi_n_954);
  not csa_tree_add_6_33_groupi_drc_bufs18826(csa_tree_add_6_33_groupi_n_425 ,csa_tree_add_6_33_groupi_n_423);
  not csa_tree_add_6_33_groupi_drc_bufs18827(csa_tree_add_6_33_groupi_n_424 ,csa_tree_add_6_33_groupi_n_423);
  not csa_tree_add_6_33_groupi_drc_bufs18828(csa_tree_add_6_33_groupi_n_423 ,csa_tree_add_6_33_groupi_n_948);
  not csa_tree_add_6_33_groupi_drc_bufs18830(csa_tree_add_6_33_groupi_n_422 ,csa_tree_add_6_33_groupi_n_420);
  not csa_tree_add_6_33_groupi_drc_bufs18831(csa_tree_add_6_33_groupi_n_421 ,csa_tree_add_6_33_groupi_n_420);
  not csa_tree_add_6_33_groupi_drc_bufs18832(csa_tree_add_6_33_groupi_n_420 ,csa_tree_add_6_33_groupi_n_927);
  not csa_tree_add_6_33_groupi_drc_bufs18834(csa_tree_add_6_33_groupi_n_419 ,csa_tree_add_6_33_groupi_n_417);
  not csa_tree_add_6_33_groupi_drc_bufs18835(csa_tree_add_6_33_groupi_n_418 ,csa_tree_add_6_33_groupi_n_417);
  not csa_tree_add_6_33_groupi_drc_bufs18836(csa_tree_add_6_33_groupi_n_417 ,csa_tree_add_6_33_groupi_n_936);
  not csa_tree_add_6_33_groupi_drc_bufs18838(csa_tree_add_6_33_groupi_n_416 ,csa_tree_add_6_33_groupi_n_414);
  not csa_tree_add_6_33_groupi_drc_bufs18839(csa_tree_add_6_33_groupi_n_415 ,csa_tree_add_6_33_groupi_n_414);
  not csa_tree_add_6_33_groupi_drc_bufs18840(csa_tree_add_6_33_groupi_n_414 ,csa_tree_add_6_33_groupi_n_936);
  not csa_tree_add_6_33_groupi_drc_bufs18842(csa_tree_add_6_33_groupi_n_413 ,csa_tree_add_6_33_groupi_n_411);
  not csa_tree_add_6_33_groupi_drc_bufs18843(csa_tree_add_6_33_groupi_n_412 ,csa_tree_add_6_33_groupi_n_411);
  not csa_tree_add_6_33_groupi_drc_bufs18844(csa_tree_add_6_33_groupi_n_411 ,csa_tree_add_6_33_groupi_n_937);
  not csa_tree_add_6_33_groupi_drc_bufs18846(csa_tree_add_6_33_groupi_n_410 ,csa_tree_add_6_33_groupi_n_408);
  not csa_tree_add_6_33_groupi_drc_bufs18847(csa_tree_add_6_33_groupi_n_409 ,csa_tree_add_6_33_groupi_n_408);
  not csa_tree_add_6_33_groupi_drc_bufs18848(csa_tree_add_6_33_groupi_n_408 ,csa_tree_add_6_33_groupi_n_937);
  not csa_tree_add_6_33_groupi_drc_bufs18850(csa_tree_add_6_33_groupi_n_407 ,csa_tree_add_6_33_groupi_n_405);
  not csa_tree_add_6_33_groupi_drc_bufs18851(csa_tree_add_6_33_groupi_n_406 ,csa_tree_add_6_33_groupi_n_405);
  not csa_tree_add_6_33_groupi_drc_bufs18852(csa_tree_add_6_33_groupi_n_405 ,csa_tree_add_6_33_groupi_n_971);
  not csa_tree_add_6_33_groupi_drc_bufs18854(csa_tree_add_6_33_groupi_n_404 ,csa_tree_add_6_33_groupi_n_402);
  not csa_tree_add_6_33_groupi_drc_bufs18855(csa_tree_add_6_33_groupi_n_403 ,csa_tree_add_6_33_groupi_n_402);
  not csa_tree_add_6_33_groupi_drc_bufs18856(csa_tree_add_6_33_groupi_n_402 ,csa_tree_add_6_33_groupi_n_971);
  not csa_tree_add_6_33_groupi_drc_bufs18858(csa_tree_add_6_33_groupi_n_401 ,csa_tree_add_6_33_groupi_n_399);
  not csa_tree_add_6_33_groupi_drc_bufs18859(csa_tree_add_6_33_groupi_n_400 ,csa_tree_add_6_33_groupi_n_399);
  not csa_tree_add_6_33_groupi_drc_bufs18860(csa_tree_add_6_33_groupi_n_399 ,csa_tree_add_6_33_groupi_n_926);
  not csa_tree_add_6_33_groupi_drc_bufs18862(csa_tree_add_6_33_groupi_n_398 ,csa_tree_add_6_33_groupi_n_396);
  not csa_tree_add_6_33_groupi_drc_bufs18863(csa_tree_add_6_33_groupi_n_397 ,csa_tree_add_6_33_groupi_n_396);
  not csa_tree_add_6_33_groupi_drc_bufs18864(csa_tree_add_6_33_groupi_n_396 ,csa_tree_add_6_33_groupi_n_938);
  not csa_tree_add_6_33_groupi_drc_bufs18866(csa_tree_add_6_33_groupi_n_395 ,csa_tree_add_6_33_groupi_n_393);
  not csa_tree_add_6_33_groupi_drc_bufs18867(csa_tree_add_6_33_groupi_n_394 ,csa_tree_add_6_33_groupi_n_393);
  not csa_tree_add_6_33_groupi_drc_bufs18868(csa_tree_add_6_33_groupi_n_393 ,csa_tree_add_6_33_groupi_n_923);
  not csa_tree_add_6_33_groupi_drc_bufs18870(csa_tree_add_6_33_groupi_n_392 ,csa_tree_add_6_33_groupi_n_390);
  not csa_tree_add_6_33_groupi_drc_bufs18871(csa_tree_add_6_33_groupi_n_391 ,csa_tree_add_6_33_groupi_n_390);
  not csa_tree_add_6_33_groupi_drc_bufs18872(csa_tree_add_6_33_groupi_n_390 ,csa_tree_add_6_33_groupi_n_923);
  not csa_tree_add_6_33_groupi_drc_bufs18874(csa_tree_add_6_33_groupi_n_389 ,csa_tree_add_6_33_groupi_n_387);
  not csa_tree_add_6_33_groupi_drc_bufs18875(csa_tree_add_6_33_groupi_n_388 ,csa_tree_add_6_33_groupi_n_387);
  not csa_tree_add_6_33_groupi_drc_bufs18876(csa_tree_add_6_33_groupi_n_387 ,csa_tree_add_6_33_groupi_n_972);
  not csa_tree_add_6_33_groupi_drc_bufs18878(csa_tree_add_6_33_groupi_n_386 ,csa_tree_add_6_33_groupi_n_384);
  not csa_tree_add_6_33_groupi_drc_bufs18879(csa_tree_add_6_33_groupi_n_385 ,csa_tree_add_6_33_groupi_n_384);
  not csa_tree_add_6_33_groupi_drc_bufs18880(csa_tree_add_6_33_groupi_n_384 ,csa_tree_add_6_33_groupi_n_972);
  not csa_tree_add_6_33_groupi_drc_bufs18882(csa_tree_add_6_33_groupi_n_383 ,csa_tree_add_6_33_groupi_n_381);
  not csa_tree_add_6_33_groupi_drc_bufs18883(csa_tree_add_6_33_groupi_n_382 ,csa_tree_add_6_33_groupi_n_381);
  not csa_tree_add_6_33_groupi_drc_bufs18884(csa_tree_add_6_33_groupi_n_381 ,csa_tree_add_6_33_groupi_n_939);
  not csa_tree_add_6_33_groupi_drc_bufs18886(csa_tree_add_6_33_groupi_n_380 ,csa_tree_add_6_33_groupi_n_378);
  not csa_tree_add_6_33_groupi_drc_bufs18887(csa_tree_add_6_33_groupi_n_379 ,csa_tree_add_6_33_groupi_n_378);
  not csa_tree_add_6_33_groupi_drc_bufs18888(csa_tree_add_6_33_groupi_n_378 ,csa_tree_add_6_33_groupi_n_939);
  not csa_tree_add_6_33_groupi_drc_bufs18890(csa_tree_add_6_33_groupi_n_377 ,csa_tree_add_6_33_groupi_n_375);
  not csa_tree_add_6_33_groupi_drc_bufs18891(csa_tree_add_6_33_groupi_n_376 ,csa_tree_add_6_33_groupi_n_375);
  not csa_tree_add_6_33_groupi_drc_bufs18892(csa_tree_add_6_33_groupi_n_375 ,csa_tree_add_6_33_groupi_n_886);
  not csa_tree_add_6_33_groupi_drc_bufs18894(csa_tree_add_6_33_groupi_n_374 ,csa_tree_add_6_33_groupi_n_372);
  not csa_tree_add_6_33_groupi_drc_bufs18895(csa_tree_add_6_33_groupi_n_373 ,csa_tree_add_6_33_groupi_n_372);
  not csa_tree_add_6_33_groupi_drc_bufs18896(csa_tree_add_6_33_groupi_n_372 ,csa_tree_add_6_33_groupi_n_921);
  not csa_tree_add_6_33_groupi_drc_bufs18898(csa_tree_add_6_33_groupi_n_371 ,csa_tree_add_6_33_groupi_n_369);
  not csa_tree_add_6_33_groupi_drc_bufs18899(csa_tree_add_6_33_groupi_n_370 ,csa_tree_add_6_33_groupi_n_369);
  not csa_tree_add_6_33_groupi_drc_bufs18900(csa_tree_add_6_33_groupi_n_369 ,csa_tree_add_6_33_groupi_n_920);
  not csa_tree_add_6_33_groupi_drc_bufs18902(csa_tree_add_6_33_groupi_n_368 ,csa_tree_add_6_33_groupi_n_366);
  not csa_tree_add_6_33_groupi_drc_bufs18903(csa_tree_add_6_33_groupi_n_367 ,csa_tree_add_6_33_groupi_n_366);
  not csa_tree_add_6_33_groupi_drc_bufs18904(csa_tree_add_6_33_groupi_n_366 ,csa_tree_add_6_33_groupi_n_920);
  not csa_tree_add_6_33_groupi_drc_bufs18906(csa_tree_add_6_33_groupi_n_365 ,csa_tree_add_6_33_groupi_n_363);
  not csa_tree_add_6_33_groupi_drc_bufs18907(csa_tree_add_6_33_groupi_n_364 ,csa_tree_add_6_33_groupi_n_363);
  not csa_tree_add_6_33_groupi_drc_bufs18908(csa_tree_add_6_33_groupi_n_363 ,csa_tree_add_6_33_groupi_n_919);
  not csa_tree_add_6_33_groupi_drc_bufs18910(csa_tree_add_6_33_groupi_n_362 ,csa_tree_add_6_33_groupi_n_360);
  not csa_tree_add_6_33_groupi_drc_bufs18911(csa_tree_add_6_33_groupi_n_361 ,csa_tree_add_6_33_groupi_n_360);
  not csa_tree_add_6_33_groupi_drc_bufs18912(csa_tree_add_6_33_groupi_n_360 ,csa_tree_add_6_33_groupi_n_919);
  not csa_tree_add_6_33_groupi_drc_bufs18914(csa_tree_add_6_33_groupi_n_359 ,csa_tree_add_6_33_groupi_n_357);
  not csa_tree_add_6_33_groupi_drc_bufs18915(csa_tree_add_6_33_groupi_n_358 ,csa_tree_add_6_33_groupi_n_357);
  not csa_tree_add_6_33_groupi_drc_bufs18916(csa_tree_add_6_33_groupi_n_357 ,csa_tree_add_6_33_groupi_n_940);
  not csa_tree_add_6_33_groupi_drc_bufs18918(csa_tree_add_6_33_groupi_n_356 ,csa_tree_add_6_33_groupi_n_354);
  not csa_tree_add_6_33_groupi_drc_bufs18919(csa_tree_add_6_33_groupi_n_355 ,csa_tree_add_6_33_groupi_n_354);
  not csa_tree_add_6_33_groupi_drc_bufs18920(csa_tree_add_6_33_groupi_n_354 ,csa_tree_add_6_33_groupi_n_940);
  not csa_tree_add_6_33_groupi_drc_bufs18922(csa_tree_add_6_33_groupi_n_353 ,csa_tree_add_6_33_groupi_n_351);
  not csa_tree_add_6_33_groupi_drc_bufs18923(csa_tree_add_6_33_groupi_n_352 ,csa_tree_add_6_33_groupi_n_351);
  not csa_tree_add_6_33_groupi_drc_bufs18924(csa_tree_add_6_33_groupi_n_351 ,csa_tree_add_6_33_groupi_n_903);
  not csa_tree_add_6_33_groupi_drc_bufs18926(csa_tree_add_6_33_groupi_n_350 ,csa_tree_add_6_33_groupi_n_348);
  not csa_tree_add_6_33_groupi_drc_bufs18927(csa_tree_add_6_33_groupi_n_349 ,csa_tree_add_6_33_groupi_n_348);
  not csa_tree_add_6_33_groupi_drc_bufs18928(csa_tree_add_6_33_groupi_n_348 ,csa_tree_add_6_33_groupi_n_941);
  not csa_tree_add_6_33_groupi_drc_bufs18930(csa_tree_add_6_33_groupi_n_347 ,csa_tree_add_6_33_groupi_n_345);
  not csa_tree_add_6_33_groupi_drc_bufs18931(csa_tree_add_6_33_groupi_n_346 ,csa_tree_add_6_33_groupi_n_345);
  not csa_tree_add_6_33_groupi_drc_bufs18932(csa_tree_add_6_33_groupi_n_345 ,csa_tree_add_6_33_groupi_n_942);
  not csa_tree_add_6_33_groupi_drc_bufs18934(csa_tree_add_6_33_groupi_n_344 ,csa_tree_add_6_33_groupi_n_342);
  not csa_tree_add_6_33_groupi_drc_bufs18935(csa_tree_add_6_33_groupi_n_343 ,csa_tree_add_6_33_groupi_n_342);
  not csa_tree_add_6_33_groupi_drc_bufs18936(csa_tree_add_6_33_groupi_n_342 ,csa_tree_add_6_33_groupi_n_942);
  not csa_tree_add_6_33_groupi_drc_bufs18938(csa_tree_add_6_33_groupi_n_341 ,csa_tree_add_6_33_groupi_n_339);
  not csa_tree_add_6_33_groupi_drc_bufs18939(csa_tree_add_6_33_groupi_n_340 ,csa_tree_add_6_33_groupi_n_339);
  not csa_tree_add_6_33_groupi_drc_bufs18940(csa_tree_add_6_33_groupi_n_339 ,csa_tree_add_6_33_groupi_n_943);
  not csa_tree_add_6_33_groupi_drc_bufs18942(csa_tree_add_6_33_groupi_n_338 ,csa_tree_add_6_33_groupi_n_336);
  not csa_tree_add_6_33_groupi_drc_bufs18943(csa_tree_add_6_33_groupi_n_337 ,csa_tree_add_6_33_groupi_n_336);
  not csa_tree_add_6_33_groupi_drc_bufs18944(csa_tree_add_6_33_groupi_n_336 ,csa_tree_add_6_33_groupi_n_943);
  not csa_tree_add_6_33_groupi_drc_bufs18946(csa_tree_add_6_33_groupi_n_335 ,csa_tree_add_6_33_groupi_n_333);
  not csa_tree_add_6_33_groupi_drc_bufs18947(csa_tree_add_6_33_groupi_n_334 ,csa_tree_add_6_33_groupi_n_333);
  not csa_tree_add_6_33_groupi_drc_bufs18948(csa_tree_add_6_33_groupi_n_333 ,csa_tree_add_6_33_groupi_n_974);
  not csa_tree_add_6_33_groupi_drc_bufs18950(csa_tree_add_6_33_groupi_n_332 ,csa_tree_add_6_33_groupi_n_330);
  not csa_tree_add_6_33_groupi_drc_bufs18951(csa_tree_add_6_33_groupi_n_331 ,csa_tree_add_6_33_groupi_n_330);
  not csa_tree_add_6_33_groupi_drc_bufs18952(csa_tree_add_6_33_groupi_n_330 ,csa_tree_add_6_33_groupi_n_974);
  not csa_tree_add_6_33_groupi_drc_bufs18954(csa_tree_add_6_33_groupi_n_329 ,csa_tree_add_6_33_groupi_n_327);
  not csa_tree_add_6_33_groupi_drc_bufs18955(csa_tree_add_6_33_groupi_n_328 ,csa_tree_add_6_33_groupi_n_327);
  not csa_tree_add_6_33_groupi_drc_bufs18956(csa_tree_add_6_33_groupi_n_327 ,csa_tree_add_6_33_groupi_n_944);
  not csa_tree_add_6_33_groupi_drc_bufs18958(csa_tree_add_6_33_groupi_n_326 ,csa_tree_add_6_33_groupi_n_324);
  not csa_tree_add_6_33_groupi_drc_bufs18959(csa_tree_add_6_33_groupi_n_325 ,csa_tree_add_6_33_groupi_n_324);
  not csa_tree_add_6_33_groupi_drc_bufs18960(csa_tree_add_6_33_groupi_n_324 ,csa_tree_add_6_33_groupi_n_944);
  not csa_tree_add_6_33_groupi_drc_bufs18962(csa_tree_add_6_33_groupi_n_323 ,csa_tree_add_6_33_groupi_n_321);
  not csa_tree_add_6_33_groupi_drc_bufs18963(csa_tree_add_6_33_groupi_n_322 ,csa_tree_add_6_33_groupi_n_321);
  not csa_tree_add_6_33_groupi_drc_bufs18964(csa_tree_add_6_33_groupi_n_321 ,csa_tree_add_6_33_groupi_n_945);
  not csa_tree_add_6_33_groupi_drc_bufs18966(csa_tree_add_6_33_groupi_n_320 ,csa_tree_add_6_33_groupi_n_318);
  not csa_tree_add_6_33_groupi_drc_bufs18967(csa_tree_add_6_33_groupi_n_319 ,csa_tree_add_6_33_groupi_n_318);
  not csa_tree_add_6_33_groupi_drc_bufs18968(csa_tree_add_6_33_groupi_n_318 ,csa_tree_add_6_33_groupi_n_945);
  not csa_tree_add_6_33_groupi_drc_bufs18970(csa_tree_add_6_33_groupi_n_317 ,csa_tree_add_6_33_groupi_n_315);
  not csa_tree_add_6_33_groupi_drc_bufs18971(csa_tree_add_6_33_groupi_n_316 ,csa_tree_add_6_33_groupi_n_315);
  not csa_tree_add_6_33_groupi_drc_bufs18972(csa_tree_add_6_33_groupi_n_315 ,csa_tree_add_6_33_groupi_n_975);
  not csa_tree_add_6_33_groupi_drc_bufs18974(csa_tree_add_6_33_groupi_n_314 ,csa_tree_add_6_33_groupi_n_312);
  not csa_tree_add_6_33_groupi_drc_bufs18975(csa_tree_add_6_33_groupi_n_313 ,csa_tree_add_6_33_groupi_n_312);
  not csa_tree_add_6_33_groupi_drc_bufs18976(csa_tree_add_6_33_groupi_n_312 ,csa_tree_add_6_33_groupi_n_975);
  not csa_tree_add_6_33_groupi_drc_bufs18978(csa_tree_add_6_33_groupi_n_311 ,csa_tree_add_6_33_groupi_n_309);
  not csa_tree_add_6_33_groupi_drc_bufs18979(csa_tree_add_6_33_groupi_n_310 ,csa_tree_add_6_33_groupi_n_309);
  not csa_tree_add_6_33_groupi_drc_bufs18980(csa_tree_add_6_33_groupi_n_309 ,csa_tree_add_6_33_groupi_n_912);
  not csa_tree_add_6_33_groupi_drc_bufs18982(csa_tree_add_6_33_groupi_n_308 ,csa_tree_add_6_33_groupi_n_306);
  not csa_tree_add_6_33_groupi_drc_bufs18983(csa_tree_add_6_33_groupi_n_307 ,csa_tree_add_6_33_groupi_n_306);
  not csa_tree_add_6_33_groupi_drc_bufs18984(csa_tree_add_6_33_groupi_n_306 ,csa_tree_add_6_33_groupi_n_912);
  not csa_tree_add_6_33_groupi_drc_bufs18986(csa_tree_add_6_33_groupi_n_305 ,csa_tree_add_6_33_groupi_n_303);
  not csa_tree_add_6_33_groupi_drc_bufs18987(csa_tree_add_6_33_groupi_n_304 ,csa_tree_add_6_33_groupi_n_303);
  not csa_tree_add_6_33_groupi_drc_bufs18988(csa_tree_add_6_33_groupi_n_303 ,csa_tree_add_6_33_groupi_n_994);
  not csa_tree_add_6_33_groupi_drc_bufs18990(csa_tree_add_6_33_groupi_n_302 ,csa_tree_add_6_33_groupi_n_300);
  not csa_tree_add_6_33_groupi_drc_bufs18991(csa_tree_add_6_33_groupi_n_301 ,csa_tree_add_6_33_groupi_n_300);
  not csa_tree_add_6_33_groupi_drc_bufs18992(csa_tree_add_6_33_groupi_n_300 ,csa_tree_add_6_33_groupi_n_911);
  not csa_tree_add_6_33_groupi_drc_bufs18994(csa_tree_add_6_33_groupi_n_299 ,csa_tree_add_6_33_groupi_n_297);
  not csa_tree_add_6_33_groupi_drc_bufs18995(csa_tree_add_6_33_groupi_n_298 ,csa_tree_add_6_33_groupi_n_297);
  not csa_tree_add_6_33_groupi_drc_bufs18996(csa_tree_add_6_33_groupi_n_297 ,csa_tree_add_6_33_groupi_n_990);
  not csa_tree_add_6_33_groupi_drc_bufs18998(csa_tree_add_6_33_groupi_n_296 ,csa_tree_add_6_33_groupi_n_294);
  not csa_tree_add_6_33_groupi_drc_bufs18999(csa_tree_add_6_33_groupi_n_295 ,csa_tree_add_6_33_groupi_n_294);
  not csa_tree_add_6_33_groupi_drc_bufs19000(csa_tree_add_6_33_groupi_n_294 ,csa_tree_add_6_33_groupi_n_990);
  not csa_tree_add_6_33_groupi_drc_bufs19002(csa_tree_add_6_33_groupi_n_293 ,csa_tree_add_6_33_groupi_n_291);
  not csa_tree_add_6_33_groupi_drc_bufs19003(csa_tree_add_6_33_groupi_n_292 ,csa_tree_add_6_33_groupi_n_291);
  not csa_tree_add_6_33_groupi_drc_bufs19004(csa_tree_add_6_33_groupi_n_291 ,csa_tree_add_6_33_groupi_n_885);
  not csa_tree_add_6_33_groupi_drc_bufs19006(csa_tree_add_6_33_groupi_n_290 ,csa_tree_add_6_33_groupi_n_288);
  not csa_tree_add_6_33_groupi_drc_bufs19007(csa_tree_add_6_33_groupi_n_289 ,csa_tree_add_6_33_groupi_n_288);
  not csa_tree_add_6_33_groupi_drc_bufs19008(csa_tree_add_6_33_groupi_n_288 ,csa_tree_add_6_33_groupi_n_885);
  not csa_tree_add_6_33_groupi_drc_bufs19010(csa_tree_add_6_33_groupi_n_287 ,csa_tree_add_6_33_groupi_n_285);
  not csa_tree_add_6_33_groupi_drc_bufs19011(csa_tree_add_6_33_groupi_n_286 ,csa_tree_add_6_33_groupi_n_285);
  not csa_tree_add_6_33_groupi_drc_bufs19012(csa_tree_add_6_33_groupi_n_285 ,csa_tree_add_6_33_groupi_n_946);
  not csa_tree_add_6_33_groupi_drc_bufs19014(csa_tree_add_6_33_groupi_n_284 ,csa_tree_add_6_33_groupi_n_282);
  not csa_tree_add_6_33_groupi_drc_bufs19015(csa_tree_add_6_33_groupi_n_283 ,csa_tree_add_6_33_groupi_n_282);
  not csa_tree_add_6_33_groupi_drc_bufs19016(csa_tree_add_6_33_groupi_n_282 ,csa_tree_add_6_33_groupi_n_946);
  not csa_tree_add_6_33_groupi_drc_bufs19018(csa_tree_add_6_33_groupi_n_281 ,csa_tree_add_6_33_groupi_n_279);
  not csa_tree_add_6_33_groupi_drc_bufs19019(csa_tree_add_6_33_groupi_n_280 ,csa_tree_add_6_33_groupi_n_279);
  not csa_tree_add_6_33_groupi_drc_bufs19020(csa_tree_add_6_33_groupi_n_279 ,csa_tree_add_6_33_groupi_n_976);
  not csa_tree_add_6_33_groupi_drc_bufs19022(csa_tree_add_6_33_groupi_n_278 ,csa_tree_add_6_33_groupi_n_276);
  not csa_tree_add_6_33_groupi_drc_bufs19023(csa_tree_add_6_33_groupi_n_277 ,csa_tree_add_6_33_groupi_n_276);
  not csa_tree_add_6_33_groupi_drc_bufs19024(csa_tree_add_6_33_groupi_n_276 ,csa_tree_add_6_33_groupi_n_947);
  not csa_tree_add_6_33_groupi_drc_bufs19026(csa_tree_add_6_33_groupi_n_275 ,csa_tree_add_6_33_groupi_n_273);
  not csa_tree_add_6_33_groupi_drc_bufs19027(csa_tree_add_6_33_groupi_n_274 ,csa_tree_add_6_33_groupi_n_273);
  not csa_tree_add_6_33_groupi_drc_bufs19028(csa_tree_add_6_33_groupi_n_273 ,csa_tree_add_6_33_groupi_n_901);
  not csa_tree_add_6_33_groupi_drc_bufs19030(csa_tree_add_6_33_groupi_n_272 ,csa_tree_add_6_33_groupi_n_270);
  not csa_tree_add_6_33_groupi_drc_bufs19031(csa_tree_add_6_33_groupi_n_271 ,csa_tree_add_6_33_groupi_n_270);
  not csa_tree_add_6_33_groupi_drc_bufs19032(csa_tree_add_6_33_groupi_n_270 ,csa_tree_add_6_33_groupi_n_947);
  not csa_tree_add_6_33_groupi_drc_bufs19034(csa_tree_add_6_33_groupi_n_269 ,csa_tree_add_6_33_groupi_n_267);
  not csa_tree_add_6_33_groupi_drc_bufs19035(csa_tree_add_6_33_groupi_n_268 ,csa_tree_add_6_33_groupi_n_267);
  not csa_tree_add_6_33_groupi_drc_bufs19036(csa_tree_add_6_33_groupi_n_267 ,csa_tree_add_6_33_groupi_n_976);
  not csa_tree_add_6_33_groupi_drc_bufs19038(csa_tree_add_6_33_groupi_n_266 ,csa_tree_add_6_33_groupi_n_264);
  not csa_tree_add_6_33_groupi_drc_bufs19039(csa_tree_add_6_33_groupi_n_265 ,csa_tree_add_6_33_groupi_n_264);
  not csa_tree_add_6_33_groupi_drc_bufs19040(csa_tree_add_6_33_groupi_n_264 ,csa_tree_add_6_33_groupi_n_899);
  not csa_tree_add_6_33_groupi_drc_bufs19042(csa_tree_add_6_33_groupi_n_263 ,csa_tree_add_6_33_groupi_n_261);
  not csa_tree_add_6_33_groupi_drc_bufs19043(csa_tree_add_6_33_groupi_n_262 ,csa_tree_add_6_33_groupi_n_261);
  not csa_tree_add_6_33_groupi_drc_bufs19044(csa_tree_add_6_33_groupi_n_261 ,csa_tree_add_6_33_groupi_n_891);
  not csa_tree_add_6_33_groupi_drc_bufs19046(csa_tree_add_6_33_groupi_n_260 ,csa_tree_add_6_33_groupi_n_258);
  not csa_tree_add_6_33_groupi_drc_bufs19047(csa_tree_add_6_33_groupi_n_259 ,csa_tree_add_6_33_groupi_n_258);
  not csa_tree_add_6_33_groupi_drc_bufs19048(csa_tree_add_6_33_groupi_n_258 ,csa_tree_add_6_33_groupi_n_985);
  not csa_tree_add_6_33_groupi_drc_bufs19050(csa_tree_add_6_33_groupi_n_257 ,csa_tree_add_6_33_groupi_n_255);
  not csa_tree_add_6_33_groupi_drc_bufs19051(csa_tree_add_6_33_groupi_n_256 ,csa_tree_add_6_33_groupi_n_255);
  not csa_tree_add_6_33_groupi_drc_bufs19052(csa_tree_add_6_33_groupi_n_255 ,csa_tree_add_6_33_groupi_n_901);
  not csa_tree_add_6_33_groupi_drc_bufs19054(csa_tree_add_6_33_groupi_n_254 ,csa_tree_add_6_33_groupi_n_252);
  not csa_tree_add_6_33_groupi_drc_bufs19055(csa_tree_add_6_33_groupi_n_253 ,csa_tree_add_6_33_groupi_n_252);
  not csa_tree_add_6_33_groupi_drc_bufs19056(csa_tree_add_6_33_groupi_n_252 ,csa_tree_add_6_33_groupi_n_999);
  not csa_tree_add_6_33_groupi_drc_bufs19058(csa_tree_add_6_33_groupi_n_251 ,csa_tree_add_6_33_groupi_n_249);
  not csa_tree_add_6_33_groupi_drc_bufs19059(csa_tree_add_6_33_groupi_n_250 ,csa_tree_add_6_33_groupi_n_249);
  not csa_tree_add_6_33_groupi_drc_bufs19060(csa_tree_add_6_33_groupi_n_249 ,csa_tree_add_6_33_groupi_n_977);
  not csa_tree_add_6_33_groupi_drc_bufs19062(csa_tree_add_6_33_groupi_n_248 ,csa_tree_add_6_33_groupi_n_246);
  not csa_tree_add_6_33_groupi_drc_bufs19063(csa_tree_add_6_33_groupi_n_247 ,csa_tree_add_6_33_groupi_n_246);
  not csa_tree_add_6_33_groupi_drc_bufs19064(csa_tree_add_6_33_groupi_n_246 ,csa_tree_add_6_33_groupi_n_999);
  not csa_tree_add_6_33_groupi_drc_bufs19066(csa_tree_add_6_33_groupi_n_245 ,csa_tree_add_6_33_groupi_n_243);
  not csa_tree_add_6_33_groupi_drc_bufs19067(csa_tree_add_6_33_groupi_n_244 ,csa_tree_add_6_33_groupi_n_243);
  not csa_tree_add_6_33_groupi_drc_bufs19068(csa_tree_add_6_33_groupi_n_243 ,csa_tree_add_6_33_groupi_n_979);
  not csa_tree_add_6_33_groupi_drc_bufs19070(csa_tree_add_6_33_groupi_n_242 ,csa_tree_add_6_33_groupi_n_240);
  not csa_tree_add_6_33_groupi_drc_bufs19071(csa_tree_add_6_33_groupi_n_241 ,csa_tree_add_6_33_groupi_n_240);
  not csa_tree_add_6_33_groupi_drc_bufs19072(csa_tree_add_6_33_groupi_n_240 ,csa_tree_add_6_33_groupi_n_965);
  not csa_tree_add_6_33_groupi_drc_bufs19074(csa_tree_add_6_33_groupi_n_239 ,csa_tree_add_6_33_groupi_n_237);
  not csa_tree_add_6_33_groupi_drc_bufs19075(csa_tree_add_6_33_groupi_n_238 ,csa_tree_add_6_33_groupi_n_237);
  not csa_tree_add_6_33_groupi_drc_bufs19076(csa_tree_add_6_33_groupi_n_237 ,csa_tree_add_6_33_groupi_n_979);
  not csa_tree_add_6_33_groupi_drc_bufs19078(csa_tree_add_6_33_groupi_n_236 ,csa_tree_add_6_33_groupi_n_234);
  not csa_tree_add_6_33_groupi_drc_bufs19079(csa_tree_add_6_33_groupi_n_235 ,csa_tree_add_6_33_groupi_n_234);
  not csa_tree_add_6_33_groupi_drc_bufs19080(csa_tree_add_6_33_groupi_n_234 ,csa_tree_add_6_33_groupi_n_911);
  not csa_tree_add_6_33_groupi_drc_bufs19082(csa_tree_add_6_33_groupi_n_233 ,csa_tree_add_6_33_groupi_n_231);
  not csa_tree_add_6_33_groupi_drc_bufs19083(csa_tree_add_6_33_groupi_n_232 ,csa_tree_add_6_33_groupi_n_231);
  not csa_tree_add_6_33_groupi_drc_bufs19084(csa_tree_add_6_33_groupi_n_231 ,csa_tree_add_6_33_groupi_n_900);
  not csa_tree_add_6_33_groupi_drc_bufs19086(csa_tree_add_6_33_groupi_n_230 ,csa_tree_add_6_33_groupi_n_228);
  not csa_tree_add_6_33_groupi_drc_bufs19087(csa_tree_add_6_33_groupi_n_229 ,csa_tree_add_6_33_groupi_n_228);
  not csa_tree_add_6_33_groupi_drc_bufs19088(csa_tree_add_6_33_groupi_n_228 ,csa_tree_add_6_33_groupi_n_893);
  not csa_tree_add_6_33_groupi_drc_bufs19090(csa_tree_add_6_33_groupi_n_227 ,csa_tree_add_6_33_groupi_n_225);
  not csa_tree_add_6_33_groupi_drc_bufs19091(csa_tree_add_6_33_groupi_n_226 ,csa_tree_add_6_33_groupi_n_225);
  not csa_tree_add_6_33_groupi_drc_bufs19092(csa_tree_add_6_33_groupi_n_225 ,csa_tree_add_6_33_groupi_n_949);
  not csa_tree_add_6_33_groupi_drc_bufs19094(csa_tree_add_6_33_groupi_n_224 ,csa_tree_add_6_33_groupi_n_222);
  not csa_tree_add_6_33_groupi_drc_bufs19095(csa_tree_add_6_33_groupi_n_223 ,csa_tree_add_6_33_groupi_n_222);
  not csa_tree_add_6_33_groupi_drc_bufs19096(csa_tree_add_6_33_groupi_n_222 ,csa_tree_add_6_33_groupi_n_949);
  not csa_tree_add_6_33_groupi_drc_bufs19098(csa_tree_add_6_33_groupi_n_221 ,csa_tree_add_6_33_groupi_n_219);
  not csa_tree_add_6_33_groupi_drc_bufs19099(csa_tree_add_6_33_groupi_n_220 ,csa_tree_add_6_33_groupi_n_219);
  not csa_tree_add_6_33_groupi_drc_bufs19100(csa_tree_add_6_33_groupi_n_219 ,csa_tree_add_6_33_groupi_n_938);
  not csa_tree_add_6_33_groupi_drc_bufs19102(csa_tree_add_6_33_groupi_n_218 ,csa_tree_add_6_33_groupi_n_216);
  not csa_tree_add_6_33_groupi_drc_bufs19103(csa_tree_add_6_33_groupi_n_217 ,csa_tree_add_6_33_groupi_n_216);
  not csa_tree_add_6_33_groupi_drc_bufs19104(csa_tree_add_6_33_groupi_n_216 ,csa_tree_add_6_33_groupi_n_950);
  not csa_tree_add_6_33_groupi_drc_bufs19106(csa_tree_add_6_33_groupi_n_215 ,csa_tree_add_6_33_groupi_n_213);
  not csa_tree_add_6_33_groupi_drc_bufs19107(csa_tree_add_6_33_groupi_n_214 ,csa_tree_add_6_33_groupi_n_213);
  not csa_tree_add_6_33_groupi_drc_bufs19108(csa_tree_add_6_33_groupi_n_213 ,csa_tree_add_6_33_groupi_n_896);
  not csa_tree_add_6_33_groupi_drc_bufs19110(csa_tree_add_6_33_groupi_n_212 ,csa_tree_add_6_33_groupi_n_210);
  not csa_tree_add_6_33_groupi_drc_bufs19111(csa_tree_add_6_33_groupi_n_211 ,csa_tree_add_6_33_groupi_n_210);
  not csa_tree_add_6_33_groupi_drc_bufs19112(csa_tree_add_6_33_groupi_n_210 ,csa_tree_add_6_33_groupi_n_896);
  not csa_tree_add_6_33_groupi_drc_bufs19114(csa_tree_add_6_33_groupi_n_209 ,csa_tree_add_6_33_groupi_n_207);
  not csa_tree_add_6_33_groupi_drc_bufs19115(csa_tree_add_6_33_groupi_n_208 ,csa_tree_add_6_33_groupi_n_207);
  not csa_tree_add_6_33_groupi_drc_bufs19116(csa_tree_add_6_33_groupi_n_207 ,csa_tree_add_6_33_groupi_n_921);
  not csa_tree_add_6_33_groupi_drc_bufs19118(csa_tree_add_6_33_groupi_n_206 ,csa_tree_add_6_33_groupi_n_204);
  not csa_tree_add_6_33_groupi_drc_bufs19119(csa_tree_add_6_33_groupi_n_205 ,csa_tree_add_6_33_groupi_n_204);
  not csa_tree_add_6_33_groupi_drc_bufs19120(csa_tree_add_6_33_groupi_n_204 ,csa_tree_add_6_33_groupi_n_897);
  not csa_tree_add_6_33_groupi_drc_bufs19122(csa_tree_add_6_33_groupi_n_203 ,csa_tree_add_6_33_groupi_n_201);
  not csa_tree_add_6_33_groupi_drc_bufs19123(csa_tree_add_6_33_groupi_n_202 ,csa_tree_add_6_33_groupi_n_201);
  not csa_tree_add_6_33_groupi_drc_bufs19124(csa_tree_add_6_33_groupi_n_201 ,csa_tree_add_6_33_groupi_n_951);
  not csa_tree_add_6_33_groupi_drc_bufs19126(csa_tree_add_6_33_groupi_n_200 ,csa_tree_add_6_33_groupi_n_198);
  not csa_tree_add_6_33_groupi_drc_bufs19127(csa_tree_add_6_33_groupi_n_199 ,csa_tree_add_6_33_groupi_n_198);
  not csa_tree_add_6_33_groupi_drc_bufs19128(csa_tree_add_6_33_groupi_n_198 ,csa_tree_add_6_33_groupi_n_951);
  not csa_tree_add_6_33_groupi_drc_bufs19130(csa_tree_add_6_33_groupi_n_197 ,csa_tree_add_6_33_groupi_n_195);
  not csa_tree_add_6_33_groupi_drc_bufs19131(csa_tree_add_6_33_groupi_n_196 ,csa_tree_add_6_33_groupi_n_195);
  not csa_tree_add_6_33_groupi_drc_bufs19132(csa_tree_add_6_33_groupi_n_195 ,csa_tree_add_6_33_groupi_n_941);
  not csa_tree_add_6_33_groupi_drc_bufs19134(csa_tree_add_6_33_groupi_n_194 ,csa_tree_add_6_33_groupi_n_192);
  not csa_tree_add_6_33_groupi_drc_bufs19135(csa_tree_add_6_33_groupi_n_193 ,csa_tree_add_6_33_groupi_n_192);
  not csa_tree_add_6_33_groupi_drc_bufs19136(csa_tree_add_6_33_groupi_n_192 ,csa_tree_add_6_33_groupi_n_978);
  not csa_tree_add_6_33_groupi_drc_bufs19138(csa_tree_add_6_33_groupi_n_191 ,csa_tree_add_6_33_groupi_n_189);
  not csa_tree_add_6_33_groupi_drc_bufs19139(csa_tree_add_6_33_groupi_n_190 ,csa_tree_add_6_33_groupi_n_189);
  not csa_tree_add_6_33_groupi_drc_bufs19140(csa_tree_add_6_33_groupi_n_189 ,csa_tree_add_6_33_groupi_n_992);
  not csa_tree_add_6_33_groupi_drc_bufs19142(csa_tree_add_6_33_groupi_n_188 ,csa_tree_add_6_33_groupi_n_186);
  not csa_tree_add_6_33_groupi_drc_bufs19143(csa_tree_add_6_33_groupi_n_187 ,csa_tree_add_6_33_groupi_n_186);
  not csa_tree_add_6_33_groupi_drc_bufs19144(csa_tree_add_6_33_groupi_n_186 ,csa_tree_add_6_33_groupi_n_992);
  not csa_tree_add_6_33_groupi_drc_bufs19146(csa_tree_add_6_33_groupi_n_185 ,csa_tree_add_6_33_groupi_n_183);
  not csa_tree_add_6_33_groupi_drc_bufs19147(csa_tree_add_6_33_groupi_n_184 ,csa_tree_add_6_33_groupi_n_183);
  not csa_tree_add_6_33_groupi_drc_bufs19148(csa_tree_add_6_33_groupi_n_183 ,csa_tree_add_6_33_groupi_n_952);
  not csa_tree_add_6_33_groupi_drc_bufs19150(csa_tree_add_6_33_groupi_n_182 ,csa_tree_add_6_33_groupi_n_180);
  not csa_tree_add_6_33_groupi_drc_bufs19151(csa_tree_add_6_33_groupi_n_181 ,csa_tree_add_6_33_groupi_n_180);
  not csa_tree_add_6_33_groupi_drc_bufs19152(csa_tree_add_6_33_groupi_n_180 ,csa_tree_add_6_33_groupi_n_1004);
  not csa_tree_add_6_33_groupi_drc_bufs19154(csa_tree_add_6_33_groupi_n_179 ,csa_tree_add_6_33_groupi_n_177);
  not csa_tree_add_6_33_groupi_drc_bufs19155(csa_tree_add_6_33_groupi_n_178 ,csa_tree_add_6_33_groupi_n_177);
  not csa_tree_add_6_33_groupi_drc_bufs19156(csa_tree_add_6_33_groupi_n_177 ,csa_tree_add_6_33_groupi_n_900);
  not csa_tree_add_6_33_groupi_drc_bufs19158(csa_tree_add_6_33_groupi_n_176 ,csa_tree_add_6_33_groupi_n_174);
  not csa_tree_add_6_33_groupi_drc_bufs19159(csa_tree_add_6_33_groupi_n_175 ,csa_tree_add_6_33_groupi_n_174);
  not csa_tree_add_6_33_groupi_drc_bufs19160(csa_tree_add_6_33_groupi_n_174 ,csa_tree_add_6_33_groupi_n_952);
  not csa_tree_add_6_33_groupi_drc_bufs19162(csa_tree_add_6_33_groupi_n_173 ,csa_tree_add_6_33_groupi_n_171);
  not csa_tree_add_6_33_groupi_drc_bufs19163(csa_tree_add_6_33_groupi_n_172 ,csa_tree_add_6_33_groupi_n_171);
  not csa_tree_add_6_33_groupi_drc_bufs19164(csa_tree_add_6_33_groupi_n_171 ,csa_tree_add_6_33_groupi_n_934);
  not csa_tree_add_6_33_groupi_drc_bufs19166(csa_tree_add_6_33_groupi_n_170 ,csa_tree_add_6_33_groupi_n_168);
  not csa_tree_add_6_33_groupi_drc_bufs19167(csa_tree_add_6_33_groupi_n_169 ,csa_tree_add_6_33_groupi_n_168);
  not csa_tree_add_6_33_groupi_drc_bufs19168(csa_tree_add_6_33_groupi_n_168 ,csa_tree_add_6_33_groupi_n_887);
  not csa_tree_add_6_33_groupi_drc_bufs19170(csa_tree_add_6_33_groupi_n_167 ,csa_tree_add_6_33_groupi_n_165);
  not csa_tree_add_6_33_groupi_drc_bufs19171(csa_tree_add_6_33_groupi_n_166 ,csa_tree_add_6_33_groupi_n_165);
  not csa_tree_add_6_33_groupi_drc_bufs19172(csa_tree_add_6_33_groupi_n_165 ,csa_tree_add_6_33_groupi_n_910);
  not csa_tree_add_6_33_groupi_drc_bufs19174(csa_tree_add_6_33_groupi_n_164 ,csa_tree_add_6_33_groupi_n_162);
  not csa_tree_add_6_33_groupi_drc_bufs19175(csa_tree_add_6_33_groupi_n_163 ,csa_tree_add_6_33_groupi_n_162);
  not csa_tree_add_6_33_groupi_drc_bufs19176(csa_tree_add_6_33_groupi_n_162 ,csa_tree_add_6_33_groupi_n_981);
  not csa_tree_add_6_33_groupi_drc_bufs19178(csa_tree_add_6_33_groupi_n_161 ,csa_tree_add_6_33_groupi_n_159);
  not csa_tree_add_6_33_groupi_drc_bufs19179(csa_tree_add_6_33_groupi_n_160 ,csa_tree_add_6_33_groupi_n_159);
  not csa_tree_add_6_33_groupi_drc_bufs19180(csa_tree_add_6_33_groupi_n_159 ,csa_tree_add_6_33_groupi_n_989);
  not csa_tree_add_6_33_groupi_drc_bufs19182(csa_tree_add_6_33_groupi_n_158 ,csa_tree_add_6_33_groupi_n_156);
  not csa_tree_add_6_33_groupi_drc_bufs19183(csa_tree_add_6_33_groupi_n_157 ,csa_tree_add_6_33_groupi_n_156);
  not csa_tree_add_6_33_groupi_drc_bufs19184(csa_tree_add_6_33_groupi_n_156 ,csa_tree_add_6_33_groupi_n_961);
  not csa_tree_add_6_33_groupi_drc_bufs19186(csa_tree_add_6_33_groupi_n_155 ,csa_tree_add_6_33_groupi_n_153);
  not csa_tree_add_6_33_groupi_drc_bufs19187(csa_tree_add_6_33_groupi_n_154 ,csa_tree_add_6_33_groupi_n_153);
  not csa_tree_add_6_33_groupi_drc_bufs19188(csa_tree_add_6_33_groupi_n_153 ,csa_tree_add_6_33_groupi_n_978);
  not csa_tree_add_6_33_groupi_drc_bufs19190(csa_tree_add_6_33_groupi_n_152 ,csa_tree_add_6_33_groupi_n_150);
  not csa_tree_add_6_33_groupi_drc_bufs19191(csa_tree_add_6_33_groupi_n_151 ,csa_tree_add_6_33_groupi_n_150);
  not csa_tree_add_6_33_groupi_drc_bufs19192(csa_tree_add_6_33_groupi_n_150 ,csa_tree_add_6_33_groupi_n_993);
  not csa_tree_add_6_33_groupi_drc_bufs19194(csa_tree_add_6_33_groupi_n_149 ,csa_tree_add_6_33_groupi_n_147);
  not csa_tree_add_6_33_groupi_drc_bufs19195(csa_tree_add_6_33_groupi_n_148 ,csa_tree_add_6_33_groupi_n_147);
  not csa_tree_add_6_33_groupi_drc_bufs19196(csa_tree_add_6_33_groupi_n_147 ,csa_tree_add_6_33_groupi_n_883);
  not csa_tree_add_6_33_groupi_drc_bufs19198(csa_tree_add_6_33_groupi_n_146 ,csa_tree_add_6_33_groupi_n_144);
  not csa_tree_add_6_33_groupi_drc_bufs19199(csa_tree_add_6_33_groupi_n_145 ,csa_tree_add_6_33_groupi_n_144);
  not csa_tree_add_6_33_groupi_drc_bufs19200(csa_tree_add_6_33_groupi_n_144 ,csa_tree_add_6_33_groupi_n_957);
  not csa_tree_add_6_33_groupi_drc_bufs19202(csa_tree_add_6_33_groupi_n_143 ,csa_tree_add_6_33_groupi_n_141);
  not csa_tree_add_6_33_groupi_drc_bufs19203(csa_tree_add_6_33_groupi_n_142 ,csa_tree_add_6_33_groupi_n_141);
  not csa_tree_add_6_33_groupi_drc_bufs19204(csa_tree_add_6_33_groupi_n_141 ,csa_tree_add_6_33_groupi_n_897);
  not csa_tree_add_6_33_groupi_drc_bufs19206(csa_tree_add_6_33_groupi_n_140 ,csa_tree_add_6_33_groupi_n_138);
  not csa_tree_add_6_33_groupi_drc_bufs19207(csa_tree_add_6_33_groupi_n_139 ,csa_tree_add_6_33_groupi_n_138);
  not csa_tree_add_6_33_groupi_drc_bufs19208(csa_tree_add_6_33_groupi_n_138 ,csa_tree_add_6_33_groupi_n_973);
  not csa_tree_add_6_33_groupi_drc_bufs19210(csa_tree_add_6_33_groupi_n_137 ,csa_tree_add_6_33_groupi_n_135);
  not csa_tree_add_6_33_groupi_drc_bufs19211(csa_tree_add_6_33_groupi_n_136 ,csa_tree_add_6_33_groupi_n_135);
  not csa_tree_add_6_33_groupi_drc_bufs19212(csa_tree_add_6_33_groupi_n_135 ,csa_tree_add_6_33_groupi_n_1005);
  not csa_tree_add_6_33_groupi_drc_bufs19214(csa_tree_add_6_33_groupi_n_134 ,csa_tree_add_6_33_groupi_n_132);
  not csa_tree_add_6_33_groupi_drc_bufs19215(csa_tree_add_6_33_groupi_n_133 ,csa_tree_add_6_33_groupi_n_132);
  not csa_tree_add_6_33_groupi_drc_bufs19216(csa_tree_add_6_33_groupi_n_132 ,csa_tree_add_6_33_groupi_n_950);
  not csa_tree_add_6_33_groupi_drc_bufs19218(csa_tree_add_6_33_groupi_n_131 ,csa_tree_add_6_33_groupi_n_129);
  not csa_tree_add_6_33_groupi_drc_bufs19219(csa_tree_add_6_33_groupi_n_130 ,csa_tree_add_6_33_groupi_n_129);
  not csa_tree_add_6_33_groupi_drc_bufs19220(csa_tree_add_6_33_groupi_n_129 ,csa_tree_add_6_33_groupi_n_889);
  not csa_tree_add_6_33_groupi_drc_bufs19222(csa_tree_add_6_33_groupi_n_128 ,csa_tree_add_6_33_groupi_n_126);
  not csa_tree_add_6_33_groupi_drc_bufs19223(csa_tree_add_6_33_groupi_n_127 ,csa_tree_add_6_33_groupi_n_126);
  not csa_tree_add_6_33_groupi_drc_bufs19224(csa_tree_add_6_33_groupi_n_126 ,csa_tree_add_6_33_groupi_n_913);
  not csa_tree_add_6_33_groupi_drc_bufs19226(csa_tree_add_6_33_groupi_n_125 ,csa_tree_add_6_33_groupi_n_123);
  not csa_tree_add_6_33_groupi_drc_bufs19227(csa_tree_add_6_33_groupi_n_124 ,csa_tree_add_6_33_groupi_n_123);
  not csa_tree_add_6_33_groupi_drc_bufs19228(csa_tree_add_6_33_groupi_n_123 ,csa_tree_add_6_33_groupi_n_909);
  not csa_tree_add_6_33_groupi_drc_bufs19230(csa_tree_add_6_33_groupi_n_122 ,csa_tree_add_6_33_groupi_n_120);
  not csa_tree_add_6_33_groupi_drc_bufs19231(csa_tree_add_6_33_groupi_n_121 ,csa_tree_add_6_33_groupi_n_120);
  not csa_tree_add_6_33_groupi_drc_bufs19232(csa_tree_add_6_33_groupi_n_120 ,csa_tree_add_6_33_groupi_n_881);
  not csa_tree_add_6_33_groupi_drc_bufs19234(csa_tree_add_6_33_groupi_n_119 ,csa_tree_add_6_33_groupi_n_117);
  not csa_tree_add_6_33_groupi_drc_bufs19235(csa_tree_add_6_33_groupi_n_118 ,csa_tree_add_6_33_groupi_n_117);
  not csa_tree_add_6_33_groupi_drc_bufs19236(csa_tree_add_6_33_groupi_n_117 ,csa_tree_add_6_33_groupi_n_898);
  not csa_tree_add_6_33_groupi_drc_bufs19238(csa_tree_add_6_33_groupi_n_116 ,csa_tree_add_6_33_groupi_n_114);
  not csa_tree_add_6_33_groupi_drc_bufs19239(csa_tree_add_6_33_groupi_n_115 ,csa_tree_add_6_33_groupi_n_114);
  not csa_tree_add_6_33_groupi_drc_bufs19240(csa_tree_add_6_33_groupi_n_114 ,csa_tree_add_6_33_groupi_n_887);
  not csa_tree_add_6_33_groupi_drc_bufs19242(csa_tree_add_6_33_groupi_n_113 ,csa_tree_add_6_33_groupi_n_111);
  not csa_tree_add_6_33_groupi_drc_bufs19243(csa_tree_add_6_33_groupi_n_112 ,csa_tree_add_6_33_groupi_n_111);
  not csa_tree_add_6_33_groupi_drc_bufs19244(csa_tree_add_6_33_groupi_n_111 ,csa_tree_add_6_33_groupi_n_902);
  not csa_tree_add_6_33_groupi_drc_bufs19246(csa_tree_add_6_33_groupi_n_110 ,csa_tree_add_6_33_groupi_n_108);
  not csa_tree_add_6_33_groupi_drc_bufs19247(csa_tree_add_6_33_groupi_n_109 ,csa_tree_add_6_33_groupi_n_108);
  not csa_tree_add_6_33_groupi_drc_bufs19248(csa_tree_add_6_33_groupi_n_108 ,csa_tree_add_6_33_groupi_n_910);
  not csa_tree_add_6_33_groupi_drc_bufs19250(csa_tree_add_6_33_groupi_n_107 ,csa_tree_add_6_33_groupi_n_105);
  not csa_tree_add_6_33_groupi_drc_bufs19251(csa_tree_add_6_33_groupi_n_106 ,csa_tree_add_6_33_groupi_n_105);
  not csa_tree_add_6_33_groupi_drc_bufs19252(csa_tree_add_6_33_groupi_n_105 ,csa_tree_add_6_33_groupi_n_886);
  not csa_tree_add_6_33_groupi_drc_bufs19254(csa_tree_add_6_33_groupi_n_104 ,csa_tree_add_6_33_groupi_n_102);
  not csa_tree_add_6_33_groupi_drc_bufs19255(csa_tree_add_6_33_groupi_n_103 ,csa_tree_add_6_33_groupi_n_102);
  not csa_tree_add_6_33_groupi_drc_bufs19256(csa_tree_add_6_33_groupi_n_102 ,csa_tree_add_6_33_groupi_n_888);
  not csa_tree_add_6_33_groupi_drc_bufs19258(csa_tree_add_6_33_groupi_n_101 ,csa_tree_add_6_33_groupi_n_99);
  not csa_tree_add_6_33_groupi_drc_bufs19259(csa_tree_add_6_33_groupi_n_100 ,csa_tree_add_6_33_groupi_n_99);
  not csa_tree_add_6_33_groupi_drc_bufs19260(csa_tree_add_6_33_groupi_n_99 ,csa_tree_add_6_33_groupi_n_894);
  not csa_tree_add_6_33_groupi_drc_bufs19262(csa_tree_add_6_33_groupi_n_98 ,csa_tree_add_6_33_groupi_n_96);
  not csa_tree_add_6_33_groupi_drc_bufs19263(csa_tree_add_6_33_groupi_n_97 ,csa_tree_add_6_33_groupi_n_96);
  not csa_tree_add_6_33_groupi_drc_bufs19264(csa_tree_add_6_33_groupi_n_96 ,csa_tree_add_6_33_groupi_n_891);
  not csa_tree_add_6_33_groupi_drc_bufs19266(csa_tree_add_6_33_groupi_n_95 ,csa_tree_add_6_33_groupi_n_93);
  not csa_tree_add_6_33_groupi_drc_bufs19267(csa_tree_add_6_33_groupi_n_94 ,csa_tree_add_6_33_groupi_n_93);
  not csa_tree_add_6_33_groupi_drc_bufs19268(csa_tree_add_6_33_groupi_n_93 ,csa_tree_add_6_33_groupi_n_930);
  not csa_tree_add_6_33_groupi_drc_bufs19270(csa_tree_add_6_33_groupi_n_92 ,csa_tree_add_6_33_groupi_n_90);
  not csa_tree_add_6_33_groupi_drc_bufs19271(csa_tree_add_6_33_groupi_n_91 ,csa_tree_add_6_33_groupi_n_90);
  not csa_tree_add_6_33_groupi_drc_bufs19272(csa_tree_add_6_33_groupi_n_90 ,csa_tree_add_6_33_groupi_n_895);
  not csa_tree_add_6_33_groupi_drc_bufs19274(csa_tree_add_6_33_groupi_n_89 ,csa_tree_add_6_33_groupi_n_87);
  not csa_tree_add_6_33_groupi_drc_bufs19275(csa_tree_add_6_33_groupi_n_88 ,csa_tree_add_6_33_groupi_n_87);
  not csa_tree_add_6_33_groupi_drc_bufs19276(csa_tree_add_6_33_groupi_n_87 ,csa_tree_add_6_33_groupi_n_878);
  not csa_tree_add_6_33_groupi_drc_bufs19278(csa_tree_add_6_33_groupi_n_86 ,csa_tree_add_6_33_groupi_n_84);
  not csa_tree_add_6_33_groupi_drc_bufs19279(csa_tree_add_6_33_groupi_n_85 ,csa_tree_add_6_33_groupi_n_84);
  not csa_tree_add_6_33_groupi_drc_bufs19280(csa_tree_add_6_33_groupi_n_84 ,csa_tree_add_6_33_groupi_n_922);
  not csa_tree_add_6_33_groupi_drc_bufs19282(csa_tree_add_6_33_groupi_n_83 ,csa_tree_add_6_33_groupi_n_81);
  not csa_tree_add_6_33_groupi_drc_bufs19283(csa_tree_add_6_33_groupi_n_82 ,csa_tree_add_6_33_groupi_n_81);
  not csa_tree_add_6_33_groupi_drc_bufs19284(csa_tree_add_6_33_groupi_n_81 ,csa_tree_add_6_33_groupi_n_882);
  not csa_tree_add_6_33_groupi_drc_bufs19286(csa_tree_add_6_33_groupi_n_80 ,csa_tree_add_6_33_groupi_n_78);
  not csa_tree_add_6_33_groupi_drc_bufs19287(csa_tree_add_6_33_groupi_n_79 ,csa_tree_add_6_33_groupi_n_78);
  not csa_tree_add_6_33_groupi_drc_bufs19288(csa_tree_add_6_33_groupi_n_78 ,csa_tree_add_6_33_groupi_n_906);
  not csa_tree_add_6_33_groupi_drc_bufs19290(csa_tree_add_6_33_groupi_n_77 ,csa_tree_add_6_33_groupi_n_75);
  not csa_tree_add_6_33_groupi_drc_bufs19291(csa_tree_add_6_33_groupi_n_76 ,csa_tree_add_6_33_groupi_n_75);
  not csa_tree_add_6_33_groupi_drc_bufs19292(csa_tree_add_6_33_groupi_n_75 ,csa_tree_add_6_33_groupi_n_879);
  not csa_tree_add_6_33_groupi_drc_bufs19294(csa_tree_add_6_33_groupi_n_74 ,csa_tree_add_6_33_groupi_n_72);
  not csa_tree_add_6_33_groupi_drc_bufs19295(csa_tree_add_6_33_groupi_n_73 ,csa_tree_add_6_33_groupi_n_72);
  not csa_tree_add_6_33_groupi_drc_bufs19296(csa_tree_add_6_33_groupi_n_72 ,csa_tree_add_6_33_groupi_n_918);
  not csa_tree_add_6_33_groupi_drc_bufs19298(csa_tree_add_6_33_groupi_n_71 ,csa_tree_add_6_33_groupi_n_69);
  not csa_tree_add_6_33_groupi_drc_bufs19299(csa_tree_add_6_33_groupi_n_70 ,csa_tree_add_6_33_groupi_n_69);
  not csa_tree_add_6_33_groupi_drc_bufs19300(csa_tree_add_6_33_groupi_n_69 ,csa_tree_add_6_33_groupi_n_899);
  not csa_tree_add_6_33_groupi_drc_bufs19302(csa_tree_add_6_33_groupi_n_68 ,csa_tree_add_6_33_groupi_n_66);
  not csa_tree_add_6_33_groupi_drc_bufs19303(csa_tree_add_6_33_groupi_n_67 ,csa_tree_add_6_33_groupi_n_66);
  not csa_tree_add_6_33_groupi_drc_bufs19304(csa_tree_add_6_33_groupi_n_66 ,csa_tree_add_6_33_groupi_n_926);
  not csa_tree_add_6_33_groupi_drc_bufs19306(csa_tree_add_6_33_groupi_n_65 ,csa_tree_add_6_33_groupi_n_63);
  not csa_tree_add_6_33_groupi_drc_bufs19307(csa_tree_add_6_33_groupi_n_64 ,csa_tree_add_6_33_groupi_n_63);
  not csa_tree_add_6_33_groupi_drc_bufs19308(csa_tree_add_6_33_groupi_n_63 ,csa_tree_add_6_33_groupi_n_890);
  not csa_tree_add_6_33_groupi_drc_bufs19310(csa_tree_add_6_33_groupi_n_62 ,csa_tree_add_6_33_groupi_n_60);
  not csa_tree_add_6_33_groupi_drc_bufs19311(csa_tree_add_6_33_groupi_n_61 ,csa_tree_add_6_33_groupi_n_60);
  not csa_tree_add_6_33_groupi_drc_bufs19312(csa_tree_add_6_33_groupi_n_60 ,csa_tree_add_6_33_groupi_n_934);
  not csa_tree_add_6_33_groupi_drc_bufs19314(csa_tree_add_6_33_groupi_n_59 ,csa_tree_add_6_33_groupi_n_57);
  not csa_tree_add_6_33_groupi_drc_bufs19315(csa_tree_add_6_33_groupi_n_58 ,csa_tree_add_6_33_groupi_n_57);
  not csa_tree_add_6_33_groupi_drc_bufs19316(csa_tree_add_6_33_groupi_n_57 ,csa_tree_add_6_33_groupi_n_883);
  not csa_tree_add_6_33_groupi_drc_bufs19318(csa_tree_add_6_33_groupi_n_56 ,csa_tree_add_6_33_groupi_n_54);
  not csa_tree_add_6_33_groupi_drc_bufs19319(csa_tree_add_6_33_groupi_n_55 ,csa_tree_add_6_33_groupi_n_54);
  not csa_tree_add_6_33_groupi_drc_bufs19320(csa_tree_add_6_33_groupi_n_54 ,csa_tree_add_6_33_groupi_n_884);
  not csa_tree_add_6_33_groupi_drc_bufs19322(csa_tree_add_6_33_groupi_n_53 ,csa_tree_add_6_33_groupi_n_51);
  not csa_tree_add_6_33_groupi_drc_bufs19323(csa_tree_add_6_33_groupi_n_52 ,csa_tree_add_6_33_groupi_n_51);
  not csa_tree_add_6_33_groupi_drc_bufs19324(csa_tree_add_6_33_groupi_n_51 ,csa_tree_add_6_33_groupi_n_914);
  not csa_tree_add_6_33_groupi_drc_bufs19326(csa_tree_add_6_33_groupi_n_50 ,csa_tree_add_6_33_groupi_n_48);
  not csa_tree_add_6_33_groupi_drc_bufs19327(csa_tree_add_6_33_groupi_n_49 ,csa_tree_add_6_33_groupi_n_48);
  not csa_tree_add_6_33_groupi_drc_bufs19328(csa_tree_add_6_33_groupi_n_48 ,csa_tree_add_6_33_groupi_n_903);
  not csa_tree_add_6_33_groupi_drc_bufs19330(csa_tree_add_6_33_groupi_n_47 ,csa_tree_add_6_33_groupi_n_45);
  not csa_tree_add_6_33_groupi_drc_bufs19331(csa_tree_add_6_33_groupi_n_46 ,csa_tree_add_6_33_groupi_n_45);
  not csa_tree_add_6_33_groupi_drc_bufs19332(csa_tree_add_6_33_groupi_n_45 ,csa_tree_add_6_33_groupi_n_880);
  not csa_tree_add_6_33_groupi_drc_bufs19334(csa_tree_add_6_33_groupi_n_44 ,csa_tree_add_6_33_groupi_n_43);
  not csa_tree_add_6_33_groupi_drc_bufs19336(csa_tree_add_6_33_groupi_n_43 ,csa_tree_add_6_33_groupi_n_812);
  not csa_tree_add_6_33_groupi_drc_bufs19338(csa_tree_add_6_33_groupi_n_42 ,csa_tree_add_6_33_groupi_n_41);
  not csa_tree_add_6_33_groupi_drc_bufs19340(csa_tree_add_6_33_groupi_n_41 ,csa_tree_add_6_33_groupi_n_773);
  not csa_tree_add_6_33_groupi_drc_bufs19342(csa_tree_add_6_33_groupi_n_40 ,csa_tree_add_6_33_groupi_n_39);
  not csa_tree_add_6_33_groupi_drc_bufs19344(csa_tree_add_6_33_groupi_n_39 ,csa_tree_add_6_33_groupi_n_776);
  not csa_tree_add_6_33_groupi_drc_bufs19346(csa_tree_add_6_33_groupi_n_38 ,csa_tree_add_6_33_groupi_n_37);
  not csa_tree_add_6_33_groupi_drc_bufs19348(csa_tree_add_6_33_groupi_n_37 ,csa_tree_add_6_33_groupi_n_779);
  not csa_tree_add_6_33_groupi_drc_bufs19350(csa_tree_add_6_33_groupi_n_36 ,csa_tree_add_6_33_groupi_n_35);
  not csa_tree_add_6_33_groupi_drc_bufs19352(csa_tree_add_6_33_groupi_n_35 ,csa_tree_add_6_33_groupi_n_782);
  not csa_tree_add_6_33_groupi_drc_bufs19354(csa_tree_add_6_33_groupi_n_34 ,csa_tree_add_6_33_groupi_n_33);
  not csa_tree_add_6_33_groupi_drc_bufs19356(csa_tree_add_6_33_groupi_n_33 ,csa_tree_add_6_33_groupi_n_785);
  not csa_tree_add_6_33_groupi_drc_bufs19358(csa_tree_add_6_33_groupi_n_32 ,csa_tree_add_6_33_groupi_n_31);
  not csa_tree_add_6_33_groupi_drc_bufs19360(csa_tree_add_6_33_groupi_n_31 ,csa_tree_add_6_33_groupi_n_788);
  not csa_tree_add_6_33_groupi_drc_bufs19362(csa_tree_add_6_33_groupi_n_30 ,csa_tree_add_6_33_groupi_n_29);
  not csa_tree_add_6_33_groupi_drc_bufs19364(csa_tree_add_6_33_groupi_n_29 ,csa_tree_add_6_33_groupi_n_791);
  not csa_tree_add_6_33_groupi_drc_bufs19366(csa_tree_add_6_33_groupi_n_28 ,csa_tree_add_6_33_groupi_n_27);
  not csa_tree_add_6_33_groupi_drc_bufs19368(csa_tree_add_6_33_groupi_n_27 ,csa_tree_add_6_33_groupi_n_794);
  not csa_tree_add_6_33_groupi_drc_bufs19370(csa_tree_add_6_33_groupi_n_26 ,csa_tree_add_6_33_groupi_n_25);
  not csa_tree_add_6_33_groupi_drc_bufs19372(csa_tree_add_6_33_groupi_n_25 ,csa_tree_add_6_33_groupi_n_797);
  not csa_tree_add_6_33_groupi_drc_bufs19374(csa_tree_add_6_33_groupi_n_24 ,csa_tree_add_6_33_groupi_n_23);
  not csa_tree_add_6_33_groupi_drc_bufs19376(csa_tree_add_6_33_groupi_n_23 ,csa_tree_add_6_33_groupi_n_800);
  not csa_tree_add_6_33_groupi_drc_bufs19378(csa_tree_add_6_33_groupi_n_22 ,csa_tree_add_6_33_groupi_n_21);
  not csa_tree_add_6_33_groupi_drc_bufs19380(csa_tree_add_6_33_groupi_n_21 ,csa_tree_add_6_33_groupi_n_803);
  not csa_tree_add_6_33_groupi_drc_bufs19382(csa_tree_add_6_33_groupi_n_20 ,csa_tree_add_6_33_groupi_n_19);
  not csa_tree_add_6_33_groupi_drc_bufs19384(csa_tree_add_6_33_groupi_n_19 ,csa_tree_add_6_33_groupi_n_806);
  not csa_tree_add_6_33_groupi_drc_bufs19386(csa_tree_add_6_33_groupi_n_18 ,csa_tree_add_6_33_groupi_n_17);
  not csa_tree_add_6_33_groupi_drc_bufs19388(csa_tree_add_6_33_groupi_n_17 ,csa_tree_add_6_33_groupi_n_809);
  xor csa_tree_add_6_33_groupi_g2(out1[61] ,csa_tree_add_6_33_groupi_n_4961 ,csa_tree_add_6_33_groupi_n_2933);
  xor csa_tree_add_6_33_groupi_g19390(out1[59] ,csa_tree_add_6_33_groupi_n_4956 ,csa_tree_add_6_33_groupi_n_3782);
  xor csa_tree_add_6_33_groupi_g19391(out1[57] ,csa_tree_add_6_33_groupi_n_4951 ,csa_tree_add_6_33_groupi_n_3926);
  xor csa_tree_add_6_33_groupi_g19392(out1[56] ,csa_tree_add_6_33_groupi_n_4949 ,csa_tree_add_6_33_groupi_n_4190);
  xor csa_tree_add_6_33_groupi_g19393(out1[55] ,csa_tree_add_6_33_groupi_n_4947 ,csa_tree_add_6_33_groupi_n_4303);
  xor csa_tree_add_6_33_groupi_g19394(out1[53] ,csa_tree_add_6_33_groupi_n_4942 ,csa_tree_add_6_33_groupi_n_4401);
  xor csa_tree_add_6_33_groupi_g19395(out1[39] ,csa_tree_add_6_33_groupi_n_4896 ,csa_tree_add_6_33_groupi_n_4792);
  xor csa_tree_add_6_33_groupi_g19396(out1[30] ,csa_tree_add_6_33_groupi_n_4868 ,csa_tree_add_6_33_groupi_n_4810);
  xor csa_tree_add_6_33_groupi_g19397(out1[25] ,csa_tree_add_6_33_groupi_n_4854 ,csa_tree_add_6_33_groupi_n_4760);
  xor csa_tree_add_6_33_groupi_g19398(out1[24] ,csa_tree_add_6_33_groupi_n_4852 ,csa_tree_add_6_33_groupi_n_4759);
  xor csa_tree_add_6_33_groupi_g19399(out1[18] ,csa_tree_add_6_33_groupi_n_4834 ,csa_tree_add_6_33_groupi_n_4673);
  xor csa_tree_add_6_33_groupi_g19400(out1[17] ,csa_tree_add_6_33_groupi_n_4832 ,csa_tree_add_6_33_groupi_n_4545);
  xor csa_tree_add_6_33_groupi_g19401(out1[16] ,csa_tree_add_6_33_groupi_n_4830 ,csa_tree_add_6_33_groupi_n_4544);
  xor csa_tree_add_6_33_groupi_g19402(out1[15] ,csa_tree_add_6_33_groupi_n_4828 ,csa_tree_add_6_33_groupi_n_4543);
  xor csa_tree_add_6_33_groupi_g19403(out1[14] ,csa_tree_add_6_33_groupi_n_4826 ,csa_tree_add_6_33_groupi_n_4391);
  xor csa_tree_add_6_33_groupi_g19404(csa_tree_add_6_33_groupi_n_1 ,csa_tree_add_6_33_groupi_n_4539 ,csa_tree_add_6_33_groupi_n_4624);
  xor csa_tree_add_6_33_groupi_g19405(csa_tree_add_6_33_groupi_n_0 ,csa_tree_add_6_33_groupi_n_3848 ,csa_tree_add_6_33_groupi_n_1007);
  not g19406(csa_tree_add_6_33_groupi_n_2013 ,csa_tree_add_6_33_groupi_n_339);
  not g19407(csa_tree_add_6_33_groupi_n_1921 ,csa_tree_add_6_33_groupi_n_297);
  buf g19408(csa_tree_add_6_33_groupi_n_2320 ,csa_tree_add_6_33_groupi_n_1320);
  buf g19409(csa_tree_add_6_33_groupi_n_2220 ,csa_tree_add_6_33_groupi_n_1539);
  buf g19410(csa_tree_add_6_33_groupi_n_2275 ,csa_tree_add_6_33_groupi_n_1265);
  buf g19411(csa_tree_add_6_33_groupi_n_2297 ,csa_tree_add_6_33_groupi_n_1547);
  buf g19412(csa_tree_add_6_33_groupi_n_2284 ,csa_tree_add_6_33_groupi_n_1285);
  buf g19413(csa_tree_add_6_33_groupi_n_2208 ,csa_tree_add_6_33_groupi_n_1598);
  buf g19414(csa_tree_add_6_33_groupi_n_2209 ,csa_tree_add_6_33_groupi_n_1313);
  buf g19415(csa_tree_add_6_33_groupi_n_2238 ,csa_tree_add_6_33_groupi_n_1568);
  buf g19416(csa_tree_add_6_33_groupi_n_2245 ,csa_tree_add_6_33_groupi_n_1279);
endmodule
