module top(in1, in2, in3, out1);
  input [3:0] in1, in2, in3;
  output [3:0] out1;
  wire [3:0] in1, in2, in3;
  wire [3:0] out1;
  wire csa_tree_ADD_TC_OP_1_groupi_n_0, csa_tree_ADD_TC_OP_1_groupi_n_1, csa_tree_ADD_TC_OP_1_groupi_n_2, csa_tree_ADD_TC_OP_1_groupi_n_3, csa_tree_ADD_TC_OP_1_groupi_n_4, csa_tree_ADD_TC_OP_1_groupi_n_5, csa_tree_ADD_TC_OP_1_groupi_n_6, csa_tree_ADD_TC_OP_1_groupi_n_7;
  wire csa_tree_ADD_TC_OP_1_groupi_n_8, csa_tree_ADD_TC_OP_1_groupi_n_9, csa_tree_ADD_TC_OP_1_groupi_n_10, csa_tree_ADD_TC_OP_1_groupi_n_11, csa_tree_ADD_TC_OP_1_groupi_n_12, csa_tree_ADD_TC_OP_1_groupi_n_13, csa_tree_ADD_TC_OP_1_groupi_n_14, csa_tree_ADD_TC_OP_1_groupi_n_15;
  wire csa_tree_ADD_TC_OP_1_groupi_n_16, csa_tree_ADD_TC_OP_1_groupi_n_17, csa_tree_ADD_TC_OP_1_groupi_n_18, csa_tree_ADD_TC_OP_1_groupi_n_19, csa_tree_ADD_TC_OP_1_groupi_n_21, csa_tree_ADD_TC_OP_1_groupi_n_22, csa_tree_ADD_TC_OP_1_groupi_n_23, csa_tree_ADD_TC_OP_1_groupi_n_24;
  wire csa_tree_ADD_TC_OP_1_groupi_n_25, csa_tree_ADD_TC_OP_1_groupi_n_26, csa_tree_ADD_TC_OP_1_groupi_n_27, csa_tree_ADD_TC_OP_1_groupi_n_29, csa_tree_ADD_TC_OP_1_groupi_n_30, csa_tree_ADD_TC_OP_1_groupi_n_31, csa_tree_ADD_TC_OP_1_groupi_n_32;
  xnor csa_tree_ADD_TC_OP_1_groupi_g111__2398(out1[3] ,csa_tree_ADD_TC_OP_1_groupi_n_29 ,csa_tree_ADD_TC_OP_1_groupi_n_32);
  xor csa_tree_ADD_TC_OP_1_groupi_g112__5107(out1[2] ,csa_tree_ADD_TC_OP_1_groupi_n_26 ,csa_tree_ADD_TC_OP_1_groupi_n_30);
  or csa_tree_ADD_TC_OP_1_groupi_g113__6260(csa_tree_ADD_TC_OP_1_groupi_n_32 ,csa_tree_ADD_TC_OP_1_groupi_n_25 ,csa_tree_ADD_TC_OP_1_groupi_n_31);
  and csa_tree_ADD_TC_OP_1_groupi_g114__4319(csa_tree_ADD_TC_OP_1_groupi_n_31 ,csa_tree_ADD_TC_OP_1_groupi_n_27 ,csa_tree_ADD_TC_OP_1_groupi_n_26);
  xnor csa_tree_ADD_TC_OP_1_groupi_g115__8428(csa_tree_ADD_TC_OP_1_groupi_n_30 ,csa_tree_ADD_TC_OP_1_groupi_n_5 ,csa_tree_ADD_TC_OP_1_groupi_n_22);
  xnor csa_tree_ADD_TC_OP_1_groupi_g116__5526(csa_tree_ADD_TC_OP_1_groupi_n_29 ,csa_tree_ADD_TC_OP_1_groupi_n_17 ,csa_tree_ADD_TC_OP_1_groupi_n_23);
  xor csa_tree_ADD_TC_OP_1_groupi_g117__6783(out1[1] ,csa_tree_ADD_TC_OP_1_groupi_n_16 ,csa_tree_ADD_TC_OP_1_groupi_n_21);
  or csa_tree_ADD_TC_OP_1_groupi_g118__3680(csa_tree_ADD_TC_OP_1_groupi_n_27 ,csa_tree_ADD_TC_OP_1_groupi_n_6 ,csa_tree_ADD_TC_OP_1_groupi_n_22);
  or csa_tree_ADD_TC_OP_1_groupi_g119__1617(csa_tree_ADD_TC_OP_1_groupi_n_26 ,csa_tree_ADD_TC_OP_1_groupi_n_19 ,csa_tree_ADD_TC_OP_1_groupi_n_24);
  and csa_tree_ADD_TC_OP_1_groupi_g120__2802(csa_tree_ADD_TC_OP_1_groupi_n_25 ,csa_tree_ADD_TC_OP_1_groupi_n_6 ,csa_tree_ADD_TC_OP_1_groupi_n_22);
  and csa_tree_ADD_TC_OP_1_groupi_g121__1705(csa_tree_ADD_TC_OP_1_groupi_n_24 ,csa_tree_ADD_TC_OP_1_groupi_n_16 ,csa_tree_ADD_TC_OP_1_groupi_n_18);
  xnor csa_tree_ADD_TC_OP_1_groupi_g122__5122(csa_tree_ADD_TC_OP_1_groupi_n_23 ,csa_tree_ADD_TC_OP_1_groupi_n_10 ,in1[3]);
  xnor csa_tree_ADD_TC_OP_1_groupi_g123__8246(csa_tree_ADD_TC_OP_1_groupi_n_22 ,csa_tree_ADD_TC_OP_1_groupi_n_9 ,in1[2]);
  xnor csa_tree_ADD_TC_OP_1_groupi_g124__7098(csa_tree_ADD_TC_OP_1_groupi_n_21 ,csa_tree_ADD_TC_OP_1_groupi_n_12 ,in2[1]);
  xnor csa_tree_ADD_TC_OP_1_groupi_g125__6131(out1[0] ,csa_tree_ADD_TC_OP_1_groupi_n_13 ,in3[0]);
  nor csa_tree_ADD_TC_OP_1_groupi_g126__1881(csa_tree_ADD_TC_OP_1_groupi_n_19 ,csa_tree_ADD_TC_OP_1_groupi_n_1 ,csa_tree_ADD_TC_OP_1_groupi_n_12);
  or csa_tree_ADD_TC_OP_1_groupi_g127__5115(csa_tree_ADD_TC_OP_1_groupi_n_18 ,in2[1] ,csa_tree_ADD_TC_OP_1_groupi_n_11);
  or csa_tree_ADD_TC_OP_1_groupi_g128__7482(csa_tree_ADD_TC_OP_1_groupi_n_17 ,csa_tree_ADD_TC_OP_1_groupi_n_7 ,csa_tree_ADD_TC_OP_1_groupi_n_15);
  or csa_tree_ADD_TC_OP_1_groupi_g129__4733(csa_tree_ADD_TC_OP_1_groupi_n_16 ,csa_tree_ADD_TC_OP_1_groupi_n_4 ,csa_tree_ADD_TC_OP_1_groupi_n_14);
  and csa_tree_ADD_TC_OP_1_groupi_g130__6161(csa_tree_ADD_TC_OP_1_groupi_n_15 ,in3[2] ,csa_tree_ADD_TC_OP_1_groupi_n_8);
  and csa_tree_ADD_TC_OP_1_groupi_g131__9315(csa_tree_ADD_TC_OP_1_groupi_n_14 ,in1[0] ,csa_tree_ADD_TC_OP_1_groupi_n_3);
  xnor csa_tree_ADD_TC_OP_1_groupi_g132__9945(csa_tree_ADD_TC_OP_1_groupi_n_13 ,in1[0] ,in2[0]);
  not csa_tree_ADD_TC_OP_1_groupi_g133(csa_tree_ADD_TC_OP_1_groupi_n_11 ,csa_tree_ADD_TC_OP_1_groupi_n_12);
  xnor csa_tree_ADD_TC_OP_1_groupi_g134__2883(csa_tree_ADD_TC_OP_1_groupi_n_12 ,in3[1] ,in1[1]);
  xnor csa_tree_ADD_TC_OP_1_groupi_g135__2346(csa_tree_ADD_TC_OP_1_groupi_n_10 ,in3[3] ,in2[3]);
  xnor csa_tree_ADD_TC_OP_1_groupi_g136__1666(csa_tree_ADD_TC_OP_1_groupi_n_9 ,in3[2] ,in2[2]);
  or csa_tree_ADD_TC_OP_1_groupi_g137__7410(csa_tree_ADD_TC_OP_1_groupi_n_8 ,in1[2] ,in2[2]);
  and csa_tree_ADD_TC_OP_1_groupi_g138__6417(csa_tree_ADD_TC_OP_1_groupi_n_7 ,in1[2] ,in2[2]);
  not csa_tree_ADD_TC_OP_1_groupi_g139(csa_tree_ADD_TC_OP_1_groupi_n_6 ,csa_tree_ADD_TC_OP_1_groupi_n_5);
  or csa_tree_ADD_TC_OP_1_groupi_g140__5477(csa_tree_ADD_TC_OP_1_groupi_n_5 ,csa_tree_ADD_TC_OP_1_groupi_n_0 ,csa_tree_ADD_TC_OP_1_groupi_n_2);
  and csa_tree_ADD_TC_OP_1_groupi_g141__2398(csa_tree_ADD_TC_OP_1_groupi_n_4 ,in3[0] ,in2[0]);
  or csa_tree_ADD_TC_OP_1_groupi_g142__5107(csa_tree_ADD_TC_OP_1_groupi_n_3 ,in3[0] ,in2[0]);
  not csa_tree_ADD_TC_OP_1_groupi_g143(csa_tree_ADD_TC_OP_1_groupi_n_2 ,in1[1]);
  not csa_tree_ADD_TC_OP_1_groupi_g144(csa_tree_ADD_TC_OP_1_groupi_n_1 ,in2[1]);
  not csa_tree_ADD_TC_OP_1_groupi_g145(csa_tree_ADD_TC_OP_1_groupi_n_0 ,in3[1]);
endmodule
