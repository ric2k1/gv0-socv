module top( n3 , n4 , n6 , n9 , n10 , n13 , n15 , n18 , n30 , n31 , n33 , n38 , n40 , n44 , n48 , n49 );
    input n3 , n4 , n9 , n13 , n15 , n30 , n31 , n38 , n40 , n44 , n48 , n49 ;
    output n6 , n10 , n18 , n33 ;
    wire n0 , n1 , n2 , n5 , n7 , n8 , n11 , n12 , n14 , n16 , n17 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n32 , n34 , n35 , n36 , n37 , n39 , n41 , n42 , n43 , n45 , n46 , n47 ;
assign n41 = ~(n49 | n48);
assign n33 = ~(n24 ^ n27);
assign n43 = n45 | n42;
assign n19 = n22 & n11;
assign n39 = n1 & n21;
assign n22 = n17 | n20;
assign n2 = ~(n35 | n39);
assign n8 = ~(n9 ^ n40);
assign n17 = ~n44;
assign n34 = n31 & n46;
assign n35 = ~(n15 | n38);
assign n45 = ~n3;
assign n18 = ~(n20 ^ n5);
assign n27 = ~(n8 ^ n47);
assign n26 = ~(n44 | n34);
assign n0 = n37 & n19;
assign n37 = ~n30;
assign n10 = ~(n23 ^ n31);
assign n12 = ~(n39 ^ n16);
assign n14 = ~(n12 | n0);
assign n46 = ~n23;
assign n20 = ~n34;
assign n42 = ~n4;
assign n28 = ~(n43 ^ n7);
assign n11 = n26 | n28;
assign n1 = ~(n49 & n48);
assign n23 = ~(n3 ^ n4);
assign n29 = n25 | n2;
assign n32 = ~(n37 | n19);
assign n21 = n43 | n41;
assign n16 = ~(n15 ^ n38);
assign n24 = ~(n29 ^ n13);
assign n36 = ~(n12 ^ n30);
assign n6 = ~(n19 ^ n36);
assign n7 = ~(n49 ^ n48);
assign n5 = ~(n28 ^ n44);
assign n47 = n32 | n14;
assign n25 = n15 & n38;
endmodule
