module top;
sub s0();
foo f0();
endmodule

module foo;
sub s0();
endmodule
