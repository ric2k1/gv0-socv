module top( n2 , n4 , n6 , n9 , n12 , n18 , n22 , n34 , n35 , n42 , n48 , n51 , n56 , n57 , n65 , n67 , n68 , n72 , n75 , n77 , n78 , n80 );
    input n2 , n4 , n12 , n18 , n22 , n34 , n35 , n51 , n57 , n67 , n72 , n75 , n78 , n80 ;
    output n6 , n9 , n42 , n48 , n56 , n65 , n68 , n77 ;
    wire n0 , n1 , n3 , n5 , n7 , n8 , n10 , n11 , n13 , n14 , n15 , n16 , n17 , n19 , n20 , n21 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n36 , n37 , n38 , n39 , n40 , n41 , n43 , n44 , n45 , n46 , n47 , n49 , n50 , n52 , n53 , n54 , n55 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n66 , n69 , n70 , n71 , n73 , n74 , n76 , n79 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 ;
assign n77 = n86 | n73;
assign n5 = ~(n45 ^ n53);
assign n9 = n61 ^ n30;
assign n40 = ~(n12 | n27);
assign n16 = ~n10;
assign n81 = ~n84;
assign n31 = n34 & n44;
assign n26 = n80 | n2;
assign n58 = n72 & n67;
assign n24 = ~n2;
assign n14 = n21 | n78;
assign n79 = n39 & n1;
assign n20 = n80 | n67;
assign n7 = ~(n84 | n76);
assign n52 = n72 & n57;
assign n50 = n28 & n36;
assign n15 = ~n45;
assign n69 = ~(n0 ^ n50);
assign n3 = ~(n72 & n4);
assign n43 = n22 & n20;
assign n27 = n53 & n16;
assign n21 = ~n4;
assign n60 = n37 | n12;
assign n1 = n55 & n70;
assign n88 = ~n67;
assign n87 = n18 & n26;
assign n48 = ~n63;
assign n71 = ~n57;
assign n6 = ~(n60 ^ n5);
assign n33 = ~(n37 | n77);
assign n59 = n35 & n25;
assign n45 = n54 & n43;
assign n55 = n52 | n64;
assign n29 = ~n75;
assign n74 = ~(n29 | n4);
assign n86 = n90 | n11;
assign n73 = n66 | n45;
assign n42 = n40 ^ n69;
assign n65 = n19 ^ n82;
assign n89 = n9 & n65;
assign n37 = ~n51;
assign n90 = n14 & n59;
assign n25 = n80 | n4;
assign n49 = n3 & n38;
assign n10 = n51 & n15;
assign n61 = ~(n12 | n7);
assign n68 = n33 | n63;
assign n70 = n11 | n47;
assign n36 = ~(n18 | n23);
assign n46 = n71 | n78;
assign n32 = ~(n90 | n1);
assign n39 = n11 | n81;
assign n13 = ~(n29 | n57);
assign n82 = n90 ^ n49;
assign n56 = n8 & n89;
assign n30 = ~(n11 ^ n55);
assign n41 = n22 | n83;
assign n54 = n88 | n78;
assign n17 = ~n72;
assign n19 = ~(n12 | n79);
assign n38 = ~(n35 | n74);
assign n11 = n46 & n31;
assign n23 = ~(n29 | n2);
assign n44 = n80 | n57;
assign n76 = n50 | n62;
assign n66 = n85 & n87;
assign n53 = n58 | n41;
assign n85 = n24 | n78;
assign n83 = ~(n29 | n67);
assign n0 = ~n66;
assign n47 = ~n76;
assign n63 = n49 | n32;
assign n62 = ~(n53 | n66);
assign n8 = n6 & n42;
assign n84 = n0 & n10;
assign n64 = n34 | n13;
assign n28 = n17 | n24;
endmodule
