module top(in1, in2, in3, in4, out1);
  input [15:0] in1, in2, in3;
  input [1:0] in4;
  output [31:0] out1;
  wire [15:0] in1, in2, in3;
  wire [1:0] in4;
  wire [31:0] out1;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_0, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_3, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_4, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_5, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_6, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_7;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_8, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_9, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_10, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_11, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_12, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_13, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_14, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_15;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_16, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_17, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_18, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_19, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_20, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_21, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_22, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_23;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_24, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_25, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_26, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_27, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_29, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_30, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_33, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_34;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_35, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_36, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_37, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_38, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_39, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_40, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_41, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_42;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_43, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_44, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_45, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_46, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_47, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_48, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_49, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_50;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_51, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_52, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_53, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_54, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_55, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_56, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_57, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_58;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_59, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_60, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_61, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_62, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_63, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_64, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_65, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_66;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_67, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_68, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_69, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_70, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_71, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_72, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_73, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_74;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_75, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_76, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_77, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_78, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_79, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_80, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_81, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_82;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_83, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_84, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_85, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_86, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_87, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_88, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_89, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_90;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_91, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_92, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_93, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_94, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_95, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_96, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_97, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_98;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_99, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_100, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_101, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_102, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_103, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_104, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_105, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_106;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_107, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_108, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_109, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_110, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_111, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_112, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_113, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_114;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_115, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_116, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_117, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_118, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_119, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_120, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_121, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_122;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_123, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_124, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_125, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_126, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_127, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_128, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_129, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_130;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_131, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_132, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_133, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_134, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_135, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_136, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_137, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_138;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_139, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_140, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_141, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_142, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_143, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_144, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_145, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_146;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_147, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_148, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_149, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_150, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_151, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_152, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_153, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_154;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_155, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_156, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_157, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_158, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_159, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_160, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_161, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_162;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_163, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_164, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_165, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_166, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_167, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_168, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_169, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_170;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_171, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_172, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_173, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_174, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_175, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_176, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_177, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_178;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_179, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_180, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_181, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_182, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_183, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_184, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_185, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_186;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_187, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_188, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_189, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_190, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_191, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_192, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_193, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_194;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_195, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_196, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_197, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_198, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_199, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_200, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_201, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_202;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_203, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_204, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_205, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_206, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_207, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_208, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_209, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_210;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_211, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_212, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_213, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_214, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_215, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_216, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_217, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_218;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_219, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_220, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_221, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_222, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_223, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_224, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_225, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_226;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_227, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_228, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_229, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_230, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_231, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_232, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_233, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_234;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_235, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_236, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_237, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_238, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_239, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_240, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_241, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_242;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_243, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_244, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_245, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_246, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_247, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_248, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_249, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_250;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_251, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_252, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_253, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_254, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_255, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_256, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_257, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_258;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_259, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_260, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_261, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_262, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_263, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_264, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_265, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_266;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_267, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_268, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_269, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_270, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_271, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_272, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_273, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_274;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_275, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_276, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_277, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_278, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_279, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_280, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_281, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_282;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_283, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_284, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_285, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_286, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_287, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_288, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_289, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_290;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_291, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_292, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_293, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_294, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_295, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_296, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_297, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_298;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_299, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_300, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_301, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_302, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_303, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_304, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_305, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_306;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_307, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_308, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_309, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_310, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_311, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_312, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_313, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_314;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_315, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_316, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_317, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_318, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_319, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_320, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_321, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_322;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_323, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_324, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_325, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_326, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_327, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_328, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_329, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_330;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_331, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_332, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_333, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_334, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_335, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_336, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_337, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_338;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_339, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_340, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_341, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_342, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_343, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_344, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_345, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_346;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_347, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_348, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_349, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_350, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_351, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_352, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_353, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_354;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_355, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_356, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_357, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_358, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_359, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_360, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_361, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_362;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_363, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_364, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_365, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_366, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_367, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_368, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_369, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_370;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_371, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_372, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_373, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_374, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_375, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_376, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_377, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_378;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_379, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_380, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_381, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_382, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_383, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_384, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_385, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_386;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_387, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_388, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_389, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_390, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_391, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_392, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_393, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_394;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_395, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_396, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_397, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_398, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_399, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_400, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_401, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_402;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_403, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_404, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_405, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_406, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_407, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_408, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_409, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_410;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_411, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_412, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_413, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_414, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_415, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_416, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_417, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_418;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_419, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_420, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_421, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_422, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_423, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_424, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_425, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_426;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_427, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_428, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_429, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_430, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_431, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_432, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_433, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_434;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_435, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_436, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_437, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_438, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_439, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_440, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_441, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_442;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_443, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_444, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_445, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_446, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_447, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_448, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_449, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_450;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_451, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_452, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_453, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_454, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_455, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_456, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_457, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_458;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_459, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_460, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_461, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_462, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_463, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_464, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_465, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_466;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_467, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_468, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_469, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_470, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_471, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_472, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_473, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_474;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_475, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_476, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_477, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_478, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_479, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_480, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_481, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_482;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_483, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_484, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_485, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_486, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_487, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_488, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_489, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_490;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_491, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_492, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_493, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_494, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_495, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_496, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_497, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_498;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_499, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_500, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_501, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_502, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_503, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_504, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_505, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_506;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_507, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_508, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_509, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_510, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_511, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_512, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_513, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_514;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_515, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_516, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_517, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_518, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_519, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_520, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_521, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_522;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_523, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_524, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_525, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_526, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_527, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_528, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_529, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_530;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_531, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_532, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_533, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_534, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_535, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_536, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_537, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_538;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_539, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_540, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_541, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_542, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_543, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_544, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_545, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_546;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_547, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_548, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_549, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_550, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_551, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_552, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_553, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_554;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_555, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_556, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_557, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_558, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_559, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_560, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_561, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_562;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_563, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_564, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_565, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_566, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_567, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_568, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_569, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_570;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_571, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_572, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_573, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_574, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_575, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_576, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_577, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_578;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_579, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_580, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_581, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_582, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_583, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_584, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_585, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_586;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_587, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_588, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_589, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_590, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_591, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_592, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_593, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_594;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_595, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_596, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_597, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_598, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_599, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_600, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_601, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_602;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_603, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_604, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_605, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_606, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_607, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_608, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_609, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_610;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_611, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_612, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_613, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_614, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_615, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_616, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_617, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_618;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_619, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_620, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_621, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_622, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_623, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_624, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_625, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_626;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_627, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_628, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_629, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_630, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_631, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_632, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_633, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_634;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_635, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_636, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_637, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_638, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_639, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_640, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_641, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_642;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_643, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_644, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_645, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_646, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_647, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_648, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_649, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_650;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_651, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_652, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_653, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_654, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_655, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_656, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_657, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_658;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_659, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_660, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_661, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_662, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_663, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_664, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_665, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_666;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_667, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_668, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_669, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_670, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_671, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_672, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_673, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_674;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_675, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_676, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_677, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_678, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_679, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_680, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_681, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_682;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_683, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_684, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_685, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_686, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_687, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_688, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_689, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_690;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_691, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_692, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_693, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_694, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_695, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_696, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_697, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_698;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_699, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_700, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_701, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_702, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_703, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_704, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_705, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_706;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_707, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_708, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_709, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_710, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_711, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_712, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_713, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_714;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_715, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_716, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_717, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_718, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_719, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_720, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_721, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_722;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_723, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_724, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_725, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_726, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_727, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_728, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_729, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_730;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_731, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_732, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_733, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_734, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_735, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_736, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_737, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_738;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_739, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_740, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_741, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_742, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_743, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_744, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_745, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_746;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_747, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_748, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_749, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_750, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_751, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_752, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_753, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_754;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_755, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_756, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_757, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_758, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_759, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_760, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_761, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_762;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_763, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_764, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_765, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_766, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_767, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_768, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_769, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_770;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_771, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_772, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_773, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_774, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_775, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_776, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_777, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_778;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_779, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_780, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_781, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_782, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_783, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_784, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_785, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_786;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_787, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_788, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_789, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_790, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_791, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_792, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_793, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_794;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_795, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_796, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_797, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_798, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_799, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_800, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_801, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_802;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_803, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_804, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_805, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_806, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_807, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_808, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_809, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_810;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_811, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_812, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_813, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_814, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_815, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_816, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_817, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_818;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_819, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_820, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_821, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_822, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_823, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_824, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_825, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_826;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_827, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_828, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_829, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_830, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_831, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_832, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_833, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_834;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_835, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_836, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_837, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_838, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_839, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_840, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_841, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_842;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_843, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_844, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_845, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_846, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_847, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_848, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_849, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_850;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_851, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_852, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_853, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_854, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_855, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_856, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_857, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_858;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_859, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_860, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_861, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_862, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_863, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_864, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_865, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_866;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_867, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_868, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_869, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_870, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_871, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_872, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_873, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_874;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_875, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_876, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_877, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_878, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_879, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_880, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_881, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_882;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_883, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_884, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_885, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_886, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_887, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_888, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_889, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_890;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_891, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_892, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_893, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_894, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_895, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_896, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_897, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_898;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_899, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_900, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_901, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_902, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_903, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_904, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_905, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_906;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_907, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_908, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_909, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_910, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_911, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_912, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_913, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_914;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_915, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_916, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_917, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_918, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_919, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_920, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_921, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_922;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_923, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_924, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_925, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_926, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_927, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_928, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_929, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_930;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_931, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_932, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_933, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_934, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_935, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_936, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_937, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_938;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_939, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_940, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_941, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_942, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_943, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_944, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_945, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_946;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_947, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_948, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_949, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_950, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_951, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_952, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_953, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_954;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_955, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_956, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_957, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_958, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_959, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_960, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_961, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_962;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_963, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_964, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_965, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_966, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_967, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_968, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_969, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_970;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_971, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_972, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_973, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_974, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_975, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_976, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_977, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_978;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_979, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_980, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_981, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_982, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_983, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_984, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_985, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_986;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_987, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_988, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_989, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_990, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_991, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_992, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_993, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_994;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_995, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_996, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_997, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_998, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_999, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1000, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1001, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1002;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1003, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1004, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1005, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1006, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1007, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1008, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1009, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1010;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1011, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1012, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1013, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1014, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1015, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1016, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1017, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1018;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1019, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1020, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1021, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1022, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1023, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1024, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1025, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1026;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1027, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1028, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1029, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1030, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1031, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1032, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1033, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1034;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1035, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1036, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1037, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1038, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1039, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1040, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1041, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1042;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1043, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1044, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1045, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1046, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1047, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1048, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1049, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1050;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1051, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1052, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1053, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1054, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1055, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1056, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1057, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1058;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1059, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1060, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1061, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1062, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1063, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1064, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1065, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1066;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1067, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1068, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1069, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1070, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1071, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1072, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1073, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1074;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1075, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1076, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1077, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1078, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1079, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1080, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1081, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1082;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1083, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1084, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1085, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1086, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1087, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1088, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1089, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1090;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1091, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1092, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1093, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1094, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1095, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1096, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1097, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1098;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1099, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1100, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1101, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1102, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1103, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1104, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1105, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1106;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1107, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1108, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1109, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1110, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1111, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1112, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1113, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1114;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1115, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1116, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1117, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1118, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1119, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1121, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1122, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1123;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1124, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1125, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1126, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1127, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1128, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1129, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1130, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1131;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1132, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1133, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1134, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1135, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1136, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1137, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1138, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1139;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1140, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1141, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1142, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1143, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1144, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1145, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1146, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1147;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1148, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1149, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1150, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1151, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1152, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1153, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1154, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1155;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1156, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1157, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1158, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1159, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1160, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1161, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1162, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1163;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1164, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1165, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1166, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1167, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1168, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1169, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1170, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1171;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1172, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1173, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1174, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1175, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1176, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1177, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1178, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1179;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1180, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1181, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1182, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1183, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1184, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1185, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1186, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1187;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1188, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1189, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1190, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1191, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1192, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1193, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1194, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1195;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1196, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1197, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1198, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1199, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1200, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1201, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1202, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1203;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1204, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1205, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1206, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1207, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1208, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1209, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1210, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1211;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1212, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1213, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1214, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1215, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1216, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1217, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1218, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1219;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1220, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1221, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1222, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1223, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1224, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1225, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1226, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1227;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1228, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1229, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1230, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1231, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1232, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1233, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1234, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1235;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1236, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1237, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1238, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1239, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1240, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1241, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1242, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1243;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1244, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1245, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1246, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1247, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1248, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1249, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1250, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1251;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1252, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1253, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1254, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1255, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1256, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1257, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1258, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1259;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1260, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1261, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1262, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1263, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1264, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1265, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1266, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1267;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1268, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1269, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1270, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1271, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1272, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1273, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1274, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1275;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1276, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1277, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1278, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1279, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1280, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1281, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1282, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1283;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1284, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1285, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1286, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1287, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1288, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1289, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1290, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1291;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1292, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1293, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1294, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1295, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1296, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1297, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1298, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1299;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1300, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1301, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1302, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1303, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1304, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1305, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1306, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1307;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1308, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1309, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1310, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1311, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1312, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1313, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1314, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1315;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1316, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1317, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1318, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1319, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1320, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1321, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1322, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1323;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1324, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1325, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1326, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1327, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1328, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1329, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1330, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1331;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1332, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1333, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1334, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1335, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1336, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1337, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1338, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1339;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1340, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1341, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1342, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1343, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1344, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1345, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1346, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1347;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1348, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1349, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1350, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1351, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1352, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1353, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1354, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1355;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1356, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1357, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1358, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1359, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1360, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1361, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1362, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1363;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1364, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1365, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1366, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1367, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1368, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1369, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1370, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1371;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1372, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1373, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1374, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1375, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1376, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1377, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1378, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1379;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1380, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1381, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1382, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1383, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1384, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1385, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1386, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1387;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1388, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1389, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1390, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1391, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1392, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1393, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1394, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1395;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1396, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1397, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1398, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1399, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1400, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1401, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1402, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1403;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1404, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1405, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1406, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1407, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1408, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1409, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1410, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1411;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1412, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1413, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1414, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1415, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1416, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1417, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1418, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1419;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1420, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1421, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1422, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1423, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1424, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1425, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1426, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1427;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1428, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1429, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1430, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1431, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1432, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1433, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1434, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1435;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1436, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1437, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1438, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1439, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1440, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1441, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1442, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1443;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1444, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1445, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1446, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1447, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1448, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1449, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1450, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1451;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1452, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1453, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1454, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1455, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1456, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1457, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1458, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1459;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1460, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1461, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1462, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1463, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1464, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1465, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1466, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1467;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1468, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1469, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1470, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1471, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1472, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1473, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1474, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1475;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1476, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1477, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1478, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1479, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1480, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1481, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1482, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1483;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1484, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1485, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1486, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1487, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1488, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1489, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1490, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1491;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1492, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1493, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1494, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1495, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1496, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1497, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1498, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1499;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1500, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1501, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1502, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1503, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1504, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1505, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1506, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1507;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1508, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1509, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1510, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1511, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1512, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1513, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1514, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1515;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1516, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1517, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1518, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1519, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1520, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1521, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1522, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1523;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1524, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1525, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1526, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1527, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1528, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1529, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1530, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1531;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1532, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1533, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1534, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1535, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1536, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1537, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1538, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1539;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1540, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1541, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1542, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1543, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1544, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1545, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1546, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1547;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1548, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1549, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1550, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1551, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1552, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1553, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1554, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1555;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1556, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1557, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1558, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1559, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1560, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1561, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1562, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1563;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1564, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1565, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1566, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1567, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1568, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1569, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1570, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1571;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1572, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1573, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1574, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1575, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1576, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1577, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1578, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1579;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1580, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1581, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1582, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1583, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1584, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1585, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1586, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1587;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1588, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1589, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1590, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1591, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1592, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1593, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1594, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1595;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1596, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1597, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1598, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1599, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1600, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1601, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1602, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1603;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1604, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1605, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1606, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1607, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1608, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1609, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1610, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1611;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1612, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1613, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1614, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1615, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1616, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1617, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1618, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1619;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1620, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1621, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1622, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1623, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1624, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1625, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1626, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1627;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1628, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1629, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1630, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1631, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1632, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1633, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1634, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1635;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1636, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1637, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1638, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1639, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1640, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1641, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1642, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1643;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1644, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1645, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1646, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1647, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1648, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1649, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1650, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1651;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1652, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1653, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1654, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1655, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1656, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1657, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1658, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1659;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1660, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1661, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1662, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1663, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1664, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1665, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1666, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1667;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1668, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1669, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1670, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1671, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1672, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1673, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1674, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1675;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1676, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1677, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1678, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1679, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1680, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1681, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1682, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1683;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1684, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1685, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1686, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1687, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1688, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1689, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1690, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1691;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1692, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1693, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1694, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1695, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1696, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1697, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1698, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1699;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1700, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1701, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1702, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1703, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1704, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1705, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1706, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1707;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1708, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1709, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1710, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1711, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1712, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1713, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1714, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1715;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1716, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1717, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1718, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1719, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1720, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1721, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1722, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1723;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1724, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1725, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1726, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1727, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1728, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1729, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1730, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1731;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1732, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1733, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1734, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1735, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1736, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1737, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1738, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1739;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1740, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1741, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1742, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1743, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1744, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1745, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1746, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1748;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1749, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1750, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1751, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1752, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1753, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1754, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1755, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1756;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1757, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1758, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1759, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1760, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1761, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1762, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1763, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1764;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1765, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1766, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1767, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1768, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1769, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1770, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1771, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1772;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1773, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1774, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1775, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1776, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1777, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1778, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1779, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1780;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1781, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1782, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1783, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1784, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1785, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1786, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1787, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1788;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1789, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1790, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1791, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1792, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1793, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1794, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1795, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1796;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1797, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1798, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1799, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1800, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1801, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1802, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1803, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1804;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1805, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1807, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1808, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1809, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1810, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1811, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1812, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1813;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1814, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1815, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1816, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1817, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1818, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1819, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1820, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1821;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1822, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1823, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1824, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1825, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1826, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1827, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1828, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1829;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1830, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1831, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1832, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1833, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1834, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1835, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1836, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1837;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1838, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1839, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1840, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1841, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1842, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1843, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1844, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1845;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1846, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1847, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1848, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1849, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1850, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1851, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1852, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1853;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1854, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1855, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1856, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1857, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1858, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1859, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1860, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1861;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1862, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1863, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1864, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1865, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1866, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1867, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1868, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1869;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1870, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1871, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1872, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1873, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1874, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1875, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1876, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1877;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1878, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1879, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1880, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1881, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1882, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1884, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1885, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1886;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1887, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1888, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1889, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1890, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1891, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1892, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1893, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1894;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1895, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1896, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1897, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1898, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1899, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1900, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1901, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1902;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1903, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1904, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1905, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1906, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1907, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1908, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1909, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1910;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1911, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1912, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1913, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1914, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1915, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1916, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1917, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1918;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1919, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1920, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1921, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1922, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1923, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1924, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1925, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1926;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1927, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1928, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1929, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1930, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1931, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1932, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1933, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1934;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1935, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1936, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1937, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1938, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1939, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1940, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1942, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1943;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1944, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1945, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1946, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1947, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1948, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1949, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1950, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1951;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1952, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1953, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1954, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1955, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1956, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1957, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1958, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1959;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1960, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1961, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1962, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1963, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1964, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1965, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1966, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1967;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1968, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1969, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1970, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1971, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1972, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1973, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1974, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1975;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1976, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1977, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1978, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1979, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1980, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1981, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1982, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1983;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1984, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1985, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1986, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1987, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1988, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1989, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1990, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1991;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1992, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1993, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1994, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1996, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1997, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1998, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1999, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2000;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2001, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2002, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2003, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2004, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2005, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2006, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2007, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2008;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2009, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2010, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2011, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2012, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2013, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2014, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2015, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2016;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2017, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2018, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2019, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2020, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2021, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2022, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2023, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2024;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2025, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2026, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2027, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2028, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2029, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2030, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2031, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2032;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2033, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2034, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2035, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2036, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2037, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2038, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2039, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2040;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2041, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2042, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2043, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2044, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2045, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2046, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2047, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2048;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2049, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2050, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2051, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2052, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2053, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2054, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2056, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2057;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2058, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2059, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2060, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2061, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2062, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2063, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2064, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2065;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2066, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2067, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2068, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2069, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2070, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2071, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2072, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2073;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2074, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2075, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2076, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2077, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2078, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2079, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2080, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2081;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2082, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2083, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2084, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2085, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2086, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2087, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2088, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2089;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2090, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2091, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2092, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2093, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2094, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2095, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2096, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2097;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2098, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2099, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2100, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2101, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2102, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2103, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2104, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2105;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2106, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2107, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2108, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2109, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2110, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2112, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2113, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2114;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2115, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2116, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2117, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2118, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2119, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2120, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2121, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2122;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2123, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2124, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2125, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2126, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2127, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2128, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2129, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2130;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2131, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2132, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2133, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2134, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2135, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2136, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2137, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2138;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2139, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2140, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2141, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2142, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2143, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2144, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2145, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2146;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2147, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2148, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2149, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2150, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2151, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2152, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2153, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2154;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2155, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2156, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2157, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2158, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2159, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2160, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2161, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2162;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2163, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2164, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2165, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2167, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2168, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2169, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2170, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2171;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2172, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2173, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2174, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2175, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2176, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2177, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2178, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2179;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2180, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2181, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2182, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2183, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2184, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2185, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2186, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2187;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2188, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2189, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2190, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2191, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2192, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2193, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2194, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2195;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2196, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2197, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2198, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2199, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2200, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2201, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2202, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2203;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2204, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2205, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2206, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2207, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2208, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2209, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2210, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2211;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2212, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2213, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2214, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2215, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2216, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2218, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2219, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2220;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2221, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2222, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2223, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2224, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2225, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2226, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2227, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2228;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2229, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2230, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2231, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2232, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2233, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2234, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2235, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2236;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2237, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2238, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2239, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2240, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2241, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2242, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2243, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2244;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2245, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2246, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2247, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2248, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2249, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2250, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2251, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2252;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2253, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2254, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2255, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2256, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2257, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2258, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2259, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2260;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2261, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2262, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2263, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2264, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2265, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2266, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2267, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2269;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2270, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2271, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2272, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2273, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2274, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2275, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2276, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2277;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2278, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2279, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2280, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2281, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2282, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2283, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2284, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2285;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2286, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2287, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2288, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2289, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2290, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2291, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2292, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2293;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2294, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2295, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2296, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2297, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2298, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2299, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2300, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2301;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2302, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2303, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2304, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2305, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2306, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2307, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2308, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2309;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2310, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2311, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2312, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2313, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2314, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2315, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2316, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2317;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2318, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2320, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2321, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2322, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2323, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2324, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2325, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2326;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2327, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2328, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2329, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2330, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2331, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2332, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2333, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2334;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2335, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2336, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2337, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2338, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2339, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2340, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2341, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2342;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2343, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2344, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2345, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2346, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2347, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2348, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2349, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2350;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2351, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2352, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2353, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2354, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2355, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2356, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2357, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2358;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2359, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2360, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2361, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2362, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2363, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2364, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2365, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2366;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2367, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2369, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2370, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2371, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2372, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2373, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2374, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2375;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2376, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2377, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2378, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2379, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2380, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2381, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2382, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2383;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2384, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2385, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2386, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2387, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2388, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2389, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2390, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2391;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2392, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2393, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2394, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2395, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2396, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2397, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2398, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2399;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2400, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2401, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2402, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2403, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2404, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2405, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2406, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2407;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2408, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2409, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2410, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2411, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2412, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2413, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2414, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2415;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2416, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2417, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2418, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2419, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2420, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2421, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2422, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2423;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2424, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2425, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2426, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2427, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2428, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2429, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2430, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2431;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2432, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2433, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2434, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2435, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2436, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2437, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2438, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2439;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2440, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2441, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2442, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2443, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2444, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2445, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2446, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2447;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2448, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2449, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2450, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2451, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2452, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2453, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2454, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2455;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2456, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2457, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2458, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2459, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2460, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2461, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2462, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2463;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2464, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2465, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2466, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2467, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2468, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2469, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2470, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2471;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2472, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2473, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2474, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2475, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2476, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2477, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2478, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2479;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2480, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2481, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2482, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2483, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2484, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2485, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2486, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2487;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2488, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2489, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2490, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2491, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2492, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2493, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2494, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2495;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2496, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2497, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2498, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2500, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2501, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2502, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2503, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2504;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2505, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2506, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2507, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2508, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2509, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2510, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2511, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2512;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2513, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2514, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2515, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2516, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2517, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2518, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2519, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2520;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2521, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2522, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2523, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2524, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2525, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2526, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2527, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2528;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2529, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2530, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2531, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2532, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2533, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2534, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2535, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2536;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2537, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2538, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2539, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2540, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2541, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2542, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2543, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2544;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2545, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2546, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2547, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2548, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2549, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2550, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2551, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2552;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2553, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2554, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2556, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2557, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2558, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2559, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2560, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2561;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2562, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2563, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2564, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2565, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2566, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2567, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2568, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2569;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2570, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2571, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2572, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2573, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2574, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2575, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2576, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2577;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2578, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2579, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2580, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2581, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2582, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2583, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2584, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2585;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2586, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2587, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2588, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2589, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2590, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2591, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2592, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2593;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2594, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2595, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2596, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2597, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2598, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2599, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2600, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2601;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2602, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2603, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2604, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2605, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2606, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2607, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2609, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2610;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2611, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2612, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2613, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2615, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2616, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2617, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2619, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2620;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2621, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2622, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2623, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2624, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2626, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2627, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2629, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2630;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2632, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2633, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2635, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2636, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2637, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2639, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2640, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2642;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2643, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2645, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2646, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2647, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2649, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2650, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2652, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2653;
  wire mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2655, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2656, mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2658, n_0, n_1, n_2, n_3, n_4;
  wire n_5, n_6, n_7, n_8, n_9, n_10, n_11, n_12;
  wire n_13, n_14, n_15, n_16, n_17, n_18, n_19, n_20;
  wire n_21, n_22, n_23, n_24, n_25, n_26, n_27, n_28;
  wire n_29, n_30, n_31, n_32, n_33, n_34, n_35, n_36;
  wire n_37, n_38, n_39, n_40, n_41, n_42, n_43, n_44;
  wire n_45, n_46, n_47, n_48, n_49, n_50, n_51, n_52;
  wire n_53, n_54, n_55, n_56, n_57, n_58, n_59, n_60;
  wire n_61, n_62, n_63, n_64, n_65, n_66, n_67, n_68;
  wire n_69, n_70, n_71, n_72, n_73, n_74, n_75, n_76;
  wire n_77, n_78, n_79, n_80, n_81, n_82, n_83, n_84;
  wire n_85, n_86, n_87, n_88, n_89, n_90, n_91, n_92;
  wire n_93, n_94, n_95, n_96, n_97, n_98, n_99, n_100;
  wire n_103, n_104, n_105, n_106, n_107, n_108, n_109, n_110;
  wire n_111, n_112, n_113, n_114, n_115, n_116, n_117, n_118;
  wire n_119, n_120, n_121, n_122, n_123, n_124, n_125, n_126;
  wire n_127, n_128, n_129, n_130, n_131, n_132, n_133, n_134;
  wire n_135, n_136, n_137, n_138, n_139, n_140, n_141, n_142;
  wire n_143, n_144, n_145, n_146, n_147, n_148, n_149, n_150;
  wire n_151, n_152, n_153, n_154, n_155, n_174, n_175, n_176;
  wire n_177, n_178, n_179, n_180, n_181, n_182, n_183, n_184;
  wire n_185, n_186, n_187, n_188, n_189, n_190, n_191, n_192;
  wire n_193, n_194, n_195, n_196, n_197, n_198, n_199, n_200;
  wire n_201, n_202, n_203, n_204, n_205;
  or g719__2398(n_192 ,n_119 ,n_136);
  or g720__5107(n_204 ,n_111 ,n_131);
  or g721__6260(n_203 ,n_120 ,n_137);
  or g722__4319(n_193 ,n_121 ,n_138);
  or g723__8428(n_205 ,n_116 ,n_129);
  or g724__5526(n_199 ,n_118 ,n_135);
  or g725__6783(n_191 ,n_134 ,n_133);
  or g726__3680(n_202 ,n_113 ,n_127);
  or g727__1617(n_196 ,n_110 ,n_126);
  or g728__2802(n_190 ,n_140 ,n_123);
  or g729__1705(n_197 ,n_112 ,n_128);
  or g730__5122(n_201 ,n_109 ,n_125);
  or g731__8246(n_198 ,n_115 ,n_130);
  or g732__7098(n_200 ,n_122 ,n_132);
  or g733__6131(n_195 ,n_108 ,n_124);
  or g734__1881(n_194 ,n_107 ,n_139);
  and g735__5115(n_140 ,in3[0] ,n_33);
  and g736__7482(n_139 ,in3[4] ,n_24);
  and g737__4733(n_138 ,in3[3] ,n_34);
  and g738__6161(n_137 ,in3[13] ,n_21);
  and g739__9315(n_136 ,in3[2] ,n_22);
  and g740__9945(n_135 ,in3[9] ,n_33);
  and g741__2883(n_134 ,in3[1] ,n_34);
  and g743__2346(n_132 ,in3[10] ,n_31);
  and g744__1666(n_131 ,in3[14] ,n_30);
  and g745__7410(n_130 ,in3[8] ,n_30);
  and g746__6417(n_129 ,in3[15] ,n_21);
  and g747__5477(n_128 ,in3[7] ,n_31);
  and g748__2398(n_127 ,in3[12] ,n_25);
  and g749__5107(n_126 ,in3[6] ,n_25);
  and g750__6260(n_125 ,in3[11] ,n_24);
  and g751__4319(n_124 ,in3[5] ,n_22);
  and g753__8428(n_122 ,in2[10] ,n_54);
  and g754__5526(n_121 ,in2[3] ,n_48);
  and g755__6783(n_120 ,in2[13] ,n_51);
  and g756__3680(n_119 ,in2[2] ,n_53);
  and g757__1617(n_118 ,in2[9] ,n_53);
  and g758__2802(n_117 ,in2[1] ,n_45);
  and g759__1705(n_116 ,in2[15] ,n_47);
  and g760__5122(n_115 ,in2[8] ,n_48);
  and g761__8246(n_114 ,in2[0] ,n_50);
  and g762__7098(n_113 ,in2[12] ,n_44);
  and g763__6131(n_112 ,in2[7] ,n_54);
  and g764__1881(n_111 ,in2[14] ,n_51);
  and g765__5115(n_110 ,in2[6] ,n_50);
  and g766__7482(n_109 ,in2[11] ,n_47);
  and g767__4733(n_108 ,in2[5] ,n_44);
  and g768__6161(n_107 ,in2[4] ,n_45);
  or g769__9315(n_179 ,n_82 ,n_97);
  or g770__9945(n_188 ,n_69 ,n_90);
  or g771__2883(n_105 ,n_66 ,n_98);
  or g772__2346(n_177 ,n_77 ,n_95);
  or g773__1666(n_176 ,n_76 ,n_94);
  or g774__7410(n_104 ,n_70 ,n_93);
  or g775__6417(n_103 ,n_73 ,n_92);
  or g778__5477(n_189 ,n_71 ,n_91);
  or g779__2398(n_178 ,n_75 ,n_96);
  or g780__5107(n_187 ,n_68 ,n_89);
  or g781__6260(n_100 ,n_67 ,n_88);
  or g782__4319(n_185 ,n_63 ,n_87);
  or g783__8428(n_184 ,n_65 ,n_86);
  or g784__5526(n_99 ,n_64 ,n_85);
  or g785__6783(n_182 ,n_72 ,n_84);
  or g786__3680(n_181 ,n_74 ,n_83);
  and g787__1617(n_106 ,n_78 ,n_81);
  and g788__2802(n_98 ,in2[6] ,n_19);
  and g789__1705(n_97 ,in2[5] ,n_28);
  and g790__5122(n_96 ,in2[4] ,n_42);
  and g791__8246(n_95 ,in2[3] ,n_39);
  and g792__7098(n_94 ,in2[2] ,n_41);
  and g793__6131(n_93 ,in2[1] ,n_27);
  and g794__1881(n_92 ,in2[0] ,n_36);
  and g795__5115(n_91 ,in2[15] ,n_17);
  and g796__7482(n_90 ,in2[14] ,n_17);
  and g797__4733(n_89 ,in2[13] ,n_28);
  and g798__6161(n_88 ,in2[12] ,n_36);
  and g799__9315(n_87 ,in2[11] ,n_39);
  and g800__9945(n_86 ,in2[10] ,n_41);
  and g801__2883(n_85 ,in2[9] ,n_27);
  and g802__2346(n_84 ,in2[8] ,n_37);
  and g803__1666(n_83 ,in2[7] ,n_16);
  and g804__7410(n_82 ,in1[5] ,in4[1]);
  not g806(n_80 ,n_78);
  not g807(n_79 ,n_78);
  and g808__6417(n_77 ,in1[3] ,in4[1]);
  and g809__5477(n_76 ,in1[2] ,in4[1]);
  and g810__2398(n_75 ,in1[4] ,in4[1]);
  and g811__5107(n_74 ,in1[7] ,in4[1]);
  and g812__6260(n_73 ,in1[0] ,in4[1]);
  and g813__4319(n_72 ,in1[8] ,in4[1]);
  and g814__8428(n_71 ,in1[15] ,in4[1]);
  and g815__5526(n_70 ,in1[1] ,in4[1]);
  and g816__6783(n_69 ,in1[14] ,in4[1]);
  and g817__3680(n_68 ,in1[13] ,in4[1]);
  and g818__1617(n_67 ,in1[12] ,in4[1]);
  and g819__2802(n_66 ,in1[6] ,in4[1]);
  and g820__1705(n_65 ,in1[10] ,in4[1]);
  and g821__5122(n_64 ,in1[9] ,in4[1]);
  and g822__8246(n_63 ,in1[11] ,in4[1]);
  or g823__7098(n_81 ,in4[1] ,in4[0]);
  or g824__6131(n_78 ,n_19 ,n_62);
  not g825(n_62 ,in4[0]);
  not g826(n_61 ,in4[1]);
  not drc_bufs851(n_141 ,n_60);
  not drc_bufs852(n_60 ,n_81);
  buf drc_bufs855(n_186 ,n_100);
  buf drc_bufs856(n_180 ,n_105);
  buf drc_bufs857(n_183 ,n_99);
  buf drc_bufs858(n_175 ,n_104);
  buf drc_bufs859(n_174 ,n_103);
  not drc_bufs865(n_59 ,n_57);
  not drc_bufs866(n_58 ,n_57);
  not drc_bufs867(n_57 ,n_61);
  not drc_bufs875(n_56 ,n_55);
  not drc_bufs877(n_55 ,n_106);
  not drc_bufs880(n_54 ,n_52);
  not drc_bufs881(n_53 ,n_52);
  not drc_bufs882(n_52 ,n_79);
  not drc_bufs884(n_51 ,n_49);
  not drc_bufs885(n_50 ,n_49);
  not drc_bufs886(n_49 ,n_79);
  not drc_bufs888(n_48 ,n_46);
  not drc_bufs889(n_47 ,n_46);
  not drc_bufs890(n_46 ,n_80);
  not drc_bufs892(n_45 ,n_43);
  not drc_bufs893(n_44 ,n_43);
  not drc_bufs894(n_43 ,n_80);
  not drc_bufs900(n_42 ,n_40);
  not drc_bufs901(n_41 ,n_40);
  not drc_bufs902(n_40 ,n_61);
  not drc_bufs905(n_39 ,n_38);
  not drc_bufs906(n_38 ,n_59);
  not drc_bufs908(n_37 ,n_35);
  not drc_bufs909(n_36 ,n_35);
  not drc_bufs910(n_35 ,n_61);
  not drc_bufs912(n_34 ,n_32);
  not drc_bufs913(n_33 ,n_32);
  not drc_bufs914(n_32 ,n_106);
  not drc_bufs916(n_31 ,n_29);
  not drc_bufs917(n_30 ,n_29);
  not drc_bufs918(n_29 ,n_106);
  not drc_bufs920(n_28 ,n_26);
  not drc_bufs921(n_27 ,n_26);
  not drc_bufs922(n_26 ,n_58);
  not drc_bufs924(n_25 ,n_23);
  not drc_bufs925(n_24 ,n_23);
  not drc_bufs926(n_23 ,n_56);
  not drc_bufs928(n_22 ,n_20);
  not drc_bufs929(n_21 ,n_20);
  not drc_bufs930(n_20 ,n_56);
  not drc_bufs932(n_19 ,n_18);
  not drc_bufs934(n_18 ,n_42);
  not drc_bufs936(n_17 ,n_15);
  not drc_bufs937(n_16 ,n_15);
  not drc_bufs938(n_15 ,n_59);
  and g428__1881(out1[22] ,n_146 ,n_11);
  and g429__5115(out1[30] ,n_154 ,n_10);
  and g430__7482(out1[28] ,n_152 ,n_5);
  and g431__4733(out1[24] ,n_148 ,n_2);
  and g432__6161(out1[23] ,n_147 ,n_8);
  and g433__9315(out1[27] ,n_151 ,n_11);
  and g434__9945(out1[31] ,n_155 ,n_4);
  and g435__2883(out1[18] ,n_142 ,n_1);
  and g436__2346(out1[29] ,n_153 ,n_7);
  and g437__1666(out1[26] ,n_150 ,n_10);
  and g438__7410(out1[20] ,n_144 ,n_5);
  and g439__6417(out1[19] ,n_143 ,n_2);
  and g440__5477(out1[25] ,n_149 ,n_7);
  and g441__2398(out1[21] ,n_145 ,n_8);
  not drc_bufs(n_14 ,n_12);
  not drc_bufs442(n_13 ,n_12);
  not drc_bufs443(n_12 ,n_141);
  not drc_bufs456(n_11 ,n_9);
  not drc_bufs457(n_10 ,n_9);
  not drc_bufs458(n_9 ,n_14);
  not drc_bufs460(n_8 ,n_6);
  not drc_bufs461(n_7 ,n_6);
  not drc_bufs462(n_6 ,n_13);
  not drc_bufs464(n_5 ,n_3);
  not drc_bufs465(n_4 ,n_3);
  not drc_bufs466(n_3 ,n_13);
  not drc_bufs468(n_2 ,n_0);
  not drc_bufs469(n_1 ,n_0);
  not drc_bufs470(n_0 ,n_14);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4560__5107(n_155 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2658 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1744);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4561__6260(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2658 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2523 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2656);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4562__4319(n_154 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2655 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2553);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4563__8428(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2656 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2521 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2655);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4564__5526(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2655 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2574 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2653);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4565__6783(n_153 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2652 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2582);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4566__3680(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2653 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2577 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2652);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4567__1617(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2652 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2576 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2650);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4568__2802(n_152 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2649 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2585);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4569__1705(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2650 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2575 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2649);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4570__5122(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2649 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2602 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2647);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4571__8246(n_151 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2645 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2607);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4572__7098(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2647 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2600 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2646);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4573(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2646 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2645);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4574__6131(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2645 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2599 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2643);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4575__1881(n_150 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2642 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2606);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4576__5115(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2643 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2598 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2642);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4577__7482(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2642 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2572 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2640);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4578__4733(n_149 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2639 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2586);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4579__6161(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2640 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2639 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2571);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4580__9315(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2639 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2596 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2637);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4581__9945(n_148 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2635 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2605);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4582__2883(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2637 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2597 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2636);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4583(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2636 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2635);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4584__2346(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2635 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2601 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2633);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4585__1666(n_147 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2632 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2604);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4586__7410(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2633 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2632 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2595);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4587__6417(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2632 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2580 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2630);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4588__5477(n_146 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2629 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2584);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4589__2398(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2630 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2573 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2629);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4590__5107(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2629 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2587 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2627);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4591__6260(n_145 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2626 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2611);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4592__4319(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2627 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2626 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2590);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4593__8428(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2626 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2594 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2624);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4594__5526(n_144 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2623 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2612);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4595__6783(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2624 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2623 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2593);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4596__3680(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2623 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2579 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2622);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4598__1617(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2622 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2578 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2621);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4600__2802(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2621 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2589 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2620);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4602__1705(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2620 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2588 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2619);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4604__5122(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2619 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2617 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2591);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4605__8246(out1[17] ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2615 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2609);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4606__7098(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2617 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2616 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2592);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4607(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2616 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2615);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4608__6131(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2615 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2570 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2613);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4609__1881(out1[16] ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2603 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2583);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4610__5115(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2613 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2603 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2556);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4611__7482(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2612 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2545 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2558);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4612__4733(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2611 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2532 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2566);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4613__6161(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2610 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2534 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2568);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4614__9315(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2609 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2539 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2562);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4615__9945(out1[15] ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2535 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2554);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4616__2883(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2607 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2559 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2537);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4617__2346(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2606 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2552 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2563);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4618__1666(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2605 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2560 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2536);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4619__7410(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2604 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2546 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2564);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4620__6417(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2602 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2537 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2559);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4621__5477(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2601 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2546 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2564);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4622__2398(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2600 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2537 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2559);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4623__5107(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2599 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2552 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2563);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4624__6260(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2598 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2552 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2563);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4625__4319(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2597 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2536 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2560);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4626__8428(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2596 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2536 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2560);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4627__5526(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2595 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2546 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2564);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4628__6783(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2594 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2544 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2558);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4629__3680(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2593 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2545 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2557);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4630__1617(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2603 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2522 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2569);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4631__2802(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2592 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2539 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2562);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4632__1705(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2591 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2538 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2561);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4633__5122(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2590 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2532 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2565);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4634__8246(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2589 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2533 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2567);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4635__7098(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2588 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2534 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2568);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4636__6131(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2587 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2531 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2566);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4637__1881(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2586 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2540 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2525);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4638__5115(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2585 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2526 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2550);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4639__7482(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2584 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2542 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2527);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4640__4733(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2583 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2517 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2528);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4641__6161(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2582 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2549 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2502);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4642__9315(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2581 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2530 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2548);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4643__9945(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2580 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2543 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2527);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4644__2883(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2579 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2529 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2547);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4645__2346(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2578 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2530 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2548);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4646__1666(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2577 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2549 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2502);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4647__7410(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2576 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2526 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2551);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4648__6417(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2575 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2526 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2551);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4649__5477(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2574 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2549 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2502);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4650__2398(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2573 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2543 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2527);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4651__5107(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2572 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2541 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2525);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4652__6260(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2571 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2541 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2525);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4653__4319(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2570 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2518 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2528);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4654__8428(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2569 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2535 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2524);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4655(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2568 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2567);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4656(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2566 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2565);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4657(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2562 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2561);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4658(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2557 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2558);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4659__5526(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2556 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2518 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2528);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4660__6783(out1[14] ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2472 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2494);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4661__3680(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2554 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2450 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2504);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4662__1617(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2553 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2520 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1716);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4663__2802(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2567 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2464 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2492);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4664__1705(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2565 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2463 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2490);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4665__5122(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2564 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2436 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2497);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4666__8246(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2563 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_23 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2496);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4667__7098(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2561 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2439 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2491);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4668__6131(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2560 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2462 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2493);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4669__1881(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2559 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2461 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2498);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4670__5115(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2558 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2437 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2495);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4671(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2551 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2550);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4672(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2547 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2548);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4673(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2544 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2545);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4674(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2543 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2542);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4675(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2541 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2540);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4676(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2538 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2539);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4677__7482(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2552 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2427 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2509);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4678__4733(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2550 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2487 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2514);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4679__6161(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2549 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1733 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2513);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4680__9315(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2548 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2483 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2512);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4681__9945(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2546 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2419 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2511);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4682__2883(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2545 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2430 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2515);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4683__2346(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2542 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2479 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2510);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4684__1666(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2540 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2471 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2508);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4685__7410(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2539 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2414 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2507);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4686__6417(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2537 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2485 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2506);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4687__5477(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2536 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2468 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2505);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4688(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2534 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2533);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4689(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2531 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2532);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4690(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2529 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2530);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4691__2398(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2524 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2450 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2503);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4692__5107(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2523 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1716 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2520);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4693__6260(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2522 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2449 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2504);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4694__4319(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2521 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1715 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2519);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4695__8428(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2535 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2516 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2465);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4696__5526(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2533 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2481 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2501);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4697__6783(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2532 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2477 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2500);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4698__3680(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2530 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2476 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2432);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4699__1617(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2528 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2473 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2431);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4700__2802(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2527 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2475 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2434);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4701__1705(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2526 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_9 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1746);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4702__5122(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2525 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2474 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2447);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4703(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2519 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2520);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4704(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2518 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2517);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4705__8246(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2516 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2472 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2466);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4706__7098(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2515 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2476 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2428);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4707__6131(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2514 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2461 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2486);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4708__1881(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2513 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1734 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_9);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4709__5115(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2512 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2482 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2464);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4710__7482(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2511 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2475 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2417);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4711__4733(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2510 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2463 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2478);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4712__6161(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2509 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2474 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2426);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4713__9315(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2508 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2462 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2470);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4714__9945(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2507 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2473 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2413);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4715__2883(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2506 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2488 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2444);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4716__2346(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2505 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2484 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2443);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4717__1666(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2520 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1603 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2489);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4718__7410(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2517 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2343 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2467);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4719(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2504 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2503);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4720__6417(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2501 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2446 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2480);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4721__5477(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2500 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2469 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2460);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4722__2398(out1[13] ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2353 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2433);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4723__5107(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2498 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1720 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2452);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4724__6260(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2497 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2406 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2443);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4725__4319(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2496 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2404 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2444);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4726__8428(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2495 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2401 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2459);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4727__5526(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2494 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2442 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2408);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4728__6783(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2493 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2454 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2376);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4729__3680(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2492 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2457 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2322);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4730__1617(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2491 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2445 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2410);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4731__2802(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2490 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2455 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2374);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4732__1705(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2503 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2458 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2367);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4733__5122(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2502 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_21 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1620);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4734__8246(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2489 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1591 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_21);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4735__7098(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2488 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2440 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2404);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4736__6131(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2487 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1720 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2451);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4737__1881(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2486 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1719 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2452);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4738__5115(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2485 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_23 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2403);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4739__7482(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2484 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2435 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2406);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4740__4733(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2483 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2456 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2322);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4741__6161(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2482 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2457 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2321);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4742__9315(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2481 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2439 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2409);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4743__9945(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2480 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2438 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2410);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4744__2883(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2479 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2455 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2374);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4745__2346(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2478 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2455 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2374);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4746__1666(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2477 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2437 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2402);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4747__7410(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2471 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2453 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2376);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4748__6417(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2470 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2454 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2375);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4749__5477(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2469 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2437 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2402);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4750__2398(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2468 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2436 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2405);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4751__5107(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2467 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2458 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2350);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4752__6260(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2466 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2441 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2408);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4753__4319(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2465 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2442 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2407);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4755__8428(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2476 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_164 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2424);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4756__5526(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2475 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_183 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2422);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4757__6783(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2474 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_172 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2425);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4758__3680(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2473 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_237 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2421);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4759__1617(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2472 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2448 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2411);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4760(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2460 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2459);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4761(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2456 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2457);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4762(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2453 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2454);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4763(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2451 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2452);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4764(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2449 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2450);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4765__2802(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2448 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2354 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2412);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4766__1705(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2447 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2378 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2364);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4767__5122(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2464 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2249 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2418);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4768__8246(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2463 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2310 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2429);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4769__7098(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2462 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2305 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2415);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4770__6131(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2461 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1497 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2420);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4771__1881(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2459 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2384 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2313);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4772__5115(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2458 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_226 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2397);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4773__7482(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2457 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_176 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2394);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4774__4733(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2455 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_154 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2398);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4775__6161(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2454 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_172 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2395);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4776__9315(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2452 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_184 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2396);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4777__9945(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2450 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2247 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2416);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4778(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2446 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2445);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4779(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2442 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2441);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4780(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2440 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_23);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4781(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2438 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2439);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4782(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2435 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2436);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4783__2883(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2434 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2366 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2380);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4784__2346(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2433 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2382 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2201);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4785__1666(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2432 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2383 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2342);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4786__7410(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2431 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2341 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2373);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4787__6417(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2445 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2385 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2266);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4788__5477(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2444 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2386 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1622);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4789__2398(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2443 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2388 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2316);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4791__5107(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2441 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2387 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2267);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4793__6260(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2439 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_752 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2389);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4794__4319(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2437 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2392 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_759);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4795__8428(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2436 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2391 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_757);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4796__5526(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2430 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2383 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2342);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4797__6783(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2429 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2384 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2308);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4798__3680(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2428 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2383 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2342);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4799__1617(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2427 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2378 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2363);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4800__2802(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2426 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2377 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2364);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4801__1705(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2425 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1653 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2369);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4802__5122(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2424 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1675 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2399);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4803__8246(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2423 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1664 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2370);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4804__7098(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2422 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1678 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2371);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4805__6131(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2421 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1452 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2400);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4806__1881(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2420 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1496 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2386);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4807__5115(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2419 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2365 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2380);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4808__7482(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2418 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2385 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2248);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4809__4733(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2417 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2366 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2379);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4810__6161(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2416 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2387 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2246);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4811__9315(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2415 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2388 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2299);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4812__9945(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2414 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2340 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2373);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4813__2883(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2413 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2341 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2372);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4814__2346(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2412 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2382 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2201);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4815__1666(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2411 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2381 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2200);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4816(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2409 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2410);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4817(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2407 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2408);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4818(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2405 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2406);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4819(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2403 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2404);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4820(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2402 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2401);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4821__7410(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2400 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_586 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_653);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4822__6417(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2399 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_592 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2352);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4823__5477(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2398 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1656 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2361);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4824__2398(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2397 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1457 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2349);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4825__5107(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2396 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1658 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2359);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4826__6260(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2395 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1668 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2360);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4827__4319(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2394 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1600 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2362);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4828__8428(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2393 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1564 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2351);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4829__5526(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2392 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1562 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2347);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4830__6783(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2391 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1563 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2344);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4831__3680(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2390 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1568 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2345);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4832__1617(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2389 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1266 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2348);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4833__2802(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2410 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2203 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2356);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4834__1705(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2408 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2196 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2346);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4835__5122(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2406 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2250 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2355);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4836__8246(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2404 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1710 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2357);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4837__7098(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2401 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2258 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2358);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4838(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2382 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2381);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4839(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2379 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2380);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4840(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2377 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2378);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4841(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2375 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2376);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4842(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2373 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2372);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4843__6131(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2371 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_589 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_653);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4844__1881(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2370 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_583 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2352);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4845__5115(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2369 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_580 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_652);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4846__7482(out1[12] ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2301 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2315);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4847__4733(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2367 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2148 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2323);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4848__6161(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2388 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_152 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2331);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4849__9315(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2387 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_150 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2329);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4850__9945(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2386 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_168 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2328);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4851__2883(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2385 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_179 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2327);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4852__2346(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2384 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_183 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2330);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4853__1666(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2383 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_5 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2265);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4854__7410(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2381 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2325 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2213);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4855__6417(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2380 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2324 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2263);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4856__5477(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2378 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2326 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1745);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4857__2398(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2376 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2291 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2314);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4858__5107(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2374 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2290 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2317);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4859__6260(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2372 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_7 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2214);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4860(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2365 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2366);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4861(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2363 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2364);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4862__4319(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2362 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1553 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2335);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4863__8428(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2361 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1449 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2337);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4864__5526(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2360 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1442 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2320);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4865__6783(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2359 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1432 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2318);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4866__3680(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2358 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_5 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2257);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4867__1617(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2357 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1732 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2326);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4868__2802(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2356 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_7 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2204);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4869__1705(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2355 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2324 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2253);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4870__5122(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2366 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2297 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2332);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4871__8246(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2364 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2303 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2338);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4872(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2354 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2353);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4873__7098(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2351 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_406 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2339);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4874__6131(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2350 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2148 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2323);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4875__1881(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2349 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1458 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2336);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4876__5115(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2348 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_394 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_658);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4877__7482(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2347 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_409 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_657);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4878__4733(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2346 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2325 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2198);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4879__6161(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2345 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_397 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_668);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4880__9315(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2344 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_400 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_658);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4881__9945(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2343 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2148 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2323);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4882__2883(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2353 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2294 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2334);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4883__2346(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2352 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1066 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2333);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4884(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2340 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2341);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4886__1666(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2338 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2291 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2302);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4887__7410(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2337 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_399 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_686);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4888__6417(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2336 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_393 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2300);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4889__5477(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2335 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_408 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_686);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4890__2398(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2334 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2293 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2301);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4891__5107(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2333 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_975 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2312);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4892__6260(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2332 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2290 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2296);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4893__4319(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2331 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1637 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2306);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4894__8428(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2330 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1645 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2309);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4895__5526(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2329 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1435 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2292);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4896__6783(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2328 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1681 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2307);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4897__3680(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2327 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1667 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2304);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4898__1617(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2342 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2197 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2298);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4899__2802(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2341 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2144 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2295);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4900__1705(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2339 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_36 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2311);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4901(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2322 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2321);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4902__5122(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2320 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_396 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2300);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4903__8246(out1[11] ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2252 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2264);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4904__7098(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2318 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_405 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_685);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4905__6131(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2317 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2274 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2222);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4906__1881(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2316 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2242 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2273);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4907__5115(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2315 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2270 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2220);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4908__7482(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2314 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1718 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2276);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4909__4733(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2313 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2240 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2271);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4910__6161(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2326 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_229 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2283);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4912__9315(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2325 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_148 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2282);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4914__9945(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2324 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_185 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2279);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4915__2883(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2323 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2278 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2161);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4916__2346(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2321 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2277 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2216);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4917(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2312 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2311);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4918__1666(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2310 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2240 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2271);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4919__7410(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2309 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1404 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2287);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4920__6417(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2308 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2240 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2271);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4921__5477(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2307 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1406 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2288);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4922__2398(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2306 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1424 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2269);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4923__5107(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2305 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2241 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2273);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4924__6260(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2304 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1331 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2285);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4925__4319(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2303 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1718 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2275);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4926__8428(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2302 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1717 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2276);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4927__5526(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2311 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1115 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2289);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4928__6783(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2299 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2242 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2272);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4929__3680(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2298 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2277 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2192);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4930__1617(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2297 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2274 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2222);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4931__2802(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2296 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2274 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2222);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4932__1705(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2295 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2278 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2143);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4933__5122(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2294 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2270 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2220);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4934__8246(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2293 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2270 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2220);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4935__7098(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2292 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1329 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2286);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4936__6131(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2301 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2244 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2284);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4937__1881(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2300 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2262 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1164);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4938__5115(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2289 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1134 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2262);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4939__7482(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2288 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_405 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_692);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4940__4733(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2287 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_399 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2251);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4941__6161(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2286 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_393 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_692);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4942__9315(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2285 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_408 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2251);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4943__9945(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2284 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2252 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2245);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4944__2883(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2283 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1676 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2261);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4945__2346(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2282 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1467 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2243);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4946__1666(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2281 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1599 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2254);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4947__7410(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2280 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1663 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2256);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4948__6417(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2279 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1677 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2255);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4949__5477(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2291 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1499 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2259);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4950__2398(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2290 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2155 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2260);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4951(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2275 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2276);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4952(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2272 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2273);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4953__5107(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2269 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_396 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_691);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4954__6260(out1[10] ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2202 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2215);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4955__4319(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2267 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2223 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2171);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4956__8428(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2266 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2218 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2170);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4957__5526(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2265 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2221 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2191);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4958__6783(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2264 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2219 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_30);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4959__3680(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2263 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2224 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2211);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4960__1617(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2278 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_203 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2230);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4961__2802(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2277 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_195 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2232);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4962__1705(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2276 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_168 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2228);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4963__5122(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2274 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_199 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2229);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4964__8246(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2273 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2227 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1621);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4965__7098(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2271 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2226 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2163);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4966__6131(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2270 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_238 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2231);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4967__1881(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2261 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1414 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2237);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4968__5115(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2260 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2226 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2153);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4969__7482(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2259 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1498 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2227);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4970__4733(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2258 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2221 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2191);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4971__6161(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2257 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2221 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2191);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4972__9315(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2256 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1330 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2234);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4973__9945(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2255 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1376 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2236);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4974__2883(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2254 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1554 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2239);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4975__2346(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2253 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2225 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2211);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4976__1666(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2262 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1121 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2238);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4977__7410(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2250 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2225 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2211);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4978__6417(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2249 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2218 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2170);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4979__5477(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2248 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2218 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2170);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4980__2398(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2247 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2223 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2171);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4981__5107(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2246 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2223 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2171);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4982__6260(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2245 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2219 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_30);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4983__4319(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2244 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2219 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_30);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4984__8428(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2243 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1345 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2235);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4985__5526(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2252 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2195 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2233);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4986__6783(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2251 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2212 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1161);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4987(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2241 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2242);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4988__3680(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2239 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_588 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_689);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4989__1617(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2238 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1116 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2212);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4990__2802(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2237 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_582 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2199);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4991__1705(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2236 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_579 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_689);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4992__5122(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2235 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_585 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2199);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4993__8246(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2234 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_591 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_688);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4994__7098(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2233 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2194 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2202);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4995__6131(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2232 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1605 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2205);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4996__1881(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2231 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1464 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2193);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4997__5115(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2230 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1651 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2210);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4998__7482(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2229 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1670 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2206);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g4999__4733(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2228 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1659 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2209);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5000__6161(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2242 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1683 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2207);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5001__9315(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2240 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2099 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2208);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5002(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2225 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2224);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5003__9945(out1[9] ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2160 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2165);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5004__2883(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2216 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2169 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2158);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5005__2346(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2215 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2173 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_29);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5006__1666(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2214 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2172 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2122);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5007__7410(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2213 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2168 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2119);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5008__6417(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2227 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_170 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2178);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5009__5477(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2226 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_197 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2177);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5010__2398(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2224 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2175 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1708);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5011__5107(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2223 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_178 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2181);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5012__6260(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2222 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2138 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2164);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5013__4319(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2221 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2176 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2106);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5014__8428(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2220 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2149 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2162);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5015__5526(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2219 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_225 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2180);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5016__6783(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2218 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_174 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2179);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5017__3680(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2210 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1377 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2184);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5018__1617(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2209 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1412 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2190);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5019__2802(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2208 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2176 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2098);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5020__1705(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2207 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1686 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2175);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5021__5122(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2206 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1399 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2188);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5022__8246(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2205 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1611 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2187);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5023__7098(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2204 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2172 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2122);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5024__6131(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2203 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2172 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2122);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5025__1881(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2212 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1103 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2189);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5026__5115(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2211 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2156 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2185);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5027(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2201 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2200);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5028__7482(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2198 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2168 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2118);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5029__4733(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2197 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2169 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2158);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5030__6161(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2196 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2167 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2119);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5031__9315(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2195 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2174 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_29);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5032__9945(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2194 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2174 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_29);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5033__2883(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2193 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1360 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2186);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5034__2346(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2192 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2169 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2158);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5035__1666(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2202 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2139 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2182);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5036__7410(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2200 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2140 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2183);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5037__6417(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2199 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2159 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1157);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5038__5477(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2190 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_402 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_680);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5039__2398(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2189 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1142 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2159);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5040__5107(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2188 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_411 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2147);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5041__6260(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2187 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_384 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_680);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5042__4319(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2186 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_390 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2147);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5043__8428(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2185 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2138 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2150);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5044__5526(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2184 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_387 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_679);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5045__6783(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2183 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2141 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2149);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5046__3680(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2182 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2142 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2160);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5047__1617(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2181 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1615 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2151);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5048__2802(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2180 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1455 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2145);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5049__1705(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2179 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1669 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2152);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5050__5122(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2178 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1652 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2157);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5051__8246(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2177 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1661 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2154);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5052__7098(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2191 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2029 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2146);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5053(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2174 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2173);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5054(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2167 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2168);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5055__6131(out1[8] ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2104 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2110);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5056__1881(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2165 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2114 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2063);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5057__5115(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2164 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1646 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2120);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5058__7482(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2163 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2082 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2121);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5059__4733(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2162 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2117 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2060);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5060__6161(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2161 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2115 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2061);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5061__9315(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2176 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_211 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2126);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5062__9945(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2175 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_228 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2124);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5063__2883(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2173 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_754 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2128);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5064__2346(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2172 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_201 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2125);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5065__1666(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2171 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2092 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2108);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5066__7410(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2170 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2091 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2107);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5068__6417(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2169 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2123 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2051);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5069__5477(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2168 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_181 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2127);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5070__2398(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2157 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1410 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2112);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5071__5107(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2156 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1646 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2120);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5072__6260(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2155 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2082 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2121);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5073__4319(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2154 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1411 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2135);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5074__8428(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2153 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2082 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2121);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5075__5526(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2152 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1422 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2137);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5076__6783(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2151 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1549 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2131);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5077__3680(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2150 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1646 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2120);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5078__1617(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2160 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2102 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2136);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5079__2802(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2159 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1106 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2129);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5080__1705(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2158 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2085 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2132);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5081__5122(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2146 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2123 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2028);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5082__8246(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2145 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1321 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2130);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5083__7098(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2144 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2115 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2061);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5084__6131(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2143 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2115 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2061);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5085__1881(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2142 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2114 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2062);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5086__5115(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2141 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2117 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2059);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5087__7482(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2140 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2116 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2060);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5088__4733(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2139 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2113 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2063);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5089__6161(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2149 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2087 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2133);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5090__9315(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2148 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2084 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2134);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5091__9945(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2147 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2103 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1160);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5092__2883(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2137 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_558 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_701);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5093__2346(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2136 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2096 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2105);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5094__1666(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2135 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_556 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2090);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5095__7410(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2134 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2088 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2092);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5096__6417(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2133 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2086 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2093);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5097__5477(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2132 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2089 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2091);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5098__2398(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2131 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_566 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_701);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5099__5107(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2130 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_552 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2090);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5100__6260(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2129 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1128 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2103);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5101__4319(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2128 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1447 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2083);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5102__8428(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2127 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1582 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2095);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5103__5526(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2126 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1574 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2094);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5104__6783(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2125 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1666 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2101);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5105__3680(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2124 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1630 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2100);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5106__1617(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2138 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1587 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2097);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5107(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2119 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2118);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5108(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2116 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2117);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5109(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2113 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2114);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5110__2802(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2112 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_564 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_700);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5111__1705(out1[7] ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2046 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2050);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5112__5122(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2110 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2067 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1998);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5113__8246(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2109 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2057 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2008);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5114__7098(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2108 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2058 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2009);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5115__6131(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2107 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2064 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2006);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5116__1881(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2106 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2026 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2065);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5117__5115(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2123 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_185 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2071);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5118__7482(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2122 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2047 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2052);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5119__4733(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2121 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_10 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1617);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5120__6161(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2120 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_205 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2070);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5122__9315(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2118 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2044 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2049);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5123__9945(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2117 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_203 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2069);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5124__2883(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2115 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_195 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2068);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5125__2346(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2114 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_751 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2072);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5126(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2105 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2104);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5127__1666(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2102 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2066 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1997);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5128__7410(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2101 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1421 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2075);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5129__6417(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2100 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1340 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2077);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5130__5477(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2099 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2026 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2065);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5131__2398(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2098 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2026 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2065);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5132__5107(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2097 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1610 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_10);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5133__6260(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2096 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2067 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1998);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5134__4319(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2095 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1533 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2074);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5135__8428(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2094 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1530 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2076);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5136__5526(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2104 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2031 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2081);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5137__6783(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2103 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1117 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2080);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5139__3680(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2089 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2064 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2006);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5140__1617(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2088 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2058 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2009);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5141__2802(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2087 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2056 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2007);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5142__1705(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2086 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2057 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2008);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5143__5122(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2085 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2064 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2006);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5144__8246(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2084 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2058 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2009);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5145__7098(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2083 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1312 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2073);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5146__6131(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2093 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2036 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2054);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5147__1881(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2092 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2033 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2079);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5148__5115(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2091 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2035 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2078);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5149__7482(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2090 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2045 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1162);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5150__4733(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2081 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2042 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2046);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5151__6161(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2080 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1100 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2045);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5152__9315(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2079 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2032 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2044);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5153__9945(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2078 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2034 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2047);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5154__2883(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2077 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_403 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_674);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5155__2346(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2076 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_412 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2037);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5156__1666(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2075 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_385 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_674);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5157__7410(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2074 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_388 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2037);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5158__6417(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2073 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_391 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_673);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5159__5477(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2072 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1439 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2027);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5160__2398(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2071 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1672 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2039);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5161__5107(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2070 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1673 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2041);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5162__6260(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2069 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1572 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2043);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5163__4319(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2068 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1650 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2040);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5164__8428(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2082 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1594 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2038);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5165(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2066 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2067);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5166(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2062 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2063);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5167(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2060 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2059);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5168(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2056 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2057);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5169__5526(out1[6] ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1975 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1992);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5170__6783(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2054 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2030 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2048);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5171__3680(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2053 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2002 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1948);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5172__1617(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2052 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2003 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1951);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5173__2802(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2051 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2010 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1989);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5174__1705(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2050 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2005 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1943);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5175__5122(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2049 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1999 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1949);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5177__8246(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2067 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_240 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2014);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5178__7098(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2065 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2011 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1619);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5179__6131(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2064 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_199 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2012);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5180__1881(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2063 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1976 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1994);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5181__5115(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2061 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1979 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1991);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5182__7482(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2059 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1977 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1993);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5183__4733(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2058 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_757 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2015);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5184__6161(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2057 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_759 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2016);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5186__9315(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2043 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1522 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2019);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5187__9945(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2042 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2005 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1943);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5188__2883(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2041 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1423 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1996);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5189__2346(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2040 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1396 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2025);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5190__1666(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2039 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1471 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2023);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5191__7410(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2038 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1593 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2011);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5192__6417(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2048 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1981 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2022);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5193__5477(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2047 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1972 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2020);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5194__2398(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2046 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1969 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2021);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5195__5107(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2045 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1119 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2024);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5196__6260(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2044 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1986 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2017);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5197__4319(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2036 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2001 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1948);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5198__8428(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2035 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2004 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1951);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5199__5526(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2034 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2004 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1951);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5200__6783(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2033 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2000 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1949);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5201__3680(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2032 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2000 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1949);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5202__1617(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2031 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2005 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1943);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5203__2802(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2030 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2002 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1947);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5204__1705(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2029 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2010 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1989);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5205__5122(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2028 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2010 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1989);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5206__8246(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2027 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1373 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2018);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5207__7098(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2037 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1990 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1165);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5208__6131(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2025 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_144 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_664);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5209__1881(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2024 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1114 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1990);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5210__5115(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2023 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_140 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1974);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5211__7482(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2022 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1983 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1976);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5212__4733(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2021 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1973 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1975);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5213__6161(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2020 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1971 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1980);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5214__9315(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2019 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_146 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_664);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5215__9945(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2018 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_138 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1974);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5216__2883(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2017 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1985 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1978);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5217__2346(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2016 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1583 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1982);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5218__1666(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2015 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1660 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1987);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5219__7410(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2014 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1438 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1968);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5220__6417(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2013 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1680 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1988);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5221__5477(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2012 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1632 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1970);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5222__2398(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2026 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1598 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1984);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5223(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2008 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2007);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5224(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2004 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2003);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5225(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2001 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2002);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5226(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2000 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1999);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5227(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1997 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1998);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5228__5107(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1996 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_142 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_663);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5229__6260(out1[5] ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1933 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1936);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5230__4319(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1994 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_8 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1897);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5231__8428(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1993 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_4 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1894);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5232__5526(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1992 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1942 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1885);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5233__6783(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1991 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1946 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1887);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5234__3680(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2011 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_209 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1955);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5235__1617(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2010 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1952 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1618);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5236__2802(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2009 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1930 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1938);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5237__1705(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2007 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1935 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1937);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5238__5122(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2006 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1932 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1940);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5239__8246(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2005 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_235 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1954);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5240__7098(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2003 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_197 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1956);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5241__6131(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2002 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_166 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1957);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5242__1881(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1999 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_158 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1953);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5243__5115(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1998 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1931 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1939);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5244__7482(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1988 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1407 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1963);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5245__4733(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1987 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1402 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1966);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5246__6161(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1986 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1944 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1893);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5247__9315(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1985 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_4 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1894);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5248__9945(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1984 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1590 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1952);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5249__2883(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1983 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_8 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1897);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5250__2346(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1982 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1528 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1961);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5251__1666(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1981 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1950 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1896);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5252__7410(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1990 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1133 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1965);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5253__6417(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1989 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1929 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1964);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5254(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1980 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1979);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5255(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1978 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1977);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5256__5477(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1973 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1942 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1885);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5257__2398(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1972 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1945 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1886);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5258__5107(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1971 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1946 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1887);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5259__6260(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1970 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1355 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_26);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5260__4319(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1969 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1942 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1885);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5261__8428(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1968 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1371 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1962);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5262__5526(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1979 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1923 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1967);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5263__6783(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1977 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1922 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1959);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5264__3680(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1976 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1920 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1958);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5265__1617(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1975 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1915 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1960);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5266__2802(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1974 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1934 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1159);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5267__1705(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1967 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1917 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1930);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5268__5122(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1966 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_72 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_703);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5269__8246(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1965 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1102 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1934);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5270__7098(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1964 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1926 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1932);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5271__6131(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1963 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_63 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1924);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5272__1881(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1962 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_80 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_703);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5273__5115(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1961 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_60 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1924);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5274__7482(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1960 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1916 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1933);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5275__4733(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1959 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1921 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1935);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5276__6161(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1958 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1919 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1931);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5277__9315(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1957 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1581 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1927);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5278__9945(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1956 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1631 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1925);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5279__2883(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1955 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1592 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1918);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5280__2346(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1954 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1437 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1914);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5281__1666(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1953 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1643 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1928);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5282(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1950 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_8);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5283(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1947 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1948);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5284(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1945 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1946);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5285(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1944 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_4);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5287__7410(out1[4] ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1877 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1880);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5288__6417(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1940 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1487 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1898);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5289__5477(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1939 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1892 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1818);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5290__2398(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1938 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1813);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5291__5107(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1937 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1889 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1816);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5292__6260(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1936 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_24 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1814);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5293__4319(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1952 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_184 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1900);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5294__8428(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1951 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1876 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1878);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5296__5526(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1949 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1873 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1881);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5297__6783(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1948 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1875 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1882);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5298__3680(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1946 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_211 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1901);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5300__1617(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1943 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1866 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1879);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5301__2802(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1942 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_594 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1903);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5302__1705(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1929 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1487 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1898);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5303__5122(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1928 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1441 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1911);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5304__8246(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1927 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1612 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1904);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5305__7098(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1926 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1487 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1898);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5306__6131(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1925 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1413 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1884);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5307__1881(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1935 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1872 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1910);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5308__5115(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1934 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1110 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1912);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5309__7482(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1933 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1867 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1907);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5310__4733(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1932 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1862 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1905);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5311__6161(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1931 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1857 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1913);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5312__9315(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1930 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1864 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1906);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5313__9945(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1923 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1890 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1813);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5314__2883(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1922 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1888 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1816);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5315__2346(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1921 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1889 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1815);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5316__1666(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1920 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1891 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1818);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5317__7410(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1919 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1892 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1817);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5318__6417(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1918 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1543 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1909);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5319__5477(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1917 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1890 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1813);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5320__2398(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1916 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1895 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1814);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5321__5107(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1915 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1895 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1814);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5322__6260(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1914 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1382 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1908);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5323__4319(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1924 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1874 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1158);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5324__8428(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1913 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1856 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1866);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5325__5526(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1912 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1112 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1874);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5326__6783(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1911 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_588 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_695);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5327__3680(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1910 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1869 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1875);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5328__1617(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1909 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_582 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1865);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5329__2802(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1908 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_585 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_695);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5330__1705(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1907 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1871 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1877);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5331__5122(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1906 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1861 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1873);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5332__8246(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1905 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1870 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1876);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5333__7098(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1904 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_591 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1865);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5334__6131(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1903 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1446 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1863);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5335__1881(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1902 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1580 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1859);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5336__5115(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1901 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1629 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1860);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5337__7482(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1900 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1586 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1858);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5338__4733(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1899 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1662 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1868);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5339(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1896 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1897);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5340(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1895 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_24);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5341(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1893 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1894);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5342(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1891 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1892);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5343(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1890 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5344(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1888 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1889);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5345(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1886 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1887);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5346__6161(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1884 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_579 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_694);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5347__9315(out1[3] ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1803 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1832);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5348__9945(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1882 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1790);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5349__2883(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1881 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_3 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1792);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5350__2346(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1880 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1842 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1781);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5351__1666(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1879 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_13 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_27);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5352__7410(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1878 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1489 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1839);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5353__6417(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1898 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_205 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1843);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5354__5477(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1897 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1801 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1831);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5356__2398(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1894 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1804 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1830);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5357__5107(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1892 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_164 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1846);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5359__6260(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1889 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_160 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1847);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5360__4319(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1887 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1805 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1834);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5361__8428(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1885 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_14 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1833);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5362__5526(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1872 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1790);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5363__6783(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1871 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1841 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1781);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5364__3680(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1870 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1489 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1839);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5365__1617(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1869 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1790);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5366__2802(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1868 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1429 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1837);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5367__1705(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1867 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1842 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1780);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5368__5122(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1877 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1810 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1852);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5369__8246(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1876 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1822 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1850);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5370__7098(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1875 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1819 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1851);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5371__6131(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1874 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1113 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1849);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5372__1881(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1873 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1821 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1855);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5373__5115(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1864 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1838 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1791);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5374__7482(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1863 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1309 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1854);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5375__4733(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1862 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1489 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1839);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5376__6161(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1861 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_3 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1792);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5377__9315(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1860 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1445 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1835);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5378__9945(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1859 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1541 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1853);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5379__2883(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1858 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1575 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1836);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5380__2346(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1857 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1840 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_27);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5381__1666(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1856 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_13 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1782);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5382__7410(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1866 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1807 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1848);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5383__6417(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1865 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1829 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1167);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5384__5477(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1855 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1820 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1804);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5385__2398(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1854 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_552 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_671);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5386__5107(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1853 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_566 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1812);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5387__6260(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1852 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1803 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1809);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5388__4319(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1851 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1826 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1801);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5389__8428(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1850 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1828 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1805);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5390__5526(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1849 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1101 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1829);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5391__6783(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1848 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1811 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1802);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5392__3680(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1847 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1633 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1823);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5393__1617(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1846 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1642 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1827);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5394__2802(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1845 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1597 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1825);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5395__1705(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1844 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1434 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1808);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5396__5122(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1843 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1601 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1824);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5397(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1842 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1841);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5398(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1840 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_13);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5399(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1838 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_3);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5400__8246(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1837 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_558 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_671);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5401__7098(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1836 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_564 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1812);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5402__6131(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1835 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_556 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_670);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5403__1881(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1834 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1292 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1786);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5404__5115(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1833 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_16 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1802);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5405__7482(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1832 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_20 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1784);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5406__4733(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1831 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_17 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_12);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5407__6161(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1830 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_15 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_6);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5409__9315(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1841 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_751 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1795);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5411__9945(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1839 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_207 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1797);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5413__2883(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1828 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1291 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1786);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5414__2346(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1827 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1378 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1798);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5415__1666(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1826 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1751 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_12);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5416__7410(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1825 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1614 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1779);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5417__6417(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1824 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1514 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1777);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5418__5477(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1823 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1417 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1778);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5419__2398(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1822 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1292 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1785);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5420__5107(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1821 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_15 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1787);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5421__6260(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1820 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1752 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_6);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5422__4319(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1819 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_17 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1789);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5423__8428(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1829 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1111 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1800);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5424(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1817 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1818);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5425(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1815 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1816);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5426__5526(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1811 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1750 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_14);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5427__6783(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1810 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_20 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1783);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5428__3680(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1809 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1749 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1784);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5429__1617(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1808 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1311 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1799);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5430__2802(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1807 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_16 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1788);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5431__1705(out1[2] ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1753 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1767);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5432__5122(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1818 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1755 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1768);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5433__8246(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1816 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_11 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1773);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5434__7098(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1814 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1757 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1775);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5435__6131(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1813 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1765 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1771);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5436__1881(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1812 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1770 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1163);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5437__5115(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1800 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1132 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1770);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5438__7482(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1799 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_390 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_677);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5439__4733(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1798 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_387 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1748);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5440__6161(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1797 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1579 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1764);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5441__9315(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1796 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1570 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1761);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5442__9945(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1795 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1443 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1760);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5443__2883(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1794 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1657 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1762);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5444__2346(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1793 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1628 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1763);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5445__1666(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1805 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1766 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1772);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5446__7410(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1804 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1759 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1774);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5447__6417(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1803 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1754 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1767);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5448__5477(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1802 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1758 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1776);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5449__2398(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1801 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1756 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1769);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5450(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1791 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1792);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5451(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1789 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_12);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5452(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1788 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_14);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5453(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1787 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_6);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5454(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1785 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1786);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5455(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1783 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1784);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5456(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1782 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_27);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5457(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1780 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1781);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5458__5107(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1779 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_411 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_677);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5459__6260(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1778 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_384 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1748);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5460__4319(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1777 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_402 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_676);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5462__8428(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1792 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1741 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1722);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5463__5526(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1790 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1737 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1725);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5467__6783(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1786 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_193 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1726);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5468__3680(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1784 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_755 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1727);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5470__1617(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1781 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1735 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1724);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5471(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1776 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1775);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5472(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1774 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1773);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5473(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1772 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1771);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5474(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1769 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1768);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5475(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1766 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1765);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5476__2802(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1764 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1548 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1712);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5477__1705(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1763 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1322 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1709);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5478__5122(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1762 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1419 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1713);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5479__8246(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1761 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1524 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1711);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5480__7098(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1760 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1358 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1714);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5481__6131(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1775 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1736 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1724);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5482__1881(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1773 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1738 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1725);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5483__5115(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1771 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1742 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1722);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5484__7482(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1770 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1129 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1731);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5485__4733(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1768 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1740 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1721);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5486__6161(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1767 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1743 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1723);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5487__9315(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1765 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_229 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1682);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5488(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1759 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_11);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5489(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1758 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1757);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5490(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1756 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1755);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5491(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1754 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1753);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5492(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1752 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_15);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5493(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1751 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_17);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5494(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1750 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_16);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5495(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1749 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_20);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5496__9945(out1[0] ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_0 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1072);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5497__2883(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1746 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1706 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1478);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5498__2346(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1745 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1705 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_921);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5499__1666(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1744 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1197 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1698);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5501__7410(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1757 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_181 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1697);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5502__6417(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1755 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_201 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1701);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5503__5477(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1753 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_594 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1700);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5508__2398(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1748 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1707 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1168);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5509(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1742 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1741);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5510(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1740 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1739);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5511(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1738 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1737);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5512(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1736 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1735);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5513__5107(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1734 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_600 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1706);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5514__6260(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1733 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_600 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1706);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5515__4319(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1732 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_909 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1705);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5516__8428(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1731 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1107 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1707);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5517__5526(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1730 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1641 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1684);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5518__6783(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1729 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1655 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1703);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5519__3680(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1728 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1571 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1702);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5520__1617(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1727 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1430 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1685);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5521__2802(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1726 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1577 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1704);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5522__1705(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1743 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1073 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1688);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5523__5122(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1741 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_979 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1690);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5524__8246(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1739 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_736 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1692);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5525__7098(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1737 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_628 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1694);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5526__6131(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1735 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_739 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1696);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5529(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1719 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1720);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5530(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1717 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1718);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5531(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1716 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1715);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5532__1881(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1714 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_394 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_683);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5533__5115(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1713 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_400 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1687);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5534__7482(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1712 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_406 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_683);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5535__4733(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1711 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_397 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1687);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5536__6161(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1710 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_909 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1705);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5537__9315(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1709 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_409 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_682);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5538__9945(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1708 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1647 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_919);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5539__2883(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1725 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_156 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1648);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5540__2346(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1724 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_178 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1625);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5541__1666(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1723 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1072 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1623);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5542__7410(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1722 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_170 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1624);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5543__6417(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1721 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_746 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1649);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5544__5477(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1720 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_18 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1479);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5545__2398(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1718 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_19 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1480);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5546__5107(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1715 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_22 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_977);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5547__6260(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1704 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1567 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1640);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5548__4319(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1703 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1398 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1638);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5549__8428(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1702 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1566 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1644);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5550__5526(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1701 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1589 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1654);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5551__6783(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1700 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1451 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1627);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5552__3680(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1699 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1609 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1679);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5553__1617(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1698 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_25 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1665);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5554__2802(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1697 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1602 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1674);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5555__1705(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1707 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1131 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1635);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5556__5122(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1706 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1503 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1671);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5557__8246(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1705 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1500 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1634);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5558(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1696 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1695);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5559(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1694 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1693);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5560(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1692 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1691);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5561(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1690 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1689);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5562(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1688 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_0);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5563__7098(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1686 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_907 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1647);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5564__6131(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1685 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1310 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1626);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5565__1881(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1684 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1361 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1636);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5566__5115(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1683 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_907 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1647);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5567__7482(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1682 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1595 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1639);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5568__4733(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1695 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_179 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1556);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5569__6161(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1693 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_162 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1558);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5570__9315(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1691 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_174 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1557);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5571__9945(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1689 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_209 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1559);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5573__2883(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1687 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1616 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1170);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5574__2346(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1681 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1354 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1513);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5575__1666(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1680 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1336 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1516);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5576__7410(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1679 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1608 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1505);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5577__6417(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1678 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1463 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1523);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5578__5477(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1677 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1436 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1512);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5579__2398(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1676 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1351 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1585);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5580__5107(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1675 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1303 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1613);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5581__6260(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1674 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1606 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1508);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5582__4319(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1673 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1368 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1545);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5583__8428(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1672 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1343 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1531);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5584__5526(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1671 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1494 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1502);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5585__6783(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1670 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1362 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1550);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5586__3680(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1669 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1374 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1551);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5587__1617(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1668 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1357 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1527);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5588__2802(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1667 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1366 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1546);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5589__1705(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1666 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1320 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1544);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5590__5122(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1665 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1493 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1504);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5591__8246(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1664 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1448 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1538);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5592__7098(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1663 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1344 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1542);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5593__6131(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1662 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1327 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1536);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5594__1881(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1661 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1334 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1521);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5595__5115(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1660 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1356 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1539);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5596__7482(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1659 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1367 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1535);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5597__4733(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1658 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1365 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1561);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5598__6161(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1657 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1349 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1540);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5599(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1656 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1350 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1511);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5600(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1655 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1342 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1565);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5601(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1654 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1584 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1506);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5602(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1653 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1459 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1526);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5603(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1652 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1341 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1518);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5604(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1651 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1325 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1532);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5605(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1650 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1346 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1520);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5606(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1649 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1469 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1588);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5607(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1648 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1300 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1607);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5608(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1645 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1332 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1517);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5609(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1644 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_78 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_698);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5610(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1643 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1324 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1537);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5611(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1642 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1308 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1529);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5612(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1641 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1328 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1569);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5613(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1640 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_64 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1555);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5614(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1639 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1573 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1507);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5615(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1638 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_73 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_698);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5616(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1637 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1353 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1547);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5617(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1636 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_61 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1555);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5618(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1635 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1130 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1616);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5619(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1634 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1492 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1501);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5620(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1633 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1319 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1534);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5621(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1632 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1405 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1552);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5622(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1631 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1339 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1515);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5623(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1630 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1418 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1519);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5624(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1629 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1369 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1510);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5625(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1628 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1315 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1525);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5626(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1627 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1347 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1509);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5627(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1626 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_81 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_697);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5628(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1625 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1298 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1596);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5629(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1624 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1297 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1576);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5630(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1623 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1304 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1604);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5634(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1622 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_598 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1484);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5635(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1621 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_596 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1482);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5636(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1620 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1491 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1478);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5637(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1619 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1488 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_235);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5638(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1618 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1485 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_241);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5639(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1617 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1486 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_755);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5640(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1647 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1105 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1578);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5641(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1646 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1495 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1171);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5642(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1615 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1313 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1370);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5643(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1614 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_456 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_962);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5644(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1613 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_438 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_935);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5645(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1612 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_486 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_929);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5646(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1611 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_414 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_944);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5647(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1610 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_148 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1486);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5648(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1609 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1470 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1428);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5649(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1608 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_742 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_624);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5650(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1607 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1460 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1425);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5651(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1606 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_743 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_609);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5652(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1605 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1359 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1427);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5653(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1604 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1219 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1466);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5654(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1603 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1490 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1478);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5655(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1602 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1453 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1380);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5656(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1601 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1318 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1403);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5657(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1600 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1317 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1454);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5658(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1599 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1337 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1416);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5659(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1598 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_234 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1485);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5660(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1597 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1306 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1426);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5661(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1596 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1462 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1450);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5662(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1595 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1461 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1444);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5663(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1594 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_240 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1488);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5664(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1593 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_234 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1488);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5665(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1592 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1305 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1420);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5666(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1591 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_977 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1491);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5667(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1590 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_237 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1485);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5668(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1589 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1465 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1415);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5669(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1588 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1456 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1299);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5670(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1587 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_150 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1486);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5671(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1586 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1379 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1440);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5672(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1585 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_450 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_953);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5673(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1584 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_617 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_608);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5674(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1583 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1375 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1316);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5675(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1582 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1364 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1381);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5676(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1581 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1335 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1363);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5677(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1580 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1338 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1333);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5678(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1579 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1314 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1408);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5679(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1578 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1099 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1495);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5680(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1577 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1348 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1401);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5681(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1576 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1468 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1433);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5682(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1575 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_459 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_947);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5683(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1574 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1326 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1400);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5684(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1573 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_617 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_605);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5685(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1572 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1307 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1372);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5686(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1571 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1352 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1409);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5687(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1570 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1323 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1397);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5688(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1569 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_498 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_930);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5689(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1568 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_475 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_956);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5690(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1567 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_498 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_948);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5691(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1566 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_572 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_957);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5692(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1565 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_509 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_938);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5693(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1564 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_37 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_950);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5694(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1563 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_570 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_939);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5695(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1562 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_507 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_932);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5696(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1561 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_468 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_954);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5697(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1560 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_187 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1296);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5698(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1559 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_232 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1294);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5699(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1558 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_191 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1301);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5700(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1557 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_189 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1295);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5701(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1556 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_231 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1302);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5702(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1616 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1104 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1431);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5703(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1554 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_450 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_941);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5704(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1553 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_468 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_936);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5705(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1552 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_480 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_959);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5706(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1551 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_441 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_945);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5707(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1550 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_414 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_963);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5708(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1549 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_441 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_932);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5709(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1548 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_489 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_950);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5710(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1547 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_426 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_959);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5711(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1546 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_426 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_933);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5712(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1545 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_477 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_951);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5713(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1544 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_417 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_941);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5714(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1543 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_486 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_951);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5715(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1542 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_532 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_933);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5716(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1541 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_459 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_936);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5717(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1540 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_489 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_942);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5718(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1539 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_480 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_942);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5719(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1538 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_438 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_954);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5720(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1537 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_516 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_945);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5721(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1536 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_540 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_913);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5722(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1535 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_514 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_915);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5723(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1534 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_456 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1386);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5724(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1533 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_417 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_911);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5725(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1532 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_518 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1475);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5726(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1531 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_477 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_960);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5727(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1530 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_522 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_960);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5728(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1529 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_548 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_935);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5729(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1528 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_560 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_930);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5730(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1527 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_546 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_963);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5731(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1526 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_526 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_917);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5732(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1525 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_575 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_911);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5733(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1524 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_512 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1394);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5734(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1523 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_530 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_944);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5735(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1522 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_577 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_929);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5736(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1521 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_534 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_962);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5737(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1520 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_550 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_939);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5738(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1519 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_528 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1390);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5739(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1518 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_542 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_953);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5740(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1517 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_520 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_913);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5741(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1516 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_568 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_948);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5742(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1515 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_536 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_957);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5743(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1514 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_562 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_915);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5744(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1513 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_524 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_947);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5745(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1512 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_538 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_917);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5746(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1511 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_554 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_938);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5747(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1510 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_544 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_956);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5748(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1509 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_391 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_661);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5749(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1508 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_388 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1395);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5750(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1507 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_403 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_661);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5751(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1506 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_385 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1395);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5752(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1505 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_412 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_660);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5753(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1504 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_980 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1478);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5755(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1503 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_628 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_598);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5756(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1502 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_734 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_650);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5757(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1501 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_745 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_596);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5758(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1500 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_745 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_648);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5759(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1499 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1481 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_648);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5760(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1498 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1065 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_919);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5761(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1497 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1483 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_650);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5762(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1496 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1064 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_921);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5763(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1555 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1293 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1169);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5764(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1490 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1491);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5765(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1483 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1484);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5766(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1481 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1482);
  buf mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5769(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1478 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1476);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5770(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1477 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1476);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5771(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1475 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1474);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5772(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1473 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_609);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5774(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1472 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1474);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5775(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1471 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_442 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_328);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5776(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1470 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_499 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_274);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5777(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1469 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_502 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_298);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5778(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1468 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_367 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_189);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5779(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1467 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1212 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1277);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5780(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1466 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_573 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_310);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5781(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1465 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_510 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_334);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5782(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1464 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1204 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1282);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5783(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1463 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_493 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_325);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5784(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1462 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_364 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_765);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5785(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1461 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_501 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_304);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5786(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1460 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_370 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_187);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5787(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1459 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_475 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_273);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5788(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1458 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_51 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_340);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5789(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1457 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1200 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1257);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5790(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1456 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_373 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_191);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5791(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1455 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1179 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1268);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5792(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1454 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_492 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_265);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5793(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1453 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_501 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_361);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5794(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1452 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1207 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1256);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5795(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1451 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1209 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1255);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5796(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1450 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_572 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_259);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5797(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1449 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_492 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_289);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5798(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1448 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_474 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_366);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5799(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1447 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1176 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1276);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5800(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1446 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1184 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1279);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5801(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1445 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_481 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_262);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5802(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1444 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_490 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_283);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5803(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1443 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1203 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1254);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5804(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1442 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_570 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_327);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5805(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1441 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_478 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_297);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5806(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1440 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_484 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_295);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5807(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1439 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1181 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1269);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5808(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1438 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1202 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1274);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5809(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1437 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1198 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1278);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5810(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1436 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_469 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_244);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5811(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1435 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1182 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1267);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5812(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1434 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1201 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1281);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5813(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1433 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_509 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_282);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5814(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1432 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_507 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_256);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5815(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1431 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1108 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1293);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5816(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1430 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1205 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1280);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5817(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1429 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_69 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_253);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5818(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1428 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_496 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_243);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5819(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1427 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_427 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_252);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5820(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1426 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_487 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_328);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5821(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1425 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_499 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_327);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5822(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1424 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_439 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_300);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5823(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1423 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_448 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_255);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5824(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1422 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_451 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_298);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5825(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1421 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_415 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_297);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5826(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1420 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_436 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_283);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5827(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1419 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_460 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_291);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5828(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1418 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_421 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_282);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5829(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1417 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_424 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_292);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5830(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1416 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_472 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_292);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5831(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1415 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_48 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_253);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5832(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1414 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_88 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_279);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5833(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1413 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_45 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_301);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5834(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1412 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_433 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_280);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5835(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1411 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_454 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_301);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5836(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1410 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_109 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_280);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5837(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1409 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_457 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_244);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5838(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1408 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_463 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_256);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5839(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1407 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_418 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_279);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5840(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1406 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_445 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_294);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5841(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1405 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_430 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_300);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5842(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1404 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_118 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_291);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5843(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1403 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_132 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_294);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5844(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1402 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_123 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_288);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5845(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1401 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_466 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_295);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5846(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1400 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_135 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_261);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5847(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1399 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_126 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_261);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5848(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1398 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_57 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_288);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5849(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1397 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_97 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_262);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5850(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1396 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_106 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_289);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5851(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1495 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1177 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1245);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5852(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1494 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1216 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1239);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5853(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1493 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1206 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1253);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5854(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1492 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1186 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1250);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5855(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1491 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1183 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1243);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5856(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1489 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1223 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1252);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5857(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1488 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1174 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1241);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5858(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1487 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1208 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1248);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5859(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1486 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1178 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1249);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5860(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1485 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1175 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1244);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5861(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1484 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1225 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1242);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5862(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1482 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1185 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1247);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5863(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1480 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1180 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1246);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5864(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1479 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1199 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1240);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5865(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1476 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1211 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1251);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5866(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1474 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1283 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1284);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5867(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1394 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1393);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5868(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1392 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_624);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5870(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1391 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1393);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5871(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1390 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1389);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5872(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1388 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_605);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5874(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1387 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1389);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5875(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1386 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1385);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5876(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1384 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_608);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5878(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1383 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1385);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5879(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1382 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_83 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_309);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5880(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1381 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_129 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_264);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5881(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1380 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_39 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_250);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5882(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1379 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_103 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_268);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5883(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1378 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_91 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_363);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5884(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1377 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_75 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_249);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5885(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1376 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_432 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_331);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5886(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1375 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_435 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_355);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5887(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1374 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_420 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_277);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5888(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1373 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_94 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_247);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5889(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1372 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_447 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_265);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5890(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1371 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_115 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_246);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5891(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1370 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_100 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_264);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5892(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1369 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_423 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_330);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5893(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1368 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_429 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_267);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5894(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1367 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_453 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_349);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5895(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1366 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_54 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_354);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5896(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1365 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_112 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_348);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5897(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1364 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_447 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_322);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5898(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1363 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_435 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_285);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5899(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1362 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_453 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_274);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5900(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1361 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_66 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_286);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5901(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1360 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_432 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_310);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5902(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1359 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_532 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_276);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5903(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1358 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_462 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_309);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5904(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1357 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_444 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_273);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5905(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1356 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_577 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_334);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5906(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1355 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_550 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_270);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5907(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1354 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_471 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_367);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5908(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1353 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_471 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_271);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5909(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1352 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_495 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_271);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5910(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1351 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_520 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_349);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5911(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1350 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_444 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_333);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5912(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1349 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_465 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_373);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5913(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1348 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_495 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_366);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5914(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1347 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_575 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_306);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5915(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1346 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_429 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_372);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5916(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1345 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_546 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_307);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5917(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1344 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_524 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_321);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5918(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1343 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_522 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_331);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5919(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1342 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_512 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_372);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5920(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1341 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_420 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_268);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5921(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1340 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_534 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_348);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5922(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1339 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_42 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_270);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5923(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1338 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_423 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_364);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5924(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1337 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_427 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_277);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5925(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1336 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_478 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_303);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5926(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1335 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_483 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_322);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5927(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1334 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_514 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_369);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5928(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1333 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_483 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_286);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5929(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1332 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_554 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_333);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5930(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1331 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_526 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_250);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5931(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1330 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_469 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_285);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5932(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1329 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_530 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_307);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5933(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1328 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_490 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_363);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5934(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1327 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_516 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_324);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5935(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1326 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_542 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_369);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5936(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1325 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_538 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_355);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5937(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1324 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_560 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_324);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5938(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1323 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_465 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_370);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5939(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1322 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_548 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_321);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5940(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1321 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_451 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_247);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5941(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1320 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_442 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_325);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5942(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1319 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_462 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_276);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5943(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1318 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_540 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_303);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5944(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1317 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_439 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_360);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5945(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1316 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_528 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_258);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5946(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1315 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_544 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_258);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5947(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1314 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_562 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_304);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5948(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1313 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_518 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_360);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5949(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1312 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_415 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_306);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5950(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1311 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_536 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_339);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5951(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1310 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_457 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_339);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5952(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1309 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_568 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_340);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5953(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1308 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_487 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_259);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5954(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1307 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_418 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_361);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5955(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1306 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_460 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_330);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5956(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1305 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_481 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_267);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5957(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1304 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_138 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_667);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5958(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1303 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_493 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_354);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5959(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1302 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_61 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_249);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5960(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1301 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_78 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_243);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5961(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1300 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_140 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1188);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5962(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1299 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_144 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_667);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5963(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1298 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_146 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1188);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5964(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1297 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_142 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_666);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5965(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1296 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_81 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_246);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5966(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1295 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_73 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_252);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5967(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1294 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_64 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_255);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5968(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1395 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1144 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1166);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5969(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1393 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1273 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1271);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5970(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1389 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1270 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1238);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5971(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1385 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1275 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1272);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5972(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1292 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1291);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5973(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1284 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_972 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1222);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5974(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1283 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_615 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1210);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5975(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1282 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_421 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_358);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5976(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1281 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_466 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_337);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5977(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1280 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_502 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_357);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5978(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1279 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_463 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_337);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5979(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1278 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_424 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_376);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5980(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1277 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_454 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_358);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5981(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1276 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_430 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_357);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5982(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1275 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_749 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1228);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5983(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1274 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_484 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_312);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5984(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1273 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_746 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1224);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5985(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1272 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_748 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1227);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5986(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1271 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_736 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1226);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5987(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1270 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1025 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1229);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5988(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1269 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_436 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_313);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5989(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1268 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_448 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_313);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5990(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1267 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_433 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_375);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5991(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1266 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_474 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_312);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5992(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1293 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1109 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1218);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5993(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1291 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_742 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_220);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5994(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1290 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1221 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1213);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5995(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1289 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1215 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1217);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5996(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1288 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1214 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1220);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5997(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1287 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1096 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1195);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5998(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1286 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1193 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1194);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g5999(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1285 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1096 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1196);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6000(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1257 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_472 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_375);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6001(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1256 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_445 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_336);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6002(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1255 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_376 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_762);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6003(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1254 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_496 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_336);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6004(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1253 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_611 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_223);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6005(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1252 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_595 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_219);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6006(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1251 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_709 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_217);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6007(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1250 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_644 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_216);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6008(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1249 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_619 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_220);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6009(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1248 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_715 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_219);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6010(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1247 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_602 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_213);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6011(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1246 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_705 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_214);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6012(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1245 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_711 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_214);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6013(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1244 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_638 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_217);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6014(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1243 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_630 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_213);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6015(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1242 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_655 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_222);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6016(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1241 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_640 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_222);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6017(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1240 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_604 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_223);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6018(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1239 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_621 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_216);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6019(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1238 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_733 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1230);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6020(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1265 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1172 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1173);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6021(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1264 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1191 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1232);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6022(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1263 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1190 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1234);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6023(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1262 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1189 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1236);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6024(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1261 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1194 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1192);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6025(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1260 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1233 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1191);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6026(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1259 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1235 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1190);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6027(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1258 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1237 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1189);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6028(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1237 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1236);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6029(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1235 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1234);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6030(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1233 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1232);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6031(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1230 ,n_186 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1154);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6032(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1229 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_903 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1155);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6033(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1228 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_901 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1145);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6034(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1227 ,n_180 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1148);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6035(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1226 ,n_183 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1152);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6036(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1225 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_107 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_343);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6037(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1224 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_905 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1149);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6038(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1223 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_379 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_232);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6039(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1222 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_597 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1124);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6040(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1221 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_734 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1137);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6041(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1220 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_166 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1140);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6042(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1219 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_382 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_761);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6044(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1217 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_158 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1139);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6045(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1216 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_110 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_352);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6046(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1215 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_737 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1141);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6047(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1214 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_749 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1127);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6048(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1213 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_152 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1138);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6049(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1212 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_127 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_319);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6050(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1211 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_76 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_351);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6051(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1210 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_965 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1125);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6052(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1209 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_86 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_381);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6053(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1208 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_121 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_342);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6054(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1207 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_52 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_316);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6055(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1206 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_119 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_351);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6056(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1205 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_49 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_315);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6057(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1204 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_101 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_346);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6058(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1203 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_58 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_345);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6059(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1202 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_46 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_382);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6060(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1201 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_98 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_346);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6061(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1200 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_113 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_381);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6062(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1199 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_136 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_352);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6063(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1198 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_70 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_316);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6064(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1236 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1146 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1147);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6065(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1234 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1156 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1153);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6066(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1197 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_52 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_34);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6067(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1232 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1150 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1151);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6068(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1231 ,n_174 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1126);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6069(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1196 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1195);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6070(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1193 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1192);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6071(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1186 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_124 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_505);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6072(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1185 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_43 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_379);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6073(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1184 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_133 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_345);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6074(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1183 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_89 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_343);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6075(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1182 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_55 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_318);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6076(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1181 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_116 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_318);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6077(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1180 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_84 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_342);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6078(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1179 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_130 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_319);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6079(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1178 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_92 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_378);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6080(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1177 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_104 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_378);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6081(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1176 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_95 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_315);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6082(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1175 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_40 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_505);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6083(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1174 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_67 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_504);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6084(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1173 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_225 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1135);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6085(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1172 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1073 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1136);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6086(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1171 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1125 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1123);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6087(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1170 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_642 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_638);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6088(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1195 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_926 ,n_175);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6089(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1194 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_241 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_971);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6090(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1192 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_748 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_965);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6091(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1191 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_737 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1082);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6092(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1190 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_733 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1080);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6093(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1189 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_739 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1081);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6094(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1169 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_636 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_715);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6095(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1168 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_719 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1006);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6096(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1167 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_707 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_711);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6097(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1166 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_613 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_969);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6098(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1165 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_646 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_644);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6099(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1164 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_611 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_630);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6100(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1163 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_626 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1000);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6101(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1162 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_717 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1003);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6102(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1161 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_634 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_709);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6103(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1160 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_713 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_997);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6104(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1159 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_632 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_705);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6105(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1158 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_607 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1015);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6106(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1157 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_623 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_991);
  xnor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6107(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1188 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_595 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1022);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6108(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1187 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_34 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1118);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6109(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1156 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1155);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6110(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1154 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1153);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6111(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1152 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1151);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6112(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1150 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1149);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6113(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1148 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1147);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6114(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1146 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1145);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6115(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1142 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_985 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_992);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6116(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1141 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_905 ,n_184);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6117(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1140 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_895 ,n_180);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6118(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1139 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_897 ,n_183);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6119(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1138 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_899 ,n_186);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6120(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1137 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_903 ,n_187);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6121(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1136 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1095 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_597);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6122(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1135 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1056 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_615);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6123(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1134 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_974 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_982);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6124(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1133 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_107 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_124);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6125(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1132 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_988 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1001);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6126(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1131 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_98 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_58);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6127(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1130 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1007 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1018);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6128(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1129 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_133 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_92);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6129(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1128 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_713 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_998);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6130(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1127 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_901 ,n_181);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6131(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1155 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1083 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_207);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6132(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1153 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_193 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_899);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6133(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1151 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_156 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1098);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6134(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1149 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_897 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_162);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6135(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1147 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_160 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1097);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6136(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1145 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_895 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_154);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6137(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1126 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_927 ,n_175);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6138(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1144 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_86 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_231);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6139(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1143 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1084 ,n_174);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6140(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1124 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1123);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6141(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1121 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_119 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_89);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6143(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1119 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_136 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_95);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6144(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1118 ,n_189 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_228);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6145(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1117 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_110 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_130);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6146(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1116 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_983 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_986);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6147(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1115 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_36 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_113);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6148(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1114 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1004 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1009);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6149(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1113 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_46 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_70);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6150(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1112 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1012 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1016);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6151(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1111 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_43 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_104);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6152(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1110 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_116 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_84);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6153(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1109 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_49 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_121);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6154(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1108 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1019 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_995);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6155(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1107 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_719 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_642);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6156(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1106 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_127 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_101);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6157(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1105 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_238 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_182);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6158(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1104 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_67 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_40);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6159(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1103 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_55 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_76);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6160(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1102 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1010 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1013);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6161(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1101 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_707 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_989);
  nor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6162(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1100 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_717 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_646);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6163(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1099 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_740 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_927);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6164(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1125 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_226 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_740);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6165(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1123 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_176 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_926);
  or mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6166(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1122 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1085 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_980);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6167(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1098 ,n_184);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6168(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1097 ,n_181);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6169(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1096 ,n_174);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6170(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1095 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_972);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6171(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1094 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_743);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6173(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1093 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_619);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6174(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1092 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_602);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6175(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1091 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_636);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6176(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1090 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_632);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6177(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1089 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_607);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6178(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1088 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_613);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6179(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1087 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_626);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6180(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1086 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_623);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6183(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1085 ,n_189);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6184(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1084 ,n_175);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6185(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1083 ,n_187);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6186(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1082 ,n_183);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6187(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1081 ,n_180);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6188(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1080 ,n_186);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6190(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1079 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_975);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6191(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1078 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_640);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6192(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1077 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_604);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6193(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1076 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_634);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6194(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1075 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_621);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6195(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1074 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_655);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6198(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1073 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1071);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6199(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1072 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1071);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6200(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1071 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_924);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6201(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1070 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_923);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6202(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1068 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_923);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6204(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1067 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_924);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g6205(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1069 ,n_176);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1052 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_727);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6206(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1051 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_728);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6207(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1050 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_727);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6208(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1049 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_728);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6209(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1048 ,n_188);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6213(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1047 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_724);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6214(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1046 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_725);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6215(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1045 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_724);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6216(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1044 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_725);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6217(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1043 ,n_185);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6221(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1042 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_721);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6222(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1041 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_722);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6223(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1040 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_721);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6224(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1039 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_722);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6225(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1038 ,n_179);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6229(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1037 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_730);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6230(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1036 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_731);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6231(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1035 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_730);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6232(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1034 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_731);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6233(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1033 ,n_182);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6328(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1032 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1030);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6329(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1031 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1030);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6330(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1030 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1059);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6486(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1029 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1028);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6488(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1028 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1054);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6491(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1027 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1026);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6493(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1026 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1057);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6496(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1025 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1023);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6497(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1024 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1023);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6498(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1023 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1055);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6500(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1022 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1020);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6501(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1021 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1020);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6502(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1020 ,n_190);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6508(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1019 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1017);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6509(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1018 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1017);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6510(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1017 ,n_193);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6512(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1016 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1014);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6513(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1015 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1014);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6514(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1014 ,n_197);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6516(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1013 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1011);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6517(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1012 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1011);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6518(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1011 ,n_198);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6520(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1010 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1008);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6521(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1009 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1008);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6522(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1008 ,n_199);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6524(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1007 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1005);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6525(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1006 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1005);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6526(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1005 ,n_194);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6528(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1004 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1002);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6529(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1003 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1002);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6530(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1002 ,n_200);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6532(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1001 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_999);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6533(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1000 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_999);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6534(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_999 ,n_195);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6536(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_998 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_996);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6537(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_997 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_996);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6538(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_996 ,n_201);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6540(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_995 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_993);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6541(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_994 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_993);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6542(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_993 ,n_192);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6544(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_992 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_990);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6545(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_991 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_990);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6546(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_990 ,n_202);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6548(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_989 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_987);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6549(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_988 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_987);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6550(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_987 ,n_196);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6552(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_986 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_984);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6553(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_985 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_984);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6554(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_984 ,n_203);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6556(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_983 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_981);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6557(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_982 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_981);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6558(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_981 ,n_204);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6570(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1053 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1067);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6572(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_980 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_978);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6573(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_979 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_978);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6574(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_978 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1058);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6576(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_977 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_976);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6578(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_976 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1477);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6644(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_975 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_973);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6645(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_974 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_973);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6646(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_973 ,n_205);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6648(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_972 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_970);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6649(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_971 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_970);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6650(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_970 ,n_177);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6668(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_969 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_967);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6669(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_968 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_967);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6670(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_967 ,n_191);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6672(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_966 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_964);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6673(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_965 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_964);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6674(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_964 ,n_178);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6676(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_963 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_961);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6677(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_962 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_961);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6678(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_961 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1392);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6680(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_960 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_958);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6681(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_959 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_958);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6682(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_958 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1062);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6684(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_957 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_955);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6685(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_956 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_955);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6686(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_955 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1391);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6688(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_954 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_952);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6689(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_953 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_952);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6690(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_952 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1388);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6692(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_951 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_949);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6693(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_950 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_949);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6694(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_949 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1061);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6696(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_948 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_946);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6697(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_947 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_946);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6698(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_946 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1387);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6700(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_945 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_943);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6701(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_944 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_943);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6702(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_943 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1384);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6704(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_942 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_940);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6705(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_941 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_940);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6706(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_940 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1060);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6708(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_939 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_937);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6709(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_938 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_937);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6710(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_937 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1383);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6712(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_936 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_934);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6713(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_935 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_934);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6714(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_934 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1473);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6716(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_933 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_931);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6717(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_932 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_931);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6718(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_931 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1063);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6720(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_930 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_928);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6721(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_929 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_928);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6722(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_928 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1472);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6724(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_927 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_925);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6725(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_926 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_925);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6726(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_925 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1053);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6728(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_924 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_922);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6729(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_923 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_922);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6730(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_922 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1069);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6733(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_921 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_920);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6734(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_920 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1484);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6737(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_919 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_918);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6738(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_918 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1482);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6745(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_917 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_916);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6747(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_916 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1394);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6749(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_915 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_914);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6751(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_914 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1390);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6753(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_913 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_912);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6755(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_912 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1386);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6757(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_911 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_910);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6759(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_910 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1475);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6949(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_909 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_908);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6950(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_908 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1483);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6953(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_907 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_906);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs6954(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_906 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1481);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7097(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_905 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_904);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7098(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_904 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1082);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7101(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_903 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_902);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7102(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_902 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1080);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7105(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_901 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_900);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7106(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_900 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1081);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7108(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_899 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_898);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7110(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_898 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1083);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7112(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_897 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_896);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7114(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_896 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1098);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7116(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_895 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_894);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7118(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_894 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1097);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7145(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_893 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_891);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7146(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_892 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_891);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7147(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_891 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1092);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7150(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_890 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_888);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7151(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_889 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_888);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7152(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_888 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1093);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7155(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_887 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_885);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7156(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_886 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_885);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7157(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_885 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1093);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7160(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_884 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_882);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7161(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_883 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_882);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7162(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_882 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1092);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7165(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_881 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_879);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7166(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_880 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_879);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7167(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_879 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1091);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7170(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_878 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_876);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7171(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_877 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_876);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7172(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_876 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1091);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7175(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_875 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_873);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7176(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_874 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_873);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7177(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_873 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1090);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7180(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_872 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_870);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7181(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_871 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_870);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7182(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_870 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1090);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7185(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_869 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_867);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7186(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_868 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_867);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7187(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_867 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1089);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7190(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_866 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_864);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7191(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_865 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_864);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7192(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_864 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1089);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7195(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_863 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_861);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7196(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_862 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_861);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7197(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_861 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1088);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7200(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_860 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_858);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7201(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_859 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_858);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7202(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_858 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1088);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7205(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_857 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_855);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7206(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_856 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_855);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7207(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_855 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1087);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7210(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_854 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_852);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7211(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_853 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_852);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7212(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_852 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1087);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7215(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_851 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_849);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7216(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_850 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_849);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7217(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_849 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1086);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7220(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_848 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_846);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7221(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_847 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_846);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7222(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_846 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1086);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7225(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_845 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_843);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7226(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_844 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_843);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7227(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_843 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1078);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7230(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_842 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_840);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7231(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_841 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_840);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7232(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_840 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1078);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7235(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_839 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_837);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7236(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_838 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_837);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7237(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_837 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1077);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7240(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_836 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_834);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7241(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_835 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_834);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7242(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_834 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1077);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7245(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_833 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_831);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7246(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_832 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_831);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7247(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_831 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1076);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7250(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_830 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_828);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7251(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_829 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_828);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7252(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_828 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1076);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7255(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_827 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_825);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7256(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_826 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_825);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7257(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_825 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1075);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7260(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_824 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_822);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7261(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_823 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_822);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7262(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_822 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1075);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7265(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_821 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_819);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7266(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_820 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_819);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7267(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_819 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1074);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7270(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_818 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_816);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7271(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_817 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_816);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7272(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_816 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1074);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7285(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_815 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_813);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7286(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_814 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_813);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7287(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_813 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1079);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7290(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_812 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_810);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7291(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_811 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_810);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7292(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_810 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1286);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7295(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_809 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_807);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7296(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_808 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_807);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7297(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_807 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1259);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7300(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_806 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_804);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7301(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_805 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_804);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7302(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_804 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1258);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7305(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_803 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_801);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7306(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_802 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_801);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7307(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_801 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1260);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7310(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_800 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_798);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7311(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_799 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_798);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7312(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_798 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1285);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7315(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_797 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_795);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7316(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_796 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_795);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7317(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_795 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1079);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7330(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_794 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_793);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7332(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_793 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1122);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7360(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_792 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_791);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7362(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_791 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1143);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7365(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_790 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_789);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7367(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_789 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1231);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7395(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_788 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_787);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7397(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_787 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1288);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7400(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_786 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_785);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7402(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_785 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1289);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7405(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_784 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_783);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7407(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_783 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1290);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7410(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_782 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_781);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7412(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_781 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1265);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7415(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_780 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_779);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7417(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_779 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1287);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7420(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_778 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_777);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7422(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_777 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1264);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7425(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_776 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_775);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7427(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_775 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1262);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7430(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_774 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_773);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7432(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_773 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1261);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7435(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_772 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_771);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7437(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_771 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1263);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7440(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_770 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_769);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7442(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_769 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1068);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7445(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_768 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_769);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7455(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_767 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_766);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7457(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_766 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1187);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7464(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_765 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_763);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7465(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_764 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_763);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7466(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_763 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1094);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7520(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_762 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_760);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7521(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_761 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_760);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7522(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_760 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1094);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7524(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_759 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_758);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7526(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_758 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1040);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7528(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_757 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_756);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7530(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_756 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1035);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7532(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_755 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_753);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7533(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_754 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_753);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7534(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_753 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1070);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7536(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_752 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_750);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7537(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_751 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_750);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7538(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_750 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1070);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7540(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_749 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_747);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7541(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_748 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_747);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7542(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_747 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1029);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7544(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_746 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_744);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7545(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_745 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_744);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7546(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_744 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1027);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7548(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_743 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_741);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7549(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_742 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_741);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7550(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_741 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1021);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7552(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_740 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_738);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7553(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_739 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_738);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7554(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_738 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1029);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7556(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_737 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_735);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7557(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_736 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_735);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7558(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_735 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1027);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7560(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_734 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_732);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7561(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_733 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_732);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7562(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_732 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1024);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7564(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_731 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_729);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7565(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_730 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_729);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7566(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_729 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1033);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7568(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_728 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_726);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7569(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_727 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_726);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7570(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_726 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1048);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7572(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_725 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_723);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7573(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_724 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_723);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7574(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_723 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1043);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7576(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_722 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_720);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7577(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_721 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_720);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7578(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_720 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1038);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7580(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_719 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_718);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7582(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_718 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1000);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7584(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_717 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_716);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7586(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_716 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_997);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7588(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_715 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_714);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7590(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_714 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_994);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7592(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_713 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_712);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7594(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_712 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_991);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7596(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_711 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_710);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7598(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_710 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_988);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7600(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_709 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_708);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7602(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_708 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_985);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7604(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_707 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_706);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7606(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_706 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1015);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7608(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_705 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_704);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7610(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_704 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1012);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7612(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_703 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_702);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7614(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_702 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1924);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7616(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_701 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_699);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7617(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_700 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_699);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7618(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_699 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2090);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7620(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_698 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_696);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7621(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_697 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_696);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7622(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_696 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1555);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7624(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_695 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_693);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7625(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_694 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_693);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7626(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_693 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1865);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7628(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_692 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_690);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7629(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_691 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_690);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7630(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_690 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2251);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7632(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_689 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_687);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7633(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_688 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_687);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7634(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_687 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2199);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7636(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_686 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_684);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7637(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_685 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_684);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7638(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_684 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2300);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7640(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_683 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_681);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7641(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_682 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_681);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7642(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_681 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1687);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7644(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_680 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_678);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7645(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_679 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_678);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7646(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_678 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2147);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7648(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_677 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_675);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7649(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_676 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_675);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7650(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_675 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1748);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7652(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_674 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_672);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7653(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_673 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_672);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7654(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_672 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2037);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7656(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_671 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_669);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7657(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_670 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_669);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7658(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_669 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1812);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7660(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_668 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1066);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7662(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1066 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2339);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7664(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_667 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_665);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7665(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_666 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_665);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7666(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_665 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1188);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7668(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_664 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_662);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7669(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_663 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_662);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7670(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_662 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1974);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7672(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_661 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_659);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7673(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_660 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_659);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7674(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_659 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1395);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7676(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_658 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_656);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7677(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_657 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_656);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7678(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_656 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2339);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7680(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_655 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_654);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7682(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_654 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1004);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7684(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_653 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_651);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7685(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_652 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_651);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7686(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_651 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2352);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7688(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_650 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_649);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7690(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_649 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1479);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7692(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_648 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_647);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7694(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_647 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1480);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7696(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_646 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_645);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7698(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_645 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1003);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7700(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_644 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_643);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7702(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_643 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1009);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7704(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_642 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_641);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7706(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_641 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1006);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7708(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_640 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_639);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7710(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_639 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1007);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7712(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_638 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_637);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7714(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_637 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1018);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7716(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_636 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_635);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7718(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_635 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1019);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7720(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_634 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_633);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7722(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_633 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_983);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7724(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_632 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_631);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7726(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_631 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1010);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7728(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_630 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_629);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7730(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_629 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_982);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7733(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_628 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_627);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7734(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_627 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1025);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7736(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_626 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_625);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7738(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_625 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_989);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7740(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_624 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1062);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7742(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1062 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1393);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7744(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_623 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_622);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7746(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_622 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_986);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7748(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_621 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_620);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7750(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_620 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_992);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7752(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_619 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_618);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7754(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_618 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1001);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7757(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_617 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_616);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7758(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_616 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1022);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7761(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_615 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_614);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7762(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_614 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_971);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7764(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_613 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_612);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7766(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_612 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_995);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7769(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_611 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_610);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7770(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_610 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_974);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7772(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_609 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1063);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7774(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1063 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1474);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7776(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_608 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1060);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7778(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1060 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1385);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7780(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_607 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_606);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7782(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_606 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1013);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7784(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_605 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1061);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7786(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1061 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1389);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7788(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_604 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_603);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7790(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_603 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_998);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7792(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_602 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_601);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7794(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_601 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1016);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7797(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_600 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_599);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7798(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_599 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1477);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7801(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_598 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1064);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7802(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1064 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1479);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7805(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_597 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1056);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7806(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1056 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_966);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7809(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_596 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1065);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7810(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1065 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1480);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7813(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_595 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1059);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7814(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1059 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_968);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7816(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_594 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_593);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7818(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_593 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1067);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7820(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_592 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_590);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7821(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_591 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_590);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7822(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_590 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1286);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7824(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_589 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_587);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7825(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_588 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_587);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7826(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_587 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1258);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7828(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_586 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_584);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7829(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_585 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_584);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7830(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_584 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1285);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7832(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_583 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_581);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7833(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_582 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_581);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7834(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_581 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1259);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7836(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_580 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_578);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7837(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_579 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_578);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7838(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_578 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1260);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7841(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_577 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_576);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7842(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_576 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_884);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7845(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_575 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_574);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7846(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_574 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_860);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7848(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_573 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_571);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7849(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_572 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_571);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7850(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_571 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1031);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7853(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_570 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_569);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7854(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_569 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_815);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7857(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_568 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_567);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7858(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_567 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_857);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7861(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_566 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_565);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7862(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_565 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_812);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7865(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_564 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_563);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7866(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_563 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_809);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7869(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_562 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_561);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7870(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_561 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_881);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7873(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_560 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_559);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7874(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_559 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_854);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7877(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_558 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_557);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7878(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_557 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_806);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7881(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_556 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_555);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7882(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_555 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_803);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7885(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_554 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_553);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7886(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_553 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_851);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7889(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_552 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_551);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7890(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_551 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_800);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7893(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_550 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_549);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7894(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_549 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_893);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7897(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_548 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_547);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7898(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_547 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_878);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7901(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_546 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_545);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7902(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_545 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_848);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7905(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_544 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_543);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7906(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_543 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_845);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7909(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_542 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_541);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7910(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_541 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_875);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7913(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_540 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_539);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7914(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_539 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_842);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7917(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_538 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_537);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7918(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_537 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_839);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7921(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_536 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_535);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7922(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_535 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_890);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7925(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_534 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_533);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7926(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_533 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_872);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7929(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_532 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_531);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7930(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_531 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_836);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7933(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_530 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_529);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7934(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_529 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_833);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7937(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_528 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_527);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7938(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_527 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_869);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7941(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_526 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_525);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7942(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_525 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_830);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7945(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_524 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_523);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7946(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_523 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_827);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7949(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_522 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_521);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7950(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_521 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_866);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7953(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_520 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_519);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7954(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_519 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_824);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7957(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_518 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_517);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7958(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_517 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_821);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7961(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_516 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_515);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7962(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_515 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_887);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7965(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_514 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_513);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7966(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_513 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_818);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7969(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_512 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_511);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7970(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_511 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_863);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7972(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_510 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_508);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7973(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_509 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_508);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7974(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_508 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1032);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7976(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_507 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_506);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7978(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_506 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_796);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7980(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_505 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_503);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7981(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_504 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_503);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7982(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_503 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1122);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7984(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_502 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_500);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7985(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_501 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_500);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7986(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_500 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1032);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7988(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_499 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_497);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7989(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_498 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_497);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7990(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_497 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1031);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7992(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_496 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_494);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7993(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_495 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_494);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7994(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_494 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_862);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7996(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_493 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_491);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7997(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_492 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_491);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs7998(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_491 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_814);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8000(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_490 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_488);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8001(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_489 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_488);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8002(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_488 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_859);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8004(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_487 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_485);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8005(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_486 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_485);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8006(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_485 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_886);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8008(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_484 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_482);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8009(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_483 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_482);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8010(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_482 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_856);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8012(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_481 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_479);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8013(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_480 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_479);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8014(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_479 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_853);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8016(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_478 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_476);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8017(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_477 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_476);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8018(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_476 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_883);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8020(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_475 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_473);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8021(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_474 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_473);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8022(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_473 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_797);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8024(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_472 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_470);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8025(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_471 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_470);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8026(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_470 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_850);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8028(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_469 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_467);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8029(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_468 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_467);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8030(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_467 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_847);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8032(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_466 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_464);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8033(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_465 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_464);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8034(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_464 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_880);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8036(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_463 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_461);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8037(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_462 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_461);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8038(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_461 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_844);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8040(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_460 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_458);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8041(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_459 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_458);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8042(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_458 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_841);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8044(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_457 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_455);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8045(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_456 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_455);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8046(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_455 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_877);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8048(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_454 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_452);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8049(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_453 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_452);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8050(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_452 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_838);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8052(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_451 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_449);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8053(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_450 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_449);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8054(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_449 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_835);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8056(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_448 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_446);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8057(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_447 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_446);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8058(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_446 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_874);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8060(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_445 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_443);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8061(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_444 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_443);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8062(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_443 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_832);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8064(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_442 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_440);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8065(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_441 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_440);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8066(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_440 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_871);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8068(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_439 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_437);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8069(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_438 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_437);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8070(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_437 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_829);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8072(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_436 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_434);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8073(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_435 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_434);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8074(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_434 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_892);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8076(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_433 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_431);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8077(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_432 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_431);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8078(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_431 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_826);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8080(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_430 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_428);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8081(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_429 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_428);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8082(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_428 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_868);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8084(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_427 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_425);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8085(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_426 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_425);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8086(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_425 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_823);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8088(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_424 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_422);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8089(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_423 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_422);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8090(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_422 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_889);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8092(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_421 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_419);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8093(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_420 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_419);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8094(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_419 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_820);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8096(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_418 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_416);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8097(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_417 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_416);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8098(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_416 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_865);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8100(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_415 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_413);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8101(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_414 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_413);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8102(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_413 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_817);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8104(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_412 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_410);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8105(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_411 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_410);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8106(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_410 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1260);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8108(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_409 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_407);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8109(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_408 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_407);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8110(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_407 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_811);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8112(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_406 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_404);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8113(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_405 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_404);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8114(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_404 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_808);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8116(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_403 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_401);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8117(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_402 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_401);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8118(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_401 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1259);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8120(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_400 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_398);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8121(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_399 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_398);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8122(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_398 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_805);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8124(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_397 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_395);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8125(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_396 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_395);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8126(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_395 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_802);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8128(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_394 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_392);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8129(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_393 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_392);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8130(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_392 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_799);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8132(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_391 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_389);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8133(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_390 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_389);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8134(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_389 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1285);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8136(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_388 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_386);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8137(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_387 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_386);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8138(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_386 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1286);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8140(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_385 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_383);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8141(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_384 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_383);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8142(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_383 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1258);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8144(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_382 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_380);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8145(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_381 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_380);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8146(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_380 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1143);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8148(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_379 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_377);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8149(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_378 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_377);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8150(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_377 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_794);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8152(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_376 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_374);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8153(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_375 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_374);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8154(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_374 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1231);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8156(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_373 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_371);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8157(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_372 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_371);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8158(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_371 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1288);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8160(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_370 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_368);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8161(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_369 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_368);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8162(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_368 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1289);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8164(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_367 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_365);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8165(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_366 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_365);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8166(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_365 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1290);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8168(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_364 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_362);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8169(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_363 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_362);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8170(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_362 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1265);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8172(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_361 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_359);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8173(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_360 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_359);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8174(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_359 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_782);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8176(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_358 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_356);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8177(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_357 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_356);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8178(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_356 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_790);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8180(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_355 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_353);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8181(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_354 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_353);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8182(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_353 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_782);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8184(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_352 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_350);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8185(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_351 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_350);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8186(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_350 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1122);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8188(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_349 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_347);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8189(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_348 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_347);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8190(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_347 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1290);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8192(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_346 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_344);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8193(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_345 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_344);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8194(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_344 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1143);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8196(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_343 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_341);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8197(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_342 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_341);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8198(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_341 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_794);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8200(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_340 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_338);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8201(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_339 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_338);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8202(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_338 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_780);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8204(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_337 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_335);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8205(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_336 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_335);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8206(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_335 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1231);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8208(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_334 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_332);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8209(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_333 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_332);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8210(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_332 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1288);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8212(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_331 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_329);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8213(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_330 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_329);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8214(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_329 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1289);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8216(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_328 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_326);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8217(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_327 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_326);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8218(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_326 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1264);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8220(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_325 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_323);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8221(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_324 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_323);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8222(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_323 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_788);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8224(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_322 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_320);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8225(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_321 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_320);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8226(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_320 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1265);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8228(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_319 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_317);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8229(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_318 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_317);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8230(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_317 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_792);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8232(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_316 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_314);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8233(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_315 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_314);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8234(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_314 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_792);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8236(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_313 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_311);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8237(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_312 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_311);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8238(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_311 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_790);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8240(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_310 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_308);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8241(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_309 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_308);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8242(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_308 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1287);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8244(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_307 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_305);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8245(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_306 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_305);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8246(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_305 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1287);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8248(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_304 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_302);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8249(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_303 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_302);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8250(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_302 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_784);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8252(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_301 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_299);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8253(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_300 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_299);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8254(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_299 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1264);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8256(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_298 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_296);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8257(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_297 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_296);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8258(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_296 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1262);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8260(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_295 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_293);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8261(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_294 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_293);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8262(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_293 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_772);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8264(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_292 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_290);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8265(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_291 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_290);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8266(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_290 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1262);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8268(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_289 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_287);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8269(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_288 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_287);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8270(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_287 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_776);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8272(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_286 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_284);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8273(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_285 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_284);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8274(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_284 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1261);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8276(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_283 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_281);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8277(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_282 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_281);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8278(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_281 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1263);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8280(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_280 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_278);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8281(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_279 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_278);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8282(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_278 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1263);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8284(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_277 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_275);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8285(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_276 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_275);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8286(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_275 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_788);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8288(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_274 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_272);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8289(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_273 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_272);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8290(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_272 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_786);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8292(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_271 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_269);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8293(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_270 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_269);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8294(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_269 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_786);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8296(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_268 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_266);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8297(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_267 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_266);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8298(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_266 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_784);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8300(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_265 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_263);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8301(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_264 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_263);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8302(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_263 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1261);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8304(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_262 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_260);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8305(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_261 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_260);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8306(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_260 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_778);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8308(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_259 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_257);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8309(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_258 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_257);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8310(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_257 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_774);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8312(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_256 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_254);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8313(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_255 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_254);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8314(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_254 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_772);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8316(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_253 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_251);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8317(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_252 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_251);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8318(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_251 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_776);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8320(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_250 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_248);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8321(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_249 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_248);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8322(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_248 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_774);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8324(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_247 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_245);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8325(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_246 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_245);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8326(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_245 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_780);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8328(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_244 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_242);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8329(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_243 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_242);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8330(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_242 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_778);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8332(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_241 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_239);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8333(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_240 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_239);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8334(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_239 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_770);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8336(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_238 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_236);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8337(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_237 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_236);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8338(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_236 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_770);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8340(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_235 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_233);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8341(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_234 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_233);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8342(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_233 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_768);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8344(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_232 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_230);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8345(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_231 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_230);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8346(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_230 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_764);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8348(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_229 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_227);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8349(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_228 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_227);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8350(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_227 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1051);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8352(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_226 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_224);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8353(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_225 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_224);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8354(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_224 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_768);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8356(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_223 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_221);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8357(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_222 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_221);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8358(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_221 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_767);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8360(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_220 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_218);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8361(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_219 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_218);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8362(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_218 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1187);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8364(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_217 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_215);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8365(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_216 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_215);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8366(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_215 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_767);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8368(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_214 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_212);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8369(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_213 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_212);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8370(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_212 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1187);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8373(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_211 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_210);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8374(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_210 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1044);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8377(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_209 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_208);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8378(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_208 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1052);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8381(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_207 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_206);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8382(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_206 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1049);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8385(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_205 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_204);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8386(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_204 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1050);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8389(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_203 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_202);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8390(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_202 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1041);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8393(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_201 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_200);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8394(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_200 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1037);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8397(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_199 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_198);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8398(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_198 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1046);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8401(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_197 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_196);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8402(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_196 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1045);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8405(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_195 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_194);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8406(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_194 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1036);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8409(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_193 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_192);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8410(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_192 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1052);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8412(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_191 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_190);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8414(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_190 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_765);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8416(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_189 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_188);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8418(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_188 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_761);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8420(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_187 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_186);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8422(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_186 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_762);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8425(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_185 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1055);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8426(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1055 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1047);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8429(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_184 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1058);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8430(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1058 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1051);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8433(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_183 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1057);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8434(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1057 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1034);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8436(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_182 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_180);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8437(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_181 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_180);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8438(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_180 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1042);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8441(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_179 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1054);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8442(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1054 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1039);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8444(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_178 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_177);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8446(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_177 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1040);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8448(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_176 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_175);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8450(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_175 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1041);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8452(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_174 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_173);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8454(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_173 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1035);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8456(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_172 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_171);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8458(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_171 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1044);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8460(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_170 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_169);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8462(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_169 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1049);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8464(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_168 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_167);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8466(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_167 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1050);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8468(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_166 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_165);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8470(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_165 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1039);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8472(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_164 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_163);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8474(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_163 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1042);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8476(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_162 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_161);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8478(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_161 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1045);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8480(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_160 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_159);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8482(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_159 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1037);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8484(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_158 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_157);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8486(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_157 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1034);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8488(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_156 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_155);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8490(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_155 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1046);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8492(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_154 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_153);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8494(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_153 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1036);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8496(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_152 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_151);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8498(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_151 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1047);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8500(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_150 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_149);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8502(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_149 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_754);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8504(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_148 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_147);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8506(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_147 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_752);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8508(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_146 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_145);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8510(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_145 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_592);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8512(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_144 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_143);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8514(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_143 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_589);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8516(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_142 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_141);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8518(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_141 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_583);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8520(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_140 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_139);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8522(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_139 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_580);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8524(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_138 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_137);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8526(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_137 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_586);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8528(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_136 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_134);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8529(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_135 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_134);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8530(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_134 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_818);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8532(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_133 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_131);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8533(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_132 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_131);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8534(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_131 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_887);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8536(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_130 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_128);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8537(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_129 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_128);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8538(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_128 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_821);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8540(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_127 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_125);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8541(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_126 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_125);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8542(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_125 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_824);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8544(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_124 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_122);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8545(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_123 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_122);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8546(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_122 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_866);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8548(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_121 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_120);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8550(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_120 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_510);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8552(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_119 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_117);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8553(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_118 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_117);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8554(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_117 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_830);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8556(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_116 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_114);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8557(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_115 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_114);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8558(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_114 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_869);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8560(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_113 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_111);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8561(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_112 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_111);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8562(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_111 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_833);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8564(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_110 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_108);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8565(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_109 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_108);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8566(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_108 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_836);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8568(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_107 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_105);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8569(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_106 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_105);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8570(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_105 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_872);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8572(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_104 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_102);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8573(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_103 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_102);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8574(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_102 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_890);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8576(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_101 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_99);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8577(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_100 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_99);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8578(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_99 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_839);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8580(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_98 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_96);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8581(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_97 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_96);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8582(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_96 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_842);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8584(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_95 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_93);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8585(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_94 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_93);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8586(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_93 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_875);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8588(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_92 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_90);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8589(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_91 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_90);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8590(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_90 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_845);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8592(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_89 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_87);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8593(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_88 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_87);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8594(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_87 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_848);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8596(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_86 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_85);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8598(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_85 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_573);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8600(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_84 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_82);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8601(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_83 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_82);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8602(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_82 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_893);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8604(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_81 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_79);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8605(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_80 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_79);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8606(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_79 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_800);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8608(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_78 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_77);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8610(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_77 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_803);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8612(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_76 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_74);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8613(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_75 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_74);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8614(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_74 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_827);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8616(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_73 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_71);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8617(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_72 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_71);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8618(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_71 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_806);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8620(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_70 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_68);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8621(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_69 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_68);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8622(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_68 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_854);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8624(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_67 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_65);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8625(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_66 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_65);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8626(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_65 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_881);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8628(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_64 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_62);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8629(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_63 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_62);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8630(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_62 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_809);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8632(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_61 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_59);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8633(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_60 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_59);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8634(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_59 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_812);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8636(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_58 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_56);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8637(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_57 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_56);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8638(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_56 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_878);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8640(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_55 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_53);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8641(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_54 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_53);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8642(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_53 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_851);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8644(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_52 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_50);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8645(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_51 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_50);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8646(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_50 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_815);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8648(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_49 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_47);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8649(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_48 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_47);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8650(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_47 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_860);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8652(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_46 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_44);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8653(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_45 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_44);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8654(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_44 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_884);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8656(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_43 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_41);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8657(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_42 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_41);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8658(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_41 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_857);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8660(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_40 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_38);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8661(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_39 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_38);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8662(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_38 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_863);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8664(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_37 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_35);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8665(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_36 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_35);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8666(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_35 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_796);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8669(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_34 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_33);
  not mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_drc_bufs8670(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_33 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_504);
  xor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g2(n_143 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2621 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2581);
  xor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g8672(n_142 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2619 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2610);
  xor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g8673(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_30 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2093 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2109);
  xor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g8674(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_29 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2048 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2053);
  xor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g8675(out1[1] ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1743 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1723);
  xor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g8676(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_27 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1721 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1739);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g8677(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_26 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_77 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_702);
  and mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g8678(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_25 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_208 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_599);
  xor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g8679(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_24 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_593 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1844);
  xor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g8680(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_23 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2390 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_210);
  xor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g8681(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_22 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1493 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_206);
  xor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g8682(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_21 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2393 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_204);
  xor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g8683(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_20 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1695 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_202);
  xor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g8684(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_19 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1492 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_200);
  xor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g8685(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_18 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1494 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_198);
  xor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g8686(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_17 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1693 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_196);
  xor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g8687(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_16 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1691 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_194);
  xor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g8688(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_15 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1689 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_192);
  xor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g8689(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_14 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_177 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1730);
  xor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g8690(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_13 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_175 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1793);
  xor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g8691(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_12 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_173 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1729);
  xor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g8692(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_11 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_171 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1699);
  xor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g8693(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_10 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_169 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2013);
  xor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g8694(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_9 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_167 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2423);
  xor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g8695(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_8 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_165 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1902);
  xor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g8696(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_7 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_163 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2280);
  xor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g8697(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_6 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_161 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1728);
  xor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g8698(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_5 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_159 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2281);
  xor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g8699(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_4 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_157 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1899);
  xor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g8700(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_3 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_155 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1796);
  xor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g8701(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_2 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_153 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1794);
  xor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g8702(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_151 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1845);
  xor mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_g8703(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_0 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1053 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1560);
  buf g8704(n_133 ,n_117);
  buf g8705(n_123 ,n_114);
  buf g8706(mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1218 ,mul_9_28_Y_mul_9_40_Y_mul_10_28_Y_mul_10_40_n_1144);
endmodule
