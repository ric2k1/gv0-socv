module top(in1, in2, in3, in4, out1);
  input [15:0] in1, in2, in3, in4;
  output [33:0] out1;
  wire [15:0] in1, in2, in3, in4;
  wire [33:0] out1;
  wire csa_tree_add_7_45_groupi_n_0, csa_tree_add_7_45_groupi_n_1, csa_tree_add_7_45_groupi_n_2, csa_tree_add_7_45_groupi_n_3, csa_tree_add_7_45_groupi_n_4, csa_tree_add_7_45_groupi_n_5, csa_tree_add_7_45_groupi_n_6, csa_tree_add_7_45_groupi_n_7;
  wire csa_tree_add_7_45_groupi_n_8, csa_tree_add_7_45_groupi_n_9, csa_tree_add_7_45_groupi_n_10, csa_tree_add_7_45_groupi_n_21, csa_tree_add_7_45_groupi_n_22, csa_tree_add_7_45_groupi_n_23, csa_tree_add_7_45_groupi_n_24, csa_tree_add_7_45_groupi_n_25;
  wire csa_tree_add_7_45_groupi_n_26, csa_tree_add_7_45_groupi_n_27, csa_tree_add_7_45_groupi_n_28, csa_tree_add_7_45_groupi_n_29, csa_tree_add_7_45_groupi_n_30, csa_tree_add_7_45_groupi_n_31, csa_tree_add_7_45_groupi_n_32, csa_tree_add_7_45_groupi_n_33;
  wire csa_tree_add_7_45_groupi_n_34, csa_tree_add_7_45_groupi_n_35, csa_tree_add_7_45_groupi_n_36, csa_tree_add_7_45_groupi_n_37, csa_tree_add_7_45_groupi_n_38, csa_tree_add_7_45_groupi_n_39, csa_tree_add_7_45_groupi_n_40, csa_tree_add_7_45_groupi_n_41;
  wire csa_tree_add_7_45_groupi_n_42, csa_tree_add_7_45_groupi_n_43, csa_tree_add_7_45_groupi_n_44, csa_tree_add_7_45_groupi_n_45, csa_tree_add_7_45_groupi_n_46, csa_tree_add_7_45_groupi_n_47, csa_tree_add_7_45_groupi_n_48, csa_tree_add_7_45_groupi_n_49;
  wire csa_tree_add_7_45_groupi_n_50, csa_tree_add_7_45_groupi_n_51, csa_tree_add_7_45_groupi_n_52, csa_tree_add_7_45_groupi_n_53, csa_tree_add_7_45_groupi_n_54, csa_tree_add_7_45_groupi_n_55, csa_tree_add_7_45_groupi_n_56, csa_tree_add_7_45_groupi_n_57;
  wire csa_tree_add_7_45_groupi_n_58, csa_tree_add_7_45_groupi_n_59, csa_tree_add_7_45_groupi_n_60, csa_tree_add_7_45_groupi_n_61, csa_tree_add_7_45_groupi_n_62, csa_tree_add_7_45_groupi_n_63, csa_tree_add_7_45_groupi_n_64, csa_tree_add_7_45_groupi_n_65;
  wire csa_tree_add_7_45_groupi_n_66, csa_tree_add_7_45_groupi_n_67, csa_tree_add_7_45_groupi_n_68, csa_tree_add_7_45_groupi_n_69, csa_tree_add_7_45_groupi_n_70, csa_tree_add_7_45_groupi_n_71, csa_tree_add_7_45_groupi_n_72, csa_tree_add_7_45_groupi_n_73;
  wire csa_tree_add_7_45_groupi_n_74, csa_tree_add_7_45_groupi_n_75, csa_tree_add_7_45_groupi_n_76, csa_tree_add_7_45_groupi_n_77, csa_tree_add_7_45_groupi_n_78, csa_tree_add_7_45_groupi_n_79, csa_tree_add_7_45_groupi_n_80, csa_tree_add_7_45_groupi_n_81;
  wire csa_tree_add_7_45_groupi_n_82, csa_tree_add_7_45_groupi_n_83, csa_tree_add_7_45_groupi_n_84, csa_tree_add_7_45_groupi_n_85, csa_tree_add_7_45_groupi_n_86, csa_tree_add_7_45_groupi_n_87, csa_tree_add_7_45_groupi_n_88, csa_tree_add_7_45_groupi_n_89;
  wire csa_tree_add_7_45_groupi_n_90, csa_tree_add_7_45_groupi_n_91, csa_tree_add_7_45_groupi_n_92, csa_tree_add_7_45_groupi_n_93, csa_tree_add_7_45_groupi_n_94, csa_tree_add_7_45_groupi_n_95, csa_tree_add_7_45_groupi_n_96, csa_tree_add_7_45_groupi_n_97;
  wire csa_tree_add_7_45_groupi_n_98, csa_tree_add_7_45_groupi_n_99, csa_tree_add_7_45_groupi_n_100, csa_tree_add_7_45_groupi_n_101, csa_tree_add_7_45_groupi_n_102, csa_tree_add_7_45_groupi_n_103, csa_tree_add_7_45_groupi_n_104, csa_tree_add_7_45_groupi_n_105;
  wire csa_tree_add_7_45_groupi_n_106, csa_tree_add_7_45_groupi_n_107, csa_tree_add_7_45_groupi_n_108, csa_tree_add_7_45_groupi_n_109, csa_tree_add_7_45_groupi_n_110, csa_tree_add_7_45_groupi_n_111, csa_tree_add_7_45_groupi_n_112, csa_tree_add_7_45_groupi_n_113;
  wire csa_tree_add_7_45_groupi_n_114, csa_tree_add_7_45_groupi_n_115, csa_tree_add_7_45_groupi_n_116, csa_tree_add_7_45_groupi_n_117, csa_tree_add_7_45_groupi_n_118, csa_tree_add_7_45_groupi_n_119, csa_tree_add_7_45_groupi_n_120, csa_tree_add_7_45_groupi_n_121;
  wire csa_tree_add_7_45_groupi_n_122, csa_tree_add_7_45_groupi_n_123, csa_tree_add_7_45_groupi_n_124, csa_tree_add_7_45_groupi_n_125, csa_tree_add_7_45_groupi_n_126, csa_tree_add_7_45_groupi_n_127, csa_tree_add_7_45_groupi_n_128, csa_tree_add_7_45_groupi_n_129;
  wire csa_tree_add_7_45_groupi_n_130, csa_tree_add_7_45_groupi_n_131, csa_tree_add_7_45_groupi_n_132, csa_tree_add_7_45_groupi_n_133, csa_tree_add_7_45_groupi_n_134, csa_tree_add_7_45_groupi_n_135, csa_tree_add_7_45_groupi_n_136, csa_tree_add_7_45_groupi_n_137;
  wire csa_tree_add_7_45_groupi_n_138, csa_tree_add_7_45_groupi_n_139, csa_tree_add_7_45_groupi_n_140, csa_tree_add_7_45_groupi_n_141, csa_tree_add_7_45_groupi_n_142, csa_tree_add_7_45_groupi_n_143, csa_tree_add_7_45_groupi_n_144, csa_tree_add_7_45_groupi_n_145;
  wire csa_tree_add_7_45_groupi_n_146, csa_tree_add_7_45_groupi_n_147, csa_tree_add_7_45_groupi_n_148, csa_tree_add_7_45_groupi_n_149, csa_tree_add_7_45_groupi_n_150, csa_tree_add_7_45_groupi_n_151, csa_tree_add_7_45_groupi_n_152, csa_tree_add_7_45_groupi_n_153;
  wire csa_tree_add_7_45_groupi_n_154, csa_tree_add_7_45_groupi_n_155, csa_tree_add_7_45_groupi_n_156, csa_tree_add_7_45_groupi_n_157, csa_tree_add_7_45_groupi_n_158, csa_tree_add_7_45_groupi_n_159, csa_tree_add_7_45_groupi_n_160, csa_tree_add_7_45_groupi_n_161;
  wire csa_tree_add_7_45_groupi_n_162, csa_tree_add_7_45_groupi_n_163, csa_tree_add_7_45_groupi_n_164, csa_tree_add_7_45_groupi_n_165, csa_tree_add_7_45_groupi_n_166, csa_tree_add_7_45_groupi_n_167, csa_tree_add_7_45_groupi_n_168, csa_tree_add_7_45_groupi_n_169;
  wire csa_tree_add_7_45_groupi_n_170, csa_tree_add_7_45_groupi_n_171, csa_tree_add_7_45_groupi_n_172, csa_tree_add_7_45_groupi_n_173, csa_tree_add_7_45_groupi_n_174, csa_tree_add_7_45_groupi_n_175, csa_tree_add_7_45_groupi_n_176, csa_tree_add_7_45_groupi_n_177;
  wire csa_tree_add_7_45_groupi_n_178, csa_tree_add_7_45_groupi_n_179, csa_tree_add_7_45_groupi_n_180, csa_tree_add_7_45_groupi_n_181, csa_tree_add_7_45_groupi_n_182, csa_tree_add_7_45_groupi_n_183, csa_tree_add_7_45_groupi_n_184, csa_tree_add_7_45_groupi_n_185;
  wire csa_tree_add_7_45_groupi_n_186, csa_tree_add_7_45_groupi_n_187, csa_tree_add_7_45_groupi_n_188, csa_tree_add_7_45_groupi_n_189, csa_tree_add_7_45_groupi_n_190, csa_tree_add_7_45_groupi_n_191, csa_tree_add_7_45_groupi_n_192, csa_tree_add_7_45_groupi_n_193;
  wire csa_tree_add_7_45_groupi_n_194, csa_tree_add_7_45_groupi_n_195, csa_tree_add_7_45_groupi_n_196, csa_tree_add_7_45_groupi_n_197, csa_tree_add_7_45_groupi_n_198, csa_tree_add_7_45_groupi_n_199, csa_tree_add_7_45_groupi_n_200, csa_tree_add_7_45_groupi_n_201;
  wire csa_tree_add_7_45_groupi_n_202, csa_tree_add_7_45_groupi_n_203, csa_tree_add_7_45_groupi_n_204, csa_tree_add_7_45_groupi_n_205, csa_tree_add_7_45_groupi_n_206, csa_tree_add_7_45_groupi_n_207, csa_tree_add_7_45_groupi_n_208, csa_tree_add_7_45_groupi_n_209;
  wire csa_tree_add_7_45_groupi_n_210, csa_tree_add_7_45_groupi_n_211, csa_tree_add_7_45_groupi_n_212, csa_tree_add_7_45_groupi_n_213, csa_tree_add_7_45_groupi_n_214, csa_tree_add_7_45_groupi_n_215, csa_tree_add_7_45_groupi_n_216, csa_tree_add_7_45_groupi_n_217;
  wire csa_tree_add_7_45_groupi_n_218, csa_tree_add_7_45_groupi_n_219, csa_tree_add_7_45_groupi_n_220, csa_tree_add_7_45_groupi_n_221, csa_tree_add_7_45_groupi_n_222, csa_tree_add_7_45_groupi_n_223, csa_tree_add_7_45_groupi_n_224, csa_tree_add_7_45_groupi_n_225;
  wire csa_tree_add_7_45_groupi_n_226, csa_tree_add_7_45_groupi_n_227, csa_tree_add_7_45_groupi_n_228, csa_tree_add_7_45_groupi_n_229, csa_tree_add_7_45_groupi_n_230, csa_tree_add_7_45_groupi_n_231, csa_tree_add_7_45_groupi_n_232, csa_tree_add_7_45_groupi_n_233;
  wire csa_tree_add_7_45_groupi_n_234, csa_tree_add_7_45_groupi_n_235, csa_tree_add_7_45_groupi_n_236, csa_tree_add_7_45_groupi_n_237, csa_tree_add_7_45_groupi_n_238, csa_tree_add_7_45_groupi_n_239, csa_tree_add_7_45_groupi_n_240, csa_tree_add_7_45_groupi_n_241;
  wire csa_tree_add_7_45_groupi_n_242, csa_tree_add_7_45_groupi_n_243, csa_tree_add_7_45_groupi_n_244, csa_tree_add_7_45_groupi_n_245, csa_tree_add_7_45_groupi_n_246, csa_tree_add_7_45_groupi_n_247, csa_tree_add_7_45_groupi_n_248, csa_tree_add_7_45_groupi_n_249;
  wire csa_tree_add_7_45_groupi_n_250, csa_tree_add_7_45_groupi_n_251, csa_tree_add_7_45_groupi_n_252, csa_tree_add_7_45_groupi_n_253, csa_tree_add_7_45_groupi_n_254, csa_tree_add_7_45_groupi_n_255, csa_tree_add_7_45_groupi_n_256, csa_tree_add_7_45_groupi_n_257;
  wire csa_tree_add_7_45_groupi_n_258, csa_tree_add_7_45_groupi_n_259, csa_tree_add_7_45_groupi_n_260, csa_tree_add_7_45_groupi_n_261, csa_tree_add_7_45_groupi_n_262, csa_tree_add_7_45_groupi_n_263, csa_tree_add_7_45_groupi_n_264, csa_tree_add_7_45_groupi_n_265;
  wire csa_tree_add_7_45_groupi_n_266, csa_tree_add_7_45_groupi_n_267, csa_tree_add_7_45_groupi_n_268, csa_tree_add_7_45_groupi_n_269, csa_tree_add_7_45_groupi_n_270, csa_tree_add_7_45_groupi_n_271, csa_tree_add_7_45_groupi_n_272, csa_tree_add_7_45_groupi_n_273;
  wire csa_tree_add_7_45_groupi_n_274, csa_tree_add_7_45_groupi_n_275, csa_tree_add_7_45_groupi_n_276, csa_tree_add_7_45_groupi_n_277, csa_tree_add_7_45_groupi_n_278, csa_tree_add_7_45_groupi_n_279, csa_tree_add_7_45_groupi_n_280, csa_tree_add_7_45_groupi_n_281;
  wire csa_tree_add_7_45_groupi_n_282, csa_tree_add_7_45_groupi_n_283, csa_tree_add_7_45_groupi_n_284, csa_tree_add_7_45_groupi_n_285, csa_tree_add_7_45_groupi_n_286, csa_tree_add_7_45_groupi_n_287, csa_tree_add_7_45_groupi_n_288, csa_tree_add_7_45_groupi_n_289;
  wire csa_tree_add_7_45_groupi_n_290, csa_tree_add_7_45_groupi_n_291, csa_tree_add_7_45_groupi_n_292, csa_tree_add_7_45_groupi_n_293, csa_tree_add_7_45_groupi_n_294, csa_tree_add_7_45_groupi_n_295, csa_tree_add_7_45_groupi_n_296, csa_tree_add_7_45_groupi_n_297;
  wire csa_tree_add_7_45_groupi_n_298, csa_tree_add_7_45_groupi_n_299, csa_tree_add_7_45_groupi_n_300, csa_tree_add_7_45_groupi_n_301, csa_tree_add_7_45_groupi_n_302, csa_tree_add_7_45_groupi_n_303, csa_tree_add_7_45_groupi_n_304, csa_tree_add_7_45_groupi_n_305;
  wire csa_tree_add_7_45_groupi_n_306, csa_tree_add_7_45_groupi_n_307, csa_tree_add_7_45_groupi_n_308, csa_tree_add_7_45_groupi_n_309, csa_tree_add_7_45_groupi_n_310, csa_tree_add_7_45_groupi_n_311, csa_tree_add_7_45_groupi_n_312, csa_tree_add_7_45_groupi_n_313;
  wire csa_tree_add_7_45_groupi_n_314, csa_tree_add_7_45_groupi_n_315, csa_tree_add_7_45_groupi_n_316, csa_tree_add_7_45_groupi_n_317, csa_tree_add_7_45_groupi_n_318, csa_tree_add_7_45_groupi_n_319, csa_tree_add_7_45_groupi_n_320, csa_tree_add_7_45_groupi_n_321;
  wire csa_tree_add_7_45_groupi_n_322, csa_tree_add_7_45_groupi_n_323, csa_tree_add_7_45_groupi_n_324, csa_tree_add_7_45_groupi_n_325, csa_tree_add_7_45_groupi_n_326, csa_tree_add_7_45_groupi_n_327, csa_tree_add_7_45_groupi_n_328, csa_tree_add_7_45_groupi_n_329;
  wire csa_tree_add_7_45_groupi_n_330, csa_tree_add_7_45_groupi_n_331, csa_tree_add_7_45_groupi_n_332, csa_tree_add_7_45_groupi_n_333, csa_tree_add_7_45_groupi_n_334, csa_tree_add_7_45_groupi_n_335, csa_tree_add_7_45_groupi_n_336, csa_tree_add_7_45_groupi_n_337;
  wire csa_tree_add_7_45_groupi_n_338, csa_tree_add_7_45_groupi_n_339, csa_tree_add_7_45_groupi_n_340, csa_tree_add_7_45_groupi_n_341, csa_tree_add_7_45_groupi_n_342, csa_tree_add_7_45_groupi_n_343, csa_tree_add_7_45_groupi_n_344, csa_tree_add_7_45_groupi_n_345;
  wire csa_tree_add_7_45_groupi_n_346, csa_tree_add_7_45_groupi_n_347, csa_tree_add_7_45_groupi_n_348, csa_tree_add_7_45_groupi_n_349, csa_tree_add_7_45_groupi_n_350, csa_tree_add_7_45_groupi_n_351, csa_tree_add_7_45_groupi_n_352, csa_tree_add_7_45_groupi_n_353;
  wire csa_tree_add_7_45_groupi_n_354, csa_tree_add_7_45_groupi_n_355, csa_tree_add_7_45_groupi_n_356, csa_tree_add_7_45_groupi_n_357, csa_tree_add_7_45_groupi_n_358, csa_tree_add_7_45_groupi_n_359, csa_tree_add_7_45_groupi_n_360, csa_tree_add_7_45_groupi_n_361;
  wire csa_tree_add_7_45_groupi_n_362, csa_tree_add_7_45_groupi_n_363, csa_tree_add_7_45_groupi_n_364, csa_tree_add_7_45_groupi_n_365, csa_tree_add_7_45_groupi_n_366, csa_tree_add_7_45_groupi_n_367, csa_tree_add_7_45_groupi_n_368, csa_tree_add_7_45_groupi_n_369;
  wire csa_tree_add_7_45_groupi_n_370, csa_tree_add_7_45_groupi_n_371, csa_tree_add_7_45_groupi_n_372, csa_tree_add_7_45_groupi_n_373, csa_tree_add_7_45_groupi_n_374, csa_tree_add_7_45_groupi_n_375, csa_tree_add_7_45_groupi_n_376, csa_tree_add_7_45_groupi_n_377;
  wire csa_tree_add_7_45_groupi_n_378, csa_tree_add_7_45_groupi_n_379, csa_tree_add_7_45_groupi_n_380, csa_tree_add_7_45_groupi_n_381, csa_tree_add_7_45_groupi_n_382, csa_tree_add_7_45_groupi_n_383, csa_tree_add_7_45_groupi_n_384, csa_tree_add_7_45_groupi_n_385;
  wire csa_tree_add_7_45_groupi_n_386, csa_tree_add_7_45_groupi_n_387, csa_tree_add_7_45_groupi_n_388, csa_tree_add_7_45_groupi_n_389, csa_tree_add_7_45_groupi_n_390, csa_tree_add_7_45_groupi_n_391, csa_tree_add_7_45_groupi_n_392, csa_tree_add_7_45_groupi_n_393;
  wire csa_tree_add_7_45_groupi_n_394, csa_tree_add_7_45_groupi_n_395, csa_tree_add_7_45_groupi_n_396, csa_tree_add_7_45_groupi_n_397, csa_tree_add_7_45_groupi_n_398, csa_tree_add_7_45_groupi_n_399, csa_tree_add_7_45_groupi_n_400, csa_tree_add_7_45_groupi_n_401;
  wire csa_tree_add_7_45_groupi_n_402, csa_tree_add_7_45_groupi_n_403, csa_tree_add_7_45_groupi_n_404, csa_tree_add_7_45_groupi_n_405, csa_tree_add_7_45_groupi_n_406, csa_tree_add_7_45_groupi_n_407, csa_tree_add_7_45_groupi_n_408, csa_tree_add_7_45_groupi_n_409;
  wire csa_tree_add_7_45_groupi_n_410, csa_tree_add_7_45_groupi_n_411, csa_tree_add_7_45_groupi_n_412, csa_tree_add_7_45_groupi_n_413, csa_tree_add_7_45_groupi_n_414, csa_tree_add_7_45_groupi_n_415, csa_tree_add_7_45_groupi_n_416, csa_tree_add_7_45_groupi_n_417;
  wire csa_tree_add_7_45_groupi_n_418, csa_tree_add_7_45_groupi_n_419, csa_tree_add_7_45_groupi_n_420, csa_tree_add_7_45_groupi_n_421, csa_tree_add_7_45_groupi_n_422, csa_tree_add_7_45_groupi_n_423, csa_tree_add_7_45_groupi_n_424, csa_tree_add_7_45_groupi_n_425;
  wire csa_tree_add_7_45_groupi_n_426, csa_tree_add_7_45_groupi_n_427, csa_tree_add_7_45_groupi_n_428, csa_tree_add_7_45_groupi_n_429, csa_tree_add_7_45_groupi_n_430, csa_tree_add_7_45_groupi_n_431, csa_tree_add_7_45_groupi_n_432, csa_tree_add_7_45_groupi_n_433;
  wire csa_tree_add_7_45_groupi_n_434, csa_tree_add_7_45_groupi_n_435, csa_tree_add_7_45_groupi_n_436, csa_tree_add_7_45_groupi_n_437, csa_tree_add_7_45_groupi_n_438, csa_tree_add_7_45_groupi_n_439, csa_tree_add_7_45_groupi_n_440, csa_tree_add_7_45_groupi_n_441;
  wire csa_tree_add_7_45_groupi_n_442, csa_tree_add_7_45_groupi_n_443, csa_tree_add_7_45_groupi_n_444, csa_tree_add_7_45_groupi_n_445, csa_tree_add_7_45_groupi_n_446, csa_tree_add_7_45_groupi_n_447, csa_tree_add_7_45_groupi_n_448, csa_tree_add_7_45_groupi_n_449;
  wire csa_tree_add_7_45_groupi_n_450, csa_tree_add_7_45_groupi_n_451, csa_tree_add_7_45_groupi_n_452, csa_tree_add_7_45_groupi_n_453, csa_tree_add_7_45_groupi_n_454, csa_tree_add_7_45_groupi_n_455, csa_tree_add_7_45_groupi_n_456, csa_tree_add_7_45_groupi_n_457;
  wire csa_tree_add_7_45_groupi_n_458, csa_tree_add_7_45_groupi_n_460, csa_tree_add_7_45_groupi_n_461, csa_tree_add_7_45_groupi_n_462, csa_tree_add_7_45_groupi_n_463, csa_tree_add_7_45_groupi_n_464, csa_tree_add_7_45_groupi_n_465, csa_tree_add_7_45_groupi_n_466;
  wire csa_tree_add_7_45_groupi_n_467, csa_tree_add_7_45_groupi_n_468, csa_tree_add_7_45_groupi_n_469, csa_tree_add_7_45_groupi_n_470, csa_tree_add_7_45_groupi_n_471, csa_tree_add_7_45_groupi_n_472, csa_tree_add_7_45_groupi_n_473, csa_tree_add_7_45_groupi_n_474;
  wire csa_tree_add_7_45_groupi_n_475, csa_tree_add_7_45_groupi_n_476, csa_tree_add_7_45_groupi_n_477, csa_tree_add_7_45_groupi_n_478, csa_tree_add_7_45_groupi_n_479, csa_tree_add_7_45_groupi_n_480, csa_tree_add_7_45_groupi_n_481, csa_tree_add_7_45_groupi_n_482;
  wire csa_tree_add_7_45_groupi_n_483, csa_tree_add_7_45_groupi_n_484, csa_tree_add_7_45_groupi_n_485, csa_tree_add_7_45_groupi_n_486, csa_tree_add_7_45_groupi_n_487, csa_tree_add_7_45_groupi_n_488, csa_tree_add_7_45_groupi_n_489, csa_tree_add_7_45_groupi_n_490;
  wire csa_tree_add_7_45_groupi_n_491, csa_tree_add_7_45_groupi_n_492, csa_tree_add_7_45_groupi_n_493, csa_tree_add_7_45_groupi_n_494, csa_tree_add_7_45_groupi_n_495, csa_tree_add_7_45_groupi_n_496, csa_tree_add_7_45_groupi_n_497, csa_tree_add_7_45_groupi_n_498;
  wire csa_tree_add_7_45_groupi_n_499, csa_tree_add_7_45_groupi_n_500, csa_tree_add_7_45_groupi_n_501, csa_tree_add_7_45_groupi_n_502, csa_tree_add_7_45_groupi_n_503, csa_tree_add_7_45_groupi_n_504, csa_tree_add_7_45_groupi_n_505, csa_tree_add_7_45_groupi_n_506;
  wire csa_tree_add_7_45_groupi_n_507, csa_tree_add_7_45_groupi_n_508, csa_tree_add_7_45_groupi_n_509, csa_tree_add_7_45_groupi_n_510, csa_tree_add_7_45_groupi_n_511, csa_tree_add_7_45_groupi_n_512, csa_tree_add_7_45_groupi_n_513, csa_tree_add_7_45_groupi_n_514;
  wire csa_tree_add_7_45_groupi_n_515, csa_tree_add_7_45_groupi_n_516, csa_tree_add_7_45_groupi_n_517, csa_tree_add_7_45_groupi_n_518, csa_tree_add_7_45_groupi_n_519, csa_tree_add_7_45_groupi_n_520, csa_tree_add_7_45_groupi_n_521, csa_tree_add_7_45_groupi_n_522;
  wire csa_tree_add_7_45_groupi_n_523, csa_tree_add_7_45_groupi_n_524, csa_tree_add_7_45_groupi_n_525, csa_tree_add_7_45_groupi_n_526, csa_tree_add_7_45_groupi_n_527, csa_tree_add_7_45_groupi_n_528, csa_tree_add_7_45_groupi_n_529, csa_tree_add_7_45_groupi_n_530;
  wire csa_tree_add_7_45_groupi_n_531, csa_tree_add_7_45_groupi_n_532, csa_tree_add_7_45_groupi_n_533, csa_tree_add_7_45_groupi_n_534, csa_tree_add_7_45_groupi_n_535, csa_tree_add_7_45_groupi_n_536, csa_tree_add_7_45_groupi_n_537, csa_tree_add_7_45_groupi_n_538;
  wire csa_tree_add_7_45_groupi_n_539, csa_tree_add_7_45_groupi_n_540, csa_tree_add_7_45_groupi_n_541, csa_tree_add_7_45_groupi_n_542, csa_tree_add_7_45_groupi_n_543, csa_tree_add_7_45_groupi_n_544, csa_tree_add_7_45_groupi_n_545, csa_tree_add_7_45_groupi_n_546;
  wire csa_tree_add_7_45_groupi_n_547, csa_tree_add_7_45_groupi_n_548, csa_tree_add_7_45_groupi_n_549, csa_tree_add_7_45_groupi_n_550, csa_tree_add_7_45_groupi_n_551, csa_tree_add_7_45_groupi_n_552, csa_tree_add_7_45_groupi_n_553, csa_tree_add_7_45_groupi_n_554;
  wire csa_tree_add_7_45_groupi_n_555, csa_tree_add_7_45_groupi_n_556, csa_tree_add_7_45_groupi_n_557, csa_tree_add_7_45_groupi_n_558, csa_tree_add_7_45_groupi_n_559, csa_tree_add_7_45_groupi_n_560, csa_tree_add_7_45_groupi_n_561, csa_tree_add_7_45_groupi_n_562;
  wire csa_tree_add_7_45_groupi_n_563, csa_tree_add_7_45_groupi_n_564, csa_tree_add_7_45_groupi_n_565, csa_tree_add_7_45_groupi_n_566, csa_tree_add_7_45_groupi_n_567, csa_tree_add_7_45_groupi_n_568, csa_tree_add_7_45_groupi_n_569, csa_tree_add_7_45_groupi_n_570;
  wire csa_tree_add_7_45_groupi_n_571, csa_tree_add_7_45_groupi_n_572, csa_tree_add_7_45_groupi_n_573, csa_tree_add_7_45_groupi_n_574, csa_tree_add_7_45_groupi_n_575, csa_tree_add_7_45_groupi_n_576, csa_tree_add_7_45_groupi_n_577, csa_tree_add_7_45_groupi_n_578;
  wire csa_tree_add_7_45_groupi_n_579, csa_tree_add_7_45_groupi_n_580, csa_tree_add_7_45_groupi_n_581, csa_tree_add_7_45_groupi_n_582, csa_tree_add_7_45_groupi_n_583, csa_tree_add_7_45_groupi_n_584, csa_tree_add_7_45_groupi_n_585, csa_tree_add_7_45_groupi_n_586;
  wire csa_tree_add_7_45_groupi_n_587, csa_tree_add_7_45_groupi_n_588, csa_tree_add_7_45_groupi_n_589, csa_tree_add_7_45_groupi_n_590, csa_tree_add_7_45_groupi_n_591, csa_tree_add_7_45_groupi_n_592, csa_tree_add_7_45_groupi_n_593, csa_tree_add_7_45_groupi_n_594;
  wire csa_tree_add_7_45_groupi_n_595, csa_tree_add_7_45_groupi_n_596, csa_tree_add_7_45_groupi_n_597, csa_tree_add_7_45_groupi_n_598, csa_tree_add_7_45_groupi_n_599, csa_tree_add_7_45_groupi_n_600, csa_tree_add_7_45_groupi_n_601, csa_tree_add_7_45_groupi_n_602;
  wire csa_tree_add_7_45_groupi_n_603, csa_tree_add_7_45_groupi_n_604, csa_tree_add_7_45_groupi_n_605, csa_tree_add_7_45_groupi_n_606, csa_tree_add_7_45_groupi_n_607, csa_tree_add_7_45_groupi_n_608, csa_tree_add_7_45_groupi_n_609, csa_tree_add_7_45_groupi_n_610;
  wire csa_tree_add_7_45_groupi_n_611, csa_tree_add_7_45_groupi_n_612, csa_tree_add_7_45_groupi_n_613, csa_tree_add_7_45_groupi_n_614, csa_tree_add_7_45_groupi_n_615, csa_tree_add_7_45_groupi_n_616, csa_tree_add_7_45_groupi_n_617, csa_tree_add_7_45_groupi_n_618;
  wire csa_tree_add_7_45_groupi_n_619, csa_tree_add_7_45_groupi_n_620, csa_tree_add_7_45_groupi_n_621, csa_tree_add_7_45_groupi_n_622, csa_tree_add_7_45_groupi_n_623, csa_tree_add_7_45_groupi_n_624, csa_tree_add_7_45_groupi_n_625, csa_tree_add_7_45_groupi_n_626;
  wire csa_tree_add_7_45_groupi_n_627, csa_tree_add_7_45_groupi_n_628, csa_tree_add_7_45_groupi_n_629, csa_tree_add_7_45_groupi_n_630, csa_tree_add_7_45_groupi_n_631, csa_tree_add_7_45_groupi_n_632, csa_tree_add_7_45_groupi_n_633, csa_tree_add_7_45_groupi_n_634;
  wire csa_tree_add_7_45_groupi_n_635, csa_tree_add_7_45_groupi_n_636, csa_tree_add_7_45_groupi_n_637, csa_tree_add_7_45_groupi_n_638, csa_tree_add_7_45_groupi_n_639, csa_tree_add_7_45_groupi_n_640, csa_tree_add_7_45_groupi_n_641, csa_tree_add_7_45_groupi_n_642;
  wire csa_tree_add_7_45_groupi_n_643, csa_tree_add_7_45_groupi_n_644, csa_tree_add_7_45_groupi_n_645, csa_tree_add_7_45_groupi_n_646, csa_tree_add_7_45_groupi_n_647, csa_tree_add_7_45_groupi_n_648, csa_tree_add_7_45_groupi_n_649, csa_tree_add_7_45_groupi_n_650;
  wire csa_tree_add_7_45_groupi_n_651, csa_tree_add_7_45_groupi_n_652, csa_tree_add_7_45_groupi_n_653, csa_tree_add_7_45_groupi_n_654, csa_tree_add_7_45_groupi_n_655, csa_tree_add_7_45_groupi_n_656, csa_tree_add_7_45_groupi_n_657, csa_tree_add_7_45_groupi_n_658;
  wire csa_tree_add_7_45_groupi_n_659, csa_tree_add_7_45_groupi_n_660, csa_tree_add_7_45_groupi_n_661, csa_tree_add_7_45_groupi_n_662, csa_tree_add_7_45_groupi_n_663, csa_tree_add_7_45_groupi_n_664, csa_tree_add_7_45_groupi_n_665, csa_tree_add_7_45_groupi_n_666;
  wire csa_tree_add_7_45_groupi_n_667, csa_tree_add_7_45_groupi_n_668, csa_tree_add_7_45_groupi_n_669, csa_tree_add_7_45_groupi_n_670, csa_tree_add_7_45_groupi_n_671, csa_tree_add_7_45_groupi_n_672, csa_tree_add_7_45_groupi_n_673, csa_tree_add_7_45_groupi_n_674;
  wire csa_tree_add_7_45_groupi_n_675, csa_tree_add_7_45_groupi_n_676, csa_tree_add_7_45_groupi_n_677, csa_tree_add_7_45_groupi_n_678, csa_tree_add_7_45_groupi_n_679, csa_tree_add_7_45_groupi_n_680, csa_tree_add_7_45_groupi_n_681, csa_tree_add_7_45_groupi_n_682;
  wire csa_tree_add_7_45_groupi_n_683, csa_tree_add_7_45_groupi_n_684, csa_tree_add_7_45_groupi_n_685, csa_tree_add_7_45_groupi_n_686, csa_tree_add_7_45_groupi_n_687, csa_tree_add_7_45_groupi_n_688, csa_tree_add_7_45_groupi_n_689, csa_tree_add_7_45_groupi_n_690;
  wire csa_tree_add_7_45_groupi_n_691, csa_tree_add_7_45_groupi_n_692, csa_tree_add_7_45_groupi_n_693, csa_tree_add_7_45_groupi_n_694, csa_tree_add_7_45_groupi_n_695, csa_tree_add_7_45_groupi_n_696, csa_tree_add_7_45_groupi_n_697, csa_tree_add_7_45_groupi_n_698;
  wire csa_tree_add_7_45_groupi_n_699, csa_tree_add_7_45_groupi_n_700, csa_tree_add_7_45_groupi_n_701, csa_tree_add_7_45_groupi_n_702, csa_tree_add_7_45_groupi_n_703, csa_tree_add_7_45_groupi_n_704, csa_tree_add_7_45_groupi_n_705, csa_tree_add_7_45_groupi_n_706;
  wire csa_tree_add_7_45_groupi_n_707, csa_tree_add_7_45_groupi_n_708, csa_tree_add_7_45_groupi_n_709, csa_tree_add_7_45_groupi_n_710, csa_tree_add_7_45_groupi_n_711, csa_tree_add_7_45_groupi_n_712, csa_tree_add_7_45_groupi_n_713, csa_tree_add_7_45_groupi_n_714;
  wire csa_tree_add_7_45_groupi_n_715, csa_tree_add_7_45_groupi_n_716, csa_tree_add_7_45_groupi_n_717, csa_tree_add_7_45_groupi_n_718, csa_tree_add_7_45_groupi_n_719, csa_tree_add_7_45_groupi_n_720, csa_tree_add_7_45_groupi_n_721, csa_tree_add_7_45_groupi_n_722;
  wire csa_tree_add_7_45_groupi_n_723, csa_tree_add_7_45_groupi_n_724, csa_tree_add_7_45_groupi_n_725, csa_tree_add_7_45_groupi_n_726, csa_tree_add_7_45_groupi_n_727, csa_tree_add_7_45_groupi_n_728, csa_tree_add_7_45_groupi_n_729, csa_tree_add_7_45_groupi_n_730;
  wire csa_tree_add_7_45_groupi_n_731, csa_tree_add_7_45_groupi_n_732, csa_tree_add_7_45_groupi_n_733, csa_tree_add_7_45_groupi_n_734, csa_tree_add_7_45_groupi_n_735, csa_tree_add_7_45_groupi_n_736, csa_tree_add_7_45_groupi_n_737, csa_tree_add_7_45_groupi_n_738;
  wire csa_tree_add_7_45_groupi_n_739, csa_tree_add_7_45_groupi_n_740, csa_tree_add_7_45_groupi_n_741, csa_tree_add_7_45_groupi_n_742, csa_tree_add_7_45_groupi_n_743, csa_tree_add_7_45_groupi_n_744, csa_tree_add_7_45_groupi_n_745, csa_tree_add_7_45_groupi_n_746;
  wire csa_tree_add_7_45_groupi_n_747, csa_tree_add_7_45_groupi_n_748, csa_tree_add_7_45_groupi_n_749, csa_tree_add_7_45_groupi_n_750, csa_tree_add_7_45_groupi_n_751, csa_tree_add_7_45_groupi_n_752, csa_tree_add_7_45_groupi_n_753, csa_tree_add_7_45_groupi_n_754;
  wire csa_tree_add_7_45_groupi_n_755, csa_tree_add_7_45_groupi_n_756, csa_tree_add_7_45_groupi_n_757, csa_tree_add_7_45_groupi_n_758, csa_tree_add_7_45_groupi_n_759, csa_tree_add_7_45_groupi_n_760, csa_tree_add_7_45_groupi_n_761, csa_tree_add_7_45_groupi_n_762;
  wire csa_tree_add_7_45_groupi_n_763, csa_tree_add_7_45_groupi_n_764, csa_tree_add_7_45_groupi_n_765, csa_tree_add_7_45_groupi_n_766, csa_tree_add_7_45_groupi_n_767, csa_tree_add_7_45_groupi_n_768, csa_tree_add_7_45_groupi_n_769, csa_tree_add_7_45_groupi_n_770;
  wire csa_tree_add_7_45_groupi_n_771, csa_tree_add_7_45_groupi_n_772, csa_tree_add_7_45_groupi_n_773, csa_tree_add_7_45_groupi_n_774, csa_tree_add_7_45_groupi_n_775, csa_tree_add_7_45_groupi_n_776, csa_tree_add_7_45_groupi_n_777, csa_tree_add_7_45_groupi_n_778;
  wire csa_tree_add_7_45_groupi_n_779, csa_tree_add_7_45_groupi_n_780, csa_tree_add_7_45_groupi_n_781, csa_tree_add_7_45_groupi_n_782, csa_tree_add_7_45_groupi_n_783, csa_tree_add_7_45_groupi_n_784, csa_tree_add_7_45_groupi_n_785, csa_tree_add_7_45_groupi_n_786;
  wire csa_tree_add_7_45_groupi_n_787, csa_tree_add_7_45_groupi_n_788, csa_tree_add_7_45_groupi_n_789, csa_tree_add_7_45_groupi_n_790, csa_tree_add_7_45_groupi_n_791, csa_tree_add_7_45_groupi_n_792, csa_tree_add_7_45_groupi_n_793, csa_tree_add_7_45_groupi_n_794;
  wire csa_tree_add_7_45_groupi_n_795, csa_tree_add_7_45_groupi_n_796, csa_tree_add_7_45_groupi_n_797, csa_tree_add_7_45_groupi_n_798, csa_tree_add_7_45_groupi_n_799, csa_tree_add_7_45_groupi_n_800, csa_tree_add_7_45_groupi_n_801, csa_tree_add_7_45_groupi_n_802;
  wire csa_tree_add_7_45_groupi_n_803, csa_tree_add_7_45_groupi_n_804, csa_tree_add_7_45_groupi_n_805, csa_tree_add_7_45_groupi_n_806, csa_tree_add_7_45_groupi_n_807, csa_tree_add_7_45_groupi_n_808, csa_tree_add_7_45_groupi_n_809, csa_tree_add_7_45_groupi_n_810;
  wire csa_tree_add_7_45_groupi_n_812, csa_tree_add_7_45_groupi_n_813, csa_tree_add_7_45_groupi_n_814, csa_tree_add_7_45_groupi_n_815, csa_tree_add_7_45_groupi_n_816, csa_tree_add_7_45_groupi_n_817, csa_tree_add_7_45_groupi_n_818, csa_tree_add_7_45_groupi_n_819;
  wire csa_tree_add_7_45_groupi_n_820, csa_tree_add_7_45_groupi_n_821, csa_tree_add_7_45_groupi_n_822, csa_tree_add_7_45_groupi_n_823, csa_tree_add_7_45_groupi_n_824, csa_tree_add_7_45_groupi_n_825, csa_tree_add_7_45_groupi_n_826, csa_tree_add_7_45_groupi_n_827;
  wire csa_tree_add_7_45_groupi_n_828, csa_tree_add_7_45_groupi_n_829, csa_tree_add_7_45_groupi_n_830, csa_tree_add_7_45_groupi_n_831, csa_tree_add_7_45_groupi_n_832, csa_tree_add_7_45_groupi_n_833, csa_tree_add_7_45_groupi_n_834, csa_tree_add_7_45_groupi_n_835;
  wire csa_tree_add_7_45_groupi_n_836, csa_tree_add_7_45_groupi_n_837, csa_tree_add_7_45_groupi_n_838, csa_tree_add_7_45_groupi_n_839, csa_tree_add_7_45_groupi_n_840, csa_tree_add_7_45_groupi_n_841, csa_tree_add_7_45_groupi_n_842, csa_tree_add_7_45_groupi_n_843;
  wire csa_tree_add_7_45_groupi_n_844, csa_tree_add_7_45_groupi_n_845, csa_tree_add_7_45_groupi_n_846, csa_tree_add_7_45_groupi_n_847, csa_tree_add_7_45_groupi_n_848, csa_tree_add_7_45_groupi_n_849, csa_tree_add_7_45_groupi_n_850, csa_tree_add_7_45_groupi_n_851;
  wire csa_tree_add_7_45_groupi_n_852, csa_tree_add_7_45_groupi_n_853, csa_tree_add_7_45_groupi_n_854, csa_tree_add_7_45_groupi_n_855, csa_tree_add_7_45_groupi_n_856, csa_tree_add_7_45_groupi_n_857, csa_tree_add_7_45_groupi_n_858, csa_tree_add_7_45_groupi_n_859;
  wire csa_tree_add_7_45_groupi_n_860, csa_tree_add_7_45_groupi_n_861, csa_tree_add_7_45_groupi_n_862, csa_tree_add_7_45_groupi_n_863, csa_tree_add_7_45_groupi_n_864, csa_tree_add_7_45_groupi_n_865, csa_tree_add_7_45_groupi_n_866, csa_tree_add_7_45_groupi_n_867;
  wire csa_tree_add_7_45_groupi_n_868, csa_tree_add_7_45_groupi_n_869, csa_tree_add_7_45_groupi_n_870, csa_tree_add_7_45_groupi_n_871, csa_tree_add_7_45_groupi_n_872, csa_tree_add_7_45_groupi_n_873, csa_tree_add_7_45_groupi_n_874, csa_tree_add_7_45_groupi_n_875;
  wire csa_tree_add_7_45_groupi_n_876, csa_tree_add_7_45_groupi_n_877, csa_tree_add_7_45_groupi_n_878, csa_tree_add_7_45_groupi_n_879, csa_tree_add_7_45_groupi_n_880, csa_tree_add_7_45_groupi_n_881, csa_tree_add_7_45_groupi_n_882, csa_tree_add_7_45_groupi_n_883;
  wire csa_tree_add_7_45_groupi_n_884, csa_tree_add_7_45_groupi_n_885, csa_tree_add_7_45_groupi_n_886, csa_tree_add_7_45_groupi_n_887, csa_tree_add_7_45_groupi_n_888, csa_tree_add_7_45_groupi_n_889, csa_tree_add_7_45_groupi_n_890, csa_tree_add_7_45_groupi_n_891;
  wire csa_tree_add_7_45_groupi_n_892, csa_tree_add_7_45_groupi_n_893, csa_tree_add_7_45_groupi_n_894, csa_tree_add_7_45_groupi_n_895, csa_tree_add_7_45_groupi_n_896, csa_tree_add_7_45_groupi_n_897, csa_tree_add_7_45_groupi_n_898, csa_tree_add_7_45_groupi_n_899;
  wire csa_tree_add_7_45_groupi_n_900, csa_tree_add_7_45_groupi_n_901, csa_tree_add_7_45_groupi_n_902, csa_tree_add_7_45_groupi_n_903, csa_tree_add_7_45_groupi_n_904, csa_tree_add_7_45_groupi_n_905, csa_tree_add_7_45_groupi_n_906, csa_tree_add_7_45_groupi_n_907;
  wire csa_tree_add_7_45_groupi_n_908, csa_tree_add_7_45_groupi_n_909, csa_tree_add_7_45_groupi_n_910, csa_tree_add_7_45_groupi_n_911, csa_tree_add_7_45_groupi_n_912, csa_tree_add_7_45_groupi_n_913, csa_tree_add_7_45_groupi_n_914, csa_tree_add_7_45_groupi_n_915;
  wire csa_tree_add_7_45_groupi_n_916, csa_tree_add_7_45_groupi_n_917, csa_tree_add_7_45_groupi_n_918, csa_tree_add_7_45_groupi_n_919, csa_tree_add_7_45_groupi_n_920, csa_tree_add_7_45_groupi_n_921, csa_tree_add_7_45_groupi_n_922, csa_tree_add_7_45_groupi_n_923;
  wire csa_tree_add_7_45_groupi_n_924, csa_tree_add_7_45_groupi_n_925, csa_tree_add_7_45_groupi_n_926, csa_tree_add_7_45_groupi_n_927, csa_tree_add_7_45_groupi_n_928, csa_tree_add_7_45_groupi_n_929, csa_tree_add_7_45_groupi_n_930, csa_tree_add_7_45_groupi_n_931;
  wire csa_tree_add_7_45_groupi_n_932, csa_tree_add_7_45_groupi_n_933, csa_tree_add_7_45_groupi_n_934, csa_tree_add_7_45_groupi_n_935, csa_tree_add_7_45_groupi_n_936, csa_tree_add_7_45_groupi_n_937, csa_tree_add_7_45_groupi_n_938, csa_tree_add_7_45_groupi_n_939;
  wire csa_tree_add_7_45_groupi_n_940, csa_tree_add_7_45_groupi_n_941, csa_tree_add_7_45_groupi_n_942, csa_tree_add_7_45_groupi_n_943, csa_tree_add_7_45_groupi_n_944, csa_tree_add_7_45_groupi_n_945, csa_tree_add_7_45_groupi_n_946, csa_tree_add_7_45_groupi_n_947;
  wire csa_tree_add_7_45_groupi_n_948, csa_tree_add_7_45_groupi_n_949, csa_tree_add_7_45_groupi_n_950, csa_tree_add_7_45_groupi_n_951, csa_tree_add_7_45_groupi_n_952, csa_tree_add_7_45_groupi_n_953, csa_tree_add_7_45_groupi_n_954, csa_tree_add_7_45_groupi_n_955;
  wire csa_tree_add_7_45_groupi_n_956, csa_tree_add_7_45_groupi_n_957, csa_tree_add_7_45_groupi_n_958, csa_tree_add_7_45_groupi_n_959, csa_tree_add_7_45_groupi_n_960, csa_tree_add_7_45_groupi_n_961, csa_tree_add_7_45_groupi_n_962, csa_tree_add_7_45_groupi_n_963;
  wire csa_tree_add_7_45_groupi_n_964, csa_tree_add_7_45_groupi_n_966, csa_tree_add_7_45_groupi_n_967, csa_tree_add_7_45_groupi_n_968, csa_tree_add_7_45_groupi_n_969, csa_tree_add_7_45_groupi_n_970, csa_tree_add_7_45_groupi_n_971, csa_tree_add_7_45_groupi_n_972;
  wire csa_tree_add_7_45_groupi_n_973, csa_tree_add_7_45_groupi_n_974, csa_tree_add_7_45_groupi_n_975, csa_tree_add_7_45_groupi_n_976, csa_tree_add_7_45_groupi_n_977, csa_tree_add_7_45_groupi_n_978, csa_tree_add_7_45_groupi_n_979, csa_tree_add_7_45_groupi_n_980;
  wire csa_tree_add_7_45_groupi_n_981, csa_tree_add_7_45_groupi_n_982, csa_tree_add_7_45_groupi_n_983, csa_tree_add_7_45_groupi_n_984, csa_tree_add_7_45_groupi_n_985, csa_tree_add_7_45_groupi_n_986, csa_tree_add_7_45_groupi_n_987, csa_tree_add_7_45_groupi_n_988;
  wire csa_tree_add_7_45_groupi_n_989, csa_tree_add_7_45_groupi_n_990, csa_tree_add_7_45_groupi_n_991, csa_tree_add_7_45_groupi_n_992, csa_tree_add_7_45_groupi_n_993, csa_tree_add_7_45_groupi_n_994, csa_tree_add_7_45_groupi_n_995, csa_tree_add_7_45_groupi_n_996;
  wire csa_tree_add_7_45_groupi_n_997, csa_tree_add_7_45_groupi_n_998, csa_tree_add_7_45_groupi_n_999, csa_tree_add_7_45_groupi_n_1000, csa_tree_add_7_45_groupi_n_1001, csa_tree_add_7_45_groupi_n_1002, csa_tree_add_7_45_groupi_n_1003, csa_tree_add_7_45_groupi_n_1004;
  wire csa_tree_add_7_45_groupi_n_1005, csa_tree_add_7_45_groupi_n_1006, csa_tree_add_7_45_groupi_n_1007, csa_tree_add_7_45_groupi_n_1008, csa_tree_add_7_45_groupi_n_1009, csa_tree_add_7_45_groupi_n_1010, csa_tree_add_7_45_groupi_n_1011, csa_tree_add_7_45_groupi_n_1012;
  wire csa_tree_add_7_45_groupi_n_1013, csa_tree_add_7_45_groupi_n_1014, csa_tree_add_7_45_groupi_n_1015, csa_tree_add_7_45_groupi_n_1016, csa_tree_add_7_45_groupi_n_1017, csa_tree_add_7_45_groupi_n_1018, csa_tree_add_7_45_groupi_n_1019, csa_tree_add_7_45_groupi_n_1020;
  wire csa_tree_add_7_45_groupi_n_1021, csa_tree_add_7_45_groupi_n_1022, csa_tree_add_7_45_groupi_n_1023, csa_tree_add_7_45_groupi_n_1024, csa_tree_add_7_45_groupi_n_1025, csa_tree_add_7_45_groupi_n_1026, csa_tree_add_7_45_groupi_n_1027, csa_tree_add_7_45_groupi_n_1028;
  wire csa_tree_add_7_45_groupi_n_1029, csa_tree_add_7_45_groupi_n_1030, csa_tree_add_7_45_groupi_n_1031, csa_tree_add_7_45_groupi_n_1032, csa_tree_add_7_45_groupi_n_1033, csa_tree_add_7_45_groupi_n_1034, csa_tree_add_7_45_groupi_n_1035, csa_tree_add_7_45_groupi_n_1036;
  wire csa_tree_add_7_45_groupi_n_1037, csa_tree_add_7_45_groupi_n_1038, csa_tree_add_7_45_groupi_n_1039, csa_tree_add_7_45_groupi_n_1040, csa_tree_add_7_45_groupi_n_1041, csa_tree_add_7_45_groupi_n_1042, csa_tree_add_7_45_groupi_n_1043, csa_tree_add_7_45_groupi_n_1044;
  wire csa_tree_add_7_45_groupi_n_1045, csa_tree_add_7_45_groupi_n_1046, csa_tree_add_7_45_groupi_n_1047, csa_tree_add_7_45_groupi_n_1048, csa_tree_add_7_45_groupi_n_1049, csa_tree_add_7_45_groupi_n_1051, csa_tree_add_7_45_groupi_n_1052, csa_tree_add_7_45_groupi_n_1053;
  wire csa_tree_add_7_45_groupi_n_1054, csa_tree_add_7_45_groupi_n_1055, csa_tree_add_7_45_groupi_n_1056, csa_tree_add_7_45_groupi_n_1057, csa_tree_add_7_45_groupi_n_1058, csa_tree_add_7_45_groupi_n_1059, csa_tree_add_7_45_groupi_n_1060, csa_tree_add_7_45_groupi_n_1061;
  wire csa_tree_add_7_45_groupi_n_1062, csa_tree_add_7_45_groupi_n_1063, csa_tree_add_7_45_groupi_n_1064, csa_tree_add_7_45_groupi_n_1065, csa_tree_add_7_45_groupi_n_1066, csa_tree_add_7_45_groupi_n_1067, csa_tree_add_7_45_groupi_n_1068, csa_tree_add_7_45_groupi_n_1069;
  wire csa_tree_add_7_45_groupi_n_1070, csa_tree_add_7_45_groupi_n_1071, csa_tree_add_7_45_groupi_n_1072, csa_tree_add_7_45_groupi_n_1073, csa_tree_add_7_45_groupi_n_1074, csa_tree_add_7_45_groupi_n_1075, csa_tree_add_7_45_groupi_n_1076, csa_tree_add_7_45_groupi_n_1077;
  wire csa_tree_add_7_45_groupi_n_1078, csa_tree_add_7_45_groupi_n_1079, csa_tree_add_7_45_groupi_n_1080, csa_tree_add_7_45_groupi_n_1081, csa_tree_add_7_45_groupi_n_1082, csa_tree_add_7_45_groupi_n_1083, csa_tree_add_7_45_groupi_n_1084, csa_tree_add_7_45_groupi_n_1085;
  wire csa_tree_add_7_45_groupi_n_1086, csa_tree_add_7_45_groupi_n_1087, csa_tree_add_7_45_groupi_n_1088, csa_tree_add_7_45_groupi_n_1089, csa_tree_add_7_45_groupi_n_1090, csa_tree_add_7_45_groupi_n_1091, csa_tree_add_7_45_groupi_n_1092, csa_tree_add_7_45_groupi_n_1093;
  wire csa_tree_add_7_45_groupi_n_1094, csa_tree_add_7_45_groupi_n_1096, csa_tree_add_7_45_groupi_n_1097, csa_tree_add_7_45_groupi_n_1098, csa_tree_add_7_45_groupi_n_1099, csa_tree_add_7_45_groupi_n_1100, csa_tree_add_7_45_groupi_n_1101, csa_tree_add_7_45_groupi_n_1102;
  wire csa_tree_add_7_45_groupi_n_1103, csa_tree_add_7_45_groupi_n_1104, csa_tree_add_7_45_groupi_n_1105, csa_tree_add_7_45_groupi_n_1106, csa_tree_add_7_45_groupi_n_1107, csa_tree_add_7_45_groupi_n_1108, csa_tree_add_7_45_groupi_n_1109, csa_tree_add_7_45_groupi_n_1110;
  wire csa_tree_add_7_45_groupi_n_1111, csa_tree_add_7_45_groupi_n_1112, csa_tree_add_7_45_groupi_n_1113, csa_tree_add_7_45_groupi_n_1114, csa_tree_add_7_45_groupi_n_1115, csa_tree_add_7_45_groupi_n_1116, csa_tree_add_7_45_groupi_n_1117, csa_tree_add_7_45_groupi_n_1118;
  wire csa_tree_add_7_45_groupi_n_1119, csa_tree_add_7_45_groupi_n_1120, csa_tree_add_7_45_groupi_n_1121, csa_tree_add_7_45_groupi_n_1122, csa_tree_add_7_45_groupi_n_1123, csa_tree_add_7_45_groupi_n_1124, csa_tree_add_7_45_groupi_n_1125, csa_tree_add_7_45_groupi_n_1126;
  wire csa_tree_add_7_45_groupi_n_1127, csa_tree_add_7_45_groupi_n_1128, csa_tree_add_7_45_groupi_n_1129, csa_tree_add_7_45_groupi_n_1130, csa_tree_add_7_45_groupi_n_1131, csa_tree_add_7_45_groupi_n_1132, csa_tree_add_7_45_groupi_n_1133, csa_tree_add_7_45_groupi_n_1134;
  wire csa_tree_add_7_45_groupi_n_1135, csa_tree_add_7_45_groupi_n_1136, csa_tree_add_7_45_groupi_n_1137, csa_tree_add_7_45_groupi_n_1138, csa_tree_add_7_45_groupi_n_1139, csa_tree_add_7_45_groupi_n_1140, csa_tree_add_7_45_groupi_n_1141, csa_tree_add_7_45_groupi_n_1142;
  wire csa_tree_add_7_45_groupi_n_1143, csa_tree_add_7_45_groupi_n_1144, csa_tree_add_7_45_groupi_n_1145, csa_tree_add_7_45_groupi_n_1146, csa_tree_add_7_45_groupi_n_1147, csa_tree_add_7_45_groupi_n_1148, csa_tree_add_7_45_groupi_n_1149, csa_tree_add_7_45_groupi_n_1150;
  wire csa_tree_add_7_45_groupi_n_1151, csa_tree_add_7_45_groupi_n_1152, csa_tree_add_7_45_groupi_n_1153, csa_tree_add_7_45_groupi_n_1154, csa_tree_add_7_45_groupi_n_1155, csa_tree_add_7_45_groupi_n_1156, csa_tree_add_7_45_groupi_n_1157, csa_tree_add_7_45_groupi_n_1158;
  wire csa_tree_add_7_45_groupi_n_1159, csa_tree_add_7_45_groupi_n_1161, csa_tree_add_7_45_groupi_n_1162, csa_tree_add_7_45_groupi_n_1163, csa_tree_add_7_45_groupi_n_1164, csa_tree_add_7_45_groupi_n_1165, csa_tree_add_7_45_groupi_n_1166, csa_tree_add_7_45_groupi_n_1167;
  wire csa_tree_add_7_45_groupi_n_1168, csa_tree_add_7_45_groupi_n_1169, csa_tree_add_7_45_groupi_n_1170, csa_tree_add_7_45_groupi_n_1171, csa_tree_add_7_45_groupi_n_1172, csa_tree_add_7_45_groupi_n_1173, csa_tree_add_7_45_groupi_n_1174, csa_tree_add_7_45_groupi_n_1175;
  wire csa_tree_add_7_45_groupi_n_1176, csa_tree_add_7_45_groupi_n_1177, csa_tree_add_7_45_groupi_n_1178, csa_tree_add_7_45_groupi_n_1179, csa_tree_add_7_45_groupi_n_1180, csa_tree_add_7_45_groupi_n_1181, csa_tree_add_7_45_groupi_n_1182, csa_tree_add_7_45_groupi_n_1183;
  wire csa_tree_add_7_45_groupi_n_1184, csa_tree_add_7_45_groupi_n_1185, csa_tree_add_7_45_groupi_n_1186, csa_tree_add_7_45_groupi_n_1187, csa_tree_add_7_45_groupi_n_1188, csa_tree_add_7_45_groupi_n_1189, csa_tree_add_7_45_groupi_n_1190, csa_tree_add_7_45_groupi_n_1191;
  wire csa_tree_add_7_45_groupi_n_1192, csa_tree_add_7_45_groupi_n_1193, csa_tree_add_7_45_groupi_n_1194, csa_tree_add_7_45_groupi_n_1195, csa_tree_add_7_45_groupi_n_1196, csa_tree_add_7_45_groupi_n_1197, csa_tree_add_7_45_groupi_n_1198, csa_tree_add_7_45_groupi_n_1199;
  wire csa_tree_add_7_45_groupi_n_1200, csa_tree_add_7_45_groupi_n_1201, csa_tree_add_7_45_groupi_n_1202, csa_tree_add_7_45_groupi_n_1203, csa_tree_add_7_45_groupi_n_1204, csa_tree_add_7_45_groupi_n_1205, csa_tree_add_7_45_groupi_n_1206, csa_tree_add_7_45_groupi_n_1207;
  wire csa_tree_add_7_45_groupi_n_1208, csa_tree_add_7_45_groupi_n_1210, csa_tree_add_7_45_groupi_n_1211, csa_tree_add_7_45_groupi_n_1212, csa_tree_add_7_45_groupi_n_1213, csa_tree_add_7_45_groupi_n_1214, csa_tree_add_7_45_groupi_n_1215, csa_tree_add_7_45_groupi_n_1216;
  wire csa_tree_add_7_45_groupi_n_1217, csa_tree_add_7_45_groupi_n_1218, csa_tree_add_7_45_groupi_n_1219, csa_tree_add_7_45_groupi_n_1220, csa_tree_add_7_45_groupi_n_1221, csa_tree_add_7_45_groupi_n_1222, csa_tree_add_7_45_groupi_n_1223, csa_tree_add_7_45_groupi_n_1224;
  wire csa_tree_add_7_45_groupi_n_1225, csa_tree_add_7_45_groupi_n_1226, csa_tree_add_7_45_groupi_n_1227, csa_tree_add_7_45_groupi_n_1228, csa_tree_add_7_45_groupi_n_1229, csa_tree_add_7_45_groupi_n_1230, csa_tree_add_7_45_groupi_n_1231, csa_tree_add_7_45_groupi_n_1232;
  wire csa_tree_add_7_45_groupi_n_1233, csa_tree_add_7_45_groupi_n_1234, csa_tree_add_7_45_groupi_n_1235, csa_tree_add_7_45_groupi_n_1236, csa_tree_add_7_45_groupi_n_1237, csa_tree_add_7_45_groupi_n_1238, csa_tree_add_7_45_groupi_n_1239, csa_tree_add_7_45_groupi_n_1240;
  wire csa_tree_add_7_45_groupi_n_1241, csa_tree_add_7_45_groupi_n_1242, csa_tree_add_7_45_groupi_n_1243, csa_tree_add_7_45_groupi_n_1244, csa_tree_add_7_45_groupi_n_1245, csa_tree_add_7_45_groupi_n_1246, csa_tree_add_7_45_groupi_n_1247, csa_tree_add_7_45_groupi_n_1248;
  wire csa_tree_add_7_45_groupi_n_1249, csa_tree_add_7_45_groupi_n_1251, csa_tree_add_7_45_groupi_n_1252, csa_tree_add_7_45_groupi_n_1253, csa_tree_add_7_45_groupi_n_1254, csa_tree_add_7_45_groupi_n_1256, csa_tree_add_7_45_groupi_n_1257, csa_tree_add_7_45_groupi_n_1258;
  wire csa_tree_add_7_45_groupi_n_1259, csa_tree_add_7_45_groupi_n_1260, csa_tree_add_7_45_groupi_n_1261, csa_tree_add_7_45_groupi_n_1263, csa_tree_add_7_45_groupi_n_1264, csa_tree_add_7_45_groupi_n_1266, csa_tree_add_7_45_groupi_n_1267, csa_tree_add_7_45_groupi_n_1269;
  wire csa_tree_add_7_45_groupi_n_1270, csa_tree_add_7_45_groupi_n_1272, csa_tree_add_7_45_groupi_n_1273, csa_tree_add_7_45_groupi_n_1275, csa_tree_add_7_45_groupi_n_1276, csa_tree_add_7_45_groupi_n_1278, csa_tree_add_7_45_groupi_n_1279, csa_tree_add_7_45_groupi_n_1281;
  buf constbuf_n1(out1[27], 1'b0);
  buf constbuf_n2(out1[28], 1'b0);
  buf constbuf_n3(out1[29], 1'b0);
  buf constbuf_n4(out1[30], 1'b0);
  buf constbuf_n5(out1[31], 1'b0);
  buf constbuf_n6(out1[32], 1'b0);
  buf constbuf_n7(out1[33], 1'b0);
  xnor csa_tree_add_7_45_groupi_g4009__2398(out1[26] ,csa_tree_add_7_45_groupi_n_1281 ,csa_tree_add_7_45_groupi_n_159);
  nor csa_tree_add_7_45_groupi_g4010__5107(csa_tree_add_7_45_groupi_n_1281 ,csa_tree_add_7_45_groupi_n_744 ,csa_tree_add_7_45_groupi_n_1279);
  xnor csa_tree_add_7_45_groupi_g4011__6260(out1[25] ,csa_tree_add_7_45_groupi_n_1278 ,csa_tree_add_7_45_groupi_n_807);
  and csa_tree_add_7_45_groupi_g4012__4319(csa_tree_add_7_45_groupi_n_1279 ,csa_tree_add_7_45_groupi_n_786 ,csa_tree_add_7_45_groupi_n_1278);
  or csa_tree_add_7_45_groupi_g4013__8428(csa_tree_add_7_45_groupi_n_1278 ,csa_tree_add_7_45_groupi_n_978 ,csa_tree_add_7_45_groupi_n_1276);
  xnor csa_tree_add_7_45_groupi_g4014__5526(out1[24] ,csa_tree_add_7_45_groupi_n_1275 ,csa_tree_add_7_45_groupi_n_1005);
  and csa_tree_add_7_45_groupi_g4015__6783(csa_tree_add_7_45_groupi_n_1276 ,csa_tree_add_7_45_groupi_n_987 ,csa_tree_add_7_45_groupi_n_1275);
  or csa_tree_add_7_45_groupi_g4016__3680(csa_tree_add_7_45_groupi_n_1275 ,csa_tree_add_7_45_groupi_n_1035 ,csa_tree_add_7_45_groupi_n_1273);
  xnor csa_tree_add_7_45_groupi_g4017__1617(out1[23] ,csa_tree_add_7_45_groupi_n_1272 ,csa_tree_add_7_45_groupi_n_1048);
  and csa_tree_add_7_45_groupi_g4018__2802(csa_tree_add_7_45_groupi_n_1273 ,csa_tree_add_7_45_groupi_n_1006 ,csa_tree_add_7_45_groupi_n_1272);
  or csa_tree_add_7_45_groupi_g4019__1705(csa_tree_add_7_45_groupi_n_1272 ,csa_tree_add_7_45_groupi_n_1073 ,csa_tree_add_7_45_groupi_n_1270);
  xnor csa_tree_add_7_45_groupi_g4020__5122(out1[22] ,csa_tree_add_7_45_groupi_n_1269 ,csa_tree_add_7_45_groupi_n_1090);
  and csa_tree_add_7_45_groupi_g4021__8246(csa_tree_add_7_45_groupi_n_1270 ,csa_tree_add_7_45_groupi_n_1071 ,csa_tree_add_7_45_groupi_n_1269);
  or csa_tree_add_7_45_groupi_g4022__7098(csa_tree_add_7_45_groupi_n_1269 ,csa_tree_add_7_45_groupi_n_1113 ,csa_tree_add_7_45_groupi_n_1267);
  xnor csa_tree_add_7_45_groupi_g4023__6131(out1[21] ,csa_tree_add_7_45_groupi_n_1266 ,csa_tree_add_7_45_groupi_n_1128);
  and csa_tree_add_7_45_groupi_g4024__1881(csa_tree_add_7_45_groupi_n_1267 ,csa_tree_add_7_45_groupi_n_1114 ,csa_tree_add_7_45_groupi_n_1266);
  or csa_tree_add_7_45_groupi_g4025__5115(csa_tree_add_7_45_groupi_n_1266 ,csa_tree_add_7_45_groupi_n_1173 ,csa_tree_add_7_45_groupi_n_1264);
  xnor csa_tree_add_7_45_groupi_g4026__7482(out1[20] ,csa_tree_add_7_45_groupi_n_1263 ,csa_tree_add_7_45_groupi_n_1183);
  and csa_tree_add_7_45_groupi_g4027__4733(csa_tree_add_7_45_groupi_n_1264 ,csa_tree_add_7_45_groupi_n_1172 ,csa_tree_add_7_45_groupi_n_1263);
  or csa_tree_add_7_45_groupi_g4028__6161(csa_tree_add_7_45_groupi_n_1263 ,csa_tree_add_7_45_groupi_n_1186 ,csa_tree_add_7_45_groupi_n_1261);
  xnor csa_tree_add_7_45_groupi_g4029__9315(out1[19] ,csa_tree_add_7_45_groupi_n_1260 ,csa_tree_add_7_45_groupi_n_1207);
  nor csa_tree_add_7_45_groupi_g4030__9945(csa_tree_add_7_45_groupi_n_1261 ,csa_tree_add_7_45_groupi_n_1260 ,csa_tree_add_7_45_groupi_n_1185);
  and csa_tree_add_7_45_groupi_g4031__2883(csa_tree_add_7_45_groupi_n_1260 ,csa_tree_add_7_45_groupi_n_1216 ,csa_tree_add_7_45_groupi_n_1259);
  or csa_tree_add_7_45_groupi_g4033__2346(csa_tree_add_7_45_groupi_n_1259 ,csa_tree_add_7_45_groupi_n_1218 ,csa_tree_add_7_45_groupi_n_1258);
  and csa_tree_add_7_45_groupi_g4035__1666(csa_tree_add_7_45_groupi_n_1258 ,csa_tree_add_7_45_groupi_n_1220 ,csa_tree_add_7_45_groupi_n_1257);
  or csa_tree_add_7_45_groupi_g4037__7410(csa_tree_add_7_45_groupi_n_1257 ,csa_tree_add_7_45_groupi_n_1215 ,csa_tree_add_7_45_groupi_n_1256);
  and csa_tree_add_7_45_groupi_g4039__6417(csa_tree_add_7_45_groupi_n_1256 ,csa_tree_add_7_45_groupi_n_1232 ,csa_tree_add_7_45_groupi_n_1254);
  xnor csa_tree_add_7_45_groupi_g4040__5477(out1[16] ,csa_tree_add_7_45_groupi_n_1253 ,csa_tree_add_7_45_groupi_n_1235);
  or csa_tree_add_7_45_groupi_g4041__2398(csa_tree_add_7_45_groupi_n_1254 ,csa_tree_add_7_45_groupi_n_1253 ,csa_tree_add_7_45_groupi_n_1227);
  and csa_tree_add_7_45_groupi_g4042__5107(csa_tree_add_7_45_groupi_n_1253 ,csa_tree_add_7_45_groupi_n_1228 ,csa_tree_add_7_45_groupi_n_1252);
  or csa_tree_add_7_45_groupi_g4044__6260(csa_tree_add_7_45_groupi_n_1252 ,csa_tree_add_7_45_groupi_n_1226 ,csa_tree_add_7_45_groupi_n_1251);
  and csa_tree_add_7_45_groupi_g4046__4319(csa_tree_add_7_45_groupi_n_1251 ,csa_tree_add_7_45_groupi_n_1230 ,csa_tree_add_7_45_groupi_n_1249);
  xnor csa_tree_add_7_45_groupi_g4047__8428(out1[14] ,csa_tree_add_7_45_groupi_n_1248 ,csa_tree_add_7_45_groupi_n_1233);
  or csa_tree_add_7_45_groupi_g4048__5526(csa_tree_add_7_45_groupi_n_1249 ,csa_tree_add_7_45_groupi_n_1231 ,csa_tree_add_7_45_groupi_n_1248);
  and csa_tree_add_7_45_groupi_g4049__6783(csa_tree_add_7_45_groupi_n_1248 ,csa_tree_add_7_45_groupi_n_1247 ,csa_tree_add_7_45_groupi_n_1214);
  or csa_tree_add_7_45_groupi_g4051__3680(csa_tree_add_7_45_groupi_n_1247 ,csa_tree_add_7_45_groupi_n_1208 ,csa_tree_add_7_45_groupi_n_1246);
  and csa_tree_add_7_45_groupi_g4053__1617(csa_tree_add_7_45_groupi_n_1246 ,csa_tree_add_7_45_groupi_n_1219 ,csa_tree_add_7_45_groupi_n_1245);
  or csa_tree_add_7_45_groupi_g4055__2802(csa_tree_add_7_45_groupi_n_1245 ,csa_tree_add_7_45_groupi_n_1217 ,csa_tree_add_7_45_groupi_n_1244);
  and csa_tree_add_7_45_groupi_g4057__1705(csa_tree_add_7_45_groupi_n_1244 ,csa_tree_add_7_45_groupi_n_1196 ,csa_tree_add_7_45_groupi_n_1243);
  or csa_tree_add_7_45_groupi_g4059__5122(csa_tree_add_7_45_groupi_n_1243 ,csa_tree_add_7_45_groupi_n_1199 ,csa_tree_add_7_45_groupi_n_1242);
  and csa_tree_add_7_45_groupi_g4061__8246(csa_tree_add_7_45_groupi_n_1242 ,csa_tree_add_7_45_groupi_n_1197 ,csa_tree_add_7_45_groupi_n_1241);
  or csa_tree_add_7_45_groupi_g4063__7098(csa_tree_add_7_45_groupi_n_1241 ,csa_tree_add_7_45_groupi_n_1198 ,csa_tree_add_7_45_groupi_n_1240);
  and csa_tree_add_7_45_groupi_g4065__6131(csa_tree_add_7_45_groupi_n_1240 ,csa_tree_add_7_45_groupi_n_1171 ,csa_tree_add_7_45_groupi_n_1239);
  or csa_tree_add_7_45_groupi_g4067__1881(csa_tree_add_7_45_groupi_n_1239 ,csa_tree_add_7_45_groupi_n_1174 ,csa_tree_add_7_45_groupi_n_1238);
  and csa_tree_add_7_45_groupi_g4069__5115(csa_tree_add_7_45_groupi_n_1238 ,csa_tree_add_7_45_groupi_n_1147 ,csa_tree_add_7_45_groupi_n_1237);
  or csa_tree_add_7_45_groupi_g4071__7482(csa_tree_add_7_45_groupi_n_1237 ,csa_tree_add_7_45_groupi_n_1146 ,csa_tree_add_7_45_groupi_n_1236);
  and csa_tree_add_7_45_groupi_g4073__4733(csa_tree_add_7_45_groupi_n_1236 ,csa_tree_add_7_45_groupi_n_1098 ,csa_tree_add_7_45_groupi_n_1229);
  xnor csa_tree_add_7_45_groupi_g4074__6161(csa_tree_add_7_45_groupi_n_1235 ,csa_tree_add_7_45_groupi_n_1202 ,csa_tree_add_7_45_groupi_n_1210);
  xnor csa_tree_add_7_45_groupi_g4075__9315(csa_tree_add_7_45_groupi_n_1234 ,csa_tree_add_7_45_groupi_n_1188 ,csa_tree_add_7_45_groupi_n_1213);
  xnor csa_tree_add_7_45_groupi_g4076__9945(csa_tree_add_7_45_groupi_n_1233 ,csa_tree_add_7_45_groupi_n_1201 ,csa_tree_add_7_45_groupi_n_1212);
  or csa_tree_add_7_45_groupi_g4078__2883(csa_tree_add_7_45_groupi_n_1232 ,csa_tree_add_7_45_groupi_n_1202 ,csa_tree_add_7_45_groupi_n_1211);
  nor csa_tree_add_7_45_groupi_g4079__2346(csa_tree_add_7_45_groupi_n_1231 ,csa_tree_add_7_45_groupi_n_1200 ,csa_tree_add_7_45_groupi_n_1212);
  or csa_tree_add_7_45_groupi_g4080__1666(csa_tree_add_7_45_groupi_n_1230 ,csa_tree_add_7_45_groupi_n_1201 ,csa_tree_add_7_45_groupi_n_9);
  or csa_tree_add_7_45_groupi_g4081__7410(csa_tree_add_7_45_groupi_n_1229 ,csa_tree_add_7_45_groupi_n_1097 ,csa_tree_add_7_45_groupi_n_1221);
  or csa_tree_add_7_45_groupi_g4082__6417(csa_tree_add_7_45_groupi_n_1228 ,csa_tree_add_7_45_groupi_n_1187 ,csa_tree_add_7_45_groupi_n_8);
  and csa_tree_add_7_45_groupi_g4083__5477(csa_tree_add_7_45_groupi_n_1227 ,csa_tree_add_7_45_groupi_n_1202 ,csa_tree_add_7_45_groupi_n_1211);
  nor csa_tree_add_7_45_groupi_g4084__2398(csa_tree_add_7_45_groupi_n_1226 ,csa_tree_add_7_45_groupi_n_1188 ,csa_tree_add_7_45_groupi_n_1213);
  xnor csa_tree_add_7_45_groupi_g4085__5107(csa_tree_add_7_45_groupi_n_1225 ,csa_tree_add_7_45_groupi_n_1154 ,csa_tree_add_7_45_groupi_n_1194);
  xnor csa_tree_add_7_45_groupi_g4086__6260(csa_tree_add_7_45_groupi_n_1224 ,csa_tree_add_7_45_groupi_n_1177 ,csa_tree_add_7_45_groupi_n_1190);
  xnor csa_tree_add_7_45_groupi_g4087__4319(csa_tree_add_7_45_groupi_n_1223 ,csa_tree_add_7_45_groupi_n_1204 ,csa_tree_add_7_45_groupi_n_1192);
  xnor csa_tree_add_7_45_groupi_g4088__8428(csa_tree_add_7_45_groupi_n_1222 ,csa_tree_add_7_45_groupi_n_1163 ,csa_tree_add_7_45_groupi_n_1191);
  or csa_tree_add_7_45_groupi_g4090__5526(csa_tree_add_7_45_groupi_n_1220 ,csa_tree_add_7_45_groupi_n_1203 ,csa_tree_add_7_45_groupi_n_10);
  or csa_tree_add_7_45_groupi_g4091__6783(csa_tree_add_7_45_groupi_n_1219 ,csa_tree_add_7_45_groupi_n_1153 ,csa_tree_add_7_45_groupi_n_1193);
  nor csa_tree_add_7_45_groupi_g4092__3680(csa_tree_add_7_45_groupi_n_1218 ,csa_tree_add_7_45_groupi_n_1163 ,csa_tree_add_7_45_groupi_n_1191);
  nor csa_tree_add_7_45_groupi_g4093__1617(csa_tree_add_7_45_groupi_n_1217 ,csa_tree_add_7_45_groupi_n_1154 ,csa_tree_add_7_45_groupi_n_1194);
  or csa_tree_add_7_45_groupi_g4094__2802(csa_tree_add_7_45_groupi_n_1216 ,csa_tree_add_7_45_groupi_n_1162 ,csa_tree_add_7_45_groupi_n_7);
  nor csa_tree_add_7_45_groupi_g4095__1705(csa_tree_add_7_45_groupi_n_1215 ,csa_tree_add_7_45_groupi_n_1204 ,csa_tree_add_7_45_groupi_n_1192);
  or csa_tree_add_7_45_groupi_g4096__5122(csa_tree_add_7_45_groupi_n_1214 ,csa_tree_add_7_45_groupi_n_1176 ,csa_tree_add_7_45_groupi_n_1189);
  and csa_tree_add_7_45_groupi_g4097__8246(csa_tree_add_7_45_groupi_n_1221 ,csa_tree_add_7_45_groupi_n_1077 ,csa_tree_add_7_45_groupi_n_1195);
  not csa_tree_add_7_45_groupi_g4098(csa_tree_add_7_45_groupi_n_1213 ,csa_tree_add_7_45_groupi_n_8);
  not csa_tree_add_7_45_groupi_g4099(csa_tree_add_7_45_groupi_n_1212 ,csa_tree_add_7_45_groupi_n_9);
  not csa_tree_add_7_45_groupi_g4100(csa_tree_add_7_45_groupi_n_1211 ,csa_tree_add_7_45_groupi_n_1210);
  xnor csa_tree_add_7_45_groupi_g4101__7098(out1[6] ,csa_tree_add_7_45_groupi_n_1181 ,csa_tree_add_7_45_groupi_n_1091);
  nor csa_tree_add_7_45_groupi_g4102__6131(csa_tree_add_7_45_groupi_n_1208 ,csa_tree_add_7_45_groupi_n_1177 ,csa_tree_add_7_45_groupi_n_1190);
  xnor csa_tree_add_7_45_groupi_g4103__1881(csa_tree_add_7_45_groupi_n_1207 ,csa_tree_add_7_45_groupi_n_1178 ,csa_tree_add_7_45_groupi_n_1166);
  xnor csa_tree_add_7_45_groupi_g4104__5115(csa_tree_add_7_45_groupi_n_1206 ,csa_tree_add_7_45_groupi_n_1180 ,csa_tree_add_7_45_groupi_n_1169);
  xnor csa_tree_add_7_45_groupi_g4105__7482(csa_tree_add_7_45_groupi_n_1205 ,csa_tree_add_7_45_groupi_n_1152 ,csa_tree_add_7_45_groupi_n_1165);
  xnor csa_tree_add_7_45_groupi_g4108__4733(csa_tree_add_7_45_groupi_n_1210 ,csa_tree_add_7_45_groupi_n_1126 ,csa_tree_add_7_45_groupi_n_1157);
  not csa_tree_add_7_45_groupi_g4109(csa_tree_add_7_45_groupi_n_1204 ,csa_tree_add_7_45_groupi_n_1203);
  not csa_tree_add_7_45_groupi_g4110(csa_tree_add_7_45_groupi_n_1200 ,csa_tree_add_7_45_groupi_n_1201);
  nor csa_tree_add_7_45_groupi_g4111__6161(csa_tree_add_7_45_groupi_n_1199 ,csa_tree_add_7_45_groupi_n_1180 ,csa_tree_add_7_45_groupi_n_1169);
  nor csa_tree_add_7_45_groupi_g4112__9315(csa_tree_add_7_45_groupi_n_1198 ,csa_tree_add_7_45_groupi_n_1152 ,csa_tree_add_7_45_groupi_n_1165);
  or csa_tree_add_7_45_groupi_g4113__9945(csa_tree_add_7_45_groupi_n_1197 ,csa_tree_add_7_45_groupi_n_1151 ,csa_tree_add_7_45_groupi_n_1164);
  or csa_tree_add_7_45_groupi_g4114__2883(csa_tree_add_7_45_groupi_n_1196 ,csa_tree_add_7_45_groupi_n_1179 ,csa_tree_add_7_45_groupi_n_1168);
  or csa_tree_add_7_45_groupi_g4115__2346(csa_tree_add_7_45_groupi_n_1195 ,csa_tree_add_7_45_groupi_n_1076 ,csa_tree_add_7_45_groupi_n_1182);
  and csa_tree_add_7_45_groupi_g4116__1666(csa_tree_add_7_45_groupi_n_1203 ,csa_tree_add_7_45_groupi_n_1142 ,csa_tree_add_7_45_groupi_n_1170);
  and csa_tree_add_7_45_groupi_g4117__7410(csa_tree_add_7_45_groupi_n_1202 ,csa_tree_add_7_45_groupi_n_1145 ,csa_tree_add_7_45_groupi_n_1159);
  and csa_tree_add_7_45_groupi_g4118__6417(csa_tree_add_7_45_groupi_n_1201 ,csa_tree_add_7_45_groupi_n_1135 ,csa_tree_add_7_45_groupi_n_1175);
  not csa_tree_add_7_45_groupi_g4119(csa_tree_add_7_45_groupi_n_1194 ,csa_tree_add_7_45_groupi_n_1193);
  not csa_tree_add_7_45_groupi_g4120(csa_tree_add_7_45_groupi_n_1192 ,csa_tree_add_7_45_groupi_n_10);
  not csa_tree_add_7_45_groupi_g4121(csa_tree_add_7_45_groupi_n_1191 ,csa_tree_add_7_45_groupi_n_7);
  not csa_tree_add_7_45_groupi_g4122(csa_tree_add_7_45_groupi_n_1190 ,csa_tree_add_7_45_groupi_n_1189);
  not csa_tree_add_7_45_groupi_g4123(csa_tree_add_7_45_groupi_n_1188 ,csa_tree_add_7_45_groupi_n_1187);
  nor csa_tree_add_7_45_groupi_g4124__5477(csa_tree_add_7_45_groupi_n_1186 ,csa_tree_add_7_45_groupi_n_1178 ,csa_tree_add_7_45_groupi_n_1167);
  and csa_tree_add_7_45_groupi_g4125__2398(csa_tree_add_7_45_groupi_n_1185 ,csa_tree_add_7_45_groupi_n_1178 ,csa_tree_add_7_45_groupi_n_1167);
  xnor csa_tree_add_7_45_groupi_g4126__5107(csa_tree_add_7_45_groupi_n_1184 ,csa_tree_add_7_45_groupi_n_1122 ,csa_tree_add_7_45_groupi_n_1140);
  xnor csa_tree_add_7_45_groupi_g4127__6260(csa_tree_add_7_45_groupi_n_1183 ,csa_tree_add_7_45_groupi_n_1099 ,csa_tree_add_7_45_groupi_n_1150);
  xnor csa_tree_add_7_45_groupi_g4128__4319(csa_tree_add_7_45_groupi_n_1193 ,csa_tree_add_7_45_groupi_n_1085 ,csa_tree_add_7_45_groupi_n_1131);
  xnor csa_tree_add_7_45_groupi_g4131__8428(csa_tree_add_7_45_groupi_n_1189 ,csa_tree_add_7_45_groupi_n_1102 ,csa_tree_add_7_45_groupi_n_1132);
  and csa_tree_add_7_45_groupi_g4132__5526(csa_tree_add_7_45_groupi_n_1187 ,csa_tree_add_7_45_groupi_n_1137 ,csa_tree_add_7_45_groupi_n_1161);
  not csa_tree_add_7_45_groupi_g4133(csa_tree_add_7_45_groupi_n_1182 ,csa_tree_add_7_45_groupi_n_1181);
  not csa_tree_add_7_45_groupi_g4134(csa_tree_add_7_45_groupi_n_1180 ,csa_tree_add_7_45_groupi_n_1179);
  not csa_tree_add_7_45_groupi_g4135(csa_tree_add_7_45_groupi_n_1177 ,csa_tree_add_7_45_groupi_n_1176);
  or csa_tree_add_7_45_groupi_g4136__6783(csa_tree_add_7_45_groupi_n_1175 ,csa_tree_add_7_45_groupi_n_1088 ,csa_tree_add_7_45_groupi_n_1133);
  nor csa_tree_add_7_45_groupi_g4137__3680(csa_tree_add_7_45_groupi_n_1174 ,csa_tree_add_7_45_groupi_n_1122 ,csa_tree_add_7_45_groupi_n_1140);
  and csa_tree_add_7_45_groupi_g4138__1617(csa_tree_add_7_45_groupi_n_1173 ,csa_tree_add_7_45_groupi_n_1099 ,csa_tree_add_7_45_groupi_n_1150);
  or csa_tree_add_7_45_groupi_g4139__2802(csa_tree_add_7_45_groupi_n_1172 ,csa_tree_add_7_45_groupi_n_1099 ,csa_tree_add_7_45_groupi_n_1150);
  or csa_tree_add_7_45_groupi_g4140__1705(csa_tree_add_7_45_groupi_n_1171 ,csa_tree_add_7_45_groupi_n_1121 ,csa_tree_add_7_45_groupi_n_1139);
  or csa_tree_add_7_45_groupi_g4141__5122(csa_tree_add_7_45_groupi_n_1170 ,csa_tree_add_7_45_groupi_n_1126 ,csa_tree_add_7_45_groupi_n_1143);
  or csa_tree_add_7_45_groupi_g4142__8246(csa_tree_add_7_45_groupi_n_1181 ,csa_tree_add_7_45_groupi_n_1081 ,csa_tree_add_7_45_groupi_n_1144);
  and csa_tree_add_7_45_groupi_g4143__7098(csa_tree_add_7_45_groupi_n_1179 ,csa_tree_add_7_45_groupi_n_1118 ,csa_tree_add_7_45_groupi_n_1141);
  and csa_tree_add_7_45_groupi_g4144__6131(csa_tree_add_7_45_groupi_n_1178 ,csa_tree_add_7_45_groupi_n_1116 ,csa_tree_add_7_45_groupi_n_1148);
  and csa_tree_add_7_45_groupi_g4145__1881(csa_tree_add_7_45_groupi_n_1176 ,csa_tree_add_7_45_groupi_n_1110 ,csa_tree_add_7_45_groupi_n_1149);
  not csa_tree_add_7_45_groupi_g4146(csa_tree_add_7_45_groupi_n_1169 ,csa_tree_add_7_45_groupi_n_1168);
  not csa_tree_add_7_45_groupi_g4147(csa_tree_add_7_45_groupi_n_1167 ,csa_tree_add_7_45_groupi_n_1166);
  not csa_tree_add_7_45_groupi_g4148(csa_tree_add_7_45_groupi_n_1165 ,csa_tree_add_7_45_groupi_n_1164);
  not csa_tree_add_7_45_groupi_g4149(csa_tree_add_7_45_groupi_n_1163 ,csa_tree_add_7_45_groupi_n_1162);
  or csa_tree_add_7_45_groupi_g4150__5115(csa_tree_add_7_45_groupi_n_1161 ,csa_tree_add_7_45_groupi_n_1123 ,csa_tree_add_7_45_groupi_n_1136);
  xnor csa_tree_add_7_45_groupi_g4151__7482(out1[5] ,csa_tree_add_7_45_groupi_n_1124 ,csa_tree_add_7_45_groupi_n_1092);
  or csa_tree_add_7_45_groupi_g4152__4733(csa_tree_add_7_45_groupi_n_1159 ,csa_tree_add_7_45_groupi_n_1108 ,csa_tree_add_7_45_groupi_n_1138);
  xnor csa_tree_add_7_45_groupi_g4153__6161(csa_tree_add_7_45_groupi_n_1158 ,csa_tree_add_7_45_groupi_n_1010 ,csa_tree_add_7_45_groupi_n_1105);
  xnor csa_tree_add_7_45_groupi_g4154__9315(csa_tree_add_7_45_groupi_n_1157 ,csa_tree_add_7_45_groupi_n_1025 ,csa_tree_add_7_45_groupi_n_1101);
  xnor csa_tree_add_7_45_groupi_g4155__9945(csa_tree_add_7_45_groupi_n_1156 ,csa_tree_add_7_45_groupi_n_1017 ,csa_tree_add_7_45_groupi_n_1107);
  xnor csa_tree_add_7_45_groupi_g4156__2883(csa_tree_add_7_45_groupi_n_1155 ,csa_tree_add_7_45_groupi_n_1084 ,csa_tree_add_7_45_groupi_n_1104);
  xnor csa_tree_add_7_45_groupi_g4157__2346(csa_tree_add_7_45_groupi_n_1168 ,csa_tree_add_7_45_groupi_n_1068 ,csa_tree_add_7_45_groupi_n_1094);
  xnor csa_tree_add_7_45_groupi_g4158__1666(csa_tree_add_7_45_groupi_n_1166 ,csa_tree_add_7_45_groupi_n_1087 ,csa_tree_add_7_45_groupi_n_1089);
  xnor csa_tree_add_7_45_groupi_g4159__7410(csa_tree_add_7_45_groupi_n_1164 ,csa_tree_add_7_45_groupi_n_1057 ,csa_tree_add_7_45_groupi_n_1093);
  and csa_tree_add_7_45_groupi_g4160__6417(csa_tree_add_7_45_groupi_n_1162 ,csa_tree_add_7_45_groupi_n_1096 ,csa_tree_add_7_45_groupi_n_1134);
  not csa_tree_add_7_45_groupi_g4161(csa_tree_add_7_45_groupi_n_1154 ,csa_tree_add_7_45_groupi_n_1153);
  not csa_tree_add_7_45_groupi_g4162(csa_tree_add_7_45_groupi_n_1152 ,csa_tree_add_7_45_groupi_n_1151);
  or csa_tree_add_7_45_groupi_g4163__5477(csa_tree_add_7_45_groupi_n_1149 ,csa_tree_add_7_45_groupi_n_1086 ,csa_tree_add_7_45_groupi_n_1109);
  or csa_tree_add_7_45_groupi_g4164__2398(csa_tree_add_7_45_groupi_n_1148 ,csa_tree_add_7_45_groupi_n_1067 ,csa_tree_add_7_45_groupi_n_1115);
  or csa_tree_add_7_45_groupi_g4165__5107(csa_tree_add_7_45_groupi_n_1147 ,csa_tree_add_7_45_groupi_n_1083 ,csa_tree_add_7_45_groupi_n_1103);
  nor csa_tree_add_7_45_groupi_g4166__6260(csa_tree_add_7_45_groupi_n_1146 ,csa_tree_add_7_45_groupi_n_1084 ,csa_tree_add_7_45_groupi_n_1104);
  or csa_tree_add_7_45_groupi_g4167__4319(csa_tree_add_7_45_groupi_n_1145 ,csa_tree_add_7_45_groupi_n_1010 ,csa_tree_add_7_45_groupi_n_1106);
  nor csa_tree_add_7_45_groupi_g4168__8428(csa_tree_add_7_45_groupi_n_1144 ,csa_tree_add_7_45_groupi_n_1055 ,csa_tree_add_7_45_groupi_n_1124);
  nor csa_tree_add_7_45_groupi_g4169__5526(csa_tree_add_7_45_groupi_n_1143 ,csa_tree_add_7_45_groupi_n_1024 ,csa_tree_add_7_45_groupi_n_1101);
  or csa_tree_add_7_45_groupi_g4170__6783(csa_tree_add_7_45_groupi_n_1142 ,csa_tree_add_7_45_groupi_n_1025 ,csa_tree_add_7_45_groupi_n_1100);
  or csa_tree_add_7_45_groupi_g4171__3680(csa_tree_add_7_45_groupi_n_1141 ,csa_tree_add_7_45_groupi_n_1043 ,csa_tree_add_7_45_groupi_n_1119);
  and csa_tree_add_7_45_groupi_g4172__1617(csa_tree_add_7_45_groupi_n_1153 ,csa_tree_add_7_45_groupi_n_1054 ,csa_tree_add_7_45_groupi_n_1117);
  and csa_tree_add_7_45_groupi_g4173__2802(csa_tree_add_7_45_groupi_n_1151 ,csa_tree_add_7_45_groupi_n_1034 ,csa_tree_add_7_45_groupi_n_1120);
  or csa_tree_add_7_45_groupi_g4174__1705(csa_tree_add_7_45_groupi_n_1150 ,csa_tree_add_7_45_groupi_n_1074 ,csa_tree_add_7_45_groupi_n_1111);
  not csa_tree_add_7_45_groupi_g4175(csa_tree_add_7_45_groupi_n_1140 ,csa_tree_add_7_45_groupi_n_1139);
  and csa_tree_add_7_45_groupi_g4176__5122(csa_tree_add_7_45_groupi_n_1138 ,csa_tree_add_7_45_groupi_n_1010 ,csa_tree_add_7_45_groupi_n_1106);
  or csa_tree_add_7_45_groupi_g4177__8246(csa_tree_add_7_45_groupi_n_1137 ,csa_tree_add_7_45_groupi_n_1017 ,csa_tree_add_7_45_groupi_n_6);
  nor csa_tree_add_7_45_groupi_g4178__7098(csa_tree_add_7_45_groupi_n_1136 ,csa_tree_add_7_45_groupi_n_1016 ,csa_tree_add_7_45_groupi_n_1107);
  or csa_tree_add_7_45_groupi_g4179__6131(csa_tree_add_7_45_groupi_n_1135 ,csa_tree_add_7_45_groupi_n_1012 ,csa_tree_add_7_45_groupi_n_5);
  or csa_tree_add_7_45_groupi_g4180__1881(csa_tree_add_7_45_groupi_n_1134 ,csa_tree_add_7_45_groupi_n_1125 ,csa_tree_add_7_45_groupi_n_1112);
  nor csa_tree_add_7_45_groupi_g4181__5115(csa_tree_add_7_45_groupi_n_1133 ,csa_tree_add_7_45_groupi_n_1013 ,csa_tree_add_7_45_groupi_n_1102);
  xnor csa_tree_add_7_45_groupi_g4182__7482(csa_tree_add_7_45_groupi_n_1132 ,csa_tree_add_7_45_groupi_n_1088 ,csa_tree_add_7_45_groupi_n_1013);
  xnor csa_tree_add_7_45_groupi_g4183__4733(csa_tree_add_7_45_groupi_n_1131 ,csa_tree_add_7_45_groupi_n_1009 ,csa_tree_add_7_45_groupi_n_1059);
  xnor csa_tree_add_7_45_groupi_g4184__6161(csa_tree_add_7_45_groupi_n_1130 ,csa_tree_add_7_45_groupi_n_970 ,csa_tree_add_7_45_groupi_n_1063);
  xnor csa_tree_add_7_45_groupi_g4185__9315(csa_tree_add_7_45_groupi_n_1129 ,csa_tree_add_7_45_groupi_n_974 ,csa_tree_add_7_45_groupi_n_1061);
  xnor csa_tree_add_7_45_groupi_g4186__9945(csa_tree_add_7_45_groupi_n_1128 ,csa_tree_add_7_45_groupi_n_1082 ,csa_tree_add_7_45_groupi_n_1064);
  xnor csa_tree_add_7_45_groupi_g4187__2883(csa_tree_add_7_45_groupi_n_1127 ,csa_tree_add_7_45_groupi_n_995 ,csa_tree_add_7_45_groupi_n_1066);
  xnor csa_tree_add_7_45_groupi_g4188__2346(csa_tree_add_7_45_groupi_n_1139 ,csa_tree_add_7_45_groupi_n_1070 ,csa_tree_add_7_45_groupi_n_1049);
  not csa_tree_add_7_45_groupi_g4191(csa_tree_add_7_45_groupi_n_1122 ,csa_tree_add_7_45_groupi_n_1121);
  or csa_tree_add_7_45_groupi_g4192__1666(csa_tree_add_7_45_groupi_n_1120 ,csa_tree_add_7_45_groupi_n_1033 ,csa_tree_add_7_45_groupi_n_1070);
  nor csa_tree_add_7_45_groupi_g4193__7410(csa_tree_add_7_45_groupi_n_1119 ,csa_tree_add_7_45_groupi_n_972 ,csa_tree_add_7_45_groupi_n_1057);
  or csa_tree_add_7_45_groupi_g4194__6417(csa_tree_add_7_45_groupi_n_1118 ,csa_tree_add_7_45_groupi_n_971 ,csa_tree_add_7_45_groupi_n_1056);
  or csa_tree_add_7_45_groupi_g4195__5477(csa_tree_add_7_45_groupi_n_1117 ,csa_tree_add_7_45_groupi_n_1053 ,csa_tree_add_7_45_groupi_n_1069);
  or csa_tree_add_7_45_groupi_g4196__2398(csa_tree_add_7_45_groupi_n_1116 ,csa_tree_add_7_45_groupi_n_970 ,csa_tree_add_7_45_groupi_n_1062);
  nor csa_tree_add_7_45_groupi_g4197__5107(csa_tree_add_7_45_groupi_n_1115 ,csa_tree_add_7_45_groupi_n_969 ,csa_tree_add_7_45_groupi_n_1063);
  or csa_tree_add_7_45_groupi_g4198__6260(csa_tree_add_7_45_groupi_n_1114 ,csa_tree_add_7_45_groupi_n_1082 ,csa_tree_add_7_45_groupi_n_1064);
  and csa_tree_add_7_45_groupi_g4199__4319(csa_tree_add_7_45_groupi_n_1113 ,csa_tree_add_7_45_groupi_n_1082 ,csa_tree_add_7_45_groupi_n_1064);
  nor csa_tree_add_7_45_groupi_g4200__8428(csa_tree_add_7_45_groupi_n_1112 ,csa_tree_add_7_45_groupi_n_973 ,csa_tree_add_7_45_groupi_n_1061);
  nor csa_tree_add_7_45_groupi_g4201__5526(csa_tree_add_7_45_groupi_n_1111 ,csa_tree_add_7_45_groupi_n_1087 ,csa_tree_add_7_45_groupi_n_1078);
  or csa_tree_add_7_45_groupi_g4202__6783(csa_tree_add_7_45_groupi_n_1110 ,csa_tree_add_7_45_groupi_n_1009 ,csa_tree_add_7_45_groupi_n_1058);
  nor csa_tree_add_7_45_groupi_g4203__3680(csa_tree_add_7_45_groupi_n_1109 ,csa_tree_add_7_45_groupi_n_1008 ,csa_tree_add_7_45_groupi_n_1059);
  and csa_tree_add_7_45_groupi_g4204__1617(csa_tree_add_7_45_groupi_n_1126 ,csa_tree_add_7_45_groupi_n_940 ,csa_tree_add_7_45_groupi_n_1052);
  and csa_tree_add_7_45_groupi_g4205__2802(csa_tree_add_7_45_groupi_n_1125 ,csa_tree_add_7_45_groupi_n_939 ,csa_tree_add_7_45_groupi_n_1080);
  and csa_tree_add_7_45_groupi_g4206__1705(csa_tree_add_7_45_groupi_n_1124 ,csa_tree_add_7_45_groupi_n_983 ,csa_tree_add_7_45_groupi_n_1072);
  and csa_tree_add_7_45_groupi_g4207__5122(csa_tree_add_7_45_groupi_n_1123 ,csa_tree_add_7_45_groupi_n_921 ,csa_tree_add_7_45_groupi_n_1075);
  and csa_tree_add_7_45_groupi_g4208__8246(csa_tree_add_7_45_groupi_n_1121 ,csa_tree_add_7_45_groupi_n_985 ,csa_tree_add_7_45_groupi_n_1079);
  not csa_tree_add_7_45_groupi_g4210(csa_tree_add_7_45_groupi_n_1107 ,csa_tree_add_7_45_groupi_n_6);
  not csa_tree_add_7_45_groupi_g4211(csa_tree_add_7_45_groupi_n_1106 ,csa_tree_add_7_45_groupi_n_1105);
  not csa_tree_add_7_45_groupi_g4212(csa_tree_add_7_45_groupi_n_1104 ,csa_tree_add_7_45_groupi_n_1103);
  not csa_tree_add_7_45_groupi_g4213(csa_tree_add_7_45_groupi_n_1102 ,csa_tree_add_7_45_groupi_n_5);
  not csa_tree_add_7_45_groupi_g4214(csa_tree_add_7_45_groupi_n_1101 ,csa_tree_add_7_45_groupi_n_1100);
  or csa_tree_add_7_45_groupi_g4215__7098(csa_tree_add_7_45_groupi_n_1098 ,csa_tree_add_7_45_groupi_n_994 ,csa_tree_add_7_45_groupi_n_1065);
  nor csa_tree_add_7_45_groupi_g4216__6131(csa_tree_add_7_45_groupi_n_1097 ,csa_tree_add_7_45_groupi_n_995 ,csa_tree_add_7_45_groupi_n_1066);
  or csa_tree_add_7_45_groupi_g4217__1881(csa_tree_add_7_45_groupi_n_1096 ,csa_tree_add_7_45_groupi_n_974 ,csa_tree_add_7_45_groupi_n_1060);
  xnor csa_tree_add_7_45_groupi_g4218__5115(out1[4] ,csa_tree_add_7_45_groupi_n_1041 ,csa_tree_add_7_45_groupi_n_1002);
  xnor csa_tree_add_7_45_groupi_g4219__7482(csa_tree_add_7_45_groupi_n_1094 ,csa_tree_add_7_45_groupi_n_1021 ,csa_tree_add_7_45_groupi_n_1037);
  xnor csa_tree_add_7_45_groupi_g4220__4733(csa_tree_add_7_45_groupi_n_1093 ,csa_tree_add_7_45_groupi_n_972 ,csa_tree_add_7_45_groupi_n_1043);
  xnor csa_tree_add_7_45_groupi_g4221__6161(csa_tree_add_7_45_groupi_n_1092 ,csa_tree_add_7_45_groupi_n_950 ,csa_tree_add_7_45_groupi_n_1018);
  xnor csa_tree_add_7_45_groupi_g4222__9315(csa_tree_add_7_45_groupi_n_1091 ,csa_tree_add_7_45_groupi_n_1011 ,csa_tree_add_7_45_groupi_n_1040);
  xnor csa_tree_add_7_45_groupi_g4223__9945(csa_tree_add_7_45_groupi_n_1090 ,csa_tree_add_7_45_groupi_n_1023 ,csa_tree_add_7_45_groupi_n_1039);
  xnor csa_tree_add_7_45_groupi_g4224__2883(csa_tree_add_7_45_groupi_n_1089 ,csa_tree_add_7_45_groupi_n_825 ,csa_tree_add_7_45_groupi_n_1014);
  and csa_tree_add_7_45_groupi_g4225__2346(csa_tree_add_7_45_groupi_n_1108 ,csa_tree_add_7_45_groupi_n_931 ,csa_tree_add_7_45_groupi_n_1051);
  xnor csa_tree_add_7_45_groupi_g4227__1666(csa_tree_add_7_45_groupi_n_1105 ,csa_tree_add_7_45_groupi_n_1045 ,csa_tree_add_7_45_groupi_n_963);
  xnor csa_tree_add_7_45_groupi_g4228__7410(csa_tree_add_7_45_groupi_n_1103 ,csa_tree_add_7_45_groupi_n_1026 ,csa_tree_add_7_45_groupi_n_1004);
  xnor csa_tree_add_7_45_groupi_g4230__6417(csa_tree_add_7_45_groupi_n_1100 ,csa_tree_add_7_45_groupi_n_1046 ,csa_tree_add_7_45_groupi_n_953);
  xnor csa_tree_add_7_45_groupi_g4231__5477(csa_tree_add_7_45_groupi_n_1099 ,csa_tree_add_7_45_groupi_n_997 ,csa_tree_add_7_45_groupi_n_1003);
  not csa_tree_add_7_45_groupi_g4232(csa_tree_add_7_45_groupi_n_1086 ,csa_tree_add_7_45_groupi_n_1085);
  not csa_tree_add_7_45_groupi_g4233(csa_tree_add_7_45_groupi_n_1083 ,csa_tree_add_7_45_groupi_n_1084);
  nor csa_tree_add_7_45_groupi_g4234__2398(csa_tree_add_7_45_groupi_n_1081 ,csa_tree_add_7_45_groupi_n_950 ,csa_tree_add_7_45_groupi_n_1019);
  or csa_tree_add_7_45_groupi_g4235__5107(csa_tree_add_7_45_groupi_n_1080 ,csa_tree_add_7_45_groupi_n_945 ,csa_tree_add_7_45_groupi_n_1046);
  or csa_tree_add_7_45_groupi_g4236__6260(csa_tree_add_7_45_groupi_n_1079 ,csa_tree_add_7_45_groupi_n_984 ,csa_tree_add_7_45_groupi_n_1027);
  and csa_tree_add_7_45_groupi_g4237__4319(csa_tree_add_7_45_groupi_n_1078 ,csa_tree_add_7_45_groupi_n_825 ,csa_tree_add_7_45_groupi_n_1015);
  or csa_tree_add_7_45_groupi_g4238__8428(csa_tree_add_7_45_groupi_n_1077 ,csa_tree_add_7_45_groupi_n_1040 ,csa_tree_add_7_45_groupi_n_1011);
  and csa_tree_add_7_45_groupi_g4239__5526(csa_tree_add_7_45_groupi_n_1076 ,csa_tree_add_7_45_groupi_n_1040 ,csa_tree_add_7_45_groupi_n_1011);
  or csa_tree_add_7_45_groupi_g4240__6783(csa_tree_add_7_45_groupi_n_1075 ,csa_tree_add_7_45_groupi_n_920 ,csa_tree_add_7_45_groupi_n_1044);
  nor csa_tree_add_7_45_groupi_g4241__3680(csa_tree_add_7_45_groupi_n_1074 ,csa_tree_add_7_45_groupi_n_825 ,csa_tree_add_7_45_groupi_n_1015);
  nor csa_tree_add_7_45_groupi_g4242__1617(csa_tree_add_7_45_groupi_n_1073 ,csa_tree_add_7_45_groupi_n_1039 ,csa_tree_add_7_45_groupi_n_1023);
  or csa_tree_add_7_45_groupi_g4243__2802(csa_tree_add_7_45_groupi_n_1072 ,csa_tree_add_7_45_groupi_n_990 ,csa_tree_add_7_45_groupi_n_1042);
  or csa_tree_add_7_45_groupi_g4244__1705(csa_tree_add_7_45_groupi_n_1071 ,csa_tree_add_7_45_groupi_n_1038 ,csa_tree_add_7_45_groupi_n_1022);
  and csa_tree_add_7_45_groupi_g4245__5122(csa_tree_add_7_45_groupi_n_1088 ,csa_tree_add_7_45_groupi_n_901 ,csa_tree_add_7_45_groupi_n_1029);
  and csa_tree_add_7_45_groupi_g4246__8246(csa_tree_add_7_45_groupi_n_1087 ,csa_tree_add_7_45_groupi_n_937 ,csa_tree_add_7_45_groupi_n_1032);
  or csa_tree_add_7_45_groupi_g4247__7098(csa_tree_add_7_45_groupi_n_1085 ,csa_tree_add_7_45_groupi_n_910 ,csa_tree_add_7_45_groupi_n_1030);
  or csa_tree_add_7_45_groupi_g4248__6131(csa_tree_add_7_45_groupi_n_1084 ,csa_tree_add_7_45_groupi_n_867 ,csa_tree_add_7_45_groupi_n_1031);
  or csa_tree_add_7_45_groupi_g4249__1881(csa_tree_add_7_45_groupi_n_1082 ,csa_tree_add_7_45_groupi_n_980 ,csa_tree_add_7_45_groupi_n_1028);
  not csa_tree_add_7_45_groupi_g4250(csa_tree_add_7_45_groupi_n_1069 ,csa_tree_add_7_45_groupi_n_1068);
  not csa_tree_add_7_45_groupi_g4252(csa_tree_add_7_45_groupi_n_1066 ,csa_tree_add_7_45_groupi_n_1065);
  not csa_tree_add_7_45_groupi_g4253(csa_tree_add_7_45_groupi_n_1062 ,csa_tree_add_7_45_groupi_n_1063);
  not csa_tree_add_7_45_groupi_g4254(csa_tree_add_7_45_groupi_n_1061 ,csa_tree_add_7_45_groupi_n_1060);
  not csa_tree_add_7_45_groupi_g4255(csa_tree_add_7_45_groupi_n_1059 ,csa_tree_add_7_45_groupi_n_1058);
  not csa_tree_add_7_45_groupi_g4256(csa_tree_add_7_45_groupi_n_1057 ,csa_tree_add_7_45_groupi_n_1056);
  and csa_tree_add_7_45_groupi_g4257__5115(csa_tree_add_7_45_groupi_n_1055 ,csa_tree_add_7_45_groupi_n_950 ,csa_tree_add_7_45_groupi_n_1019);
  or csa_tree_add_7_45_groupi_g4258__7482(csa_tree_add_7_45_groupi_n_1054 ,csa_tree_add_7_45_groupi_n_1021 ,csa_tree_add_7_45_groupi_n_1036);
  nor csa_tree_add_7_45_groupi_g4259__4733(csa_tree_add_7_45_groupi_n_1053 ,csa_tree_add_7_45_groupi_n_1020 ,csa_tree_add_7_45_groupi_n_1037);
  or csa_tree_add_7_45_groupi_g4260__6161(csa_tree_add_7_45_groupi_n_1052 ,csa_tree_add_7_45_groupi_n_935 ,csa_tree_add_7_45_groupi_n_1045);
  or csa_tree_add_7_45_groupi_g4261__9315(csa_tree_add_7_45_groupi_n_1051 ,csa_tree_add_7_45_groupi_n_927 ,csa_tree_add_7_45_groupi_n_1047);
  xnor csa_tree_add_7_45_groupi_g4262__9945(out1[3] ,csa_tree_add_7_45_groupi_n_952 ,csa_tree_add_7_45_groupi_n_956);
  xnor csa_tree_add_7_45_groupi_g4263__2883(csa_tree_add_7_45_groupi_n_1049 ,csa_tree_add_7_45_groupi_n_837 ,csa_tree_add_7_45_groupi_n_993);
  xnor csa_tree_add_7_45_groupi_g4264__2346(csa_tree_add_7_45_groupi_n_1048 ,csa_tree_add_7_45_groupi_n_916 ,csa_tree_add_7_45_groupi_n_991);
  xnor csa_tree_add_7_45_groupi_g4265__1666(csa_tree_add_7_45_groupi_n_1070 ,csa_tree_add_7_45_groupi_n_799 ,csa_tree_add_7_45_groupi_n_955);
  xnor csa_tree_add_7_45_groupi_g4266__7410(csa_tree_add_7_45_groupi_n_1068 ,csa_tree_add_7_45_groupi_n_975 ,csa_tree_add_7_45_groupi_n_957);
  and csa_tree_add_7_45_groupi_g4267__6417(csa_tree_add_7_45_groupi_n_1067 ,csa_tree_add_7_45_groupi_n_923 ,csa_tree_add_7_45_groupi_n_1007);
  xnor csa_tree_add_7_45_groupi_g4268__5477(csa_tree_add_7_45_groupi_n_1065 ,csa_tree_add_7_45_groupi_n_976 ,csa_tree_add_7_45_groupi_n_891);
  xnor csa_tree_add_7_45_groupi_g4269__2398(csa_tree_add_7_45_groupi_n_1064 ,csa_tree_add_7_45_groupi_n_951 ,csa_tree_add_7_45_groupi_n_958);
  xnor csa_tree_add_7_45_groupi_g4270__5107(csa_tree_add_7_45_groupi_n_1063 ,csa_tree_add_7_45_groupi_n_1000 ,csa_tree_add_7_45_groupi_n_960);
  xnor csa_tree_add_7_45_groupi_g4271__6260(csa_tree_add_7_45_groupi_n_1060 ,csa_tree_add_7_45_groupi_n_998 ,csa_tree_add_7_45_groupi_n_961);
  xnor csa_tree_add_7_45_groupi_g4272__4319(csa_tree_add_7_45_groupi_n_1058 ,csa_tree_add_7_45_groupi_n_996 ,csa_tree_add_7_45_groupi_n_959);
  xnor csa_tree_add_7_45_groupi_g4273__8428(csa_tree_add_7_45_groupi_n_1056 ,csa_tree_add_7_45_groupi_n_876 ,csa_tree_add_7_45_groupi_n_964);
  not csa_tree_add_7_45_groupi_g4276(csa_tree_add_7_45_groupi_n_1042 ,csa_tree_add_7_45_groupi_n_1041);
  not csa_tree_add_7_45_groupi_g4277(csa_tree_add_7_45_groupi_n_1038 ,csa_tree_add_7_45_groupi_n_1039);
  not csa_tree_add_7_45_groupi_g4278(csa_tree_add_7_45_groupi_n_1037 ,csa_tree_add_7_45_groupi_n_1036);
  and csa_tree_add_7_45_groupi_g4279__5526(csa_tree_add_7_45_groupi_n_1035 ,csa_tree_add_7_45_groupi_n_916 ,csa_tree_add_7_45_groupi_n_991);
  or csa_tree_add_7_45_groupi_g4280__6783(csa_tree_add_7_45_groupi_n_1034 ,csa_tree_add_7_45_groupi_n_836 ,csa_tree_add_7_45_groupi_n_992);
  nor csa_tree_add_7_45_groupi_g4281__3680(csa_tree_add_7_45_groupi_n_1033 ,csa_tree_add_7_45_groupi_n_837 ,csa_tree_add_7_45_groupi_n_993);
  or csa_tree_add_7_45_groupi_g4282__1617(csa_tree_add_7_45_groupi_n_1032 ,csa_tree_add_7_45_groupi_n_932 ,csa_tree_add_7_45_groupi_n_1001);
  and csa_tree_add_7_45_groupi_g4283__2802(csa_tree_add_7_45_groupi_n_1031 ,csa_tree_add_7_45_groupi_n_861 ,csa_tree_add_7_45_groupi_n_976);
  nor csa_tree_add_7_45_groupi_g4284__1705(csa_tree_add_7_45_groupi_n_1030 ,csa_tree_add_7_45_groupi_n_975 ,csa_tree_add_7_45_groupi_n_909);
  or csa_tree_add_7_45_groupi_g4285__5122(csa_tree_add_7_45_groupi_n_1029 ,csa_tree_add_7_45_groupi_n_996 ,csa_tree_add_7_45_groupi_n_900);
  and csa_tree_add_7_45_groupi_g4286__8246(csa_tree_add_7_45_groupi_n_1028 ,csa_tree_add_7_45_groupi_n_997 ,csa_tree_add_7_45_groupi_n_977);
  and csa_tree_add_7_45_groupi_g4287__7098(csa_tree_add_7_45_groupi_n_1047 ,csa_tree_add_7_45_groupi_n_914 ,csa_tree_add_7_45_groupi_n_981);
  and csa_tree_add_7_45_groupi_g4288__6131(csa_tree_add_7_45_groupi_n_1046 ,csa_tree_add_7_45_groupi_n_908 ,csa_tree_add_7_45_groupi_n_968);
  and csa_tree_add_7_45_groupi_g4289__1881(csa_tree_add_7_45_groupi_n_1045 ,csa_tree_add_7_45_groupi_n_906 ,csa_tree_add_7_45_groupi_n_966);
  and csa_tree_add_7_45_groupi_g4290__5115(csa_tree_add_7_45_groupi_n_1044 ,csa_tree_add_7_45_groupi_n_904 ,csa_tree_add_7_45_groupi_n_967);
  and csa_tree_add_7_45_groupi_g4291__7482(csa_tree_add_7_45_groupi_n_1043 ,csa_tree_add_7_45_groupi_n_941 ,csa_tree_add_7_45_groupi_n_988);
  or csa_tree_add_7_45_groupi_g4292__4733(csa_tree_add_7_45_groupi_n_1041 ,csa_tree_add_7_45_groupi_n_924 ,csa_tree_add_7_45_groupi_n_982);
  and csa_tree_add_7_45_groupi_g4293__6161(csa_tree_add_7_45_groupi_n_1040 ,csa_tree_add_7_45_groupi_n_928 ,csa_tree_add_7_45_groupi_n_979);
  and csa_tree_add_7_45_groupi_g4294__9315(csa_tree_add_7_45_groupi_n_1039 ,csa_tree_add_7_45_groupi_n_915 ,csa_tree_add_7_45_groupi_n_989);
  and csa_tree_add_7_45_groupi_g4295__9945(csa_tree_add_7_45_groupi_n_1036 ,csa_tree_add_7_45_groupi_n_944 ,csa_tree_add_7_45_groupi_n_986);
  not csa_tree_add_7_45_groupi_g4296(csa_tree_add_7_45_groupi_n_1027 ,csa_tree_add_7_45_groupi_n_1026);
  not csa_tree_add_7_45_groupi_g4297(csa_tree_add_7_45_groupi_n_1025 ,csa_tree_add_7_45_groupi_n_1024);
  not csa_tree_add_7_45_groupi_g4298(csa_tree_add_7_45_groupi_n_1023 ,csa_tree_add_7_45_groupi_n_1022);
  not csa_tree_add_7_45_groupi_g4299(csa_tree_add_7_45_groupi_n_1021 ,csa_tree_add_7_45_groupi_n_1020);
  not csa_tree_add_7_45_groupi_g4300(csa_tree_add_7_45_groupi_n_1019 ,csa_tree_add_7_45_groupi_n_1018);
  not csa_tree_add_7_45_groupi_g4301(csa_tree_add_7_45_groupi_n_1017 ,csa_tree_add_7_45_groupi_n_1016);
  not csa_tree_add_7_45_groupi_g4302(csa_tree_add_7_45_groupi_n_1015 ,csa_tree_add_7_45_groupi_n_1014);
  not csa_tree_add_7_45_groupi_g4303(csa_tree_add_7_45_groupi_n_1013 ,csa_tree_add_7_45_groupi_n_1012);
  not csa_tree_add_7_45_groupi_g4304(csa_tree_add_7_45_groupi_n_1009 ,csa_tree_add_7_45_groupi_n_1008);
  or csa_tree_add_7_45_groupi_g4305__2883(csa_tree_add_7_45_groupi_n_1007 ,csa_tree_add_7_45_groupi_n_926 ,csa_tree_add_7_45_groupi_n_999);
  or csa_tree_add_7_45_groupi_g4306__2346(csa_tree_add_7_45_groupi_n_1006 ,csa_tree_add_7_45_groupi_n_916 ,csa_tree_add_7_45_groupi_n_991);
  xnor csa_tree_add_7_45_groupi_g4307__1666(csa_tree_add_7_45_groupi_n_1005 ,csa_tree_add_7_45_groupi_n_949 ,csa_tree_add_7_45_groupi_n_704);
  xnor csa_tree_add_7_45_groupi_g4308__7410(csa_tree_add_7_45_groupi_n_1004 ,csa_tree_add_7_45_groupi_n_947 ,csa_tree_add_7_45_groupi_n_833);
  xnor csa_tree_add_7_45_groupi_g4309__6417(csa_tree_add_7_45_groupi_n_1003 ,csa_tree_add_7_45_groupi_n_750 ,csa_tree_add_7_45_groupi_n_917);
  xnor csa_tree_add_7_45_groupi_g4310__5477(csa_tree_add_7_45_groupi_n_1002 ,csa_tree_add_7_45_groupi_n_789 ,csa_tree_add_7_45_groupi_n_919);
  xnor csa_tree_add_7_45_groupi_g4311__2398(csa_tree_add_7_45_groupi_n_1026 ,csa_tree_add_7_45_groupi_n_804 ,csa_tree_add_7_45_groupi_n_893);
  xnor csa_tree_add_7_45_groupi_g4312__5107(csa_tree_add_7_45_groupi_n_1024 ,csa_tree_add_7_45_groupi_n_770 ,csa_tree_add_7_45_groupi_n_896);
  xnor csa_tree_add_7_45_groupi_g4313__6260(csa_tree_add_7_45_groupi_n_1022 ,csa_tree_add_7_45_groupi_n_776 ,csa_tree_add_7_45_groupi_n_894);
  xnor csa_tree_add_7_45_groupi_g4314__4319(csa_tree_add_7_45_groupi_n_1020 ,csa_tree_add_7_45_groupi_n_753 ,csa_tree_add_7_45_groupi_n_897);
  xnor csa_tree_add_7_45_groupi_g4315__8428(csa_tree_add_7_45_groupi_n_1018 ,csa_tree_add_7_45_groupi_n_819 ,csa_tree_add_7_45_groupi_n_889);
  xnor csa_tree_add_7_45_groupi_g4316__5526(csa_tree_add_7_45_groupi_n_1016 ,csa_tree_add_7_45_groupi_n_848 ,csa_tree_add_7_45_groupi_n_888);
  xnor csa_tree_add_7_45_groupi_g4317__6783(csa_tree_add_7_45_groupi_n_1014 ,csa_tree_add_7_45_groupi_n_887 ,csa_tree_add_7_45_groupi_n_895);
  xnor csa_tree_add_7_45_groupi_g4318__3680(csa_tree_add_7_45_groupi_n_1012 ,csa_tree_add_7_45_groupi_n_827 ,csa_tree_add_7_45_groupi_n_892);
  xnor csa_tree_add_7_45_groupi_g4319__1617(csa_tree_add_7_45_groupi_n_1011 ,csa_tree_add_7_45_groupi_n_849 ,csa_tree_add_7_45_groupi_n_890);
  xnor csa_tree_add_7_45_groupi_g4320__2802(csa_tree_add_7_45_groupi_n_1010 ,csa_tree_add_7_45_groupi_n_814 ,csa_tree_add_7_45_groupi_n_899);
  xnor csa_tree_add_7_45_groupi_g4321__1705(csa_tree_add_7_45_groupi_n_1008 ,csa_tree_add_7_45_groupi_n_843 ,csa_tree_add_7_45_groupi_n_898);
  not csa_tree_add_7_45_groupi_g4322(csa_tree_add_7_45_groupi_n_1001 ,csa_tree_add_7_45_groupi_n_1000);
  not csa_tree_add_7_45_groupi_g4323(csa_tree_add_7_45_groupi_n_999 ,csa_tree_add_7_45_groupi_n_998);
  not csa_tree_add_7_45_groupi_g4324(csa_tree_add_7_45_groupi_n_995 ,csa_tree_add_7_45_groupi_n_994);
  not csa_tree_add_7_45_groupi_g4325(csa_tree_add_7_45_groupi_n_992 ,csa_tree_add_7_45_groupi_n_993);
  nor csa_tree_add_7_45_groupi_g4326__5122(csa_tree_add_7_45_groupi_n_990 ,csa_tree_add_7_45_groupi_n_789 ,csa_tree_add_7_45_groupi_n_919);
  or csa_tree_add_7_45_groupi_g4327__8246(csa_tree_add_7_45_groupi_n_989 ,csa_tree_add_7_45_groupi_n_951 ,csa_tree_add_7_45_groupi_n_942);
  or csa_tree_add_7_45_groupi_g4328__7098(csa_tree_add_7_45_groupi_n_988 ,csa_tree_add_7_45_groupi_n_799 ,csa_tree_add_7_45_groupi_n_938);
  or csa_tree_add_7_45_groupi_g4329__6131(csa_tree_add_7_45_groupi_n_987 ,csa_tree_add_7_45_groupi_n_59 ,csa_tree_add_7_45_groupi_n_948);
  or csa_tree_add_7_45_groupi_g4330__1881(csa_tree_add_7_45_groupi_n_986 ,csa_tree_add_7_45_groupi_n_800 ,csa_tree_add_7_45_groupi_n_943);
  or csa_tree_add_7_45_groupi_g4331__5115(csa_tree_add_7_45_groupi_n_985 ,csa_tree_add_7_45_groupi_n_947 ,csa_tree_add_7_45_groupi_n_832);
  nor csa_tree_add_7_45_groupi_g4332__7482(csa_tree_add_7_45_groupi_n_984 ,csa_tree_add_7_45_groupi_n_946 ,csa_tree_add_7_45_groupi_n_833);
  or csa_tree_add_7_45_groupi_g4333__4733(csa_tree_add_7_45_groupi_n_983 ,csa_tree_add_7_45_groupi_n_788 ,csa_tree_add_7_45_groupi_n_918);
  and csa_tree_add_7_45_groupi_g4334__6161(csa_tree_add_7_45_groupi_n_982 ,csa_tree_add_7_45_groupi_n_952 ,csa_tree_add_7_45_groupi_n_922);
  or csa_tree_add_7_45_groupi_g4335__9315(csa_tree_add_7_45_groupi_n_981 ,csa_tree_add_7_45_groupi_n_795 ,csa_tree_add_7_45_groupi_n_913);
  and csa_tree_add_7_45_groupi_g4336__9945(csa_tree_add_7_45_groupi_n_980 ,csa_tree_add_7_45_groupi_n_750 ,csa_tree_add_7_45_groupi_n_917);
  or csa_tree_add_7_45_groupi_g4337__2883(csa_tree_add_7_45_groupi_n_979 ,csa_tree_add_7_45_groupi_n_802 ,csa_tree_add_7_45_groupi_n_933);
  nor csa_tree_add_7_45_groupi_g4338__2346(csa_tree_add_7_45_groupi_n_978 ,csa_tree_add_7_45_groupi_n_36 ,csa_tree_add_7_45_groupi_n_949);
  or csa_tree_add_7_45_groupi_g4339__1666(csa_tree_add_7_45_groupi_n_977 ,csa_tree_add_7_45_groupi_n_750 ,csa_tree_add_7_45_groupi_n_917);
  or csa_tree_add_7_45_groupi_g4340__7410(csa_tree_add_7_45_groupi_n_1000 ,csa_tree_add_7_45_groupi_n_858 ,csa_tree_add_7_45_groupi_n_930);
  or csa_tree_add_7_45_groupi_g4341__6417(csa_tree_add_7_45_groupi_n_998 ,csa_tree_add_7_45_groupi_n_855 ,csa_tree_add_7_45_groupi_n_911);
  or csa_tree_add_7_45_groupi_g4342__5477(csa_tree_add_7_45_groupi_n_997 ,csa_tree_add_7_45_groupi_n_865 ,csa_tree_add_7_45_groupi_n_912);
  and csa_tree_add_7_45_groupi_g4343__2398(csa_tree_add_7_45_groupi_n_996 ,csa_tree_add_7_45_groupi_n_871 ,csa_tree_add_7_45_groupi_n_934);
  and csa_tree_add_7_45_groupi_g4344__5107(csa_tree_add_7_45_groupi_n_994 ,csa_tree_add_7_45_groupi_n_866 ,csa_tree_add_7_45_groupi_n_929);
  or csa_tree_add_7_45_groupi_g4345__6260(csa_tree_add_7_45_groupi_n_993 ,csa_tree_add_7_45_groupi_n_853 ,csa_tree_add_7_45_groupi_n_936);
  or csa_tree_add_7_45_groupi_g4346__4319(csa_tree_add_7_45_groupi_n_991 ,csa_tree_add_7_45_groupi_n_869 ,csa_tree_add_7_45_groupi_n_925);
  not csa_tree_add_7_45_groupi_g4347(csa_tree_add_7_45_groupi_n_974 ,csa_tree_add_7_45_groupi_n_973);
  not csa_tree_add_7_45_groupi_g4348(csa_tree_add_7_45_groupi_n_972 ,csa_tree_add_7_45_groupi_n_971);
  not csa_tree_add_7_45_groupi_g4349(csa_tree_add_7_45_groupi_n_970 ,csa_tree_add_7_45_groupi_n_969);
  or csa_tree_add_7_45_groupi_g4350__8428(csa_tree_add_7_45_groupi_n_968 ,csa_tree_add_7_45_groupi_n_801 ,csa_tree_add_7_45_groupi_n_907);
  or csa_tree_add_7_45_groupi_g4351__5526(csa_tree_add_7_45_groupi_n_967 ,csa_tree_add_7_45_groupi_n_803 ,csa_tree_add_7_45_groupi_n_903);
  or csa_tree_add_7_45_groupi_g4352__6783(csa_tree_add_7_45_groupi_n_966 ,csa_tree_add_7_45_groupi_n_798 ,csa_tree_add_7_45_groupi_n_905);
  xnor csa_tree_add_7_45_groupi_g4353__3680(out1[2] ,csa_tree_add_7_45_groupi_n_805 ,csa_tree_add_7_45_groupi_n_810);
  xnor csa_tree_add_7_45_groupi_g4354__1617(csa_tree_add_7_45_groupi_n_964 ,csa_tree_add_7_45_groupi_n_800 ,csa_tree_add_7_45_groupi_n_839);
  xnor csa_tree_add_7_45_groupi_g4355__2802(csa_tree_add_7_45_groupi_n_963 ,csa_tree_add_7_45_groupi_n_874 ,csa_tree_add_7_45_groupi_n_821);
  xnor csa_tree_add_7_45_groupi_g4356__1705(csa_tree_add_7_45_groupi_n_962 ,csa_tree_add_7_45_groupi_n_878 ,csa_tree_add_7_45_groupi_n_818);
  xnor csa_tree_add_7_45_groupi_g4357__5122(csa_tree_add_7_45_groupi_n_961 ,csa_tree_add_7_45_groupi_n_882 ,csa_tree_add_7_45_groupi_n_829);
  xnor csa_tree_add_7_45_groupi_g4358__8246(csa_tree_add_7_45_groupi_n_960 ,csa_tree_add_7_45_groupi_n_822 ,csa_tree_add_7_45_groupi_n_793);
  xnor csa_tree_add_7_45_groupi_g4359__7098(csa_tree_add_7_45_groupi_n_959 ,csa_tree_add_7_45_groupi_n_880 ,csa_tree_add_7_45_groupi_n_831);
  xnor csa_tree_add_7_45_groupi_g4360__6131(csa_tree_add_7_45_groupi_n_958 ,csa_tree_add_7_45_groupi_n_755 ,csa_tree_add_7_45_groupi_n_841);
  xnor csa_tree_add_7_45_groupi_g4361__1881(csa_tree_add_7_45_groupi_n_957 ,csa_tree_add_7_45_groupi_n_823 ,csa_tree_add_7_45_groupi_n_4);
  xnor csa_tree_add_7_45_groupi_g4362__5115(csa_tree_add_7_45_groupi_n_956 ,csa_tree_add_7_45_groupi_n_702 ,csa_tree_add_7_45_groupi_n_846);
  xnor csa_tree_add_7_45_groupi_g4363__7482(csa_tree_add_7_45_groupi_n_955 ,csa_tree_add_7_45_groupi_n_765 ,csa_tree_add_7_45_groupi_n_835);
  xnor csa_tree_add_7_45_groupi_g4364__4733(csa_tree_add_7_45_groupi_n_954 ,csa_tree_add_7_45_groupi_n_884 ,csa_tree_add_7_45_groupi_n_816);
  xnor csa_tree_add_7_45_groupi_g4365__6161(csa_tree_add_7_45_groupi_n_953 ,csa_tree_add_7_45_groupi_n_886 ,csa_tree_add_7_45_groupi_n_845);
  xnor csa_tree_add_7_45_groupi_g4366__9315(csa_tree_add_7_45_groupi_n_976 ,csa_tree_add_7_45_groupi_n_733 ,csa_tree_add_7_45_groupi_n_806);
  and csa_tree_add_7_45_groupi_g4367__9945(csa_tree_add_7_45_groupi_n_975 ,csa_tree_add_7_45_groupi_n_851 ,csa_tree_add_7_45_groupi_n_902);
  xnor csa_tree_add_7_45_groupi_g4368__2883(csa_tree_add_7_45_groupi_n_973 ,csa_tree_add_7_45_groupi_n_761 ,csa_tree_add_7_45_groupi_n_808);
  xnor csa_tree_add_7_45_groupi_g4369__2346(csa_tree_add_7_45_groupi_n_971 ,csa_tree_add_7_45_groupi_n_769 ,csa_tree_add_7_45_groupi_n_0);
  xnor csa_tree_add_7_45_groupi_g4370__1666(csa_tree_add_7_45_groupi_n_969 ,csa_tree_add_7_45_groupi_n_616 ,csa_tree_add_7_45_groupi_n_809);
  not csa_tree_add_7_45_groupi_g4371(csa_tree_add_7_45_groupi_n_948 ,csa_tree_add_7_45_groupi_n_949);
  not csa_tree_add_7_45_groupi_g4372(csa_tree_add_7_45_groupi_n_947 ,csa_tree_add_7_45_groupi_n_946);
  nor csa_tree_add_7_45_groupi_g4373__7410(csa_tree_add_7_45_groupi_n_945 ,csa_tree_add_7_45_groupi_n_886 ,csa_tree_add_7_45_groupi_n_845);
  or csa_tree_add_7_45_groupi_g4374__6417(csa_tree_add_7_45_groupi_n_944 ,csa_tree_add_7_45_groupi_n_875 ,csa_tree_add_7_45_groupi_n_838);
  nor csa_tree_add_7_45_groupi_g4375__5477(csa_tree_add_7_45_groupi_n_943 ,csa_tree_add_7_45_groupi_n_876 ,csa_tree_add_7_45_groupi_n_839);
  nor csa_tree_add_7_45_groupi_g4376__2398(csa_tree_add_7_45_groupi_n_942 ,csa_tree_add_7_45_groupi_n_755 ,csa_tree_add_7_45_groupi_n_840);
  or csa_tree_add_7_45_groupi_g4377__5107(csa_tree_add_7_45_groupi_n_941 ,csa_tree_add_7_45_groupi_n_764 ,csa_tree_add_7_45_groupi_n_834);
  or csa_tree_add_7_45_groupi_g4378__6260(csa_tree_add_7_45_groupi_n_940 ,csa_tree_add_7_45_groupi_n_873 ,csa_tree_add_7_45_groupi_n_821);
  or csa_tree_add_7_45_groupi_g4379__4319(csa_tree_add_7_45_groupi_n_939 ,csa_tree_add_7_45_groupi_n_885 ,csa_tree_add_7_45_groupi_n_844);
  nor csa_tree_add_7_45_groupi_g4380__8428(csa_tree_add_7_45_groupi_n_938 ,csa_tree_add_7_45_groupi_n_765 ,csa_tree_add_7_45_groupi_n_835);
  or csa_tree_add_7_45_groupi_g4381__5526(csa_tree_add_7_45_groupi_n_937 ,csa_tree_add_7_45_groupi_n_793 ,csa_tree_add_7_45_groupi_n_822);
  and csa_tree_add_7_45_groupi_g4382__6783(csa_tree_add_7_45_groupi_n_936 ,csa_tree_add_7_45_groupi_n_804 ,csa_tree_add_7_45_groupi_n_852);
  nor csa_tree_add_7_45_groupi_g4383__3680(csa_tree_add_7_45_groupi_n_935 ,csa_tree_add_7_45_groupi_n_874 ,csa_tree_add_7_45_groupi_n_820);
  or csa_tree_add_7_45_groupi_g4384__1617(csa_tree_add_7_45_groupi_n_934 ,csa_tree_add_7_45_groupi_n_774 ,csa_tree_add_7_45_groupi_n_812);
  and csa_tree_add_7_45_groupi_g4385__2802(csa_tree_add_7_45_groupi_n_933 ,csa_tree_add_7_45_groupi_n_3 ,csa_tree_add_7_45_groupi_n_819);
  and csa_tree_add_7_45_groupi_g4386__1705(csa_tree_add_7_45_groupi_n_932 ,csa_tree_add_7_45_groupi_n_793 ,csa_tree_add_7_45_groupi_n_822);
  or csa_tree_add_7_45_groupi_g4387__5122(csa_tree_add_7_45_groupi_n_931 ,csa_tree_add_7_45_groupi_n_877 ,csa_tree_add_7_45_groupi_n_818);
  and csa_tree_add_7_45_groupi_g4388__8246(csa_tree_add_7_45_groupi_n_930 ,csa_tree_add_7_45_groupi_n_741 ,csa_tree_add_7_45_groupi_n_862);
  or csa_tree_add_7_45_groupi_g4389__7098(csa_tree_add_7_45_groupi_n_929 ,csa_tree_add_7_45_groupi_n_864 ,csa_tree_add_7_45_groupi_n_850);
  or csa_tree_add_7_45_groupi_g4390__6131(csa_tree_add_7_45_groupi_n_928 ,csa_tree_add_7_45_groupi_n_3 ,csa_tree_add_7_45_groupi_n_819);
  nor csa_tree_add_7_45_groupi_g4391__1881(csa_tree_add_7_45_groupi_n_927 ,csa_tree_add_7_45_groupi_n_878 ,csa_tree_add_7_45_groupi_n_817);
  nor csa_tree_add_7_45_groupi_g4392__5115(csa_tree_add_7_45_groupi_n_926 ,csa_tree_add_7_45_groupi_n_882 ,csa_tree_add_7_45_groupi_n_828);
  and csa_tree_add_7_45_groupi_g4393__7482(csa_tree_add_7_45_groupi_n_925 ,csa_tree_add_7_45_groupi_n_776 ,csa_tree_add_7_45_groupi_n_859);
  and csa_tree_add_7_45_groupi_g4394__4733(csa_tree_add_7_45_groupi_n_924 ,csa_tree_add_7_45_groupi_n_702 ,csa_tree_add_7_45_groupi_n_846);
  or csa_tree_add_7_45_groupi_g4395__6161(csa_tree_add_7_45_groupi_n_923 ,csa_tree_add_7_45_groupi_n_881 ,csa_tree_add_7_45_groupi_n_829);
  or csa_tree_add_7_45_groupi_g4396__9315(csa_tree_add_7_45_groupi_n_922 ,csa_tree_add_7_45_groupi_n_702 ,csa_tree_add_7_45_groupi_n_846);
  or csa_tree_add_7_45_groupi_g4397__9945(csa_tree_add_7_45_groupi_n_921 ,csa_tree_add_7_45_groupi_n_883 ,csa_tree_add_7_45_groupi_n_816);
  nor csa_tree_add_7_45_groupi_g4398__2883(csa_tree_add_7_45_groupi_n_920 ,csa_tree_add_7_45_groupi_n_884 ,csa_tree_add_7_45_groupi_n_815);
  or csa_tree_add_7_45_groupi_g4399__2346(csa_tree_add_7_45_groupi_n_952 ,csa_tree_add_7_45_groupi_n_782 ,csa_tree_add_7_45_groupi_n_856);
  and csa_tree_add_7_45_groupi_g4400__1666(csa_tree_add_7_45_groupi_n_951 ,csa_tree_add_7_45_groupi_n_655 ,csa_tree_add_7_45_groupi_n_868);
  and csa_tree_add_7_45_groupi_g4401__7410(csa_tree_add_7_45_groupi_n_950 ,csa_tree_add_7_45_groupi_n_652 ,csa_tree_add_7_45_groupi_n_863);
  and csa_tree_add_7_45_groupi_g4402__6417(csa_tree_add_7_45_groupi_n_949 ,csa_tree_add_7_45_groupi_n_725 ,csa_tree_add_7_45_groupi_n_860);
  or csa_tree_add_7_45_groupi_g4403__5477(csa_tree_add_7_45_groupi_n_946 ,csa_tree_add_7_45_groupi_n_778 ,csa_tree_add_7_45_groupi_n_870);
  not csa_tree_add_7_45_groupi_g4404(csa_tree_add_7_45_groupi_n_918 ,csa_tree_add_7_45_groupi_n_919);
  or csa_tree_add_7_45_groupi_g4405__2398(csa_tree_add_7_45_groupi_n_915 ,csa_tree_add_7_45_groupi_n_754 ,csa_tree_add_7_45_groupi_n_841);
  or csa_tree_add_7_45_groupi_g4406__5107(csa_tree_add_7_45_groupi_n_914 ,csa_tree_add_7_45_groupi_n_759 ,csa_tree_add_7_45_groupi_n_826);
  nor csa_tree_add_7_45_groupi_g4407__6260(csa_tree_add_7_45_groupi_n_913 ,csa_tree_add_7_45_groupi_n_760 ,csa_tree_add_7_45_groupi_n_827);
  and csa_tree_add_7_45_groupi_g4408__4319(csa_tree_add_7_45_groupi_n_912 ,csa_tree_add_7_45_groupi_n_872 ,csa_tree_add_7_45_groupi_n_887);
  nor csa_tree_add_7_45_groupi_g4409__8428(csa_tree_add_7_45_groupi_n_911 ,csa_tree_add_7_45_groupi_n_797 ,csa_tree_add_7_45_groupi_n_854);
  nor csa_tree_add_7_45_groupi_g4410__5526(csa_tree_add_7_45_groupi_n_910 ,csa_tree_add_7_45_groupi_n_824 ,csa_tree_add_7_45_groupi_n_4);
  and csa_tree_add_7_45_groupi_g4411__6783(csa_tree_add_7_45_groupi_n_909 ,csa_tree_add_7_45_groupi_n_824 ,csa_tree_add_7_45_groupi_n_4);
  or csa_tree_add_7_45_groupi_g4412__3680(csa_tree_add_7_45_groupi_n_908 ,csa_tree_add_7_45_groupi_n_751 ,csa_tree_add_7_45_groupi_n_813);
  nor csa_tree_add_7_45_groupi_g4413__1617(csa_tree_add_7_45_groupi_n_907 ,csa_tree_add_7_45_groupi_n_752 ,csa_tree_add_7_45_groupi_n_814);
  or csa_tree_add_7_45_groupi_g4414__2802(csa_tree_add_7_45_groupi_n_906 ,csa_tree_add_7_45_groupi_n_763 ,csa_tree_add_7_45_groupi_n_847);
  nor csa_tree_add_7_45_groupi_g4415__1705(csa_tree_add_7_45_groupi_n_905 ,csa_tree_add_7_45_groupi_n_762 ,csa_tree_add_7_45_groupi_n_848);
  or csa_tree_add_7_45_groupi_g4416__5122(csa_tree_add_7_45_groupi_n_904 ,csa_tree_add_7_45_groupi_n_758 ,csa_tree_add_7_45_groupi_n_842);
  nor csa_tree_add_7_45_groupi_g4417__8246(csa_tree_add_7_45_groupi_n_903 ,csa_tree_add_7_45_groupi_n_757 ,csa_tree_add_7_45_groupi_n_843);
  or csa_tree_add_7_45_groupi_g4418__7098(csa_tree_add_7_45_groupi_n_902 ,csa_tree_add_7_45_groupi_n_740 ,csa_tree_add_7_45_groupi_n_857);
  or csa_tree_add_7_45_groupi_g4419__6131(csa_tree_add_7_45_groupi_n_901 ,csa_tree_add_7_45_groupi_n_879 ,csa_tree_add_7_45_groupi_n_830);
  nor csa_tree_add_7_45_groupi_g4420__1881(csa_tree_add_7_45_groupi_n_900 ,csa_tree_add_7_45_groupi_n_880 ,csa_tree_add_7_45_groupi_n_831);
  xnor csa_tree_add_7_45_groupi_g4421__5115(csa_tree_add_7_45_groupi_n_899 ,csa_tree_add_7_45_groupi_n_801 ,csa_tree_add_7_45_groupi_n_752);
  xnor csa_tree_add_7_45_groupi_g4422__7482(csa_tree_add_7_45_groupi_n_898 ,csa_tree_add_7_45_groupi_n_758 ,csa_tree_add_7_45_groupi_n_803);
  xnor csa_tree_add_7_45_groupi_g4423__4733(csa_tree_add_7_45_groupi_n_897 ,csa_tree_add_7_45_groupi_n_617 ,csa_tree_add_7_45_groupi_n_774);
  xnor csa_tree_add_7_45_groupi_g4424__6161(csa_tree_add_7_45_groupi_n_896 ,csa_tree_add_7_45_groupi_n_796 ,csa_tree_add_7_45_groupi_n_756);
  xnor csa_tree_add_7_45_groupi_g4425__9315(csa_tree_add_7_45_groupi_n_895 ,csa_tree_add_7_45_groupi_n_619 ,csa_tree_add_7_45_groupi_n_790);
  xnor csa_tree_add_7_45_groupi_g4426__9945(csa_tree_add_7_45_groupi_n_894 ,csa_tree_add_7_45_groupi_n_771 ,csa_tree_add_7_45_groupi_n_426);
  xnor csa_tree_add_7_45_groupi_g4427__2883(csa_tree_add_7_45_groupi_n_893 ,csa_tree_add_7_45_groupi_n_622 ,csa_tree_add_7_45_groupi_n_2);
  xnor csa_tree_add_7_45_groupi_g4428__2346(csa_tree_add_7_45_groupi_n_892 ,csa_tree_add_7_45_groupi_n_795 ,csa_tree_add_7_45_groupi_n_760);
  xnor csa_tree_add_7_45_groupi_g4429__1666(csa_tree_add_7_45_groupi_n_891 ,csa_tree_add_7_45_groupi_n_773 ,csa_tree_add_7_45_groupi_n_767);
  xnor csa_tree_add_7_45_groupi_g4430__7410(csa_tree_add_7_45_groupi_n_890 ,csa_tree_add_7_45_groupi_n_792 ,csa_tree_add_7_45_groupi_n_749);
  xor csa_tree_add_7_45_groupi_g4431__6417(csa_tree_add_7_45_groupi_n_889 ,csa_tree_add_7_45_groupi_n_802 ,csa_tree_add_7_45_groupi_n_3);
  xnor csa_tree_add_7_45_groupi_g4432__5477(csa_tree_add_7_45_groupi_n_888 ,csa_tree_add_7_45_groupi_n_763 ,csa_tree_add_7_45_groupi_n_798);
  xnor csa_tree_add_7_45_groupi_g4433__2398(csa_tree_add_7_45_groupi_n_919 ,csa_tree_add_7_45_groupi_n_777 ,csa_tree_add_7_45_groupi_n_679);
  xnor csa_tree_add_7_45_groupi_g4434__5107(csa_tree_add_7_45_groupi_n_917 ,csa_tree_add_7_45_groupi_n_775 ,csa_tree_add_7_45_groupi_n_691);
  xnor csa_tree_add_7_45_groupi_g4435__6260(csa_tree_add_7_45_groupi_n_916 ,csa_tree_add_7_45_groupi_n_794 ,csa_tree_add_7_45_groupi_n_743);
  not csa_tree_add_7_45_groupi_g4436(csa_tree_add_7_45_groupi_n_885 ,csa_tree_add_7_45_groupi_n_886);
  not csa_tree_add_7_45_groupi_g4437(csa_tree_add_7_45_groupi_n_883 ,csa_tree_add_7_45_groupi_n_884);
  not csa_tree_add_7_45_groupi_g4438(csa_tree_add_7_45_groupi_n_881 ,csa_tree_add_7_45_groupi_n_882);
  not csa_tree_add_7_45_groupi_g4439(csa_tree_add_7_45_groupi_n_880 ,csa_tree_add_7_45_groupi_n_879);
  not csa_tree_add_7_45_groupi_g4440(csa_tree_add_7_45_groupi_n_877 ,csa_tree_add_7_45_groupi_n_878);
  not csa_tree_add_7_45_groupi_g4441(csa_tree_add_7_45_groupi_n_876 ,csa_tree_add_7_45_groupi_n_875);
  not csa_tree_add_7_45_groupi_g4442(csa_tree_add_7_45_groupi_n_873 ,csa_tree_add_7_45_groupi_n_874);
  or csa_tree_add_7_45_groupi_g4443__4319(csa_tree_add_7_45_groupi_n_872 ,csa_tree_add_7_45_groupi_n_619 ,csa_tree_add_7_45_groupi_n_790);
  or csa_tree_add_7_45_groupi_g4444__8428(csa_tree_add_7_45_groupi_n_871 ,csa_tree_add_7_45_groupi_n_618 ,csa_tree_add_7_45_groupi_n_753);
  and csa_tree_add_7_45_groupi_g4445__5526(csa_tree_add_7_45_groupi_n_870 ,csa_tree_add_7_45_groupi_n_733 ,csa_tree_add_7_45_groupi_n_787);
  and csa_tree_add_7_45_groupi_g4446__6783(csa_tree_add_7_45_groupi_n_869 ,csa_tree_add_7_45_groupi_n_52 ,csa_tree_add_7_45_groupi_n_771);
  or csa_tree_add_7_45_groupi_g4447__3680(csa_tree_add_7_45_groupi_n_868 ,csa_tree_add_7_45_groupi_n_644 ,csa_tree_add_7_45_groupi_n_775);
  nor csa_tree_add_7_45_groupi_g4448__1617(csa_tree_add_7_45_groupi_n_867 ,csa_tree_add_7_45_groupi_n_772 ,csa_tree_add_7_45_groupi_n_767);
  or csa_tree_add_7_45_groupi_g4449__2802(csa_tree_add_7_45_groupi_n_866 ,csa_tree_add_7_45_groupi_n_791 ,csa_tree_add_7_45_groupi_n_749);
  and csa_tree_add_7_45_groupi_g4450__1705(csa_tree_add_7_45_groupi_n_865 ,csa_tree_add_7_45_groupi_n_619 ,csa_tree_add_7_45_groupi_n_790);
  nor csa_tree_add_7_45_groupi_g4451__5122(csa_tree_add_7_45_groupi_n_864 ,csa_tree_add_7_45_groupi_n_792 ,csa_tree_add_7_45_groupi_n_748);
  or csa_tree_add_7_45_groupi_g4452__8246(csa_tree_add_7_45_groupi_n_863 ,csa_tree_add_7_45_groupi_n_608 ,csa_tree_add_7_45_groupi_n_777);
  or csa_tree_add_7_45_groupi_g4453__7098(csa_tree_add_7_45_groupi_n_862 ,csa_tree_add_7_45_groupi_n_730 ,csa_tree_add_7_45_groupi_n_1);
  or csa_tree_add_7_45_groupi_g4454__6131(csa_tree_add_7_45_groupi_n_861 ,csa_tree_add_7_45_groupi_n_773 ,csa_tree_add_7_45_groupi_n_766);
  or csa_tree_add_7_45_groupi_g4455__1881(csa_tree_add_7_45_groupi_n_860 ,csa_tree_add_7_45_groupi_n_714 ,csa_tree_add_7_45_groupi_n_794);
  or csa_tree_add_7_45_groupi_g4456__5115(csa_tree_add_7_45_groupi_n_859 ,csa_tree_add_7_45_groupi_n_426 ,csa_tree_add_7_45_groupi_n_771);
  nor csa_tree_add_7_45_groupi_g4457__7482(csa_tree_add_7_45_groupi_n_858 ,csa_tree_add_7_45_groupi_n_731 ,csa_tree_add_7_45_groupi_n_761);
  nor csa_tree_add_7_45_groupi_g4458__4733(csa_tree_add_7_45_groupi_n_857 ,csa_tree_add_7_45_groupi_n_705 ,csa_tree_add_7_45_groupi_n_769);
  nor csa_tree_add_7_45_groupi_g4459__6161(csa_tree_add_7_45_groupi_n_856 ,csa_tree_add_7_45_groupi_n_805 ,csa_tree_add_7_45_groupi_n_784);
  and csa_tree_add_7_45_groupi_g4460__9315(csa_tree_add_7_45_groupi_n_855 ,csa_tree_add_7_45_groupi_n_770 ,csa_tree_add_7_45_groupi_n_756);
  nor csa_tree_add_7_45_groupi_g4461__9945(csa_tree_add_7_45_groupi_n_854 ,csa_tree_add_7_45_groupi_n_770 ,csa_tree_add_7_45_groupi_n_756);
  and csa_tree_add_7_45_groupi_g4462__2883(csa_tree_add_7_45_groupi_n_853 ,csa_tree_add_7_45_groupi_n_622 ,csa_tree_add_7_45_groupi_n_2);
  or csa_tree_add_7_45_groupi_g4463__2346(csa_tree_add_7_45_groupi_n_852 ,csa_tree_add_7_45_groupi_n_622 ,csa_tree_add_7_45_groupi_n_2);
  or csa_tree_add_7_45_groupi_g4464__1666(csa_tree_add_7_45_groupi_n_851 ,csa_tree_add_7_45_groupi_n_60 ,csa_tree_add_7_45_groupi_n_768);
  or csa_tree_add_7_45_groupi_g4465__7410(csa_tree_add_7_45_groupi_n_887 ,csa_tree_add_7_45_groupi_n_701 ,csa_tree_add_7_45_groupi_n_745);
  or csa_tree_add_7_45_groupi_g4466__6417(csa_tree_add_7_45_groupi_n_886 ,csa_tree_add_7_45_groupi_n_593 ,csa_tree_add_7_45_groupi_n_779);
  or csa_tree_add_7_45_groupi_g4467__5477(csa_tree_add_7_45_groupi_n_884 ,csa_tree_add_7_45_groupi_n_626 ,csa_tree_add_7_45_groupi_n_746);
  or csa_tree_add_7_45_groupi_g4468__2398(csa_tree_add_7_45_groupi_n_882 ,csa_tree_add_7_45_groupi_n_628 ,csa_tree_add_7_45_groupi_n_783);
  and csa_tree_add_7_45_groupi_g4469__5107(csa_tree_add_7_45_groupi_n_879 ,csa_tree_add_7_45_groupi_n_605 ,csa_tree_add_7_45_groupi_n_747);
  or csa_tree_add_7_45_groupi_g4470__6260(csa_tree_add_7_45_groupi_n_878 ,csa_tree_add_7_45_groupi_n_637 ,csa_tree_add_7_45_groupi_n_781);
  and csa_tree_add_7_45_groupi_g4471__4319(csa_tree_add_7_45_groupi_n_875 ,csa_tree_add_7_45_groupi_n_666 ,csa_tree_add_7_45_groupi_n_785);
  or csa_tree_add_7_45_groupi_g4472__8428(csa_tree_add_7_45_groupi_n_874 ,csa_tree_add_7_45_groupi_n_656 ,csa_tree_add_7_45_groupi_n_780);
  not csa_tree_add_7_45_groupi_g4473(csa_tree_add_7_45_groupi_n_850 ,csa_tree_add_7_45_groupi_n_849);
  not csa_tree_add_7_45_groupi_g4474(csa_tree_add_7_45_groupi_n_847 ,csa_tree_add_7_45_groupi_n_848);
  not csa_tree_add_7_45_groupi_g4475(csa_tree_add_7_45_groupi_n_844 ,csa_tree_add_7_45_groupi_n_845);
  not csa_tree_add_7_45_groupi_g4476(csa_tree_add_7_45_groupi_n_842 ,csa_tree_add_7_45_groupi_n_843);
  not csa_tree_add_7_45_groupi_g4477(csa_tree_add_7_45_groupi_n_841 ,csa_tree_add_7_45_groupi_n_840);
  not csa_tree_add_7_45_groupi_g4478(csa_tree_add_7_45_groupi_n_838 ,csa_tree_add_7_45_groupi_n_839);
  not csa_tree_add_7_45_groupi_g4479(csa_tree_add_7_45_groupi_n_837 ,csa_tree_add_7_45_groupi_n_836);
  not csa_tree_add_7_45_groupi_g4480(csa_tree_add_7_45_groupi_n_834 ,csa_tree_add_7_45_groupi_n_835);
  not csa_tree_add_7_45_groupi_g4481(csa_tree_add_7_45_groupi_n_832 ,csa_tree_add_7_45_groupi_n_833);
  not csa_tree_add_7_45_groupi_g4482(csa_tree_add_7_45_groupi_n_831 ,csa_tree_add_7_45_groupi_n_830);
  not csa_tree_add_7_45_groupi_g4483(csa_tree_add_7_45_groupi_n_828 ,csa_tree_add_7_45_groupi_n_829);
  not csa_tree_add_7_45_groupi_g4484(csa_tree_add_7_45_groupi_n_826 ,csa_tree_add_7_45_groupi_n_827);
  not csa_tree_add_7_45_groupi_g4485(csa_tree_add_7_45_groupi_n_824 ,csa_tree_add_7_45_groupi_n_823);
  not csa_tree_add_7_45_groupi_g4486(csa_tree_add_7_45_groupi_n_820 ,csa_tree_add_7_45_groupi_n_821);
  not csa_tree_add_7_45_groupi_g4487(csa_tree_add_7_45_groupi_n_817 ,csa_tree_add_7_45_groupi_n_818);
  not csa_tree_add_7_45_groupi_g4488(csa_tree_add_7_45_groupi_n_815 ,csa_tree_add_7_45_groupi_n_816);
  not csa_tree_add_7_45_groupi_g4489(csa_tree_add_7_45_groupi_n_813 ,csa_tree_add_7_45_groupi_n_814);
  and csa_tree_add_7_45_groupi_g4490__5526(csa_tree_add_7_45_groupi_n_812 ,csa_tree_add_7_45_groupi_n_618 ,csa_tree_add_7_45_groupi_n_753);
  xnor csa_tree_add_7_45_groupi_g4491__6783(out1[1] ,csa_tree_add_7_45_groupi_n_410 ,csa_tree_add_7_45_groupi_n_688);
  xnor csa_tree_add_7_45_groupi_g4492__3680(csa_tree_add_7_45_groupi_n_810 ,csa_tree_add_7_45_groupi_n_370 ,csa_tree_add_7_45_groupi_n_703);
  xnor csa_tree_add_7_45_groupi_g4493__1617(csa_tree_add_7_45_groupi_n_809 ,csa_tree_add_7_45_groupi_n_560 ,csa_tree_add_7_45_groupi_n_739);
  xnor csa_tree_add_7_45_groupi_g4494__2802(csa_tree_add_7_45_groupi_n_808 ,csa_tree_add_7_45_groupi_n_741 ,csa_tree_add_7_45_groupi_n_731);
  xnor csa_tree_add_7_45_groupi_g4495__1705(csa_tree_add_7_45_groupi_n_807 ,csa_tree_add_7_45_groupi_n_732 ,csa_tree_add_7_45_groupi_n_51);
  xnor csa_tree_add_7_45_groupi_g4496__5122(csa_tree_add_7_45_groupi_n_806 ,csa_tree_add_7_45_groupi_n_707 ,csa_tree_add_7_45_groupi_n_519);
  xnor csa_tree_add_7_45_groupi_g4498__8246(csa_tree_add_7_45_groupi_n_849 ,csa_tree_add_7_45_groupi_n_623 ,csa_tree_add_7_45_groupi_n_689);
  xnor csa_tree_add_7_45_groupi_g4499__7098(csa_tree_add_7_45_groupi_n_848 ,csa_tree_add_7_45_groupi_n_503 ,csa_tree_add_7_45_groupi_n_682);
  xnor csa_tree_add_7_45_groupi_g4500__6131(csa_tree_add_7_45_groupi_n_846 ,csa_tree_add_7_45_groupi_n_624 ,csa_tree_add_7_45_groupi_n_676);
  xnor csa_tree_add_7_45_groupi_g4501__1881(csa_tree_add_7_45_groupi_n_845 ,csa_tree_add_7_45_groupi_n_742 ,csa_tree_add_7_45_groupi_n_674);
  xnor csa_tree_add_7_45_groupi_g4502__5115(csa_tree_add_7_45_groupi_n_843 ,csa_tree_add_7_45_groupi_n_481 ,csa_tree_add_7_45_groupi_n_681);
  xnor csa_tree_add_7_45_groupi_g4504__7482(csa_tree_add_7_45_groupi_n_840 ,csa_tree_add_7_45_groupi_n_571 ,csa_tree_add_7_45_groupi_n_678);
  xnor csa_tree_add_7_45_groupi_g4505__4733(csa_tree_add_7_45_groupi_n_839 ,csa_tree_add_7_45_groupi_n_466 ,csa_tree_add_7_45_groupi_n_697);
  xnor csa_tree_add_7_45_groupi_g4506__6161(csa_tree_add_7_45_groupi_n_836 ,csa_tree_add_7_45_groupi_n_735 ,csa_tree_add_7_45_groupi_n_675);
  xnor csa_tree_add_7_45_groupi_g4507__9315(csa_tree_add_7_45_groupi_n_835 ,csa_tree_add_7_45_groupi_n_523 ,csa_tree_add_7_45_groupi_n_693);
  xnor csa_tree_add_7_45_groupi_g4508__9945(csa_tree_add_7_45_groupi_n_833 ,csa_tree_add_7_45_groupi_n_524 ,csa_tree_add_7_45_groupi_n_695);
  xnor csa_tree_add_7_45_groupi_g4509__2883(csa_tree_add_7_45_groupi_n_830 ,csa_tree_add_7_45_groupi_n_708 ,csa_tree_add_7_45_groupi_n_686);
  xnor csa_tree_add_7_45_groupi_g4510__2346(csa_tree_add_7_45_groupi_n_829 ,csa_tree_add_7_45_groupi_n_494 ,csa_tree_add_7_45_groupi_n_692);
  xnor csa_tree_add_7_45_groupi_g4511__1666(csa_tree_add_7_45_groupi_n_827 ,csa_tree_add_7_45_groupi_n_499 ,csa_tree_add_7_45_groupi_n_685);
  xnor csa_tree_add_7_45_groupi_g4512__7410(csa_tree_add_7_45_groupi_n_825 ,csa_tree_add_7_45_groupi_n_625 ,csa_tree_add_7_45_groupi_n_696);
  xnor csa_tree_add_7_45_groupi_g4513__6417(csa_tree_add_7_45_groupi_n_823 ,csa_tree_add_7_45_groupi_n_500 ,csa_tree_add_7_45_groupi_n_684);
  xnor csa_tree_add_7_45_groupi_g4514__5477(csa_tree_add_7_45_groupi_n_822 ,csa_tree_add_7_45_groupi_n_520 ,csa_tree_add_7_45_groupi_n_677);
  xnor csa_tree_add_7_45_groupi_g4515__2398(csa_tree_add_7_45_groupi_n_821 ,csa_tree_add_7_45_groupi_n_734 ,csa_tree_add_7_45_groupi_n_694);
  xnor csa_tree_add_7_45_groupi_g4516__5107(csa_tree_add_7_45_groupi_n_819 ,csa_tree_add_7_45_groupi_n_409 ,csa_tree_add_7_45_groupi_n_680);
  xnor csa_tree_add_7_45_groupi_g4517__6260(csa_tree_add_7_45_groupi_n_818 ,csa_tree_add_7_45_groupi_n_736 ,csa_tree_add_7_45_groupi_n_687);
  xnor csa_tree_add_7_45_groupi_g4518__4319(csa_tree_add_7_45_groupi_n_816 ,csa_tree_add_7_45_groupi_n_738 ,csa_tree_add_7_45_groupi_n_690);
  xnor csa_tree_add_7_45_groupi_g4519__8428(csa_tree_add_7_45_groupi_n_814 ,csa_tree_add_7_45_groupi_n_471 ,csa_tree_add_7_45_groupi_n_683);
  not csa_tree_add_7_45_groupi_g4520(csa_tree_add_7_45_groupi_n_797 ,csa_tree_add_7_45_groupi_n_796);
  not csa_tree_add_7_45_groupi_g4521(csa_tree_add_7_45_groupi_n_791 ,csa_tree_add_7_45_groupi_n_792);
  not csa_tree_add_7_45_groupi_g4522(csa_tree_add_7_45_groupi_n_788 ,csa_tree_add_7_45_groupi_n_789);
  or csa_tree_add_7_45_groupi_g4523__5526(csa_tree_add_7_45_groupi_n_787 ,csa_tree_add_7_45_groupi_n_518 ,csa_tree_add_7_45_groupi_n_706);
  or csa_tree_add_7_45_groupi_g4524__6783(csa_tree_add_7_45_groupi_n_786 ,csa_tree_add_7_45_groupi_n_51 ,csa_tree_add_7_45_groupi_n_732);
  or csa_tree_add_7_45_groupi_g4525__3680(csa_tree_add_7_45_groupi_n_785 ,csa_tree_add_7_45_groupi_n_665 ,csa_tree_add_7_45_groupi_n_735);
  and csa_tree_add_7_45_groupi_g4526__1617(csa_tree_add_7_45_groupi_n_784 ,csa_tree_add_7_45_groupi_n_371 ,csa_tree_add_7_45_groupi_n_703);
  and csa_tree_add_7_45_groupi_g4527__2802(csa_tree_add_7_45_groupi_n_783 ,csa_tree_add_7_45_groupi_n_614 ,csa_tree_add_7_45_groupi_n_742);
  nor csa_tree_add_7_45_groupi_g4528__1705(csa_tree_add_7_45_groupi_n_782 ,csa_tree_add_7_45_groupi_n_371 ,csa_tree_add_7_45_groupi_n_703);
  and csa_tree_add_7_45_groupi_g4529__5122(csa_tree_add_7_45_groupi_n_781 ,csa_tree_add_7_45_groupi_n_609 ,csa_tree_add_7_45_groupi_n_738);
  and csa_tree_add_7_45_groupi_g4530__8246(csa_tree_add_7_45_groupi_n_780 ,csa_tree_add_7_45_groupi_n_612 ,csa_tree_add_7_45_groupi_n_736);
  and csa_tree_add_7_45_groupi_g4531__7098(csa_tree_add_7_45_groupi_n_779 ,csa_tree_add_7_45_groupi_n_671 ,csa_tree_add_7_45_groupi_n_734);
  nor csa_tree_add_7_45_groupi_g4532__6131(csa_tree_add_7_45_groupi_n_778 ,csa_tree_add_7_45_groupi_n_519 ,csa_tree_add_7_45_groupi_n_707);
  and csa_tree_add_7_45_groupi_g4533__1881(csa_tree_add_7_45_groupi_n_805 ,csa_tree_add_7_45_groupi_n_673 ,csa_tree_add_7_45_groupi_n_716);
  or csa_tree_add_7_45_groupi_g4534__5115(csa_tree_add_7_45_groupi_n_804 ,csa_tree_add_7_45_groupi_n_649 ,csa_tree_add_7_45_groupi_n_724);
  and csa_tree_add_7_45_groupi_g4535__7482(csa_tree_add_7_45_groupi_n_803 ,csa_tree_add_7_45_groupi_n_639 ,csa_tree_add_7_45_groupi_n_715);
  and csa_tree_add_7_45_groupi_g4536__4733(csa_tree_add_7_45_groupi_n_802 ,csa_tree_add_7_45_groupi_n_634 ,csa_tree_add_7_45_groupi_n_719);
  and csa_tree_add_7_45_groupi_g4537__6161(csa_tree_add_7_45_groupi_n_801 ,csa_tree_add_7_45_groupi_n_664 ,csa_tree_add_7_45_groupi_n_728);
  and csa_tree_add_7_45_groupi_g4538__9315(csa_tree_add_7_45_groupi_n_800 ,csa_tree_add_7_45_groupi_n_662 ,csa_tree_add_7_45_groupi_n_727);
  and csa_tree_add_7_45_groupi_g4539__9945(csa_tree_add_7_45_groupi_n_799 ,csa_tree_add_7_45_groupi_n_654 ,csa_tree_add_7_45_groupi_n_726);
  and csa_tree_add_7_45_groupi_g4540__2883(csa_tree_add_7_45_groupi_n_798 ,csa_tree_add_7_45_groupi_n_646 ,csa_tree_add_7_45_groupi_n_722);
  or csa_tree_add_7_45_groupi_g4541__2346(csa_tree_add_7_45_groupi_n_796 ,csa_tree_add_7_45_groupi_n_607 ,csa_tree_add_7_45_groupi_n_713);
  and csa_tree_add_7_45_groupi_g4542__1666(csa_tree_add_7_45_groupi_n_795 ,csa_tree_add_7_45_groupi_n_595 ,csa_tree_add_7_45_groupi_n_717);
  and csa_tree_add_7_45_groupi_g4543__7410(csa_tree_add_7_45_groupi_n_794 ,csa_tree_add_7_45_groupi_n_610 ,csa_tree_add_7_45_groupi_n_721);
  and csa_tree_add_7_45_groupi_g4544__6417(csa_tree_add_7_45_groupi_n_793 ,csa_tree_add_7_45_groupi_n_667 ,csa_tree_add_7_45_groupi_n_723);
  or csa_tree_add_7_45_groupi_g4545__5477(csa_tree_add_7_45_groupi_n_792 ,csa_tree_add_7_45_groupi_n_638 ,csa_tree_add_7_45_groupi_n_720);
  or csa_tree_add_7_45_groupi_g4546__2398(csa_tree_add_7_45_groupi_n_790 ,csa_tree_add_7_45_groupi_n_606 ,csa_tree_add_7_45_groupi_n_712);
  or csa_tree_add_7_45_groupi_g4547__5107(csa_tree_add_7_45_groupi_n_789 ,csa_tree_add_7_45_groupi_n_632 ,csa_tree_add_7_45_groupi_n_718);
  not csa_tree_add_7_45_groupi_g4548(csa_tree_add_7_45_groupi_n_772 ,csa_tree_add_7_45_groupi_n_773);
  not csa_tree_add_7_45_groupi_g4549(csa_tree_add_7_45_groupi_n_769 ,csa_tree_add_7_45_groupi_n_768);
  not csa_tree_add_7_45_groupi_g4550(csa_tree_add_7_45_groupi_n_766 ,csa_tree_add_7_45_groupi_n_767);
  not csa_tree_add_7_45_groupi_g4551(csa_tree_add_7_45_groupi_n_765 ,csa_tree_add_7_45_groupi_n_764);
  not csa_tree_add_7_45_groupi_g4552(csa_tree_add_7_45_groupi_n_763 ,csa_tree_add_7_45_groupi_n_762);
  not csa_tree_add_7_45_groupi_g4553(csa_tree_add_7_45_groupi_n_761 ,csa_tree_add_7_45_groupi_n_1);
  not csa_tree_add_7_45_groupi_g4554(csa_tree_add_7_45_groupi_n_760 ,csa_tree_add_7_45_groupi_n_759);
  not csa_tree_add_7_45_groupi_g4555(csa_tree_add_7_45_groupi_n_758 ,csa_tree_add_7_45_groupi_n_757);
  not csa_tree_add_7_45_groupi_g4556(csa_tree_add_7_45_groupi_n_754 ,csa_tree_add_7_45_groupi_n_755);
  not csa_tree_add_7_45_groupi_g4557(csa_tree_add_7_45_groupi_n_752 ,csa_tree_add_7_45_groupi_n_751);
  not csa_tree_add_7_45_groupi_g4558(csa_tree_add_7_45_groupi_n_748 ,csa_tree_add_7_45_groupi_n_749);
  or csa_tree_add_7_45_groupi_g4559__6260(csa_tree_add_7_45_groupi_n_747 ,csa_tree_add_7_45_groupi_n_603 ,csa_tree_add_7_45_groupi_n_737);
  and csa_tree_add_7_45_groupi_g4560__4319(csa_tree_add_7_45_groupi_n_746 ,csa_tree_add_7_45_groupi_n_708 ,csa_tree_add_7_45_groupi_n_651);
  and csa_tree_add_7_45_groupi_g4561__8428(csa_tree_add_7_45_groupi_n_745 ,csa_tree_add_7_45_groupi_n_739 ,csa_tree_add_7_45_groupi_n_710);
  and csa_tree_add_7_45_groupi_g4562__5526(csa_tree_add_7_45_groupi_n_744 ,csa_tree_add_7_45_groupi_n_159 ,csa_tree_add_7_45_groupi_n_732);
  xnor csa_tree_add_7_45_groupi_g4563__6783(csa_tree_add_7_45_groupi_n_743 ,csa_tree_add_7_45_groupi_n_436 ,csa_tree_add_7_45_groupi_n_621);
  xnor csa_tree_add_7_45_groupi_g4564__3680(csa_tree_add_7_45_groupi_n_777 ,csa_tree_add_7_45_groupi_n_482 ,csa_tree_add_7_45_groupi_n_588);
  or csa_tree_add_7_45_groupi_g4565__1617(csa_tree_add_7_45_groupi_n_776 ,csa_tree_add_7_45_groupi_n_597 ,csa_tree_add_7_45_groupi_n_700);
  xnor csa_tree_add_7_45_groupi_g4566__2802(csa_tree_add_7_45_groupi_n_775 ,csa_tree_add_7_45_groupi_n_504 ,csa_tree_add_7_45_groupi_n_587);
  and csa_tree_add_7_45_groupi_g4567__1705(csa_tree_add_7_45_groupi_n_774 ,csa_tree_add_7_45_groupi_n_596 ,csa_tree_add_7_45_groupi_n_711);
  xnor csa_tree_add_7_45_groupi_g4568__5122(csa_tree_add_7_45_groupi_n_773 ,csa_tree_add_7_45_groupi_n_562 ,csa_tree_add_7_45_groupi_n_577);
  xnor csa_tree_add_7_45_groupi_g4569__8246(csa_tree_add_7_45_groupi_n_771 ,csa_tree_add_7_45_groupi_n_467 ,csa_tree_add_7_45_groupi_n_584);
  xnor csa_tree_add_7_45_groupi_g4570__7098(csa_tree_add_7_45_groupi_n_770 ,csa_tree_add_7_45_groupi_n_437 ,csa_tree_add_7_45_groupi_n_590);
  xnor csa_tree_add_7_45_groupi_g4571__6131(csa_tree_add_7_45_groupi_n_768 ,csa_tree_add_7_45_groupi_n_400 ,csa_tree_add_7_45_groupi_n_579);
  and csa_tree_add_7_45_groupi_g4572__1881(csa_tree_add_7_45_groupi_n_767 ,csa_tree_add_7_45_groupi_n_642 ,csa_tree_add_7_45_groupi_n_699);
  xnor csa_tree_add_7_45_groupi_g4573__5115(csa_tree_add_7_45_groupi_n_764 ,csa_tree_add_7_45_groupi_n_416 ,csa_tree_add_7_45_groupi_n_582);
  xnor csa_tree_add_7_45_groupi_g4575__7482(csa_tree_add_7_45_groupi_n_762 ,csa_tree_add_7_45_groupi_n_403 ,csa_tree_add_7_45_groupi_n_581);
  xnor csa_tree_add_7_45_groupi_g4577__4733(csa_tree_add_7_45_groupi_n_759 ,csa_tree_add_7_45_groupi_n_415 ,csa_tree_add_7_45_groupi_n_591);
  xnor csa_tree_add_7_45_groupi_g4578__6161(csa_tree_add_7_45_groupi_n_757 ,csa_tree_add_7_45_groupi_n_411 ,csa_tree_add_7_45_groupi_n_576);
  xnor csa_tree_add_7_45_groupi_g4579__9315(csa_tree_add_7_45_groupi_n_756 ,csa_tree_add_7_45_groupi_n_374 ,csa_tree_add_7_45_groupi_n_578);
  or csa_tree_add_7_45_groupi_g4580__9945(csa_tree_add_7_45_groupi_n_755 ,csa_tree_add_7_45_groupi_n_594 ,csa_tree_add_7_45_groupi_n_709);
  xnor csa_tree_add_7_45_groupi_g4581__2883(csa_tree_add_7_45_groupi_n_753 ,csa_tree_add_7_45_groupi_n_404 ,csa_tree_add_7_45_groupi_n_585);
  xnor csa_tree_add_7_45_groupi_g4582__2346(csa_tree_add_7_45_groupi_n_751 ,csa_tree_add_7_45_groupi_n_405 ,csa_tree_add_7_45_groupi_n_583);
  or csa_tree_add_7_45_groupi_g4583__1666(csa_tree_add_7_45_groupi_n_750 ,csa_tree_add_7_45_groupi_n_633 ,csa_tree_add_7_45_groupi_n_729);
  xnor csa_tree_add_7_45_groupi_g4584__7410(csa_tree_add_7_45_groupi_n_749 ,csa_tree_add_7_45_groupi_n_373 ,csa_tree_add_7_45_groupi_n_586);
  not csa_tree_add_7_45_groupi_g4586(csa_tree_add_7_45_groupi_n_731 ,csa_tree_add_7_45_groupi_n_730);
  and csa_tree_add_7_45_groupi_g4587__6417(csa_tree_add_7_45_groupi_n_729 ,csa_tree_add_7_45_groupi_n_625 ,csa_tree_add_7_45_groupi_n_648);
  or csa_tree_add_7_45_groupi_g4588__5477(csa_tree_add_7_45_groupi_n_728 ,csa_tree_add_7_45_groupi_n_444 ,csa_tree_add_7_45_groupi_n_661);
  or csa_tree_add_7_45_groupi_g4589__2398(csa_tree_add_7_45_groupi_n_727 ,csa_tree_add_7_45_groupi_n_523 ,csa_tree_add_7_45_groupi_n_658);
  or csa_tree_add_7_45_groupi_g4590__5107(csa_tree_add_7_45_groupi_n_726 ,csa_tree_add_7_45_groupi_n_524 ,csa_tree_add_7_45_groupi_n_653);
  or csa_tree_add_7_45_groupi_g4591__6260(csa_tree_add_7_45_groupi_n_725 ,csa_tree_add_7_45_groupi_n_435 ,csa_tree_add_7_45_groupi_n_621);
  nor csa_tree_add_7_45_groupi_g4592__4319(csa_tree_add_7_45_groupi_n_724 ,csa_tree_add_7_45_groupi_n_451 ,csa_tree_add_7_45_groupi_n_657);
  or csa_tree_add_7_45_groupi_g4593__8428(csa_tree_add_7_45_groupi_n_723 ,csa_tree_add_7_45_groupi_n_521 ,csa_tree_add_7_45_groupi_n_647);
  or csa_tree_add_7_45_groupi_g4594__5526(csa_tree_add_7_45_groupi_n_722 ,csa_tree_add_7_45_groupi_n_442 ,csa_tree_add_7_45_groupi_n_643);
  or csa_tree_add_7_45_groupi_g4595__6783(csa_tree_add_7_45_groupi_n_721 ,csa_tree_add_7_45_groupi_n_445 ,csa_tree_add_7_45_groupi_n_660);
  nor csa_tree_add_7_45_groupi_g4596__3680(csa_tree_add_7_45_groupi_n_720 ,csa_tree_add_7_45_groupi_n_409 ,csa_tree_add_7_45_groupi_n_636);
  or csa_tree_add_7_45_groupi_g4597__1617(csa_tree_add_7_45_groupi_n_719 ,csa_tree_add_7_45_groupi_n_449 ,csa_tree_add_7_45_groupi_n_627);
  and csa_tree_add_7_45_groupi_g4598__2802(csa_tree_add_7_45_groupi_n_718 ,csa_tree_add_7_45_groupi_n_631 ,csa_tree_add_7_45_groupi_n_624);
  or csa_tree_add_7_45_groupi_g4599__1705(csa_tree_add_7_45_groupi_n_717 ,csa_tree_add_7_45_groupi_n_452 ,csa_tree_add_7_45_groupi_n_629);
  or csa_tree_add_7_45_groupi_g4600__5122(csa_tree_add_7_45_groupi_n_716 ,csa_tree_add_7_45_groupi_n_410 ,csa_tree_add_7_45_groupi_n_672);
  or csa_tree_add_7_45_groupi_g4601__8246(csa_tree_add_7_45_groupi_n_715 ,csa_tree_add_7_45_groupi_n_450 ,csa_tree_add_7_45_groupi_n_611);
  nor csa_tree_add_7_45_groupi_g4602__7098(csa_tree_add_7_45_groupi_n_714 ,csa_tree_add_7_45_groupi_n_436 ,csa_tree_add_7_45_groupi_n_620);
  and csa_tree_add_7_45_groupi_g4603__6131(csa_tree_add_7_45_groupi_n_713 ,csa_tree_add_7_45_groupi_n_402 ,csa_tree_add_7_45_groupi_n_602);
  nor csa_tree_add_7_45_groupi_g4604__1881(csa_tree_add_7_45_groupi_n_712 ,csa_tree_add_7_45_groupi_n_520 ,csa_tree_add_7_45_groupi_n_600);
  or csa_tree_add_7_45_groupi_g4605__5115(csa_tree_add_7_45_groupi_n_711 ,csa_tree_add_7_45_groupi_n_522 ,csa_tree_add_7_45_groupi_n_592);
  or csa_tree_add_7_45_groupi_g4606__7482(csa_tree_add_7_45_groupi_n_710 ,csa_tree_add_7_45_groupi_n_559 ,csa_tree_add_7_45_groupi_n_615);
  and csa_tree_add_7_45_groupi_g4607__4733(csa_tree_add_7_45_groupi_n_709 ,csa_tree_add_7_45_groupi_n_447 ,csa_tree_add_7_45_groupi_n_659);
  or csa_tree_add_7_45_groupi_g4608__6161(csa_tree_add_7_45_groupi_n_742 ,csa_tree_add_7_45_groupi_n_531 ,csa_tree_add_7_45_groupi_n_613);
  or csa_tree_add_7_45_groupi_g4609__9315(csa_tree_add_7_45_groupi_n_741 ,csa_tree_add_7_45_groupi_n_544 ,csa_tree_add_7_45_groupi_n_635);
  and csa_tree_add_7_45_groupi_g4610__9945(csa_tree_add_7_45_groupi_n_740 ,csa_tree_add_7_45_groupi_n_534 ,csa_tree_add_7_45_groupi_n_668);
  or csa_tree_add_7_45_groupi_g4611__2883(csa_tree_add_7_45_groupi_n_739 ,csa_tree_add_7_45_groupi_n_533 ,csa_tree_add_7_45_groupi_n_669);
  or csa_tree_add_7_45_groupi_g4612__2346(csa_tree_add_7_45_groupi_n_738 ,csa_tree_add_7_45_groupi_n_540 ,csa_tree_add_7_45_groupi_n_630);
  and csa_tree_add_7_45_groupi_g4613__1666(csa_tree_add_7_45_groupi_n_737 ,csa_tree_add_7_45_groupi_n_542 ,csa_tree_add_7_45_groupi_n_601);
  or csa_tree_add_7_45_groupi_g4614__7410(csa_tree_add_7_45_groupi_n_736 ,csa_tree_add_7_45_groupi_n_528 ,csa_tree_add_7_45_groupi_n_650);
  and csa_tree_add_7_45_groupi_g4615__6417(csa_tree_add_7_45_groupi_n_735 ,csa_tree_add_7_45_groupi_n_553 ,csa_tree_add_7_45_groupi_n_663);
  or csa_tree_add_7_45_groupi_g4616__5477(csa_tree_add_7_45_groupi_n_734 ,csa_tree_add_7_45_groupi_n_554 ,csa_tree_add_7_45_groupi_n_670);
  or csa_tree_add_7_45_groupi_g4617__2398(csa_tree_add_7_45_groupi_n_733 ,csa_tree_add_7_45_groupi_n_547 ,csa_tree_add_7_45_groupi_n_645);
  or csa_tree_add_7_45_groupi_g4618__5107(csa_tree_add_7_45_groupi_n_732 ,csa_tree_add_7_45_groupi_n_422 ,csa_tree_add_7_45_groupi_n_599);
  or csa_tree_add_7_45_groupi_g4619__6260(csa_tree_add_7_45_groupi_n_730 ,csa_tree_add_7_45_groupi_n_549 ,csa_tree_add_7_45_groupi_n_641);
  not csa_tree_add_7_45_groupi_g4620(csa_tree_add_7_45_groupi_n_706 ,csa_tree_add_7_45_groupi_n_707);
  nor csa_tree_add_7_45_groupi_g4623__4319(csa_tree_add_7_45_groupi_n_701 ,csa_tree_add_7_45_groupi_n_560 ,csa_tree_add_7_45_groupi_n_616);
  nor csa_tree_add_7_45_groupi_g4624__8428(csa_tree_add_7_45_groupi_n_700 ,csa_tree_add_7_45_groupi_n_446 ,csa_tree_add_7_45_groupi_n_604);
  or csa_tree_add_7_45_groupi_g4625__5526(csa_tree_add_7_45_groupi_n_699 ,csa_tree_add_7_45_groupi_n_623 ,csa_tree_add_7_45_groupi_n_640);
  xnor csa_tree_add_7_45_groupi_g4626__6783(csa_tree_add_7_45_groupi_n_698 ,csa_tree_add_7_45_groupi_n_469 ,csa_tree_add_7_45_groupi_n_490);
  xnor csa_tree_add_7_45_groupi_g4627__3680(csa_tree_add_7_45_groupi_n_697 ,csa_tree_add_7_45_groupi_n_522 ,csa_tree_add_7_45_groupi_n_515);
  xnor csa_tree_add_7_45_groupi_g4628__1617(csa_tree_add_7_45_groupi_n_696 ,csa_tree_add_7_45_groupi_n_492 ,csa_tree_add_7_45_groupi_n_488);
  xnor csa_tree_add_7_45_groupi_g4629__2802(csa_tree_add_7_45_groupi_n_695 ,csa_tree_add_7_45_groupi_n_511 ,csa_tree_add_7_45_groupi_n_574);
  xnor csa_tree_add_7_45_groupi_g4630__1705(csa_tree_add_7_45_groupi_n_694 ,csa_tree_add_7_45_groupi_n_462 ,csa_tree_add_7_45_groupi_n_513);
  xnor csa_tree_add_7_45_groupi_g4631__5122(csa_tree_add_7_45_groupi_n_693 ,csa_tree_add_7_45_groupi_n_502 ,csa_tree_add_7_45_groupi_n_569);
  xnor csa_tree_add_7_45_groupi_g4632__8246(csa_tree_add_7_45_groupi_n_692 ,csa_tree_add_7_45_groupi_n_521 ,csa_tree_add_7_45_groupi_n_300);
  xnor csa_tree_add_7_45_groupi_g4633__7098(csa_tree_add_7_45_groupi_n_691 ,csa_tree_add_7_45_groupi_n_294 ,csa_tree_add_7_45_groupi_n_558);
  xnor csa_tree_add_7_45_groupi_g4634__6131(csa_tree_add_7_45_groupi_n_690 ,csa_tree_add_7_45_groupi_n_484 ,csa_tree_add_7_45_groupi_n_461);
  xnor csa_tree_add_7_45_groupi_g4635__1881(csa_tree_add_7_45_groupi_n_689 ,csa_tree_add_7_45_groupi_n_486 ,csa_tree_add_7_45_groupi_n_498);
  xnor csa_tree_add_7_45_groupi_g4636__5115(csa_tree_add_7_45_groupi_n_688 ,csa_tree_add_7_45_groupi_n_477 ,in3[0]);
  xnor csa_tree_add_7_45_groupi_g4637__7482(csa_tree_add_7_45_groupi_n_687 ,csa_tree_add_7_45_groupi_n_496 ,csa_tree_add_7_45_groupi_n_564);
  xnor csa_tree_add_7_45_groupi_g4638__4733(csa_tree_add_7_45_groupi_n_686 ,csa_tree_add_7_45_groupi_n_476 ,csa_tree_add_7_45_groupi_n_507);
  xor csa_tree_add_7_45_groupi_g4639__6161(csa_tree_add_7_45_groupi_n_685 ,csa_tree_add_7_45_groupi_n_509 ,csa_tree_add_7_45_groupi_n_442);
  xor csa_tree_add_7_45_groupi_g4640__9315(csa_tree_add_7_45_groupi_n_684 ,csa_tree_add_7_45_groupi_n_479 ,csa_tree_add_7_45_groupi_n_450);
  xnor csa_tree_add_7_45_groupi_g4641__9945(csa_tree_add_7_45_groupi_n_683 ,csa_tree_add_7_45_groupi_n_402 ,csa_tree_add_7_45_groupi_n_473);
  xor csa_tree_add_7_45_groupi_g4642__2883(csa_tree_add_7_45_groupi_n_682 ,csa_tree_add_7_45_groupi_n_512 ,csa_tree_add_7_45_groupi_n_444);
  xor csa_tree_add_7_45_groupi_g4643__2346(csa_tree_add_7_45_groupi_n_681 ,csa_tree_add_7_45_groupi_n_464 ,csa_tree_add_7_45_groupi_n_452);
  xnor csa_tree_add_7_45_groupi_g4644__1666(csa_tree_add_7_45_groupi_n_680 ,csa_tree_add_7_45_groupi_n_567 ,csa_tree_add_7_45_groupi_n_570);
  xnor csa_tree_add_7_45_groupi_g4645__7410(csa_tree_add_7_45_groupi_n_679 ,csa_tree_add_7_45_groupi_n_561 ,csa_tree_add_7_45_groupi_n_516);
  xnor csa_tree_add_7_45_groupi_g4646__6417(csa_tree_add_7_45_groupi_n_678 ,csa_tree_add_7_45_groupi_n_480 ,csa_tree_add_7_45_groupi_n_446);
  xnor csa_tree_add_7_45_groupi_g4647__5477(csa_tree_add_7_45_groupi_n_677 ,csa_tree_add_7_45_groupi_n_508 ,csa_tree_add_7_45_groupi_n_55);
  xnor csa_tree_add_7_45_groupi_g4648__2398(csa_tree_add_7_45_groupi_n_676 ,csa_tree_add_7_45_groupi_n_493 ,csa_tree_add_7_45_groupi_n_161);
  xnor csa_tree_add_7_45_groupi_g4649__5107(csa_tree_add_7_45_groupi_n_675 ,csa_tree_add_7_45_groupi_n_478 ,csa_tree_add_7_45_groupi_n_566);
  xnor csa_tree_add_7_45_groupi_g4650__6260(csa_tree_add_7_45_groupi_n_674 ,csa_tree_add_7_45_groupi_n_474 ,csa_tree_add_7_45_groupi_n_565);
  or csa_tree_add_7_45_groupi_g4651__4319(csa_tree_add_7_45_groupi_n_708 ,csa_tree_add_7_45_groupi_n_546 ,csa_tree_add_7_45_groupi_n_598);
  xnor csa_tree_add_7_45_groupi_g4652__8428(csa_tree_add_7_45_groupi_n_707 ,csa_tree_add_7_45_groupi_n_408 ,csa_tree_add_7_45_groupi_n_527);
  xnor csa_tree_add_7_45_groupi_g4653__5526(csa_tree_add_7_45_groupi_n_705 ,csa_tree_add_7_45_groupi_n_406 ,csa_tree_add_7_45_groupi_n_457);
  xnor csa_tree_add_7_45_groupi_g4654__6783(csa_tree_add_7_45_groupi_n_704 ,csa_tree_add_7_45_groupi_n_575 ,csa_tree_add_7_45_groupi_n_525);
  xnor csa_tree_add_7_45_groupi_g4655__3680(csa_tree_add_7_45_groupi_n_703 ,csa_tree_add_7_45_groupi_n_401 ,csa_tree_add_7_45_groupi_n_526);
  xnor csa_tree_add_7_45_groupi_g4656__1617(csa_tree_add_7_45_groupi_n_702 ,csa_tree_add_7_45_groupi_n_170 ,csa_tree_add_7_45_groupi_n_458);
  or csa_tree_add_7_45_groupi_g4657__2802(csa_tree_add_7_45_groupi_n_673 ,csa_tree_add_7_45_groupi_n_108 ,csa_tree_add_7_45_groupi_n_477);
  and csa_tree_add_7_45_groupi_g4658__1705(csa_tree_add_7_45_groupi_n_672 ,csa_tree_add_7_45_groupi_n_108 ,csa_tree_add_7_45_groupi_n_477);
  or csa_tree_add_7_45_groupi_g4659__5122(csa_tree_add_7_45_groupi_n_671 ,csa_tree_add_7_45_groupi_n_513 ,csa_tree_add_7_45_groupi_n_463);
  and csa_tree_add_7_45_groupi_g4660__8246(csa_tree_add_7_45_groupi_n_670 ,csa_tree_add_7_45_groupi_n_403 ,csa_tree_add_7_45_groupi_n_529);
  and csa_tree_add_7_45_groupi_g4661__7098(csa_tree_add_7_45_groupi_n_669 ,csa_tree_add_7_45_groupi_n_443 ,csa_tree_add_7_45_groupi_n_532);
  or csa_tree_add_7_45_groupi_g4662__6131(csa_tree_add_7_45_groupi_n_668 ,csa_tree_add_7_45_groupi_n_417 ,csa_tree_add_7_45_groupi_n_555);
  or csa_tree_add_7_45_groupi_g4663__1881(csa_tree_add_7_45_groupi_n_667 ,csa_tree_add_7_45_groupi_n_300 ,csa_tree_add_7_45_groupi_n_494);
  or csa_tree_add_7_45_groupi_g4664__5115(csa_tree_add_7_45_groupi_n_666 ,csa_tree_add_7_45_groupi_n_566 ,csa_tree_add_7_45_groupi_n_478);
  and csa_tree_add_7_45_groupi_g4665__7482(csa_tree_add_7_45_groupi_n_665 ,csa_tree_add_7_45_groupi_n_566 ,csa_tree_add_7_45_groupi_n_478);
  or csa_tree_add_7_45_groupi_g4666__4733(csa_tree_add_7_45_groupi_n_664 ,csa_tree_add_7_45_groupi_n_512 ,csa_tree_add_7_45_groupi_n_503);
  or csa_tree_add_7_45_groupi_g4667__6161(csa_tree_add_7_45_groupi_n_663 ,csa_tree_add_7_45_groupi_n_412 ,csa_tree_add_7_45_groupi_n_552);
  or csa_tree_add_7_45_groupi_g4668__9315(csa_tree_add_7_45_groupi_n_662 ,csa_tree_add_7_45_groupi_n_568 ,csa_tree_add_7_45_groupi_n_502);
  and csa_tree_add_7_45_groupi_g4669__9945(csa_tree_add_7_45_groupi_n_661 ,csa_tree_add_7_45_groupi_n_512 ,csa_tree_add_7_45_groupi_n_503);
  and csa_tree_add_7_45_groupi_g4670__2883(csa_tree_add_7_45_groupi_n_660 ,csa_tree_add_7_45_groupi_n_296 ,csa_tree_add_7_45_groupi_n_467);
  or csa_tree_add_7_45_groupi_g4671__2346(csa_tree_add_7_45_groupi_n_659 ,csa_tree_add_7_45_groupi_n_391 ,csa_tree_add_7_45_groupi_n_505);
  nor csa_tree_add_7_45_groupi_g4672__1666(csa_tree_add_7_45_groupi_n_658 ,csa_tree_add_7_45_groupi_n_569 ,csa_tree_add_7_45_groupi_n_501);
  nor csa_tree_add_7_45_groupi_g4673__7410(csa_tree_add_7_45_groupi_n_657 ,csa_tree_add_7_45_groupi_n_233 ,csa_tree_add_7_45_groupi_n_562);
  nor csa_tree_add_7_45_groupi_g4674__6417(csa_tree_add_7_45_groupi_n_656 ,csa_tree_add_7_45_groupi_n_563 ,csa_tree_add_7_45_groupi_n_496);
  or csa_tree_add_7_45_groupi_g4675__5477(csa_tree_add_7_45_groupi_n_655 ,csa_tree_add_7_45_groupi_n_293 ,csa_tree_add_7_45_groupi_n_49);
  or csa_tree_add_7_45_groupi_g4676__2398(csa_tree_add_7_45_groupi_n_654 ,csa_tree_add_7_45_groupi_n_573 ,csa_tree_add_7_45_groupi_n_511);
  nor csa_tree_add_7_45_groupi_g4677__5107(csa_tree_add_7_45_groupi_n_653 ,csa_tree_add_7_45_groupi_n_574 ,csa_tree_add_7_45_groupi_n_510);
  or csa_tree_add_7_45_groupi_g4678__6260(csa_tree_add_7_45_groupi_n_652 ,csa_tree_add_7_45_groupi_n_561 ,csa_tree_add_7_45_groupi_n_517);
  or csa_tree_add_7_45_groupi_g4679__4319(csa_tree_add_7_45_groupi_n_651 ,csa_tree_add_7_45_groupi_n_507 ,csa_tree_add_7_45_groupi_n_475);
  and csa_tree_add_7_45_groupi_g4680__8428(csa_tree_add_7_45_groupi_n_650 ,csa_tree_add_7_45_groupi_n_415 ,csa_tree_add_7_45_groupi_n_538);
  and csa_tree_add_7_45_groupi_g4681__5526(csa_tree_add_7_45_groupi_n_649 ,csa_tree_add_7_45_groupi_n_38 ,csa_tree_add_7_45_groupi_n_562);
  or csa_tree_add_7_45_groupi_g4682__6783(csa_tree_add_7_45_groupi_n_648 ,csa_tree_add_7_45_groupi_n_488 ,csa_tree_add_7_45_groupi_n_491);
  and csa_tree_add_7_45_groupi_g4683__3680(csa_tree_add_7_45_groupi_n_647 ,csa_tree_add_7_45_groupi_n_300 ,csa_tree_add_7_45_groupi_n_494);
  or csa_tree_add_7_45_groupi_g4684__1617(csa_tree_add_7_45_groupi_n_646 ,csa_tree_add_7_45_groupi_n_509 ,csa_tree_add_7_45_groupi_n_499);
  and csa_tree_add_7_45_groupi_g4685__2802(csa_tree_add_7_45_groupi_n_645 ,csa_tree_add_7_45_groupi_n_413 ,csa_tree_add_7_45_groupi_n_550);
  nor csa_tree_add_7_45_groupi_g4686__1705(csa_tree_add_7_45_groupi_n_644 ,csa_tree_add_7_45_groupi_n_294 ,csa_tree_add_7_45_groupi_n_58);
  and csa_tree_add_7_45_groupi_g4687__5122(csa_tree_add_7_45_groupi_n_643 ,csa_tree_add_7_45_groupi_n_509 ,csa_tree_add_7_45_groupi_n_499);
  or csa_tree_add_7_45_groupi_g4688__8246(csa_tree_add_7_45_groupi_n_642 ,csa_tree_add_7_45_groupi_n_497 ,csa_tree_add_7_45_groupi_n_486);
  nor csa_tree_add_7_45_groupi_g4689__7098(csa_tree_add_7_45_groupi_n_641 ,csa_tree_add_7_45_groupi_n_448 ,csa_tree_add_7_45_groupi_n_537);
  nor csa_tree_add_7_45_groupi_g4690__6131(csa_tree_add_7_45_groupi_n_640 ,csa_tree_add_7_45_groupi_n_498 ,csa_tree_add_7_45_groupi_n_485);
  or csa_tree_add_7_45_groupi_g4691__1881(csa_tree_add_7_45_groupi_n_639 ,csa_tree_add_7_45_groupi_n_500 ,csa_tree_add_7_45_groupi_n_479);
  and csa_tree_add_7_45_groupi_g4692__5115(csa_tree_add_7_45_groupi_n_638 ,csa_tree_add_7_45_groupi_n_567 ,csa_tree_add_7_45_groupi_n_570);
  nor csa_tree_add_7_45_groupi_g4693__7482(csa_tree_add_7_45_groupi_n_637 ,csa_tree_add_7_45_groupi_n_460 ,csa_tree_add_7_45_groupi_n_484);
  nor csa_tree_add_7_45_groupi_g4694__4733(csa_tree_add_7_45_groupi_n_636 ,csa_tree_add_7_45_groupi_n_567 ,csa_tree_add_7_45_groupi_n_570);
  nor csa_tree_add_7_45_groupi_g4695__6161(csa_tree_add_7_45_groupi_n_635 ,csa_tree_add_7_45_groupi_n_441 ,csa_tree_add_7_45_groupi_n_548);
  or csa_tree_add_7_45_groupi_g4696__9315(csa_tree_add_7_45_groupi_n_634 ,csa_tree_add_7_45_groupi_n_292 ,csa_tree_add_7_45_groupi_n_482);
  nor csa_tree_add_7_45_groupi_g4697__9945(csa_tree_add_7_45_groupi_n_633 ,csa_tree_add_7_45_groupi_n_487 ,csa_tree_add_7_45_groupi_n_492);
  and csa_tree_add_7_45_groupi_g4698__2883(csa_tree_add_7_45_groupi_n_632 ,csa_tree_add_7_45_groupi_n_53 ,csa_tree_add_7_45_groupi_n_493);
  or csa_tree_add_7_45_groupi_g4699__2346(csa_tree_add_7_45_groupi_n_631 ,csa_tree_add_7_45_groupi_n_161 ,csa_tree_add_7_45_groupi_n_493);
  and csa_tree_add_7_45_groupi_g4700__1666(csa_tree_add_7_45_groupi_n_630 ,csa_tree_add_7_45_groupi_n_411 ,csa_tree_add_7_45_groupi_n_551);
  and csa_tree_add_7_45_groupi_g4701__7410(csa_tree_add_7_45_groupi_n_629 ,csa_tree_add_7_45_groupi_n_464 ,csa_tree_add_7_45_groupi_n_481);
  and csa_tree_add_7_45_groupi_g4702__6417(csa_tree_add_7_45_groupi_n_628 ,csa_tree_add_7_45_groupi_n_565 ,csa_tree_add_7_45_groupi_n_474);
  and csa_tree_add_7_45_groupi_g4703__5477(csa_tree_add_7_45_groupi_n_627 ,csa_tree_add_7_45_groupi_n_292 ,csa_tree_add_7_45_groupi_n_482);
  nor csa_tree_add_7_45_groupi_g4704__2398(csa_tree_add_7_45_groupi_n_626 ,csa_tree_add_7_45_groupi_n_506 ,csa_tree_add_7_45_groupi_n_476);
  not csa_tree_add_7_45_groupi_g4705(csa_tree_add_7_45_groupi_n_620 ,csa_tree_add_7_45_groupi_n_621);
  not csa_tree_add_7_45_groupi_g4706(csa_tree_add_7_45_groupi_n_618 ,csa_tree_add_7_45_groupi_n_617);
  not csa_tree_add_7_45_groupi_g4707(csa_tree_add_7_45_groupi_n_615 ,csa_tree_add_7_45_groupi_n_616);
  or csa_tree_add_7_45_groupi_g4708__5107(csa_tree_add_7_45_groupi_n_614 ,csa_tree_add_7_45_groupi_n_474 ,csa_tree_add_7_45_groupi_n_565);
  and csa_tree_add_7_45_groupi_g4709__6260(csa_tree_add_7_45_groupi_n_613 ,csa_tree_add_7_45_groupi_n_405 ,csa_tree_add_7_45_groupi_n_530);
  or csa_tree_add_7_45_groupi_g4710__4319(csa_tree_add_7_45_groupi_n_612 ,csa_tree_add_7_45_groupi_n_564 ,csa_tree_add_7_45_groupi_n_495);
  and csa_tree_add_7_45_groupi_g4711__8428(csa_tree_add_7_45_groupi_n_611 ,csa_tree_add_7_45_groupi_n_500 ,csa_tree_add_7_45_groupi_n_479);
  or csa_tree_add_7_45_groupi_g4712__5526(csa_tree_add_7_45_groupi_n_610 ,csa_tree_add_7_45_groupi_n_296 ,csa_tree_add_7_45_groupi_n_467);
  or csa_tree_add_7_45_groupi_g4713__6783(csa_tree_add_7_45_groupi_n_609 ,csa_tree_add_7_45_groupi_n_461 ,csa_tree_add_7_45_groupi_n_483);
  and csa_tree_add_7_45_groupi_g4714__3680(csa_tree_add_7_45_groupi_n_608 ,csa_tree_add_7_45_groupi_n_561 ,csa_tree_add_7_45_groupi_n_517);
  nor csa_tree_add_7_45_groupi_g4715__1617(csa_tree_add_7_45_groupi_n_607 ,csa_tree_add_7_45_groupi_n_473 ,csa_tree_add_7_45_groupi_n_471);
  and csa_tree_add_7_45_groupi_g4716__2802(csa_tree_add_7_45_groupi_n_606 ,csa_tree_add_7_45_groupi_n_55 ,csa_tree_add_7_45_groupi_n_508);
  or csa_tree_add_7_45_groupi_g4717__1705(csa_tree_add_7_45_groupi_n_605 ,csa_tree_add_7_45_groupi_n_489 ,csa_tree_add_7_45_groupi_n_469);
  and csa_tree_add_7_45_groupi_g4718__5122(csa_tree_add_7_45_groupi_n_604 ,csa_tree_add_7_45_groupi_n_480 ,csa_tree_add_7_45_groupi_n_572);
  nor csa_tree_add_7_45_groupi_g4719__8246(csa_tree_add_7_45_groupi_n_603 ,csa_tree_add_7_45_groupi_n_490 ,csa_tree_add_7_45_groupi_n_468);
  or csa_tree_add_7_45_groupi_g4720__7098(csa_tree_add_7_45_groupi_n_602 ,csa_tree_add_7_45_groupi_n_472 ,csa_tree_add_7_45_groupi_n_470);
  or csa_tree_add_7_45_groupi_g4721__6131(csa_tree_add_7_45_groupi_n_601 ,csa_tree_add_7_45_groupi_n_400 ,csa_tree_add_7_45_groupi_n_541);
  nor csa_tree_add_7_45_groupi_g4722__1881(csa_tree_add_7_45_groupi_n_600 ,csa_tree_add_7_45_groupi_n_234 ,csa_tree_add_7_45_groupi_n_508);
  and csa_tree_add_7_45_groupi_g4723__5115(csa_tree_add_7_45_groupi_n_599 ,csa_tree_add_7_45_groupi_n_425 ,csa_tree_add_7_45_groupi_n_575);
  and csa_tree_add_7_45_groupi_g4724__7482(csa_tree_add_7_45_groupi_n_598 ,csa_tree_add_7_45_groupi_n_404 ,csa_tree_add_7_45_groupi_n_545);
  nor csa_tree_add_7_45_groupi_g4725__4733(csa_tree_add_7_45_groupi_n_597 ,csa_tree_add_7_45_groupi_n_480 ,csa_tree_add_7_45_groupi_n_572);
  or csa_tree_add_7_45_groupi_g4726__6161(csa_tree_add_7_45_groupi_n_596 ,csa_tree_add_7_45_groupi_n_514 ,csa_tree_add_7_45_groupi_n_466);
  or csa_tree_add_7_45_groupi_g4727__9315(csa_tree_add_7_45_groupi_n_595 ,csa_tree_add_7_45_groupi_n_464 ,csa_tree_add_7_45_groupi_n_481);
  and csa_tree_add_7_45_groupi_g4728__9945(csa_tree_add_7_45_groupi_n_594 ,csa_tree_add_7_45_groupi_n_391 ,csa_tree_add_7_45_groupi_n_505);
  and csa_tree_add_7_45_groupi_g4729__2883(csa_tree_add_7_45_groupi_n_593 ,csa_tree_add_7_45_groupi_n_513 ,csa_tree_add_7_45_groupi_n_463);
  nor csa_tree_add_7_45_groupi_g4730__2346(csa_tree_add_7_45_groupi_n_592 ,csa_tree_add_7_45_groupi_n_515 ,csa_tree_add_7_45_groupi_n_465);
  xnor csa_tree_add_7_45_groupi_g4731__1666(csa_tree_add_7_45_groupi_n_591 ,csa_tree_add_7_45_groupi_n_395 ,csa_tree_add_7_45_groupi_n_430);
  xor csa_tree_add_7_45_groupi_g4732__7410(csa_tree_add_7_45_groupi_n_590 ,csa_tree_add_7_45_groupi_n_441 ,in2[13]);
  xnor csa_tree_add_7_45_groupi_g4733__6417(csa_tree_add_7_45_groupi_n_589 ,csa_tree_add_7_45_groupi_n_171 ,csa_tree_add_7_45_groupi_n_434);
  xnor csa_tree_add_7_45_groupi_g4734__5477(csa_tree_add_7_45_groupi_n_588 ,csa_tree_add_7_45_groupi_n_449 ,csa_tree_add_7_45_groupi_n_292);
  xnor csa_tree_add_7_45_groupi_g4735__2398(csa_tree_add_7_45_groupi_n_587 ,csa_tree_add_7_45_groupi_n_391 ,csa_tree_add_7_45_groupi_n_447);
  xnor csa_tree_add_7_45_groupi_g4736__5107(csa_tree_add_7_45_groupi_n_586 ,csa_tree_add_7_45_groupi_n_413 ,csa_tree_add_7_45_groupi_n_390);
  xnor csa_tree_add_7_45_groupi_g4737__6260(csa_tree_add_7_45_groupi_n_585 ,csa_tree_add_7_45_groupi_n_165 ,csa_tree_add_7_45_groupi_n_439);
  xor csa_tree_add_7_45_groupi_g4738__4319(csa_tree_add_7_45_groupi_n_584 ,csa_tree_add_7_45_groupi_n_445 ,csa_tree_add_7_45_groupi_n_296);
  xnor csa_tree_add_7_45_groupi_g4739__8428(csa_tree_add_7_45_groupi_n_583 ,csa_tree_add_7_45_groupi_n_399 ,csa_tree_add_7_45_groupi_n_393);
  xnor csa_tree_add_7_45_groupi_g4740__5526(csa_tree_add_7_45_groupi_n_582 ,csa_tree_add_7_45_groupi_n_163 ,csa_tree_add_7_45_groupi_n_432);
  xnor csa_tree_add_7_45_groupi_g4741__6783(csa_tree_add_7_45_groupi_n_581 ,csa_tree_add_7_45_groupi_n_440 ,csa_tree_add_7_45_groupi_n_427);
  xnor csa_tree_add_7_45_groupi_g4742__3680(csa_tree_add_7_45_groupi_n_580 ,csa_tree_add_7_45_groupi_n_387 ,csa_tree_add_7_45_groupi_n_443);
  xnor csa_tree_add_7_45_groupi_g4743__1617(csa_tree_add_7_45_groupi_n_579 ,csa_tree_add_7_45_groupi_n_397 ,csa_tree_add_7_45_groupi_n_385);
  xnor csa_tree_add_7_45_groupi_g4744__2802(csa_tree_add_7_45_groupi_n_578 ,csa_tree_add_7_45_groupi_n_448 ,csa_tree_add_7_45_groupi_n_428);
  xor csa_tree_add_7_45_groupi_g4745__1705(csa_tree_add_7_45_groupi_n_577 ,csa_tree_add_7_45_groupi_n_451 ,csa_tree_add_7_45_groupi_n_38);
  xnor csa_tree_add_7_45_groupi_g4746__5122(csa_tree_add_7_45_groupi_n_576 ,csa_tree_add_7_45_groupi_n_433 ,csa_tree_add_7_45_groupi_n_388);
  or csa_tree_add_7_45_groupi_g4747__8246(csa_tree_add_7_45_groupi_n_625 ,csa_tree_add_7_45_groupi_n_349 ,csa_tree_add_7_45_groupi_n_557);
  or csa_tree_add_7_45_groupi_g4748__7098(csa_tree_add_7_45_groupi_n_624 ,csa_tree_add_7_45_groupi_n_423 ,csa_tree_add_7_45_groupi_n_556);
  and csa_tree_add_7_45_groupi_g4749__6131(csa_tree_add_7_45_groupi_n_623 ,csa_tree_add_7_45_groupi_n_357 ,csa_tree_add_7_45_groupi_n_535);
  or csa_tree_add_7_45_groupi_g4750__1881(csa_tree_add_7_45_groupi_n_622 ,csa_tree_add_7_45_groupi_n_420 ,csa_tree_add_7_45_groupi_n_536);
  xnor csa_tree_add_7_45_groupi_g4751__5115(csa_tree_add_7_45_groupi_n_621 ,csa_tree_add_7_45_groupi_n_307 ,csa_tree_add_7_45_groupi_n_376);
  or csa_tree_add_7_45_groupi_g4752__7482(csa_tree_add_7_45_groupi_n_619 ,csa_tree_add_7_45_groupi_n_543 ,csa_tree_add_7_45_groupi_n_558);
  or csa_tree_add_7_45_groupi_g4753__4733(csa_tree_add_7_45_groupi_n_617 ,csa_tree_add_7_45_groupi_n_382 ,csa_tree_add_7_45_groupi_n_539);
  xnor csa_tree_add_7_45_groupi_g4754__6161(csa_tree_add_7_45_groupi_n_616 ,csa_tree_add_7_45_groupi_n_407 ,csa_tree_add_7_45_groupi_n_377);
  not csa_tree_add_7_45_groupi_g4756(csa_tree_add_7_45_groupi_n_573 ,csa_tree_add_7_45_groupi_n_574);
  not csa_tree_add_7_45_groupi_g4757(csa_tree_add_7_45_groupi_n_572 ,csa_tree_add_7_45_groupi_n_571);
  not csa_tree_add_7_45_groupi_g4758(csa_tree_add_7_45_groupi_n_568 ,csa_tree_add_7_45_groupi_n_569);
  not csa_tree_add_7_45_groupi_g4759(csa_tree_add_7_45_groupi_n_563 ,csa_tree_add_7_45_groupi_n_564);
  not csa_tree_add_7_45_groupi_g4760(csa_tree_add_7_45_groupi_n_559 ,csa_tree_add_7_45_groupi_n_560);
  and csa_tree_add_7_45_groupi_g4762__9315(csa_tree_add_7_45_groupi_n_557 ,csa_tree_add_7_45_groupi_n_346 ,csa_tree_add_7_45_groupi_n_407);
  and csa_tree_add_7_45_groupi_g4763__9945(csa_tree_add_7_45_groupi_n_556 ,csa_tree_add_7_45_groupi_n_401 ,csa_tree_add_7_45_groupi_n_379);
  nor csa_tree_add_7_45_groupi_g4764__2883(csa_tree_add_7_45_groupi_n_555 ,csa_tree_add_7_45_groupi_n_162 ,csa_tree_add_7_45_groupi_n_432);
  and csa_tree_add_7_45_groupi_g4765__2346(csa_tree_add_7_45_groupi_n_554 ,csa_tree_add_7_45_groupi_n_440 ,csa_tree_add_7_45_groupi_n_427);
  or csa_tree_add_7_45_groupi_g4766__1666(csa_tree_add_7_45_groupi_n_553 ,csa_tree_add_7_45_groupi_n_171 ,csa_tree_add_7_45_groupi_n_434);
  and csa_tree_add_7_45_groupi_g4767__7410(csa_tree_add_7_45_groupi_n_552 ,csa_tree_add_7_45_groupi_n_171 ,csa_tree_add_7_45_groupi_n_434);
  or csa_tree_add_7_45_groupi_g4768__6417(csa_tree_add_7_45_groupi_n_551 ,csa_tree_add_7_45_groupi_n_433 ,csa_tree_add_7_45_groupi_n_388);
  or csa_tree_add_7_45_groupi_g4769__5477(csa_tree_add_7_45_groupi_n_550 ,csa_tree_add_7_45_groupi_n_373 ,csa_tree_add_7_45_groupi_n_389);
  nor csa_tree_add_7_45_groupi_g4770__2398(csa_tree_add_7_45_groupi_n_549 ,csa_tree_add_7_45_groupi_n_375 ,csa_tree_add_7_45_groupi_n_428);
  nor csa_tree_add_7_45_groupi_g4771__5107(csa_tree_add_7_45_groupi_n_548 ,in2[13] ,csa_tree_add_7_45_groupi_n_437);
  nor csa_tree_add_7_45_groupi_g4772__6260(csa_tree_add_7_45_groupi_n_547 ,csa_tree_add_7_45_groupi_n_372 ,csa_tree_add_7_45_groupi_n_390);
  nor csa_tree_add_7_45_groupi_g4773__4319(csa_tree_add_7_45_groupi_n_546 ,csa_tree_add_7_45_groupi_n_165 ,csa_tree_add_7_45_groupi_n_438);
  or csa_tree_add_7_45_groupi_g4774__8428(csa_tree_add_7_45_groupi_n_545 ,csa_tree_add_7_45_groupi_n_164 ,csa_tree_add_7_45_groupi_n_439);
  and csa_tree_add_7_45_groupi_g4775__5526(csa_tree_add_7_45_groupi_n_544 ,in2[13] ,csa_tree_add_7_45_groupi_n_437);
  and csa_tree_add_7_45_groupi_g4776__6783(csa_tree_add_7_45_groupi_n_543 ,csa_tree_add_7_45_groupi_n_453 ,csa_tree_add_7_45_groupi_n_456);
  or csa_tree_add_7_45_groupi_g4777__3680(csa_tree_add_7_45_groupi_n_542 ,csa_tree_add_7_45_groupi_n_396 ,csa_tree_add_7_45_groupi_n_384);
  nor csa_tree_add_7_45_groupi_g4778__1617(csa_tree_add_7_45_groupi_n_541 ,csa_tree_add_7_45_groupi_n_397 ,csa_tree_add_7_45_groupi_n_385);
  and csa_tree_add_7_45_groupi_g4779__2802(csa_tree_add_7_45_groupi_n_540 ,csa_tree_add_7_45_groupi_n_433 ,csa_tree_add_7_45_groupi_n_388);
  and csa_tree_add_7_45_groupi_g4780__1705(csa_tree_add_7_45_groupi_n_539 ,csa_tree_add_7_45_groupi_n_406 ,csa_tree_add_7_45_groupi_n_381);
  or csa_tree_add_7_45_groupi_g4781__5122(csa_tree_add_7_45_groupi_n_538 ,csa_tree_add_7_45_groupi_n_395 ,csa_tree_add_7_45_groupi_n_429);
  and csa_tree_add_7_45_groupi_g4782__8246(csa_tree_add_7_45_groupi_n_537 ,csa_tree_add_7_45_groupi_n_375 ,csa_tree_add_7_45_groupi_n_428);
  and csa_tree_add_7_45_groupi_g4783__7098(csa_tree_add_7_45_groupi_n_536 ,csa_tree_add_7_45_groupi_n_408 ,csa_tree_add_7_45_groupi_n_424);
  or csa_tree_add_7_45_groupi_g4784__6131(csa_tree_add_7_45_groupi_n_535 ,csa_tree_add_7_45_groupi_n_356 ,csa_tree_add_7_45_groupi_n_414);
  or csa_tree_add_7_45_groupi_g4785__1881(csa_tree_add_7_45_groupi_n_534 ,csa_tree_add_7_45_groupi_n_163 ,csa_tree_add_7_45_groupi_n_431);
  nor csa_tree_add_7_45_groupi_g4786__5115(csa_tree_add_7_45_groupi_n_533 ,csa_tree_add_7_45_groupi_n_37 ,csa_tree_add_7_45_groupi_n_387);
  or csa_tree_add_7_45_groupi_g4787__7482(csa_tree_add_7_45_groupi_n_532 ,csa_tree_add_7_45_groupi_n_160 ,csa_tree_add_7_45_groupi_n_386);
  nor csa_tree_add_7_45_groupi_g4788__4733(csa_tree_add_7_45_groupi_n_531 ,csa_tree_add_7_45_groupi_n_398 ,csa_tree_add_7_45_groupi_n_393);
  or csa_tree_add_7_45_groupi_g4789__6161(csa_tree_add_7_45_groupi_n_530 ,csa_tree_add_7_45_groupi_n_399 ,csa_tree_add_7_45_groupi_n_392);
  or csa_tree_add_7_45_groupi_g4790__9315(csa_tree_add_7_45_groupi_n_529 ,csa_tree_add_7_45_groupi_n_440 ,csa_tree_add_7_45_groupi_n_427);
  nor csa_tree_add_7_45_groupi_g4791__9945(csa_tree_add_7_45_groupi_n_528 ,csa_tree_add_7_45_groupi_n_394 ,csa_tree_add_7_45_groupi_n_430);
  xnor csa_tree_add_7_45_groupi_g4792__2883(csa_tree_add_7_45_groupi_n_527 ,csa_tree_add_7_45_groupi_n_291 ,in1[0]);
  xnor csa_tree_add_7_45_groupi_g4793__2346(csa_tree_add_7_45_groupi_n_526 ,csa_tree_add_7_45_groupi_n_303 ,in4[0]);
  xnor csa_tree_add_7_45_groupi_g4794__1666(csa_tree_add_7_45_groupi_n_525 ,csa_tree_add_7_45_groupi_n_167 ,csa_tree_add_7_45_groupi_n_299);
  or csa_tree_add_7_45_groupi_g4795__7410(csa_tree_add_7_45_groupi_n_575 ,csa_tree_add_7_45_groupi_n_347 ,csa_tree_add_7_45_groupi_n_383);
  xnor csa_tree_add_7_45_groupi_g4796__6417(csa_tree_add_7_45_groupi_n_574 ,csa_tree_add_7_45_groupi_n_258 ,in2[5]);
  or csa_tree_add_7_45_groupi_g4797__5477(csa_tree_add_7_45_groupi_n_571 ,csa_tree_add_7_45_groupi_n_418 ,csa_tree_add_7_45_groupi_n_57);
  xnor csa_tree_add_7_45_groupi_g4798__2398(csa_tree_add_7_45_groupi_n_570 ,csa_tree_add_7_45_groupi_n_278 ,in1[3]);
  xnor csa_tree_add_7_45_groupi_g4799__5107(csa_tree_add_7_45_groupi_n_569 ,csa_tree_add_7_45_groupi_n_253 ,in4[5]);
  xnor csa_tree_add_7_45_groupi_g4800__6260(csa_tree_add_7_45_groupi_n_567 ,csa_tree_add_7_45_groupi_n_269 ,in4[1]);
  and csa_tree_add_7_45_groupi_g4801__4319(csa_tree_add_7_45_groupi_n_566 ,csa_tree_add_7_45_groupi_n_137 ,csa_tree_add_7_45_groupi_n_419);
  xnor csa_tree_add_7_45_groupi_g4802__8428(csa_tree_add_7_45_groupi_n_565 ,csa_tree_add_7_45_groupi_n_262 ,in4[7]);
  xnor csa_tree_add_7_45_groupi_g4803__5526(csa_tree_add_7_45_groupi_n_564 ,csa_tree_add_7_45_groupi_n_245 ,in4[10]);
  xnor csa_tree_add_7_45_groupi_g4804__6783(csa_tree_add_7_45_groupi_n_562 ,csa_tree_add_7_45_groupi_n_280 ,in1[5]);
  and csa_tree_add_7_45_groupi_g4805__3680(csa_tree_add_7_45_groupi_n_561 ,csa_tree_add_7_45_groupi_n_359 ,csa_tree_add_7_45_groupi_n_421);
  and csa_tree_add_7_45_groupi_g4806__1617(csa_tree_add_7_45_groupi_n_560 ,csa_tree_add_7_45_groupi_n_125 ,csa_tree_add_7_45_groupi_n_380);
  and csa_tree_add_7_45_groupi_g4807__2802(csa_tree_add_7_45_groupi_n_558 ,csa_tree_add_7_45_groupi_n_454 ,csa_tree_add_7_45_groupi_n_455);
  not csa_tree_add_7_45_groupi_g4808(csa_tree_add_7_45_groupi_n_518 ,csa_tree_add_7_45_groupi_n_519);
  not csa_tree_add_7_45_groupi_g4809(csa_tree_add_7_45_groupi_n_517 ,csa_tree_add_7_45_groupi_n_516);
  not csa_tree_add_7_45_groupi_g4810(csa_tree_add_7_45_groupi_n_514 ,csa_tree_add_7_45_groupi_n_515);
  not csa_tree_add_7_45_groupi_g4811(csa_tree_add_7_45_groupi_n_510 ,csa_tree_add_7_45_groupi_n_511);
  not csa_tree_add_7_45_groupi_g4812(csa_tree_add_7_45_groupi_n_506 ,csa_tree_add_7_45_groupi_n_507);
  not csa_tree_add_7_45_groupi_g4813(csa_tree_add_7_45_groupi_n_505 ,csa_tree_add_7_45_groupi_n_504);
  not csa_tree_add_7_45_groupi_g4814(csa_tree_add_7_45_groupi_n_501 ,csa_tree_add_7_45_groupi_n_502);
  not csa_tree_add_7_45_groupi_g4815(csa_tree_add_7_45_groupi_n_497 ,csa_tree_add_7_45_groupi_n_498);
  not csa_tree_add_7_45_groupi_g4816(csa_tree_add_7_45_groupi_n_495 ,csa_tree_add_7_45_groupi_n_496);
  not csa_tree_add_7_45_groupi_g4817(csa_tree_add_7_45_groupi_n_491 ,csa_tree_add_7_45_groupi_n_492);
  not csa_tree_add_7_45_groupi_g4818(csa_tree_add_7_45_groupi_n_489 ,csa_tree_add_7_45_groupi_n_490);
  not csa_tree_add_7_45_groupi_g4819(csa_tree_add_7_45_groupi_n_487 ,csa_tree_add_7_45_groupi_n_488);
  not csa_tree_add_7_45_groupi_g4820(csa_tree_add_7_45_groupi_n_485 ,csa_tree_add_7_45_groupi_n_486);
  not csa_tree_add_7_45_groupi_g4821(csa_tree_add_7_45_groupi_n_483 ,csa_tree_add_7_45_groupi_n_484);
  not csa_tree_add_7_45_groupi_g4822(csa_tree_add_7_45_groupi_n_475 ,csa_tree_add_7_45_groupi_n_476);
  not csa_tree_add_7_45_groupi_g4823(csa_tree_add_7_45_groupi_n_472 ,csa_tree_add_7_45_groupi_n_473);
  not csa_tree_add_7_45_groupi_g4824(csa_tree_add_7_45_groupi_n_470 ,csa_tree_add_7_45_groupi_n_471);
  not csa_tree_add_7_45_groupi_g4825(csa_tree_add_7_45_groupi_n_468 ,csa_tree_add_7_45_groupi_n_469);
  not csa_tree_add_7_45_groupi_g4826(csa_tree_add_7_45_groupi_n_465 ,csa_tree_add_7_45_groupi_n_466);
  not csa_tree_add_7_45_groupi_g4827(csa_tree_add_7_45_groupi_n_463 ,csa_tree_add_7_45_groupi_n_462);
  not csa_tree_add_7_45_groupi_g4828(csa_tree_add_7_45_groupi_n_460 ,csa_tree_add_7_45_groupi_n_461);
  xnor csa_tree_add_7_45_groupi_g4829__1705(out1[0] ,csa_tree_add_7_45_groupi_n_283 ,in1[0]);
  xnor csa_tree_add_7_45_groupi_g4830__5122(csa_tree_add_7_45_groupi_n_458 ,csa_tree_add_7_45_groupi_n_306 ,in2[0]);
  xnor csa_tree_add_7_45_groupi_g4831__8246(csa_tree_add_7_45_groupi_n_457 ,csa_tree_add_7_45_groupi_n_305 ,in1[10]);
  xnor csa_tree_add_7_45_groupi_g4832__7098(csa_tree_add_7_45_groupi_n_524 ,csa_tree_add_7_45_groupi_n_308 ,csa_tree_add_7_45_groupi_n_250);
  xnor csa_tree_add_7_45_groupi_g4833__6131(csa_tree_add_7_45_groupi_n_523 ,csa_tree_add_7_45_groupi_n_268 ,in1[9]);
  xnor csa_tree_add_7_45_groupi_g4834__1881(csa_tree_add_7_45_groupi_n_522 ,csa_tree_add_7_45_groupi_n_256 ,in2[4]);
  xnor csa_tree_add_7_45_groupi_g4835__5115(csa_tree_add_7_45_groupi_n_521 ,csa_tree_add_7_45_groupi_n_297 ,in4[8]);
  xnor csa_tree_add_7_45_groupi_g4836__7482(csa_tree_add_7_45_groupi_n_520 ,csa_tree_add_7_45_groupi_n_301 ,in4[9]);
  xnor csa_tree_add_7_45_groupi_g4837__4733(csa_tree_add_7_45_groupi_n_519 ,csa_tree_add_7_45_groupi_n_257 ,in2[1]);
  xnor csa_tree_add_7_45_groupi_g4838__6161(csa_tree_add_7_45_groupi_n_516 ,csa_tree_add_7_45_groupi_n_172 ,csa_tree_add_7_45_groupi_n_277);
  xnor csa_tree_add_7_45_groupi_g4839__9315(csa_tree_add_7_45_groupi_n_515 ,csa_tree_add_7_45_groupi_n_252 ,in2[1]);
  xnor csa_tree_add_7_45_groupi_g4840__9945(csa_tree_add_7_45_groupi_n_513 ,csa_tree_add_7_45_groupi_n_244 ,in4[11]);
  xnor csa_tree_add_7_45_groupi_g4841__2883(csa_tree_add_7_45_groupi_n_512 ,csa_tree_add_7_45_groupi_n_281 ,in4[6]);
  xnor csa_tree_add_7_45_groupi_g4842__2346(csa_tree_add_7_45_groupi_n_511 ,csa_tree_add_7_45_groupi_n_282 ,in4[6]);
  xnor csa_tree_add_7_45_groupi_g4843__1666(csa_tree_add_7_45_groupi_n_509 ,csa_tree_add_7_45_groupi_n_284 ,in4[5]);
  xnor csa_tree_add_7_45_groupi_g4844__7410(csa_tree_add_7_45_groupi_n_508 ,csa_tree_add_7_45_groupi_n_247 ,in1[11]);
  xnor csa_tree_add_7_45_groupi_g4845__6417(csa_tree_add_7_45_groupi_n_507 ,csa_tree_add_7_45_groupi_n_260 ,in4[8]);
  xnor csa_tree_add_7_45_groupi_g4846__5477(csa_tree_add_7_45_groupi_n_504 ,csa_tree_add_7_45_groupi_n_265 ,in2[14]);
  xnor csa_tree_add_7_45_groupi_g4847__2398(csa_tree_add_7_45_groupi_n_503 ,csa_tree_add_7_45_groupi_n_297 ,in4[12]);
  xnor csa_tree_add_7_45_groupi_g4848__5107(csa_tree_add_7_45_groupi_n_502 ,csa_tree_add_7_45_groupi_n_285 ,in4[1]);
  xnor csa_tree_add_7_45_groupi_g4849__6260(csa_tree_add_7_45_groupi_n_500 ,csa_tree_add_7_45_groupi_n_272 ,in4[3]);
  xnor csa_tree_add_7_45_groupi_g4850__4319(csa_tree_add_7_45_groupi_n_499 ,csa_tree_add_7_45_groupi_n_295 ,in4[11]);
  xnor csa_tree_add_7_45_groupi_g4851__8428(csa_tree_add_7_45_groupi_n_498 ,csa_tree_add_7_45_groupi_n_266 ,in4[2]);
  xnor csa_tree_add_7_45_groupi_g4852__5526(csa_tree_add_7_45_groupi_n_496 ,csa_tree_add_7_45_groupi_n_267 ,in1[14]);
  xnor csa_tree_add_7_45_groupi_g4853__6783(csa_tree_add_7_45_groupi_n_494 ,csa_tree_add_7_45_groupi_n_309 ,csa_tree_add_7_45_groupi_n_249);
  xnor csa_tree_add_7_45_groupi_g4854__3680(csa_tree_add_7_45_groupi_n_493 ,csa_tree_add_7_45_groupi_n_289 ,in4[1]);
  xnor csa_tree_add_7_45_groupi_g4855__1617(csa_tree_add_7_45_groupi_n_492 ,csa_tree_add_7_45_groupi_n_271 ,in2[10]);
  xnor csa_tree_add_7_45_groupi_g4856__2802(csa_tree_add_7_45_groupi_n_490 ,csa_tree_add_7_45_groupi_n_254 ,in4[7]);
  xnor csa_tree_add_7_45_groupi_g4857__1705(csa_tree_add_7_45_groupi_n_488 ,csa_tree_add_7_45_groupi_n_251 ,in1[12]);
  xnor csa_tree_add_7_45_groupi_g4858__5122(csa_tree_add_7_45_groupi_n_486 ,csa_tree_add_7_45_groupi_n_275 ,in2[3]);
  xnor csa_tree_add_7_45_groupi_g4859__8246(csa_tree_add_7_45_groupi_n_484 ,csa_tree_add_7_45_groupi_n_263 ,in1[13]);
  xnor csa_tree_add_7_45_groupi_g4860__7098(csa_tree_add_7_45_groupi_n_482 ,csa_tree_add_7_45_groupi_n_279 ,in4[2]);
  xnor csa_tree_add_7_45_groupi_g4861__6131(csa_tree_add_7_45_groupi_n_481 ,csa_tree_add_7_45_groupi_n_259 ,in4[10]);
  xnor csa_tree_add_7_45_groupi_g4862__1881(csa_tree_add_7_45_groupi_n_480 ,csa_tree_add_7_45_groupi_n_301 ,in1[14]);
  xnor csa_tree_add_7_45_groupi_g4863__5115(csa_tree_add_7_45_groupi_n_479 ,csa_tree_add_7_45_groupi_n_264 ,in1[11]);
  xnor csa_tree_add_7_45_groupi_g4864__7482(csa_tree_add_7_45_groupi_n_478 ,csa_tree_add_7_45_groupi_n_287 ,in4[7]);
  xnor csa_tree_add_7_45_groupi_g4865__4733(csa_tree_add_7_45_groupi_n_477 ,csa_tree_add_7_45_groupi_n_255 ,in1[1]);
  xnor csa_tree_add_7_45_groupi_g4866__6161(csa_tree_add_7_45_groupi_n_476 ,csa_tree_add_7_45_groupi_n_261 ,in1[12]);
  xnor csa_tree_add_7_45_groupi_g4867__9315(csa_tree_add_7_45_groupi_n_474 ,csa_tree_add_7_45_groupi_n_295 ,in1[14]);
  xnor csa_tree_add_7_45_groupi_g4868__9945(csa_tree_add_7_45_groupi_n_473 ,csa_tree_add_7_45_groupi_n_274 ,in4[7]);
  xnor csa_tree_add_7_45_groupi_g4869__2883(csa_tree_add_7_45_groupi_n_471 ,csa_tree_add_7_45_groupi_n_273 ,in4[13]);
  xnor csa_tree_add_7_45_groupi_g4870__2346(csa_tree_add_7_45_groupi_n_469 ,csa_tree_add_7_45_groupi_n_288 ,in4[9]);
  xnor csa_tree_add_7_45_groupi_g4871__1666(csa_tree_add_7_45_groupi_n_467 ,csa_tree_add_7_45_groupi_n_173 ,csa_tree_add_7_45_groupi_n_246);
  xnor csa_tree_add_7_45_groupi_g4872__7410(csa_tree_add_7_45_groupi_n_466 ,csa_tree_add_7_45_groupi_n_286 ,in1[3]);
  xnor csa_tree_add_7_45_groupi_g4873__6417(csa_tree_add_7_45_groupi_n_464 ,csa_tree_add_7_45_groupi_n_276 ,in4[4]);
  xnor csa_tree_add_7_45_groupi_g4874__5477(csa_tree_add_7_45_groupi_n_462 ,csa_tree_add_7_45_groupi_n_270 ,in1[15]);
  xnor csa_tree_add_7_45_groupi_g4875__2398(csa_tree_add_7_45_groupi_n_461 ,csa_tree_add_7_45_groupi_n_248 ,in4[9]);
  not csa_tree_add_7_45_groupi_g4876(csa_tree_add_7_45_groupi_n_456 ,csa_tree_add_7_45_groupi_n_455);
  not csa_tree_add_7_45_groupi_g4877(csa_tree_add_7_45_groupi_n_454 ,csa_tree_add_7_45_groupi_n_453);
  not csa_tree_add_7_45_groupi_g4878(csa_tree_add_7_45_groupi_n_438 ,csa_tree_add_7_45_groupi_n_439);
  not csa_tree_add_7_45_groupi_g4879(csa_tree_add_7_45_groupi_n_435 ,csa_tree_add_7_45_groupi_n_436);
  not csa_tree_add_7_45_groupi_g4880(csa_tree_add_7_45_groupi_n_432 ,csa_tree_add_7_45_groupi_n_431);
  not csa_tree_add_7_45_groupi_g4881(csa_tree_add_7_45_groupi_n_430 ,csa_tree_add_7_45_groupi_n_429);
  or csa_tree_add_7_45_groupi_g4883__5107(csa_tree_add_7_45_groupi_n_425 ,csa_tree_add_7_45_groupi_n_166 ,csa_tree_add_7_45_groupi_n_299);
  or csa_tree_add_7_45_groupi_g4884__6260(csa_tree_add_7_45_groupi_n_424 ,in1[0] ,csa_tree_add_7_45_groupi_n_290);
  nor csa_tree_add_7_45_groupi_g4885__4319(csa_tree_add_7_45_groupi_n_423 ,csa_tree_add_7_45_groupi_n_63 ,csa_tree_add_7_45_groupi_n_303);
  nor csa_tree_add_7_45_groupi_g4886__8428(csa_tree_add_7_45_groupi_n_422 ,csa_tree_add_7_45_groupi_n_167 ,csa_tree_add_7_45_groupi_n_298);
  or csa_tree_add_7_45_groupi_g4887__5526(csa_tree_add_7_45_groupi_n_421 ,csa_tree_add_7_45_groupi_n_360 ,csa_tree_add_7_45_groupi_n_306);
  nor csa_tree_add_7_45_groupi_g4888__6783(csa_tree_add_7_45_groupi_n_420 ,csa_tree_add_7_45_groupi_n_83 ,csa_tree_add_7_45_groupi_n_291);
  or csa_tree_add_7_45_groupi_g4889__3680(csa_tree_add_7_45_groupi_n_419 ,csa_tree_add_7_45_groupi_n_144 ,csa_tree_add_7_45_groupi_n_308);
  nor csa_tree_add_7_45_groupi_g4890__1617(csa_tree_add_7_45_groupi_n_418 ,csa_tree_add_7_45_groupi_n_240 ,csa_tree_add_7_45_groupi_n_310);
  and csa_tree_add_7_45_groupi_g4891__2802(csa_tree_add_7_45_groupi_n_455 ,csa_tree_add_7_45_groupi_n_155 ,csa_tree_add_7_45_groupi_n_318);
  or csa_tree_add_7_45_groupi_g4892__1705(csa_tree_add_7_45_groupi_n_453 ,csa_tree_add_7_45_groupi_n_176 ,csa_tree_add_7_45_groupi_n_350);
  and csa_tree_add_7_45_groupi_g4893__5122(csa_tree_add_7_45_groupi_n_452 ,csa_tree_add_7_45_groupi_n_212 ,csa_tree_add_7_45_groupi_n_319);
  and csa_tree_add_7_45_groupi_g4894__8246(csa_tree_add_7_45_groupi_n_451 ,csa_tree_add_7_45_groupi_n_131 ,csa_tree_add_7_45_groupi_n_367);
  and csa_tree_add_7_45_groupi_g4895__7098(csa_tree_add_7_45_groupi_n_450 ,csa_tree_add_7_45_groupi_n_207 ,csa_tree_add_7_45_groupi_n_316);
  and csa_tree_add_7_45_groupi_g4896__6131(csa_tree_add_7_45_groupi_n_449 ,csa_tree_add_7_45_groupi_n_239 ,csa_tree_add_7_45_groupi_n_353);
  and csa_tree_add_7_45_groupi_g4897__1881(csa_tree_add_7_45_groupi_n_448 ,csa_tree_add_7_45_groupi_n_126 ,csa_tree_add_7_45_groupi_n_324);
  or csa_tree_add_7_45_groupi_g4898__5115(csa_tree_add_7_45_groupi_n_447 ,csa_tree_add_7_45_groupi_n_175 ,csa_tree_add_7_45_groupi_n_351);
  and csa_tree_add_7_45_groupi_g4899__7482(csa_tree_add_7_45_groupi_n_446 ,csa_tree_add_7_45_groupi_n_132 ,csa_tree_add_7_45_groupi_n_314);
  and csa_tree_add_7_45_groupi_g4900__4733(csa_tree_add_7_45_groupi_n_445 ,csa_tree_add_7_45_groupi_n_229 ,csa_tree_add_7_45_groupi_n_329);
  and csa_tree_add_7_45_groupi_g4901__6161(csa_tree_add_7_45_groupi_n_444 ,csa_tree_add_7_45_groupi_n_205 ,csa_tree_add_7_45_groupi_n_315);
  or csa_tree_add_7_45_groupi_g4902__9315(csa_tree_add_7_45_groupi_n_443 ,csa_tree_add_7_45_groupi_n_136 ,csa_tree_add_7_45_groupi_n_345);
  and csa_tree_add_7_45_groupi_g4903__9945(csa_tree_add_7_45_groupi_n_442 ,csa_tree_add_7_45_groupi_n_191 ,csa_tree_add_7_45_groupi_n_334);
  and csa_tree_add_7_45_groupi_g4904__2883(csa_tree_add_7_45_groupi_n_441 ,csa_tree_add_7_45_groupi_n_174 ,csa_tree_add_7_45_groupi_n_365);
  or csa_tree_add_7_45_groupi_g4905__2346(csa_tree_add_7_45_groupi_n_440 ,csa_tree_add_7_45_groupi_n_200 ,csa_tree_add_7_45_groupi_n_317);
  or csa_tree_add_7_45_groupi_g4906__1666(csa_tree_add_7_45_groupi_n_439 ,csa_tree_add_7_45_groupi_n_152 ,csa_tree_add_7_45_groupi_n_355);
  or csa_tree_add_7_45_groupi_g4907__7410(csa_tree_add_7_45_groupi_n_437 ,csa_tree_add_7_45_groupi_n_197 ,csa_tree_add_7_45_groupi_n_336);
  or csa_tree_add_7_45_groupi_g4908__6417(csa_tree_add_7_45_groupi_n_436 ,csa_tree_add_7_45_groupi_n_153 ,csa_tree_add_7_45_groupi_n_335);
  and csa_tree_add_7_45_groupi_g4909__5477(csa_tree_add_7_45_groupi_n_434 ,csa_tree_add_7_45_groupi_n_208 ,csa_tree_add_7_45_groupi_n_352);
  or csa_tree_add_7_45_groupi_g4910__2398(csa_tree_add_7_45_groupi_n_433 ,csa_tree_add_7_45_groupi_n_201 ,csa_tree_add_7_45_groupi_n_332);
  and csa_tree_add_7_45_groupi_g4911__5107(csa_tree_add_7_45_groupi_n_431 ,csa_tree_add_7_45_groupi_n_185 ,csa_tree_add_7_45_groupi_n_342);
  or csa_tree_add_7_45_groupi_g4912__6260(csa_tree_add_7_45_groupi_n_429 ,csa_tree_add_7_45_groupi_n_149 ,csa_tree_add_7_45_groupi_n_325);
  and csa_tree_add_7_45_groupi_g4913__4319(csa_tree_add_7_45_groupi_n_428 ,csa_tree_add_7_45_groupi_n_213 ,csa_tree_add_7_45_groupi_n_344);
  or csa_tree_add_7_45_groupi_g4914__8428(csa_tree_add_7_45_groupi_n_427 ,csa_tree_add_7_45_groupi_n_133 ,csa_tree_add_7_45_groupi_n_323);
  or csa_tree_add_7_45_groupi_g4915__5526(csa_tree_add_7_45_groupi_n_426 ,csa_tree_add_7_45_groupi_n_241 ,csa_tree_add_7_45_groupi_n_311);
  not csa_tree_add_7_45_groupi_g4916(csa_tree_add_7_45_groupi_n_417 ,csa_tree_add_7_45_groupi_n_416);
  not csa_tree_add_7_45_groupi_g4919(csa_tree_add_7_45_groupi_n_398 ,csa_tree_add_7_45_groupi_n_399);
  not csa_tree_add_7_45_groupi_g4920(csa_tree_add_7_45_groupi_n_396 ,csa_tree_add_7_45_groupi_n_397);
  not csa_tree_add_7_45_groupi_g4921(csa_tree_add_7_45_groupi_n_394 ,csa_tree_add_7_45_groupi_n_395);
  not csa_tree_add_7_45_groupi_g4922(csa_tree_add_7_45_groupi_n_393 ,csa_tree_add_7_45_groupi_n_392);
  not csa_tree_add_7_45_groupi_g4923(csa_tree_add_7_45_groupi_n_389 ,csa_tree_add_7_45_groupi_n_390);
  not csa_tree_add_7_45_groupi_g4924(csa_tree_add_7_45_groupi_n_387 ,csa_tree_add_7_45_groupi_n_386);
  not csa_tree_add_7_45_groupi_g4925(csa_tree_add_7_45_groupi_n_384 ,csa_tree_add_7_45_groupi_n_385);
  and csa_tree_add_7_45_groupi_g4926__6783(csa_tree_add_7_45_groupi_n_383 ,csa_tree_add_7_45_groupi_n_348 ,csa_tree_add_7_45_groupi_n_307);
  nor csa_tree_add_7_45_groupi_g4927__3680(csa_tree_add_7_45_groupi_n_382 ,in1[10] ,csa_tree_add_7_45_groupi_n_305);
  or csa_tree_add_7_45_groupi_g4928__1617(csa_tree_add_7_45_groupi_n_381 ,csa_tree_add_7_45_groupi_n_74 ,csa_tree_add_7_45_groupi_n_304);
  or csa_tree_add_7_45_groupi_g4929__2802(csa_tree_add_7_45_groupi_n_380 ,csa_tree_add_7_45_groupi_n_181 ,csa_tree_add_7_45_groupi_n_309);
  or csa_tree_add_7_45_groupi_g4930__1705(csa_tree_add_7_45_groupi_n_379 ,in4[0] ,csa_tree_add_7_45_groupi_n_302);
  xnor csa_tree_add_7_45_groupi_g4931__5122(csa_tree_add_7_45_groupi_n_378 ,csa_tree_add_7_45_groupi_n_237 ,in2[2]);
  xnor csa_tree_add_7_45_groupi_g4932__8246(csa_tree_add_7_45_groupi_n_377 ,csa_tree_add_7_45_groupi_n_169 ,in2[9]);
  xnor csa_tree_add_7_45_groupi_g4933__7098(csa_tree_add_7_45_groupi_n_376 ,csa_tree_add_7_45_groupi_n_236 ,in2[14]);
  or csa_tree_add_7_45_groupi_g4934__6131(csa_tree_add_7_45_groupi_n_416 ,csa_tree_add_7_45_groupi_n_127 ,csa_tree_add_7_45_groupi_n_361);
  or csa_tree_add_7_45_groupi_g4935__1881(csa_tree_add_7_45_groupi_n_415 ,csa_tree_add_7_45_groupi_n_157 ,csa_tree_add_7_45_groupi_n_364);
  and csa_tree_add_7_45_groupi_g4936__5115(csa_tree_add_7_45_groupi_n_414 ,csa_tree_add_7_45_groupi_n_138 ,csa_tree_add_7_45_groupi_n_333);
  or csa_tree_add_7_45_groupi_g4937__7482(csa_tree_add_7_45_groupi_n_413 ,csa_tree_add_7_45_groupi_n_128 ,csa_tree_add_7_45_groupi_n_366);
  and csa_tree_add_7_45_groupi_g4938__4733(csa_tree_add_7_45_groupi_n_412 ,csa_tree_add_7_45_groupi_n_124 ,csa_tree_add_7_45_groupi_n_340);
  or csa_tree_add_7_45_groupi_g4939__6161(csa_tree_add_7_45_groupi_n_411 ,csa_tree_add_7_45_groupi_n_148 ,csa_tree_add_7_45_groupi_n_339);
  and csa_tree_add_7_45_groupi_g4940__9315(csa_tree_add_7_45_groupi_n_410 ,csa_tree_add_7_45_groupi_n_223 ,csa_tree_add_7_45_groupi_n_358);
  and csa_tree_add_7_45_groupi_g4941__9945(csa_tree_add_7_45_groupi_n_409 ,csa_tree_add_7_45_groupi_n_227 ,csa_tree_add_7_45_groupi_n_331);
  or csa_tree_add_7_45_groupi_g4942__2883(csa_tree_add_7_45_groupi_n_408 ,csa_tree_add_7_45_groupi_n_215 ,csa_tree_add_7_45_groupi_n_337);
  or csa_tree_add_7_45_groupi_g4943__2346(csa_tree_add_7_45_groupi_n_407 ,csa_tree_add_7_45_groupi_n_231 ,csa_tree_add_7_45_groupi_n_322);
  or csa_tree_add_7_45_groupi_g4944__1666(csa_tree_add_7_45_groupi_n_406 ,csa_tree_add_7_45_groupi_n_219 ,csa_tree_add_7_45_groupi_n_312);
  or csa_tree_add_7_45_groupi_g4945__7410(csa_tree_add_7_45_groupi_n_405 ,csa_tree_add_7_45_groupi_n_176 ,csa_tree_add_7_45_groupi_n_363);
  or csa_tree_add_7_45_groupi_g4946__6417(csa_tree_add_7_45_groupi_n_404 ,csa_tree_add_7_45_groupi_n_118 ,csa_tree_add_7_45_groupi_n_341);
  or csa_tree_add_7_45_groupi_g4947__5477(csa_tree_add_7_45_groupi_n_403 ,csa_tree_add_7_45_groupi_n_180 ,csa_tree_add_7_45_groupi_n_368);
  or csa_tree_add_7_45_groupi_g4948__2398(csa_tree_add_7_45_groupi_n_402 ,csa_tree_add_7_45_groupi_n_209 ,csa_tree_add_7_45_groupi_n_320);
  or csa_tree_add_7_45_groupi_g4949__5107(csa_tree_add_7_45_groupi_n_401 ,csa_tree_add_7_45_groupi_n_238 ,csa_tree_add_7_45_groupi_n_338);
  and csa_tree_add_7_45_groupi_g4950__6260(csa_tree_add_7_45_groupi_n_400 ,csa_tree_add_7_45_groupi_n_129 ,csa_tree_add_7_45_groupi_n_326);
  or csa_tree_add_7_45_groupi_g4951__4319(csa_tree_add_7_45_groupi_n_399 ,csa_tree_add_7_45_groupi_n_189 ,csa_tree_add_7_45_groupi_n_321);
  or csa_tree_add_7_45_groupi_g4952__8428(csa_tree_add_7_45_groupi_n_397 ,csa_tree_add_7_45_groupi_n_196 ,csa_tree_add_7_45_groupi_n_313);
  or csa_tree_add_7_45_groupi_g4953__5526(csa_tree_add_7_45_groupi_n_395 ,csa_tree_add_7_45_groupi_n_198 ,csa_tree_add_7_45_groupi_n_343);
  or csa_tree_add_7_45_groupi_g4954__6783(csa_tree_add_7_45_groupi_n_392 ,csa_tree_add_7_45_groupi_n_142 ,csa_tree_add_7_45_groupi_n_369);
  or csa_tree_add_7_45_groupi_g4955__3680(csa_tree_add_7_45_groupi_n_391 ,csa_tree_add_7_45_groupi_n_190 ,csa_tree_add_7_45_groupi_n_330);
  and csa_tree_add_7_45_groupi_g4956__1617(csa_tree_add_7_45_groupi_n_390 ,csa_tree_add_7_45_groupi_n_216 ,csa_tree_add_7_45_groupi_n_354);
  or csa_tree_add_7_45_groupi_g4957__2802(csa_tree_add_7_45_groupi_n_388 ,csa_tree_add_7_45_groupi_n_130 ,csa_tree_add_7_45_groupi_n_327);
  or csa_tree_add_7_45_groupi_g4958__1705(csa_tree_add_7_45_groupi_n_386 ,csa_tree_add_7_45_groupi_n_147 ,csa_tree_add_7_45_groupi_n_328);
  or csa_tree_add_7_45_groupi_g4959__5122(csa_tree_add_7_45_groupi_n_385 ,csa_tree_add_7_45_groupi_n_151 ,csa_tree_add_7_45_groupi_n_362);
  not csa_tree_add_7_45_groupi_g4960(csa_tree_add_7_45_groupi_n_375 ,csa_tree_add_7_45_groupi_n_374);
  not csa_tree_add_7_45_groupi_g4961(csa_tree_add_7_45_groupi_n_372 ,csa_tree_add_7_45_groupi_n_373);
  not csa_tree_add_7_45_groupi_g4962(csa_tree_add_7_45_groupi_n_371 ,csa_tree_add_7_45_groupi_n_370);
  nor csa_tree_add_7_45_groupi_g4963__8246(csa_tree_add_7_45_groupi_n_369 ,in2[8] ,csa_tree_add_7_45_groupi_n_182);
  and csa_tree_add_7_45_groupi_g4964__7098(csa_tree_add_7_45_groupi_n_368 ,in3[13] ,csa_tree_add_7_45_groupi_n_119);
  or csa_tree_add_7_45_groupi_g4965__6131(csa_tree_add_7_45_groupi_n_367 ,csa_tree_add_7_45_groupi_n_111 ,csa_tree_add_7_45_groupi_n_117);
  and csa_tree_add_7_45_groupi_g4966__1881(csa_tree_add_7_45_groupi_n_366 ,in3[5] ,csa_tree_add_7_45_groupi_n_122);
  or csa_tree_add_7_45_groupi_g4967__5115(csa_tree_add_7_45_groupi_n_365 ,csa_tree_add_7_45_groupi_n_109 ,csa_tree_add_7_45_groupi_n_179);
  and csa_tree_add_7_45_groupi_g4968__7482(csa_tree_add_7_45_groupi_n_364 ,in3[12] ,csa_tree_add_7_45_groupi_n_184);
  and csa_tree_add_7_45_groupi_g4969__4733(csa_tree_add_7_45_groupi_n_363 ,in3[14] ,csa_tree_add_7_45_groupi_n_177);
  and csa_tree_add_7_45_groupi_g4970__6161(csa_tree_add_7_45_groupi_n_362 ,in3[9] ,csa_tree_add_7_45_groupi_n_139);
  nor csa_tree_add_7_45_groupi_g4971__9315(csa_tree_add_7_45_groupi_n_361 ,csa_tree_add_7_45_groupi_n_86 ,csa_tree_add_7_45_groupi_n_116);
  and csa_tree_add_7_45_groupi_g4972__9945(csa_tree_add_7_45_groupi_n_360 ,csa_tree_add_7_45_groupi_n_103 ,csa_tree_add_7_45_groupi_n_170);
  or csa_tree_add_7_45_groupi_g4973__2883(csa_tree_add_7_45_groupi_n_359 ,csa_tree_add_7_45_groupi_n_103 ,csa_tree_add_7_45_groupi_n_170);
  or csa_tree_add_7_45_groupi_g4974__2346(csa_tree_add_7_45_groupi_n_358 ,in3[0] ,csa_tree_add_7_45_groupi_n_214);
  or csa_tree_add_7_45_groupi_g4975__1666(csa_tree_add_7_45_groupi_n_357 ,csa_tree_add_7_45_groupi_n_79 ,csa_tree_add_7_45_groupi_n_237);
  and csa_tree_add_7_45_groupi_g4976__7410(csa_tree_add_7_45_groupi_n_356 ,csa_tree_add_7_45_groupi_n_79 ,csa_tree_add_7_45_groupi_n_237);
  nor csa_tree_add_7_45_groupi_g4977__6417(csa_tree_add_7_45_groupi_n_355 ,csa_tree_add_7_45_groupi_n_98 ,csa_tree_add_7_45_groupi_n_146);
  or csa_tree_add_7_45_groupi_g4978__5477(csa_tree_add_7_45_groupi_n_354 ,in1[3] ,csa_tree_add_7_45_groupi_n_222);
  or csa_tree_add_7_45_groupi_g4979__2398(csa_tree_add_7_45_groupi_n_353 ,in1[3] ,csa_tree_add_7_45_groupi_n_243);
  or csa_tree_add_7_45_groupi_g4980__5107(csa_tree_add_7_45_groupi_n_352 ,in1[5] ,csa_tree_add_7_45_groupi_n_203);
  nor csa_tree_add_7_45_groupi_g4981__6260(csa_tree_add_7_45_groupi_n_351 ,csa_tree_add_7_45_groupi_n_78 ,csa_tree_add_7_45_groupi_n_179);
  nor csa_tree_add_7_45_groupi_g4982__4319(csa_tree_add_7_45_groupi_n_350 ,csa_tree_add_7_45_groupi_n_94 ,csa_tree_add_7_45_groupi_n_178);
  nor csa_tree_add_7_45_groupi_g4983__8428(csa_tree_add_7_45_groupi_n_349 ,csa_tree_add_7_45_groupi_n_77 ,csa_tree_add_7_45_groupi_n_169);
  or csa_tree_add_7_45_groupi_g4984__5526(csa_tree_add_7_45_groupi_n_348 ,in2[14] ,csa_tree_add_7_45_groupi_n_235);
  nor csa_tree_add_7_45_groupi_g4985__6783(csa_tree_add_7_45_groupi_n_347 ,csa_tree_add_7_45_groupi_n_96 ,csa_tree_add_7_45_groupi_n_236);
  or csa_tree_add_7_45_groupi_g4986__3680(csa_tree_add_7_45_groupi_n_346 ,in2[9] ,csa_tree_add_7_45_groupi_n_168);
  nor csa_tree_add_7_45_groupi_g4987__1617(csa_tree_add_7_45_groupi_n_345 ,csa_tree_add_7_45_groupi_n_69 ,csa_tree_add_7_45_groupi_n_134);
  or csa_tree_add_7_45_groupi_g4988__2802(csa_tree_add_7_45_groupi_n_344 ,csa_tree_add_7_45_groupi_n_80 ,csa_tree_add_7_45_groupi_n_224);
  and csa_tree_add_7_45_groupi_g4989__1705(csa_tree_add_7_45_groupi_n_343 ,in2[3] ,csa_tree_add_7_45_groupi_n_202);
  or csa_tree_add_7_45_groupi_g4990__5122(csa_tree_add_7_45_groupi_n_342 ,in2[2] ,csa_tree_add_7_45_groupi_n_120);
  nor csa_tree_add_7_45_groupi_g4991__8246(csa_tree_add_7_45_groupi_n_341 ,in2[4] ,csa_tree_add_7_45_groupi_n_143);
  or csa_tree_add_7_45_groupi_g4992__7098(csa_tree_add_7_45_groupi_n_340 ,in2[1] ,csa_tree_add_7_45_groupi_n_141);
  and csa_tree_add_7_45_groupi_g4993__6131(csa_tree_add_7_45_groupi_n_339 ,in3[11] ,csa_tree_add_7_45_groupi_n_154);
  and csa_tree_add_7_45_groupi_g4994__1881(csa_tree_add_7_45_groupi_n_338 ,in3[1] ,csa_tree_add_7_45_groupi_n_242);
  and csa_tree_add_7_45_groupi_g4995__5115(csa_tree_add_7_45_groupi_n_337 ,in2[3] ,csa_tree_add_7_45_groupi_n_217);
  and csa_tree_add_7_45_groupi_g4996__7482(csa_tree_add_7_45_groupi_n_336 ,in1[8] ,csa_tree_add_7_45_groupi_n_206);
  nor csa_tree_add_7_45_groupi_g4997__4733(csa_tree_add_7_45_groupi_n_335 ,csa_tree_add_7_45_groupi_n_173 ,csa_tree_add_7_45_groupi_n_135);
  or csa_tree_add_7_45_groupi_g4998__6161(csa_tree_add_7_45_groupi_n_334 ,csa_tree_add_7_45_groupi_n_82 ,csa_tree_add_7_45_groupi_n_186);
  or csa_tree_add_7_45_groupi_g4999__9315(csa_tree_add_7_45_groupi_n_333 ,in1[4] ,csa_tree_add_7_45_groupi_n_121);
  and csa_tree_add_7_45_groupi_g5000__9945(csa_tree_add_7_45_groupi_n_332 ,in2[2] ,csa_tree_add_7_45_groupi_n_199);
  or csa_tree_add_7_45_groupi_g5001__2883(csa_tree_add_7_45_groupi_n_331 ,csa_tree_add_7_45_groupi_n_172 ,csa_tree_add_7_45_groupi_n_228);
  and csa_tree_add_7_45_groupi_g5002__2346(csa_tree_add_7_45_groupi_n_330 ,in2[10] ,csa_tree_add_7_45_groupi_n_187);
  or csa_tree_add_7_45_groupi_g5003__1666(csa_tree_add_7_45_groupi_n_329 ,csa_tree_add_7_45_groupi_n_107 ,csa_tree_add_7_45_groupi_n_226);
  and csa_tree_add_7_45_groupi_g5004__7410(csa_tree_add_7_45_groupi_n_328 ,in2[7] ,csa_tree_add_7_45_groupi_n_145);
  nor csa_tree_add_7_45_groupi_g5005__6417(csa_tree_add_7_45_groupi_n_327 ,in2[5] ,csa_tree_add_7_45_groupi_n_211);
  or csa_tree_add_7_45_groupi_g5006__5477(csa_tree_add_7_45_groupi_n_326 ,in2[3] ,csa_tree_add_7_45_groupi_n_140);
  nor csa_tree_add_7_45_groupi_g5007__2398(csa_tree_add_7_45_groupi_n_325 ,in2[6] ,csa_tree_add_7_45_groupi_n_150);
  or csa_tree_add_7_45_groupi_g5008__5107(csa_tree_add_7_45_groupi_n_324 ,in2[9] ,csa_tree_add_7_45_groupi_n_221);
  nor csa_tree_add_7_45_groupi_g5009__6260(csa_tree_add_7_45_groupi_n_323 ,in2[7] ,csa_tree_add_7_45_groupi_n_158);
  and csa_tree_add_7_45_groupi_g5010__4319(csa_tree_add_7_45_groupi_n_322 ,in2[8] ,csa_tree_add_7_45_groupi_n_230);
  and csa_tree_add_7_45_groupi_g5011__8428(csa_tree_add_7_45_groupi_n_321 ,in2[5] ,csa_tree_add_7_45_groupi_n_188);
  and csa_tree_add_7_45_groupi_g5012__5526(csa_tree_add_7_45_groupi_n_320 ,in1[7] ,csa_tree_add_7_45_groupi_n_193);
  or csa_tree_add_7_45_groupi_g5013__6783(csa_tree_add_7_45_groupi_n_319 ,csa_tree_add_7_45_groupi_n_99 ,csa_tree_add_7_45_groupi_n_210);
  or csa_tree_add_7_45_groupi_g5014__3680(csa_tree_add_7_45_groupi_n_318 ,in2[12] ,csa_tree_add_7_45_groupi_n_115);
  and csa_tree_add_7_45_groupi_g5015__1617(csa_tree_add_7_45_groupi_n_317 ,in2[4] ,csa_tree_add_7_45_groupi_n_194);
  or csa_tree_add_7_45_groupi_g5016__2802(csa_tree_add_7_45_groupi_n_316 ,csa_tree_add_7_45_groupi_n_84 ,csa_tree_add_7_45_groupi_n_192);
  or csa_tree_add_7_45_groupi_g5017__1705(csa_tree_add_7_45_groupi_n_315 ,csa_tree_add_7_45_groupi_n_85 ,csa_tree_add_7_45_groupi_n_204);
  or csa_tree_add_7_45_groupi_g5018__5122(csa_tree_add_7_45_groupi_n_314 ,in2[14] ,csa_tree_add_7_45_groupi_n_156);
  and csa_tree_add_7_45_groupi_g5019__8246(csa_tree_add_7_45_groupi_n_313 ,in1[2] ,csa_tree_add_7_45_groupi_n_195);
  and csa_tree_add_7_45_groupi_g5020__7098(csa_tree_add_7_45_groupi_n_312 ,in2[0] ,csa_tree_add_7_45_groupi_n_225);
  or csa_tree_add_7_45_groupi_g5021__6131(csa_tree_add_7_45_groupi_n_374 ,csa_tree_add_7_45_groupi_n_183 ,csa_tree_add_7_45_groupi_n_37);
  or csa_tree_add_7_45_groupi_g5022__1881(csa_tree_add_7_45_groupi_n_373 ,csa_tree_add_7_45_groupi_n_232 ,csa_tree_add_7_45_groupi_n_220);
  or csa_tree_add_7_45_groupi_g5023__5115(csa_tree_add_7_45_groupi_n_370 ,csa_tree_add_7_45_groupi_n_56 ,csa_tree_add_7_45_groupi_n_123);
  not csa_tree_add_7_45_groupi_g5024(csa_tree_add_7_45_groupi_n_311 ,csa_tree_add_7_45_groupi_n_310);
  not csa_tree_add_7_45_groupi_g5025(csa_tree_add_7_45_groupi_n_304 ,csa_tree_add_7_45_groupi_n_305);
  not csa_tree_add_7_45_groupi_g5026(csa_tree_add_7_45_groupi_n_302 ,csa_tree_add_7_45_groupi_n_303);
  not csa_tree_add_7_45_groupi_g5027(csa_tree_add_7_45_groupi_n_298 ,csa_tree_add_7_45_groupi_n_299);
  not csa_tree_add_7_45_groupi_g5028(csa_tree_add_7_45_groupi_n_293 ,csa_tree_add_7_45_groupi_n_294);
  not csa_tree_add_7_45_groupi_g5029(csa_tree_add_7_45_groupi_n_291 ,csa_tree_add_7_45_groupi_n_290);
  xnor csa_tree_add_7_45_groupi_g5030__7482(csa_tree_add_7_45_groupi_n_289 ,in1[3] ,in1[1]);
  xnor csa_tree_add_7_45_groupi_g5031__4733(csa_tree_add_7_45_groupi_n_288 ,in2[8] ,in2[5]);
  xnor csa_tree_add_7_45_groupi_g5032__6161(csa_tree_add_7_45_groupi_n_287 ,in2[6] ,in2[3]);
  xnor csa_tree_add_7_45_groupi_g5033__9315(csa_tree_add_7_45_groupi_n_286 ,in4[6] ,in1[8]);
  xnor csa_tree_add_7_45_groupi_g5034__9945(csa_tree_add_7_45_groupi_n_285 ,in1[7] ,in1[2]);
  xnor csa_tree_add_7_45_groupi_g5035__2883(csa_tree_add_7_45_groupi_n_284 ,in1[11] ,in1[6]);
  xnor csa_tree_add_7_45_groupi_g5036__2346(csa_tree_add_7_45_groupi_n_283 ,in4[0] ,in3[0]);
  xnor csa_tree_add_7_45_groupi_g5037__1666(csa_tree_add_7_45_groupi_n_282 ,in4[0] ,in2[2]);
  xnor csa_tree_add_7_45_groupi_g5038__7410(csa_tree_add_7_45_groupi_n_281 ,in1[12] ,in1[7]);
  xnor csa_tree_add_7_45_groupi_g5039__6417(csa_tree_add_7_45_groupi_n_280 ,in4[5] ,in1[7]);
  xnor csa_tree_add_7_45_groupi_g5040__5477(csa_tree_add_7_45_groupi_n_279 ,in4[0] ,in1[4]);
  xnor csa_tree_add_7_45_groupi_g5041__2398(csa_tree_add_7_45_groupi_n_278 ,in4[3] ,in1[5]);
  xnor csa_tree_add_7_45_groupi_g5042__5107(csa_tree_add_7_45_groupi_n_277 ,in1[2] ,in2[1]);
  xnor csa_tree_add_7_45_groupi_g5043__6260(csa_tree_add_7_45_groupi_n_276 ,in1[10] ,in1[5]);
  xnor csa_tree_add_7_45_groupi_g5044__4319(csa_tree_add_7_45_groupi_n_275 ,in4[4] ,in1[4]);
  xnor csa_tree_add_7_45_groupi_g5045__8428(csa_tree_add_7_45_groupi_n_274 ,in1[13] ,in1[8]);
  xnor csa_tree_add_7_45_groupi_g5046__5526(csa_tree_add_7_45_groupi_n_273 ,in2[12] ,in2[9]);
  xnor csa_tree_add_7_45_groupi_g5047__6783(csa_tree_add_7_45_groupi_n_272 ,in1[9] ,in1[4]);
  xnor csa_tree_add_7_45_groupi_g5048__3680(csa_tree_add_7_45_groupi_n_271 ,in4[10] ,in2[13]);
  xnor csa_tree_add_7_45_groupi_g5049__1617(csa_tree_add_7_45_groupi_n_270 ,in4[6] ,in2[6]);
  xnor csa_tree_add_7_45_groupi_g5050__2802(csa_tree_add_7_45_groupi_n_269 ,in4[5] ,in3[5]);
  xnor csa_tree_add_7_45_groupi_g5051__1705(csa_tree_add_7_45_groupi_n_268 ,in4[0] ,in2[0]);
  xnor csa_tree_add_7_45_groupi_g5052__5122(csa_tree_add_7_45_groupi_n_267 ,in4[5] ,in2[5]);
  xnor csa_tree_add_7_45_groupi_g5053__8246(csa_tree_add_7_45_groupi_n_266 ,in4[6] ,in3[6]);
  xnor csa_tree_add_7_45_groupi_g5054__7098(csa_tree_add_7_45_groupi_n_265 ,in4[12] ,in4[11]);
  xnor csa_tree_add_7_45_groupi_g5055__6131(csa_tree_add_7_45_groupi_n_264 ,in4[2] ,in2[2]);
  xnor csa_tree_add_7_45_groupi_g5056__1881(csa_tree_add_7_45_groupi_n_263 ,in4[4] ,in2[4]);
  xnor csa_tree_add_7_45_groupi_g5057__5115(csa_tree_add_7_45_groupi_n_262 ,in4[14] ,in4[12]);
  xnor csa_tree_add_7_45_groupi_g5058__7482(csa_tree_add_7_45_groupi_n_261 ,in4[3] ,in2[3]);
  xnor csa_tree_add_7_45_groupi_g5059__4733(csa_tree_add_7_45_groupi_n_260 ,in4[12] ,in3[12]);
  xnor csa_tree_add_7_45_groupi_g5060__6161(csa_tree_add_7_45_groupi_n_310 ,in4[13] ,in4[12]);
  xnor csa_tree_add_7_45_groupi_g5061__9315(csa_tree_add_7_45_groupi_n_259 ,in2[9] ,in2[6]);
  xnor csa_tree_add_7_45_groupi_g5062__9945(csa_tree_add_7_45_groupi_n_258 ,in4[4] ,in1[1]);
  xnor csa_tree_add_7_45_groupi_g5063__2883(csa_tree_add_7_45_groupi_n_257 ,in4[3] ,in2[4]);
  xnor csa_tree_add_7_45_groupi_g5064__2346(csa_tree_add_7_45_groupi_n_256 ,in4[2] ,in2[7]);
  xnor csa_tree_add_7_45_groupi_g5065__1666(csa_tree_add_7_45_groupi_n_255 ,in4[1] ,in3[1]);
  xnor csa_tree_add_7_45_groupi_g5066__7410(csa_tree_add_7_45_groupi_n_254 ,in4[11] ,in3[11]);
  xnor csa_tree_add_7_45_groupi_g5067__6417(csa_tree_add_7_45_groupi_n_253 ,in4[9] ,in3[9]);
  xnor csa_tree_add_7_45_groupi_g5068__5477(csa_tree_add_7_45_groupi_n_252 ,in4[8] ,in4[1]);
  xnor csa_tree_add_7_45_groupi_g5069__2398(csa_tree_add_7_45_groupi_n_251 ,in4[15] ,in4[11]);
  xnor csa_tree_add_7_45_groupi_g5070__5107(csa_tree_add_7_45_groupi_n_250 ,in1[8] ,in1[6]);
  xnor csa_tree_add_7_45_groupi_g5071__6260(csa_tree_add_7_45_groupi_n_249 ,in1[10] ,in2[14]);
  xnor csa_tree_add_7_45_groupi_g5072__4319(csa_tree_add_7_45_groupi_n_248 ,in4[13] ,in3[13]);
  xnor csa_tree_add_7_45_groupi_g5073__8428(csa_tree_add_7_45_groupi_n_247 ,in4[14] ,in4[10]);
  xnor csa_tree_add_7_45_groupi_g5074__5526(csa_tree_add_7_45_groupi_n_246 ,in1[15] ,in2[13]);
  xnor csa_tree_add_7_45_groupi_g5075__6783(csa_tree_add_7_45_groupi_n_245 ,in4[14] ,in3[14]);
  xnor csa_tree_add_7_45_groupi_g5076__3680(csa_tree_add_7_45_groupi_n_244 ,in4[15] ,in3[15]);
  xnor csa_tree_add_7_45_groupi_g5077__1617(csa_tree_add_7_45_groupi_n_309 ,in4[15] ,in4[13]);
  xnor csa_tree_add_7_45_groupi_g5078__2802(csa_tree_add_7_45_groupi_n_308 ,in4[8] ,in3[8]);
  xnor csa_tree_add_7_45_groupi_g5079__1705(csa_tree_add_7_45_groupi_n_307 ,in4[15] ,in4[14]);
  xnor csa_tree_add_7_45_groupi_g5080__5122(csa_tree_add_7_45_groupi_n_306 ,in4[3] ,in3[3]);
  xnor csa_tree_add_7_45_groupi_g5081__8246(csa_tree_add_7_45_groupi_n_305 ,in4[10] ,in3[10]);
  xnor csa_tree_add_7_45_groupi_g5082__7098(csa_tree_add_7_45_groupi_n_303 ,in4[2] ,in3[2]);
  xnor csa_tree_add_7_45_groupi_g5083__6131(csa_tree_add_7_45_groupi_n_301 ,in2[15] ,in2[12]);
  and csa_tree_add_7_45_groupi_g5084__1881(csa_tree_add_7_45_groupi_n_300 ,csa_tree_add_7_45_groupi_n_234 ,csa_tree_add_7_45_groupi_n_218);
  xnor csa_tree_add_7_45_groupi_g5085__5115(csa_tree_add_7_45_groupi_n_299 ,in4[15] ,in2[15]);
  xnor csa_tree_add_7_45_groupi_g5086__7482(csa_tree_add_7_45_groupi_n_297 ,in2[11] ,in2[8]);
  xnor csa_tree_add_7_45_groupi_g5087__4733(csa_tree_add_7_45_groupi_n_296 ,in4[14] ,in4[13]);
  xnor csa_tree_add_7_45_groupi_g5088__6161(csa_tree_add_7_45_groupi_n_295 ,in2[10] ,in2[7]);
  xnor csa_tree_add_7_45_groupi_g5089__9315(csa_tree_add_7_45_groupi_n_294 ,in1[13] ,in2[11]);
  xnor csa_tree_add_7_45_groupi_g5090__9945(csa_tree_add_7_45_groupi_n_292 ,in4[4] ,in3[4]);
  xnor csa_tree_add_7_45_groupi_g5091__2883(csa_tree_add_7_45_groupi_n_290 ,csa_tree_add_7_45_groupi_n_69 ,in3[7]);
  not csa_tree_add_7_45_groupi_g5092(csa_tree_add_7_45_groupi_n_243 ,csa_tree_add_7_45_groupi_n_242);
  not csa_tree_add_7_45_groupi_g5093(csa_tree_add_7_45_groupi_n_241 ,csa_tree_add_7_45_groupi_n_240);
  not csa_tree_add_7_45_groupi_g5094(csa_tree_add_7_45_groupi_n_239 ,csa_tree_add_7_45_groupi_n_238);
  not csa_tree_add_7_45_groupi_g5095(csa_tree_add_7_45_groupi_n_235 ,csa_tree_add_7_45_groupi_n_236);
  not csa_tree_add_7_45_groupi_g5096(csa_tree_add_7_45_groupi_n_233 ,csa_tree_add_7_45_groupi_n_232);
  nor csa_tree_add_7_45_groupi_g5097__2346(csa_tree_add_7_45_groupi_n_231 ,csa_tree_add_7_45_groupi_n_91 ,in2[11]);
  or csa_tree_add_7_45_groupi_g5098__1666(csa_tree_add_7_45_groupi_n_230 ,csa_tree_add_7_45_groupi_n_104 ,in4[8]);
  or csa_tree_add_7_45_groupi_g5099__7410(csa_tree_add_7_45_groupi_n_229 ,csa_tree_add_7_45_groupi_n_75 ,in2[15]);
  and csa_tree_add_7_45_groupi_g5100__6417(csa_tree_add_7_45_groupi_n_228 ,in1[2] ,csa_tree_add_7_45_groupi_n_98);
  or csa_tree_add_7_45_groupi_g5101__5477(csa_tree_add_7_45_groupi_n_227 ,csa_tree_add_7_45_groupi_n_98 ,in1[2]);
  nor csa_tree_add_7_45_groupi_g5102__2398(csa_tree_add_7_45_groupi_n_226 ,csa_tree_add_7_45_groupi_n_106 ,in1[14]);
  or csa_tree_add_7_45_groupi_g5103__5107(csa_tree_add_7_45_groupi_n_225 ,csa_tree_add_7_45_groupi_n_97 ,in4[0]);
  nor csa_tree_add_7_45_groupi_g5104__6260(csa_tree_add_7_45_groupi_n_224 ,csa_tree_add_7_45_groupi_n_100 ,in4[6]);
  or csa_tree_add_7_45_groupi_g5105__4319(csa_tree_add_7_45_groupi_n_223 ,csa_tree_add_7_45_groupi_n_63 ,in1[0]);
  nor csa_tree_add_7_45_groupi_g5106__8428(csa_tree_add_7_45_groupi_n_222 ,csa_tree_add_7_45_groupi_n_82 ,in4[3]);
  nor csa_tree_add_7_45_groupi_g5107__5526(csa_tree_add_7_45_groupi_n_221 ,in4[13] ,in2[12]);
  nor csa_tree_add_7_45_groupi_g5108__6783(csa_tree_add_7_45_groupi_n_220 ,in1[6] ,in2[0]);
  nor csa_tree_add_7_45_groupi_g5109__3680(csa_tree_add_7_45_groupi_n_219 ,csa_tree_add_7_45_groupi_n_32 ,in1[9]);
  or csa_tree_add_7_45_groupi_g5110__1617(csa_tree_add_7_45_groupi_n_218 ,csa_tree_add_7_45_groupi_n_67 ,in1[15]);
  or csa_tree_add_7_45_groupi_g5111__2802(csa_tree_add_7_45_groupi_n_217 ,csa_tree_add_7_45_groupi_n_99 ,in4[4]);
  or csa_tree_add_7_45_groupi_g5112__1705(csa_tree_add_7_45_groupi_n_216 ,csa_tree_add_7_45_groupi_n_89 ,in1[5]);
  and csa_tree_add_7_45_groupi_g5113__5122(csa_tree_add_7_45_groupi_n_215 ,in4[4] ,csa_tree_add_7_45_groupi_n_99);
  nor csa_tree_add_7_45_groupi_g5114__8246(csa_tree_add_7_45_groupi_n_214 ,csa_tree_add_7_45_groupi_n_83 ,in4[0]);
  or csa_tree_add_7_45_groupi_g5115__7098(csa_tree_add_7_45_groupi_n_213 ,csa_tree_add_7_45_groupi_n_62 ,in1[15]);
  or csa_tree_add_7_45_groupi_g5116__6131(csa_tree_add_7_45_groupi_n_212 ,csa_tree_add_7_45_groupi_n_42 ,in1[9]);
  nor csa_tree_add_7_45_groupi_g5117__1881(csa_tree_add_7_45_groupi_n_211 ,in4[9] ,in2[8]);
  nor csa_tree_add_7_45_groupi_g5118__5115(csa_tree_add_7_45_groupi_n_210 ,csa_tree_add_7_45_groupi_n_97 ,in4[3]);
  nor csa_tree_add_7_45_groupi_g5119__7482(csa_tree_add_7_45_groupi_n_209 ,csa_tree_add_7_45_groupi_n_62 ,in1[12]);
  or csa_tree_add_7_45_groupi_g5120__4733(csa_tree_add_7_45_groupi_n_208 ,csa_tree_add_7_45_groupi_n_28 ,in1[7]);
  or csa_tree_add_7_45_groupi_g5121__6161(csa_tree_add_7_45_groupi_n_207 ,csa_tree_add_7_45_groupi_n_23 ,in1[8]);
  or csa_tree_add_7_45_groupi_g5122__9315(csa_tree_add_7_45_groupi_n_206 ,csa_tree_add_7_45_groupi_n_76 ,in4[7]);
  or csa_tree_add_7_45_groupi_g5123__9945(csa_tree_add_7_45_groupi_n_205 ,csa_tree_add_7_45_groupi_n_28 ,in1[11]);
  nor csa_tree_add_7_45_groupi_g5124__2883(csa_tree_add_7_45_groupi_n_204 ,csa_tree_add_7_45_groupi_n_46 ,in4[5]);
  nor csa_tree_add_7_45_groupi_g5125__2346(csa_tree_add_7_45_groupi_n_203 ,csa_tree_add_7_45_groupi_n_95 ,in4[5]);
  or csa_tree_add_7_45_groupi_g5126__1666(csa_tree_add_7_45_groupi_n_202 ,csa_tree_add_7_45_groupi_n_44 ,in4[3]);
  and csa_tree_add_7_45_groupi_g5127__7410(csa_tree_add_7_45_groupi_n_201 ,in4[2] ,csa_tree_add_7_45_groupi_n_46);
  nor csa_tree_add_7_45_groupi_g5128__6417(csa_tree_add_7_45_groupi_n_200 ,csa_tree_add_7_45_groupi_n_65 ,in1[13]);
  or csa_tree_add_7_45_groupi_g5129__5477(csa_tree_add_7_45_groupi_n_199 ,csa_tree_add_7_45_groupi_n_94 ,in4[2]);
  and csa_tree_add_7_45_groupi_g5130__2398(csa_tree_add_7_45_groupi_n_198 ,in4[3] ,csa_tree_add_7_45_groupi_n_78);
  nor csa_tree_add_7_45_groupi_g5131__5107(csa_tree_add_7_45_groupi_n_197 ,csa_tree_add_7_45_groupi_n_35 ,in1[13]);
  nor csa_tree_add_7_45_groupi_g5132__6260(csa_tree_add_7_45_groupi_n_196 ,csa_tree_add_7_45_groupi_n_90 ,in1[7]);
  or csa_tree_add_7_45_groupi_g5133__4319(csa_tree_add_7_45_groupi_n_195 ,csa_tree_add_7_45_groupi_n_95 ,in4[1]);
  or csa_tree_add_7_45_groupi_g5134__8428(csa_tree_add_7_45_groupi_n_194 ,csa_tree_add_7_45_groupi_n_76 ,in4[4]);
  or csa_tree_add_7_45_groupi_g5135__5526(csa_tree_add_7_45_groupi_n_193 ,csa_tree_add_7_45_groupi_n_44 ,in4[6]);
  nor csa_tree_add_7_45_groupi_g5136__6783(csa_tree_add_7_45_groupi_n_192 ,csa_tree_add_7_45_groupi_n_93 ,in4[6]);
  or csa_tree_add_7_45_groupi_g5137__3680(csa_tree_add_7_45_groupi_n_191 ,csa_tree_add_7_45_groupi_n_65 ,in1[10]);
  nor csa_tree_add_7_45_groupi_g5138__1617(csa_tree_add_7_45_groupi_n_190 ,csa_tree_add_7_45_groupi_n_70 ,in2[13]);
  nor csa_tree_add_7_45_groupi_g5139__2802(csa_tree_add_7_45_groupi_n_189 ,csa_tree_add_7_45_groupi_n_61 ,in1[14]);
  or csa_tree_add_7_45_groupi_g5140__1705(csa_tree_add_7_45_groupi_n_188 ,csa_tree_add_7_45_groupi_n_75 ,in4[5]);
  or csa_tree_add_7_45_groupi_g5141__5122(csa_tree_add_7_45_groupi_n_187 ,csa_tree_add_7_45_groupi_n_73 ,in4[10]);
  nor csa_tree_add_7_45_groupi_g5142__8246(csa_tree_add_7_45_groupi_n_186 ,csa_tree_add_7_45_groupi_n_74 ,in4[4]);
  or csa_tree_add_7_45_groupi_g5143__7098(csa_tree_add_7_45_groupi_n_185 ,csa_tree_add_7_45_groupi_n_23 ,csa_tree_add_7_45_groupi_n_31);
  or csa_tree_add_7_45_groupi_g5144__6131(csa_tree_add_7_45_groupi_n_184 ,in4[12] ,in4[8]);
  and csa_tree_add_7_45_groupi_g5145__1881(csa_tree_add_7_45_groupi_n_183 ,in4[8] ,in1[9]);
  nor csa_tree_add_7_45_groupi_g5146__5115(csa_tree_add_7_45_groupi_n_182 ,in4[12] ,in2[11]);
  nor csa_tree_add_7_45_groupi_g5147__7482(csa_tree_add_7_45_groupi_n_181 ,in1[10] ,in2[14]);
  and csa_tree_add_7_45_groupi_g5148__4733(csa_tree_add_7_45_groupi_n_180 ,in4[13] ,in4[9]);
  or csa_tree_add_7_45_groupi_g5149__6161(csa_tree_add_7_45_groupi_n_242 ,csa_tree_add_7_45_groupi_n_101 ,in4[1]);
  and csa_tree_add_7_45_groupi_g5150__9315(csa_tree_add_7_45_groupi_n_240 ,csa_tree_add_7_45_groupi_n_76 ,csa_tree_add_7_45_groupi_n_104);
  and csa_tree_add_7_45_groupi_g5151__9945(csa_tree_add_7_45_groupi_n_238 ,in4[1] ,csa_tree_add_7_45_groupi_n_101);
  or csa_tree_add_7_45_groupi_g5152__2883(csa_tree_add_7_45_groupi_n_237 ,csa_tree_add_7_45_groupi_n_48 ,csa_tree_add_7_45_groupi_n_114);
  or csa_tree_add_7_45_groupi_g5153__2346(csa_tree_add_7_45_groupi_n_236 ,csa_tree_add_7_45_groupi_n_92 ,csa_tree_add_7_45_groupi_n_71);
  or csa_tree_add_7_45_groupi_g5154__1666(csa_tree_add_7_45_groupi_n_234 ,csa_tree_add_7_45_groupi_n_100 ,in4[9]);
  and csa_tree_add_7_45_groupi_g5155__7410(csa_tree_add_7_45_groupi_n_232 ,in1[6] ,in2[0]);
  not csa_tree_add_7_45_groupi_g5156(csa_tree_add_7_45_groupi_n_178 ,csa_tree_add_7_45_groupi_n_177);
  not csa_tree_add_7_45_groupi_g5157(csa_tree_add_7_45_groupi_n_175 ,csa_tree_add_7_45_groupi_n_174);
  not csa_tree_add_7_45_groupi_g5158(csa_tree_add_7_45_groupi_n_168 ,csa_tree_add_7_45_groupi_n_169);
  not csa_tree_add_7_45_groupi_g5159(csa_tree_add_7_45_groupi_n_166 ,csa_tree_add_7_45_groupi_n_167);
  not csa_tree_add_7_45_groupi_g5160(csa_tree_add_7_45_groupi_n_164 ,csa_tree_add_7_45_groupi_n_165);
  not csa_tree_add_7_45_groupi_g5161(csa_tree_add_7_45_groupi_n_162 ,csa_tree_add_7_45_groupi_n_163);
  nor csa_tree_add_7_45_groupi_g5164__6417(csa_tree_add_7_45_groupi_n_158 ,in4[11] ,in2[10]);
  and csa_tree_add_7_45_groupi_g5165__5477(csa_tree_add_7_45_groupi_n_157 ,in4[12] ,in4[8]);
  nor csa_tree_add_7_45_groupi_g5166__2398(csa_tree_add_7_45_groupi_n_156 ,in4[12] ,in4[11]);
  or csa_tree_add_7_45_groupi_g5167__5107(csa_tree_add_7_45_groupi_n_155 ,csa_tree_add_7_45_groupi_n_67 ,csa_tree_add_7_45_groupi_n_106);
  or csa_tree_add_7_45_groupi_g5168__6260(csa_tree_add_7_45_groupi_n_154 ,in4[11] ,in4[7]);
  nor csa_tree_add_7_45_groupi_g5169__4319(csa_tree_add_7_45_groupi_n_153 ,csa_tree_add_7_45_groupi_n_100 ,csa_tree_add_7_45_groupi_n_73);
  nor csa_tree_add_7_45_groupi_g5170__8428(csa_tree_add_7_45_groupi_n_152 ,csa_tree_add_7_45_groupi_n_91 ,csa_tree_add_7_45_groupi_n_90);
  nor csa_tree_add_7_45_groupi_g5171__5526(csa_tree_add_7_45_groupi_n_151 ,csa_tree_add_7_45_groupi_n_67 ,csa_tree_add_7_45_groupi_n_29);
  nor csa_tree_add_7_45_groupi_g5172__6783(csa_tree_add_7_45_groupi_n_150 ,in4[10] ,in2[9]);
  nor csa_tree_add_7_45_groupi_g5173__3680(csa_tree_add_7_45_groupi_n_149 ,csa_tree_add_7_45_groupi_n_70 ,csa_tree_add_7_45_groupi_n_77);
  and csa_tree_add_7_45_groupi_g5174__1617(csa_tree_add_7_45_groupi_n_148 ,in4[11] ,in4[7]);
  nor csa_tree_add_7_45_groupi_g5175__2802(csa_tree_add_7_45_groupi_n_147 ,in1[14] ,in2[10]);
  nor csa_tree_add_7_45_groupi_g5176__1705(csa_tree_add_7_45_groupi_n_146 ,in4[8] ,in4[1]);
  or csa_tree_add_7_45_groupi_g5177__5122(csa_tree_add_7_45_groupi_n_145 ,csa_tree_add_7_45_groupi_n_75 ,csa_tree_add_7_45_groupi_n_102);
  nor csa_tree_add_7_45_groupi_g5178__8246(csa_tree_add_7_45_groupi_n_144 ,csa_tree_add_7_45_groupi_n_93 ,csa_tree_add_7_45_groupi_n_85);
  nor csa_tree_add_7_45_groupi_g5179__7098(csa_tree_add_7_45_groupi_n_143 ,in4[2] ,in2[7]);
  and csa_tree_add_7_45_groupi_g5180__6131(csa_tree_add_7_45_groupi_n_142 ,in4[12] ,in2[11]);
  nor csa_tree_add_7_45_groupi_g5181__1881(csa_tree_add_7_45_groupi_n_141 ,in4[3] ,in2[4]);
  nor csa_tree_add_7_45_groupi_g5182__5115(csa_tree_add_7_45_groupi_n_140 ,in4[7] ,in2[6]);
  or csa_tree_add_7_45_groupi_g5183__7482(csa_tree_add_7_45_groupi_n_139 ,in4[9] ,in4[5]);
  or csa_tree_add_7_45_groupi_g5184__4733(csa_tree_add_7_45_groupi_n_138 ,csa_tree_add_7_45_groupi_n_64 ,csa_tree_add_7_45_groupi_n_31);
  or csa_tree_add_7_45_groupi_g5185__6161(csa_tree_add_7_45_groupi_n_137 ,in1[8] ,in1[6]);
  and csa_tree_add_7_45_groupi_g5186__9315(csa_tree_add_7_45_groupi_n_136 ,in4[14] ,in4[12]);
  nor csa_tree_add_7_45_groupi_g5187__9945(csa_tree_add_7_45_groupi_n_135 ,in1[15] ,in2[13]);
  nor csa_tree_add_7_45_groupi_g5188__2883(csa_tree_add_7_45_groupi_n_134 ,in4[14] ,in4[12]);
  and csa_tree_add_7_45_groupi_g5189__2346(csa_tree_add_7_45_groupi_n_133 ,in4[11] ,in2[10]);
  or csa_tree_add_7_45_groupi_g5190__1666(csa_tree_add_7_45_groupi_n_132 ,csa_tree_add_7_45_groupi_n_66 ,csa_tree_add_7_45_groupi_n_68);
  or csa_tree_add_7_45_groupi_g5191__7410(csa_tree_add_7_45_groupi_n_131 ,csa_tree_add_7_45_groupi_n_22 ,csa_tree_add_7_45_groupi_n_64);
  and csa_tree_add_7_45_groupi_g5192__6417(csa_tree_add_7_45_groupi_n_130 ,in4[9] ,in2[8]);
  or csa_tree_add_7_45_groupi_g5193__5477(csa_tree_add_7_45_groupi_n_129 ,csa_tree_add_7_45_groupi_n_34 ,csa_tree_add_7_45_groupi_n_80);
  nor csa_tree_add_7_45_groupi_g5194__2398(csa_tree_add_7_45_groupi_n_128 ,csa_tree_add_7_45_groupi_n_61 ,csa_tree_add_7_45_groupi_n_90);
  nor csa_tree_add_7_45_groupi_g5195__5107(csa_tree_add_7_45_groupi_n_127 ,csa_tree_add_7_45_groupi_n_48 ,csa_tree_add_7_45_groupi_n_101);
  or csa_tree_add_7_45_groupi_g5196__6260(csa_tree_add_7_45_groupi_n_126 ,csa_tree_add_7_45_groupi_n_40 ,csa_tree_add_7_45_groupi_n_107);
  or csa_tree_add_7_45_groupi_g5197__4319(csa_tree_add_7_45_groupi_n_125 ,csa_tree_add_7_45_groupi_n_74 ,csa_tree_add_7_45_groupi_n_96);
  or csa_tree_add_7_45_groupi_g5198__8428(csa_tree_add_7_45_groupi_n_124 ,csa_tree_add_7_45_groupi_n_42 ,csa_tree_add_7_45_groupi_n_81);
  nor csa_tree_add_7_45_groupi_g5199__5526(csa_tree_add_7_45_groupi_n_123 ,in1[2] ,in1[0]);
  or csa_tree_add_7_45_groupi_g5200__6783(csa_tree_add_7_45_groupi_n_122 ,in4[5] ,in4[1]);
  nor csa_tree_add_7_45_groupi_g5201__3680(csa_tree_add_7_45_groupi_n_121 ,in4[2] ,in4[0]);
  nor csa_tree_add_7_45_groupi_g5202__1617(csa_tree_add_7_45_groupi_n_120 ,in4[6] ,in4[0]);
  or csa_tree_add_7_45_groupi_g5203__2802(csa_tree_add_7_45_groupi_n_119 ,in4[13] ,in4[9]);
  and csa_tree_add_7_45_groupi_g5204__1705(csa_tree_add_7_45_groupi_n_118 ,in4[2] ,in2[7]);
  nor csa_tree_add_7_45_groupi_g5205__5122(csa_tree_add_7_45_groupi_n_117 ,in4[6] ,in4[2]);
  nor csa_tree_add_7_45_groupi_g5206__8246(csa_tree_add_7_45_groupi_n_116 ,in4[4] ,in1[1]);
  nor csa_tree_add_7_45_groupi_g5207__7098(csa_tree_add_7_45_groupi_n_115 ,in4[9] ,in2[15]);
  and csa_tree_add_7_45_groupi_g5208__6131(csa_tree_add_7_45_groupi_n_179 ,csa_tree_add_7_45_groupi_n_72 ,csa_tree_add_7_45_groupi_n_68);
  or csa_tree_add_7_45_groupi_g5209__1881(csa_tree_add_7_45_groupi_n_177 ,in4[14] ,in4[10]);
  and csa_tree_add_7_45_groupi_g5210__5115(csa_tree_add_7_45_groupi_n_176 ,in4[14] ,in4[10]);
  or csa_tree_add_7_45_groupi_g5211__7482(csa_tree_add_7_45_groupi_n_174 ,csa_tree_add_7_45_groupi_n_26 ,csa_tree_add_7_45_groupi_n_68);
  or csa_tree_add_7_45_groupi_g5212__4733(csa_tree_add_7_45_groupi_n_173 ,csa_tree_add_7_45_groupi_n_40 ,csa_tree_add_7_45_groupi_n_66);
  or csa_tree_add_7_45_groupi_g5213__6161(csa_tree_add_7_45_groupi_n_172 ,csa_tree_add_7_45_groupi_n_89 ,csa_tree_add_7_45_groupi_n_87);
  or csa_tree_add_7_45_groupi_g5214(csa_tree_add_7_45_groupi_n_171 ,csa_tree_add_7_45_groupi_n_34 ,csa_tree_add_7_45_groupi_n_112);
  or csa_tree_add_7_45_groupi_g5215(csa_tree_add_7_45_groupi_n_170 ,csa_tree_add_7_45_groupi_n_64 ,csa_tree_add_7_45_groupi_n_88);
  or csa_tree_add_7_45_groupi_g5216(csa_tree_add_7_45_groupi_n_169 ,csa_tree_add_7_45_groupi_n_26 ,csa_tree_add_7_45_groupi_n_71);
  and csa_tree_add_7_45_groupi_g5217(csa_tree_add_7_45_groupi_n_167 ,csa_tree_add_7_45_groupi_n_72 ,csa_tree_add_7_45_groupi_n_92);
  or csa_tree_add_7_45_groupi_g5218(csa_tree_add_7_45_groupi_n_165 ,csa_tree_add_7_45_groupi_n_70 ,csa_tree_add_7_45_groupi_n_113);
  or csa_tree_add_7_45_groupi_g5219(csa_tree_add_7_45_groupi_n_163 ,csa_tree_add_7_45_groupi_n_91 ,csa_tree_add_7_45_groupi_n_110);
  or csa_tree_add_7_45_groupi_g5220(csa_tree_add_7_45_groupi_n_161 ,csa_tree_add_7_45_groupi_n_105 ,csa_tree_add_7_45_groupi_n_83);
  or csa_tree_add_7_45_groupi_g5221(csa_tree_add_7_45_groupi_n_160 ,in4[8] ,in1[9]);
  and csa_tree_add_7_45_groupi_g5222(csa_tree_add_7_45_groupi_n_159 ,csa_tree_add_7_45_groupi_n_25 ,csa_tree_add_7_45_groupi_n_106);
  not csa_tree_add_7_45_groupi_g5223(csa_tree_add_7_45_groupi_n_114 ,in3[4]);
  not csa_tree_add_7_45_groupi_g5224(csa_tree_add_7_45_groupi_n_113 ,in3[10]);
  not csa_tree_add_7_45_groupi_g5225(csa_tree_add_7_45_groupi_n_112 ,in3[7]);
  not csa_tree_add_7_45_groupi_g5226(csa_tree_add_7_45_groupi_n_111 ,in3[6]);
  not csa_tree_add_7_45_groupi_g5227(csa_tree_add_7_45_groupi_n_110 ,in3[8]);
  not csa_tree_add_7_45_groupi_g5228(csa_tree_add_7_45_groupi_n_109 ,in3[15]);
  not csa_tree_add_7_45_groupi_g5229(csa_tree_add_7_45_groupi_n_108 ,in3[0]);
  not csa_tree_add_7_45_groupi_g5230(csa_tree_add_7_45_groupi_n_107 ,in2[12]);
  not csa_tree_add_7_45_groupi_g5231(csa_tree_add_7_45_groupi_n_106 ,in2[15]);
  not csa_tree_add_7_45_groupi_g5232(csa_tree_add_7_45_groupi_n_105 ,in1[2]);
  not csa_tree_add_7_45_groupi_g5233(csa_tree_add_7_45_groupi_n_104 ,in2[11]);
  not csa_tree_add_7_45_groupi_g5234(csa_tree_add_7_45_groupi_n_103 ,in2[0]);
  not csa_tree_add_7_45_groupi_g5235(csa_tree_add_7_45_groupi_n_102 ,in2[10]);
  not csa_tree_add_7_45_groupi_g5236(csa_tree_add_7_45_groupi_n_101 ,in1[1]);
  not csa_tree_add_7_45_groupi_g5237(csa_tree_add_7_45_groupi_n_100 ,in1[15]);
  not csa_tree_add_7_45_groupi_g5238(csa_tree_add_7_45_groupi_n_99 ,in1[4]);
  not csa_tree_add_7_45_groupi_g5239(csa_tree_add_7_45_groupi_n_98 ,in2[1]);
  not csa_tree_add_7_45_groupi_g5240(csa_tree_add_7_45_groupi_n_97 ,in1[9]);
  not csa_tree_add_7_45_groupi_g5241(csa_tree_add_7_45_groupi_n_96 ,in2[14]);
  not csa_tree_add_7_45_groupi_g5242(csa_tree_add_7_45_groupi_n_95 ,in1[7]);
  not csa_tree_add_7_45_groupi_g5243(csa_tree_add_7_45_groupi_n_94 ,in1[11]);
  not csa_tree_add_7_45_groupi_g5244(csa_tree_add_7_45_groupi_n_93 ,in1[8]);
  not csa_tree_add_7_45_groupi_g5245(csa_tree_add_7_45_groupi_n_92 ,in4[14]);
  not csa_tree_add_7_45_groupi_g5246(csa_tree_add_7_45_groupi_n_91 ,in4[8]);
  not csa_tree_add_7_45_groupi_g5247(csa_tree_add_7_45_groupi_n_90 ,in4[1]);
  not csa_tree_add_7_45_groupi_g5248(csa_tree_add_7_45_groupi_n_89 ,in4[3]);
  not csa_tree_add_7_45_groupi_g5249(csa_tree_add_7_45_groupi_n_88 ,in3[2]);
  not csa_tree_add_7_45_groupi_g5250(csa_tree_add_7_45_groupi_n_87 ,in3[3]);
  not csa_tree_add_7_45_groupi_g5251(csa_tree_add_7_45_groupi_n_86 ,in2[5]);
  not csa_tree_add_7_45_groupi_g5252(csa_tree_add_7_45_groupi_n_85 ,in1[6]);
  not csa_tree_add_7_45_groupi_g5253(csa_tree_add_7_45_groupi_n_84 ,in1[3]);
  not csa_tree_add_7_45_groupi_g5254(csa_tree_add_7_45_groupi_n_83 ,in1[0]);
  not csa_tree_add_7_45_groupi_g5255(csa_tree_add_7_45_groupi_n_82 ,in1[5]);
  not csa_tree_add_7_45_groupi_g5256(csa_tree_add_7_45_groupi_n_81 ,in2[4]);
  not csa_tree_add_7_45_groupi_g5257(csa_tree_add_7_45_groupi_n_80 ,in2[6]);
  not csa_tree_add_7_45_groupi_g5258(csa_tree_add_7_45_groupi_n_79 ,in2[2]);
  not csa_tree_add_7_45_groupi_g5259(csa_tree_add_7_45_groupi_n_78 ,in1[12]);
  not csa_tree_add_7_45_groupi_g5260(csa_tree_add_7_45_groupi_n_77 ,in2[9]);
  not csa_tree_add_7_45_groupi_g5261(csa_tree_add_7_45_groupi_n_76 ,in1[13]);
  not csa_tree_add_7_45_groupi_g5262(csa_tree_add_7_45_groupi_n_75 ,in1[14]);
  not csa_tree_add_7_45_groupi_g5263(csa_tree_add_7_45_groupi_n_74 ,in1[10]);
  not csa_tree_add_7_45_groupi_g5264(csa_tree_add_7_45_groupi_n_73 ,in2[13]);
  not csa_tree_add_7_45_groupi_g5265(csa_tree_add_7_45_groupi_n_72 ,in4[15]);
  not csa_tree_add_7_45_groupi_g5266(csa_tree_add_7_45_groupi_n_71 ,in4[13]);
  not csa_tree_add_7_45_groupi_g5267(csa_tree_add_7_45_groupi_n_70 ,in4[10]);
  not csa_tree_add_7_45_groupi_g5268(csa_tree_add_7_45_groupi_n_69 ,in4[7]);
  not csa_tree_add_7_45_groupi_g5269(csa_tree_add_7_45_groupi_n_68 ,in4[11]);
  not csa_tree_add_7_45_groupi_g5270(csa_tree_add_7_45_groupi_n_67 ,in4[9]);
  not csa_tree_add_7_45_groupi_g5271(csa_tree_add_7_45_groupi_n_66 ,in4[12]);
  not csa_tree_add_7_45_groupi_g5272(csa_tree_add_7_45_groupi_n_65 ,in4[4]);
  not csa_tree_add_7_45_groupi_g5273(csa_tree_add_7_45_groupi_n_64 ,in4[2]);
  not csa_tree_add_7_45_groupi_g5274(csa_tree_add_7_45_groupi_n_63 ,in4[0]);
  not csa_tree_add_7_45_groupi_g5275(csa_tree_add_7_45_groupi_n_62 ,in4[6]);
  not csa_tree_add_7_45_groupi_g5276(csa_tree_add_7_45_groupi_n_61 ,in4[5]);
  not csa_tree_add_7_45_groupi_drc_bufs5297(csa_tree_add_7_45_groupi_n_55 ,csa_tree_add_7_45_groupi_n_54);
  not csa_tree_add_7_45_groupi_drc_bufs5298(csa_tree_add_7_45_groupi_n_54 ,csa_tree_add_7_45_groupi_n_234);
  not csa_tree_add_7_45_groupi_drc_bufs5301(csa_tree_add_7_45_groupi_n_53 ,csa_tree_add_7_45_groupi_n_56);
  not csa_tree_add_7_45_groupi_drc_bufs5302(csa_tree_add_7_45_groupi_n_56 ,csa_tree_add_7_45_groupi_n_161);
  not csa_tree_add_7_45_groupi_drc_bufs5305(csa_tree_add_7_45_groupi_n_52 ,csa_tree_add_7_45_groupi_n_57);
  not csa_tree_add_7_45_groupi_drc_bufs5306(csa_tree_add_7_45_groupi_n_57 ,csa_tree_add_7_45_groupi_n_426);
  not csa_tree_add_7_45_groupi_drc_bufs5309(csa_tree_add_7_45_groupi_n_51 ,csa_tree_add_7_45_groupi_n_50);
  not csa_tree_add_7_45_groupi_drc_bufs5310(csa_tree_add_7_45_groupi_n_50 ,csa_tree_add_7_45_groupi_n_159);
  not csa_tree_add_7_45_groupi_drc_bufs5313(csa_tree_add_7_45_groupi_n_49 ,csa_tree_add_7_45_groupi_n_58);
  not csa_tree_add_7_45_groupi_drc_bufs5314(csa_tree_add_7_45_groupi_n_58 ,csa_tree_add_7_45_groupi_n_558);
  not csa_tree_add_7_45_groupi_drc_bufs5317(csa_tree_add_7_45_groupi_n_48 ,csa_tree_add_7_45_groupi_n_47);
  not csa_tree_add_7_45_groupi_drc_bufs5318(csa_tree_add_7_45_groupi_n_47 ,csa_tree_add_7_45_groupi_n_65);
  not csa_tree_add_7_45_groupi_drc_bufs5321(csa_tree_add_7_45_groupi_n_46 ,csa_tree_add_7_45_groupi_n_45);
  not csa_tree_add_7_45_groupi_drc_bufs5322(csa_tree_add_7_45_groupi_n_45 ,csa_tree_add_7_45_groupi_n_94);
  not csa_tree_add_7_45_groupi_drc_bufs5325(csa_tree_add_7_45_groupi_n_44 ,csa_tree_add_7_45_groupi_n_43);
  not csa_tree_add_7_45_groupi_drc_bufs5326(csa_tree_add_7_45_groupi_n_43 ,csa_tree_add_7_45_groupi_n_78);
  not csa_tree_add_7_45_groupi_drc_bufs5329(csa_tree_add_7_45_groupi_n_42 ,csa_tree_add_7_45_groupi_n_41);
  not csa_tree_add_7_45_groupi_drc_bufs5330(csa_tree_add_7_45_groupi_n_41 ,csa_tree_add_7_45_groupi_n_89);
  not csa_tree_add_7_45_groupi_drc_bufs5333(csa_tree_add_7_45_groupi_n_40 ,csa_tree_add_7_45_groupi_n_39);
  not csa_tree_add_7_45_groupi_drc_bufs5334(csa_tree_add_7_45_groupi_n_39 ,csa_tree_add_7_45_groupi_n_71);
  not csa_tree_add_7_45_groupi_drc_bufs5336(csa_tree_add_7_45_groupi_n_38 ,csa_tree_add_7_45_groupi_n_232);
  not csa_tree_add_7_45_groupi_drc_bufs5340(csa_tree_add_7_45_groupi_n_37 ,csa_tree_add_7_45_groupi_n_160);
  not csa_tree_add_7_45_groupi_drc_bufs5346(csa_tree_add_7_45_groupi_n_60 ,csa_tree_add_7_45_groupi_n_705);
  not csa_tree_add_7_45_groupi_drc_bufs5349(csa_tree_add_7_45_groupi_n_36 ,csa_tree_add_7_45_groupi_n_59);
  not csa_tree_add_7_45_groupi_drc_bufs5350(csa_tree_add_7_45_groupi_n_59 ,csa_tree_add_7_45_groupi_n_704);
  not csa_tree_add_7_45_groupi_drc_bufs5352(csa_tree_add_7_45_groupi_n_35 ,csa_tree_add_7_45_groupi_n_33);
  not csa_tree_add_7_45_groupi_drc_bufs5353(csa_tree_add_7_45_groupi_n_34 ,csa_tree_add_7_45_groupi_n_33);
  not csa_tree_add_7_45_groupi_drc_bufs5354(csa_tree_add_7_45_groupi_n_33 ,csa_tree_add_7_45_groupi_n_69);
  not csa_tree_add_7_45_groupi_drc_bufs5356(csa_tree_add_7_45_groupi_n_32 ,csa_tree_add_7_45_groupi_n_30);
  not csa_tree_add_7_45_groupi_drc_bufs5357(csa_tree_add_7_45_groupi_n_31 ,csa_tree_add_7_45_groupi_n_30);
  not csa_tree_add_7_45_groupi_drc_bufs5358(csa_tree_add_7_45_groupi_n_30 ,csa_tree_add_7_45_groupi_n_63);
  not csa_tree_add_7_45_groupi_drc_bufs5360(csa_tree_add_7_45_groupi_n_29 ,csa_tree_add_7_45_groupi_n_27);
  not csa_tree_add_7_45_groupi_drc_bufs5361(csa_tree_add_7_45_groupi_n_28 ,csa_tree_add_7_45_groupi_n_27);
  not csa_tree_add_7_45_groupi_drc_bufs5362(csa_tree_add_7_45_groupi_n_27 ,csa_tree_add_7_45_groupi_n_61);
  not csa_tree_add_7_45_groupi_drc_bufs5364(csa_tree_add_7_45_groupi_n_26 ,csa_tree_add_7_45_groupi_n_24);
  not csa_tree_add_7_45_groupi_drc_bufs5365(csa_tree_add_7_45_groupi_n_25 ,csa_tree_add_7_45_groupi_n_24);
  not csa_tree_add_7_45_groupi_drc_bufs5366(csa_tree_add_7_45_groupi_n_24 ,csa_tree_add_7_45_groupi_n_72);
  not csa_tree_add_7_45_groupi_drc_bufs5368(csa_tree_add_7_45_groupi_n_23 ,csa_tree_add_7_45_groupi_n_21);
  not csa_tree_add_7_45_groupi_drc_bufs5369(csa_tree_add_7_45_groupi_n_22 ,csa_tree_add_7_45_groupi_n_21);
  not csa_tree_add_7_45_groupi_drc_bufs5370(csa_tree_add_7_45_groupi_n_21 ,csa_tree_add_7_45_groupi_n_62);
  xor csa_tree_add_7_45_groupi_g2(out1[18] ,csa_tree_add_7_45_groupi_n_1258 ,csa_tree_add_7_45_groupi_n_1222);
  xor csa_tree_add_7_45_groupi_g5372(out1[17] ,csa_tree_add_7_45_groupi_n_1256 ,csa_tree_add_7_45_groupi_n_1223);
  xor csa_tree_add_7_45_groupi_g5373(out1[15] ,csa_tree_add_7_45_groupi_n_1251 ,csa_tree_add_7_45_groupi_n_1234);
  xor csa_tree_add_7_45_groupi_g5374(out1[13] ,csa_tree_add_7_45_groupi_n_1246 ,csa_tree_add_7_45_groupi_n_1224);
  xor csa_tree_add_7_45_groupi_g5375(out1[12] ,csa_tree_add_7_45_groupi_n_1244 ,csa_tree_add_7_45_groupi_n_1225);
  xor csa_tree_add_7_45_groupi_g5376(out1[11] ,csa_tree_add_7_45_groupi_n_1242 ,csa_tree_add_7_45_groupi_n_1206);
  xor csa_tree_add_7_45_groupi_g5377(out1[10] ,csa_tree_add_7_45_groupi_n_1240 ,csa_tree_add_7_45_groupi_n_1205);
  xor csa_tree_add_7_45_groupi_g5378(out1[9] ,csa_tree_add_7_45_groupi_n_1238 ,csa_tree_add_7_45_groupi_n_1184);
  xor csa_tree_add_7_45_groupi_g5379(out1[8] ,csa_tree_add_7_45_groupi_n_1236 ,csa_tree_add_7_45_groupi_n_1155);
  xor csa_tree_add_7_45_groupi_g5380(out1[7] ,csa_tree_add_7_45_groupi_n_1221 ,csa_tree_add_7_45_groupi_n_1127);
  xor csa_tree_add_7_45_groupi_g5381(csa_tree_add_7_45_groupi_n_10 ,csa_tree_add_7_45_groupi_n_1125 ,csa_tree_add_7_45_groupi_n_1129);
  xor csa_tree_add_7_45_groupi_g5382(csa_tree_add_7_45_groupi_n_9 ,csa_tree_add_7_45_groupi_n_1123 ,csa_tree_add_7_45_groupi_n_1156);
  xor csa_tree_add_7_45_groupi_g5383(csa_tree_add_7_45_groupi_n_8 ,csa_tree_add_7_45_groupi_n_1108 ,csa_tree_add_7_45_groupi_n_1158);
  xor csa_tree_add_7_45_groupi_g5384(csa_tree_add_7_45_groupi_n_7 ,csa_tree_add_7_45_groupi_n_1067 ,csa_tree_add_7_45_groupi_n_1130);
  xor csa_tree_add_7_45_groupi_g5385(csa_tree_add_7_45_groupi_n_6 ,csa_tree_add_7_45_groupi_n_1047 ,csa_tree_add_7_45_groupi_n_962);
  xor csa_tree_add_7_45_groupi_g5386(csa_tree_add_7_45_groupi_n_5 ,csa_tree_add_7_45_groupi_n_1044 ,csa_tree_add_7_45_groupi_n_954);
  xor csa_tree_add_7_45_groupi_g5387(csa_tree_add_7_45_groupi_n_4 ,csa_tree_add_7_45_groupi_n_737 ,csa_tree_add_7_45_groupi_n_698);
  xor csa_tree_add_7_45_groupi_g5388(csa_tree_add_7_45_groupi_n_3 ,csa_tree_add_7_45_groupi_n_414 ,csa_tree_add_7_45_groupi_n_378);
  xor csa_tree_add_7_45_groupi_g5389(csa_tree_add_7_45_groupi_n_2 ,csa_tree_add_7_45_groupi_n_412 ,csa_tree_add_7_45_groupi_n_589);
  xor csa_tree_add_7_45_groupi_g5390(csa_tree_add_7_45_groupi_n_1 ,csa_tree_add_7_45_groupi_n_580 ,csa_tree_add_7_45_groupi_n_160);
  xor csa_tree_add_7_45_groupi_g5391(csa_tree_add_7_45_groupi_n_0 ,csa_tree_add_7_45_groupi_n_740 ,csa_tree_add_7_45_groupi_n_60);
endmodule
