// Benchmark "top" written by ABC on Mon Jun 12 20:57:39 2023

module top ( 
    \1_n1 , \1_n1013 , \1_n1014 , \1_n1025 , \1_n1030 , \1_n1042 ,
    \1_n1049 , \1_n1052 , \1_n1058 , \1_n1065 , \1_n107 , \1_n1070 ,
    \1_n1091 , \1_n1093 , \1_n1098 , \1_n1099 , \1_n1108 , \1_n1121 ,
    \1_n1131 , \1_n1134 , \1_n1143 , \1_n1146 , \1_n1150 , \1_n1161 ,
    \1_n1162 , \1_n1165 , \1_n1170 , \1_n1184 , \1_n1187 , \1_n1189 ,
    \1_n120 , \1_n1223 , \1_n1240 , \1_n1243 , \1_n1251 , \1_n1253 ,
    \1_n1255 , \1_n1276 , \1_n128 , \1_n1280 , \1_n1303 , \1_n1310 ,
    \1_n1311 , \1_n1331 , \1_n1335 , \1_n1339 , \1_n135 , \1_n1361 ,
    \1_n1366 , \1_n137 , \1_n1373 , \1_n1378 , \1_n1389 , \1_n1396 ,
    \1_n1398 , \1_n1407 , \1_n1409 , \1_n1412 , \1_n1413 , \1_n1418 ,
    \1_n1422 , \1_n1425 , \1_n1438 , \1_n145 , \1_n147 , \1_n1475 ,
    \1_n1479 , \1_n1485 , \1_n1508 , \1_n1511 , \1_n1515 , \1_n1518 ,
    \1_n1530 , \1_n1545 , \1_n1549 , \1_n1551 , \1_n1555 , \1_n1562 ,
    \1_n1575 , \1_n1580 , \1_n1581 , \1_n1596 , \1_n1606 , \1_n1620 ,
    \1_n1630 , \1_n1648 , \1_n1655 , \1_n1676 , \1_n182 , \1_n184 ,
    \1_n198 , \1_n209 , \1_n220 , \1_n222 , \1_n230 , \1_n233 , \1_n268 ,
    \1_n283 , \1_n289 , \1_n290 , \1_n293 , \1_n296 , \1_n325 , \1_n330 ,
    \1_n342 , \1_n356 , \1_n362 , \1_n365 , \1_n373 , \1_n386 , \1_n403 ,
    \1_n415 , \1_n418 , \1_n421 , \1_n432 , \1_n468 , \1_n478 , \1_n481 ,
    \1_n490 , \1_n507 , \1_n514 , \1_n526 , \1_n532 , \1_n574 , \1_n576 ,
    \1_n579 , \1_n588 , \1_n596 , \1_n605 , \1_n615 , \1_n629 , \1_n635 ,
    \1_n646 , \1_n654 , \1_n664 , \1_n67 , \1_n677 , \1_n69 , \1_n704 ,
    \1_n710 , \1_n716 , \1_n726 , \1_n727 , \1_n737 , \1_n750 , \1_n751 ,
    \1_n765 , \1_n769 , \1_n793 , \1_n794 , \1_n797 , \1_n818 , \1_n824 ,
    \1_n829 , \1_n835 , \1_n837 , \1_n84 , \1_n842 , \1_n848 , \1_n851 ,
    \1_n857 , \1_n859 , \1_n869 , \1_n877 , \1_n9 , \1_n901 , \1_n909 ,
    \1_n923 , \1_n933 , \1_n934 , \1_n938 , \1_n950 , \1_n956 , \1_n96 ,
    \1_n973 , \1_n974 , \1_n989 , \1_n990 , \2_n1016 , \2_n1033 ,
    \2_n1039 , \2_n1043 , \2_n1058 , \2_n1088 , \2_n1095 , \2_n1097 ,
    \2_n1100 , \2_n1119 , \2_n1125 , \2_n1135 , \2_n1150 , \2_n1172 ,
    \2_n1175 , \2_n1177 , \2_n1180 , \2_n1181 , \2_n1182 , \2_n119 ,
    \2_n12 , \2_n1205 , \2_n1207 , \2_n1219 , \2_n1227 , \2_n1238 ,
    \2_n1279 , \2_n128 , \2_n1281 , \2_n1288 , \2_n1299 , \2_n132 ,
    \2_n1338 , \2_n1353 , \2_n1357 , \2_n1361 , \2_n1362 , \2_n1363 ,
    \2_n1366 , \2_n1391 , \2_n1396 , \2_n1402 , \2_n1406 , \2_n1408 ,
    \2_n1426 , \2_n1427 , \2_n1435 , \2_n1436 , \2_n1454 , \2_n1463 ,
    \2_n1471 , \2_n1485 , \2_n1498 , \2_n1503 , \2_n1515 , \2_n1518 ,
    \2_n1519 , \2_n1534 , \2_n1540 , \2_n1553 , \2_n1568 , \2_n157 ,
    \2_n1575 , \2_n1598 , \2_n1613 , \2_n1632 , \2_n1633 , \2_n1649 ,
    \2_n1655 , \2_n1660 , \2_n1663 , \2_n1674 , \2_n1675 , \2_n1700 ,
    \2_n1707 , \2_n1729 , \2_n1740 , \2_n1743 , \2_n1753 , \2_n1755 ,
    \2_n1756 , \2_n1768 , \2_n1788 , \2_n179 , \2_n1790 , \2_n186 ,
    \2_n187 , \2_n19 , \2_n190 , \2_n228 , \2_n236 , \2_n238 , \2_n239 ,
    \2_n257 , \2_n261 , \2_n270 , \2_n288 , \2_n297 , \2_n307 , \2_n319 ,
    \2_n321 , \2_n326 , \2_n33 , \2_n335 , \2_n342 , \2_n371 , \2_n377 ,
    \2_n378 , \2_n38 , \2_n380 , \2_n384 , \2_n386 , \2_n387 , \2_n389 ,
    \2_n39 , \2_n403 , \2_n448 , \2_n457 , \2_n482 , \2_n488 , \2_n495 ,
    \2_n504 , \2_n516 , \2_n520 , \2_n530 , \2_n541 , \2_n544 , \2_n560 ,
    \2_n564 , \2_n565 , \2_n566 , \2_n579 , \2_n591 , \2_n60 , \2_n600 ,
    \2_n601 , \2_n606 , \2_n617 , \2_n627 , \2_n636 , \2_n64 , \2_n643 ,
    \2_n668 , \2_n676 , \2_n697 , \2_n7 , \2_n708 , \2_n714 , \2_n715 ,
    \2_n721 , \2_n754 , \2_n758 , \2_n760 , \2_n77 , \2_n779 , \2_n801 ,
    \2_n807 , \2_n813 , \2_n830 , \2_n84 , \2_n841 , \2_n850 , \2_n887 ,
    \2_n894 , \2_n9 , \2_n912 , \2_n917 , \2_n918 , \2_n92 , \2_n937 ,
    \2_n946 , \2_n955 , \2_n961 , \2_n962 , \2_n966 , \2_n971 , \2_n984 ,
    \2_n999 ,
    \1_n1019 , \1_n1021 , \1_n1023 , \1_n1026 , \1_n1032 , \1_n1036 ,
    \1_n1039 , \1_n1043 , \1_n110 , \1_n1117 , \1_n1122 , \1_n1138 ,
    \1_n1151 , \1_n1157 , \1_n1160 , \1_n117 , \1_n1177 , \1_n1192 ,
    \1_n1194 , \1_n1198 , \1_n1239 , \1_n1275 , \1_n1314 , \1_n1375 ,
    \1_n1392 , \1_n1411 , \1_n142 , \1_n1442 , \1_n1454 , \1_n1474 ,
    \1_n1478 , \1_n150 , \1_n1512 , \1_n1531 , \1_n154 , \1_n1542 ,
    \1_n1547 , \1_n1552 , \1_n1556 , \1_n1574 , \1_n1589 , \1_n1594 ,
    \1_n1601 , \1_n1604 , \1_n1628 , \1_n1629 , \1_n1631 , \1_n1645 ,
    \1_n1665 , \1_n167 , \1_n1671 , \1_n170 , \1_n172 , \1_n190 , \1_n204 ,
    \1_n21 , \1_n210 , \1_n231 , \1_n232 , \1_n24 , \1_n240 , \1_n253 ,
    \1_n265 , \1_n269 , \1_n291 , \1_n292 , \1_n313 , \1_n32 , \1_n324 ,
    \1_n336 , \1_n347 , \1_n350 , \1_n363 , \1_n364 , \1_n368 , \1_n383 ,
    \1_n388 , \1_n427 , \1_n434 , \1_n476 , \1_n480 , \1_n489 , \1_n506 ,
    \1_n524 , \1_n54 , \1_n543 , \1_n565 , \1_n598 , \1_n608 , \1_n61 ,
    \1_n614 , \1_n618 , \1_n623 , \1_n633 , \1_n64 , \1_n640 , \1_n656 ,
    \1_n663 , \1_n675 , \1_n676 , \1_n678 , \1_n691 , \1_n693 , \1_n717 ,
    \1_n722 , \1_n740 , \1_n76 , \1_n785 , \1_n786 , \1_n790 , \1_n8 ,
    \1_n800 , \1_n814 , \1_n821 , \1_n83 , \1_n836 , \1_n840 , \1_n845 ,
    \1_n887 , \1_n894 , \1_n928 , \1_n964 , \1_n97 , \2_n101 , \2_n1027 ,
    \2_n1044 , \2_n1047 , \2_n1050 , \2_n1065 , \2_n107 , \2_n1087 ,
    \2_n1096 , \2_n1110 , \2_n112 , \2_n1140 , \2_n1163 , \2_n117 ,
    \2_n1186 , \2_n1224 , \2_n123 , \2_n1233 , \2_n1269 , \2_n1270 ,
    \2_n129 , \2_n1297 , \2_n130 , \2_n1314 , \2_n1322 , \2_n1346 ,
    \2_n1355 , \2_n1370 , \2_n1377 , \2_n1378 , \2_n1390 , \2_n1409 ,
    \2_n1414 , \2_n1425 , \2_n1462 , \2_n1464 , \2_n1491 , \2_n1495 ,
    \2_n1510 , \2_n1511 , \2_n1543 , \2_n158 , \2_n1584 , \2_n1587 ,
    \2_n1631 , \2_n165 , \2_n1654 , \2_n1657 , \2_n1676 , \2_n168 ,
    \2_n1682 , \2_n1697 , \2_n1698 , \2_n1708 , \2_n1710 , \2_n1721 ,
    \2_n173 , \2_n1733 , \2_n1761 , \2_n1780 , \2_n1784 , \2_n1793 ,
    \2_n1794 , \2_n18 , \2_n193 , \2_n211 , \2_n222 , \2_n235 , \2_n245 ,
    \2_n249 , \2_n259 , \2_n262 , \2_n264 , \2_n315 , \2_n320 , \2_n337 ,
    \2_n357 , \2_n361 , \2_n370 , \2_n375 , \2_n379 , \2_n381 , \2_n413 ,
    \2_n417 , \2_n454 , \2_n456 , \2_n476 , \2_n487 , \2_n542 , \2_n547 ,
    \2_n56 , \2_n567 , \2_n574 , \2_n596 , \2_n61 , \2_n611 , \2_n623 ,
    \2_n635 , \2_n649 , \2_n66 , \2_n661 , \2_n67 , \2_n673 , \2_n722 ,
    \2_n75 , \2_n765 , \2_n776 , \2_n786 , \2_n793 , \2_n824 , \2_n83 ,
    \2_n840 , \2_n845 , \2_n849 , \2_n860 , \2_n878 , \2_n882 , \2_n889 ,
    \2_n944 , \2_n951 , \2_n964 , \2_n967 , \2_n974   );
  input  \1_n1 , \1_n1013 , \1_n1014 , \1_n1025 , \1_n1030 , \1_n1042 ,
    \1_n1049 , \1_n1052 , \1_n1058 , \1_n1065 , \1_n107 , \1_n1070 ,
    \1_n1091 , \1_n1093 , \1_n1098 , \1_n1099 , \1_n1108 , \1_n1121 ,
    \1_n1131 , \1_n1134 , \1_n1143 , \1_n1146 , \1_n1150 , \1_n1161 ,
    \1_n1162 , \1_n1165 , \1_n1170 , \1_n1184 , \1_n1187 , \1_n1189 ,
    \1_n120 , \1_n1223 , \1_n1240 , \1_n1243 , \1_n1251 , \1_n1253 ,
    \1_n1255 , \1_n1276 , \1_n128 , \1_n1280 , \1_n1303 , \1_n1310 ,
    \1_n1311 , \1_n1331 , \1_n1335 , \1_n1339 , \1_n135 , \1_n1361 ,
    \1_n1366 , \1_n137 , \1_n1373 , \1_n1378 , \1_n1389 , \1_n1396 ,
    \1_n1398 , \1_n1407 , \1_n1409 , \1_n1412 , \1_n1413 , \1_n1418 ,
    \1_n1422 , \1_n1425 , \1_n1438 , \1_n145 , \1_n147 , \1_n1475 ,
    \1_n1479 , \1_n1485 , \1_n1508 , \1_n1511 , \1_n1515 , \1_n1518 ,
    \1_n1530 , \1_n1545 , \1_n1549 , \1_n1551 , \1_n1555 , \1_n1562 ,
    \1_n1575 , \1_n1580 , \1_n1581 , \1_n1596 , \1_n1606 , \1_n1620 ,
    \1_n1630 , \1_n1648 , \1_n1655 , \1_n1676 , \1_n182 , \1_n184 ,
    \1_n198 , \1_n209 , \1_n220 , \1_n222 , \1_n230 , \1_n233 , \1_n268 ,
    \1_n283 , \1_n289 , \1_n290 , \1_n293 , \1_n296 , \1_n325 , \1_n330 ,
    \1_n342 , \1_n356 , \1_n362 , \1_n365 , \1_n373 , \1_n386 , \1_n403 ,
    \1_n415 , \1_n418 , \1_n421 , \1_n432 , \1_n468 , \1_n478 , \1_n481 ,
    \1_n490 , \1_n507 , \1_n514 , \1_n526 , \1_n532 , \1_n574 , \1_n576 ,
    \1_n579 , \1_n588 , \1_n596 , \1_n605 , \1_n615 , \1_n629 , \1_n635 ,
    \1_n646 , \1_n654 , \1_n664 , \1_n67 , \1_n677 , \1_n69 , \1_n704 ,
    \1_n710 , \1_n716 , \1_n726 , \1_n727 , \1_n737 , \1_n750 , \1_n751 ,
    \1_n765 , \1_n769 , \1_n793 , \1_n794 , \1_n797 , \1_n818 , \1_n824 ,
    \1_n829 , \1_n835 , \1_n837 , \1_n84 , \1_n842 , \1_n848 , \1_n851 ,
    \1_n857 , \1_n859 , \1_n869 , \1_n877 , \1_n9 , \1_n901 , \1_n909 ,
    \1_n923 , \1_n933 , \1_n934 , \1_n938 , \1_n950 , \1_n956 , \1_n96 ,
    \1_n973 , \1_n974 , \1_n989 , \1_n990 , \2_n1016 , \2_n1033 ,
    \2_n1039 , \2_n1043 , \2_n1058 , \2_n1088 , \2_n1095 , \2_n1097 ,
    \2_n1100 , \2_n1119 , \2_n1125 , \2_n1135 , \2_n1150 , \2_n1172 ,
    \2_n1175 , \2_n1177 , \2_n1180 , \2_n1181 , \2_n1182 , \2_n119 ,
    \2_n12 , \2_n1205 , \2_n1207 , \2_n1219 , \2_n1227 , \2_n1238 ,
    \2_n1279 , \2_n128 , \2_n1281 , \2_n1288 , \2_n1299 , \2_n132 ,
    \2_n1338 , \2_n1353 , \2_n1357 , \2_n1361 , \2_n1362 , \2_n1363 ,
    \2_n1366 , \2_n1391 , \2_n1396 , \2_n1402 , \2_n1406 , \2_n1408 ,
    \2_n1426 , \2_n1427 , \2_n1435 , \2_n1436 , \2_n1454 , \2_n1463 ,
    \2_n1471 , \2_n1485 , \2_n1498 , \2_n1503 , \2_n1515 , \2_n1518 ,
    \2_n1519 , \2_n1534 , \2_n1540 , \2_n1553 , \2_n1568 , \2_n157 ,
    \2_n1575 , \2_n1598 , \2_n1613 , \2_n1632 , \2_n1633 , \2_n1649 ,
    \2_n1655 , \2_n1660 , \2_n1663 , \2_n1674 , \2_n1675 , \2_n1700 ,
    \2_n1707 , \2_n1729 , \2_n1740 , \2_n1743 , \2_n1753 , \2_n1755 ,
    \2_n1756 , \2_n1768 , \2_n1788 , \2_n179 , \2_n1790 , \2_n186 ,
    \2_n187 , \2_n19 , \2_n190 , \2_n228 , \2_n236 , \2_n238 , \2_n239 ,
    \2_n257 , \2_n261 , \2_n270 , \2_n288 , \2_n297 , \2_n307 , \2_n319 ,
    \2_n321 , \2_n326 , \2_n33 , \2_n335 , \2_n342 , \2_n371 , \2_n377 ,
    \2_n378 , \2_n38 , \2_n380 , \2_n384 , \2_n386 , \2_n387 , \2_n389 ,
    \2_n39 , \2_n403 , \2_n448 , \2_n457 , \2_n482 , \2_n488 , \2_n495 ,
    \2_n504 , \2_n516 , \2_n520 , \2_n530 , \2_n541 , \2_n544 , \2_n560 ,
    \2_n564 , \2_n565 , \2_n566 , \2_n579 , \2_n591 , \2_n60 , \2_n600 ,
    \2_n601 , \2_n606 , \2_n617 , \2_n627 , \2_n636 , \2_n64 , \2_n643 ,
    \2_n668 , \2_n676 , \2_n697 , \2_n7 , \2_n708 , \2_n714 , \2_n715 ,
    \2_n721 , \2_n754 , \2_n758 , \2_n760 , \2_n77 , \2_n779 , \2_n801 ,
    \2_n807 , \2_n813 , \2_n830 , \2_n84 , \2_n841 , \2_n850 , \2_n887 ,
    \2_n894 , \2_n9 , \2_n912 , \2_n917 , \2_n918 , \2_n92 , \2_n937 ,
    \2_n946 , \2_n955 , \2_n961 , \2_n962 , \2_n966 , \2_n971 , \2_n984 ,
    \2_n999 ;
  output \1_n1019 , \1_n1021 , \1_n1023 , \1_n1026 , \1_n1032 , \1_n1036 ,
    \1_n1039 , \1_n1043 , \1_n110 , \1_n1117 , \1_n1122 , \1_n1138 ,
    \1_n1151 , \1_n1157 , \1_n1160 , \1_n117 , \1_n1177 , \1_n1192 ,
    \1_n1194 , \1_n1198 , \1_n1239 , \1_n1275 , \1_n1314 , \1_n1375 ,
    \1_n1392 , \1_n1411 , \1_n142 , \1_n1442 , \1_n1454 , \1_n1474 ,
    \1_n1478 , \1_n150 , \1_n1512 , \1_n1531 , \1_n154 , \1_n1542 ,
    \1_n1547 , \1_n1552 , \1_n1556 , \1_n1574 , \1_n1589 , \1_n1594 ,
    \1_n1601 , \1_n1604 , \1_n1628 , \1_n1629 , \1_n1631 , \1_n1645 ,
    \1_n1665 , \1_n167 , \1_n1671 , \1_n170 , \1_n172 , \1_n190 , \1_n204 ,
    \1_n21 , \1_n210 , \1_n231 , \1_n232 , \1_n24 , \1_n240 , \1_n253 ,
    \1_n265 , \1_n269 , \1_n291 , \1_n292 , \1_n313 , \1_n32 , \1_n324 ,
    \1_n336 , \1_n347 , \1_n350 , \1_n363 , \1_n364 , \1_n368 , \1_n383 ,
    \1_n388 , \1_n427 , \1_n434 , \1_n476 , \1_n480 , \1_n489 , \1_n506 ,
    \1_n524 , \1_n54 , \1_n543 , \1_n565 , \1_n598 , \1_n608 , \1_n61 ,
    \1_n614 , \1_n618 , \1_n623 , \1_n633 , \1_n64 , \1_n640 , \1_n656 ,
    \1_n663 , \1_n675 , \1_n676 , \1_n678 , \1_n691 , \1_n693 , \1_n717 ,
    \1_n722 , \1_n740 , \1_n76 , \1_n785 , \1_n786 , \1_n790 , \1_n8 ,
    \1_n800 , \1_n814 , \1_n821 , \1_n83 , \1_n836 , \1_n840 , \1_n845 ,
    \1_n887 , \1_n894 , \1_n928 , \1_n964 , \1_n97 , \2_n101 , \2_n1027 ,
    \2_n1044 , \2_n1047 , \2_n1050 , \2_n1065 , \2_n107 , \2_n1087 ,
    \2_n1096 , \2_n1110 , \2_n112 , \2_n1140 , \2_n1163 , \2_n117 ,
    \2_n1186 , \2_n1224 , \2_n123 , \2_n1233 , \2_n1269 , \2_n1270 ,
    \2_n129 , \2_n1297 , \2_n130 , \2_n1314 , \2_n1322 , \2_n1346 ,
    \2_n1355 , \2_n1370 , \2_n1377 , \2_n1378 , \2_n1390 , \2_n1409 ,
    \2_n1414 , \2_n1425 , \2_n1462 , \2_n1464 , \2_n1491 , \2_n1495 ,
    \2_n1510 , \2_n1511 , \2_n1543 , \2_n158 , \2_n1584 , \2_n1587 ,
    \2_n1631 , \2_n165 , \2_n1654 , \2_n1657 , \2_n1676 , \2_n168 ,
    \2_n1682 , \2_n1697 , \2_n1698 , \2_n1708 , \2_n1710 , \2_n1721 ,
    \2_n173 , \2_n1733 , \2_n1761 , \2_n1780 , \2_n1784 , \2_n1793 ,
    \2_n1794 , \2_n18 , \2_n193 , \2_n211 , \2_n222 , \2_n235 , \2_n245 ,
    \2_n249 , \2_n259 , \2_n262 , \2_n264 , \2_n315 , \2_n320 , \2_n337 ,
    \2_n357 , \2_n361 , \2_n370 , \2_n375 , \2_n379 , \2_n381 , \2_n413 ,
    \2_n417 , \2_n454 , \2_n456 , \2_n476 , \2_n487 , \2_n542 , \2_n547 ,
    \2_n56 , \2_n567 , \2_n574 , \2_n596 , \2_n61 , \2_n611 , \2_n623 ,
    \2_n635 , \2_n649 , \2_n66 , \2_n661 , \2_n67 , \2_n673 , \2_n722 ,
    \2_n75 , \2_n765 , \2_n776 , \2_n786 , \2_n793 , \2_n824 , \2_n83 ,
    \2_n840 , \2_n845 , \2_n849 , \2_n860 , \2_n878 , \2_n882 , \2_n889 ,
    \2_n944 , \2_n951 , \2_n964 , \2_n967 , \2_n974 ;
  wire new_n603_, new_n604_, new_n605_, new_n606_, new_n607_, new_n608_,
    new_n609_, new_n610_, new_n611_, new_n612_, new_n613_, new_n614_,
    new_n615_, new_n616_, new_n617_, new_n618_, new_n619_, new_n620_,
    new_n621_, new_n622_, new_n623_, new_n624_, new_n625_, new_n626_,
    new_n627_, new_n628_, new_n629_, new_n630_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n794_, new_n796_, new_n797_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n841_, new_n842_,
    new_n843_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n964_, new_n965_, new_n966_, new_n967_, new_n968_, new_n969_,
    new_n970_, new_n971_, new_n972_, new_n973_, new_n974_, new_n975_,
    new_n976_, new_n977_, new_n978_, new_n979_, new_n980_, new_n981_,
    new_n982_, new_n983_, new_n984_, new_n985_, new_n986_, new_n987_,
    new_n988_, new_n989_, new_n990_, new_n991_, new_n992_, new_n993_,
    new_n994_, new_n995_, new_n996_, new_n997_, new_n998_, new_n999_,
    new_n1000_, new_n1001_, new_n1002_, new_n1003_, new_n1004_, new_n1005_,
    new_n1006_, new_n1007_, new_n1008_, new_n1009_, new_n1010_, new_n1011_,
    new_n1012_, new_n1013_, new_n1014_, new_n1015_, new_n1016_, new_n1017_,
    new_n1018_, new_n1019_, new_n1020_, new_n1021_, new_n1022_, new_n1023_,
    new_n1024_, new_n1025_, new_n1026_, new_n1027_, new_n1028_, new_n1029_,
    new_n1030_, new_n1031_, new_n1032_, new_n1033_, new_n1034_, new_n1035_,
    new_n1036_, new_n1037_, new_n1038_, new_n1039_, new_n1040_, new_n1041_,
    new_n1042_, new_n1043_, new_n1044_, new_n1045_, new_n1046_, new_n1047_,
    new_n1048_, new_n1049_, new_n1050_, new_n1051_, new_n1052_, new_n1053_,
    new_n1054_, new_n1055_, new_n1056_, new_n1057_, new_n1058_, new_n1059_,
    new_n1060_, new_n1061_, new_n1062_, new_n1063_, new_n1064_, new_n1065_,
    new_n1066_, new_n1067_, new_n1068_, new_n1069_, new_n1070_, new_n1071_,
    new_n1072_, new_n1073_, new_n1074_, new_n1075_, new_n1076_, new_n1077_,
    new_n1078_, new_n1079_, new_n1080_, new_n1081_, new_n1082_, new_n1083_,
    new_n1084_, new_n1085_, new_n1086_, new_n1087_, new_n1088_, new_n1089_,
    new_n1090_, new_n1091_, new_n1092_, new_n1093_, new_n1094_, new_n1095_,
    new_n1096_, new_n1097_, new_n1098_, new_n1099_, new_n1100_, new_n1101_,
    new_n1102_, new_n1103_, new_n1104_, new_n1105_, new_n1106_, new_n1107_,
    new_n1108_, new_n1109_, new_n1110_, new_n1111_, new_n1112_, new_n1113_,
    new_n1114_, new_n1115_, new_n1116_, new_n1117_, new_n1118_, new_n1119_,
    new_n1120_, new_n1121_, new_n1122_, new_n1123_, new_n1124_, new_n1125_,
    new_n1126_, new_n1127_, new_n1128_, new_n1129_, new_n1130_, new_n1131_,
    new_n1132_, new_n1133_, new_n1134_, new_n1135_, new_n1136_, new_n1137_,
    new_n1138_, new_n1139_, new_n1140_, new_n1141_, new_n1142_, new_n1143_,
    new_n1144_, new_n1145_, new_n1146_, new_n1147_, new_n1148_, new_n1149_,
    new_n1150_, new_n1151_, new_n1152_, new_n1153_, new_n1154_, new_n1155_,
    new_n1156_, new_n1157_, new_n1158_, new_n1159_, new_n1160_, new_n1161_,
    new_n1162_, new_n1163_, new_n1164_, new_n1165_, new_n1166_, new_n1167_,
    new_n1168_, new_n1169_, new_n1170_, new_n1171_, new_n1172_, new_n1173_,
    new_n1174_, new_n1175_, new_n1176_, new_n1177_, new_n1178_, new_n1179_,
    new_n1180_, new_n1181_, new_n1182_, new_n1183_, new_n1184_, new_n1185_,
    new_n1186_, new_n1187_, new_n1188_, new_n1189_, new_n1190_, new_n1191_,
    new_n1192_, new_n1193_, new_n1194_, new_n1195_, new_n1196_, new_n1197_,
    new_n1198_, new_n1199_, new_n1200_, new_n1201_, new_n1202_, new_n1203_,
    new_n1204_, new_n1205_, new_n1206_, new_n1207_, new_n1208_, new_n1209_,
    new_n1210_, new_n1211_, new_n1212_, new_n1213_, new_n1214_, new_n1215_,
    new_n1216_, new_n1217_, new_n1219_, new_n1220_, new_n1221_, new_n1222_,
    new_n1223_, new_n1224_, new_n1225_, new_n1226_, new_n1227_, new_n1228_,
    new_n1229_, new_n1230_, new_n1231_, new_n1232_, new_n1233_, new_n1234_,
    new_n1235_, new_n1236_, new_n1237_, new_n1238_, new_n1239_, new_n1240_,
    new_n1241_, new_n1242_, new_n1243_, new_n1244_, new_n1245_, new_n1246_,
    new_n1247_, new_n1248_, new_n1249_, new_n1250_, new_n1251_, new_n1252_,
    new_n1253_, new_n1255_, new_n1256_, new_n1257_, new_n1258_, new_n1259_,
    new_n1260_, new_n1261_, new_n1262_, new_n1263_, new_n1264_, new_n1266_,
    new_n1267_, new_n1268_, new_n1269_, new_n1270_, new_n1271_, new_n1272_,
    new_n1273_, new_n1274_, new_n1275_, new_n1276_, new_n1277_, new_n1278_,
    new_n1279_, new_n1280_, new_n1281_, new_n1282_, new_n1283_, new_n1284_,
    new_n1285_, new_n1287_, new_n1288_, new_n1289_, new_n1290_, new_n1291_,
    new_n1292_, new_n1293_, new_n1294_, new_n1295_, new_n1296_, new_n1297_,
    new_n1298_, new_n1299_, new_n1300_, new_n1301_, new_n1302_, new_n1304_,
    new_n1305_, new_n1306_, new_n1310_, new_n1311_, new_n1312_, new_n1313_,
    new_n1314_, new_n1315_, new_n1317_, new_n1318_, new_n1320_, new_n1321_,
    new_n1322_, new_n1323_, new_n1324_, new_n1325_, new_n1326_, new_n1327_,
    new_n1328_, new_n1329_, new_n1330_, new_n1331_, new_n1332_, new_n1333_,
    new_n1334_, new_n1335_, new_n1336_, new_n1337_, new_n1338_, new_n1339_,
    new_n1340_, new_n1341_, new_n1342_, new_n1343_, new_n1344_, new_n1345_,
    new_n1346_, new_n1347_, new_n1348_, new_n1349_, new_n1350_, new_n1351_,
    new_n1352_, new_n1353_, new_n1354_, new_n1355_, new_n1356_, new_n1357_,
    new_n1358_, new_n1359_, new_n1360_, new_n1361_, new_n1362_, new_n1363_,
    new_n1364_, new_n1365_, new_n1366_, new_n1367_, new_n1368_, new_n1369_,
    new_n1370_, new_n1371_, new_n1372_, new_n1373_, new_n1374_, new_n1375_,
    new_n1376_, new_n1377_, new_n1378_, new_n1379_, new_n1380_, new_n1382_,
    new_n1383_, new_n1385_, new_n1386_, new_n1387_, new_n1388_, new_n1389_,
    new_n1391_, new_n1392_, new_n1393_, new_n1394_, new_n1395_, new_n1396_,
    new_n1397_, new_n1398_, new_n1399_, new_n1400_, new_n1402_, new_n1403_,
    new_n1404_, new_n1406_, new_n1407_, new_n1408_, new_n1409_, new_n1410_,
    new_n1411_, new_n1412_, new_n1413_, new_n1414_, new_n1415_, new_n1416_,
    new_n1417_, new_n1418_, new_n1419_, new_n1420_, new_n1421_, new_n1422_,
    new_n1423_, new_n1424_, new_n1425_, new_n1426_, new_n1427_, new_n1428_,
    new_n1429_, new_n1430_, new_n1431_, new_n1432_, new_n1434_, new_n1435_,
    new_n1436_, new_n1437_, new_n1438_, new_n1439_, new_n1440_, new_n1442_,
    new_n1443_, new_n1444_, new_n1445_, new_n1446_, new_n1447_, new_n1448_,
    new_n1449_, new_n1450_, new_n1451_, new_n1452_, new_n1453_, new_n1454_,
    new_n1455_, new_n1456_, new_n1457_, new_n1458_, new_n1459_, new_n1460_,
    new_n1461_, new_n1462_, new_n1463_, new_n1464_, new_n1465_, new_n1466_,
    new_n1468_, new_n1469_, new_n1470_, new_n1471_, new_n1472_, new_n1473_,
    new_n1475_, new_n1476_, new_n1477_, new_n1478_, new_n1480_, new_n1481_,
    new_n1482_, new_n1483_, new_n1484_, new_n1486_, new_n1487_, new_n1488_,
    new_n1489_, new_n1490_, new_n1491_, new_n1492_, new_n1494_, new_n1495_,
    new_n1497_, new_n1498_, new_n1500_, new_n1501_, new_n1502_, new_n1503_,
    new_n1504_, new_n1506_, new_n1507_, new_n1508_, new_n1509_, new_n1510_,
    new_n1511_, new_n1512_, new_n1514_, new_n1515_, new_n1516_, new_n1519_,
    new_n1520_, new_n1521_, new_n1522_, new_n1523_, new_n1524_, new_n1526_,
    new_n1527_, new_n1528_, new_n1529_, new_n1531_, new_n1532_, new_n1533_,
    new_n1534_, new_n1535_, new_n1536_, new_n1537_, new_n1539_, new_n1540_,
    new_n1541_, new_n1542_, new_n1544_, new_n1545_, new_n1546_, new_n1547_,
    new_n1548_, new_n1549_, new_n1550_, new_n1552_, new_n1553_, new_n1554_,
    new_n1555_, new_n1556_, new_n1557_, new_n1558_, new_n1559_, new_n1560_,
    new_n1561_, new_n1562_, new_n1563_, new_n1564_, new_n1566_, new_n1567_,
    new_n1569_, new_n1570_, new_n1571_, new_n1572_, new_n1574_, new_n1575_,
    new_n1576_, new_n1577_, new_n1578_, new_n1579_, new_n1581_, new_n1582_,
    new_n1583_, new_n1584_, new_n1585_, new_n1586_, new_n1587_, new_n1589_,
    new_n1590_, new_n1591_, new_n1592_, new_n1593_, new_n1594_, new_n1595_,
    new_n1597_, new_n1598_, new_n1599_, new_n1600_, new_n1601_, new_n1602_,
    new_n1603_, new_n1605_, new_n1607_, new_n1608_, new_n1609_, new_n1610_,
    new_n1612_, new_n1613_, new_n1614_, new_n1615_, new_n1616_, new_n1617_,
    new_n1619_, new_n1620_, new_n1621_, new_n1622_, new_n1623_, new_n1624_,
    new_n1625_, new_n1626_, new_n1627_, new_n1628_, new_n1629_, new_n1630_,
    new_n1631_, new_n1632_, new_n1633_, new_n1634_, new_n1635_, new_n1636_,
    new_n1637_, new_n1638_, new_n1639_, new_n1640_, new_n1641_, new_n1642_,
    new_n1643_, new_n1644_, new_n1646_, new_n1647_, new_n1648_, new_n1649_,
    new_n1650_, new_n1651_, new_n1652_, new_n1653_, new_n1654_, new_n1655_,
    new_n1656_, new_n1657_, new_n1658_, new_n1659_, new_n1660_, new_n1661_,
    new_n1662_, new_n1663_, new_n1664_, new_n1665_, new_n1666_, new_n1667_,
    new_n1668_, new_n1669_, new_n1670_, new_n1671_, new_n1672_, new_n1673_,
    new_n1674_, new_n1676_, new_n1677_, new_n1678_, new_n1679_, new_n1680_,
    new_n1681_, new_n1682_, new_n1683_, new_n1685_, new_n1686_, new_n1688_,
    new_n1689_, new_n1690_, new_n1691_, new_n1693_, new_n1694_, new_n1696_,
    new_n1697_, new_n1698_, new_n1699_, new_n1700_, new_n1701_, new_n1702_,
    new_n1703_, new_n1704_, new_n1705_, new_n1706_, new_n1707_, new_n1708_,
    new_n1709_, new_n1710_, new_n1711_, new_n1712_, new_n1713_, new_n1714_,
    new_n1715_, new_n1716_, new_n1717_, new_n1718_, new_n1719_, new_n1720_,
    new_n1721_, new_n1724_, new_n1725_, new_n1726_, new_n1727_, new_n1728_,
    new_n1729_, new_n1730_, new_n1731_, new_n1733_, new_n1734_, new_n1736_,
    new_n1738_, new_n1739_, new_n1740_, new_n1742_, new_n1743_, new_n1744_,
    new_n1745_, new_n1746_, new_n1747_, new_n1748_, new_n1750_, new_n1751_,
    new_n1752_, new_n1753_, new_n1754_, new_n1755_, new_n1756_, new_n1760_,
    new_n1761_, new_n1762_, new_n1763_, new_n1764_, new_n1765_, new_n1766_,
    new_n1767_, new_n1768_, new_n1769_, new_n1770_, new_n1771_, new_n1772_,
    new_n1773_, new_n1774_, new_n1775_, new_n1776_, new_n1777_, new_n1778_,
    new_n1779_, new_n1780_, new_n1781_, new_n1782_, new_n1783_, new_n1785_,
    new_n1786_, new_n1787_, new_n1788_, new_n1789_, new_n1791_, new_n1792_,
    new_n1793_, new_n1795_, new_n1796_, new_n1797_, new_n1798_, new_n1799_,
    new_n1800_, new_n1802_, new_n1803_, new_n1804_, new_n1805_, new_n1806_,
    new_n1807_, new_n1808_, new_n1810_, new_n1811_, new_n1812_, new_n1813_,
    new_n1814_, new_n1815_, new_n1817_, new_n1818_, new_n1819_, new_n1820_,
    new_n1821_, new_n1822_, new_n1823_, new_n1825_, new_n1826_, new_n1827_,
    new_n1828_, new_n1829_, new_n1830_, new_n1832_, new_n1833_, new_n1834_,
    new_n1835_, new_n1836_, new_n1837_, new_n1838_, new_n1840_, new_n1841_,
    new_n1842_, new_n1843_, new_n1844_, new_n1845_, new_n1846_, new_n1848_,
    new_n1849_, new_n1850_, new_n1851_, new_n1852_, new_n1853_, new_n1855_,
    new_n1856_, new_n1857_, new_n1859_, new_n1860_, new_n1861_, new_n1862_,
    new_n1863_, new_n1864_, new_n1866_, new_n1867_, new_n1868_, new_n1869_,
    new_n1870_, new_n1871_, new_n1873_, new_n1874_, new_n1875_, new_n1876_,
    new_n1877_, new_n1878_, new_n1879_, new_n1881_, new_n1882_, new_n1883_,
    new_n1884_, new_n1885_, new_n1886_, new_n1889_, new_n1890_, new_n1891_,
    new_n1892_, new_n1893_, new_n1894_, new_n1895_, new_n1897_, new_n1898_,
    new_n1899_, new_n1900_, new_n1901_, new_n1902_, new_n1904_, new_n1905_,
    new_n1906_, new_n1909_, new_n1910_, new_n1911_, new_n1912_, new_n1913_,
    new_n1914_, new_n1916_, new_n1917_, new_n1918_, new_n1919_, new_n1920_,
    new_n1921_, new_n1922_, new_n1925_, new_n1926_, new_n1927_, new_n1928_,
    new_n1929_, new_n1930_, new_n1932_, new_n1933_, new_n1934_, new_n1935_,
    new_n1936_, new_n1937_, new_n1938_, new_n1939_, new_n1940_, new_n1941_,
    new_n1942_, new_n1943_, new_n1944_, new_n1945_, new_n1946_, new_n1947_,
    new_n1948_, new_n1949_, new_n1950_, new_n1951_, new_n1952_, new_n1953_,
    new_n1954_, new_n1955_, new_n1956_, new_n1957_, new_n1958_, new_n1959_,
    new_n1960_, new_n1961_, new_n1962_, new_n1963_, new_n1964_, new_n1965_,
    new_n1966_, new_n1967_, new_n1968_, new_n1969_, new_n1970_, new_n1971_,
    new_n1972_, new_n1973_, new_n1974_, new_n1975_, new_n1976_, new_n1977_,
    new_n1978_, new_n1979_, new_n1980_, new_n1981_, new_n1982_, new_n1983_,
    new_n1984_, new_n1985_, new_n1986_, new_n1987_, new_n1988_, new_n1989_,
    new_n1990_, new_n1991_, new_n1992_, new_n1993_, new_n1994_, new_n1995_,
    new_n1996_, new_n1997_, new_n1998_, new_n1999_, new_n2000_, new_n2001_,
    new_n2002_, new_n2003_, new_n2004_, new_n2005_, new_n2006_, new_n2007_,
    new_n2008_, new_n2009_, new_n2010_, new_n2011_, new_n2012_, new_n2013_,
    new_n2014_, new_n2015_, new_n2016_, new_n2017_, new_n2018_, new_n2019_,
    new_n2020_, new_n2021_, new_n2022_, new_n2024_, new_n2025_, new_n2026_,
    new_n2028_, new_n2029_, new_n2030_, new_n2031_, new_n2032_, new_n2033_,
    new_n2034_, new_n2035_, new_n2036_, new_n2037_, new_n2038_, new_n2039_,
    new_n2040_, new_n2041_, new_n2042_, new_n2043_, new_n2044_, new_n2045_,
    new_n2046_, new_n2047_, new_n2048_, new_n2049_, new_n2050_, new_n2051_,
    new_n2052_, new_n2053_, new_n2054_, new_n2055_, new_n2056_, new_n2057_,
    new_n2058_, new_n2059_, new_n2060_, new_n2061_, new_n2062_, new_n2063_,
    new_n2064_, new_n2065_, new_n2066_, new_n2067_, new_n2068_, new_n2069_,
    new_n2070_, new_n2071_, new_n2072_, new_n2073_, new_n2074_, new_n2075_,
    new_n2076_, new_n2077_, new_n2078_, new_n2079_, new_n2080_, new_n2081_,
    new_n2082_, new_n2083_, new_n2084_, new_n2085_, new_n2086_, new_n2087_,
    new_n2088_, new_n2089_, new_n2090_, new_n2091_, new_n2092_, new_n2093_,
    new_n2094_, new_n2095_, new_n2096_, new_n2097_, new_n2098_, new_n2099_,
    new_n2100_, new_n2101_, new_n2102_, new_n2103_, new_n2104_, new_n2105_,
    new_n2106_, new_n2107_, new_n2108_, new_n2109_, new_n2110_, new_n2111_,
    new_n2112_, new_n2113_, new_n2114_, new_n2115_, new_n2116_, new_n2117_,
    new_n2118_, new_n2119_, new_n2120_, new_n2121_, new_n2122_, new_n2123_,
    new_n2124_, new_n2125_, new_n2126_, new_n2127_, new_n2128_, new_n2129_,
    new_n2130_, new_n2131_, new_n2132_, new_n2133_, new_n2134_, new_n2135_,
    new_n2136_, new_n2137_, new_n2138_, new_n2139_, new_n2140_, new_n2142_,
    new_n2143_, new_n2144_, new_n2147_, new_n2148_, new_n2149_, new_n2150_,
    new_n2151_, new_n2152_, new_n2153_, new_n2154_, new_n2155_, new_n2156_,
    new_n2157_, new_n2158_, new_n2159_, new_n2160_, new_n2161_, new_n2162_,
    new_n2163_, new_n2164_, new_n2165_, new_n2166_, new_n2167_, new_n2168_,
    new_n2169_, new_n2170_, new_n2171_, new_n2173_, new_n2174_, new_n2175_,
    new_n2176_, new_n2177_, new_n2178_, new_n2179_, new_n2180_, new_n2181_,
    new_n2182_, new_n2183_, new_n2184_, new_n2185_, new_n2186_, new_n2187_,
    new_n2188_, new_n2189_, new_n2190_, new_n2191_, new_n2192_, new_n2193_,
    new_n2194_, new_n2195_, new_n2197_, new_n2198_, new_n2199_, new_n2200_,
    new_n2202_, new_n2203_, new_n2204_, new_n2205_, new_n2206_, new_n2207_,
    new_n2208_, new_n2209_, new_n2210_, new_n2211_, new_n2212_, new_n2213_,
    new_n2214_, new_n2215_, new_n2216_, new_n2217_, new_n2218_, new_n2219_,
    new_n2220_, new_n2221_, new_n2222_, new_n2223_, new_n2224_, new_n2225_,
    new_n2226_, new_n2227_, new_n2228_, new_n2229_, new_n2230_, new_n2231_,
    new_n2232_, new_n2233_, new_n2234_, new_n2235_, new_n2236_, new_n2237_,
    new_n2238_, new_n2239_, new_n2240_, new_n2241_, new_n2242_, new_n2243_,
    new_n2244_, new_n2245_, new_n2246_, new_n2247_, new_n2248_, new_n2249_,
    new_n2250_, new_n2251_, new_n2252_, new_n2253_, new_n2254_, new_n2255_,
    new_n2256_, new_n2257_, new_n2258_, new_n2259_, new_n2260_, new_n2261_,
    new_n2262_, new_n2263_, new_n2264_, new_n2265_, new_n2266_, new_n2267_,
    new_n2268_, new_n2269_, new_n2270_, new_n2271_, new_n2272_, new_n2273_,
    new_n2274_, new_n2275_, new_n2276_, new_n2277_, new_n2278_, new_n2279_,
    new_n2280_, new_n2281_, new_n2282_, new_n2283_, new_n2284_, new_n2285_,
    new_n2286_, new_n2287_, new_n2288_, new_n2289_, new_n2290_, new_n2291_,
    new_n2292_, new_n2293_, new_n2294_, new_n2295_, new_n2296_, new_n2297_,
    new_n2298_, new_n2299_, new_n2300_, new_n2301_, new_n2302_, new_n2303_,
    new_n2304_, new_n2305_, new_n2306_, new_n2307_, new_n2308_, new_n2309_,
    new_n2310_, new_n2311_, new_n2312_, new_n2313_, new_n2314_, new_n2315_,
    new_n2316_, new_n2317_, new_n2318_, new_n2319_, new_n2320_, new_n2321_,
    new_n2322_, new_n2323_, new_n2324_, new_n2325_, new_n2326_, new_n2327_,
    new_n2328_, new_n2329_, new_n2330_, new_n2331_, new_n2332_, new_n2333_,
    new_n2334_, new_n2335_, new_n2336_, new_n2337_, new_n2338_, new_n2339_,
    new_n2340_, new_n2341_, new_n2342_, new_n2343_, new_n2344_, new_n2345_,
    new_n2346_, new_n2347_, new_n2348_, new_n2349_, new_n2350_, new_n2351_,
    new_n2352_, new_n2353_, new_n2354_, new_n2355_, new_n2356_, new_n2357_,
    new_n2358_, new_n2359_, new_n2360_, new_n2361_, new_n2362_, new_n2363_,
    new_n2364_, new_n2365_, new_n2366_, new_n2367_, new_n2368_, new_n2369_,
    new_n2370_, new_n2371_, new_n2372_, new_n2373_, new_n2374_, new_n2375_,
    new_n2376_, new_n2377_, new_n2378_, new_n2379_, new_n2380_, new_n2381_,
    new_n2382_, new_n2383_, new_n2384_, new_n2385_, new_n2386_, new_n2387_,
    new_n2388_, new_n2389_, new_n2390_, new_n2391_, new_n2392_, new_n2393_,
    new_n2394_, new_n2395_, new_n2396_, new_n2397_, new_n2398_, new_n2399_,
    new_n2400_, new_n2401_, new_n2402_, new_n2403_, new_n2404_, new_n2405_,
    new_n2406_, new_n2407_, new_n2408_, new_n2409_, new_n2410_, new_n2411_,
    new_n2412_, new_n2413_, new_n2414_, new_n2415_, new_n2416_, new_n2417_,
    new_n2418_, new_n2419_, new_n2420_, new_n2421_, new_n2422_, new_n2423_,
    new_n2424_, new_n2425_, new_n2426_, new_n2427_, new_n2428_, new_n2429_,
    new_n2430_, new_n2431_, new_n2432_, new_n2433_, new_n2434_, new_n2435_,
    new_n2436_, new_n2437_, new_n2438_, new_n2439_, new_n2440_, new_n2441_,
    new_n2442_, new_n2443_, new_n2444_, new_n2445_, new_n2446_, new_n2447_,
    new_n2448_, new_n2449_, new_n2450_, new_n2451_, new_n2452_, new_n2453_,
    new_n2454_, new_n2455_, new_n2456_, new_n2457_, new_n2458_, new_n2459_,
    new_n2460_, new_n2461_, new_n2462_, new_n2463_, new_n2464_, new_n2465_,
    new_n2466_, new_n2467_, new_n2468_, new_n2469_, new_n2470_, new_n2471_,
    new_n2472_, new_n2473_, new_n2474_, new_n2475_, new_n2476_, new_n2477_,
    new_n2478_, new_n2479_, new_n2480_, new_n2481_, new_n2482_, new_n2483_,
    new_n2484_, new_n2485_, new_n2486_, new_n2487_, new_n2488_, new_n2489_,
    new_n2490_, new_n2491_, new_n2492_, new_n2493_, new_n2494_, new_n2495_,
    new_n2496_, new_n2497_, new_n2498_, new_n2499_, new_n2500_, new_n2501_,
    new_n2502_, new_n2503_, new_n2504_, new_n2505_, new_n2506_, new_n2507_,
    new_n2508_, new_n2509_, new_n2510_, new_n2511_, new_n2512_, new_n2513_,
    new_n2514_, new_n2515_, new_n2516_, new_n2517_, new_n2518_, new_n2519_,
    new_n2520_, new_n2521_, new_n2522_, new_n2523_, new_n2524_, new_n2525_,
    new_n2526_, new_n2527_, new_n2528_, new_n2529_, new_n2530_, new_n2531_,
    new_n2532_, new_n2533_, new_n2534_, new_n2535_, new_n2536_, new_n2537_,
    new_n2538_, new_n2539_, new_n2540_, new_n2541_, new_n2542_, new_n2543_,
    new_n2544_, new_n2545_, new_n2546_, new_n2547_, new_n2548_, new_n2549_,
    new_n2550_, new_n2551_, new_n2552_, new_n2553_, new_n2554_, new_n2555_,
    new_n2556_, new_n2557_, new_n2558_, new_n2559_, new_n2560_, new_n2561_,
    new_n2562_, new_n2563_, new_n2564_, new_n2565_, new_n2566_, new_n2567_,
    new_n2568_, new_n2569_, new_n2570_, new_n2571_, new_n2572_, new_n2573_,
    new_n2574_, new_n2575_, new_n2576_, new_n2577_, new_n2578_, new_n2579_,
    new_n2580_, new_n2581_, new_n2582_, new_n2583_, new_n2584_, new_n2585_,
    new_n2586_, new_n2587_, new_n2588_, new_n2589_, new_n2590_, new_n2591_,
    new_n2592_, new_n2593_, new_n2594_, new_n2595_, new_n2596_, new_n2597_,
    new_n2598_, new_n2599_, new_n2600_, new_n2602_, new_n2603_, new_n2604_,
    new_n2605_, new_n2606_, new_n2607_, new_n2608_, new_n2609_, new_n2610_,
    new_n2611_, new_n2612_, new_n2613_, new_n2614_, new_n2615_, new_n2616_,
    new_n2617_, new_n2618_, new_n2619_, new_n2620_, new_n2621_, new_n2622_,
    new_n2623_, new_n2624_, new_n2625_, new_n2626_, new_n2627_, new_n2628_,
    new_n2629_, new_n2630_, new_n2631_, new_n2632_, new_n2633_, new_n2634_,
    new_n2635_, new_n2636_, new_n2637_, new_n2638_, new_n2639_, new_n2640_,
    new_n2641_, new_n2642_, new_n2643_, new_n2644_, new_n2645_, new_n2646_,
    new_n2647_, new_n2648_, new_n2649_, new_n2650_, new_n2651_, new_n2652_,
    new_n2653_, new_n2654_, new_n2655_, new_n2656_, new_n2657_, new_n2658_,
    new_n2659_, new_n2660_, new_n2661_, new_n2662_, new_n2663_, new_n2664_,
    new_n2665_, new_n2666_, new_n2667_, new_n2668_, new_n2669_, new_n2670_,
    new_n2671_, new_n2673_, new_n2674_, new_n2675_, new_n2676_, new_n2677_,
    new_n2678_, new_n2679_, new_n2680_, new_n2681_, new_n2682_, new_n2683_,
    new_n2684_, new_n2685_, new_n2686_, new_n2687_, new_n2689_, new_n2690_,
    new_n2691_, new_n2692_, new_n2693_, new_n2694_, new_n2695_, new_n2696_,
    new_n2697_, new_n2698_, new_n2699_, new_n2700_, new_n2701_, new_n2702_,
    new_n2703_, new_n2704_, new_n2705_, new_n2706_, new_n2707_, new_n2708_,
    new_n2709_, new_n2711_, new_n2712_, new_n2713_, new_n2714_, new_n2715_,
    new_n2716_, new_n2717_, new_n2718_, new_n2719_, new_n2720_, new_n2721_,
    new_n2722_, new_n2723_, new_n2724_, new_n2725_, new_n2727_, new_n2728_,
    new_n2729_, new_n2731_, new_n2732_, new_n2733_, new_n2734_, new_n2735_,
    new_n2736_, new_n2737_, new_n2738_, new_n2739_, new_n2740_, new_n2741_,
    new_n2745_, new_n2746_, new_n2747_, new_n2748_, new_n2749_, new_n2750_,
    new_n2751_, new_n2752_, new_n2753_, new_n2754_, new_n2755_, new_n2756_,
    new_n2757_, new_n2758_, new_n2759_, new_n2760_, new_n2761_, new_n2762_,
    new_n2763_, new_n2764_, new_n2766_, new_n2767_, new_n2768_, new_n2769_,
    new_n2770_, new_n2771_, new_n2772_, new_n2773_, new_n2774_, new_n2775_,
    new_n2776_, new_n2777_, new_n2778_, new_n2779_, new_n2780_, new_n2781_,
    new_n2782_, new_n2784_, new_n2785_, new_n2786_, new_n2787_, new_n2789_,
    new_n2790_, new_n2791_, new_n2792_, new_n2793_, new_n2794_, new_n2795_,
    new_n2796_, new_n2797_, new_n2798_, new_n2799_, new_n2800_, new_n2801_,
    new_n2802_, new_n2803_, new_n2804_, new_n2805_, new_n2807_, new_n2808_,
    new_n2809_, new_n2810_, new_n2811_, new_n2812_, new_n2813_, new_n2814_,
    new_n2815_, new_n2816_, new_n2817_, new_n2818_, new_n2819_, new_n2820_,
    new_n2821_, new_n2823_, new_n2824_, new_n2825_, new_n2826_, new_n2827_,
    new_n2828_, new_n2829_, new_n2830_, new_n2831_, new_n2832_, new_n2833_,
    new_n2834_, new_n2835_, new_n2836_, new_n2837_, new_n2838_, new_n2839_,
    new_n2840_, new_n2841_, new_n2842_, new_n2843_, new_n2844_, new_n2845_,
    new_n2846_, new_n2847_, new_n2849_, new_n2850_, new_n2851_, new_n2852_,
    new_n2853_, new_n2854_, new_n2856_, new_n2857_, new_n2858_, new_n2859_,
    new_n2860_, new_n2861_, new_n2862_, new_n2863_, new_n2864_, new_n2865_,
    new_n2866_, new_n2867_, new_n2868_, new_n2869_, new_n2871_, new_n2872_,
    new_n2873_, new_n2874_, new_n2875_, new_n2876_, new_n2877_, new_n2878_,
    new_n2879_, new_n2881_, new_n2882_, new_n2883_, new_n2885_, new_n2886_,
    new_n2888_, new_n2889_, new_n2890_, new_n2891_, new_n2892_, new_n2893_,
    new_n2894_, new_n2895_, new_n2896_, new_n2897_, new_n2898_, new_n2900_,
    new_n2901_, new_n2902_, new_n2903_, new_n2904_, new_n2905_, new_n2906_,
    new_n2907_, new_n2908_, new_n2909_, new_n2910_, new_n2911_, new_n2912_,
    new_n2913_, new_n2914_, new_n2915_, new_n2916_, new_n2917_, new_n2918_,
    new_n2919_, new_n2920_, new_n2921_, new_n2922_, new_n2923_, new_n2924_,
    new_n2925_, new_n2927_, new_n2928_, new_n2929_, new_n2930_, new_n2931_,
    new_n2932_, new_n2933_, new_n2934_, new_n2935_, new_n2937_, new_n2938_,
    new_n2939_, new_n2941_, new_n2942_, new_n2943_, new_n2944_, new_n2945_,
    new_n2946_, new_n2947_, new_n2948_, new_n2949_, new_n2950_, new_n2953_,
    new_n2954_, new_n2955_, new_n2956_, new_n2957_, new_n2958_, new_n2959_,
    new_n2961_, new_n2962_, new_n2963_, new_n2964_, new_n2965_, new_n2966_,
    new_n2967_, new_n2968_, new_n2969_, new_n2970_, new_n2971_, new_n2974_,
    new_n2975_, new_n2976_, new_n2977_, new_n2978_, new_n2979_, new_n2980_,
    new_n2981_, new_n2982_, new_n2983_, new_n2985_, new_n2986_, new_n2987_,
    new_n2988_, new_n2989_, new_n2990_, new_n2991_, new_n2992_, new_n2993_,
    new_n2994_, new_n2995_, new_n2996_, new_n2997_, new_n2998_, new_n2999_,
    new_n3000_, new_n3001_, new_n3002_, new_n3003_, new_n3004_, new_n3005_,
    new_n3006_, new_n3007_, new_n3009_, new_n3010_, new_n3011_, new_n3012_,
    new_n3013_, new_n3014_, new_n3015_, new_n3016_, new_n3017_, new_n3018_,
    new_n3019_, new_n3020_, new_n3021_, new_n3022_, new_n3023_, new_n3025_,
    new_n3026_, new_n3027_, new_n3028_, new_n3029_, new_n3030_, new_n3031_,
    new_n3032_, new_n3033_, new_n3035_, new_n3036_, new_n3037_, new_n3039_,
    new_n3040_, new_n3041_, new_n3042_, new_n3043_, new_n3044_, new_n3045_,
    new_n3046_, new_n3047_, new_n3048_, new_n3049_, new_n3052_, new_n3053_,
    new_n3054_, new_n3055_, new_n3056_, new_n3057_, new_n3058_, new_n3059_,
    new_n3060_, new_n3061_, new_n3062_, new_n3063_, new_n3064_, new_n3065_,
    new_n3066_, new_n3067_, new_n3068_, new_n3069_, new_n3070_, new_n3071_,
    new_n3072_, new_n3074_, new_n3075_, new_n3076_, new_n3077_, new_n3078_,
    new_n3079_, new_n3081_, new_n3082_, new_n3083_, new_n3084_, new_n3085_,
    new_n3086_, new_n3087_, new_n3089_, new_n3091_, new_n3092_, new_n3093_,
    new_n3094_, new_n3095_, new_n3096_, new_n3097_, new_n3099_, new_n3100_,
    new_n3102_, new_n3103_, new_n3104_, new_n3105_, new_n3106_, new_n3107_,
    new_n3108_, new_n3109_, new_n3110_, new_n3111_, new_n3112_, new_n3114_,
    new_n3115_, new_n3116_, new_n3117_, new_n3118_, new_n3119_, new_n3120_,
    new_n3121_, new_n3122_, new_n3123_, new_n3126_, new_n3127_, new_n3128_,
    new_n3129_, new_n3130_, new_n3131_, new_n3132_, new_n3133_, new_n3134_,
    new_n3135_, new_n3136_, new_n3138_, new_n3139_, new_n3140_, new_n3141_,
    new_n3142_, new_n3143_, new_n3144_, new_n3145_, new_n3146_, new_n3147_,
    new_n3148_, new_n3150_, new_n3151_, new_n3152_, new_n3153_, new_n3154_,
    new_n3155_, new_n3156_, new_n3157_, new_n3158_, new_n3159_, new_n3161_,
    new_n3162_, new_n3163_, new_n3164_, new_n3165_, new_n3166_, new_n3167_,
    new_n3168_, new_n3169_, new_n3170_, new_n3172_, new_n3173_, new_n3174_,
    new_n3175_, new_n3176_, new_n3177_, new_n3178_, new_n3179_, new_n3180_,
    new_n3181_, new_n3182_, new_n3184_, new_n3185_, new_n3186_, new_n3187_,
    new_n3189_, new_n3190_, new_n3191_, new_n3192_, new_n3193_, new_n3194_,
    new_n3195_, new_n3196_, new_n3197_, new_n3198_, new_n3199_, new_n3201_,
    new_n3202_, new_n3203_, new_n3204_, new_n3205_, new_n3206_, new_n3207_,
    new_n3208_, new_n3209_, new_n3210_, new_n3211_, new_n3213_, new_n3214_,
    new_n3215_, new_n3216_, new_n3217_, new_n3218_, new_n3219_, new_n3220_,
    new_n3221_, new_n3222_, new_n3223_, new_n3224_, new_n3225_, new_n3226_,
    new_n3227_, new_n3228_, new_n3229_, new_n3230_, new_n3231_, new_n3232_,
    new_n3233_, new_n3234_, new_n3235_, new_n3236_, new_n3237_, new_n3238_,
    new_n3239_, new_n3241_, new_n3242_, new_n3243_, new_n3244_, new_n3245_,
    new_n3246_, new_n3247_, new_n3248_, new_n3249_, new_n3250_, new_n3251_,
    new_n3252_, new_n3253_, new_n3254_, new_n3255_, new_n3256_, new_n3257_,
    new_n3258_, new_n3259_, new_n3260_, new_n3261_, new_n3262_, new_n3263_,
    new_n3264_, new_n3265_, new_n3266_, new_n3267_, new_n3268_, new_n3269_,
    new_n3270_, new_n3271_, new_n3273_, new_n3274_, new_n3275_, new_n3276_,
    new_n3277_, new_n3278_, new_n3279_, new_n3280_, new_n3281_, new_n3282_,
    new_n3283_, new_n3284_, new_n3285_, new_n3286_, new_n3287_, new_n3288_,
    new_n3289_, new_n3290_, new_n3291_, new_n3292_, new_n3293_, new_n3294_,
    new_n3295_, new_n3296_, new_n3297_, new_n3298_, new_n3300_, new_n3301_,
    new_n3302_, new_n3303_, new_n3305_, new_n3306_, new_n3307_, new_n3308_,
    new_n3309_, new_n3310_, new_n3311_, new_n3312_, new_n3313_, new_n3314_,
    new_n3315_, new_n3317_, new_n3318_, new_n3319_, new_n3320_, new_n3321_,
    new_n3322_, new_n3323_, new_n3324_, new_n3325_, new_n3326_, new_n3327_,
    new_n3329_, new_n3330_, new_n3331_, new_n3332_, new_n3333_, new_n3335_,
    new_n3336_, new_n3337_, new_n3338_, new_n3340_, new_n3341_, new_n3342_,
    new_n3343_, new_n3344_, new_n3345_, new_n3346_, new_n3347_, new_n3348_,
    new_n3349_, new_n3351_, new_n3352_, new_n3353_, new_n3354_, new_n3355_,
    new_n3356_, new_n3357_, new_n3358_, new_n3359_, new_n3360_, new_n3362_,
    new_n3363_, new_n3364_, new_n3365_, new_n3366_, new_n3367_, new_n3368_,
    new_n3369_, new_n3370_, new_n3371_, new_n3373_, new_n3374_, new_n3375_,
    new_n3376_, new_n3378_, new_n3379_, new_n3380_, new_n3381_, new_n3382_,
    new_n3383_, new_n3384_, new_n3385_, new_n3386_, new_n3387_, new_n3388_,
    new_n3390_, new_n3391_, new_n3392_, new_n3393_, new_n3394_, new_n3395_,
    new_n3396_, new_n3397_, new_n3398_, new_n3399_, new_n3400_, new_n3403_,
    new_n3404_, new_n3405_, new_n3406_, new_n3407_, new_n3408_, new_n3409_,
    new_n3410_, new_n3411_, new_n3412_, new_n3414_, new_n3415_, new_n3416_,
    new_n3418_, new_n3419_, new_n3420_, new_n3421_, new_n3422_, new_n3423_,
    new_n3424_, new_n3425_, new_n3426_, new_n3427_, new_n3429_, new_n3430_,
    new_n3431_, new_n3432_, new_n3434_, new_n3435_, new_n3436_, new_n3437_,
    new_n3438_, new_n3439_, new_n3440_, new_n3441_, new_n3442_, new_n3443_,
    new_n3446_, new_n3447_, new_n3448_, new_n3449_, new_n3450_, new_n3451_,
    new_n3452_, new_n3453_, new_n3454_, new_n3455_, new_n3457_, new_n3458_,
    new_n3459_, new_n3460_, new_n3461_, new_n3462_, new_n3463_, new_n3464_,
    new_n3465_, new_n3466_, new_n3467_, new_n3469_, new_n3470_, new_n3471_,
    new_n3472_, new_n3473_, new_n3474_, new_n3475_, new_n3476_, new_n3477_,
    new_n3478_, new_n3480_, new_n3481_, new_n3482_, new_n3483_, new_n3484_,
    new_n3485_, new_n3486_, new_n3487_, new_n3488_, new_n3489_, new_n3491_,
    new_n3492_, new_n3493_, new_n3494_, new_n3495_, new_n3496_, new_n3497_,
    new_n3498_, new_n3499_, new_n3500_, new_n3502_, new_n3503_, new_n3505_,
    new_n3506_, new_n3507_, new_n3508_, new_n3509_, new_n3510_, new_n3511_,
    new_n3512_, new_n3513_, new_n3514_, new_n3515_, new_n3517_, new_n3518_,
    new_n3519_, new_n3521_, new_n3522_, new_n3523_, new_n3524_;
  assign new_n603_ = \1_n1551  & \1_n1655 ;
  assign new_n604_ = ~\1_n526  & new_n603_;
  assign new_n605_ = ~\1_n1551  & \1_n1655 ;
  assign new_n606_ = ~\1_n532  & \1_n1065 ;
  assign new_n607_ = \1_n1475  & new_n606_;
  assign new_n608_ = \1_n325  & \1_n677 ;
  assign new_n609_ = \1_n507  & ~\1_n677 ;
  assign new_n610_ = ~new_n608_ & ~new_n609_;
  assign new_n611_ = ~\1_n1240  & ~new_n610_;
  assign new_n612_ = ~\1_n677  & ~\1_n1311 ;
  assign new_n613_ = ~\1_n198  & \1_n677 ;
  assign new_n614_ = ~new_n612_ & ~new_n613_;
  assign new_n615_ = \1_n1240  & ~new_n614_;
  assign new_n616_ = ~new_n611_ & ~new_n615_;
  assign new_n617_ = ~\1_n532  & ~\1_n1065 ;
  assign new_n618_ = ~new_n616_ & new_n617_;
  assign new_n619_ = ~new_n607_ & ~new_n618_;
  assign new_n620_ = \1_n373  & \1_n1243 ;
  assign new_n621_ = \1_n677  & ~\1_n1243 ;
  assign new_n622_ = ~new_n620_ & ~new_n621_;
  assign new_n623_ = \1_n1240  & new_n622_;
  assign new_n624_ = ~\1_n1240  & ~new_n622_;
  assign new_n625_ = ~new_n623_ & ~new_n624_;
  assign new_n626_ = \1_n137  & \1_n1243 ;
  assign new_n627_ = \1_n859  & ~\1_n1243 ;
  assign new_n628_ = ~new_n626_ & ~new_n627_;
  assign new_n629_ = \1_n184  & new_n628_;
  assign new_n630_ = ~\1_n184  & ~new_n628_;
  assign new_n631_ = ~new_n629_ & ~new_n630_;
  assign new_n632_ = \1_n1243  & \1_n1331 ;
  assign new_n633_ = \1_n824  & ~\1_n1243 ;
  assign new_n634_ = ~new_n632_ & ~new_n633_;
  assign new_n635_ = \1_n1530  & ~new_n634_;
  assign new_n636_ = \1_n737  & \1_n1243 ;
  assign new_n637_ = \1_n135  & ~\1_n1243 ;
  assign new_n638_ = ~new_n636_ & ~new_n637_;
  assign new_n639_ = \1_n765  & ~new_n638_;
  assign new_n640_ = \1_n1530  & new_n634_;
  assign new_n641_ = ~\1_n1530  & ~new_n634_;
  assign new_n642_ = ~new_n640_ & ~new_n641_;
  assign new_n643_ = new_n639_ & ~new_n642_;
  assign new_n644_ = ~new_n635_ & ~new_n643_;
  assign new_n645_ = ~new_n631_ & ~new_n644_;
  assign new_n646_ = \1_n184  & ~new_n628_;
  assign new_n647_ = ~new_n645_ & ~new_n646_;
  assign new_n648_ = \1_n765  & new_n638_;
  assign new_n649_ = ~\1_n765  & ~new_n638_;
  assign new_n650_ = ~new_n648_ & ~new_n649_;
  assign new_n651_ = ~new_n642_ & ~new_n650_;
  assign new_n652_ = ~new_n631_ & new_n651_;
  assign new_n653_ = new_n647_ & ~new_n652_;
  assign new_n654_ = \1_n579  & \1_n1243 ;
  assign new_n655_ = \1_n1143  & ~\1_n1243 ;
  assign new_n656_ = ~new_n654_ & ~new_n655_;
  assign new_n657_ = \1_n1108  & new_n656_;
  assign new_n658_ = ~\1_n1108  & ~new_n656_;
  assign new_n659_ = ~new_n657_ & ~new_n658_;
  assign new_n660_ = \1_n1243  & \1_n1407 ;
  assign new_n661_ = \1_n956  & ~\1_n1243 ;
  assign new_n662_ = ~new_n660_ & ~new_n661_;
  assign new_n663_ = \1_n1479  & ~new_n662_;
  assign new_n664_ = \1_n1479  & new_n662_;
  assign new_n665_ = ~\1_n1479  & ~new_n662_;
  assign new_n666_ = ~new_n664_ & ~new_n665_;
  assign new_n667_ = \1_n69  & \1_n1243 ;
  assign new_n668_ = ~\1_n1243  & \1_n1251 ;
  assign new_n669_ = ~new_n667_ & ~new_n668_;
  assign new_n670_ = \1_n147  & ~new_n669_;
  assign new_n671_ = \1_n356  & \1_n1243 ;
  assign new_n672_ = \1_n1030  & ~\1_n1243 ;
  assign new_n673_ = ~new_n671_ & ~new_n672_;
  assign new_n674_ = \1_n938  & ~new_n673_;
  assign new_n675_ = \1_n107  & \1_n1243 ;
  assign new_n676_ = \1_n209  & ~\1_n1243 ;
  assign new_n677_ = ~new_n675_ & ~new_n676_;
  assign new_n678_ = \1_n950  & ~new_n677_;
  assign new_n679_ = \1_n938  & new_n673_;
  assign new_n680_ = ~\1_n938  & ~new_n673_;
  assign new_n681_ = ~new_n679_ & ~new_n680_;
  assign new_n682_ = new_n678_ & ~new_n681_;
  assign new_n683_ = ~new_n674_ & ~new_n682_;
  assign new_n684_ = \1_n147  & new_n669_;
  assign new_n685_ = ~\1_n147  & ~new_n669_;
  assign new_n686_ = ~new_n684_ & ~new_n685_;
  assign new_n687_ = ~new_n683_ & ~new_n686_;
  assign new_n688_ = ~new_n670_ & ~new_n687_;
  assign new_n689_ = ~new_n666_ & ~new_n688_;
  assign new_n690_ = ~new_n663_ & ~new_n689_;
  assign new_n691_ = ~new_n659_ & ~new_n690_;
  assign new_n692_ = \1_n1108  & ~new_n656_;
  assign new_n693_ = ~new_n691_ & ~new_n692_;
  assign new_n694_ = \1_n950  & new_n677_;
  assign new_n695_ = ~\1_n950  & ~new_n677_;
  assign new_n696_ = ~new_n694_ & ~new_n695_;
  assign new_n697_ = ~new_n681_ & ~new_n696_;
  assign new_n698_ = ~new_n686_ & new_n697_;
  assign new_n699_ = ~new_n666_ & new_n698_;
  assign new_n700_ = \1_n857  & new_n699_;
  assign new_n701_ = ~new_n659_ & new_n700_;
  assign new_n702_ = new_n693_ & ~new_n701_;
  assign new_n703_ = new_n647_ & new_n702_;
  assign new_n704_ = ~new_n653_ & ~new_n703_;
  assign new_n705_ = ~new_n625_ & new_n704_;
  assign new_n706_ = new_n625_ & ~new_n704_;
  assign new_n707_ = ~new_n705_ & ~new_n706_;
  assign new_n708_ = \1_n532  & ~\1_n1065 ;
  assign new_n709_ = new_n707_ & new_n708_;
  assign \1_n1645  = ~new_n619_ | new_n709_;
  assign new_n711_ = new_n605_ & ~\1_n1645 ;
  assign new_n712_ = ~new_n604_ & ~new_n711_;
  assign new_n713_ = \1_n1551  & ~\1_n1655 ;
  assign new_n714_ = ~\1_n362  & new_n713_;
  assign new_n715_ = ~\1_n1551  & ~\1_n1655 ;
  assign new_n716_ = \1_n664  & new_n606_;
  assign new_n717_ = \1_n325  & \1_n629 ;
  assign new_n718_ = \1_n507  & ~\1_n629 ;
  assign new_n719_ = ~new_n717_ & ~new_n718_;
  assign new_n720_ = new_n617_ & ~new_n719_;
  assign new_n721_ = ~new_n716_ & ~new_n720_;
  assign new_n722_ = \1_n842  & \1_n1606 ;
  assign new_n723_ = \1_n629  & ~\1_n1606 ;
  assign new_n724_ = ~new_n722_ & ~new_n723_;
  assign new_n725_ = \1_n1335  & ~\1_n1606 ;
  assign new_n726_ = \1_n1170  & \1_n1606 ;
  assign new_n727_ = ~new_n725_ & ~new_n726_;
  assign new_n728_ = \1_n1223  & \1_n1606 ;
  assign new_n729_ = \1_n490  & ~\1_n1606 ;
  assign new_n730_ = ~new_n728_ & ~new_n729_;
  assign new_n731_ = \1_n1165  & ~new_n730_;
  assign new_n732_ = \1_n1025  & \1_n1606 ;
  assign new_n733_ = \1_n654  & ~\1_n1606 ;
  assign new_n734_ = ~new_n732_ & ~new_n733_;
  assign new_n735_ = \1_n1389  & ~new_n734_;
  assign new_n736_ = \1_n1165  & new_n730_;
  assign new_n737_ = ~\1_n1165  & ~new_n730_;
  assign new_n738_ = ~new_n736_ & ~new_n737_;
  assign new_n739_ = new_n735_ & ~new_n738_;
  assign new_n740_ = ~new_n731_ & ~new_n739_;
  assign new_n741_ = ~\1_n574  & \1_n1606 ;
  assign new_n742_ = \1_n1545  & ~new_n741_;
  assign new_n743_ = ~\1_n1545  & new_n741_;
  assign new_n744_ = ~new_n742_ & ~new_n743_;
  assign new_n745_ = \1_n481  & \1_n1606 ;
  assign new_n746_ = \1_n646  & ~\1_n1606 ;
  assign new_n747_ = ~new_n745_ & ~new_n746_;
  assign new_n748_ = \1_n1378  & new_n747_;
  assign new_n749_ = ~\1_n1378  & ~new_n747_;
  assign new_n750_ = ~new_n748_ & ~new_n749_;
  assign new_n751_ = \1_n1596  & \1_n1606 ;
  assign new_n752_ = \1_n1518  & ~\1_n1606 ;
  assign new_n753_ = ~new_n751_ & ~new_n752_;
  assign new_n754_ = \1_n769  & new_n753_;
  assign new_n755_ = ~\1_n769  & ~new_n753_;
  assign new_n756_ = ~new_n754_ & ~new_n755_;
  assign new_n757_ = ~new_n750_ & ~new_n756_;
  assign new_n758_ = new_n744_ & new_n757_;
  assign new_n759_ = \1_n727  & \1_n1606 ;
  assign new_n760_ = \1_n1058  & ~\1_n1606 ;
  assign new_n761_ = ~new_n759_ & ~new_n760_;
  assign new_n762_ = \1_n403  & new_n761_;
  assign new_n763_ = ~\1_n403  & ~new_n761_;
  assign new_n764_ = ~new_n762_ & ~new_n763_;
  assign new_n765_ = new_n758_ & ~new_n764_;
  assign new_n766_ = \1_n1013  & \1_n1606 ;
  assign new_n767_ = \1_n1161  & ~\1_n1606 ;
  assign new_n768_ = ~new_n766_ & ~new_n767_;
  assign new_n769_ = new_n765_ & new_n768_;
  assign new_n770_ = \1_n1555  & new_n769_;
  assign new_n771_ = \1_n769  & ~new_n753_;
  assign new_n772_ = \1_n1378  & ~new_n747_;
  assign new_n773_ = ~new_n756_ & new_n772_;
  assign new_n774_ = ~new_n771_ & ~new_n773_;
  assign new_n775_ = new_n744_ & ~new_n774_;
  assign new_n776_ = ~new_n742_ & ~new_n775_;
  assign new_n777_ = new_n758_ & ~new_n768_;
  assign new_n778_ = new_n776_ & ~new_n777_;
  assign new_n779_ = ~new_n764_ & ~new_n778_;
  assign new_n780_ = \1_n403  & ~new_n761_;
  assign new_n781_ = ~new_n779_ & ~new_n780_;
  assign new_n782_ = ~new_n770_ & new_n781_;
  assign new_n783_ = new_n740_ & new_n782_;
  assign new_n784_ = \1_n1389  & new_n734_;
  assign new_n785_ = ~\1_n1389  & ~new_n734_;
  assign new_n786_ = ~new_n784_ & ~new_n785_;
  assign new_n787_ = ~new_n738_ & ~new_n786_;
  assign new_n788_ = new_n740_ & ~new_n787_;
  assign new_n789_ = ~new_n783_ & ~new_n788_;
  assign new_n790_ = new_n727_ & ~new_n789_;
  assign new_n791_ = new_n724_ & new_n790_;
  assign new_n792_ = ~new_n724_ & ~new_n790_;
  assign \1_n693  = new_n791_ | new_n792_;
  assign new_n794_ = new_n708_ & \1_n693 ;
  assign \1_n1478  = ~new_n721_ | new_n794_;
  assign new_n796_ = new_n715_ & ~\1_n1478 ;
  assign new_n797_ = ~new_n714_ & ~new_n796_;
  assign \1_n21  = ~new_n712_ | ~new_n797_;
  assign new_n799_ = ~\1_n84  & \1_n726 ;
  assign new_n800_ = ~\1_n468  & new_n799_;
  assign new_n801_ = ~\1_n84  & ~\1_n726 ;
  assign new_n802_ = \1_n230  & \1_n1545 ;
  assign new_n803_ = ~\1_n1425  & ~\1_n1545 ;
  assign new_n804_ = ~new_n802_ & ~new_n803_;
  assign new_n805_ = new_n617_ & ~new_n804_;
  assign new_n806_ = \1_n1189  & new_n606_;
  assign new_n807_ = ~new_n805_ & ~new_n806_;
  assign new_n808_ = \1_n1555  & new_n757_;
  assign new_n809_ = new_n757_ & ~new_n768_;
  assign new_n810_ = new_n774_ & ~new_n809_;
  assign new_n811_ = ~new_n808_ & new_n810_;
  assign new_n812_ = ~new_n744_ & new_n811_;
  assign new_n813_ = new_n744_ & ~new_n811_;
  assign new_n814_ = ~new_n812_ & ~new_n813_;
  assign new_n815_ = new_n708_ & new_n814_;
  assign \1_n1157  = ~new_n807_ | new_n815_;
  assign new_n817_ = new_n801_ & ~\1_n1157 ;
  assign new_n818_ = ~new_n800_ & ~new_n817_;
  assign new_n819_ = \1_n84  & \1_n726 ;
  assign new_n820_ = ~\1_n934  & new_n819_;
  assign new_n821_ = \1_n84  & ~\1_n726 ;
  assign new_n822_ = \1_n751  & new_n606_;
  assign new_n823_ = \1_n230  & \1_n956 ;
  assign new_n824_ = \1_n365  & ~\1_n956 ;
  assign new_n825_ = ~new_n823_ & ~new_n824_;
  assign new_n826_ = \1_n1479  & ~new_n825_;
  assign new_n827_ = ~\1_n956  & ~\1_n1255 ;
  assign new_n828_ = \1_n956  & ~\1_n1425 ;
  assign new_n829_ = ~new_n827_ & ~new_n828_;
  assign new_n830_ = ~\1_n1479  & ~new_n829_;
  assign new_n831_ = ~new_n826_ & ~new_n830_;
  assign new_n832_ = new_n617_ & ~new_n831_;
  assign new_n833_ = ~new_n822_ & ~new_n832_;
  assign new_n834_ = \1_n857  & new_n698_;
  assign new_n835_ = new_n688_ & ~new_n834_;
  assign new_n836_ = ~new_n666_ & ~new_n835_;
  assign new_n837_ = new_n666_ & new_n835_;
  assign new_n838_ = ~new_n836_ & ~new_n837_;
  assign new_n839_ = new_n708_ & new_n838_;
  assign \1_n928  = ~new_n833_ | new_n839_;
  assign new_n841_ = new_n821_ & ~\1_n928 ;
  assign new_n842_ = ~new_n820_ & ~new_n841_;
  assign new_n843_ = new_n818_ & new_n842_;
  assign \1_n24  = ~\1_n1310  | ~new_n843_;
  assign new_n845_ = ~\1_n989  & \1_n1413 ;
  assign new_n846_ = \1_n1121  & new_n845_;
  assign new_n847_ = \1_n837  & \1_n1065 ;
  assign new_n848_ = \1_n1311  & ~\1_n1335 ;
  assign new_n849_ = \1_n198  & \1_n1335 ;
  assign new_n850_ = ~new_n848_ & ~new_n849_;
  assign new_n851_ = new_n719_ & new_n850_;
  assign new_n852_ = ~new_n719_ & ~new_n850_;
  assign new_n853_ = ~new_n851_ & ~new_n852_;
  assign new_n854_ = \1_n325  & \1_n654 ;
  assign new_n855_ = \1_n507  & ~\1_n654 ;
  assign new_n856_ = ~new_n854_ & ~new_n855_;
  assign new_n857_ = ~\1_n1389  & ~new_n856_;
  assign new_n858_ = ~\1_n654  & ~\1_n1311 ;
  assign new_n859_ = ~\1_n198  & \1_n654 ;
  assign new_n860_ = ~new_n858_ & ~new_n859_;
  assign new_n861_ = \1_n1389  & ~new_n860_;
  assign new_n862_ = ~new_n857_ & ~new_n861_;
  assign new_n863_ = \1_n325  & \1_n490 ;
  assign new_n864_ = ~\1_n490  & \1_n507 ;
  assign new_n865_ = ~new_n863_ & ~new_n864_;
  assign new_n866_ = ~\1_n1165  & ~new_n865_;
  assign new_n867_ = ~\1_n490  & ~\1_n1311 ;
  assign new_n868_ = ~\1_n198  & \1_n490 ;
  assign new_n869_ = ~new_n867_ & ~new_n868_;
  assign new_n870_ = \1_n1165  & ~new_n869_;
  assign new_n871_ = ~new_n866_ & ~new_n870_;
  assign new_n872_ = new_n862_ & ~new_n871_;
  assign new_n873_ = ~new_n862_ & new_n871_;
  assign new_n874_ = ~new_n872_ & ~new_n873_;
  assign new_n875_ = new_n853_ & ~new_n874_;
  assign new_n876_ = ~new_n853_ & new_n874_;
  assign new_n877_ = ~new_n875_ & ~new_n876_;
  assign new_n878_ = \1_n325  & ~\1_n1545 ;
  assign new_n879_ = ~\1_n198  & \1_n1545 ;
  assign new_n880_ = ~new_n878_ & ~new_n879_;
  assign new_n881_ = \1_n325  & \1_n1058 ;
  assign new_n882_ = \1_n507  & ~\1_n1058 ;
  assign new_n883_ = ~new_n881_ & ~new_n882_;
  assign new_n884_ = ~\1_n403  & ~new_n883_;
  assign new_n885_ = ~\1_n1058  & ~\1_n1311 ;
  assign new_n886_ = ~\1_n198  & \1_n1058 ;
  assign new_n887_ = ~new_n885_ & ~new_n886_;
  assign new_n888_ = \1_n403  & ~new_n887_;
  assign new_n889_ = ~new_n884_ & ~new_n888_;
  assign new_n890_ = ~new_n880_ & new_n889_;
  assign new_n891_ = new_n880_ & ~new_n889_;
  assign new_n892_ = ~new_n890_ & ~new_n891_;
  assign new_n893_ = \1_n198  & \1_n1161 ;
  assign new_n894_ = ~\1_n1161  & \1_n1311 ;
  assign new_n895_ = ~new_n893_ & ~new_n894_;
  assign new_n896_ = \1_n325  & \1_n1518 ;
  assign new_n897_ = \1_n507  & ~\1_n1518 ;
  assign new_n898_ = ~new_n896_ & ~new_n897_;
  assign new_n899_ = ~\1_n769  & ~new_n898_;
  assign new_n900_ = ~\1_n1311  & ~\1_n1518 ;
  assign new_n901_ = ~\1_n198  & \1_n1518 ;
  assign new_n902_ = ~new_n900_ & ~new_n901_;
  assign new_n903_ = \1_n769  & ~new_n902_;
  assign new_n904_ = ~new_n899_ & ~new_n903_;
  assign new_n905_ = \1_n325  & \1_n646 ;
  assign new_n906_ = \1_n507  & ~\1_n646 ;
  assign new_n907_ = ~new_n905_ & ~new_n906_;
  assign new_n908_ = ~\1_n1378  & ~new_n907_;
  assign new_n909_ = ~\1_n646  & ~\1_n1311 ;
  assign new_n910_ = ~\1_n198  & \1_n646 ;
  assign new_n911_ = ~new_n909_ & ~new_n910_;
  assign new_n912_ = \1_n1378  & ~new_n911_;
  assign new_n913_ = ~new_n908_ & ~new_n912_;
  assign new_n914_ = ~new_n904_ & ~new_n913_;
  assign new_n915_ = new_n904_ & new_n913_;
  assign new_n916_ = ~new_n914_ & ~new_n915_;
  assign new_n917_ = new_n895_ & new_n916_;
  assign new_n918_ = ~new_n895_ & ~new_n916_;
  assign new_n919_ = ~new_n917_ & ~new_n918_;
  assign new_n920_ = ~new_n892_ & new_n919_;
  assign new_n921_ = new_n892_ & ~new_n919_;
  assign new_n922_ = ~new_n920_ & ~new_n921_;
  assign new_n923_ = ~new_n877_ & new_n922_;
  assign new_n924_ = new_n877_ & ~new_n922_;
  assign new_n925_ = ~new_n923_ & ~new_n924_;
  assign new_n926_ = new_n617_ & ~new_n925_;
  assign new_n927_ = ~new_n750_ & ~new_n768_;
  assign new_n928_ = ~new_n772_ & ~new_n927_;
  assign new_n929_ = new_n744_ & ~new_n764_;
  assign new_n930_ = ~new_n744_ & new_n764_;
  assign new_n931_ = ~new_n929_ & ~new_n930_;
  assign new_n932_ = new_n928_ & new_n931_;
  assign new_n933_ = ~new_n928_ & ~new_n931_;
  assign new_n934_ = ~new_n932_ & ~new_n933_;
  assign new_n935_ = ~new_n768_ & new_n810_;
  assign new_n936_ = new_n768_ & ~new_n810_;
  assign new_n937_ = ~new_n935_ & ~new_n936_;
  assign new_n938_ = ~new_n934_ & new_n937_;
  assign new_n939_ = new_n934_ & ~new_n937_;
  assign new_n940_ = ~new_n938_ & ~new_n939_;
  assign new_n941_ = new_n750_ & new_n768_;
  assign new_n942_ = ~new_n927_ & ~new_n941_;
  assign new_n943_ = ~new_n756_ & new_n942_;
  assign new_n944_ = new_n756_ & ~new_n942_;
  assign new_n945_ = ~new_n943_ & ~new_n944_;
  assign new_n946_ = ~new_n778_ & new_n945_;
  assign new_n947_ = new_n778_ & ~new_n945_;
  assign new_n948_ = ~new_n946_ & ~new_n947_;
  assign new_n949_ = ~new_n940_ & new_n948_;
  assign new_n950_ = new_n940_ & ~new_n948_;
  assign new_n951_ = ~new_n949_ & ~new_n950_;
  assign new_n952_ = ~\1_n1  & ~new_n951_;
  assign new_n953_ = ~new_n750_ & new_n768_;
  assign new_n954_ = new_n928_ & ~new_n953_;
  assign new_n955_ = ~new_n757_ & new_n774_;
  assign new_n956_ = ~new_n758_ & new_n776_;
  assign new_n957_ = ~new_n955_ & new_n956_;
  assign new_n958_ = new_n955_ & ~new_n956_;
  assign new_n959_ = ~new_n957_ & ~new_n958_;
  assign new_n960_ = ~new_n945_ & new_n959_;
  assign new_n961_ = new_n945_ & ~new_n959_;
  assign new_n962_ = ~new_n960_ & ~new_n961_;
  assign new_n963_ = ~new_n931_ & new_n962_;
  assign new_n964_ = new_n931_ & ~new_n962_;
  assign new_n965_ = ~new_n963_ & ~new_n964_;
  assign new_n966_ = ~new_n954_ & new_n965_;
  assign new_n967_ = new_n954_ & ~new_n965_;
  assign new_n968_ = ~new_n966_ & ~new_n967_;
  assign new_n969_ = \1_n1  & new_n968_;
  assign new_n970_ = ~new_n952_ & ~new_n969_;
  assign new_n971_ = new_n724_ & new_n727_;
  assign new_n972_ = ~new_n724_ & ~new_n727_;
  assign new_n973_ = ~new_n971_ & ~new_n972_;
  assign new_n974_ = new_n740_ & new_n973_;
  assign new_n975_ = ~new_n740_ & ~new_n973_;
  assign new_n976_ = ~new_n974_ & ~new_n975_;
  assign new_n977_ = new_n738_ & new_n786_;
  assign new_n978_ = ~new_n787_ & ~new_n977_;
  assign new_n979_ = new_n727_ & new_n740_;
  assign new_n980_ = ~new_n735_ & new_n979_;
  assign new_n981_ = new_n735_ & ~new_n979_;
  assign new_n982_ = ~new_n980_ & ~new_n981_;
  assign new_n983_ = new_n978_ & ~new_n982_;
  assign new_n984_ = ~new_n978_ & new_n982_;
  assign new_n985_ = ~new_n983_ & ~new_n984_;
  assign new_n986_ = ~new_n976_ & new_n985_;
  assign new_n987_ = new_n976_ & ~new_n985_;
  assign new_n988_ = ~new_n986_ & ~new_n987_;
  assign new_n989_ = \1_n1  & new_n769_;
  assign new_n990_ = new_n781_ & ~new_n989_;
  assign new_n991_ = ~new_n988_ & new_n990_;
  assign new_n992_ = ~new_n788_ & ~new_n973_;
  assign new_n993_ = new_n788_ & new_n973_;
  assign new_n994_ = ~new_n992_ & ~new_n993_;
  assign new_n995_ = ~new_n735_ & new_n786_;
  assign new_n996_ = new_n727_ & new_n788_;
  assign new_n997_ = ~new_n995_ & new_n996_;
  assign new_n998_ = new_n995_ & ~new_n996_;
  assign new_n999_ = ~new_n997_ & ~new_n998_;
  assign new_n1000_ = new_n978_ & new_n999_;
  assign new_n1001_ = ~new_n978_ & ~new_n999_;
  assign new_n1002_ = ~new_n1000_ & ~new_n1001_;
  assign new_n1003_ = ~new_n994_ & new_n1002_;
  assign new_n1004_ = new_n994_ & ~new_n1002_;
  assign new_n1005_ = ~new_n1003_ & ~new_n1004_;
  assign new_n1006_ = ~new_n990_ & new_n1005_;
  assign new_n1007_ = ~new_n991_ & ~new_n1006_;
  assign new_n1008_ = ~new_n970_ & ~new_n1007_;
  assign new_n1009_ = new_n970_ & new_n1007_;
  assign new_n1010_ = ~new_n1008_ & ~new_n1009_;
  assign new_n1011_ = new_n708_ & ~new_n1010_;
  assign new_n1012_ = ~new_n926_ & ~new_n1011_;
  assign new_n1013_ = ~new_n847_ & new_n1012_;
  assign new_n1014_ = ~\1_n989  & ~\1_n1413 ;
  assign new_n1015_ = ~new_n1013_ & new_n1014_;
  assign new_n1016_ = ~new_n846_ & ~new_n1015_;
  assign new_n1017_ = \1_n989  & \1_n1413 ;
  assign new_n1018_ = \1_n1515  & new_n1017_;
  assign new_n1019_ = \1_n901  & \1_n1065 ;
  assign new_n1020_ = \1_n325  & \1_n824 ;
  assign new_n1021_ = \1_n507  & ~\1_n824 ;
  assign new_n1022_ = ~new_n1020_ & ~new_n1021_;
  assign new_n1023_ = ~\1_n1530  & ~new_n1022_;
  assign new_n1024_ = ~\1_n824  & ~\1_n1311 ;
  assign new_n1025_ = ~\1_n198  & \1_n824 ;
  assign new_n1026_ = ~new_n1024_ & ~new_n1025_;
  assign new_n1027_ = \1_n1530  & ~new_n1026_;
  assign new_n1028_ = ~new_n1023_ & ~new_n1027_;
  assign new_n1029_ = \1_n135  & \1_n325 ;
  assign new_n1030_ = ~\1_n135  & \1_n507 ;
  assign new_n1031_ = ~new_n1029_ & ~new_n1030_;
  assign new_n1032_ = ~\1_n765  & ~new_n1031_;
  assign new_n1033_ = ~\1_n135  & ~\1_n1311 ;
  assign new_n1034_ = \1_n135  & ~\1_n198 ;
  assign new_n1035_ = ~new_n1033_ & ~new_n1034_;
  assign new_n1036_ = \1_n765  & ~new_n1035_;
  assign new_n1037_ = ~new_n1032_ & ~new_n1036_;
  assign new_n1038_ = ~new_n1028_ & ~new_n1037_;
  assign new_n1039_ = new_n1028_ & new_n1037_;
  assign new_n1040_ = ~new_n1038_ & ~new_n1039_;
  assign new_n1041_ = \1_n325  & \1_n859 ;
  assign new_n1042_ = \1_n507  & ~\1_n859 ;
  assign new_n1043_ = ~new_n1041_ & ~new_n1042_;
  assign new_n1044_ = ~\1_n184  & ~new_n1043_;
  assign new_n1045_ = ~\1_n859  & ~\1_n1311 ;
  assign new_n1046_ = ~\1_n198  & \1_n859 ;
  assign new_n1047_ = ~new_n1045_ & ~new_n1046_;
  assign new_n1048_ = \1_n184  & ~new_n1047_;
  assign new_n1049_ = ~new_n1044_ & ~new_n1048_;
  assign new_n1050_ = new_n616_ & new_n1049_;
  assign new_n1051_ = ~new_n616_ & ~new_n1049_;
  assign new_n1052_ = ~new_n1050_ & ~new_n1051_;
  assign new_n1053_ = ~new_n1040_ & new_n1052_;
  assign new_n1054_ = new_n1040_ & ~new_n1052_;
  assign new_n1055_ = ~new_n1053_ & ~new_n1054_;
  assign new_n1056_ = \1_n325  & \1_n1143 ;
  assign new_n1057_ = \1_n507  & ~\1_n1143 ;
  assign new_n1058_ = ~new_n1056_ & ~new_n1057_;
  assign new_n1059_ = ~\1_n1108  & ~new_n1058_;
  assign new_n1060_ = ~\1_n1143  & ~\1_n1311 ;
  assign new_n1061_ = ~\1_n198  & \1_n1143 ;
  assign new_n1062_ = ~new_n1060_ & ~new_n1061_;
  assign new_n1063_ = \1_n1108  & ~new_n1062_;
  assign new_n1064_ = ~new_n1059_ & ~new_n1063_;
  assign new_n1065_ = \1_n325  & \1_n956 ;
  assign new_n1066_ = \1_n507  & ~\1_n956 ;
  assign new_n1067_ = ~new_n1065_ & ~new_n1066_;
  assign new_n1068_ = ~\1_n1479  & ~new_n1067_;
  assign new_n1069_ = ~\1_n956  & ~\1_n1311 ;
  assign new_n1070_ = ~\1_n198  & \1_n956 ;
  assign new_n1071_ = ~new_n1069_ & ~new_n1070_;
  assign new_n1072_ = \1_n1479  & ~new_n1071_;
  assign new_n1073_ = ~new_n1068_ & ~new_n1072_;
  assign new_n1074_ = ~new_n1064_ & new_n1073_;
  assign new_n1075_ = new_n1064_ & ~new_n1073_;
  assign new_n1076_ = ~new_n1074_ & ~new_n1075_;
  assign new_n1077_ = \1_n209  & \1_n325 ;
  assign new_n1078_ = ~\1_n209  & \1_n507 ;
  assign new_n1079_ = ~new_n1077_ & ~new_n1078_;
  assign new_n1080_ = ~\1_n950  & ~new_n1079_;
  assign new_n1081_ = ~\1_n209  & ~\1_n1311 ;
  assign new_n1082_ = ~\1_n198  & \1_n209 ;
  assign new_n1083_ = ~new_n1081_ & ~new_n1082_;
  assign new_n1084_ = \1_n950  & ~new_n1083_;
  assign new_n1085_ = ~new_n1080_ & ~new_n1084_;
  assign new_n1086_ = \1_n325  & \1_n1251 ;
  assign new_n1087_ = \1_n507  & ~\1_n1251 ;
  assign new_n1088_ = ~new_n1086_ & ~new_n1087_;
  assign new_n1089_ = ~\1_n147  & ~new_n1088_;
  assign new_n1090_ = ~\1_n1251  & ~\1_n1311 ;
  assign new_n1091_ = ~\1_n198  & \1_n1251 ;
  assign new_n1092_ = ~new_n1090_ & ~new_n1091_;
  assign new_n1093_ = \1_n147  & ~new_n1092_;
  assign new_n1094_ = ~new_n1089_ & ~new_n1093_;
  assign new_n1095_ = \1_n325  & \1_n1030 ;
  assign new_n1096_ = \1_n507  & ~\1_n1030 ;
  assign new_n1097_ = ~new_n1095_ & ~new_n1096_;
  assign new_n1098_ = ~\1_n938  & ~new_n1097_;
  assign new_n1099_ = ~\1_n1030  & ~\1_n1311 ;
  assign new_n1100_ = ~\1_n198  & \1_n1030 ;
  assign new_n1101_ = ~new_n1099_ & ~new_n1100_;
  assign new_n1102_ = \1_n938  & ~new_n1101_;
  assign new_n1103_ = ~new_n1098_ & ~new_n1102_;
  assign new_n1104_ = ~new_n1094_ & ~new_n1103_;
  assign new_n1105_ = new_n1094_ & new_n1103_;
  assign new_n1106_ = ~new_n1104_ & ~new_n1105_;
  assign new_n1107_ = ~new_n1085_ & new_n1106_;
  assign new_n1108_ = new_n1085_ & ~new_n1106_;
  assign new_n1109_ = ~new_n1107_ & ~new_n1108_;
  assign new_n1110_ = ~new_n1076_ & new_n1109_;
  assign new_n1111_ = new_n1076_ & ~new_n1109_;
  assign new_n1112_ = ~new_n1110_ & ~new_n1111_;
  assign new_n1113_ = ~new_n1055_ & new_n1112_;
  assign new_n1114_ = new_n1055_ & ~new_n1112_;
  assign new_n1115_ = ~new_n1113_ & ~new_n1114_;
  assign new_n1116_ = new_n617_ & ~new_n1115_;
  assign new_n1117_ = ~new_n659_ & ~new_n666_;
  assign new_n1118_ = new_n659_ & new_n666_;
  assign new_n1119_ = ~new_n1117_ & ~new_n1118_;
  assign new_n1120_ = new_n683_ & ~new_n1119_;
  assign new_n1121_ = ~new_n683_ & new_n1119_;
  assign new_n1122_ = ~new_n1120_ & ~new_n1121_;
  assign new_n1123_ = new_n678_ & ~new_n688_;
  assign new_n1124_ = ~new_n678_ & new_n688_;
  assign new_n1125_ = ~new_n1123_ & ~new_n1124_;
  assign new_n1126_ = ~new_n1122_ & new_n1125_;
  assign new_n1127_ = new_n1122_ & ~new_n1125_;
  assign new_n1128_ = ~new_n1126_ & ~new_n1127_;
  assign new_n1129_ = ~new_n690_ & new_n696_;
  assign new_n1130_ = new_n690_ & ~new_n696_;
  assign new_n1131_ = ~new_n1129_ & ~new_n1130_;
  assign new_n1132_ = new_n681_ & new_n686_;
  assign new_n1133_ = ~new_n681_ & ~new_n686_;
  assign new_n1134_ = ~new_n1132_ & ~new_n1133_;
  assign new_n1135_ = ~new_n1131_ & ~new_n1134_;
  assign new_n1136_ = new_n1131_ & new_n1134_;
  assign new_n1137_ = ~new_n1135_ & ~new_n1136_;
  assign new_n1138_ = ~new_n1128_ & new_n1137_;
  assign new_n1139_ = new_n1128_ & ~new_n1137_;
  assign new_n1140_ = ~new_n1138_ & ~new_n1139_;
  assign new_n1141_ = ~\1_n283  & ~new_n1140_;
  assign new_n1142_ = new_n683_ & ~new_n697_;
  assign new_n1143_ = ~new_n659_ & ~new_n686_;
  assign new_n1144_ = new_n659_ & new_n686_;
  assign new_n1145_ = ~new_n1143_ & ~new_n1144_;
  assign new_n1146_ = ~new_n1142_ & ~new_n1145_;
  assign new_n1147_ = new_n1142_ & new_n1145_;
  assign new_n1148_ = ~new_n1146_ & ~new_n1147_;
  assign new_n1149_ = new_n688_ & ~new_n698_;
  assign new_n1150_ = ~new_n678_ & new_n696_;
  assign new_n1151_ = ~new_n1149_ & ~new_n1150_;
  assign new_n1152_ = new_n1149_ & new_n1150_;
  assign new_n1153_ = ~new_n1151_ & ~new_n1152_;
  assign new_n1154_ = ~new_n1148_ & new_n1153_;
  assign new_n1155_ = new_n1148_ & ~new_n1153_;
  assign new_n1156_ = ~new_n1154_ & ~new_n1155_;
  assign new_n1157_ = ~new_n666_ & new_n681_;
  assign new_n1158_ = new_n666_ & ~new_n681_;
  assign new_n1159_ = ~new_n1157_ & ~new_n1158_;
  assign new_n1160_ = ~new_n699_ & new_n1130_;
  assign new_n1161_ = ~new_n1129_ & ~new_n1160_;
  assign new_n1162_ = ~new_n1159_ & ~new_n1161_;
  assign new_n1163_ = new_n1159_ & new_n1161_;
  assign new_n1164_ = ~new_n1162_ & ~new_n1163_;
  assign new_n1165_ = ~new_n1156_ & new_n1164_;
  assign new_n1166_ = new_n1156_ & ~new_n1164_;
  assign new_n1167_ = ~new_n1165_ & ~new_n1166_;
  assign new_n1168_ = \1_n283  & new_n1167_;
  assign new_n1169_ = ~new_n1141_ & ~new_n1168_;
  assign new_n1170_ = \1_n283  & new_n699_;
  assign new_n1171_ = ~new_n659_ & new_n1170_;
  assign new_n1172_ = new_n693_ & ~new_n1171_;
  assign new_n1173_ = ~new_n625_ & new_n631_;
  assign new_n1174_ = new_n625_ & ~new_n631_;
  assign new_n1175_ = ~new_n1173_ & ~new_n1174_;
  assign new_n1176_ = new_n644_ & new_n1175_;
  assign new_n1177_ = ~new_n644_ & ~new_n1175_;
  assign new_n1178_ = ~new_n1176_ & ~new_n1177_;
  assign new_n1179_ = ~new_n642_ & new_n650_;
  assign new_n1180_ = new_n642_ & ~new_n650_;
  assign new_n1181_ = ~new_n1179_ & ~new_n1180_;
  assign new_n1182_ = new_n639_ & new_n647_;
  assign new_n1183_ = ~new_n639_ & ~new_n647_;
  assign new_n1184_ = ~new_n1182_ & ~new_n1183_;
  assign new_n1185_ = ~new_n1181_ & ~new_n1184_;
  assign new_n1186_ = new_n1181_ & new_n1184_;
  assign new_n1187_ = ~new_n1185_ & ~new_n1186_;
  assign new_n1188_ = new_n1178_ & new_n1187_;
  assign new_n1189_ = ~new_n1178_ & ~new_n1187_;
  assign new_n1190_ = ~new_n1188_ & ~new_n1189_;
  assign new_n1191_ = new_n1172_ & new_n1190_;
  assign new_n1192_ = new_n644_ & ~new_n651_;
  assign new_n1193_ = ~new_n1175_ & new_n1192_;
  assign new_n1194_ = new_n1175_ & ~new_n1192_;
  assign new_n1195_ = ~new_n1193_ & ~new_n1194_;
  assign new_n1196_ = ~new_n639_ & new_n650_;
  assign new_n1197_ = ~new_n653_ & new_n1196_;
  assign new_n1198_ = new_n653_ & ~new_n1196_;
  assign new_n1199_ = ~new_n1197_ & ~new_n1198_;
  assign new_n1200_ = ~new_n1181_ & ~new_n1199_;
  assign new_n1201_ = new_n1181_ & new_n1199_;
  assign new_n1202_ = ~new_n1200_ & ~new_n1201_;
  assign new_n1203_ = ~new_n1195_ & new_n1202_;
  assign new_n1204_ = new_n1195_ & ~new_n1202_;
  assign new_n1205_ = ~new_n1203_ & ~new_n1204_;
  assign new_n1206_ = ~new_n1172_ & ~new_n1205_;
  assign new_n1207_ = ~new_n1191_ & ~new_n1206_;
  assign new_n1208_ = ~new_n1169_ & ~new_n1207_;
  assign new_n1209_ = new_n1169_ & new_n1207_;
  assign new_n1210_ = ~new_n1208_ & ~new_n1209_;
  assign new_n1211_ = new_n708_ & ~new_n1210_;
  assign new_n1212_ = ~new_n1116_ & ~new_n1211_;
  assign new_n1213_ = ~new_n1019_ & new_n1212_;
  assign new_n1214_ = \1_n989  & ~\1_n1413 ;
  assign new_n1215_ = ~new_n1213_ & new_n1214_;
  assign new_n1216_ = ~new_n1018_ & ~new_n1215_;
  assign new_n1217_ = new_n1016_ & new_n1216_;
  assign \1_n32  = \1_n24 ;
  assign new_n1219_ = ~\1_n1555  & new_n768_;
  assign new_n1220_ = new_n750_ & ~new_n1219_;
  assign new_n1221_ = ~\1_n1555  & new_n953_;
  assign new_n1222_ = ~new_n1220_ & ~new_n1221_;
  assign new_n1223_ = \1_n1555  & new_n768_;
  assign new_n1224_ = ~\1_n1555  & ~new_n768_;
  assign new_n1225_ = ~new_n1223_ & ~new_n1224_;
  assign new_n1226_ = \1_n1555  & ~new_n750_;
  assign new_n1227_ = new_n928_ & ~new_n1226_;
  assign new_n1228_ = ~new_n756_ & ~new_n1227_;
  assign new_n1229_ = new_n756_ & new_n1227_;
  assign new_n1230_ = ~new_n1228_ & ~new_n1229_;
  assign new_n1231_ = \1_n1555  & new_n758_;
  assign new_n1232_ = new_n778_ & ~new_n1231_;
  assign new_n1233_ = ~new_n764_ & ~new_n1232_;
  assign new_n1234_ = new_n764_ & new_n1232_;
  assign new_n1235_ = ~new_n1233_ & ~new_n1234_;
  assign new_n1236_ = ~new_n782_ & ~new_n786_;
  assign new_n1237_ = new_n782_ & new_n786_;
  assign new_n1238_ = ~new_n1236_ & ~new_n1237_;
  assign new_n1239_ = ~new_n735_ & new_n782_;
  assign new_n1240_ = ~new_n995_ & ~new_n1239_;
  assign new_n1241_ = ~new_n738_ & ~new_n1240_;
  assign new_n1242_ = new_n738_ & new_n1240_;
  assign new_n1243_ = ~new_n1241_ & ~new_n1242_;
  assign new_n1244_ = new_n727_ & new_n789_;
  assign new_n1245_ = ~new_n727_ & ~new_n789_;
  assign new_n1246_ = ~new_n1244_ & ~new_n1245_;
  assign new_n1247_ = new_n1243_ & ~new_n1246_;
  assign new_n1248_ = ~new_n1238_ & new_n1247_;
  assign new_n1249_ = ~new_n1235_ & new_n1248_;
  assign new_n1250_ = ~new_n814_ & new_n1249_;
  assign new_n1251_ = ~new_n1230_ & new_n1250_;
  assign new_n1252_ = ~new_n1225_ & new_n1251_;
  assign new_n1253_ = new_n1222_ & new_n1252_;
  assign \1_n54  = \1_n693  | ~new_n1253_;
  assign new_n1255_ = \1_n182  & \1_n877 ;
  assign new_n1256_ = ~\1_n923  & new_n1255_;
  assign new_n1257_ = ~\1_n182  & ~\1_n877 ;
  assign new_n1258_ = new_n1013_ & new_n1257_;
  assign new_n1259_ = ~new_n1256_ & ~new_n1258_;
  assign new_n1260_ = ~\1_n182  & \1_n877 ;
  assign new_n1261_ = ~\1_n1280  & new_n1260_;
  assign new_n1262_ = \1_n182  & ~\1_n877 ;
  assign new_n1263_ = new_n1213_ & new_n1262_;
  assign new_n1264_ = ~new_n1261_ & ~new_n1263_;
  assign \1_n64  = ~new_n1259_ | ~new_n1264_;
  assign new_n1266_ = ~\1_n1511  & new_n819_;
  assign new_n1267_ = \1_n1418  & new_n606_;
  assign new_n1268_ = \1_n230  & \1_n1251 ;
  assign new_n1269_ = \1_n365  & ~\1_n1251 ;
  assign new_n1270_ = ~new_n1268_ & ~new_n1269_;
  assign new_n1271_ = \1_n147  & ~new_n1270_;
  assign new_n1272_ = ~\1_n1251  & ~\1_n1255 ;
  assign new_n1273_ = \1_n1251  & ~\1_n1425 ;
  assign new_n1274_ = ~new_n1272_ & ~new_n1273_;
  assign new_n1275_ = ~\1_n147  & ~new_n1274_;
  assign new_n1276_ = ~new_n1271_ & ~new_n1275_;
  assign new_n1277_ = new_n617_ & ~new_n1276_;
  assign new_n1278_ = ~new_n1267_ & ~new_n1277_;
  assign new_n1279_ = \1_n857  & ~new_n696_;
  assign new_n1280_ = ~new_n681_ & new_n1279_;
  assign new_n1281_ = new_n683_ & ~new_n1280_;
  assign new_n1282_ = new_n686_ & new_n1281_;
  assign new_n1283_ = ~new_n686_ & ~new_n1281_;
  assign new_n1284_ = ~new_n1282_ & ~new_n1283_;
  assign new_n1285_ = new_n708_ & new_n1284_;
  assign \1_n1589  = ~new_n1278_ | new_n1285_;
  assign new_n1287_ = new_n821_ & ~\1_n1589 ;
  assign new_n1288_ = ~new_n1266_ & ~new_n1287_;
  assign new_n1289_ = ~\1_n909  & new_n799_;
  assign new_n1290_ = \1_n1049  & new_n606_;
  assign new_n1291_ = \1_n230  & \1_n1518 ;
  assign new_n1292_ = \1_n365  & ~\1_n1518 ;
  assign new_n1293_ = ~new_n1291_ & ~new_n1292_;
  assign new_n1294_ = \1_n769  & ~new_n1293_;
  assign new_n1295_ = ~\1_n1255  & ~\1_n1518 ;
  assign new_n1296_ = ~\1_n1425  & \1_n1518 ;
  assign new_n1297_ = ~new_n1295_ & ~new_n1296_;
  assign new_n1298_ = ~\1_n769  & ~new_n1297_;
  assign new_n1299_ = ~new_n1294_ & ~new_n1298_;
  assign new_n1300_ = new_n617_ & ~new_n1299_;
  assign new_n1301_ = ~new_n1290_ & ~new_n1300_;
  assign new_n1302_ = new_n708_ & new_n1230_;
  assign \1_n1177  = ~new_n1301_ | new_n1302_;
  assign new_n1304_ = new_n801_ & ~\1_n1177 ;
  assign new_n1305_ = ~new_n1289_ & ~new_n1304_;
  assign new_n1306_ = new_n1288_ & new_n1305_;
  assign \1_n76  = \1_n24 ;
  assign \1_n167  = \1_n421  & \1_n1412 ;
  assign \1_n83  = \1_n415  & \1_n167 ;
  assign new_n1310_ = ~\1_n933  & new_n1260_;
  assign new_n1311_ = new_n1262_ & ~\1_n1589 ;
  assign new_n1312_ = ~new_n1310_ & ~new_n1311_;
  assign new_n1313_ = ~\1_n1042  & new_n1255_;
  assign new_n1314_ = new_n1257_ & ~\1_n1177 ;
  assign new_n1315_ = ~new_n1313_ & ~new_n1314_;
  assign \1_n97  = ~new_n1312_ | ~new_n1315_;
  assign new_n1317_ = new_n769_ & new_n787_;
  assign new_n1318_ = new_n724_ & new_n1317_;
  assign \1_n110  = ~new_n727_ | ~new_n1318_;
  assign new_n1320_ = \1_n230  & \1_n1030 ;
  assign new_n1321_ = \1_n365  & ~\1_n1030 ;
  assign new_n1322_ = ~new_n1320_ & ~new_n1321_;
  assign new_n1323_ = \1_n938  & ~new_n1322_;
  assign new_n1324_ = ~\1_n1030  & ~\1_n1255 ;
  assign new_n1325_ = \1_n1030  & ~\1_n1425 ;
  assign new_n1326_ = ~new_n1324_ & ~new_n1325_;
  assign new_n1327_ = ~\1_n938  & ~new_n1326_;
  assign new_n1328_ = ~new_n1323_ & ~new_n1327_;
  assign new_n1329_ = \1_n209  & \1_n230 ;
  assign new_n1330_ = ~\1_n209  & \1_n365 ;
  assign new_n1331_ = ~new_n1329_ & ~new_n1330_;
  assign new_n1332_ = \1_n950  & ~new_n1331_;
  assign new_n1333_ = ~\1_n209  & ~\1_n1255 ;
  assign new_n1334_ = \1_n209  & ~\1_n1425 ;
  assign new_n1335_ = ~new_n1333_ & ~new_n1334_;
  assign new_n1336_ = ~\1_n950  & ~new_n1335_;
  assign new_n1337_ = ~new_n1332_ & ~new_n1336_;
  assign new_n1338_ = \1_n230  & \1_n1143 ;
  assign new_n1339_ = \1_n365  & ~\1_n1143 ;
  assign new_n1340_ = ~new_n1338_ & ~new_n1339_;
  assign new_n1341_ = \1_n1108  & ~new_n1340_;
  assign new_n1342_ = ~\1_n1143  & ~\1_n1255 ;
  assign new_n1343_ = \1_n1143  & ~\1_n1425 ;
  assign new_n1344_ = ~new_n1342_ & ~new_n1343_;
  assign new_n1345_ = ~\1_n1108  & ~new_n1344_;
  assign new_n1346_ = ~new_n1341_ & ~new_n1345_;
  assign new_n1347_ = \1_n135  & \1_n230 ;
  assign new_n1348_ = ~\1_n135  & \1_n365 ;
  assign new_n1349_ = ~new_n1347_ & ~new_n1348_;
  assign new_n1350_ = \1_n765  & ~new_n1349_;
  assign new_n1351_ = ~\1_n135  & ~\1_n1255 ;
  assign new_n1352_ = \1_n135  & ~\1_n1425 ;
  assign new_n1353_ = ~new_n1351_ & ~new_n1352_;
  assign new_n1354_ = ~\1_n765  & ~new_n1353_;
  assign new_n1355_ = ~new_n1350_ & ~new_n1354_;
  assign new_n1356_ = ~\1_n824  & ~\1_n1255 ;
  assign new_n1357_ = \1_n824  & ~\1_n1425 ;
  assign new_n1358_ = ~new_n1356_ & ~new_n1357_;
  assign new_n1359_ = ~\1_n1530  & ~new_n1358_;
  assign new_n1360_ = \1_n365  & ~\1_n824 ;
  assign new_n1361_ = \1_n230  & \1_n824 ;
  assign new_n1362_ = ~new_n1360_ & ~new_n1361_;
  assign new_n1363_ = \1_n1530  & ~new_n1362_;
  assign new_n1364_ = ~new_n1359_ & ~new_n1363_;
  assign new_n1365_ = ~\1_n859  & ~\1_n1255 ;
  assign new_n1366_ = \1_n859  & ~\1_n1425 ;
  assign new_n1367_ = ~new_n1365_ & ~new_n1366_;
  assign new_n1368_ = ~\1_n184  & ~new_n1367_;
  assign new_n1369_ = \1_n365  & ~\1_n859 ;
  assign new_n1370_ = \1_n230  & \1_n859 ;
  assign new_n1371_ = ~new_n1369_ & ~new_n1370_;
  assign new_n1372_ = \1_n184  & ~new_n1371_;
  assign new_n1373_ = ~new_n1368_ & ~new_n1372_;
  assign new_n1374_ = new_n1364_ & new_n1373_;
  assign new_n1375_ = new_n1355_ & new_n1374_;
  assign new_n1376_ = new_n1346_ & new_n1375_;
  assign new_n1377_ = new_n831_ & new_n1376_;
  assign new_n1378_ = new_n1276_ & new_n1377_;
  assign new_n1379_ = new_n1337_ & new_n1378_;
  assign new_n1380_ = new_n1328_ & new_n1379_;
  assign \1_n117  = ~new_n616_ | ~new_n1380_;
  assign new_n1382_ = ~new_n625_ & new_n652_;
  assign new_n1383_ = new_n699_ & new_n1382_;
  assign \1_n142  = new_n659_ | ~new_n1383_;
  assign new_n1385_ = ~\1_n1146  & new_n799_;
  assign new_n1386_ = \1_n1580  & new_n606_;
  assign new_n1387_ = new_n617_ & ~new_n862_;
  assign new_n1388_ = ~new_n1386_ & ~new_n1387_;
  assign new_n1389_ = new_n708_ & new_n1238_;
  assign \1_n434  = ~new_n1388_ | new_n1389_;
  assign new_n1391_ = new_n801_ & ~\1_n434 ;
  assign new_n1392_ = ~new_n1385_ & ~new_n1391_;
  assign new_n1393_ = ~\1_n1398  & new_n819_;
  assign new_n1394_ = \1_n233  & new_n606_;
  assign new_n1395_ = new_n617_ & ~new_n1355_;
  assign new_n1396_ = ~new_n1394_ & ~new_n1395_;
  assign new_n1397_ = ~new_n650_ & ~new_n702_;
  assign new_n1398_ = new_n650_ & new_n702_;
  assign new_n1399_ = ~new_n1397_ & ~new_n1398_;
  assign new_n1400_ = new_n708_ & new_n1399_;
  assign \1_n675  = ~new_n1396_ | new_n1400_;
  assign new_n1402_ = new_n821_ & ~\1_n675 ;
  assign new_n1403_ = ~new_n1393_ & ~new_n1402_;
  assign new_n1404_ = new_n1392_ & new_n1403_;
  assign \1_n150  = \1_n24 ;
  assign new_n1406_ = ~new_n678_ & ~new_n1279_;
  assign new_n1407_ = ~new_n681_ & ~new_n1406_;
  assign new_n1408_ = new_n681_ & new_n1406_;
  assign new_n1409_ = ~new_n1407_ & ~new_n1408_;
  assign new_n1410_ = ~\1_n857  & new_n696_;
  assign new_n1411_ = ~new_n1279_ & ~new_n1410_;
  assign new_n1412_ = new_n690_ & ~new_n700_;
  assign new_n1413_ = ~new_n659_ & ~new_n1412_;
  assign new_n1414_ = new_n659_ & new_n1412_;
  assign new_n1415_ = ~new_n1413_ & ~new_n1414_;
  assign new_n1416_ = ~new_n639_ & new_n702_;
  assign new_n1417_ = ~new_n1196_ & ~new_n1416_;
  assign new_n1418_ = new_n642_ & ~new_n1417_;
  assign new_n1419_ = ~new_n642_ & new_n1417_;
  assign new_n1420_ = ~new_n1418_ & ~new_n1419_;
  assign new_n1421_ = ~new_n702_ & ~new_n1192_;
  assign new_n1422_ = new_n644_ & ~new_n1421_;
  assign new_n1423_ = ~new_n631_ & new_n1422_;
  assign new_n1424_ = new_n631_ & ~new_n1422_;
  assign new_n1425_ = ~new_n1423_ & ~new_n1424_;
  assign new_n1426_ = ~new_n707_ & new_n1425_;
  assign new_n1427_ = ~new_n1420_ & new_n1426_;
  assign new_n1428_ = ~new_n1399_ & new_n1427_;
  assign new_n1429_ = ~new_n1415_ & new_n1428_;
  assign new_n1430_ = ~new_n838_ & new_n1429_;
  assign new_n1431_ = ~new_n1284_ & new_n1430_;
  assign new_n1432_ = ~new_n1411_ & new_n1431_;
  assign \1_n170  = new_n1409_ | ~new_n1432_;
  assign new_n1434_ = \1_n1121  & new_n799_;
  assign new_n1435_ = new_n801_ & ~new_n1013_;
  assign new_n1436_ = ~new_n1434_ & ~new_n1435_;
  assign new_n1437_ = \1_n1515  & new_n819_;
  assign new_n1438_ = new_n821_ & ~new_n1213_;
  assign new_n1439_ = ~new_n1437_ & ~new_n1438_;
  assign new_n1440_ = new_n1436_ & new_n1439_;
  assign \1_n172  = \1_n24 ;
  assign new_n1442_ = \1_n230  & \1_n1058 ;
  assign new_n1443_ = \1_n365  & ~\1_n1058 ;
  assign new_n1444_ = ~new_n1442_ & ~new_n1443_;
  assign new_n1445_ = \1_n403  & ~new_n1444_;
  assign new_n1446_ = ~\1_n1058  & ~\1_n1255 ;
  assign new_n1447_ = \1_n1058  & ~\1_n1425 ;
  assign new_n1448_ = ~new_n1446_ & ~new_n1447_;
  assign new_n1449_ = ~\1_n403  & ~new_n1448_;
  assign new_n1450_ = ~new_n1445_ & ~new_n1449_;
  assign new_n1451_ = ~\1_n646  & ~\1_n1255 ;
  assign new_n1452_ = \1_n646  & ~\1_n1425 ;
  assign new_n1453_ = ~new_n1451_ & ~new_n1452_;
  assign new_n1454_ = ~\1_n1378  & ~new_n1453_;
  assign new_n1455_ = \1_n365  & ~\1_n646 ;
  assign new_n1456_ = \1_n230  & \1_n646 ;
  assign new_n1457_ = ~new_n1455_ & ~new_n1456_;
  assign new_n1458_ = \1_n1378  & ~new_n1457_;
  assign new_n1459_ = ~new_n1454_ & ~new_n1458_;
  assign new_n1460_ = new_n804_ & new_n1459_;
  assign new_n1461_ = new_n1299_ & new_n1460_;
  assign new_n1462_ = new_n1450_ & new_n1461_;
  assign new_n1463_ = ~new_n895_ & new_n1462_;
  assign new_n1464_ = ~new_n850_ & new_n1463_;
  assign new_n1465_ = new_n862_ & new_n1464_;
  assign new_n1466_ = new_n871_ & new_n1465_;
  assign \1_n190  = ~new_n719_ | ~new_n1466_;
  assign new_n1468_ = ~\1_n362  & new_n1260_;
  assign new_n1469_ = ~\1_n1645  & new_n1262_;
  assign new_n1470_ = ~new_n1468_ & ~new_n1469_;
  assign new_n1471_ = ~\1_n526  & new_n1255_;
  assign new_n1472_ = ~\1_n1478  & new_n1257_;
  assign new_n1473_ = ~new_n1471_ & ~new_n1472_;
  assign \1_n204  = ~new_n1470_ | ~new_n1473_;
  assign new_n1475_ = \1_n635  & new_n606_;
  assign new_n1476_ = new_n617_ & ~new_n1459_;
  assign new_n1477_ = ~new_n1475_ & ~new_n1476_;
  assign new_n1478_ = new_n708_ & ~new_n1222_;
  assign \1_n210  = ~new_n1477_ | new_n1478_;
  assign new_n1480_ = ~\1_n1014  & new_n1255_;
  assign new_n1481_ = \1_n1620  & new_n606_;
  assign new_n1482_ = new_n617_ & ~new_n1450_;
  assign new_n1483_ = ~new_n1481_ & ~new_n1482_;
  assign new_n1484_ = new_n708_ & new_n1235_;
  assign \1_n1665  = ~new_n1483_ | new_n1484_;
  assign new_n1486_ = new_n1257_ & ~\1_n1665 ;
  assign new_n1487_ = ~new_n1480_ & ~new_n1486_;
  assign new_n1488_ = ~\1_n596  & new_n1260_;
  assign new_n1489_ = \1_n432  & new_n606_;
  assign new_n1490_ = new_n617_ & ~new_n1346_;
  assign new_n1491_ = ~new_n1489_ & ~new_n1490_;
  assign new_n1492_ = new_n708_ & new_n1415_;
  assign \1_n1039  = ~new_n1491_ | new_n1492_;
  assign new_n1494_ = new_n1262_ & ~\1_n1039 ;
  assign new_n1495_ = ~new_n1488_ & ~new_n1494_;
  assign \1_n231  = ~new_n1487_ | ~new_n1495_;
  assign new_n1497_ = ~new_n781_ & new_n787_;
  assign new_n1498_ = new_n979_ & ~new_n1497_;
  assign \1_n232  = new_n724_ & new_n1498_;
  assign new_n1500_ = ~\1_n289  & new_n799_;
  assign new_n1501_ = \1_n1131  & new_n606_;
  assign new_n1502_ = new_n617_ & ~new_n871_;
  assign new_n1503_ = ~new_n1501_ & ~new_n1502_;
  assign new_n1504_ = new_n708_ & ~new_n1243_;
  assign \1_n640  = ~new_n1503_ | new_n1504_;
  assign new_n1506_ = new_n801_ & ~\1_n640 ;
  assign new_n1507_ = ~new_n1500_ & ~new_n1506_;
  assign new_n1508_ = ~\1_n1485  & new_n819_;
  assign new_n1509_ = \1_n973  & new_n606_;
  assign new_n1510_ = new_n617_ & ~new_n1364_;
  assign new_n1511_ = ~new_n1509_ & ~new_n1510_;
  assign new_n1512_ = new_n708_ & new_n1420_;
  assign \1_n964  = ~new_n1511_ | new_n1512_;
  assign new_n1514_ = new_n821_ & ~\1_n964 ;
  assign new_n1515_ = ~new_n1508_ & ~new_n1514_;
  assign new_n1516_ = new_n1507_ & new_n1515_;
  assign \1_n240  = \1_n24 ;
  assign \1_n265  = ~\1_n220  | \1_n797 ;
  assign new_n1519_ = ~\1_n290  & new_n1255_;
  assign new_n1520_ = new_n1257_ & ~\1_n434 ;
  assign new_n1521_ = ~new_n1519_ & ~new_n1520_;
  assign new_n1522_ = ~\1_n818  & new_n1260_;
  assign new_n1523_ = new_n1262_ & ~\1_n675 ;
  assign new_n1524_ = ~new_n1522_ & ~new_n1523_;
  assign \1_n269  = ~new_n1521_ | ~new_n1524_;
  assign new_n1526_ = \1_n716  & new_n606_;
  assign new_n1527_ = new_n617_ & new_n895_;
  assign new_n1528_ = ~new_n1526_ & ~new_n1527_;
  assign new_n1529_ = new_n708_ & new_n1225_;
  assign \1_n291  = ~new_n1528_ | new_n1529_;
  assign new_n1531_ = ~\1_n1146  & new_n845_;
  assign new_n1532_ = new_n1014_ & ~\1_n434 ;
  assign new_n1533_ = ~new_n1531_ & ~new_n1532_;
  assign new_n1534_ = ~\1_n1398  & new_n1017_;
  assign new_n1535_ = new_n1214_ & ~\1_n675 ;
  assign new_n1536_ = ~new_n1534_ & ~new_n1535_;
  assign new_n1537_ = new_n1533_ & new_n1536_;
  assign \1_n313  = \1_n24 ;
  assign new_n1539_ = \1_n1508  & new_n606_;
  assign new_n1540_ = new_n617_ & ~new_n1373_;
  assign new_n1541_ = ~new_n1539_ & ~new_n1540_;
  assign new_n1542_ = new_n708_ & ~new_n1425_;
  assign \1_n336  = ~new_n1541_ | new_n1542_;
  assign new_n1544_ = ~\1_n386  & new_n799_;
  assign new_n1545_ = new_n801_ & ~\1_n1665 ;
  assign new_n1546_ = ~new_n1544_ & ~new_n1545_;
  assign new_n1547_ = ~\1_n605  & new_n819_;
  assign new_n1548_ = new_n821_ & ~\1_n1039 ;
  assign new_n1549_ = ~new_n1547_ & ~new_n1548_;
  assign new_n1550_ = new_n1546_ & new_n1549_;
  assign \1_n347  = \1_n24 ;
  assign new_n1552_ = \1_n1276  & \1_n1396 ;
  assign new_n1553_ = \1_n120  & ~\1_n664 ;
  assign new_n1554_ = ~\1_n120  & new_n719_;
  assign new_n1555_ = ~new_n1553_ & ~new_n1554_;
  assign new_n1556_ = ~\1_n869  & ~new_n1555_;
  assign new_n1557_ = ~new_n1552_ & ~new_n1556_;
  assign new_n1558_ = \1_n835  & new_n724_;
  assign new_n1559_ = ~\1_n835  & ~new_n724_;
  assign new_n1560_ = ~new_n1558_ & ~new_n1559_;
  assign new_n1561_ = ~\1_n120  & ~new_n1560_;
  assign new_n1562_ = \1_n120  & ~\1_n693 ;
  assign new_n1563_ = ~new_n1561_ & ~new_n1562_;
  assign new_n1564_ = \1_n869  & ~new_n1563_;
  assign \1_n363  = ~new_n1557_ | new_n1564_;
  assign new_n1566_ = ~\1_n693  & new_n1560_;
  assign new_n1567_ = \1_n693  & ~new_n1560_;
  assign \1_n368  = ~new_n1566_ & ~new_n1567_;
  assign new_n1569_ = ~\1_n514  & \1_n167 ;
  assign new_n1570_ = \1_n576  & new_n1569_;
  assign new_n1571_ = \1_n514  & \1_n167 ;
  assign new_n1572_ = \1_n1052  & new_n1571_;
  assign \1_n383  = new_n1570_ | new_n1572_;
  assign new_n1574_ = ~\1_n9  & new_n713_;
  assign new_n1575_ = new_n715_ & ~\1_n1157 ;
  assign new_n1576_ = ~new_n1574_ & ~new_n1575_;
  assign new_n1577_ = ~\1_n1162  & new_n603_;
  assign new_n1578_ = new_n605_ & ~\1_n928 ;
  assign new_n1579_ = ~new_n1577_ & ~new_n1578_;
  assign \1_n427  = ~new_n1576_ | ~new_n1579_;
  assign new_n1581_ = ~\1_n386  & new_n845_;
  assign new_n1582_ = new_n1014_ & ~\1_n1665 ;
  assign new_n1583_ = ~new_n1581_ & ~new_n1582_;
  assign new_n1584_ = ~\1_n605  & new_n1017_;
  assign new_n1585_ = new_n1214_ & ~\1_n1039 ;
  assign new_n1586_ = ~new_n1584_ & ~new_n1585_;
  assign new_n1587_ = new_n1583_ & new_n1586_;
  assign \1_n506  = \1_n24 ;
  assign new_n1589_ = ~\1_n1091  & new_n819_;
  assign new_n1590_ = ~\1_n1645  & new_n821_;
  assign new_n1591_ = ~new_n1589_ & ~new_n1590_;
  assign new_n1592_ = ~\1_n418  & new_n799_;
  assign new_n1593_ = ~\1_n1478  & new_n801_;
  assign new_n1594_ = ~new_n1592_ & ~new_n1593_;
  assign new_n1595_ = new_n1591_ & new_n1594_;
  assign \1_n524  = \1_n24 ;
  assign new_n1597_ = ~\1_n1511  & new_n1017_;
  assign new_n1598_ = new_n1214_ & ~\1_n1589 ;
  assign new_n1599_ = ~new_n1597_ & ~new_n1598_;
  assign new_n1600_ = ~\1_n909  & new_n845_;
  assign new_n1601_ = new_n1014_ & ~\1_n1177 ;
  assign new_n1602_ = ~new_n1600_ & ~new_n1601_;
  assign new_n1603_ = new_n1599_ & new_n1602_;
  assign \1_n543  = \1_n24 ;
  assign new_n1605_ = ~\1_n1366  & new_n606_;
  assign \1_n598  = ~new_n1212_ | new_n1605_;
  assign new_n1607_ = new_n647_ & new_n693_;
  assign new_n1608_ = ~new_n653_ & ~new_n1607_;
  assign new_n1609_ = ~new_n625_ & new_n1608_;
  assign new_n1610_ = \1_n1240  & ~new_n622_;
  assign \1_n623  = ~new_n1609_ & ~new_n1610_;
  assign new_n1612_ = ~\1_n596  & new_n713_;
  assign new_n1613_ = new_n715_ & ~\1_n1665 ;
  assign new_n1614_ = ~new_n1612_ & ~new_n1613_;
  assign new_n1615_ = ~\1_n1014  & new_n603_;
  assign new_n1616_ = new_n605_ & ~\1_n1039 ;
  assign new_n1617_ = ~new_n1615_ & ~new_n1616_;
  assign \1_n633  = ~new_n1614_ | ~new_n1617_;
  assign new_n1619_ = ~new_n730_ & new_n734_;
  assign new_n1620_ = new_n730_ & ~new_n734_;
  assign new_n1621_ = ~new_n1619_ & ~new_n1620_;
  assign new_n1622_ = ~new_n973_ & new_n1621_;
  assign new_n1623_ = new_n973_ & ~new_n1621_;
  assign new_n1624_ = ~new_n1622_ & ~new_n1623_;
  assign new_n1625_ = ~new_n741_ & ~new_n761_;
  assign new_n1626_ = new_n741_ & new_n761_;
  assign new_n1627_ = ~new_n1625_ & ~new_n1626_;
  assign new_n1628_ = \1_n588  & \1_n1606 ;
  assign new_n1629_ = \1_n1575  & ~\1_n1606 ;
  assign new_n1630_ = ~new_n1628_ & ~new_n1629_;
  assign new_n1631_ = ~new_n768_ & new_n1630_;
  assign new_n1632_ = new_n768_ & ~new_n1630_;
  assign new_n1633_ = ~new_n1631_ & ~new_n1632_;
  assign new_n1634_ = new_n747_ & ~new_n753_;
  assign new_n1635_ = ~new_n747_ & new_n753_;
  assign new_n1636_ = ~new_n1634_ & ~new_n1635_;
  assign new_n1637_ = ~new_n1633_ & new_n1636_;
  assign new_n1638_ = new_n1633_ & ~new_n1636_;
  assign new_n1639_ = ~new_n1637_ & ~new_n1638_;
  assign new_n1640_ = ~new_n1627_ & new_n1639_;
  assign new_n1641_ = new_n1627_ & ~new_n1639_;
  assign new_n1642_ = ~new_n1640_ & ~new_n1641_;
  assign new_n1643_ = new_n1624_ & new_n1642_;
  assign new_n1644_ = ~new_n1624_ & ~new_n1642_;
  assign \1_n656  = new_n1643_ | new_n1644_;
  assign new_n1646_ = ~new_n622_ & new_n628_;
  assign new_n1647_ = new_n622_ & ~new_n628_;
  assign new_n1648_ = ~new_n1646_ & ~new_n1647_;
  assign new_n1649_ = ~new_n634_ & new_n638_;
  assign new_n1650_ = new_n634_ & ~new_n638_;
  assign new_n1651_ = ~new_n1649_ & ~new_n1650_;
  assign new_n1652_ = ~new_n1648_ & new_n1651_;
  assign new_n1653_ = new_n1648_ & ~new_n1651_;
  assign new_n1654_ = ~new_n1652_ & ~new_n1653_;
  assign new_n1655_ = ~new_n656_ & new_n662_;
  assign new_n1656_ = new_n656_ & ~new_n662_;
  assign new_n1657_ = ~new_n1655_ & ~new_n1656_;
  assign new_n1658_ = \1_n1243  & \1_n1253 ;
  assign new_n1659_ = \1_n268  & ~\1_n1243 ;
  assign new_n1660_ = ~new_n1658_ & ~new_n1659_;
  assign new_n1661_ = new_n677_ & ~new_n1660_;
  assign new_n1662_ = ~new_n677_ & new_n1660_;
  assign new_n1663_ = ~new_n1661_ & ~new_n1662_;
  assign new_n1664_ = ~new_n669_ & new_n673_;
  assign new_n1665_ = new_n669_ & ~new_n673_;
  assign new_n1666_ = ~new_n1664_ & ~new_n1665_;
  assign new_n1667_ = ~new_n1663_ & new_n1666_;
  assign new_n1668_ = new_n1663_ & ~new_n1666_;
  assign new_n1669_ = ~new_n1667_ & ~new_n1668_;
  assign new_n1670_ = ~new_n1657_ & new_n1669_;
  assign new_n1671_ = new_n1657_ & ~new_n1669_;
  assign new_n1672_ = ~new_n1670_ & ~new_n1671_;
  assign new_n1673_ = ~new_n1654_ & new_n1672_;
  assign new_n1674_ = new_n1654_ & ~new_n1672_;
  assign \1_n676  = ~new_n1673_ & ~new_n1674_;
  assign new_n1676_ = ~\1_n1184  & new_n713_;
  assign new_n1677_ = new_n715_ & ~\1_n291 ;
  assign new_n1678_ = ~new_n1676_ & ~new_n1677_;
  assign new_n1679_ = ~\1_n1361  & new_n603_;
  assign new_n1680_ = \1_n1339  & new_n606_;
  assign new_n1681_ = new_n617_ & ~new_n1337_;
  assign new_n1682_ = ~new_n1680_ & ~new_n1681_;
  assign new_n1683_ = new_n708_ & new_n1411_;
  assign \1_n1601  = ~new_n1682_ | new_n1683_;
  assign new_n1685_ = new_n605_ & ~\1_n1601 ;
  assign new_n1686_ = ~new_n1679_ & ~new_n1685_;
  assign \1_n691  = ~new_n1678_ | ~new_n1686_;
  assign new_n1688_ = \1_n145  & new_n606_;
  assign new_n1689_ = new_n617_ & new_n850_;
  assign new_n1690_ = ~new_n1688_ & ~new_n1689_;
  assign new_n1691_ = new_n708_ & new_n1246_;
  assign \1_n722  = ~new_n1690_ | new_n1691_;
  assign new_n1693_ = \1_n1648  & new_n1569_;
  assign new_n1694_ = \1_n1549  & new_n1571_;
  assign \1_n1026  = new_n1693_ | new_n1694_;
  assign new_n1696_ = \1_n677  & ~\1_n859 ;
  assign new_n1697_ = ~\1_n677  & \1_n859 ;
  assign new_n1698_ = ~new_n1696_ & ~new_n1697_;
  assign new_n1699_ = ~\1_n135  & \1_n824 ;
  assign new_n1700_ = \1_n135  & ~\1_n824 ;
  assign new_n1701_ = ~new_n1699_ & ~new_n1700_;
  assign new_n1702_ = ~new_n1698_ & new_n1701_;
  assign new_n1703_ = new_n1698_ & ~new_n1701_;
  assign new_n1704_ = ~new_n1702_ & ~new_n1703_;
  assign new_n1705_ = ~\1_n956  & \1_n1143 ;
  assign new_n1706_ = \1_n956  & ~\1_n1143 ;
  assign new_n1707_ = ~new_n1705_ & ~new_n1706_;
  assign new_n1708_ = ~\1_n1030  & \1_n1251 ;
  assign new_n1709_ = \1_n1030  & ~\1_n1251 ;
  assign new_n1710_ = ~new_n1708_ & ~new_n1709_;
  assign new_n1711_ = \1_n209  & ~\1_n268 ;
  assign new_n1712_ = ~\1_n209  & \1_n268 ;
  assign new_n1713_ = ~new_n1711_ & ~new_n1712_;
  assign new_n1714_ = ~new_n1710_ & new_n1713_;
  assign new_n1715_ = new_n1710_ & ~new_n1713_;
  assign new_n1716_ = ~new_n1714_ & ~new_n1715_;
  assign new_n1717_ = ~new_n1707_ & new_n1716_;
  assign new_n1718_ = new_n1707_ & ~new_n1716_;
  assign new_n1719_ = ~new_n1717_ & ~new_n1718_;
  assign new_n1720_ = ~new_n1704_ & new_n1719_;
  assign new_n1721_ = new_n1704_ & ~new_n1719_;
  assign \1_n785  = ~new_n1720_ & ~new_n1721_;
  assign \1_n790  = ~\1_n128  | ~\1_n1562 ;
  assign new_n1724_ = ~\1_n793  & new_n713_;
  assign new_n1725_ = new_n715_ & ~\1_n210 ;
  assign new_n1726_ = ~new_n1724_ & ~new_n1725_;
  assign new_n1727_ = ~\1_n1676  & new_n603_;
  assign new_n1728_ = \1_n1303  & new_n606_;
  assign new_n1729_ = new_n617_ & ~new_n1328_;
  assign new_n1730_ = ~new_n1728_ & ~new_n1729_;
  assign new_n1731_ = new_n708_ & new_n1409_;
  assign \1_n887  = ~new_n1730_ | new_n1731_;
  assign new_n1733_ = new_n605_ & ~\1_n887 ;
  assign new_n1734_ = ~new_n1727_ & ~new_n1733_;
  assign \1_n814  = ~new_n1726_ | ~new_n1734_;
  assign new_n1736_ = ~\1_n222  & new_n606_;
  assign \1_n821  = ~new_n1012_ | new_n1736_;
  assign new_n1738_ = ~\1_n704  & new_n1569_;
  assign new_n1739_ = ~\1_n1438  & new_n1571_;
  assign new_n1740_ = ~new_n1738_ & ~new_n1739_;
  assign \1_n836  = ~\1_n1150  | ~new_n1740_;
  assign new_n1742_ = ~\1_n851  & new_n819_;
  assign new_n1743_ = new_n821_ & ~\1_n336 ;
  assign new_n1744_ = ~new_n1742_ & ~new_n1743_;
  assign new_n1745_ = ~\1_n615  & new_n799_;
  assign new_n1746_ = new_n801_ & ~\1_n722 ;
  assign new_n1747_ = ~new_n1745_ & ~new_n1746_;
  assign new_n1748_ = new_n1744_ & new_n1747_;
  assign \1_n840  = \1_n24 ;
  assign new_n1750_ = ~\1_n710  & new_n799_;
  assign new_n1751_ = new_n801_ & ~\1_n291 ;
  assign new_n1752_ = ~new_n1750_ & ~new_n1751_;
  assign new_n1753_ = ~\1_n1187  & new_n819_;
  assign new_n1754_ = new_n821_ & ~\1_n1601 ;
  assign new_n1755_ = ~new_n1753_ & ~new_n1754_;
  assign new_n1756_ = new_n1752_ & new_n1755_;
  assign \1_n894  = \1_n24 ;
  assign \1_n1032  = ~\1_n293  | ~\1_n750 ;
  assign \1_n1631  = \1_n296  & \1_n1409 ;
  assign new_n1760_ = ~\1_n1032  & \1_n1631 ;
  assign new_n1761_ = \1_n629  & ~\1_n1335 ;
  assign new_n1762_ = ~\1_n629  & \1_n1335 ;
  assign new_n1763_ = ~new_n1761_ & ~new_n1762_;
  assign new_n1764_ = \1_n490  & ~\1_n654 ;
  assign new_n1765_ = ~\1_n490  & \1_n654 ;
  assign new_n1766_ = ~new_n1764_ & ~new_n1765_;
  assign new_n1767_ = ~new_n1763_ & new_n1766_;
  assign new_n1768_ = new_n1763_ & ~new_n1766_;
  assign new_n1769_ = ~new_n1767_ & ~new_n1768_;
  assign new_n1770_ = ~\1_n646  & \1_n1518 ;
  assign new_n1771_ = \1_n646  & ~\1_n1518 ;
  assign new_n1772_ = ~new_n1770_ & ~new_n1771_;
  assign new_n1773_ = \1_n1161  & ~\1_n1575 ;
  assign new_n1774_ = ~\1_n1161  & \1_n1575 ;
  assign new_n1775_ = ~new_n1773_ & ~new_n1774_;
  assign new_n1776_ = ~new_n1772_ & new_n1775_;
  assign new_n1777_ = new_n1772_ & ~new_n1775_;
  assign new_n1778_ = ~new_n1776_ & ~new_n1777_;
  assign new_n1779_ = \1_n1058  & ~new_n1778_;
  assign new_n1780_ = ~\1_n1058  & new_n1778_;
  assign new_n1781_ = ~new_n1779_ & ~new_n1780_;
  assign new_n1782_ = ~new_n1769_ & new_n1781_;
  assign new_n1783_ = new_n1769_ & ~new_n1781_;
  assign \1_n1411  = ~new_n1782_ & ~new_n1783_;
  assign new_n1785_ = new_n1760_ & \1_n1411 ;
  assign new_n1786_ = \1_n785  & new_n1785_;
  assign new_n1787_ = \1_n656  & new_n1786_;
  assign new_n1788_ = \1_n676  & new_n1787_;
  assign new_n1789_ = \1_n1630  & new_n1788_;
  assign \1_n1019  = ~\1_n829  | ~new_n1789_;
  assign new_n1791_ = ~\1_n330  & new_n1569_;
  assign new_n1792_ = ~\1_n990  & new_n1571_;
  assign new_n1793_ = ~new_n1791_ & ~new_n1792_;
  assign \1_n1021  = \1_n836 ;
  assign new_n1795_ = ~\1_n1676  & new_n1255_;
  assign new_n1796_ = new_n1257_ & ~\1_n210 ;
  assign new_n1797_ = ~new_n1795_ & ~new_n1796_;
  assign new_n1798_ = ~\1_n793  & new_n1260_;
  assign new_n1799_ = new_n1262_ & ~\1_n887 ;
  assign new_n1800_ = ~new_n1798_ & ~new_n1799_;
  assign \1_n1036  = ~new_n1797_ | ~new_n1800_;
  assign new_n1802_ = ~\1_n710  & new_n845_;
  assign new_n1803_ = new_n1014_ & ~\1_n291 ;
  assign new_n1804_ = ~new_n1802_ & ~new_n1803_;
  assign new_n1805_ = ~\1_n1187  & new_n1017_;
  assign new_n1806_ = new_n1214_ & ~\1_n1601 ;
  assign new_n1807_ = ~new_n1805_ & ~new_n1806_;
  assign new_n1808_ = new_n1804_ & new_n1807_;
  assign \1_n1043  = \1_n24 ;
  assign new_n1810_ = ~\1_n1361  & new_n1255_;
  assign new_n1811_ = new_n1257_ & ~\1_n291 ;
  assign new_n1812_ = ~new_n1810_ & ~new_n1811_;
  assign new_n1813_ = ~\1_n1184  & new_n1260_;
  assign new_n1814_ = new_n1262_ & ~\1_n1601 ;
  assign new_n1815_ = ~new_n1813_ & ~new_n1814_;
  assign \1_n1122  = ~new_n1812_ | ~new_n1815_;
  assign new_n1817_ = ~\1_n342  & new_n799_;
  assign new_n1818_ = new_n801_ & ~\1_n210 ;
  assign new_n1819_ = ~new_n1817_ & ~new_n1818_;
  assign new_n1820_ = ~\1_n1093  & new_n819_;
  assign new_n1821_ = new_n821_ & ~\1_n887 ;
  assign new_n1822_ = ~new_n1820_ & ~new_n1821_;
  assign new_n1823_ = new_n1819_ & new_n1822_;
  assign \1_n1138  = \1_n24 ;
  assign new_n1825_ = ~\1_n1373  & new_n603_;
  assign new_n1826_ = new_n605_ & ~\1_n336 ;
  assign new_n1827_ = ~new_n1825_ & ~new_n1826_;
  assign new_n1828_ = ~\1_n67  & new_n713_;
  assign new_n1829_ = new_n715_ & ~\1_n722 ;
  assign new_n1830_ = ~new_n1828_ & ~new_n1829_;
  assign \1_n1151  = ~new_n1827_ | ~new_n1830_;
  assign new_n1832_ = ~\1_n289  & new_n845_;
  assign new_n1833_ = new_n1014_ & ~\1_n640 ;
  assign new_n1834_ = ~new_n1832_ & ~new_n1833_;
  assign new_n1835_ = ~\1_n1485  & new_n1017_;
  assign new_n1836_ = new_n1214_ & ~\1_n964 ;
  assign new_n1837_ = ~new_n1835_ & ~new_n1836_;
  assign new_n1838_ = new_n1834_ & new_n1837_;
  assign \1_n1160  = \1_n24 ;
  assign new_n1840_ = ~\1_n342  & new_n845_;
  assign new_n1841_ = new_n1014_ & ~\1_n210 ;
  assign new_n1842_ = ~new_n1840_ & ~new_n1841_;
  assign new_n1843_ = ~\1_n1093  & new_n1017_;
  assign new_n1844_ = new_n1214_ & ~\1_n887 ;
  assign new_n1845_ = ~new_n1843_ & ~new_n1844_;
  assign new_n1846_ = new_n1842_ & new_n1845_;
  assign \1_n1194  = \1_n24 ;
  assign new_n1848_ = ~\1_n1042  & new_n603_;
  assign new_n1849_ = new_n605_ & ~\1_n1589 ;
  assign new_n1850_ = ~new_n1848_ & ~new_n1849_;
  assign new_n1851_ = ~\1_n933  & new_n713_;
  assign new_n1852_ = new_n715_ & ~\1_n1177 ;
  assign new_n1853_ = ~new_n1851_ & ~new_n1852_;
  assign \1_n1198  = ~new_n1850_ | ~new_n1853_;
  assign new_n1855_ = ~\1_n1070  & new_n1569_;
  assign new_n1856_ = ~\1_n1422  & new_n1571_;
  assign new_n1857_ = ~new_n1855_ & ~new_n1856_;
  assign \1_n1239  = \1_n836 ;
  assign new_n1859_ = ~\1_n818  & new_n713_;
  assign new_n1860_ = new_n715_ & ~\1_n434 ;
  assign new_n1861_ = ~new_n1859_ & ~new_n1860_;
  assign new_n1862_ = ~\1_n290  & new_n603_;
  assign new_n1863_ = new_n605_ & ~\1_n675 ;
  assign new_n1864_ = ~new_n1862_ & ~new_n1863_;
  assign \1_n1275  = ~new_n1861_ | ~new_n1864_;
  assign new_n1866_ = ~\1_n1162  & new_n1255_;
  assign new_n1867_ = ~\1_n1157  & new_n1257_;
  assign new_n1868_ = ~new_n1866_ & ~new_n1867_;
  assign new_n1869_ = ~\1_n9  & new_n1260_;
  assign new_n1870_ = ~\1_n928  & new_n1262_;
  assign new_n1871_ = ~new_n1869_ & ~new_n1870_;
  assign \1_n1314  = ~new_n1868_ | ~new_n1871_;
  assign new_n1873_ = ~\1_n468  & new_n845_;
  assign new_n1874_ = ~\1_n1157  & new_n1014_;
  assign new_n1875_ = ~new_n1873_ & ~new_n1874_;
  assign new_n1876_ = ~\1_n934  & new_n1017_;
  assign new_n1877_ = ~\1_n928  & new_n1214_;
  assign new_n1878_ = ~new_n1876_ & ~new_n1877_;
  assign new_n1879_ = new_n1875_ & new_n1878_;
  assign \1_n1375  = \1_n24 ;
  assign new_n1881_ = ~\1_n67  & new_n1260_;
  assign new_n1882_ = new_n1262_ & ~\1_n336 ;
  assign new_n1883_ = ~new_n1881_ & ~new_n1882_;
  assign new_n1884_ = ~\1_n1373  & new_n1255_;
  assign new_n1885_ = new_n1257_ & ~\1_n722 ;
  assign new_n1886_ = ~new_n1884_ & ~new_n1885_;
  assign \1_n1392  = ~new_n1883_ | ~new_n1886_;
  assign \1_n1454  = ~\1_n1099  & \1_n1412 ;
  assign new_n1889_ = ~\1_n1091  & new_n1017_;
  assign new_n1890_ = ~\1_n1645  & new_n1214_;
  assign new_n1891_ = ~new_n1889_ & ~new_n1890_;
  assign new_n1892_ = ~\1_n418  & new_n845_;
  assign new_n1893_ = ~\1_n1478  & new_n1014_;
  assign new_n1894_ = ~new_n1892_ & ~new_n1893_;
  assign new_n1895_ = new_n1891_ & new_n1894_;
  assign \1_n1474  = \1_n24 ;
  assign new_n1897_ = ~\1_n1581  & new_n1255_;
  assign new_n1898_ = new_n1257_ & ~\1_n640 ;
  assign new_n1899_ = ~new_n1897_ & ~new_n1898_;
  assign new_n1900_ = ~\1_n848  & new_n1260_;
  assign new_n1901_ = new_n1262_ & ~\1_n964 ;
  assign new_n1902_ = ~new_n1900_ & ~new_n1901_;
  assign \1_n1512  = ~new_n1899_ | ~new_n1902_;
  assign new_n1904_ = ~\1_n1098  & new_n1569_;
  assign new_n1905_ = ~\1_n974  & new_n1571_;
  assign new_n1906_ = ~new_n1904_ & ~new_n1905_;
  assign \1_n1531  = \1_n836 ;
  assign \1_n1574  = ~\1_n96  | ~\1_n1150 ;
  assign new_n1909_ = ~\1_n1280  & new_n713_;
  assign new_n1910_ = new_n715_ & new_n1013_;
  assign new_n1911_ = ~new_n1909_ & ~new_n1910_;
  assign new_n1912_ = ~\1_n923  & new_n603_;
  assign new_n1913_ = new_n605_ & new_n1213_;
  assign new_n1914_ = ~new_n1912_ & ~new_n1913_;
  assign \1_n1594  = ~new_n1911_ | ~new_n1914_;
  assign new_n1916_ = ~\1_n851  & new_n1017_;
  assign new_n1917_ = new_n1214_ & ~\1_n336 ;
  assign new_n1918_ = ~new_n1916_ & ~new_n1917_;
  assign new_n1919_ = ~\1_n615  & new_n845_;
  assign new_n1920_ = new_n1014_ & ~\1_n722 ;
  assign new_n1921_ = ~new_n1919_ & ~new_n1920_;
  assign new_n1922_ = new_n1918_ & new_n1921_;
  assign \1_n1604  = \1_n24 ;
  assign \1_n1628  = \1_n794  & \1_n167 ;
  assign new_n1925_ = ~\1_n848  & new_n713_;
  assign new_n1926_ = new_n715_ & ~\1_n640 ;
  assign new_n1927_ = ~new_n1925_ & ~new_n1926_;
  assign new_n1928_ = ~\1_n1581  & new_n603_;
  assign new_n1929_ = new_n605_ & ~\1_n964 ;
  assign new_n1930_ = ~new_n1928_ & ~new_n1929_;
  assign \1_n1671  = ~new_n1927_ | ~new_n1930_;
  assign new_n1932_ = \2_n186  & \2_n754 ;
  assign new_n1933_ = \2_n560  & new_n1932_;
  assign new_n1934_ = \2_n1177  & \2_n186 ;
  assign new_n1935_ = ~\2_n560  & new_n1934_;
  assign new_n1936_ = ~new_n1933_ & ~new_n1935_;
  assign new_n1937_ = \2_n482  & ~\2_n579 ;
  assign new_n1938_ = \2_n261  & new_n1937_;
  assign new_n1939_ = \2_n288  & \2_n807 ;
  assign new_n1940_ = ~\2_n288  & \2_n714 ;
  assign new_n1941_ = ~new_n1939_ & ~new_n1940_;
  assign new_n1942_ = ~\2_n579  & ~new_n1941_;
  assign new_n1943_ = ~\2_n261  & new_n1942_;
  assign new_n1944_ = \2_n600  & \2_n971 ;
  assign new_n1945_ = \2_n1518  & ~\2_n600 ;
  assign new_n1946_ = ~new_n1944_ & ~new_n1945_;
  assign new_n1947_ = \2_n1426  & \2_n600 ;
  assign new_n1948_ = ~\2_n600  & \2_n966 ;
  assign new_n1949_ = ~new_n1947_ & ~new_n1948_;
  assign new_n1950_ = \2_n326  & ~new_n1949_;
  assign new_n1951_ = new_n1946_ & ~new_n1950_;
  assign new_n1952_ = \2_n600  & \2_n894 ;
  assign new_n1953_ = ~\2_n600  & \2_n946 ;
  assign new_n1954_ = ~new_n1952_ & ~new_n1953_;
  assign new_n1955_ = \2_n1406  & ~new_n1954_;
  assign new_n1956_ = \2_n326  & new_n1949_;
  assign new_n1957_ = ~\2_n326  & ~new_n1949_;
  assign new_n1958_ = ~new_n1956_ & ~new_n1957_;
  assign new_n1959_ = new_n1955_ & ~new_n1958_;
  assign new_n1960_ = new_n1951_ & ~new_n1959_;
  assign new_n1961_ = \2_n389  & \2_n600 ;
  assign new_n1962_ = \2_n288  & ~\2_n600 ;
  assign new_n1963_ = ~new_n1961_ & ~new_n1962_;
  assign new_n1964_ = new_n1960_ & new_n1963_;
  assign new_n1965_ = ~new_n1960_ & ~new_n1963_;
  assign new_n1966_ = ~new_n1964_ & ~new_n1965_;
  assign new_n1967_ = ~\2_n1568  & \2_n600 ;
  assign new_n1968_ = \2_n238  & ~new_n1967_;
  assign new_n1969_ = ~\2_n238  & new_n1967_;
  assign new_n1970_ = ~new_n1968_ & ~new_n1969_;
  assign new_n1971_ = \2_n1707  & \2_n600 ;
  assign new_n1972_ = \2_n380  & ~\2_n600 ;
  assign new_n1973_ = ~new_n1971_ & ~new_n1972_;
  assign new_n1974_ = \2_n1391  & new_n1973_;
  assign new_n1975_ = ~\2_n1391  & ~new_n1973_;
  assign new_n1976_ = ~new_n1974_ & ~new_n1975_;
  assign new_n1977_ = new_n1970_ & ~new_n1976_;
  assign new_n1978_ = \2_n600  & \2_n937 ;
  assign new_n1979_ = \2_n1435  & ~\2_n600 ;
  assign new_n1980_ = ~new_n1978_ & ~new_n1979_;
  assign new_n1981_ = \2_n1016  & new_n1980_;
  assign new_n1982_ = ~\2_n1016  & ~new_n1980_;
  assign new_n1983_ = ~new_n1981_ & ~new_n1982_;
  assign new_n1984_ = \2_n1338  & \2_n600 ;
  assign new_n1985_ = \2_n1515  & ~\2_n600 ;
  assign new_n1986_ = ~new_n1984_ & ~new_n1985_;
  assign new_n1987_ = \2_n448  & \2_n600 ;
  assign new_n1988_ = \2_n1043  & ~\2_n600 ;
  assign new_n1989_ = ~new_n1987_ & ~new_n1988_;
  assign new_n1990_ = \2_n1125  & new_n1989_;
  assign new_n1991_ = ~\2_n1125  & ~new_n1989_;
  assign new_n1992_ = ~new_n1990_ & ~new_n1991_;
  assign new_n1993_ = new_n1986_ & ~new_n1992_;
  assign new_n1994_ = ~new_n1983_ & new_n1993_;
  assign new_n1995_ = new_n1977_ & new_n1994_;
  assign new_n1996_ = \2_n1788  & new_n1995_;
  assign new_n1997_ = ~new_n1986_ & ~new_n1992_;
  assign new_n1998_ = ~new_n1983_ & new_n1997_;
  assign new_n1999_ = new_n1977_ & new_n1998_;
  assign new_n2000_ = \2_n1391  & ~new_n1973_;
  assign new_n2001_ = new_n1968_ & ~new_n1976_;
  assign new_n2002_ = ~new_n2000_ & ~new_n2001_;
  assign new_n2003_ = \2_n1016  & ~new_n1980_;
  assign new_n2004_ = new_n1970_ & new_n2003_;
  assign new_n2005_ = \2_n1125  & ~new_n1989_;
  assign new_n2006_ = ~new_n1983_ & new_n2005_;
  assign new_n2007_ = new_n1970_ & new_n2006_;
  assign new_n2008_ = ~new_n2004_ & ~new_n2007_;
  assign new_n2009_ = ~new_n1976_ & ~new_n2008_;
  assign new_n2010_ = new_n2002_ & ~new_n2009_;
  assign new_n2011_ = ~new_n1999_ & new_n2010_;
  assign new_n2012_ = ~new_n1996_ & new_n2011_;
  assign new_n2013_ = ~new_n1966_ & new_n2012_;
  assign new_n2014_ = \2_n1406  & new_n1954_;
  assign new_n2015_ = ~\2_n1406  & ~new_n1954_;
  assign new_n2016_ = ~new_n2014_ & ~new_n2015_;
  assign new_n2017_ = ~new_n1958_ & ~new_n2016_;
  assign new_n2018_ = new_n1960_ & ~new_n2017_;
  assign new_n2019_ = ~new_n1963_ & new_n2018_;
  assign new_n2020_ = new_n1963_ & ~new_n2018_;
  assign new_n2021_ = ~new_n2012_ & ~new_n2020_;
  assign new_n2022_ = ~new_n2019_ & new_n2021_;
  assign \2_n1793  = ~new_n2013_ & ~new_n2022_;
  assign new_n2024_ = \2_n579  & ~\2_n1793 ;
  assign new_n2025_ = ~\2_n261  & new_n2024_;
  assign new_n2026_ = ~new_n1943_ & ~new_n2025_;
  assign \2_n1027  = ~new_n1938_ & new_n2026_;
  assign new_n2028_ = ~\2_n186  & ~\2_n1027 ;
  assign new_n2029_ = ~\2_n560  & new_n2028_;
  assign new_n2030_ = ~\2_n579  & \2_n850 ;
  assign new_n2031_ = \2_n261  & new_n2030_;
  assign new_n2032_ = \2_n591  & \2_n708 ;
  assign new_n2033_ = \2_n1227  & ~\2_n708 ;
  assign new_n2034_ = ~new_n2032_ & ~new_n2033_;
  assign new_n2035_ = \2_n60  & ~new_n2034_;
  assign new_n2036_ = \2_n708  & \2_n807 ;
  assign new_n2037_ = ~\2_n708  & \2_n714 ;
  assign new_n2038_ = ~\2_n60  & ~new_n2037_;
  assign new_n2039_ = ~new_n2036_ & new_n2038_;
  assign new_n2040_ = ~new_n2035_ & ~new_n2039_;
  assign new_n2041_ = ~\2_n579  & new_n2040_;
  assign new_n2042_ = ~\2_n261  & new_n2041_;
  assign new_n2043_ = \2_n1408  & \2_n504 ;
  assign new_n2044_ = ~\2_n504  & \2_n708 ;
  assign new_n2045_ = ~new_n2043_ & ~new_n2044_;
  assign new_n2046_ = \2_n60  & new_n2045_;
  assign new_n2047_ = ~\2_n60  & ~new_n2045_;
  assign new_n2048_ = ~new_n2046_ & ~new_n2047_;
  assign new_n2049_ = \2_n504  & \2_n801 ;
  assign new_n2050_ = \2_n1660  & ~\2_n504 ;
  assign new_n2051_ = ~new_n2049_ & ~new_n2050_;
  assign new_n2052_ = \2_n1575  & ~new_n2051_;
  assign new_n2053_ = \2_n1575  & new_n2051_;
  assign new_n2054_ = ~\2_n1575  & ~new_n2051_;
  assign new_n2055_ = ~new_n2053_ & ~new_n2054_;
  assign new_n2056_ = \2_n1485  & \2_n504 ;
  assign new_n2057_ = \2_n1172  & ~\2_n504 ;
  assign new_n2058_ = ~new_n2056_ & ~new_n2057_;
  assign new_n2059_ = \2_n697  & ~new_n2058_;
  assign new_n2060_ = \2_n504  & \2_n917 ;
  assign new_n2061_ = \2_n1553  & ~\2_n504 ;
  assign new_n2062_ = ~new_n2060_ & ~new_n2061_;
  assign new_n2063_ = \2_n1755  & ~new_n2062_;
  assign new_n2064_ = \2_n697  & new_n2058_;
  assign new_n2065_ = ~\2_n697  & ~new_n2058_;
  assign new_n2066_ = ~new_n2064_ & ~new_n2065_;
  assign new_n2067_ = new_n2063_ & ~new_n2066_;
  assign new_n2068_ = ~new_n2059_ & ~new_n2067_;
  assign new_n2069_ = ~new_n2055_ & ~new_n2068_;
  assign new_n2070_ = ~new_n2052_ & ~new_n2069_;
  assign new_n2071_ = new_n2048_ & ~new_n2070_;
  assign new_n2072_ = ~new_n2048_ & new_n2070_;
  assign new_n2073_ = ~new_n2071_ & ~new_n2072_;
  assign new_n2074_ = \2_n1436  & \2_n504 ;
  assign new_n2075_ = \2_n319  & ~\2_n504 ;
  assign new_n2076_ = ~new_n2074_ & ~new_n2075_;
  assign new_n2077_ = \2_n1402  & ~new_n2076_;
  assign new_n2078_ = ~\2_n1402  & new_n2076_;
  assign new_n2079_ = ~new_n2077_ & ~new_n2078_;
  assign new_n2080_ = \2_n504  & \2_n887 ;
  assign new_n2081_ = \2_n1729  & ~\2_n504 ;
  assign new_n2082_ = ~new_n2080_ & ~new_n2081_;
  assign new_n2083_ = \2_n1135  & new_n2082_;
  assign new_n2084_ = ~\2_n1135  & ~new_n2082_;
  assign new_n2085_ = ~new_n2083_ & ~new_n2084_;
  assign new_n2086_ = \2_n504  & \2_n961 ;
  assign new_n2087_ = \2_n1238  & ~\2_n504 ;
  assign new_n2088_ = ~new_n2086_ & ~new_n2087_;
  assign new_n2089_ = \2_n1100  & ~new_n2088_;
  assign new_n2090_ = ~\2_n1100  & new_n2088_;
  assign new_n2091_ = ~new_n2089_ & ~new_n2090_;
  assign new_n2092_ = ~new_n2085_ & new_n2091_;
  assign new_n2093_ = \2_n1632  & \2_n504 ;
  assign new_n2094_ = \2_n1498  & ~\2_n504 ;
  assign new_n2095_ = ~new_n2093_ & ~new_n2094_;
  assign new_n2096_ = \2_n1039  & new_n2095_;
  assign new_n2097_ = ~\2_n1039  & ~new_n2095_;
  assign new_n2098_ = ~new_n2096_ & ~new_n2097_;
  assign new_n2099_ = \2_n1396  & \2_n504 ;
  assign new_n2100_ = ~\2_n504  & \2_n617 ;
  assign new_n2101_ = ~new_n2099_ & ~new_n2100_;
  assign new_n2102_ = \2_n39  & new_n2101_;
  assign new_n2103_ = ~\2_n39  & ~new_n2101_;
  assign new_n2104_ = ~new_n2102_ & ~new_n2103_;
  assign new_n2105_ = ~new_n2098_ & ~new_n2104_;
  assign new_n2106_ = new_n2092_ & new_n2105_;
  assign new_n2107_ = new_n2079_ & new_n2106_;
  assign new_n2108_ = \2_n1279  & new_n2107_;
  assign new_n2109_ = new_n2079_ & ~new_n2085_;
  assign new_n2110_ = \2_n39  & ~new_n2101_;
  assign new_n2111_ = ~new_n2098_ & new_n2110_;
  assign new_n2112_ = new_n2091_ & new_n2111_;
  assign new_n2113_ = new_n2109_ & new_n2112_;
  assign new_n2114_ = \2_n1135  & ~new_n2082_;
  assign new_n2115_ = new_n2077_ & ~new_n2085_;
  assign new_n2116_ = ~new_n2114_ & ~new_n2115_;
  assign new_n2117_ = new_n2079_ & new_n2089_;
  assign new_n2118_ = \2_n1039  & ~new_n2095_;
  assign new_n2119_ = new_n2091_ & new_n2118_;
  assign new_n2120_ = new_n2079_ & new_n2119_;
  assign new_n2121_ = ~new_n2117_ & ~new_n2120_;
  assign new_n2122_ = ~new_n2085_ & ~new_n2121_;
  assign new_n2123_ = new_n2116_ & ~new_n2122_;
  assign new_n2124_ = ~new_n2113_ & new_n2123_;
  assign new_n2125_ = ~new_n2108_ & new_n2124_;
  assign new_n2126_ = ~new_n2073_ & new_n2125_;
  assign new_n2127_ = \2_n1755  & new_n2062_;
  assign new_n2128_ = ~\2_n1755  & ~new_n2062_;
  assign new_n2129_ = ~new_n2127_ & ~new_n2128_;
  assign new_n2130_ = ~new_n2066_ & ~new_n2129_;
  assign new_n2131_ = ~new_n2055_ & new_n2130_;
  assign new_n2132_ = new_n2070_ & ~new_n2131_;
  assign new_n2133_ = ~new_n2048_ & ~new_n2132_;
  assign new_n2134_ = new_n2048_ & new_n2132_;
  assign new_n2135_ = ~new_n2125_ & ~new_n2134_;
  assign new_n2136_ = ~new_n2133_ & new_n2135_;
  assign new_n2137_ = ~new_n2126_ & ~new_n2136_;
  assign new_n2138_ = \2_n579  & ~new_n2137_;
  assign new_n2139_ = ~\2_n261  & new_n2138_;
  assign new_n2140_ = ~new_n2042_ & ~new_n2139_;
  assign \2_n123  = ~new_n2031_ & new_n2140_;
  assign new_n2142_ = ~\2_n186  & ~\2_n123 ;
  assign new_n2143_ = \2_n560  & new_n2142_;
  assign new_n2144_ = ~new_n2029_ & ~new_n2143_;
  assign \2_n101  = ~new_n1936_ | ~new_n2144_;
  assign \2_n1047  = \2_n457  & \2_n92 ;
  assign new_n2147_ = \2_n627  & \2_n7 ;
  assign new_n2148_ = \2_n378  & new_n2147_;
  assign new_n2149_ = \2_n1180  & \2_n627 ;
  assign new_n2150_ = ~\2_n378  & new_n2149_;
  assign new_n2151_ = ~new_n2148_ & ~new_n2150_;
  assign new_n2152_ = ~\2_n579  & \2_n668 ;
  assign new_n2153_ = \2_n261  & new_n2152_;
  assign new_n2154_ = \2_n1043  & \2_n1288 ;
  assign new_n2155_ = ~\2_n1043  & \2_n721 ;
  assign new_n2156_ = \2_n1125  & ~new_n2155_;
  assign new_n2157_ = ~new_n2154_ & new_n2156_;
  assign new_n2158_ = \2_n1043  & \2_n77 ;
  assign new_n2159_ = ~\2_n1043  & \2_n1519 ;
  assign new_n2160_ = ~new_n2158_ & ~new_n2159_;
  assign new_n2161_ = ~\2_n1125  & ~new_n2160_;
  assign new_n2162_ = ~new_n2157_ & ~new_n2161_;
  assign new_n2163_ = ~\2_n579  & new_n2162_;
  assign new_n2164_ = ~\2_n261  & new_n2163_;
  assign new_n2165_ = ~\2_n1788  & new_n1986_;
  assign new_n2166_ = ~new_n1992_ & new_n2165_;
  assign new_n2167_ = new_n1992_ & ~new_n2165_;
  assign new_n2168_ = ~new_n2166_ & ~new_n2167_;
  assign new_n2169_ = \2_n579  & ~new_n2168_;
  assign new_n2170_ = ~\2_n261  & new_n2169_;
  assign new_n2171_ = ~new_n2164_ & ~new_n2170_;
  assign \2_n168  = ~new_n2153_ & new_n2171_;
  assign new_n2173_ = ~\2_n627  & ~\2_n168 ;
  assign new_n2174_ = ~\2_n378  & new_n2173_;
  assign new_n2175_ = \2_n1633  & ~\2_n579 ;
  assign new_n2176_ = \2_n261  & new_n2175_;
  assign new_n2177_ = ~\2_n1288  & \2_n1498 ;
  assign new_n2178_ = ~\2_n1498  & ~\2_n721 ;
  assign new_n2179_ = ~new_n2177_ & ~new_n2178_;
  assign new_n2180_ = \2_n1039  & ~new_n2179_;
  assign new_n2181_ = \2_n1498  & ~\2_n77 ;
  assign new_n2182_ = ~\2_n1498  & ~\2_n1519 ;
  assign new_n2183_ = ~\2_n1039  & ~new_n2182_;
  assign new_n2184_ = ~new_n2181_ & new_n2183_;
  assign new_n2185_ = ~new_n2180_ & ~new_n2184_;
  assign new_n2186_ = ~\2_n579  & new_n2185_;
  assign new_n2187_ = ~\2_n261  & new_n2186_;
  assign new_n2188_ = \2_n1279  & ~new_n2104_;
  assign new_n2189_ = ~new_n2110_ & ~new_n2188_;
  assign new_n2190_ = ~new_n2098_ & ~new_n2189_;
  assign new_n2191_ = new_n2098_ & new_n2189_;
  assign new_n2192_ = ~new_n2190_ & ~new_n2191_;
  assign new_n2193_ = \2_n579  & new_n2192_;
  assign new_n2194_ = ~\2_n261  & new_n2193_;
  assign new_n2195_ = ~new_n2187_ & ~new_n2194_;
  assign \2_n1346  = ~new_n2176_ & new_n2195_;
  assign new_n2197_ = ~\2_n627  & ~\2_n1346 ;
  assign new_n2198_ = \2_n378  & new_n2197_;
  assign new_n2199_ = ~new_n2174_ & ~new_n2198_;
  assign new_n2200_ = new_n2151_ & new_n2199_;
  assign \2_n1050  = \2_n1534  & ~new_n2200_;
  assign new_n2202_ = \2_n1205  & \2_n962 ;
  assign new_n2203_ = \2_n228  & new_n2202_;
  assign new_n2204_ = \2_n1205  & \2_n1663 ;
  assign new_n2205_ = ~\2_n228  & new_n2204_;
  assign new_n2206_ = ~new_n2203_ & ~new_n2205_;
  assign new_n2207_ = \2_n261  & \2_n321 ;
  assign new_n2208_ = ~\2_n591  & \2_n946 ;
  assign new_n2209_ = ~\2_n1227  & ~\2_n946 ;
  assign new_n2210_ = \2_n1406  & ~new_n2209_;
  assign new_n2211_ = ~new_n2208_ & new_n2210_;
  assign new_n2212_ = ~\2_n807  & \2_n946 ;
  assign new_n2213_ = ~\2_n714  & ~\2_n946 ;
  assign new_n2214_ = ~new_n2212_ & ~new_n2213_;
  assign new_n2215_ = ~\2_n1406  & ~new_n2214_;
  assign new_n2216_ = ~new_n2211_ & ~new_n2215_;
  assign new_n2217_ = ~\2_n591  & \2_n966 ;
  assign new_n2218_ = ~\2_n1227  & ~\2_n966 ;
  assign new_n2219_ = \2_n326  & ~new_n2218_;
  assign new_n2220_ = ~new_n2217_ & new_n2219_;
  assign new_n2221_ = ~\2_n807  & \2_n966 ;
  assign new_n2222_ = ~\2_n714  & ~\2_n966 ;
  assign new_n2223_ = ~new_n2221_ & ~new_n2222_;
  assign new_n2224_ = ~\2_n326  & ~new_n2223_;
  assign new_n2225_ = ~new_n2220_ & ~new_n2224_;
  assign new_n2226_ = ~new_n2216_ & new_n2225_;
  assign new_n2227_ = new_n2216_ & ~new_n2225_;
  assign new_n2228_ = ~new_n2226_ & ~new_n2227_;
  assign new_n2229_ = \2_n1518  & \2_n591 ;
  assign new_n2230_ = \2_n1227  & ~\2_n1518 ;
  assign new_n2231_ = ~new_n2229_ & ~new_n2230_;
  assign new_n2232_ = new_n1941_ & new_n2231_;
  assign new_n2233_ = ~new_n1941_ & ~new_n2231_;
  assign new_n2234_ = ~new_n2232_ & ~new_n2233_;
  assign new_n2235_ = ~new_n2228_ & new_n2234_;
  assign new_n2236_ = new_n2228_ & ~new_n2234_;
  assign new_n2237_ = ~new_n2235_ & ~new_n2236_;
  assign new_n2238_ = ~\2_n238  & \2_n807 ;
  assign new_n2239_ = \2_n238  & ~\2_n591 ;
  assign new_n2240_ = ~new_n2238_ & ~new_n2239_;
  assign new_n2241_ = \2_n380  & ~\2_n591 ;
  assign new_n2242_ = ~\2_n1227  & ~\2_n380 ;
  assign new_n2243_ = \2_n1391  & ~new_n2242_;
  assign new_n2244_ = ~new_n2241_ & new_n2243_;
  assign new_n2245_ = \2_n380  & ~\2_n807 ;
  assign new_n2246_ = ~\2_n380  & ~\2_n714 ;
  assign new_n2247_ = ~new_n2245_ & ~new_n2246_;
  assign new_n2248_ = ~\2_n1391  & ~new_n2247_;
  assign new_n2249_ = ~new_n2244_ & ~new_n2248_;
  assign new_n2250_ = ~new_n2240_ & new_n2249_;
  assign new_n2251_ = new_n2240_ & ~new_n2249_;
  assign new_n2252_ = ~new_n2250_ & ~new_n2251_;
  assign new_n2253_ = \2_n1515  & \2_n591 ;
  assign new_n2254_ = \2_n1227  & ~\2_n1515 ;
  assign new_n2255_ = ~new_n2253_ & ~new_n2254_;
  assign new_n2256_ = \2_n1435  & ~\2_n591 ;
  assign new_n2257_ = ~\2_n1227  & ~\2_n1435 ;
  assign new_n2258_ = \2_n1016  & ~new_n2257_;
  assign new_n2259_ = ~new_n2256_ & new_n2258_;
  assign new_n2260_ = \2_n1435  & ~\2_n807 ;
  assign new_n2261_ = ~\2_n1435  & ~\2_n714 ;
  assign new_n2262_ = ~new_n2260_ & ~new_n2261_;
  assign new_n2263_ = ~\2_n1016  & ~new_n2262_;
  assign new_n2264_ = ~new_n2259_ & ~new_n2263_;
  assign new_n2265_ = \2_n1043  & \2_n591 ;
  assign new_n2266_ = ~\2_n1043  & \2_n1227 ;
  assign new_n2267_ = ~new_n2265_ & ~new_n2266_;
  assign new_n2268_ = \2_n1125  & ~new_n2267_;
  assign new_n2269_ = \2_n1043  & \2_n807 ;
  assign new_n2270_ = ~\2_n1043  & \2_n714 ;
  assign new_n2271_ = ~\2_n1125  & ~new_n2270_;
  assign new_n2272_ = ~new_n2269_ & new_n2271_;
  assign new_n2273_ = ~new_n2268_ & ~new_n2272_;
  assign new_n2274_ = ~new_n2264_ & ~new_n2273_;
  assign new_n2275_ = new_n2264_ & new_n2273_;
  assign new_n2276_ = ~new_n2274_ & ~new_n2275_;
  assign new_n2277_ = new_n2255_ & new_n2276_;
  assign new_n2278_ = ~new_n2255_ & ~new_n2276_;
  assign new_n2279_ = ~new_n2277_ & ~new_n2278_;
  assign new_n2280_ = ~new_n2252_ & new_n2279_;
  assign new_n2281_ = new_n2252_ & ~new_n2279_;
  assign new_n2282_ = ~new_n2280_ & ~new_n2281_;
  assign new_n2283_ = ~new_n2237_ & ~new_n2282_;
  assign new_n2284_ = new_n2237_ & new_n2282_;
  assign new_n2285_ = ~\2_n579  & ~new_n2284_;
  assign new_n2286_ = ~new_n2283_ & new_n2285_;
  assign new_n2287_ = new_n1946_ & ~new_n1963_;
  assign new_n2288_ = ~new_n1946_ & new_n1963_;
  assign new_n2289_ = ~new_n2287_ & ~new_n2288_;
  assign new_n2290_ = ~new_n1950_ & ~new_n1959_;
  assign new_n2291_ = ~new_n2289_ & ~new_n2290_;
  assign new_n2292_ = new_n2289_ & new_n2290_;
  assign new_n2293_ = ~new_n2291_ & ~new_n2292_;
  assign new_n2294_ = new_n1958_ & ~new_n2016_;
  assign new_n2295_ = ~new_n1958_ & new_n2016_;
  assign new_n2296_ = ~new_n2294_ & ~new_n2295_;
  assign new_n2297_ = ~new_n1955_ & new_n1960_;
  assign new_n2298_ = new_n1955_ & ~new_n1960_;
  assign new_n2299_ = ~new_n2297_ & ~new_n2298_;
  assign new_n2300_ = ~new_n2296_ & new_n2299_;
  assign new_n2301_ = new_n2296_ & ~new_n2299_;
  assign new_n2302_ = ~new_n2300_ & ~new_n2301_;
  assign new_n2303_ = ~new_n2293_ & new_n2302_;
  assign new_n2304_ = new_n2293_ & ~new_n2302_;
  assign new_n2305_ = ~new_n2303_ & ~new_n2304_;
  assign new_n2306_ = new_n2011_ & new_n2305_;
  assign new_n2307_ = ~\2_n1366  & ~new_n2306_;
  assign new_n2308_ = ~new_n2017_ & new_n2290_;
  assign new_n2309_ = ~new_n2289_ & new_n2308_;
  assign new_n2310_ = new_n2289_ & ~new_n2308_;
  assign new_n2311_ = ~new_n2309_ & ~new_n2310_;
  assign new_n2312_ = ~new_n1955_ & new_n2016_;
  assign new_n2313_ = ~new_n2018_ & ~new_n2312_;
  assign new_n2314_ = new_n2018_ & new_n2312_;
  assign new_n2315_ = ~new_n2313_ & ~new_n2314_;
  assign new_n2316_ = ~new_n2296_ & new_n2315_;
  assign new_n2317_ = new_n2296_ & ~new_n2315_;
  assign new_n2318_ = ~new_n2316_ & ~new_n2317_;
  assign new_n2319_ = ~new_n2311_ & new_n2318_;
  assign new_n2320_ = new_n2311_ & ~new_n2318_;
  assign new_n2321_ = ~new_n2319_ & ~new_n2320_;
  assign new_n2322_ = ~new_n2011_ & new_n2321_;
  assign new_n2323_ = new_n2307_ & ~new_n2322_;
  assign new_n2324_ = ~new_n1995_ & new_n2011_;
  assign new_n2325_ = ~new_n2305_ & new_n2324_;
  assign new_n2326_ = ~new_n2321_ & ~new_n2324_;
  assign new_n2327_ = ~new_n2325_ & ~new_n2326_;
  assign new_n2328_ = \2_n1366  & ~new_n2327_;
  assign new_n2329_ = ~new_n2323_ & ~new_n2328_;
  assign new_n2330_ = ~new_n1997_ & ~new_n2005_;
  assign new_n2331_ = ~new_n2003_ & ~new_n2006_;
  assign new_n2332_ = ~new_n1998_ & new_n2331_;
  assign new_n2333_ = new_n2330_ & new_n2332_;
  assign new_n2334_ = ~new_n2330_ & ~new_n2332_;
  assign new_n2335_ = ~new_n2333_ & ~new_n2334_;
  assign new_n2336_ = ~new_n1970_ & new_n1976_;
  assign new_n2337_ = ~new_n1977_ & ~new_n2336_;
  assign new_n2338_ = new_n1970_ & new_n1998_;
  assign new_n2339_ = ~new_n1968_ & new_n2008_;
  assign new_n2340_ = ~new_n2338_ & new_n2339_;
  assign new_n2341_ = ~new_n1983_ & new_n2340_;
  assign new_n2342_ = new_n1983_ & ~new_n2340_;
  assign new_n2343_ = ~new_n2341_ & ~new_n2342_;
  assign new_n2344_ = ~new_n1992_ & new_n2343_;
  assign new_n2345_ = new_n1992_ & ~new_n2343_;
  assign new_n2346_ = ~new_n2344_ & ~new_n2345_;
  assign new_n2347_ = ~new_n2337_ & new_n2346_;
  assign new_n2348_ = new_n2337_ & ~new_n2346_;
  assign new_n2349_ = ~new_n2347_ & ~new_n2348_;
  assign new_n2350_ = ~new_n2335_ & new_n2349_;
  assign new_n2351_ = new_n2335_ & ~new_n2349_;
  assign new_n2352_ = ~\2_n1366  & ~new_n2351_;
  assign new_n2353_ = ~new_n2350_ & new_n2352_;
  assign new_n2354_ = ~new_n1993_ & new_n2330_;
  assign new_n2355_ = ~new_n1983_ & new_n2354_;
  assign new_n2356_ = new_n1983_ & ~new_n2354_;
  assign new_n2357_ = ~new_n2355_ & ~new_n2356_;
  assign new_n2358_ = ~new_n2337_ & new_n2357_;
  assign new_n2359_ = new_n2337_ & ~new_n2357_;
  assign new_n2360_ = ~new_n2358_ & ~new_n2359_;
  assign new_n2361_ = ~new_n1994_ & new_n2332_;
  assign new_n2362_ = new_n1970_ & new_n1994_;
  assign new_n2363_ = new_n2340_ & ~new_n2362_;
  assign new_n2364_ = new_n2361_ & ~new_n2363_;
  assign new_n2365_ = ~new_n2361_ & new_n2363_;
  assign new_n2366_ = ~new_n2364_ & ~new_n2365_;
  assign new_n2367_ = new_n1986_ & new_n1992_;
  assign new_n2368_ = ~new_n1997_ & ~new_n2367_;
  assign new_n2369_ = ~new_n2366_ & new_n2368_;
  assign new_n2370_ = new_n2366_ & ~new_n2368_;
  assign new_n2371_ = ~new_n2369_ & ~new_n2370_;
  assign new_n2372_ = ~new_n2360_ & new_n2371_;
  assign new_n2373_ = new_n2360_ & ~new_n2371_;
  assign new_n2374_ = ~new_n2372_ & ~new_n2373_;
  assign new_n2375_ = \2_n1366  & new_n2374_;
  assign new_n2376_ = ~new_n2353_ & ~new_n2375_;
  assign new_n2377_ = new_n2329_ & ~new_n2376_;
  assign new_n2378_ = ~new_n2329_ & new_n2376_;
  assign new_n2379_ = ~new_n2377_ & ~new_n2378_;
  assign new_n2380_ = \2_n579  & ~new_n2379_;
  assign new_n2381_ = ~\2_n261  & ~new_n2380_;
  assign new_n2382_ = ~new_n2286_ & new_n2381_;
  assign new_n2383_ = ~new_n2207_ & ~new_n2382_;
  assign new_n2384_ = ~\2_n1205  & ~new_n2383_;
  assign new_n2385_ = ~\2_n228  & new_n2384_;
  assign new_n2386_ = \2_n261  & \2_n520 ;
  assign new_n2387_ = \2_n1660  & ~\2_n591 ;
  assign new_n2388_ = ~\2_n1227  & ~\2_n1660 ;
  assign new_n2389_ = \2_n1575  & ~new_n2388_;
  assign new_n2390_ = ~new_n2387_ & new_n2389_;
  assign new_n2391_ = \2_n1660  & ~\2_n807 ;
  assign new_n2392_ = ~\2_n1660  & ~\2_n714 ;
  assign new_n2393_ = ~new_n2391_ & ~new_n2392_;
  assign new_n2394_ = ~\2_n1575  & ~new_n2393_;
  assign new_n2395_ = ~new_n2390_ & ~new_n2394_;
  assign new_n2396_ = new_n2040_ & new_n2395_;
  assign new_n2397_ = ~new_n2040_ & ~new_n2395_;
  assign new_n2398_ = ~new_n2396_ & ~new_n2397_;
  assign new_n2399_ = \2_n1553  & ~\2_n591 ;
  assign new_n2400_ = ~\2_n1227  & ~\2_n1553 ;
  assign new_n2401_ = \2_n1755  & ~new_n2400_;
  assign new_n2402_ = ~new_n2399_ & new_n2401_;
  assign new_n2403_ = \2_n1553  & ~\2_n807 ;
  assign new_n2404_ = ~\2_n1553  & ~\2_n714 ;
  assign new_n2405_ = ~new_n2403_ & ~new_n2404_;
  assign new_n2406_ = ~\2_n1755  & ~new_n2405_;
  assign new_n2407_ = ~new_n2402_ & ~new_n2406_;
  assign new_n2408_ = \2_n1172  & ~\2_n591 ;
  assign new_n2409_ = ~\2_n1172  & ~\2_n1227 ;
  assign new_n2410_ = \2_n697  & ~new_n2409_;
  assign new_n2411_ = ~new_n2408_ & new_n2410_;
  assign new_n2412_ = \2_n1172  & ~\2_n807 ;
  assign new_n2413_ = ~\2_n1172  & ~\2_n714 ;
  assign new_n2414_ = ~new_n2412_ & ~new_n2413_;
  assign new_n2415_ = ~\2_n697  & ~new_n2414_;
  assign new_n2416_ = ~new_n2411_ & ~new_n2415_;
  assign new_n2417_ = ~new_n2407_ & new_n2416_;
  assign new_n2418_ = new_n2407_ & ~new_n2416_;
  assign new_n2419_ = ~new_n2417_ & ~new_n2418_;
  assign new_n2420_ = ~new_n2398_ & new_n2419_;
  assign new_n2421_ = new_n2398_ & ~new_n2419_;
  assign new_n2422_ = ~new_n2420_ & ~new_n2421_;
  assign new_n2423_ = \2_n1498  & ~\2_n591 ;
  assign new_n2424_ = ~\2_n1227  & ~\2_n1498 ;
  assign new_n2425_ = \2_n1039  & ~new_n2424_;
  assign new_n2426_ = ~new_n2423_ & new_n2425_;
  assign new_n2427_ = \2_n1498  & ~\2_n807 ;
  assign new_n2428_ = ~\2_n1498  & ~\2_n714 ;
  assign new_n2429_ = ~new_n2427_ & ~new_n2428_;
  assign new_n2430_ = ~\2_n1039  & ~new_n2429_;
  assign new_n2431_ = ~new_n2426_ & ~new_n2430_;
  assign new_n2432_ = \2_n1238  & ~\2_n591 ;
  assign new_n2433_ = ~\2_n1227  & ~\2_n1238 ;
  assign new_n2434_ = \2_n1100  & ~new_n2433_;
  assign new_n2435_ = ~new_n2432_ & new_n2434_;
  assign new_n2436_ = \2_n1238  & ~\2_n807 ;
  assign new_n2437_ = ~\2_n1238  & ~\2_n714 ;
  assign new_n2438_ = ~new_n2436_ & ~new_n2437_;
  assign new_n2439_ = ~\2_n1100  & ~new_n2438_;
  assign new_n2440_ = ~new_n2435_ & ~new_n2439_;
  assign new_n2441_ = ~new_n2431_ & new_n2440_;
  assign new_n2442_ = new_n2431_ & ~new_n2440_;
  assign new_n2443_ = ~new_n2441_ & ~new_n2442_;
  assign new_n2444_ = \2_n591  & \2_n617 ;
  assign new_n2445_ = \2_n1227  & ~\2_n617 ;
  assign new_n2446_ = ~new_n2444_ & ~new_n2445_;
  assign new_n2447_ = \2_n39  & ~new_n2446_;
  assign new_n2448_ = \2_n617  & \2_n807 ;
  assign new_n2449_ = ~\2_n617  & \2_n714 ;
  assign new_n2450_ = ~\2_n39  & ~new_n2449_;
  assign new_n2451_ = ~new_n2448_ & new_n2450_;
  assign new_n2452_ = ~new_n2447_ & ~new_n2451_;
  assign new_n2453_ = ~new_n2443_ & ~new_n2452_;
  assign new_n2454_ = new_n2443_ & new_n2452_;
  assign new_n2455_ = ~new_n2453_ & ~new_n2454_;
  assign new_n2456_ = \2_n1729  & \2_n591 ;
  assign new_n2457_ = \2_n1227  & ~\2_n1729 ;
  assign new_n2458_ = ~new_n2456_ & ~new_n2457_;
  assign new_n2459_ = \2_n1135  & ~new_n2458_;
  assign new_n2460_ = \2_n1729  & \2_n807 ;
  assign new_n2461_ = ~\2_n1729  & \2_n714 ;
  assign new_n2462_ = ~\2_n1135  & ~new_n2461_;
  assign new_n2463_ = ~new_n2460_ & new_n2462_;
  assign new_n2464_ = ~new_n2459_ & ~new_n2463_;
  assign new_n2465_ = \2_n319  & \2_n591 ;
  assign new_n2466_ = \2_n1227  & ~\2_n319 ;
  assign new_n2467_ = ~new_n2465_ & ~new_n2466_;
  assign new_n2468_ = \2_n1402  & ~new_n2467_;
  assign new_n2469_ = \2_n319  & \2_n807 ;
  assign new_n2470_ = ~\2_n319  & \2_n714 ;
  assign new_n2471_ = ~\2_n1402  & ~new_n2470_;
  assign new_n2472_ = ~new_n2469_ & new_n2471_;
  assign new_n2473_ = ~new_n2468_ & ~new_n2472_;
  assign new_n2474_ = new_n2464_ & ~new_n2473_;
  assign new_n2475_ = ~new_n2464_ & new_n2473_;
  assign new_n2476_ = ~new_n2474_ & ~new_n2475_;
  assign new_n2477_ = ~new_n2455_ & new_n2476_;
  assign new_n2478_ = new_n2455_ & ~new_n2476_;
  assign new_n2479_ = ~new_n2477_ & ~new_n2478_;
  assign new_n2480_ = new_n2422_ & ~new_n2479_;
  assign new_n2481_ = ~new_n2422_ & new_n2479_;
  assign new_n2482_ = ~\2_n579  & ~new_n2481_;
  assign new_n2483_ = ~new_n2480_ & new_n2482_;
  assign new_n2484_ = new_n2079_ & new_n2112_;
  assign new_n2485_ = ~new_n2077_ & new_n2121_;
  assign new_n2486_ = ~new_n2484_ & new_n2485_;
  assign new_n2487_ = ~new_n2104_ & new_n2486_;
  assign new_n2488_ = new_n2104_ & ~new_n2486_;
  assign new_n2489_ = ~new_n2487_ & ~new_n2488_;
  assign new_n2490_ = ~new_n2091_ & ~new_n2098_;
  assign new_n2491_ = new_n2091_ & new_n2098_;
  assign new_n2492_ = ~new_n2490_ & ~new_n2491_;
  assign new_n2493_ = ~new_n2489_ & new_n2492_;
  assign new_n2494_ = new_n2489_ & ~new_n2492_;
  assign new_n2495_ = ~new_n2493_ & ~new_n2494_;
  assign new_n2496_ = ~new_n2089_ & ~new_n2119_;
  assign new_n2497_ = ~new_n2112_ & new_n2496_;
  assign new_n2498_ = ~new_n2110_ & new_n2497_;
  assign new_n2499_ = new_n2110_ & ~new_n2497_;
  assign new_n2500_ = ~new_n2498_ & ~new_n2499_;
  assign new_n2501_ = ~new_n2111_ & ~new_n2118_;
  assign new_n2502_ = ~new_n2079_ & ~new_n2085_;
  assign new_n2503_ = new_n2079_ & new_n2085_;
  assign new_n2504_ = ~new_n2502_ & ~new_n2503_;
  assign new_n2505_ = new_n2501_ & new_n2504_;
  assign new_n2506_ = ~new_n2501_ & ~new_n2504_;
  assign new_n2507_ = ~new_n2505_ & ~new_n2506_;
  assign new_n2508_ = ~new_n2500_ & new_n2507_;
  assign new_n2509_ = new_n2500_ & ~new_n2507_;
  assign new_n2510_ = ~new_n2508_ & ~new_n2509_;
  assign new_n2511_ = ~new_n2495_ & new_n2510_;
  assign new_n2512_ = new_n2495_ & ~new_n2510_;
  assign new_n2513_ = ~new_n2511_ & ~new_n2512_;
  assign new_n2514_ = ~\2_n1175  & ~new_n2513_;
  assign new_n2515_ = ~new_n2079_ & ~new_n2098_;
  assign new_n2516_ = new_n2079_ & new_n2098_;
  assign new_n2517_ = ~new_n2515_ & ~new_n2516_;
  assign new_n2518_ = new_n2091_ & new_n2105_;
  assign new_n2519_ = new_n2079_ & new_n2518_;
  assign new_n2520_ = new_n2486_ & ~new_n2519_;
  assign new_n2521_ = ~new_n2104_ & ~new_n2520_;
  assign new_n2522_ = new_n2104_ & new_n2520_;
  assign new_n2523_ = ~new_n2521_ & ~new_n2522_;
  assign new_n2524_ = ~new_n2517_ & new_n2523_;
  assign new_n2525_ = new_n2517_ & ~new_n2523_;
  assign new_n2526_ = ~new_n2524_ & ~new_n2525_;
  assign new_n2527_ = ~new_n2105_ & new_n2501_;
  assign new_n2528_ = ~new_n2085_ & ~new_n2091_;
  assign new_n2529_ = new_n2085_ & new_n2091_;
  assign new_n2530_ = ~new_n2528_ & ~new_n2529_;
  assign new_n2531_ = ~new_n2527_ & new_n2530_;
  assign new_n2532_ = new_n2527_ & ~new_n2530_;
  assign new_n2533_ = ~new_n2531_ & ~new_n2532_;
  assign new_n2534_ = new_n2497_ & ~new_n2518_;
  assign new_n2535_ = new_n2104_ & ~new_n2110_;
  assign new_n2536_ = ~new_n2534_ & ~new_n2535_;
  assign new_n2537_ = new_n2534_ & new_n2535_;
  assign new_n2538_ = ~new_n2536_ & ~new_n2537_;
  assign new_n2539_ = ~new_n2533_ & new_n2538_;
  assign new_n2540_ = new_n2533_ & ~new_n2538_;
  assign new_n2541_ = ~new_n2539_ & ~new_n2540_;
  assign new_n2542_ = new_n2526_ & ~new_n2541_;
  assign new_n2543_ = ~new_n2526_ & new_n2541_;
  assign new_n2544_ = \2_n1175  & ~new_n2543_;
  assign new_n2545_ = ~new_n2542_ & new_n2544_;
  assign new_n2546_ = ~new_n2514_ & ~new_n2545_;
  assign new_n2547_ = new_n2048_ & ~new_n2055_;
  assign new_n2548_ = ~new_n2048_ & new_n2055_;
  assign new_n2549_ = ~new_n2547_ & ~new_n2548_;
  assign new_n2550_ = ~new_n2068_ & ~new_n2549_;
  assign new_n2551_ = new_n2068_ & new_n2549_;
  assign new_n2552_ = ~new_n2550_ & ~new_n2551_;
  assign new_n2553_ = new_n2066_ & ~new_n2129_;
  assign new_n2554_ = ~new_n2066_ & new_n2129_;
  assign new_n2555_ = ~new_n2553_ & ~new_n2554_;
  assign new_n2556_ = ~new_n2063_ & new_n2070_;
  assign new_n2557_ = new_n2063_ & ~new_n2070_;
  assign new_n2558_ = ~new_n2556_ & ~new_n2557_;
  assign new_n2559_ = ~new_n2555_ & new_n2558_;
  assign new_n2560_ = new_n2555_ & ~new_n2558_;
  assign new_n2561_ = ~new_n2559_ & ~new_n2560_;
  assign new_n2562_ = ~new_n2552_ & new_n2561_;
  assign new_n2563_ = new_n2552_ & ~new_n2561_;
  assign new_n2564_ = ~new_n2562_ & ~new_n2563_;
  assign new_n2565_ = new_n2124_ & new_n2564_;
  assign new_n2566_ = ~\2_n1175  & ~new_n2565_;
  assign new_n2567_ = new_n2068_ & ~new_n2130_;
  assign new_n2568_ = new_n2549_ & ~new_n2567_;
  assign new_n2569_ = ~new_n2549_ & new_n2567_;
  assign new_n2570_ = ~new_n2568_ & ~new_n2569_;
  assign new_n2571_ = ~new_n2063_ & new_n2129_;
  assign new_n2572_ = new_n2132_ & ~new_n2571_;
  assign new_n2573_ = ~new_n2132_ & new_n2571_;
  assign new_n2574_ = ~new_n2572_ & ~new_n2573_;
  assign new_n2575_ = ~new_n2555_ & new_n2574_;
  assign new_n2576_ = new_n2555_ & ~new_n2574_;
  assign new_n2577_ = ~new_n2575_ & ~new_n2576_;
  assign new_n2578_ = ~new_n2570_ & new_n2577_;
  assign new_n2579_ = new_n2570_ & ~new_n2577_;
  assign new_n2580_ = ~new_n2578_ & ~new_n2579_;
  assign new_n2581_ = ~new_n2124_ & ~new_n2580_;
  assign new_n2582_ = new_n2566_ & ~new_n2581_;
  assign new_n2583_ = new_n2109_ & new_n2518_;
  assign new_n2584_ = new_n2124_ & ~new_n2583_;
  assign new_n2585_ = ~new_n2564_ & new_n2584_;
  assign new_n2586_ = new_n2580_ & ~new_n2584_;
  assign new_n2587_ = ~new_n2585_ & ~new_n2586_;
  assign new_n2588_ = \2_n1175  & ~new_n2587_;
  assign new_n2589_ = ~new_n2582_ & ~new_n2588_;
  assign new_n2590_ = ~new_n2546_ & ~new_n2589_;
  assign new_n2591_ = new_n2546_ & new_n2589_;
  assign new_n2592_ = ~new_n2590_ & ~new_n2591_;
  assign new_n2593_ = \2_n579  & new_n2592_;
  assign new_n2594_ = ~\2_n261  & ~new_n2593_;
  assign new_n2595_ = ~new_n2483_ & new_n2594_;
  assign new_n2596_ = ~new_n2386_ & ~new_n2595_;
  assign new_n2597_ = ~\2_n1205  & ~new_n2596_;
  assign new_n2598_ = \2_n228  & new_n2597_;
  assign new_n2599_ = ~new_n2385_ & ~new_n2598_;
  assign new_n2600_ = new_n2206_ & new_n2599_;
  assign \2_n1065  = \2_n1050 ;
  assign new_n2602_ = \2_n1238  & \2_n1288 ;
  assign new_n2603_ = ~\2_n1238  & \2_n721 ;
  assign new_n2604_ = \2_n1100  & ~new_n2603_;
  assign new_n2605_ = ~new_n2602_ & new_n2604_;
  assign new_n2606_ = \2_n1238  & \2_n77 ;
  assign new_n2607_ = ~\2_n1238  & \2_n1519 ;
  assign new_n2608_ = ~new_n2606_ & ~new_n2607_;
  assign new_n2609_ = ~\2_n1100  & ~new_n2608_;
  assign new_n2610_ = ~new_n2605_ & ~new_n2609_;
  assign new_n2611_ = \2_n1172  & ~\2_n1288 ;
  assign new_n2612_ = ~\2_n1172  & ~\2_n721 ;
  assign new_n2613_ = ~new_n2611_ & ~new_n2612_;
  assign new_n2614_ = \2_n697  & ~new_n2613_;
  assign new_n2615_ = \2_n1172  & ~\2_n77 ;
  assign new_n2616_ = ~\2_n1172  & ~\2_n1519 ;
  assign new_n2617_ = ~\2_n697  & ~new_n2616_;
  assign new_n2618_ = ~new_n2615_ & new_n2617_;
  assign new_n2619_ = ~new_n2614_ & ~new_n2618_;
  assign new_n2620_ = ~new_n2610_ & ~new_n2619_;
  assign new_n2621_ = \2_n1288  & \2_n1729 ;
  assign new_n2622_ = ~\2_n1729  & \2_n721 ;
  assign new_n2623_ = \2_n1135  & ~new_n2622_;
  assign new_n2624_ = ~new_n2621_ & new_n2623_;
  assign new_n2625_ = \2_n1729  & \2_n77 ;
  assign new_n2626_ = \2_n1519  & ~\2_n1729 ;
  assign new_n2627_ = ~new_n2625_ & ~new_n2626_;
  assign new_n2628_ = ~\2_n1135  & ~new_n2627_;
  assign new_n2629_ = ~new_n2624_ & ~new_n2628_;
  assign new_n2630_ = ~\2_n1288  & \2_n1553 ;
  assign new_n2631_ = ~\2_n1553  & ~\2_n721 ;
  assign new_n2632_ = ~new_n2630_ & ~new_n2631_;
  assign new_n2633_ = \2_n1755  & ~new_n2632_;
  assign new_n2634_ = \2_n1553  & ~\2_n77 ;
  assign new_n2635_ = ~\2_n1519  & ~\2_n1553 ;
  assign new_n2636_ = ~\2_n1755  & ~new_n2635_;
  assign new_n2637_ = ~new_n2634_ & new_n2636_;
  assign new_n2638_ = ~new_n2633_ & ~new_n2637_;
  assign new_n2639_ = ~new_n2629_ & ~new_n2638_;
  assign new_n2640_ = new_n2620_ & new_n2639_;
  assign new_n2641_ = \2_n1288  & \2_n1660 ;
  assign new_n2642_ = ~\2_n1660  & \2_n721 ;
  assign new_n2643_ = \2_n1575  & ~new_n2642_;
  assign new_n2644_ = ~new_n2641_ & new_n2643_;
  assign new_n2645_ = \2_n1660  & \2_n77 ;
  assign new_n2646_ = \2_n1519  & ~\2_n1660 ;
  assign new_n2647_ = ~new_n2645_ & ~new_n2646_;
  assign new_n2648_ = ~\2_n1575  & ~new_n2647_;
  assign new_n2649_ = ~new_n2644_ & ~new_n2648_;
  assign new_n2650_ = \2_n1288  & \2_n319 ;
  assign new_n2651_ = ~\2_n319  & \2_n721 ;
  assign new_n2652_ = \2_n1402  & ~new_n2651_;
  assign new_n2653_ = ~new_n2650_ & new_n2652_;
  assign new_n2654_ = \2_n319  & \2_n77 ;
  assign new_n2655_ = \2_n1519  & ~\2_n319 ;
  assign new_n2656_ = ~new_n2654_ & ~new_n2655_;
  assign new_n2657_ = ~\2_n1402  & ~new_n2656_;
  assign new_n2658_ = ~new_n2653_ & ~new_n2657_;
  assign new_n2659_ = ~new_n2649_ & ~new_n2658_;
  assign new_n2660_ = ~\2_n1288  & \2_n617 ;
  assign new_n2661_ = ~\2_n617  & ~\2_n721 ;
  assign new_n2662_ = ~new_n2660_ & ~new_n2661_;
  assign new_n2663_ = \2_n39  & ~new_n2662_;
  assign new_n2664_ = \2_n617  & ~\2_n77 ;
  assign new_n2665_ = ~\2_n1519  & ~\2_n617 ;
  assign new_n2666_ = ~\2_n39  & ~new_n2665_;
  assign new_n2667_ = ~new_n2664_ & new_n2666_;
  assign new_n2668_ = ~new_n2663_ & ~new_n2667_;
  assign new_n2669_ = ~new_n2185_ & ~new_n2668_;
  assign new_n2670_ = new_n2659_ & new_n2669_;
  assign new_n2671_ = new_n2640_ & new_n2670_;
  assign \2_n107  = ~new_n2040_ & new_n2671_;
  assign new_n2673_ = \2_n386  & ~\2_n579 ;
  assign new_n2674_ = \2_n261  & new_n2673_;
  assign new_n2675_ = ~\2_n579  & new_n2649_;
  assign new_n2676_ = ~\2_n261  & new_n2675_;
  assign new_n2677_ = new_n2055_ & new_n2068_;
  assign new_n2678_ = new_n2125_ & ~new_n2677_;
  assign new_n2679_ = ~new_n2069_ & new_n2678_;
  assign new_n2680_ = ~new_n2055_ & new_n2567_;
  assign new_n2681_ = new_n2055_ & ~new_n2567_;
  assign new_n2682_ = ~new_n2680_ & ~new_n2681_;
  assign new_n2683_ = ~new_n2125_ & ~new_n2682_;
  assign new_n2684_ = ~new_n2679_ & ~new_n2683_;
  assign new_n2685_ = \2_n579  & ~new_n2684_;
  assign new_n2686_ = ~\2_n261  & new_n2685_;
  assign new_n2687_ = ~new_n2676_ & ~new_n2686_;
  assign \2_n1087  = ~new_n2674_ & new_n2687_;
  assign new_n2689_ = \2_n307  & \2_n565 ;
  assign new_n2690_ = \2_n377  & new_n2689_;
  assign new_n2691_ = \2_n1540  & \2_n307 ;
  assign new_n2692_ = ~\2_n377  & new_n2691_;
  assign new_n2693_ = ~new_n2690_ & ~new_n2692_;
  assign new_n2694_ = \2_n1361  & ~\2_n579 ;
  assign new_n2695_ = \2_n261  & new_n2694_;
  assign new_n2696_ = \2_n1288  & \2_n238 ;
  assign new_n2697_ = ~\2_n238  & ~\2_n77 ;
  assign new_n2698_ = ~new_n2696_ & ~new_n2697_;
  assign new_n2699_ = ~\2_n579  & ~new_n2698_;
  assign new_n2700_ = ~\2_n261  & new_n2699_;
  assign new_n2701_ = \2_n1788  & new_n1993_;
  assign new_n2702_ = ~new_n1983_ & new_n2701_;
  assign new_n2703_ = new_n2332_ & ~new_n2702_;
  assign new_n2704_ = ~new_n1970_ & new_n2703_;
  assign new_n2705_ = new_n1970_ & ~new_n2703_;
  assign new_n2706_ = ~new_n2704_ & ~new_n2705_;
  assign new_n2707_ = \2_n579  & new_n2706_;
  assign new_n2708_ = ~\2_n261  & new_n2707_;
  assign new_n2709_ = ~new_n2700_ & ~new_n2708_;
  assign \2_n487  = ~new_n2695_ & new_n2709_;
  assign new_n2711_ = ~\2_n307  & ~\2_n487 ;
  assign new_n2712_ = ~\2_n377  & new_n2711_;
  assign new_n2713_ = ~\2_n579  & \2_n999 ;
  assign new_n2714_ = \2_n261  & new_n2713_;
  assign new_n2715_ = ~\2_n579  & new_n2658_;
  assign new_n2716_ = ~\2_n261  & new_n2715_;
  assign new_n2717_ = ~new_n2098_ & new_n2188_;
  assign new_n2718_ = new_n2091_ & new_n2717_;
  assign new_n2719_ = new_n2497_ & ~new_n2718_;
  assign new_n2720_ = new_n2079_ & ~new_n2719_;
  assign new_n2721_ = ~new_n2079_ & new_n2719_;
  assign new_n2722_ = ~new_n2720_ & ~new_n2721_;
  assign new_n2723_ = \2_n579  & new_n2722_;
  assign new_n2724_ = ~\2_n261  & new_n2723_;
  assign new_n2725_ = ~new_n2716_ & ~new_n2724_;
  assign \2_n1710  = ~new_n2714_ & new_n2725_;
  assign new_n2727_ = ~\2_n307  & ~\2_n1710 ;
  assign new_n2728_ = \2_n377  & new_n2727_;
  assign new_n2729_ = ~new_n2712_ & ~new_n2728_;
  assign \2_n1096  = ~new_n2693_ | ~new_n2729_;
  assign new_n2731_ = ~\2_n579  & \2_n9 ;
  assign new_n2732_ = \2_n261  & new_n2731_;
  assign new_n2733_ = ~\2_n579  & new_n2610_;
  assign new_n2734_ = ~\2_n261  & new_n2733_;
  assign new_n2735_ = new_n2501_ & ~new_n2717_;
  assign new_n2736_ = new_n2091_ & new_n2735_;
  assign new_n2737_ = ~new_n2091_ & ~new_n2735_;
  assign new_n2738_ = ~new_n2736_ & ~new_n2737_;
  assign new_n2739_ = \2_n579  & ~new_n2738_;
  assign new_n2740_ = ~\2_n261  & new_n2739_;
  assign new_n2741_ = ~new_n2734_ & ~new_n2740_;
  assign \2_n1110  = ~new_n2732_ & new_n2741_;
  assign \2_n117  = ~\2_n601  | ~\2_n841 ;
  assign \2_n1163  = ~\2_n1463  | \2_n117 ;
  assign new_n2745_ = \2_n335  & \2_n627 ;
  assign new_n2746_ = \2_n378  & new_n2745_;
  assign new_n2747_ = \2_n270  & \2_n627 ;
  assign new_n2748_ = ~\2_n378  & new_n2747_;
  assign new_n2749_ = ~new_n2746_ & ~new_n2748_;
  assign new_n2750_ = \2_n1182  & ~\2_n579 ;
  assign new_n2751_ = \2_n261  & new_n2750_;
  assign new_n2752_ = ~\2_n579  & new_n2225_;
  assign new_n2753_ = ~\2_n261  & new_n2752_;
  assign new_n2754_ = ~new_n1955_ & new_n1958_;
  assign new_n2755_ = ~new_n1959_ & new_n2012_;
  assign new_n2756_ = ~new_n2754_ & new_n2755_;
  assign new_n2757_ = ~new_n1958_ & ~new_n2312_;
  assign new_n2758_ = new_n1958_ & new_n2312_;
  assign new_n2759_ = ~new_n2757_ & ~new_n2758_;
  assign new_n2760_ = ~new_n2012_ & new_n2759_;
  assign new_n2761_ = ~new_n2756_ & ~new_n2760_;
  assign new_n2762_ = \2_n579  & ~new_n2761_;
  assign new_n2763_ = ~\2_n261  & new_n2762_;
  assign new_n2764_ = ~new_n2753_ & ~new_n2763_;
  assign \2_n882  = ~new_n2751_ & new_n2764_;
  assign new_n2766_ = ~\2_n627  & ~\2_n882 ;
  assign new_n2767_ = ~\2_n378  & new_n2766_;
  assign new_n2768_ = ~\2_n579  & \2_n779 ;
  assign new_n2769_ = \2_n261  & new_n2768_;
  assign new_n2770_ = ~\2_n579  & new_n2619_;
  assign new_n2771_ = ~\2_n261  & new_n2770_;
  assign new_n2772_ = ~new_n2063_ & new_n2066_;
  assign new_n2773_ = ~new_n2067_ & new_n2125_;
  assign new_n2774_ = ~new_n2772_ & new_n2773_;
  assign new_n2775_ = ~new_n2066_ & ~new_n2571_;
  assign new_n2776_ = new_n2066_ & new_n2571_;
  assign new_n2777_ = ~new_n2775_ & ~new_n2776_;
  assign new_n2778_ = ~new_n2125_ & new_n2777_;
  assign new_n2779_ = ~new_n2774_ & ~new_n2778_;
  assign new_n2780_ = \2_n579  & ~new_n2779_;
  assign new_n2781_ = ~\2_n261  & new_n2780_;
  assign new_n2782_ = ~new_n2771_ & ~new_n2781_;
  assign \2_n456  = ~new_n2769_ & new_n2782_;
  assign new_n2784_ = ~\2_n627  & ~\2_n456 ;
  assign new_n2785_ = \2_n378  & new_n2784_;
  assign new_n2786_ = ~new_n2767_ & ~new_n2785_;
  assign new_n2787_ = new_n2749_ & new_n2786_;
  assign \2_n1186  = \2_n1050 ;
  assign new_n2789_ = ~\2_n1279  & new_n2104_;
  assign new_n2790_ = ~new_n2188_ & ~new_n2789_;
  assign new_n2791_ = ~new_n2192_ & ~new_n2790_;
  assign new_n2792_ = ~new_n2722_ & new_n2738_;
  assign new_n2793_ = new_n2791_ & new_n2792_;
  assign new_n2794_ = new_n2079_ & new_n2718_;
  assign new_n2795_ = new_n2486_ & ~new_n2794_;
  assign new_n2796_ = ~new_n2085_ & ~new_n2795_;
  assign new_n2797_ = new_n2085_ & new_n2795_;
  assign new_n2798_ = ~new_n2796_ & ~new_n2797_;
  assign new_n2799_ = new_n2125_ & new_n2129_;
  assign new_n2800_ = ~new_n2125_ & ~new_n2129_;
  assign new_n2801_ = ~new_n2799_ & ~new_n2800_;
  assign new_n2802_ = ~new_n2798_ & ~new_n2801_;
  assign new_n2803_ = new_n2137_ & new_n2684_;
  assign new_n2804_ = new_n2802_ & new_n2803_;
  assign new_n2805_ = new_n2793_ & new_n2804_;
  assign \2_n1224  = new_n2779_ & new_n2805_;
  assign new_n2807_ = \2_n1357  & \2_n1649 ;
  assign new_n2808_ = ~\2_n342  & ~new_n1941_;
  assign new_n2809_ = ~\2_n495  & new_n2808_;
  assign new_n2810_ = \2_n1790  & new_n1963_;
  assign new_n2811_ = ~\2_n1790  & ~new_n1963_;
  assign new_n2812_ = ~new_n2810_ & ~new_n2811_;
  assign new_n2813_ = ~\2_n342  & new_n2812_;
  assign new_n2814_ = \2_n495  & new_n2813_;
  assign new_n2815_ = ~new_n2809_ & ~new_n2814_;
  assign new_n2816_ = \2_n342  & \2_n482 ;
  assign new_n2817_ = ~\2_n495  & new_n2816_;
  assign new_n2818_ = \2_n342  & ~\2_n1793 ;
  assign new_n2819_ = \2_n495  & new_n2818_;
  assign new_n2820_ = ~new_n2817_ & ~new_n2819_;
  assign new_n2821_ = new_n2815_ & new_n2820_;
  assign \2_n1269  = ~new_n2807_ & ~new_n2821_;
  assign new_n2823_ = \2_n1205  & \2_n606 ;
  assign new_n2824_ = \2_n228  & new_n2823_;
  assign new_n2825_ = \2_n1205  & \2_n387 ;
  assign new_n2826_ = ~\2_n228  & new_n2825_;
  assign new_n2827_ = ~new_n2824_ & ~new_n2826_;
  assign new_n2828_ = \2_n1740  & ~\2_n579 ;
  assign new_n2829_ = \2_n261  & new_n2828_;
  assign new_n2830_ = \2_n1288  & \2_n1435 ;
  assign new_n2831_ = ~\2_n1435  & \2_n721 ;
  assign new_n2832_ = \2_n1016  & ~new_n2831_;
  assign new_n2833_ = ~new_n2830_ & new_n2832_;
  assign new_n2834_ = \2_n1435  & \2_n77 ;
  assign new_n2835_ = ~\2_n1435  & \2_n1519 ;
  assign new_n2836_ = ~new_n2834_ & ~new_n2835_;
  assign new_n2837_ = ~\2_n1016  & ~new_n2836_;
  assign new_n2838_ = ~new_n2833_ & ~new_n2837_;
  assign new_n2839_ = ~\2_n579  & new_n2838_;
  assign new_n2840_ = ~\2_n261  & new_n2839_;
  assign new_n2841_ = new_n2330_ & ~new_n2701_;
  assign new_n2842_ = ~new_n1983_ & ~new_n2841_;
  assign new_n2843_ = new_n1983_ & new_n2841_;
  assign new_n2844_ = ~new_n2842_ & ~new_n2843_;
  assign new_n2845_ = \2_n579  & new_n2844_;
  assign new_n2846_ = ~\2_n261  & new_n2845_;
  assign new_n2847_ = ~new_n2840_ & ~new_n2846_;
  assign \2_n1314  = ~new_n2829_ & new_n2847_;
  assign new_n2849_ = ~\2_n1205  & ~\2_n1314 ;
  assign new_n2850_ = ~\2_n228  & new_n2849_;
  assign new_n2851_ = ~\2_n1205  & ~\2_n1110 ;
  assign new_n2852_ = \2_n228  & new_n2851_;
  assign new_n2853_ = ~new_n2850_ & ~new_n2852_;
  assign new_n2854_ = new_n2827_ & new_n2853_;
  assign \2_n1270  = \2_n1050 ;
  assign new_n2856_ = \2_n186  & \2_n676 ;
  assign new_n2857_ = \2_n560  & new_n2856_;
  assign new_n2858_ = \2_n1207  & \2_n186 ;
  assign new_n2859_ = ~\2_n560  & new_n2858_;
  assign new_n2860_ = ~new_n2857_ & ~new_n2859_;
  assign new_n2861_ = \2_n1753  & ~\2_n579 ;
  assign new_n2862_ = \2_n261  & new_n2861_;
  assign new_n2863_ = ~\2_n579  & new_n2255_;
  assign new_n2864_ = ~\2_n261  & new_n2863_;
  assign new_n2865_ = \2_n1788  & ~new_n1986_;
  assign new_n2866_ = ~new_n2165_ & ~new_n2865_;
  assign new_n2867_ = \2_n579  & ~new_n2866_;
  assign new_n2868_ = ~\2_n261  & new_n2867_;
  assign new_n2869_ = ~new_n2864_ & ~new_n2868_;
  assign \2_n454  = ~new_n2862_ & new_n2869_;
  assign new_n2871_ = ~\2_n186  & ~\2_n454 ;
  assign new_n2872_ = ~\2_n560  & new_n2871_;
  assign new_n2873_ = \2_n190  & ~\2_n579 ;
  assign new_n2874_ = \2_n261  & new_n2873_;
  assign new_n2875_ = ~\2_n579  & new_n2668_;
  assign new_n2876_ = ~\2_n261  & new_n2875_;
  assign new_n2877_ = \2_n579  & new_n2790_;
  assign new_n2878_ = ~\2_n261  & new_n2877_;
  assign new_n2879_ = ~new_n2876_ & ~new_n2878_;
  assign \2_n259  = ~new_n2874_ & new_n2879_;
  assign new_n2881_ = ~\2_n186  & ~\2_n259 ;
  assign new_n2882_ = \2_n560  & new_n2881_;
  assign new_n2883_ = ~new_n2872_ & ~new_n2882_;
  assign \2_n1297  = ~new_n2860_ | ~new_n2883_;
  assign new_n2885_ = new_n1946_ & ~new_n2011_;
  assign new_n2886_ = new_n2017_ & new_n2885_;
  assign \2_n130  = ~new_n1964_ | new_n2886_;
  assign new_n2888_ = \2_n627  & \2_n962 ;
  assign new_n2889_ = \2_n378  & new_n2888_;
  assign new_n2890_ = \2_n1663  & \2_n627 ;
  assign new_n2891_ = ~\2_n378  & new_n2890_;
  assign new_n2892_ = ~new_n2889_ & ~new_n2891_;
  assign new_n2893_ = ~\2_n627  & ~new_n2383_;
  assign new_n2894_ = ~\2_n378  & new_n2893_;
  assign new_n2895_ = ~\2_n627  & ~new_n2596_;
  assign new_n2896_ = \2_n378  & new_n2895_;
  assign new_n2897_ = ~new_n2894_ & ~new_n2896_;
  assign new_n2898_ = new_n2892_ & new_n2897_;
  assign \2_n1322  = \2_n1050 ;
  assign new_n2900_ = \2_n1119  & \2_n307 ;
  assign new_n2901_ = \2_n377  & new_n2900_;
  assign new_n2902_ = \2_n239  & \2_n307 ;
  assign new_n2903_ = ~\2_n377  & new_n2902_;
  assign new_n2904_ = ~new_n2901_ & ~new_n2903_;
  assign new_n2905_ = \2_n1095  & ~\2_n579 ;
  assign new_n2906_ = \2_n261  & new_n2905_;
  assign new_n2907_ = ~\2_n1288  & \2_n380 ;
  assign new_n2908_ = ~\2_n380  & ~\2_n721 ;
  assign new_n2909_ = ~new_n2907_ & ~new_n2908_;
  assign new_n2910_ = \2_n1391  & ~new_n2909_;
  assign new_n2911_ = \2_n380  & ~\2_n77 ;
  assign new_n2912_ = ~\2_n1519  & ~\2_n380 ;
  assign new_n2913_ = ~\2_n1391  & ~new_n2912_;
  assign new_n2914_ = ~new_n2911_ & new_n2913_;
  assign new_n2915_ = ~new_n2910_ & ~new_n2914_;
  assign new_n2916_ = ~\2_n579  & new_n2915_;
  assign new_n2917_ = ~\2_n261  & new_n2916_;
  assign new_n2918_ = new_n1970_ & new_n2702_;
  assign new_n2919_ = new_n2340_ & ~new_n2918_;
  assign new_n2920_ = ~new_n1976_ & ~new_n2919_;
  assign new_n2921_ = new_n1976_ & new_n2919_;
  assign new_n2922_ = ~new_n2920_ & ~new_n2921_;
  assign new_n2923_ = \2_n579  & new_n2922_;
  assign new_n2924_ = ~\2_n261  & new_n2923_;
  assign new_n2925_ = ~new_n2917_ & ~new_n2924_;
  assign \2_n1495  = ~new_n2906_ & new_n2925_;
  assign new_n2927_ = ~\2_n307  & ~\2_n1495 ;
  assign new_n2928_ = ~\2_n377  & new_n2927_;
  assign new_n2929_ = \2_n157  & ~\2_n579 ;
  assign new_n2930_ = \2_n261  & new_n2929_;
  assign new_n2931_ = ~\2_n579  & new_n2629_;
  assign new_n2932_ = ~\2_n261  & new_n2931_;
  assign new_n2933_ = \2_n579  & new_n2798_;
  assign new_n2934_ = ~\2_n261  & new_n2933_;
  assign new_n2935_ = ~new_n2932_ & ~new_n2934_;
  assign \2_n1631  = ~new_n2930_ & new_n2935_;
  assign new_n2937_ = ~\2_n307  & ~\2_n1631 ;
  assign new_n2938_ = \2_n377  & new_n2937_;
  assign new_n2939_ = ~new_n2928_ & ~new_n2938_;
  assign \2_n1377  = ~new_n2904_ | ~new_n2939_;
  assign new_n2941_ = \2_n307  & \2_n676 ;
  assign new_n2942_ = \2_n377  & new_n2941_;
  assign new_n2943_ = \2_n1207  & \2_n307 ;
  assign new_n2944_ = ~\2_n377  & new_n2943_;
  assign new_n2945_ = ~new_n2942_ & ~new_n2944_;
  assign new_n2946_ = ~\2_n307  & ~\2_n454 ;
  assign new_n2947_ = ~\2_n377  & new_n2946_;
  assign new_n2948_ = ~\2_n307  & ~\2_n259 ;
  assign new_n2949_ = \2_n377  & new_n2948_;
  assign new_n2950_ = ~new_n2947_ & ~new_n2949_;
  assign \2_n1390  = ~new_n2945_ | ~new_n2950_;
  assign \2_n1409  = \2_n1427  | ~\2_n841 ;
  assign new_n2953_ = \2_n60  & ~new_n2045_;
  assign new_n2954_ = ~new_n2048_ & new_n2052_;
  assign new_n2955_ = ~new_n2953_ & ~new_n2954_;
  assign new_n2956_ = ~new_n2048_ & new_n2069_;
  assign new_n2957_ = ~new_n2048_ & new_n2131_;
  assign new_n2958_ = ~new_n2124_ & new_n2957_;
  assign new_n2959_ = ~new_n2956_ & ~new_n2958_;
  assign \2_n1414  = ~new_n2955_ | ~new_n2959_;
  assign new_n2961_ = \2_n1205  & \2_n830 ;
  assign new_n2962_ = \2_n228  & new_n2961_;
  assign new_n2963_ = \2_n1033  & \2_n1205 ;
  assign new_n2964_ = ~\2_n228  & new_n2963_;
  assign new_n2965_ = ~new_n2962_ & ~new_n2964_;
  assign new_n2966_ = ~\2_n1205  & ~\2_n1027 ;
  assign new_n2967_ = ~\2_n228  & new_n2966_;
  assign new_n2968_ = ~\2_n1205  & ~\2_n123 ;
  assign new_n2969_ = \2_n228  & new_n2968_;
  assign new_n2970_ = ~new_n2967_ & ~new_n2969_;
  assign new_n2971_ = new_n2965_ & new_n2970_;
  assign \2_n1462  = \2_n1050 ;
  assign \2_n1491  = ~\2_n119  | ~\2_n1768 ;
  assign new_n2974_ = \2_n1119  & \2_n186 ;
  assign new_n2975_ = \2_n560  & new_n2974_;
  assign new_n2976_ = \2_n186  & \2_n239 ;
  assign new_n2977_ = ~\2_n560  & new_n2976_;
  assign new_n2978_ = ~new_n2975_ & ~new_n2977_;
  assign new_n2979_ = ~\2_n186  & ~\2_n1495 ;
  assign new_n2980_ = ~\2_n560  & new_n2979_;
  assign new_n2981_ = ~\2_n186  & ~\2_n1631 ;
  assign new_n2982_ = \2_n560  & new_n2981_;
  assign new_n2983_ = ~new_n2980_ & ~new_n2982_;
  assign \2_n1510  = ~new_n2978_ | ~new_n2983_;
  assign new_n2985_ = ~\2_n1515  & \2_n643 ;
  assign new_n2986_ = \2_n1515  & ~\2_n643 ;
  assign new_n2987_ = ~new_n2985_ & ~new_n2986_;
  assign new_n2988_ = \2_n1043  & ~\2_n1435 ;
  assign new_n2989_ = ~\2_n1043  & \2_n1435 ;
  assign new_n2990_ = ~new_n2988_ & ~new_n2989_;
  assign new_n2991_ = ~new_n2987_ & new_n2990_;
  assign new_n2992_ = new_n2987_ & ~new_n2990_;
  assign new_n2993_ = ~new_n2991_ & ~new_n2992_;
  assign new_n2994_ = \2_n380  & ~new_n2993_;
  assign new_n2995_ = ~\2_n380  & new_n2993_;
  assign new_n2996_ = ~new_n2994_ & ~new_n2995_;
  assign new_n2997_ = \2_n946  & ~\2_n966 ;
  assign new_n2998_ = ~\2_n946  & \2_n966 ;
  assign new_n2999_ = ~new_n2997_ & ~new_n2998_;
  assign new_n3000_ = \2_n1518  & ~\2_n288 ;
  assign new_n3001_ = ~\2_n1518  & \2_n288 ;
  assign new_n3002_ = ~new_n3000_ & ~new_n3001_;
  assign new_n3003_ = ~new_n2999_ & new_n3002_;
  assign new_n3004_ = new_n2999_ & ~new_n3002_;
  assign new_n3005_ = ~new_n3003_ & ~new_n3004_;
  assign new_n3006_ = ~new_n2996_ & new_n3005_;
  assign new_n3007_ = new_n2996_ & ~new_n3005_;
  assign \2_n1511  = new_n3006_ | new_n3007_;
  assign new_n3009_ = \2_n19  & \2_n307 ;
  assign new_n3010_ = \2_n377  & new_n3009_;
  assign new_n3011_ = \2_n307  & \2_n955 ;
  assign new_n3012_ = ~\2_n377  & new_n3011_;
  assign new_n3013_ = ~new_n3010_ & ~new_n3012_;
  assign new_n3014_ = \2_n1097  & ~\2_n579 ;
  assign new_n3015_ = \2_n261  & new_n3014_;
  assign new_n3016_ = ~\2_n579  & new_n2216_;
  assign new_n3017_ = ~\2_n261  & new_n3016_;
  assign new_n3018_ = ~new_n2012_ & ~new_n2016_;
  assign new_n3019_ = new_n2012_ & new_n2016_;
  assign new_n3020_ = ~new_n3018_ & ~new_n3019_;
  assign new_n3021_ = \2_n579  & new_n3020_;
  assign new_n3022_ = ~\2_n261  & new_n3021_;
  assign new_n3023_ = ~new_n3017_ & ~new_n3022_;
  assign \2_n964  = ~new_n3015_ & new_n3023_;
  assign new_n3025_ = ~\2_n307  & ~\2_n964 ;
  assign new_n3026_ = ~\2_n377  & new_n3025_;
  assign new_n3027_ = ~\2_n579  & \2_n984 ;
  assign new_n3028_ = \2_n261  & new_n3027_;
  assign new_n3029_ = ~\2_n579  & new_n2638_;
  assign new_n3030_ = ~\2_n261  & new_n3029_;
  assign new_n3031_ = \2_n579  & new_n2801_;
  assign new_n3032_ = ~\2_n261  & new_n3031_;
  assign new_n3033_ = ~new_n3030_ & ~new_n3032_;
  assign \2_n370  = ~new_n3028_ & new_n3033_;
  assign new_n3035_ = ~\2_n307  & ~\2_n370 ;
  assign new_n3036_ = \2_n377  & new_n3035_;
  assign new_n3037_ = ~new_n3026_ & ~new_n3036_;
  assign \2_n1543  = ~new_n3013_ | ~new_n3037_;
  assign new_n3039_ = \2_n627  & \2_n830 ;
  assign new_n3040_ = \2_n378  & new_n3039_;
  assign new_n3041_ = \2_n1033  & \2_n627 ;
  assign new_n3042_ = ~\2_n378  & new_n3041_;
  assign new_n3043_ = ~new_n3040_ & ~new_n3042_;
  assign new_n3044_ = ~\2_n627  & ~\2_n1027 ;
  assign new_n3045_ = ~\2_n378  & new_n3044_;
  assign new_n3046_ = ~\2_n627  & ~\2_n123 ;
  assign new_n3047_ = \2_n378  & new_n3046_;
  assign new_n3048_ = ~new_n3045_ & ~new_n3047_;
  assign new_n3049_ = new_n3043_ & new_n3048_;
  assign \2_n158  = \2_n1050 ;
  assign \2_n1584  = \2_n1613  & \2_n912 ;
  assign new_n3052_ = \2_n1205  & \2_n1353 ;
  assign new_n3053_ = \2_n228  & new_n3052_;
  assign new_n3054_ = \2_n1205  & \2_n530 ;
  assign new_n3055_ = ~\2_n228  & new_n3054_;
  assign new_n3056_ = ~new_n3053_ & ~new_n3055_;
  assign new_n3057_ = ~\2_n579  & \2_n813 ;
  assign new_n3058_ = \2_n261  & new_n3057_;
  assign new_n3059_ = ~\2_n579  & new_n2231_;
  assign new_n3060_ = ~\2_n261  & new_n3059_;
  assign new_n3061_ = new_n1946_ & ~new_n2290_;
  assign new_n3062_ = ~new_n1946_ & new_n2290_;
  assign new_n3063_ = new_n2012_ & ~new_n3062_;
  assign new_n3064_ = ~new_n3061_ & new_n3063_;
  assign new_n3065_ = new_n1946_ & new_n2308_;
  assign new_n3066_ = ~new_n1946_ & ~new_n2308_;
  assign new_n3067_ = ~new_n3065_ & ~new_n3066_;
  assign new_n3068_ = ~new_n2012_ & ~new_n3067_;
  assign new_n3069_ = ~new_n3064_ & ~new_n3068_;
  assign new_n3070_ = \2_n579  & ~new_n3069_;
  assign new_n3071_ = ~\2_n261  & new_n3070_;
  assign new_n3072_ = ~new_n3060_ & ~new_n3071_;
  assign \2_n75  = ~new_n3058_ & new_n3072_;
  assign new_n3074_ = ~\2_n1205  & ~\2_n75 ;
  assign new_n3075_ = ~\2_n228  & new_n3074_;
  assign new_n3076_ = ~\2_n1205  & ~\2_n1087 ;
  assign new_n3077_ = \2_n228  & new_n3076_;
  assign new_n3078_ = ~new_n3075_ & ~new_n3077_;
  assign new_n3079_ = new_n3056_ & new_n3078_;
  assign \2_n1587  = \2_n1050 ;
  assign new_n3081_ = new_n2168_ & ~new_n2844_;
  assign new_n3082_ = ~new_n2706_ & ~new_n2922_;
  assign new_n3083_ = new_n3081_ & new_n3082_;
  assign new_n3084_ = new_n2866_ & ~new_n3020_;
  assign new_n3085_ = \2_n1793  & new_n3069_;
  assign new_n3086_ = new_n3084_ & new_n3085_;
  assign new_n3087_ = new_n3083_ & new_n3086_;
  assign \2_n165  = new_n2761_ & new_n3087_;
  assign new_n3089_ = new_n2107_ & new_n2131_;
  assign \2_n1698  = ~new_n2048_ & new_n3089_;
  assign new_n3091_ = ~new_n2231_ & ~new_n2255_;
  assign new_n3092_ = new_n1941_ & ~new_n2162_;
  assign new_n3093_ = new_n3091_ & new_n3092_;
  assign new_n3094_ = ~new_n2216_ & ~new_n2838_;
  assign new_n3095_ = ~new_n2225_ & ~new_n2915_;
  assign new_n3096_ = new_n3094_ & new_n3095_;
  assign new_n3097_ = new_n3093_ & new_n3096_;
  assign \2_n1708  = new_n2698_ & new_n3097_;
  assign new_n3099_ = new_n1946_ & new_n1963_;
  assign new_n3100_ = new_n1995_ & new_n2017_;
  assign \2_n1721  = new_n3099_ & new_n3100_;
  assign new_n3102_ = \2_n606  & \2_n627 ;
  assign new_n3103_ = \2_n378  & new_n3102_;
  assign new_n3104_ = \2_n387  & \2_n627 ;
  assign new_n3105_ = ~\2_n378  & new_n3104_;
  assign new_n3106_ = ~new_n3103_ & ~new_n3105_;
  assign new_n3107_ = ~\2_n627  & ~\2_n1314 ;
  assign new_n3108_ = ~\2_n378  & new_n3107_;
  assign new_n3109_ = ~\2_n627  & ~\2_n1110 ;
  assign new_n3110_ = \2_n378  & new_n3109_;
  assign new_n3111_ = ~new_n3108_ & ~new_n3110_;
  assign new_n3112_ = new_n3106_ & new_n3111_;
  assign \2_n1733  = \2_n1050 ;
  assign new_n3114_ = \2_n179  & \2_n186 ;
  assign new_n3115_ = \2_n560  & new_n3114_;
  assign new_n3116_ = \2_n186  & \2_n760 ;
  assign new_n3117_ = ~\2_n560  & new_n3116_;
  assign new_n3118_ = ~new_n3115_ & ~new_n3117_;
  assign new_n3119_ = ~\2_n186  & ~\2_n168 ;
  assign new_n3120_ = ~\2_n560  & new_n3119_;
  assign new_n3121_ = ~\2_n186  & ~\2_n1346 ;
  assign new_n3122_ = \2_n560  & new_n3121_;
  assign new_n3123_ = ~new_n3120_ & ~new_n3122_;
  assign \2_n1761  = ~new_n3118_ | ~new_n3123_;
  assign \2_n1780  = \2_n1058  & \2_n84 ;
  assign new_n3126_ = \2_n1205  & \2_n236 ;
  assign new_n3127_ = \2_n228  & new_n3126_;
  assign new_n3128_ = \2_n1205  & \2_n1743 ;
  assign new_n3129_ = ~\2_n228  & new_n3128_;
  assign new_n3130_ = ~new_n3127_ & ~new_n3129_;
  assign new_n3131_ = ~\2_n1205  & ~\2_n1495 ;
  assign new_n3132_ = ~\2_n228  & new_n3131_;
  assign new_n3133_ = ~\2_n1205  & ~\2_n1631 ;
  assign new_n3134_ = \2_n228  & new_n3133_;
  assign new_n3135_ = ~new_n3132_ & ~new_n3134_;
  assign new_n3136_ = new_n3130_ & new_n3135_;
  assign \2_n1784  = \2_n1050 ;
  assign new_n3138_ = \2_n1205  & \2_n1362 ;
  assign new_n3139_ = \2_n228  & new_n3138_;
  assign new_n3140_ = \2_n1205  & \2_n1598 ;
  assign new_n3141_ = ~\2_n228  & new_n3140_;
  assign new_n3142_ = ~new_n3139_ & ~new_n3141_;
  assign new_n3143_ = ~\2_n1205  & ~\2_n487 ;
  assign new_n3144_ = ~\2_n228  & new_n3143_;
  assign new_n3145_ = ~\2_n1205  & ~\2_n1710 ;
  assign new_n3146_ = \2_n228  & new_n3145_;
  assign new_n3147_ = ~new_n3144_ & ~new_n3146_;
  assign new_n3148_ = new_n3142_ & new_n3147_;
  assign \2_n1794  = \2_n1050 ;
  assign new_n3150_ = \2_n186  & \2_n19 ;
  assign new_n3151_ = \2_n560  & new_n3150_;
  assign new_n3152_ = \2_n186  & \2_n955 ;
  assign new_n3153_ = ~\2_n560  & new_n3152_;
  assign new_n3154_ = ~new_n3151_ & ~new_n3153_;
  assign new_n3155_ = ~\2_n186  & ~\2_n964 ;
  assign new_n3156_ = ~\2_n560  & new_n3155_;
  assign new_n3157_ = ~\2_n186  & ~\2_n370 ;
  assign new_n3158_ = \2_n560  & new_n3157_;
  assign new_n3159_ = ~new_n3156_ & ~new_n3158_;
  assign \2_n18  = ~new_n3154_ | ~new_n3159_;
  assign new_n3161_ = \2_n186  & \2_n297 ;
  assign new_n3162_ = \2_n560  & new_n3161_;
  assign new_n3163_ = \2_n186  & \2_n384 ;
  assign new_n3164_ = ~\2_n560  & new_n3163_;
  assign new_n3165_ = ~new_n3162_ & ~new_n3164_;
  assign new_n3166_ = ~\2_n186  & ~\2_n75 ;
  assign new_n3167_ = ~\2_n560  & new_n3166_;
  assign new_n3168_ = ~\2_n186  & ~\2_n1087 ;
  assign new_n3169_ = \2_n560  & new_n3168_;
  assign new_n3170_ = ~new_n3167_ & ~new_n3169_;
  assign \2_n211  = ~new_n3165_ | ~new_n3170_;
  assign new_n3172_ = \2_n627  & \2_n715 ;
  assign new_n3173_ = \2_n378  & new_n3172_;
  assign new_n3174_ = \2_n128  & \2_n627 ;
  assign new_n3175_ = ~\2_n378  & new_n3174_;
  assign new_n3176_ = ~new_n3173_ & ~new_n3175_;
  assign new_n3177_ = ~\2_n627  & ~\2_n964 ;
  assign new_n3178_ = ~\2_n378  & new_n3177_;
  assign new_n3179_ = ~\2_n627  & ~\2_n370 ;
  assign new_n3180_ = \2_n378  & new_n3179_;
  assign new_n3181_ = ~new_n3178_ & ~new_n3180_;
  assign new_n3182_ = new_n3176_ & new_n3181_;
  assign \2_n222  = \2_n1050 ;
  assign new_n3184_ = \2_n1088  & \2_n1281 ;
  assign new_n3185_ = \2_n1219  & ~\2_n1281 ;
  assign new_n3186_ = ~new_n3184_ & ~new_n3185_;
  assign new_n3187_ = ~\2_n117  & new_n3186_;
  assign \2_n245  = \2_n1584 ;
  assign new_n3189_ = \2_n236  & \2_n627 ;
  assign new_n3190_ = \2_n378  & new_n3189_;
  assign new_n3191_ = \2_n1743  & \2_n627 ;
  assign new_n3192_ = ~\2_n378  & new_n3191_;
  assign new_n3193_ = ~new_n3190_ & ~new_n3192_;
  assign new_n3194_ = ~\2_n627  & ~\2_n1495 ;
  assign new_n3195_ = ~\2_n378  & new_n3194_;
  assign new_n3196_ = ~\2_n627  & ~\2_n1631 ;
  assign new_n3197_ = \2_n378  & new_n3196_;
  assign new_n3198_ = ~new_n3195_ & ~new_n3197_;
  assign new_n3199_ = new_n3193_ & new_n3198_;
  assign \2_n249  = \2_n1050 ;
  assign new_n3201_ = \2_n627  & \2_n758 ;
  assign new_n3202_ = \2_n378  & new_n3201_;
  assign new_n3203_ = \2_n1675  & \2_n627 ;
  assign new_n3204_ = ~\2_n378  & new_n3203_;
  assign new_n3205_ = ~new_n3202_ & ~new_n3204_;
  assign new_n3206_ = ~\2_n627  & ~\2_n454 ;
  assign new_n3207_ = ~\2_n378  & new_n3206_;
  assign new_n3208_ = ~\2_n627  & ~\2_n259 ;
  assign new_n3209_ = \2_n378  & new_n3208_;
  assign new_n3210_ = ~new_n3207_ & ~new_n3209_;
  assign new_n3211_ = new_n3205_ & new_n3210_;
  assign \2_n262  = \2_n1050 ;
  assign new_n3213_ = \2_n1503  & \2_n1047 ;
  assign new_n3214_ = \2_n1674  & ~\2_n617 ;
  assign new_n3215_ = ~\2_n1674  & \2_n617 ;
  assign new_n3216_ = ~new_n3214_ & ~new_n3215_;
  assign new_n3217_ = ~\2_n1238  & \2_n1498 ;
  assign new_n3218_ = \2_n1238  & ~\2_n1498 ;
  assign new_n3219_ = ~new_n3217_ & ~new_n3218_;
  assign new_n3220_ = ~new_n3216_ & new_n3219_;
  assign new_n3221_ = new_n3216_ & ~new_n3219_;
  assign new_n3222_ = ~new_n3220_ & ~new_n3221_;
  assign new_n3223_ = ~\2_n1729  & \2_n319 ;
  assign new_n3224_ = \2_n1729  & ~\2_n319 ;
  assign new_n3225_ = ~new_n3223_ & ~new_n3224_;
  assign new_n3226_ = ~new_n3222_ & new_n3225_;
  assign new_n3227_ = new_n3222_ & ~new_n3225_;
  assign new_n3228_ = ~new_n3226_ & ~new_n3227_;
  assign new_n3229_ = ~\2_n1172  & \2_n1553 ;
  assign new_n3230_ = \2_n1172  & ~\2_n1553 ;
  assign new_n3231_ = ~new_n3229_ & ~new_n3230_;
  assign new_n3232_ = \2_n1660  & ~\2_n708 ;
  assign new_n3233_ = ~\2_n1660  & \2_n708 ;
  assign new_n3234_ = ~new_n3232_ & ~new_n3233_;
  assign new_n3235_ = ~new_n3231_ & new_n3234_;
  assign new_n3236_ = new_n3231_ & ~new_n3234_;
  assign new_n3237_ = ~new_n3235_ & ~new_n3236_;
  assign new_n3238_ = ~new_n3228_ & new_n3237_;
  assign new_n3239_ = new_n3228_ & ~new_n3237_;
  assign \2_n878  = new_n3238_ | new_n3239_;
  assign new_n3241_ = \2_n516  & ~\2_n878 ;
  assign new_n3242_ = \2_n119  & new_n3241_;
  assign new_n3243_ = \2_n504  & \2_n64 ;
  assign new_n3244_ = \2_n1674  & ~\2_n504 ;
  assign new_n3245_ = ~new_n3243_ & ~new_n3244_;
  assign new_n3246_ = new_n2101_ & ~new_n3245_;
  assign new_n3247_ = ~new_n2101_ & new_n3245_;
  assign new_n3248_ = ~new_n3246_ & ~new_n3247_;
  assign new_n3249_ = ~new_n2088_ & new_n2095_;
  assign new_n3250_ = new_n2088_ & ~new_n2095_;
  assign new_n3251_ = ~new_n3249_ & ~new_n3250_;
  assign new_n3252_ = ~new_n3248_ & new_n3251_;
  assign new_n3253_ = new_n3248_ & ~new_n3251_;
  assign new_n3254_ = ~new_n3252_ & ~new_n3253_;
  assign new_n3255_ = ~new_n2076_ & new_n2082_;
  assign new_n3256_ = new_n2076_ & ~new_n2082_;
  assign new_n3257_ = ~new_n3255_ & ~new_n3256_;
  assign new_n3258_ = ~new_n3254_ & new_n3257_;
  assign new_n3259_ = new_n3254_ & ~new_n3257_;
  assign new_n3260_ = ~new_n3258_ & ~new_n3259_;
  assign new_n3261_ = new_n2058_ & ~new_n2062_;
  assign new_n3262_ = ~new_n2058_ & new_n2062_;
  assign new_n3263_ = ~new_n3261_ & ~new_n3262_;
  assign new_n3264_ = new_n2045_ & ~new_n2051_;
  assign new_n3265_ = ~new_n2045_ & new_n2051_;
  assign new_n3266_ = ~new_n3264_ & ~new_n3265_;
  assign new_n3267_ = ~new_n3263_ & new_n3266_;
  assign new_n3268_ = new_n3263_ & ~new_n3266_;
  assign new_n3269_ = ~new_n3267_ & ~new_n3268_;
  assign new_n3270_ = ~new_n3260_ & new_n3269_;
  assign new_n3271_ = new_n3260_ & ~new_n3269_;
  assign \2_n547  = new_n3270_ | new_n3271_;
  assign new_n3273_ = new_n1949_ & ~new_n1954_;
  assign new_n3274_ = ~new_n1949_ & new_n1954_;
  assign new_n3275_ = ~new_n3273_ & ~new_n3274_;
  assign new_n3276_ = ~new_n2289_ & new_n3275_;
  assign new_n3277_ = new_n2289_ & ~new_n3275_;
  assign new_n3278_ = ~new_n3276_ & ~new_n3277_;
  assign new_n3279_ = ~new_n1967_ & ~new_n1973_;
  assign new_n3280_ = new_n1967_ & new_n1973_;
  assign new_n3281_ = ~new_n3279_ & ~new_n3280_;
  assign new_n3282_ = \2_n541  & \2_n600 ;
  assign new_n3283_ = ~\2_n600  & \2_n643 ;
  assign new_n3284_ = ~new_n3282_ & ~new_n3283_;
  assign new_n3285_ = new_n1986_ & ~new_n3284_;
  assign new_n3286_ = ~new_n1986_ & new_n3284_;
  assign new_n3287_ = ~new_n3285_ & ~new_n3286_;
  assign new_n3288_ = new_n1980_ & ~new_n1989_;
  assign new_n3289_ = ~new_n1980_ & new_n1989_;
  assign new_n3290_ = ~new_n3288_ & ~new_n3289_;
  assign new_n3291_ = ~new_n3287_ & new_n3290_;
  assign new_n3292_ = new_n3287_ & ~new_n3290_;
  assign new_n3293_ = ~new_n3291_ & ~new_n3292_;
  assign new_n3294_ = ~new_n3281_ & new_n3293_;
  assign new_n3295_ = new_n3281_ & ~new_n3293_;
  assign new_n3296_ = ~new_n3294_ & ~new_n3295_;
  assign new_n3297_ = ~new_n3278_ & new_n3296_;
  assign new_n3298_ = new_n3278_ & ~new_n3296_;
  assign \2_n320  = ~new_n3297_ & ~new_n3298_;
  assign new_n3300_ = ~\2_n1511  & ~\2_n320 ;
  assign new_n3301_ = ~\2_n547  & new_n3300_;
  assign new_n3302_ = new_n3242_ & new_n3301_;
  assign new_n3303_ = \2_n1768  & new_n3302_;
  assign \2_n264  = new_n3213_ & new_n3303_;
  assign new_n3305_ = \2_n1205  & \2_n335 ;
  assign new_n3306_ = \2_n228  & new_n3305_;
  assign new_n3307_ = \2_n1205  & \2_n270 ;
  assign new_n3308_ = ~\2_n228  & new_n3307_;
  assign new_n3309_ = ~new_n3306_ & ~new_n3308_;
  assign new_n3310_ = ~\2_n1205  & ~\2_n882 ;
  assign new_n3311_ = ~\2_n228  & new_n3310_;
  assign new_n3312_ = ~\2_n1205  & ~\2_n456 ;
  assign new_n3313_ = \2_n228  & new_n3312_;
  assign new_n3314_ = ~new_n3311_ & ~new_n3313_;
  assign new_n3315_ = new_n3309_ & new_n3314_;
  assign \2_n315  = \2_n1050 ;
  assign new_n3317_ = \2_n1205  & \2_n758 ;
  assign new_n3318_ = \2_n228  & new_n3317_;
  assign new_n3319_ = \2_n1205  & \2_n1675 ;
  assign new_n3320_ = ~\2_n228  & new_n3319_;
  assign new_n3321_ = ~new_n3318_ & ~new_n3320_;
  assign new_n3322_ = ~\2_n1205  & ~\2_n454 ;
  assign new_n3323_ = ~\2_n228  & new_n3322_;
  assign new_n3324_ = ~\2_n1205  & ~\2_n259 ;
  assign new_n3325_ = \2_n228  & new_n3324_;
  assign new_n3326_ = ~new_n3323_ & ~new_n3325_;
  assign new_n3327_ = new_n3321_ & new_n3326_;
  assign \2_n337  = \2_n1050 ;
  assign new_n3329_ = \2_n261  & \2_n579 ;
  assign new_n3330_ = \2_n132  & \2_n261 ;
  assign new_n3331_ = ~new_n3329_ & ~new_n3330_;
  assign new_n3332_ = ~\2_n261  & new_n2483_;
  assign new_n3333_ = ~new_n2593_ & ~new_n3332_;
  assign \2_n361  = ~new_n3331_ | ~new_n3333_;
  assign new_n3335_ = \2_n1281  & \2_n636 ;
  assign new_n3336_ = ~\2_n1281  & \2_n371 ;
  assign new_n3337_ = ~new_n3335_ & ~new_n3336_;
  assign new_n3338_ = ~\2_n117  & new_n3337_;
  assign \2_n379  = \2_n1584 ;
  assign new_n3340_ = \2_n186  & \2_n564 ;
  assign new_n3341_ = \2_n560  & new_n3340_;
  assign new_n3342_ = \2_n1655  & \2_n186 ;
  assign new_n3343_ = ~\2_n560  & new_n3342_;
  assign new_n3344_ = ~new_n3341_ & ~new_n3343_;
  assign new_n3345_ = ~\2_n186  & ~\2_n1314 ;
  assign new_n3346_ = ~\2_n560  & new_n3345_;
  assign new_n3347_ = ~\2_n186  & ~\2_n1110 ;
  assign new_n3348_ = \2_n560  & new_n3347_;
  assign new_n3349_ = ~new_n3346_ & ~new_n3348_;
  assign \2_n381  = ~new_n3344_ | ~new_n3349_;
  assign new_n3351_ = \2_n1150  & \2_n307 ;
  assign new_n3352_ = \2_n377  & new_n3351_;
  assign new_n3353_ = \2_n307  & \2_n488 ;
  assign new_n3354_ = ~\2_n377  & new_n3353_;
  assign new_n3355_ = ~new_n3352_ & ~new_n3354_;
  assign new_n3356_ = ~\2_n307  & ~\2_n882 ;
  assign new_n3357_ = ~\2_n377  & new_n3356_;
  assign new_n3358_ = ~\2_n307  & ~\2_n456 ;
  assign new_n3359_ = \2_n377  & new_n3358_;
  assign new_n3360_ = ~new_n3357_ & ~new_n3359_;
  assign \2_n413  = ~new_n3355_ | ~new_n3360_;
  assign new_n3362_ = \2_n307  & \2_n754 ;
  assign new_n3363_ = \2_n377  & new_n3362_;
  assign new_n3364_ = \2_n1177  & \2_n307 ;
  assign new_n3365_ = ~\2_n377  & new_n3364_;
  assign new_n3366_ = ~new_n3363_ & ~new_n3365_;
  assign new_n3367_ = ~\2_n307  & ~\2_n1027 ;
  assign new_n3368_ = ~\2_n377  & new_n3367_;
  assign new_n3369_ = ~\2_n307  & ~\2_n123 ;
  assign new_n3370_ = \2_n377  & new_n3369_;
  assign new_n3371_ = ~new_n3368_ & ~new_n3370_;
  assign \2_n417  = ~new_n3366_ | ~new_n3371_;
  assign new_n3373_ = \2_n12  & \2_n1281 ;
  assign new_n3374_ = ~\2_n117  & ~new_n3373_;
  assign new_n3375_ = \2_n1181  & ~\2_n1281 ;
  assign new_n3376_ = new_n3374_ & ~new_n3375_;
  assign \2_n476  = \2_n1584 ;
  assign new_n3378_ = \2_n1205  & \2_n7 ;
  assign new_n3379_ = \2_n228  & new_n3378_;
  assign new_n3380_ = \2_n1180  & \2_n1205 ;
  assign new_n3381_ = ~\2_n228  & new_n3380_;
  assign new_n3382_ = ~new_n3379_ & ~new_n3381_;
  assign new_n3383_ = ~\2_n1205  & ~\2_n168 ;
  assign new_n3384_ = ~\2_n228  & new_n3383_;
  assign new_n3385_ = ~\2_n1205  & ~\2_n1346 ;
  assign new_n3386_ = \2_n228  & new_n3385_;
  assign new_n3387_ = ~new_n3384_ & ~new_n3386_;
  assign new_n3388_ = new_n3382_ & new_n3387_;
  assign \2_n56  = \2_n1050 ;
  assign new_n3390_ = \2_n1362  & \2_n627 ;
  assign new_n3391_ = \2_n378  & new_n3390_;
  assign new_n3392_ = \2_n1598  & \2_n627 ;
  assign new_n3393_ = ~\2_n378  & new_n3392_;
  assign new_n3394_ = ~new_n3391_ & ~new_n3393_;
  assign new_n3395_ = ~\2_n627  & ~\2_n487 ;
  assign new_n3396_ = ~\2_n378  & new_n3395_;
  assign new_n3397_ = ~\2_n627  & ~\2_n1710 ;
  assign new_n3398_ = \2_n378  & new_n3397_;
  assign new_n3399_ = ~new_n3396_ & ~new_n3398_;
  assign new_n3400_ = new_n3394_ & new_n3399_;
  assign \2_n567  = \2_n1050 ;
  assign \2_n574  = ~\2_n1454  | \2_n117 ;
  assign new_n3403_ = \2_n1150  & \2_n186 ;
  assign new_n3404_ = \2_n560  & new_n3403_;
  assign new_n3405_ = \2_n186  & \2_n488 ;
  assign new_n3406_ = ~\2_n560  & new_n3405_;
  assign new_n3407_ = ~new_n3404_ & ~new_n3406_;
  assign new_n3408_ = ~\2_n186  & ~\2_n882 ;
  assign new_n3409_ = ~\2_n560  & new_n3408_;
  assign new_n3410_ = ~\2_n186  & ~\2_n456 ;
  assign new_n3411_ = \2_n560  & new_n3410_;
  assign new_n3412_ = ~new_n3409_ & ~new_n3411_;
  assign \2_n596  = ~new_n3407_ | ~new_n3412_;
  assign new_n3414_ = \2_n1281  & ~\2_n1363 ;
  assign new_n3415_ = ~\2_n1281  & ~\2_n257 ;
  assign new_n3416_ = ~\2_n117  & ~new_n3415_;
  assign \2_n623  = new_n3414_ | ~new_n3416_;
  assign new_n3418_ = \2_n187  & \2_n307 ;
  assign new_n3419_ = \2_n377  & new_n3418_;
  assign new_n3420_ = \2_n1756  & \2_n307 ;
  assign new_n3421_ = ~\2_n377  & new_n3420_;
  assign new_n3422_ = ~new_n3419_ & ~new_n3421_;
  assign new_n3423_ = ~\2_n307  & ~new_n2383_;
  assign new_n3424_ = ~\2_n377  & new_n3423_;
  assign new_n3425_ = ~\2_n307  & ~new_n2596_;
  assign new_n3426_ = \2_n377  & new_n3425_;
  assign new_n3427_ = ~new_n3424_ & ~new_n3426_;
  assign \2_n635  = ~new_n3422_ | ~new_n3427_;
  assign new_n3429_ = \2_n1281  & \2_n403 ;
  assign new_n3430_ = ~\2_n1281  & \2_n1299 ;
  assign new_n3431_ = ~new_n3429_ & ~new_n3430_;
  assign new_n3432_ = ~\2_n117  & new_n3431_;
  assign \2_n649  = \2_n1584 ;
  assign new_n3434_ = \2_n186  & \2_n187 ;
  assign new_n3435_ = \2_n560  & new_n3434_;
  assign new_n3436_ = \2_n1756  & \2_n186 ;
  assign new_n3437_ = ~\2_n560  & new_n3436_;
  assign new_n3438_ = ~new_n3435_ & ~new_n3437_;
  assign new_n3439_ = ~\2_n186  & ~new_n2383_;
  assign new_n3440_ = ~\2_n560  & new_n3439_;
  assign new_n3441_ = ~\2_n186  & ~new_n2596_;
  assign new_n3442_ = \2_n560  & new_n3441_;
  assign new_n3443_ = ~new_n3440_ & ~new_n3442_;
  assign \2_n661  = ~new_n3438_ | ~new_n3443_;
  assign \2_n67  = \2_n1471  & ~\2_n544 ;
  assign new_n3446_ = \2_n297  & \2_n307 ;
  assign new_n3447_ = \2_n377  & new_n3446_;
  assign new_n3448_ = \2_n307  & \2_n384 ;
  assign new_n3449_ = ~\2_n377  & new_n3448_;
  assign new_n3450_ = ~new_n3447_ & ~new_n3449_;
  assign new_n3451_ = ~\2_n307  & ~\2_n75 ;
  assign new_n3452_ = ~\2_n377  & new_n3451_;
  assign new_n3453_ = ~\2_n307  & ~\2_n1087 ;
  assign new_n3454_ = \2_n377  & new_n3453_;
  assign new_n3455_ = ~new_n3452_ & ~new_n3454_;
  assign \2_n722  = ~new_n3450_ | ~new_n3455_;
  assign new_n3457_ = \2_n1205  & \2_n715 ;
  assign new_n3458_ = \2_n228  & new_n3457_;
  assign new_n3459_ = \2_n1205  & \2_n128 ;
  assign new_n3460_ = ~\2_n228  & new_n3459_;
  assign new_n3461_ = ~new_n3458_ & ~new_n3460_;
  assign new_n3462_ = ~\2_n1205  & ~\2_n964 ;
  assign new_n3463_ = ~\2_n228  & new_n3462_;
  assign new_n3464_ = ~\2_n1205  & ~\2_n370 ;
  assign new_n3465_ = \2_n228  & new_n3464_;
  assign new_n3466_ = ~new_n3463_ & ~new_n3465_;
  assign new_n3467_ = new_n3461_ & new_n3466_;
  assign \2_n786  = \2_n1050 ;
  assign new_n3469_ = \2_n307  & \2_n564 ;
  assign new_n3470_ = \2_n377  & new_n3469_;
  assign new_n3471_ = \2_n1655  & \2_n307 ;
  assign new_n3472_ = ~\2_n377  & new_n3471_;
  assign new_n3473_ = ~new_n3470_ & ~new_n3472_;
  assign new_n3474_ = ~\2_n307  & ~\2_n1314 ;
  assign new_n3475_ = ~\2_n377  & new_n3474_;
  assign new_n3476_ = ~\2_n307  & ~\2_n1110 ;
  assign new_n3477_ = \2_n377  & new_n3476_;
  assign new_n3478_ = ~new_n3475_ & ~new_n3477_;
  assign \2_n824  = ~new_n3473_ | ~new_n3478_;
  assign new_n3480_ = \2_n186  & \2_n565 ;
  assign new_n3481_ = \2_n560  & new_n3480_;
  assign new_n3482_ = \2_n1540  & \2_n186 ;
  assign new_n3483_ = ~\2_n560  & new_n3482_;
  assign new_n3484_ = ~new_n3481_ & ~new_n3483_;
  assign new_n3485_ = ~\2_n186  & ~\2_n487 ;
  assign new_n3486_ = ~\2_n560  & new_n3485_;
  assign new_n3487_ = ~\2_n186  & ~\2_n1710 ;
  assign new_n3488_ = \2_n560  & new_n3487_;
  assign new_n3489_ = ~new_n3486_ & ~new_n3488_;
  assign \2_n83  = ~new_n3484_ | ~new_n3489_;
  assign new_n3491_ = \2_n179  & \2_n307 ;
  assign new_n3492_ = \2_n377  & new_n3491_;
  assign new_n3493_ = \2_n307  & \2_n760 ;
  assign new_n3494_ = ~\2_n377  & new_n3493_;
  assign new_n3495_ = ~new_n3492_ & ~new_n3494_;
  assign new_n3496_ = ~\2_n307  & ~\2_n168 ;
  assign new_n3497_ = ~\2_n377  & new_n3496_;
  assign new_n3498_ = ~\2_n307  & ~\2_n1346 ;
  assign new_n3499_ = \2_n377  & new_n3498_;
  assign new_n3500_ = ~new_n3497_ & ~new_n3499_;
  assign \2_n840  = ~new_n3495_ | ~new_n3500_;
  assign new_n3502_ = ~\2_n1793  & new_n2812_;
  assign new_n3503_ = \2_n1793  & ~new_n2812_;
  assign \2_n889  = ~new_n3502_ & ~new_n3503_;
  assign new_n3505_ = \2_n1353  & \2_n627 ;
  assign new_n3506_ = \2_n378  & new_n3505_;
  assign new_n3507_ = \2_n530  & \2_n627 ;
  assign new_n3508_ = ~\2_n378  & new_n3507_;
  assign new_n3509_ = ~new_n3506_ & ~new_n3508_;
  assign new_n3510_ = ~\2_n627  & ~\2_n75 ;
  assign new_n3511_ = ~\2_n378  & new_n3510_;
  assign new_n3512_ = ~\2_n627  & ~\2_n1087 ;
  assign new_n3513_ = \2_n378  & new_n3512_;
  assign new_n3514_ = ~new_n3511_ & ~new_n3513_;
  assign new_n3515_ = new_n3509_ & new_n3514_;
  assign \2_n944  = \2_n1050 ;
  assign new_n3517_ = \2_n1281  & ~\2_n38 ;
  assign new_n3518_ = ~\2_n1281  & ~\2_n1700 ;
  assign new_n3519_ = ~\2_n117  & ~new_n3518_;
  assign \2_n951  = new_n3517_ | ~new_n3519_;
  assign new_n3521_ = \2_n261  & \2_n33 ;
  assign new_n3522_ = ~new_n3329_ & ~new_n3521_;
  assign new_n3523_ = ~\2_n261  & new_n2286_;
  assign new_n3524_ = ~new_n2380_ & ~new_n3523_;
  assign \2_n974  = ~new_n3522_ | ~new_n3524_;
  assign \1_n1547  = ~\1_n842 ;
  assign \1_n1629  = ~\1_n1310 ;
  assign \1_n292  = ~\1_n1134 ;
  assign \1_n350  = ~\1_n128 ;
  assign \1_n476  = ~\1_n1150 ;
  assign \1_n618  = ~\1_n797 ;
  assign \1_n800  = ~\1_n629 ;
  assign \2_n1044  = ~\2_n918 ;
  assign \2_n112  = ~\2_n448 ;
  assign \2_n1140  = ~\2_n1568 ;
  assign \2_n1370  = ~\2_n92 ;
  assign \2_n1464  = ~\2_n389 ;
  assign \2_n1654  = ~\2_n457 ;
  assign \2_n1676  = ~\2_n1338 ;
  assign \2_n193  = ~\2_n937 ;
  assign \2_n357  = ~\2_n566 ;
  assign \2_n61  = ~\2_n1503 ;
  assign \2_n849  = ~\2_n516 ;
  assign \1_n1023  = \1_n1630 ;
  assign \1_n1117  = \1_n110 ;
  assign \1_n1192  = \1_n1134 ;
  assign \1_n1442  = \1_n574 ;
  assign \1_n154  = \1_n478 ;
  assign \1_n1542  = \1_n750 ;
  assign \1_n1552  = \1_n154 ;
  assign \1_n1556  = \1_n1019 ;
  assign \1_n253  = \1_n481 ;
  assign \1_n324  = \1_n1032 ;
  assign \1_n364  = \1_n842 ;
  assign \1_n388  = \1_n1013 ;
  assign \1_n480  = \1_n232 ;
  assign \1_n489  = \1_n350 ;
  assign \1_n565  = \1_n1547 ;
  assign \1_n608  = \1_n1596 ;
  assign \1_n61  = \1_n489 ;
  assign \1_n614  = \1_n142 ;
  assign \1_n663  = \1_n489 ;
  assign \1_n678  = \1_n623 ;
  assign \1_n717  = \1_n1192 ;
  assign \1_n740  = \1_n1026 ;
  assign \1_n786  = \1_n154 ;
  assign \1_n8  = \1_n476 ;
  assign \1_n845  = \1_n489 ;
  assign \2_n1233  = \2_n1044 ;
  assign \2_n129  = \2_n566 ;
  assign \2_n1355  = \2_n288 ;
  assign \2_n1378  = \2_n84 ;
  assign \2_n1425  = \2_n1050 ;
  assign \2_n1657  = \2_n389 ;
  assign \2_n1682  = \2_n130 ;
  assign \2_n1697  = \2_n1414 ;
  assign \2_n173  = \2_n1378 ;
  assign \2_n235  = \2_n1721 ;
  assign \2_n375  = \2_n1378 ;
  assign \2_n542  = \2_n1378 ;
  assign \2_n611  = \2_n1378 ;
  assign \2_n66  = \2_n1657 ;
  assign \2_n673  = \2_n1698 ;
  assign \2_n765  = \2_n1233 ;
  assign \2_n776  = \2_n1584 ;
  assign \2_n793  = \2_n544 ;
  assign \2_n845  = \2_n1584 ;
  assign \2_n860  = \2_n623 ;
  assign \2_n967  = \2_n357 ;
endmodule


