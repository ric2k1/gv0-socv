module top( n4 , n14 , n23 , n25 , n28 , n32 , n34 , n38 , n40 , n50 , n55 , n58 , n59 , n60 , n63 , n65 );
    input n4 , n23 , n25 , n28 , n32 , n38 , n50 , n55 , n58 , n60 , n63 , n65 ;
    output n14 , n34 , n40 , n59 ;
    wire n0 , n1 , n2 , n3 , n5 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n24 , n26 , n27 , n29 , n30 , n31 , n33 , n35 , n36 , n37 , n39 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n51 , n52 , n53 , n54 , n56 , n57 , n61 , n62 , n64 , n66 , n67 , n68 ;
assign n49 = ~(n47 | n13);
assign n12 = ~(n1 ^ n47);
assign n57 = ~(n8 ^ n23);
assign n62 = ~(n0 | n45);
assign n56 = n37 | n44;
assign n22 = ~(n32 & n60);
assign n44 = ~n25;
assign n47 = n3 | n19;
assign n46 = n65 | n61;
assign n33 = n53 | n31;
assign n31 = n3 | n44;
assign n66 = n37 | n36;
assign n2 = ~n58;
assign n11 = ~n7;
assign n51 = ~n32;
assign n9 = ~n5;
assign n68 = ~(n26 ^ n21);
assign n7 = n51 | n44;
assign n42 = ~(n23 | n52);
assign n43 = n27 | n64;
assign n64 = ~(n42 | n8);
assign n35 = ~(n41 ^ n68);
assign n52 = ~n33;
assign n29 = n9 | n24;
assign n21 = n15 | n44;
assign n40 = ~(n30 | n52);
assign n16 = n10 & n7;
assign n53 = ~n4;
assign n45 = n43 & n46;
assign n24 = ~(n56 ^ n12);
assign n15 = ~n55;
assign n26 = n3 | n2;
assign n19 = ~n60;
assign n27 = n23 & n52;
assign n30 = ~(n4 | n39);
assign n37 = ~n63;
assign n48 = ~(n62 ^ n28);
assign n36 = ~n38;
assign n13 = n1 & n56;
assign n39 = ~n31;
assign n18 = ~(n6 ^ n48);
assign n8 = n16 | n5;
assign n67 = ~(n17 | n49);
assign n17 = ~(n1 | n56);
assign n20 = ~(n61 ^ n65);
assign n5 = n54 & n11;
assign n0 = n65 & n61;
assign n14 = ~(n43 ^ n20);
assign n41 = ~(n22 ^ n66);
assign n10 = ~n54;
assign n61 = ~(n5 ^ n24);
assign n1 = n51 | n36;
assign n54 = n50 & n38;
assign n59 = ~(n35 ^ n18);
assign n6 = ~(n67 ^ n29);
assign n3 = ~n50;
assign n34 = ~(n33 ^ n57);
endmodule
