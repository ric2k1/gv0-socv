module alu4_lev2(pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, 
	pi10, pi11, pi12, pi13, po0, po1, po2, po3, po4, po5, po6, po7);

input pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, 
	pi10, pi11, pi12, pi13;

output po0, po1, po2, po3, po4, po5, po6, po7;

wire n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, 
	n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, 
	n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, 
	n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, 
	n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, 
	n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, 
	n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, 
	n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, 
	n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, 
	n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, 
	n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, 
	n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, 
	n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, 
	n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, 
	n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, 
	n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, 
	n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, 
	n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, 
	n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, 
	n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, 
	n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, 
	n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, 
	n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, 
	n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, 
	n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, 
	n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, 
	n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, 
	n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, 
	n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, 
	n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, 
	n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, 
	n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, 
	n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, 
	n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, 
	n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, 
	n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, 
	n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, 
	n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, 
	n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, 
	n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, 
	n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, 
	n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, 
	n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, 
	n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, 
	n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, 
	n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, 
	n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, 
	n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, 
	n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, 
	n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, 
	n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, 
	n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, 
	n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, 
	n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, 
	n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, 
	n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, 
	n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, 
	n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, 
	n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, 
	n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, 
	n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, 
	n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, 
	n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, 
	n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, 
	n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, 
	n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, 
	n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, 
	n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, 
	n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, 
	n1395, n1396;

  AN2 U712 ( .A(n705), .B(po4), .Z(po7));
  OR2 U713 ( .A(n706), .B(n707), .Z(n705));
  AN2 U714 ( .A(n708), .B(n709), .Z(n707));
  OR2 U715 ( .A(n710), .B(n711), .Z(n708));
  AN2 U716 ( .A(n712), .B(n713), .Z(n711));
  AN2 U717 ( .A(n714), .B(n715), .Z(n710));
  AN2 U718 ( .A(n716), .B(n717), .Z(n714));
  AN2 U719 ( .A(n718), .B(n719), .Z(n706));
  OR2 U720 ( .A(n720), .B(n712), .Z(n719));
  OR2 U721 ( .A(n721), .B(n722), .Z(n712));
  AN2 U722 ( .A(n723), .B(n724), .Z(n722));
  AN2 U723 ( .A(n725), .B(n726), .Z(n721));
  OR2 U724 ( .A(n724), .B(n727), .Z(n726));
  AN2 U725 ( .A(n727), .B(n723), .Z(n720));
  OR2 U726 ( .A(n728), .B(n729), .Z(po6));
  AN2 U727 ( .A(pi13), .B(n730), .Z(n729));
  OR2 U728 ( .A(n731), .B(n732), .Z(n730));
  OR2 U729 ( .A(n733), .B(n734), .Z(n732));
  OR2 U730 ( .A(n735), .B(n736), .Z(n734));
  AN2 U731 ( .A(n737), .B(n738), .Z(n736));
  OR2 U732 ( .A(n739), .B(n740), .Z(n737));
  OR2 U733 ( .A(n741), .B(n742), .Z(n740));
  AN2 U734 ( .A(n743), .B(n744), .Z(n742));
  OR2 U735 ( .A(n745), .B(n746), .Z(n743));
  AN2 U736 ( .A(pi03), .B(n747), .Z(n745));
  AN2 U737 ( .A(n748), .B(n749), .Z(n741));
  AN2 U738 ( .A(n750), .B(n751), .Z(n748));
  AN2 U739 ( .A(pi11), .B(n752), .Z(n735));
  OR2 U740 ( .A(n753), .B(n754), .Z(n752));
  OR2 U741 ( .A(n755), .B(n756), .Z(n754));
  AN2 U742 ( .A(n757), .B(n747), .Z(n756));
  OR2 U743 ( .A(n758), .B(n759), .Z(n757));
  IV2 U744 ( .A(n760), .Z(n755));
  AN2 U745 ( .A(n761), .B(n762), .Z(n753));
  OR2 U746 ( .A(n763), .B(po5), .Z(n762));
  AN2 U747 ( .A(n764), .B(n765), .Z(n763));
  AN2 U748 ( .A(n766), .B(n767), .Z(n733));
  OR2 U749 ( .A(n768), .B(n769), .Z(n767));
  AN2 U750 ( .A(n770), .B(n771), .Z(n768));
  IV2 U751 ( .A(n772), .Z(n766));
  OR2 U752 ( .A(n773), .B(n774), .Z(n731));
  AN2 U753 ( .A(n775), .B(n776), .Z(n774));
  AN2 U754 ( .A(n777), .B(n778), .Z(n775));
  AN2 U755 ( .A(n779), .B(n780), .Z(n773));
  AN2 U756 ( .A(n781), .B(n782), .Z(n779));
  AN2 U757 ( .A(n783), .B(n781), .Z(n728));
  AN2 U758 ( .A(n782), .B(n784), .Z(n783));
  OR2 U759 ( .A(n785), .B(n786), .Z(po3));
  OR2 U760 ( .A(n787), .B(n788), .Z(n786));
  OR2 U761 ( .A(n789), .B(n790), .Z(n788));
  OR2 U762 ( .A(n791), .B(n792), .Z(n790));
  AN2 U763 ( .A(n793), .B(n782), .Z(n792));
  AN2 U764 ( .A(n794), .B(n795), .Z(n791));
  OR2 U765 ( .A(n796), .B(n797), .Z(n789));
  IV2 U766 ( .A(n798), .Z(n797));
  OR2 U767 ( .A(n799), .B(n778), .Z(n798));
  AN2 U768 ( .A(n778), .B(n799), .Z(n796));
  OR2 U769 ( .A(n800), .B(n801), .Z(n799));
  IV2 U770 ( .A(n802), .Z(n778));
  OR2 U771 ( .A(n803), .B(n804), .Z(n802));
  AN2 U772 ( .A(n805), .B(n806), .Z(n803));
  AN2 U773 ( .A(n807), .B(n808), .Z(n806));
  AN2 U774 ( .A(n809), .B(n810), .Z(n808));
  OR2 U775 ( .A(pi11), .B(n811), .Z(n810));
  AN2 U776 ( .A(n812), .B(n813), .Z(n811));
  AN2 U777 ( .A(n814), .B(n815), .Z(n813));
  OR2 U778 ( .A(n782), .B(n816), .Z(n815));
  OR2 U779 ( .A(n817), .B(n818), .Z(n814));
  OR2 U780 ( .A(n819), .B(n820), .Z(n818));
  AN2 U781 ( .A(n750), .B(n821), .Z(n820));
  AN2 U782 ( .A(n749), .B(n747), .Z(n819));
  IV2 U783 ( .A(n821), .Z(n749));
  AN2 U784 ( .A(n822), .B(n823), .Z(n812));
  OR2 U785 ( .A(n824), .B(n825), .Z(n823));
  OR2 U786 ( .A(n826), .B(n827), .Z(n822));
  AN2 U787 ( .A(pi10), .B(n828), .Z(n826));
  OR2 U788 ( .A(n829), .B(n830), .Z(n828));
  OR2 U789 ( .A(n831), .B(n738), .Z(n809));
  AN2 U790 ( .A(n832), .B(n833), .Z(n831));
  AN2 U791 ( .A(n834), .B(n760), .Z(n833));
  OR2 U792 ( .A(n817), .B(n835), .Z(n760));
  OR2 U793 ( .A(pi03), .B(n836), .Z(n835));
  OR2 U794 ( .A(n817), .B(n837), .Z(n834));
  OR2 U795 ( .A(n715), .B(n827), .Z(n837));
  IV2 U796 ( .A(n836), .Z(n715));
  AN2 U797 ( .A(n838), .B(n839), .Z(n832));
  OR2 U798 ( .A(n765), .B(n840), .Z(n839));
  OR2 U799 ( .A(n841), .B(n825), .Z(n840));
  OR2 U800 ( .A(n816), .B(n842), .Z(n838));
  OR2 U801 ( .A(n843), .B(n844), .Z(n842));
  AN2 U802 ( .A(n845), .B(n846), .Z(n844));
  OR2 U803 ( .A(n847), .B(n848), .Z(n845));
  AN2 U804 ( .A(n758), .B(n747), .Z(n848));
  IV2 U805 ( .A(n849), .Z(n758));
  AN2 U806 ( .A(n750), .B(n849), .Z(n847));
  AN2 U807 ( .A(n849), .B(n759), .Z(n843));
  OR2 U808 ( .A(n850), .B(n851), .Z(n849));
  AN2 U809 ( .A(n852), .B(n853), .Z(n850));
  IV2 U810 ( .A(n854), .Z(n816));
  AN2 U811 ( .A(n855), .B(n856), .Z(n807));
  OR2 U812 ( .A(n857), .B(n858), .Z(n856));
  OR2 U813 ( .A(n859), .B(n860), .Z(n858));
  AN2 U814 ( .A(n861), .B(n739), .Z(n859));
  OR2 U815 ( .A(n862), .B(n863), .Z(n739));
  AN2 U816 ( .A(n759), .B(n795), .Z(n862));
  OR2 U817 ( .A(n846), .B(n864), .Z(n861));
  IV2 U818 ( .A(n865), .Z(n864));
  AN2 U819 ( .A(n795), .B(n863), .Z(n865));
  IV2 U820 ( .A(n759), .Z(n846));
  OR2 U821 ( .A(n866), .B(n867), .Z(n759));
  AN2 U822 ( .A(n868), .B(po5), .Z(n867));
  AN2 U823 ( .A(n750), .B(n869), .Z(n866));
  OR2 U824 ( .A(n825), .B(n870), .Z(n855));
  OR2 U825 ( .A(n871), .B(n872), .Z(n870));
  AN2 U826 ( .A(n764), .B(n873), .Z(n872));
  IV2 U827 ( .A(po5), .Z(n873));
  AN2 U828 ( .A(n841), .B(po4), .Z(n871));
  OR2 U829 ( .A(n874), .B(po5), .Z(po4));
  IV2 U830 ( .A(n764), .Z(n841));
  OR2 U831 ( .A(n875), .B(n724), .Z(n764));
  AN2 U832 ( .A(n876), .B(n877), .Z(n875));
  AN2 U833 ( .A(n878), .B(n879), .Z(n805));
  AN2 U834 ( .A(n880), .B(n881), .Z(n879));
  OR2 U835 ( .A(n782), .B(n882), .Z(n881));
  OR2 U836 ( .A(n781), .B(n883), .Z(n882));
  IV2 U837 ( .A(n884), .Z(n781));
  OR2 U838 ( .A(n795), .B(n885), .Z(n880));
  AN2 U839 ( .A(n886), .B(n887), .Z(n878));
  OR2 U840 ( .A(pi03), .B(n888), .Z(n887));
  AN2 U841 ( .A(n889), .B(n890), .Z(n888));
  IV2 U842 ( .A(n891), .Z(n890));
  AN2 U843 ( .A(n830), .B(n892), .Z(n891));
  OR2 U844 ( .A(n893), .B(n894), .Z(n830));
  IV2 U845 ( .A(n895), .Z(n894));
  OR2 U846 ( .A(n746), .B(n750), .Z(n895));
  AN2 U847 ( .A(n750), .B(n746), .Z(n893));
  OR2 U848 ( .A(n896), .B(n897), .Z(n746));
  AN2 U849 ( .A(pi02), .B(n898), .Z(n896));
  IV2 U850 ( .A(n747), .Z(n750));
  OR2 U851 ( .A(n899), .B(n900), .Z(n747));
  AN2 U852 ( .A(n901), .B(n771), .Z(n900));
  OR2 U853 ( .A(pi03), .B(n795), .Z(n771));
  AN2 U854 ( .A(n902), .B(n903), .Z(n899));
  OR2 U855 ( .A(n904), .B(n905), .Z(n903));
  OR2 U856 ( .A(n906), .B(n907), .Z(n905));
  AN2 U857 ( .A(n782), .B(n892), .Z(n907));
  AN2 U858 ( .A(n769), .B(n751), .Z(n906));
  AN2 U859 ( .A(po5), .B(n908), .Z(n904));
  OR2 U860 ( .A(n909), .B(n772), .Z(n889));
  AN2 U861 ( .A(n910), .B(n911), .Z(n909));
  OR2 U862 ( .A(n912), .B(n795), .Z(n911));
  OR2 U863 ( .A(n782), .B(n770), .Z(n910));
  OR2 U864 ( .A(n827), .B(n913), .Z(n886));
  OR2 U865 ( .A(n914), .B(n772), .Z(n913));
  OR2 U866 ( .A(n915), .B(n916), .Z(n914));
  AN2 U867 ( .A(n912), .B(n795), .Z(n916));
  IV2 U868 ( .A(n770), .Z(n912));
  AN2 U869 ( .A(n782), .B(n770), .Z(n915));
  OR2 U870 ( .A(n917), .B(n918), .Z(n770));
  AN2 U871 ( .A(n919), .B(n920), .Z(n917));
  IV2 U872 ( .A(n795), .Z(n782));
  OR2 U873 ( .A(n921), .B(n922), .Z(n787));
  AN2 U874 ( .A(n923), .B(n824), .Z(n922));
  AN2 U875 ( .A(n924), .B(n925), .Z(n923));
  OR2 U876 ( .A(n926), .B(n927), .Z(n925));
  AN2 U877 ( .A(pi11), .B(pi03), .Z(n926));
  AN2 U878 ( .A(pi07), .B(n928), .Z(n921));
  OR2 U879 ( .A(n929), .B(n930), .Z(n928));
  AN2 U880 ( .A(n931), .B(n804), .Z(n929));
  OR2 U881 ( .A(n932), .B(n933), .Z(n931));
  AN2 U882 ( .A(n854), .B(n795), .Z(n933));
  AN2 U883 ( .A(n934), .B(n827), .Z(n932));
  OR2 U884 ( .A(n935), .B(n936), .Z(n785));
  OR2 U885 ( .A(n937), .B(n938), .Z(n936));
  AN2 U886 ( .A(n939), .B(n940), .Z(n938));
  OR2 U887 ( .A(n941), .B(n942), .Z(n940));
  OR2 U888 ( .A(n769), .B(n943), .Z(n942));
  AN2 U889 ( .A(n874), .B(n944), .Z(n943));
  AN2 U890 ( .A(n795), .B(pi03), .Z(n769));
  OR2 U891 ( .A(n945), .B(n946), .Z(n795));
  OR2 U892 ( .A(n947), .B(n948), .Z(n946));
  AN2 U893 ( .A(n949), .B(n824), .Z(n948));
  AN2 U894 ( .A(n950), .B(n765), .Z(n947));
  IV2 U895 ( .A(n874), .Z(n765));
  OR2 U896 ( .A(n951), .B(n952), .Z(n945));
  OR2 U897 ( .A(n953), .B(n954), .Z(n952));
  AN2 U898 ( .A(n955), .B(n827), .Z(n954));
  OR2 U899 ( .A(n956), .B(n957), .Z(n955));
  AN2 U900 ( .A(n958), .B(n784), .Z(n956));
  AN2 U901 ( .A(pi07), .B(n959), .Z(n958));
  AN2 U902 ( .A(po5), .B(n960), .Z(n953));
  OR2 U903 ( .A(n961), .B(n962), .Z(n960));
  AN2 U904 ( .A(n892), .B(n963), .Z(n962));
  AN2 U905 ( .A(n964), .B(n965), .Z(n961));
  AN2 U906 ( .A(pi13), .B(n966), .Z(n951));
  OR2 U907 ( .A(n967), .B(n968), .Z(n966));
  OR2 U908 ( .A(n969), .B(n970), .Z(n968));
  AN2 U909 ( .A(n971), .B(pi02), .Z(n970));
  AN2 U910 ( .A(n972), .B(n973), .Z(n969));
  AN2 U911 ( .A(n974), .B(n975), .Z(n972));
  OR2 U912 ( .A(n874), .B(n959), .Z(n975));
  AN2 U913 ( .A(n827), .B(n824), .Z(n874));
  IV2 U914 ( .A(pi03), .Z(n827));
  OR2 U915 ( .A(n964), .B(n976), .Z(n974));
  AN2 U916 ( .A(pi03), .B(n824), .Z(n976));
  IV2 U917 ( .A(pi07), .Z(n824));
  IV2 U918 ( .A(n959), .Z(n964));
  OR2 U919 ( .A(n977), .B(n978), .Z(n959));
  AN2 U920 ( .A(n979), .B(pi02), .Z(n978));
  AN2 U921 ( .A(n980), .B(n717), .Z(n977));
  OR2 U922 ( .A(n979), .B(pi02), .Z(n980));
  AN2 U923 ( .A(n981), .B(po5), .Z(n967));
  AN2 U924 ( .A(po5), .B(n982), .Z(n941));
  AN2 U925 ( .A(pi03), .B(pi07), .Z(po5));
  AN2 U926 ( .A(n983), .B(pi03), .Z(n935));
  OR2 U927 ( .A(n984), .B(n985), .Z(po2));
  OR2 U928 ( .A(n986), .B(n987), .Z(n985));
  OR2 U929 ( .A(n988), .B(n989), .Z(n987));
  OR2 U930 ( .A(n990), .B(n991), .Z(n989));
  AN2 U931 ( .A(n793), .B(n992), .Z(n991));
  AN2 U932 ( .A(n794), .B(n993), .Z(n990));
  OR2 U933 ( .A(n994), .B(n995), .Z(n988));
  AN2 U934 ( .A(n777), .B(n801), .Z(n995));
  IV2 U935 ( .A(n800), .Z(n777));
  AN2 U936 ( .A(n776), .B(n800), .Z(n994));
  OR2 U937 ( .A(n996), .B(n804), .Z(n800));
  AN2 U938 ( .A(n997), .B(n998), .Z(n996));
  AN2 U939 ( .A(n999), .B(n1000), .Z(n998));
  AN2 U940 ( .A(n1001), .B(n1002), .Z(n1000));
  OR2 U941 ( .A(n1003), .B(n817), .Z(n1002));
  AN2 U942 ( .A(n1004), .B(n836), .Z(n1003));
  OR2 U943 ( .A(pi00), .B(n1005), .Z(n836));
  OR2 U944 ( .A(pi02), .B(pi01), .Z(n1005));
  AN2 U945 ( .A(n1006), .B(n1007), .Z(n1004));
  OR2 U946 ( .A(pi11), .B(n1008), .Z(n1007));
  AN2 U947 ( .A(n1009), .B(n821), .Z(n1008));
  OR2 U948 ( .A(n898), .B(n1010), .Z(n821));
  OR2 U949 ( .A(n1011), .B(n851), .Z(n1009));
  AN2 U950 ( .A(n1012), .B(n1013), .Z(n1011));
  OR2 U951 ( .A(n738), .B(n1014), .Z(n1006));
  OR2 U952 ( .A(n1015), .B(n1016), .Z(n1014));
  AN2 U953 ( .A(n713), .B(n1017), .Z(n1015));
  OR2 U954 ( .A(n1018), .B(n1019), .Z(n1001));
  OR2 U955 ( .A(n744), .B(n1020), .Z(n1019));
  OR2 U956 ( .A(n1021), .B(n1022), .Z(n1018));
  AN2 U957 ( .A(n717), .B(n1023), .Z(n1022));
  AN2 U958 ( .A(n863), .B(n1024), .Z(n1021));
  OR2 U959 ( .A(n1025), .B(n1026), .Z(n1024));
  OR2 U960 ( .A(n992), .B(n852), .Z(n1026));
  IV2 U961 ( .A(n1027), .Z(n1025));
  OR2 U962 ( .A(n1028), .B(n1027), .Z(n863));
  OR2 U963 ( .A(n1029), .B(n1030), .Z(n1027));
  AN2 U964 ( .A(n1031), .B(n1032), .Z(n1029));
  AN2 U965 ( .A(n1033), .B(n993), .Z(n1028));
  AN2 U966 ( .A(n885), .B(n1034), .Z(n999));
  OR2 U967 ( .A(n825), .B(n1035), .Z(n1034));
  OR2 U968 ( .A(n1036), .B(n1037), .Z(n1035));
  AN2 U969 ( .A(n1038), .B(n1039), .Z(n1037));
  IV2 U970 ( .A(n724), .Z(n1039));
  OR2 U971 ( .A(n877), .B(n738), .Z(n1038));
  IV2 U972 ( .A(n876), .Z(n1036));
  OR2 U973 ( .A(n1040), .B(n884), .Z(n885));
  OR2 U974 ( .A(n1041), .B(n1042), .Z(n884));
  OR2 U975 ( .A(n993), .B(n1032), .Z(n1042));
  AN2 U976 ( .A(n1043), .B(n1044), .Z(n997));
  AN2 U977 ( .A(n1045), .B(n1046), .Z(n1044));
  OR2 U978 ( .A(pi02), .B(n1047), .Z(n1046));
  AN2 U979 ( .A(n1048), .B(n1049), .Z(n1047));
  OR2 U980 ( .A(n876), .B(n1050), .Z(n1049));
  OR2 U981 ( .A(n717), .B(n825), .Z(n1050));
  AN2 U982 ( .A(n1051), .B(n1052), .Z(n1048));
  OR2 U983 ( .A(n1053), .B(n1054), .Z(n1052));
  OR2 U984 ( .A(n1055), .B(n772), .Z(n1051));
  AN2 U985 ( .A(n1056), .B(n1057), .Z(n1055));
  OR2 U986 ( .A(n1058), .B(n993), .Z(n1057));
  OR2 U987 ( .A(n992), .B(n919), .Z(n1056));
  OR2 U988 ( .A(n1059), .B(n1016), .Z(n1045));
  AN2 U989 ( .A(n1060), .B(n1061), .Z(n1059));
  AN2 U990 ( .A(n1062), .B(n1063), .Z(n1061));
  OR2 U991 ( .A(n876), .B(n1064), .Z(n1062));
  OR2 U992 ( .A(pi06), .B(n825), .Z(n1064));
  OR2 U993 ( .A(n1065), .B(n725), .Z(n876));
  AN2 U994 ( .A(n718), .B(n1066), .Z(n1065));
  AN2 U995 ( .A(n1067), .B(n1068), .Z(n1060));
  OR2 U996 ( .A(n772), .B(n1069), .Z(n1068));
  OR2 U997 ( .A(n1070), .B(n1071), .Z(n1069));
  AN2 U998 ( .A(n1058), .B(n993), .Z(n1071));
  IV2 U999 ( .A(n919), .Z(n1058));
  AN2 U1000 ( .A(n992), .B(n919), .Z(n1070));
  OR2 U1001 ( .A(n1072), .B(n1073), .Z(n919));
  AN2 U1002 ( .A(n1074), .B(n1075), .Z(n1072));
  OR2 U1003 ( .A(n1054), .B(n1076), .Z(n1067));
  IV2 U1004 ( .A(n1053), .Z(n1076));
  AN2 U1005 ( .A(n1077), .B(n1078), .Z(n1053));
  OR2 U1006 ( .A(n897), .B(n851), .Z(n1078));
  IV2 U1007 ( .A(n1079), .Z(n1077));
  AN2 U1008 ( .A(n851), .B(n897), .Z(n1079));
  OR2 U1009 ( .A(n1080), .B(n1081), .Z(n897));
  AN2 U1010 ( .A(pi01), .B(n1082), .Z(n1080));
  AN2 U1011 ( .A(n1083), .B(n1084), .Z(n1043));
  OR2 U1012 ( .A(pi10), .B(n1085), .Z(n1084));
  OR2 U1013 ( .A(n1086), .B(n1087), .Z(n1085));
  AN2 U1014 ( .A(n1088), .B(n1089), .Z(n1087));
  AN2 U1015 ( .A(n852), .B(n898), .Z(n1088));
  IV2 U1016 ( .A(n1033), .Z(n852));
  AN2 U1017 ( .A(n1090), .B(n853), .Z(n1086));
  IV2 U1018 ( .A(n1089), .Z(n853));
  AN2 U1019 ( .A(n1091), .B(n1082), .Z(n1089));
  OR2 U1020 ( .A(n1031), .B(n1092), .Z(n1091));
  OR2 U1021 ( .A(n851), .B(n1033), .Z(n1090));
  OR2 U1022 ( .A(n1093), .B(n1094), .Z(n1033));
  AN2 U1023 ( .A(n868), .B(n724), .Z(n1094));
  AN2 U1024 ( .A(n851), .B(n869), .Z(n1093));
  IV2 U1025 ( .A(n898), .Z(n851));
  OR2 U1026 ( .A(n1095), .B(n1096), .Z(n898));
  AN2 U1027 ( .A(n901), .B(n920), .Z(n1096));
  OR2 U1028 ( .A(pi02), .B(n993), .Z(n920));
  AN2 U1029 ( .A(n902), .B(n1097), .Z(n1095));
  OR2 U1030 ( .A(n1098), .B(n1099), .Z(n1097));
  OR2 U1031 ( .A(n1100), .B(n1101), .Z(n1099));
  AN2 U1032 ( .A(n992), .B(n892), .Z(n1101));
  AN2 U1033 ( .A(n918), .B(n751), .Z(n1100));
  AN2 U1034 ( .A(n908), .B(n724), .Z(n1098));
  OR2 U1035 ( .A(n1102), .B(n992), .Z(n1083));
  IV2 U1036 ( .A(n993), .Z(n992));
  AN2 U1037 ( .A(n1103), .B(n1104), .Z(n1102));
  OR2 U1038 ( .A(n883), .B(n1105), .Z(n1104));
  IV2 U1039 ( .A(n1106), .Z(n883));
  IV2 U1040 ( .A(n801), .Z(n776));
  OR2 U1041 ( .A(n1107), .B(n1108), .Z(n801));
  OR2 U1042 ( .A(pi12), .B(n1109), .Z(n1108));
  OR2 U1043 ( .A(n1110), .B(n1111), .Z(n986));
  AN2 U1044 ( .A(n1112), .B(n717), .Z(n1111));
  AN2 U1045 ( .A(n924), .B(n1113), .Z(n1112));
  OR2 U1046 ( .A(n1114), .B(n927), .Z(n1113));
  AN2 U1047 ( .A(pi11), .B(pi02), .Z(n1114));
  AN2 U1048 ( .A(pi06), .B(n1115), .Z(n1110));
  OR2 U1049 ( .A(n1116), .B(n930), .Z(n1115));
  AN2 U1050 ( .A(n1117), .B(n804), .Z(n1116));
  OR2 U1051 ( .A(n1118), .B(n1119), .Z(n1117));
  AN2 U1052 ( .A(n854), .B(n993), .Z(n1119));
  AN2 U1053 ( .A(n934), .B(n1016), .Z(n1118));
  OR2 U1054 ( .A(n1120), .B(n1121), .Z(n984));
  OR2 U1055 ( .A(n937), .B(n1122), .Z(n1121));
  AN2 U1056 ( .A(n939), .B(n1123), .Z(n1122));
  OR2 U1057 ( .A(n1124), .B(n1125), .Z(n1123));
  OR2 U1058 ( .A(n918), .B(n1126), .Z(n1125));
  AN2 U1059 ( .A(n724), .B(n982), .Z(n1126));
  AN2 U1060 ( .A(n993), .B(pi02), .Z(n918));
  OR2 U1061 ( .A(n1127), .B(n1128), .Z(n993));
  OR2 U1062 ( .A(n1129), .B(n1130), .Z(n1128));
  AN2 U1063 ( .A(n949), .B(n717), .Z(n1130));
  AN2 U1064 ( .A(n950), .B(n877), .Z(n1129));
  IV2 U1065 ( .A(n727), .Z(n877));
  OR2 U1066 ( .A(n1131), .B(n1132), .Z(n1127));
  OR2 U1067 ( .A(n1133), .B(n1134), .Z(n1132));
  AN2 U1068 ( .A(n1135), .B(n1016), .Z(n1134));
  OR2 U1069 ( .A(n1136), .B(n957), .Z(n1135));
  AN2 U1070 ( .A(n1137), .B(n979), .Z(n1136));
  AN2 U1071 ( .A(n784), .B(pi06), .Z(n1137));
  AN2 U1072 ( .A(n724), .B(n1138), .Z(n1133));
  OR2 U1073 ( .A(n1139), .B(n1140), .Z(n1138));
  AN2 U1074 ( .A(n965), .B(n1141), .Z(n1139));
  AN2 U1075 ( .A(pi02), .B(pi06), .Z(n724));
  AN2 U1076 ( .A(pi13), .B(n1142), .Z(n1131));
  OR2 U1077 ( .A(n1143), .B(n1144), .Z(n1142));
  AN2 U1078 ( .A(n971), .B(pi01), .Z(n1144));
  AN2 U1079 ( .A(n1145), .B(n973), .Z(n1143));
  AN2 U1080 ( .A(n1146), .B(n1147), .Z(n1145));
  OR2 U1081 ( .A(n727), .B(n979), .Z(n1147));
  IV2 U1082 ( .A(n1141), .Z(n979));
  OR2 U1083 ( .A(n1148), .B(n1141), .Z(n1146));
  OR2 U1084 ( .A(n1149), .B(n1150), .Z(n1141));
  AN2 U1085 ( .A(n1151), .B(n1017), .Z(n1150));
  AN2 U1086 ( .A(pi05), .B(n1152), .Z(n1149));
  OR2 U1087 ( .A(n1151), .B(n1017), .Z(n1152));
  AN2 U1088 ( .A(pi02), .B(n717), .Z(n1148));
  AN2 U1089 ( .A(n944), .B(n727), .Z(n1124));
  AN2 U1090 ( .A(n1016), .B(n717), .Z(n727));
  IV2 U1091 ( .A(pi06), .Z(n717));
  IV2 U1092 ( .A(pi02), .Z(n1016));
  AN2 U1093 ( .A(n983), .B(pi02), .Z(n1120));
  OR2 U1094 ( .A(n1153), .B(n1154), .Z(po1));
  OR2 U1095 ( .A(n1155), .B(n1156), .Z(n1154));
  OR2 U1096 ( .A(n1157), .B(n1158), .Z(n1156));
  OR2 U1097 ( .A(n1159), .B(n1160), .Z(n1158));
  AN2 U1098 ( .A(n793), .B(n1105), .Z(n1160));
  AN2 U1099 ( .A(n794), .B(n1032), .Z(n1159));
  OR2 U1100 ( .A(n1161), .B(n1162), .Z(n1157));
  AN2 U1101 ( .A(n1163), .B(n1107), .Z(n1162));
  IV2 U1102 ( .A(n1164), .Z(n1161));
  OR2 U1103 ( .A(n1107), .B(n1163), .Z(n1164));
  AN2 U1104 ( .A(n1165), .B(n1166), .Z(n1163));
  OR2 U1105 ( .A(n1167), .B(n804), .Z(n1107));
  AN2 U1106 ( .A(n1168), .B(n1169), .Z(n1167));
  AN2 U1107 ( .A(n1170), .B(n1171), .Z(n1169));
  OR2 U1108 ( .A(n817), .B(n1172), .Z(n1171));
  OR2 U1109 ( .A(pi11), .B(n1173), .Z(n1172));
  AN2 U1110 ( .A(n1010), .B(n1174), .Z(n1173));
  OR2 U1111 ( .A(n1012), .B(n1013), .Z(n1174));
  OR2 U1112 ( .A(n1175), .B(n1082), .Z(n1010));
  AN2 U1113 ( .A(n1176), .B(n1177), .Z(n1170));
  OR2 U1114 ( .A(pi10), .B(n1178), .Z(n1177));
  OR2 U1115 ( .A(n1179), .B(n1180), .Z(n1178));
  AN2 U1116 ( .A(n1181), .B(n1031), .Z(n1180));
  IV2 U1117 ( .A(n1182), .Z(n1179));
  OR2 U1118 ( .A(n1181), .B(n1031), .Z(n1182));
  OR2 U1119 ( .A(n1183), .B(n1184), .Z(n1181));
  AN2 U1120 ( .A(n1185), .B(n1082), .Z(n1184));
  AN2 U1121 ( .A(n1012), .B(n1092), .Z(n1183));
  OR2 U1122 ( .A(n825), .B(n1186), .Z(n1176));
  OR2 U1123 ( .A(n1187), .B(n1188), .Z(n1186));
  AN2 U1124 ( .A(n1189), .B(n1190), .Z(n1187));
  IV2 U1125 ( .A(n725), .Z(n1190));
  OR2 U1126 ( .A(n1066), .B(n738), .Z(n1189));
  AN2 U1127 ( .A(n1191), .B(n1192), .Z(n1168));
  AN2 U1128 ( .A(n1193), .B(n1194), .Z(n1192));
  OR2 U1129 ( .A(n1195), .B(n1017), .Z(n1194));
  AN2 U1130 ( .A(n1196), .B(n1197), .Z(n1195));
  AN2 U1131 ( .A(n1198), .B(n1199), .Z(n1197));
  OR2 U1132 ( .A(pi05), .B(n1200), .Z(n1199));
  AN2 U1133 ( .A(n1201), .B(n1063), .Z(n1198));
  OR2 U1134 ( .A(n1202), .B(n772), .Z(n1201));
  AN2 U1135 ( .A(n1203), .B(n1204), .Z(n1202));
  OR2 U1136 ( .A(n1074), .B(n1032), .Z(n1204));
  OR2 U1137 ( .A(n1105), .B(n1205), .Z(n1203));
  AN2 U1138 ( .A(n1206), .B(n1207), .Z(n1196));
  OR2 U1139 ( .A(n1208), .B(n1054), .Z(n1207));
  AN2 U1140 ( .A(n1209), .B(n1210), .Z(n1208));
  OR2 U1141 ( .A(n1081), .B(n1082), .Z(n1210));
  OR2 U1142 ( .A(n1012), .B(n1211), .Z(n1209));
  IV2 U1143 ( .A(n1081), .Z(n1211));
  OR2 U1144 ( .A(n817), .B(n1212), .Z(n1206));
  OR2 U1145 ( .A(n713), .B(n738), .Z(n1212));
  OR2 U1146 ( .A(pi01), .B(n1213), .Z(n1193));
  AN2 U1147 ( .A(n1214), .B(n1215), .Z(n1213));
  AN2 U1148 ( .A(n1216), .B(n1217), .Z(n1215));
  OR2 U1149 ( .A(n1054), .B(n1218), .Z(n1216));
  OR2 U1150 ( .A(n1012), .B(n1081), .Z(n1218));
  AN2 U1151 ( .A(pi00), .B(n1175), .Z(n1081));
  OR2 U1152 ( .A(pi08), .B(n1020), .Z(n1054));
  AN2 U1153 ( .A(n1219), .B(n1220), .Z(n1214));
  OR2 U1154 ( .A(n772), .B(n1221), .Z(n1220));
  OR2 U1155 ( .A(n1222), .B(n1223), .Z(n1221));
  AN2 U1156 ( .A(n1074), .B(n1032), .Z(n1223));
  AN2 U1157 ( .A(n1105), .B(n1205), .Z(n1222));
  OR2 U1158 ( .A(n1224), .B(n738), .Z(n772));
  AN2 U1159 ( .A(n1225), .B(n829), .Z(n1224));
  OR2 U1160 ( .A(n751), .B(n1023), .Z(n1225));
  OR2 U1161 ( .A(n716), .B(n1200), .Z(n1219));
  OR2 U1162 ( .A(n718), .B(n825), .Z(n1200));
  IV2 U1163 ( .A(n761), .Z(n825));
  AN2 U1164 ( .A(n1226), .B(n1227), .Z(n1191));
  OR2 U1165 ( .A(n1228), .B(n1229), .Z(n1227));
  OR2 U1166 ( .A(n1020), .B(n1230), .Z(n1229));
  OR2 U1167 ( .A(n1231), .B(n1232), .Z(n1230));
  AN2 U1168 ( .A(n1233), .B(n1234), .Z(n1232));
  AN2 U1169 ( .A(n1235), .B(n1031), .Z(n1233));
  OR2 U1170 ( .A(n1030), .B(n1032), .Z(n1235));
  AN2 U1171 ( .A(n1092), .B(n1041), .Z(n1030));
  IV2 U1172 ( .A(n1236), .Z(n1231));
  OR2 U1173 ( .A(n1234), .B(n1031), .Z(n1236));
  OR2 U1174 ( .A(n1237), .B(n1238), .Z(n1031));
  AN2 U1175 ( .A(n868), .B(n725), .Z(n1238));
  AN2 U1176 ( .A(n1012), .B(n869), .Z(n1237));
  IV2 U1177 ( .A(n1082), .Z(n1012));
  OR2 U1178 ( .A(n1239), .B(n1240), .Z(n1082));
  AN2 U1179 ( .A(n901), .B(n1075), .Z(n1240));
  OR2 U1180 ( .A(pi01), .B(n1032), .Z(n1075));
  AN2 U1181 ( .A(n902), .B(n1241), .Z(n1239));
  OR2 U1182 ( .A(n1242), .B(n1243), .Z(n1241));
  OR2 U1183 ( .A(n1244), .B(n1245), .Z(n1243));
  AN2 U1184 ( .A(n1105), .B(n892), .Z(n1245));
  AN2 U1185 ( .A(n1073), .B(n751), .Z(n1244));
  AN2 U1186 ( .A(n908), .B(n725), .Z(n1242));
  OR2 U1187 ( .A(n1185), .B(n1246), .Z(n1234));
  OR2 U1188 ( .A(n1247), .B(n1105), .Z(n1246));
  IV2 U1189 ( .A(n1248), .Z(n1020));
  OR2 U1190 ( .A(n1249), .B(n744), .Z(n1228));
  AN2 U1191 ( .A(n716), .B(n1023), .Z(n1249));
  AN2 U1192 ( .A(n1250), .B(n1251), .Z(n1226));
  OR2 U1193 ( .A(n1105), .B(n1103), .Z(n1251));
  IV2 U1194 ( .A(n1252), .Z(n1103));
  OR2 U1195 ( .A(n1253), .B(n1254), .Z(n1252));
  AN2 U1196 ( .A(n1106), .B(n1041), .Z(n1254));
  OR2 U1197 ( .A(n1255), .B(n780), .Z(n1106));
  AN2 U1198 ( .A(n973), .B(n738), .Z(n1255));
  AN2 U1199 ( .A(n854), .B(n738), .Z(n1253));
  IV2 U1200 ( .A(n1032), .Z(n1105));
  OR2 U1201 ( .A(n1032), .B(n1256), .Z(n1250));
  OR2 U1202 ( .A(n1040), .B(n1041), .Z(n1256));
  IV2 U1203 ( .A(n1257), .Z(n1040));
  OR2 U1204 ( .A(n1258), .B(n1259), .Z(n1155));
  AN2 U1205 ( .A(n1260), .B(n716), .Z(n1259));
  AN2 U1206 ( .A(n924), .B(n1261), .Z(n1260));
  OR2 U1207 ( .A(n1262), .B(n927), .Z(n1261));
  AN2 U1208 ( .A(pi11), .B(pi01), .Z(n1262));
  AN2 U1209 ( .A(pi05), .B(n1263), .Z(n1258));
  OR2 U1210 ( .A(n1264), .B(n930), .Z(n1263));
  AN2 U1211 ( .A(n1265), .B(n804), .Z(n1264));
  OR2 U1212 ( .A(n1266), .B(n1267), .Z(n1265));
  AN2 U1213 ( .A(n854), .B(n1032), .Z(n1267));
  AN2 U1214 ( .A(n934), .B(n1017), .Z(n1266));
  AN2 U1215 ( .A(pi11), .B(n761), .Z(n934));
  OR2 U1216 ( .A(n1268), .B(n1269), .Z(n1153));
  OR2 U1217 ( .A(n937), .B(n1270), .Z(n1269));
  AN2 U1218 ( .A(n939), .B(n1271), .Z(n1270));
  OR2 U1219 ( .A(n1272), .B(n1273), .Z(n1271));
  OR2 U1220 ( .A(n1073), .B(n1274), .Z(n1273));
  AN2 U1221 ( .A(n725), .B(n982), .Z(n1274));
  AN2 U1222 ( .A(n1032), .B(pi01), .Z(n1073));
  OR2 U1223 ( .A(n1275), .B(n1276), .Z(n1032));
  OR2 U1224 ( .A(n1277), .B(n1278), .Z(n1276));
  AN2 U1225 ( .A(n949), .B(n716), .Z(n1278));
  AN2 U1226 ( .A(n950), .B(n1066), .Z(n1277));
  IV2 U1227 ( .A(n723), .Z(n1066));
  OR2 U1228 ( .A(n1279), .B(n1280), .Z(n1275));
  OR2 U1229 ( .A(n1281), .B(n1282), .Z(n1280));
  AN2 U1230 ( .A(n1283), .B(n1017), .Z(n1282));
  OR2 U1231 ( .A(n1284), .B(n957), .Z(n1283));
  AN2 U1232 ( .A(n1285), .B(n784), .Z(n1284));
  AN2 U1233 ( .A(pi05), .B(n1286), .Z(n1285));
  AN2 U1234 ( .A(n725), .B(n1287), .Z(n1281));
  OR2 U1235 ( .A(n1288), .B(n1140), .Z(n1287));
  AN2 U1236 ( .A(n965), .B(n1151), .Z(n1288));
  AN2 U1237 ( .A(n744), .B(n902), .Z(n965));
  AN2 U1238 ( .A(pi01), .B(pi05), .Z(n725));
  AN2 U1239 ( .A(pi13), .B(n1289), .Z(n1279));
  OR2 U1240 ( .A(n1290), .B(n1291), .Z(n1289));
  AN2 U1241 ( .A(n971), .B(pi00), .Z(n1291));
  AN2 U1242 ( .A(n892), .B(n1292), .Z(n971));
  AN2 U1243 ( .A(pi10), .B(pi11), .Z(n1292));
  AN2 U1244 ( .A(n1293), .B(n973), .Z(n1290));
  AN2 U1245 ( .A(n1294), .B(n1295), .Z(n1293));
  OR2 U1246 ( .A(n723), .B(n1286), .Z(n1295));
  IV2 U1247 ( .A(n1151), .Z(n1286));
  OR2 U1248 ( .A(n1151), .B(n1296), .Z(n1294));
  AN2 U1249 ( .A(pi01), .B(n716), .Z(n1296));
  AN2 U1250 ( .A(n944), .B(n723), .Z(n1272));
  AN2 U1251 ( .A(n1017), .B(n716), .Z(n723));
  IV2 U1252 ( .A(pi05), .Z(n716));
  IV2 U1253 ( .A(pi01), .Z(n1017));
  AN2 U1254 ( .A(n983), .B(pi01), .Z(n1268));
  AN2 U1255 ( .A(pi11), .B(n1297), .Z(n983));
  OR2 U1256 ( .A(n1298), .B(n1299), .Z(po0));
  OR2 U1257 ( .A(n1300), .B(n1301), .Z(n1299));
  OR2 U1258 ( .A(n1302), .B(n1303), .Z(n1301));
  OR2 U1259 ( .A(n1304), .B(n1305), .Z(n1303));
  AN2 U1260 ( .A(n793), .B(n1247), .Z(n1305));
  AN2 U1261 ( .A(n924), .B(n1306), .Z(n793));
  IV2 U1262 ( .A(n1307), .Z(n1306));
  OR2 U1263 ( .A(n854), .B(n1308), .Z(n1307));
  AN2 U1264 ( .A(pi08), .B(n1063), .Z(n1308));
  IV2 U1265 ( .A(n1309), .Z(n1063));
  AN2 U1266 ( .A(n794), .B(n1041), .Z(n1304));
  AN2 U1267 ( .A(n1310), .B(n924), .Z(n794));
  OR2 U1268 ( .A(pi11), .B(n854), .Z(n1310));
  AN2 U1269 ( .A(pi11), .B(n1311), .Z(n1302));
  OR2 U1270 ( .A(n1312), .B(n1313), .Z(n1311));
  OR2 U1271 ( .A(n1314), .B(n1315), .Z(n1313));
  AN2 U1272 ( .A(n924), .B(n1316), .Z(n1315));
  AN2 U1273 ( .A(n1317), .B(n761), .Z(n1314));
  AN2 U1274 ( .A(n1023), .B(n908), .Z(n761));
  AN2 U1275 ( .A(n1151), .B(n804), .Z(n1317));
  AN2 U1276 ( .A(n1297), .B(pi00), .Z(n1312));
  AN2 U1277 ( .A(n804), .B(n1318), .Z(n1297));
  OR2 U1278 ( .A(pi10), .B(n892), .Z(n1318));
  OR2 U1279 ( .A(n1319), .B(n1320), .Z(n1300));
  AN2 U1280 ( .A(n1321), .B(n709), .Z(n1320));
  AN2 U1281 ( .A(n927), .B(n924), .Z(n1321));
  AN2 U1282 ( .A(pi04), .B(n1322), .Z(n1319));
  OR2 U1283 ( .A(n1323), .B(n930), .Z(n1322));
  AN2 U1284 ( .A(n939), .B(n1324), .Z(n930));
  AN2 U1285 ( .A(n744), .B(pi11), .Z(n1324));
  AN2 U1286 ( .A(n957), .B(n1041), .Z(n1323));
  OR2 U1287 ( .A(n1325), .B(n1326), .Z(n1298));
  OR2 U1288 ( .A(n937), .B(n1327), .Z(n1326));
  AN2 U1289 ( .A(pi13), .B(n1328), .Z(n1327));
  OR2 U1290 ( .A(n1329), .B(n1330), .Z(n1328));
  AN2 U1291 ( .A(n1109), .B(n1166), .Z(n1330));
  IV2 U1292 ( .A(pi12), .Z(n1166));
  IV2 U1293 ( .A(n1165), .Z(n1109));
  AN2 U1294 ( .A(pi12), .B(n1165), .Z(n1329));
  OR2 U1295 ( .A(n1331), .B(n1332), .Z(n1165));
  AN2 U1296 ( .A(pi13), .B(n1333), .Z(n1332));
  OR2 U1297 ( .A(n1334), .B(n1335), .Z(n1333));
  OR2 U1298 ( .A(n1336), .B(n1337), .Z(n1335));
  AN2 U1299 ( .A(n1247), .B(n1257), .Z(n1337));
  OR2 U1300 ( .A(n1338), .B(n780), .Z(n1257));
  AN2 U1301 ( .A(n1023), .B(n751), .Z(n780));
  AN2 U1302 ( .A(n944), .B(pi09), .Z(n1338));
  AN2 U1303 ( .A(pi11), .B(n1339), .Z(n1336));
  OR2 U1304 ( .A(n1340), .B(n1341), .Z(n1339));
  OR2 U1305 ( .A(n1342), .B(n1343), .Z(n1341));
  AN2 U1306 ( .A(n1344), .B(pi00), .Z(n1343));
  AN2 U1307 ( .A(n1345), .B(n1247), .Z(n1344));
  AN2 U1308 ( .A(pi10), .B(n1346), .Z(n1345));
  AN2 U1309 ( .A(n1041), .B(n713), .Z(n1342));
  IV2 U1310 ( .A(n1217), .Z(n1340));
  OR2 U1311 ( .A(pi00), .B(n817), .Z(n1217));
  OR2 U1312 ( .A(n1023), .B(n1346), .Z(n817));
  OR2 U1313 ( .A(n1347), .B(n1348), .Z(n1334));
  OR2 U1314 ( .A(n1349), .B(n1350), .Z(n1348));
  AN2 U1315 ( .A(n1316), .B(n1023), .Z(n1350));
  AN2 U1316 ( .A(n854), .B(n1351), .Z(n1349));
  OR2 U1317 ( .A(n1352), .B(n1353), .Z(n1351));
  AN2 U1318 ( .A(pi00), .B(n738), .Z(n1353));
  AN2 U1319 ( .A(pi09), .B(n1041), .Z(n1352));
  AN2 U1320 ( .A(n1248), .B(n1354), .Z(n1347));
  OR2 U1321 ( .A(n1355), .B(n1356), .Z(n1354));
  OR2 U1322 ( .A(n1357), .B(n1358), .Z(n1356));
  AN2 U1323 ( .A(n1185), .B(n1041), .Z(n1358));
  IV2 U1324 ( .A(n1092), .Z(n1185));
  AN2 U1325 ( .A(n1247), .B(n1092), .Z(n1357));
  OR2 U1326 ( .A(n1359), .B(n1360), .Z(n1092));
  AN2 U1327 ( .A(n868), .B(n718), .Z(n1360));
  AN2 U1328 ( .A(n1023), .B(n901), .Z(n868));
  AN2 U1329 ( .A(n973), .B(pi11), .Z(n901));
  AN2 U1330 ( .A(n869), .B(n1013), .Z(n1359));
  AN2 U1331 ( .A(n1361), .B(n927), .Z(n869));
  AN2 U1332 ( .A(n963), .B(pi08), .Z(n927));
  IV2 U1333 ( .A(n1041), .Z(n1247));
  AN2 U1334 ( .A(n1175), .B(n713), .Z(n1355));
  IV2 U1335 ( .A(n1013), .Z(n1175));
  AN2 U1336 ( .A(n1361), .B(n738), .Z(n1248));
  AN2 U1337 ( .A(n1362), .B(n751), .Z(n1331));
  AN2 U1338 ( .A(n902), .B(n1013), .Z(n1362));
  OR2 U1339 ( .A(n1363), .B(n1364), .Z(n1013));
  IV2 U1340 ( .A(n902), .Z(n1364));
  AN2 U1341 ( .A(n1365), .B(n1366), .Z(n1363));
  OR2 U1342 ( .A(n1188), .B(n857), .Z(n1366));
  IV2 U1343 ( .A(n908), .Z(n857));
  IV2 U1344 ( .A(n718), .Z(n1188));
  AN2 U1345 ( .A(n1367), .B(n1368), .Z(n1365));
  OR2 U1346 ( .A(n1346), .B(n1205), .Z(n1368));
  IV2 U1347 ( .A(n1074), .Z(n1205));
  IV2 U1348 ( .A(n751), .Z(n1346));
  OR2 U1349 ( .A(n829), .B(n1041), .Z(n1367));
  IV2 U1350 ( .A(n892), .Z(n829));
  AN2 U1351 ( .A(n1309), .B(n1369), .Z(n937));
  AN2 U1352 ( .A(pi13), .B(n751), .Z(n1369));
  AN2 U1353 ( .A(n939), .B(n1370), .Z(n1325));
  OR2 U1354 ( .A(n1371), .B(n1372), .Z(n1370));
  OR2 U1355 ( .A(n1074), .B(n1373), .Z(n1372));
  AN2 U1356 ( .A(n1374), .B(n944), .Z(n1373));
  AN2 U1357 ( .A(n713), .B(n709), .Z(n1374));
  AN2 U1358 ( .A(n1041), .B(pi00), .Z(n1074));
  OR2 U1359 ( .A(n1375), .B(n1376), .Z(n1041));
  OR2 U1360 ( .A(n1377), .B(n1378), .Z(n1376));
  OR2 U1361 ( .A(n1379), .B(n1380), .Z(n1378));
  AN2 U1362 ( .A(n949), .B(n709), .Z(n1380));
  OR2 U1363 ( .A(n1381), .B(n1382), .Z(n949));
  OR2 U1364 ( .A(n1383), .B(n1384), .Z(n1382));
  AN2 U1365 ( .A(n751), .B(n963), .Z(n1384));
  AN2 U1366 ( .A(n1385), .B(n860), .Z(n1383));
  IV2 U1367 ( .A(n963), .Z(n860));
  AN2 U1368 ( .A(n1386), .B(n924), .Z(n1381));
  AN2 U1369 ( .A(n804), .B(n1361), .Z(n924));
  AN2 U1370 ( .A(pi08), .B(pi10), .Z(n1386));
  AN2 U1371 ( .A(n718), .B(n1140), .Z(n1379));
  OR2 U1372 ( .A(n1387), .B(n981), .Z(n1140));
  AN2 U1373 ( .A(pi11), .B(n1388), .Z(n981));
  AN2 U1374 ( .A(n1023), .B(n1389), .Z(n1388));
  OR2 U1375 ( .A(n751), .B(n892), .Z(n1389));
  AN2 U1376 ( .A(n744), .B(n1361), .Z(n892));
  AN2 U1377 ( .A(pi09), .B(pi08), .Z(n751));
  AN2 U1378 ( .A(n944), .B(n1361), .Z(n1387));
  AN2 U1379 ( .A(n744), .B(n963), .Z(n944));
  AN2 U1380 ( .A(n784), .B(n1151), .Z(n1377));
  AN2 U1381 ( .A(n713), .B(pi04), .Z(n1151));
  AN2 U1382 ( .A(n973), .B(n902), .Z(n784));
  AN2 U1383 ( .A(n963), .B(pi13), .Z(n902));
  AN2 U1384 ( .A(n738), .B(pi10), .Z(n963));
  OR2 U1385 ( .A(n1390), .B(n1391), .Z(n1375));
  OR2 U1386 ( .A(n1392), .B(n1393), .Z(n1391));
  AN2 U1387 ( .A(n950), .B(n1394), .Z(n1393));
  OR2 U1388 ( .A(pi00), .B(pi04), .Z(n1394));
  AN2 U1389 ( .A(n1395), .B(n908), .Z(n950));
  AN2 U1390 ( .A(n1361), .B(pi08), .Z(n908));
  IV2 U1391 ( .A(pi09), .Z(n1361));
  OR2 U1392 ( .A(pi13), .B(n1309), .Z(n1395));
  AN2 U1393 ( .A(n1023), .B(n738), .Z(n1309));
  IV2 U1394 ( .A(pi11), .Z(n738));
  AN2 U1395 ( .A(n1385), .B(n1316), .Z(n1392));
  AN2 U1396 ( .A(n709), .B(pi00), .Z(n1316));
  IV2 U1397 ( .A(pi04), .Z(n709));
  AN2 U1398 ( .A(n973), .B(pi13), .Z(n1385));
  AN2 U1399 ( .A(n744), .B(pi09), .Z(n973));
  AN2 U1400 ( .A(n957), .B(n713), .Z(n1390));
  IV2 U1401 ( .A(pi00), .Z(n713));
  AN2 U1402 ( .A(n804), .B(n854), .Z(n957));
  AN2 U1403 ( .A(n744), .B(n1023), .Z(n854));
  IV2 U1404 ( .A(pi10), .Z(n1023));
  AN2 U1405 ( .A(n718), .B(n982), .Z(n1371));
  OR2 U1406 ( .A(n1396), .B(pi11), .Z(n982));
  AN2 U1407 ( .A(pi10), .B(n744), .Z(n1396));
  IV2 U1408 ( .A(pi08), .Z(n744));
  AN2 U1409 ( .A(pi00), .B(pi04), .Z(n718));
  AN2 U1410 ( .A(n804), .B(pi09), .Z(n939));
  IV2 U1411 ( .A(pi13), .Z(n804));

endmodule

module IV2(A,  Z);
  input A;
  output Z;

  assign Z = ~A;
endmodule

module AN2(A,  B,  Z);
  input A,  B;
  output Z;

  assign Z = A & B;
endmodule

module OR2(A,  B,  Z);
  input A,  B;
  output Z;

  assign Z = A | B;
endmodule
