module a #(p = 0)
();
endmodule

