module top( 1_n1 , 1_n8 , 1_n9 , 1_n21 , 1_n24 , 1_n32 , 1_n54 , 1_n61 , 1_n64 , 1_n67 , 1_n69 , 1_n76 , 1_n83 , 1_n84 , 1_n96 , 1_n97 , 1_n107 , 1_n110 , 1_n117 , 1_n120 , 1_n128 , 1_n135 , 1_n137 , 1_n142 , 1_n145 , 1_n147 , 1_n150 , 1_n154 , 1_n167 , 1_n170 , 1_n172 , 1_n182 , 1_n184 , 1_n190 , 1_n198 , 1_n204 , 1_n209 , 1_n210 , 1_n220 , 1_n222 , 1_n230 , 1_n231 , 1_n232 , 1_n233 , 1_n240 , 1_n253 , 1_n265 , 1_n268 , 1_n269 , 1_n283 , 1_n289 , 1_n290 , 1_n291 , 1_n292 , 1_n293 , 1_n296 , 1_n313 , 1_n324 , 1_n325 , 1_n330 , 1_n336 , 1_n342 , 1_n347 , 1_n350 , 1_n356 , 1_n362 , 1_n363 , 1_n364 , 1_n365 , 1_n368 , 1_n373 , 1_n383 , 1_n386 , 1_n388 , 1_n403 , 1_n415 , 1_n418 , 1_n421 , 1_n427 , 1_n432 , 1_n434 , 1_n468 , 1_n476 , 1_n478 , 1_n480 , 1_n481 , 1_n489 , 1_n490 , 1_n506 , 1_n507 , 1_n514 , 1_n524 , 1_n526 , 1_n532 , 1_n543 , 1_n565 , 1_n574 , 1_n576 , 1_n579 , 1_n588 , 1_n596 , 1_n598 , 1_n605 , 1_n608 , 1_n614 , 1_n615 , 1_n618 , 1_n623 , 1_n629 , 1_n633 , 1_n635 , 1_n640 , 1_n646 , 1_n654 , 1_n656 , 1_n663 , 1_n664 , 1_n675 , 1_n676 , 1_n677 , 1_n678 , 1_n691 , 1_n693 , 1_n704 , 1_n710 , 1_n716 , 1_n717 , 1_n722 , 1_n726 , 1_n727 , 1_n737 , 1_n740 , 1_n750 , 1_n751 , 1_n765 , 1_n769 , 1_n785 , 1_n786 , 1_n790 , 1_n793 , 1_n794 , 1_n797 , 1_n800 , 1_n814 , 1_n818 , 1_n821 , 1_n824 , 1_n829 , 1_n835 , 1_n836 , 1_n837 , 1_n840 , 1_n842 , 1_n845 , 1_n848 , 1_n851 , 1_n857 , 1_n859 , 1_n869 , 1_n877 , 1_n887 , 1_n894 , 1_n901 , 1_n909 , 1_n923 , 1_n928 , 1_n933 , 1_n934 , 1_n938 , 1_n950 , 1_n956 , 1_n964 , 1_n973 , 1_n974 , 1_n989 , 1_n990 , 1_n1013 , 1_n1014 , 1_n1019 , 1_n1021 , 1_n1023 , 1_n1025 , 1_n1026 , 1_n1030 , 1_n1032 , 1_n1036 , 1_n1039 , 1_n1042 , 1_n1043 , 1_n1049 , 1_n1052 , 1_n1058 , 1_n1065 , 1_n1070 , 1_n1091 , 1_n1093 , 1_n1098 , 1_n1099 , 1_n1108 , 1_n1117 , 1_n1121 , 1_n1122 , 1_n1131 , 1_n1134 , 1_n1138 , 1_n1143 , 1_n1146 , 1_n1150 , 1_n1151 , 1_n1157 , 1_n1160 , 1_n1161 , 1_n1162 , 1_n1165 , 1_n1170 , 1_n1177 , 1_n1184 , 1_n1187 , 1_n1189 , 1_n1192 , 1_n1194 , 1_n1198 , 1_n1223 , 1_n1239 , 1_n1240 , 1_n1243 , 1_n1251 , 1_n1253 , 1_n1255 , 1_n1275 , 1_n1276 , 1_n1280 , 1_n1303 , 1_n1310 , 1_n1311 , 1_n1314 , 1_n1331 , 1_n1335 , 1_n1339 , 1_n1361 , 1_n1366 , 1_n1373 , 1_n1375 , 1_n1378 , 1_n1389 , 1_n1392 , 1_n1396 , 1_n1398 , 1_n1407 , 1_n1409 , 1_n1411 , 1_n1412 , 1_n1413 , 1_n1418 , 1_n1422 , 1_n1425 , 1_n1438 , 1_n1442 , 1_n1454 , 1_n1474 , 1_n1475 , 1_n1478 , 1_n1479 , 1_n1485 , 1_n1508 , 1_n1511 , 1_n1512 , 1_n1515 , 1_n1518 , 1_n1530 , 1_n1531 , 1_n1542 , 1_n1545 , 1_n1547 , 1_n1549 , 1_n1551 , 1_n1552 , 1_n1555 , 1_n1556 , 1_n1562 , 1_n1574 , 1_n1575 , 1_n1580 , 1_n1581 , 1_n1589 , 1_n1594 , 1_n1596 , 1_n1601 , 1_n1604 , 1_n1606 , 1_n1620 , 1_n1628 , 1_n1629 , 1_n1630 , 1_n1631 , 1_n1645 , 1_n1648 , 1_n1655 , 1_n1665 , 1_n1671 , 1_n1676 );
    input 1_n1 , 1_n9 , 1_n67 , 1_n69 , 1_n84 , 1_n96 , 1_n107 , 1_n120 , 1_n128 , 1_n135 , 1_n137 , 1_n145 , 1_n147 , 1_n182 , 1_n184 , 1_n198 , 1_n209 , 1_n220 , 1_n222 , 1_n230 , 1_n233 , 1_n268 , 1_n283 , 1_n289 , 1_n290 , 1_n293 , 1_n296 , 1_n325 , 1_n330 , 1_n342 , 1_n356 , 1_n362 , 1_n365 , 1_n373 , 1_n386 , 1_n403 , 1_n415 , 1_n418 , 1_n421 , 1_n432 , 1_n468 , 1_n478 , 1_n481 , 1_n490 , 1_n507 , 1_n514 , 1_n526 , 1_n532 , 1_n574 , 1_n576 , 1_n579 , 1_n588 , 1_n596 , 1_n605 , 1_n615 , 1_n629 , 1_n635 , 1_n646 , 1_n654 , 1_n664 , 1_n677 , 1_n704 , 1_n710 , 1_n716 , 1_n726 , 1_n727 , 1_n737 , 1_n750 , 1_n751 , 1_n765 , 1_n769 , 1_n793 , 1_n794 , 1_n797 , 1_n818 , 1_n824 , 1_n829 , 1_n835 , 1_n837 , 1_n842 , 1_n848 , 1_n851 , 1_n857 , 1_n859 , 1_n869 , 1_n877 , 1_n901 , 1_n909 , 1_n923 , 1_n933 , 1_n934 , 1_n938 , 1_n950 , 1_n956 , 1_n973 , 1_n974 , 1_n989 , 1_n990 , 1_n1013 , 1_n1014 , 1_n1025 , 1_n1030 , 1_n1042 , 1_n1049 , 1_n1052 , 1_n1058 , 1_n1065 , 1_n1070 , 1_n1091 , 1_n1093 , 1_n1098 , 1_n1099 , 1_n1108 , 1_n1121 , 1_n1131 , 1_n1134 , 1_n1143 , 1_n1146 , 1_n1150 , 1_n1161 , 1_n1162 , 1_n1165 , 1_n1170 , 1_n1184 , 1_n1187 , 1_n1189 , 1_n1223 , 1_n1240 , 1_n1243 , 1_n1251 , 1_n1253 , 1_n1255 , 1_n1276 , 1_n1280 , 1_n1303 , 1_n1310 , 1_n1311 , 1_n1331 , 1_n1335 , 1_n1339 , 1_n1361 , 1_n1366 , 1_n1373 , 1_n1378 , 1_n1389 , 1_n1396 , 1_n1398 , 1_n1407 , 1_n1409 , 1_n1412 , 1_n1413 , 1_n1418 , 1_n1422 , 1_n1425 , 1_n1438 , 1_n1475 , 1_n1479 , 1_n1485 , 1_n1508 , 1_n1511 , 1_n1515 , 1_n1518 , 1_n1530 , 1_n1545 , 1_n1549 , 1_n1551 , 1_n1555 , 1_n1562 , 1_n1575 , 1_n1580 , 1_n1581 , 1_n1596 , 1_n1606 , 1_n1620 , 1_n1630 , 1_n1648 , 1_n1655 , 1_n1676 ;
    output 1_n8 , 1_n21 , 1_n24 , 1_n32 , 1_n54 , 1_n61 , 1_n64 , 1_n76 , 1_n83 , 1_n97 , 1_n110 , 1_n117 , 1_n142 , 1_n150 , 1_n154 , 1_n167 , 1_n170 , 1_n172 , 1_n190 , 1_n204 , 1_n210 , 1_n231 , 1_n232 , 1_n240 , 1_n253 , 1_n265 , 1_n269 , 1_n291 , 1_n292 , 1_n313 , 1_n324 , 1_n336 , 1_n347 , 1_n350 , 1_n363 , 1_n364 , 1_n368 , 1_n383 , 1_n388 , 1_n427 , 1_n434 , 1_n476 , 1_n480 , 1_n489 , 1_n506 , 1_n524 , 1_n543 , 1_n565 , 1_n598 , 1_n608 , 1_n614 , 1_n618 , 1_n623 , 1_n633 , 1_n640 , 1_n656 , 1_n663 , 1_n675 , 1_n676 , 1_n678 , 1_n691 , 1_n693 , 1_n717 , 1_n722 , 1_n740 , 1_n785 , 1_n786 , 1_n790 , 1_n800 , 1_n814 , 1_n821 , 1_n836 , 1_n840 , 1_n845 , 1_n887 , 1_n894 , 1_n928 , 1_n964 , 1_n1019 , 1_n1021 , 1_n1023 , 1_n1026 , 1_n1032 , 1_n1036 , 1_n1039 , 1_n1043 , 1_n1117 , 1_n1122 , 1_n1138 , 1_n1151 , 1_n1157 , 1_n1160 , 1_n1177 , 1_n1192 , 1_n1194 , 1_n1198 , 1_n1239 , 1_n1275 , 1_n1314 , 1_n1375 , 1_n1392 , 1_n1411 , 1_n1442 , 1_n1454 , 1_n1474 , 1_n1478 , 1_n1512 , 1_n1531 , 1_n1542 , 1_n1547 , 1_n1552 , 1_n1556 , 1_n1574 , 1_n1589 , 1_n1594 , 1_n1601 , 1_n1604 , 1_n1628 , 1_n1629 , 1_n1631 , 1_n1645 , 1_n1665 , 1_n1671 ;
    wire 1_n0 , 1_n2 , 1_n3 , 1_n4 , 1_n5 , 1_n6 , 1_n7 , 1_n10 , 1_n11 , 1_n12 , 1_n13 , 1_n14 , 1_n15 , 1_n16 , 1_n17 , 1_n18 , 1_n19 , 1_n20 , 1_n22 , 1_n23 , 1_n25 , 1_n26 , 1_n27 , 1_n28 , 1_n29 , 1_n30 , 1_n31 , 1_n33 , 1_n34 , 1_n35 , 1_n36 , 1_n37 , 1_n38 , 1_n39 , 1_n40 , 1_n41 , 1_n42 , 1_n43 , 1_n44 , 1_n45 , 1_n46 , 1_n47 , 1_n48 , 1_n49 , 1_n50 , 1_n51 , 1_n52 , 1_n53 , 1_n55 , 1_n56 , 1_n57 , 1_n58 , 1_n59 , 1_n60 , 1_n62 , 1_n63 , 1_n65 , 1_n66 , 1_n68 , 1_n70 , 1_n71 , 1_n72 , 1_n73 , 1_n74 , 1_n75 , 1_n77 , 1_n78 , 1_n79 , 1_n80 , 1_n81 , 1_n82 , 1_n85 , 1_n86 , 1_n87 , 1_n88 , 1_n89 , 1_n90 , 1_n91 , 1_n92 , 1_n93 , 1_n94 , 1_n95 , 1_n98 , 1_n99 , 1_n100 , 1_n101 , 1_n102 , 1_n103 , 1_n104 , 1_n105 , 1_n106 , 1_n108 , 1_n109 , 1_n111 , 1_n112 , 1_n113 , 1_n114 , 1_n115 , 1_n116 , 1_n118 , 1_n119 , 1_n121 , 1_n122 , 1_n123 , 1_n124 , 1_n125 , 1_n126 , 1_n127 , 1_n129 , 1_n130 , 1_n131 , 1_n132 , 1_n133 , 1_n134 , 1_n136 , 1_n138 , 1_n139 , 1_n140 , 1_n141 , 1_n143 , 1_n144 , 1_n146 , 1_n148 , 1_n149 , 1_n151 , 1_n152 , 1_n153 , 1_n155 , 1_n156 , 1_n157 , 1_n158 , 1_n159 , 1_n160 , 1_n161 , 1_n162 , 1_n163 , 1_n164 , 1_n165 , 1_n166 , 1_n168 , 1_n169 , 1_n171 , 1_n173 , 1_n174 , 1_n175 , 1_n176 , 1_n177 , 1_n178 , 1_n179 , 1_n180 , 1_n181 , 1_n183 , 1_n185 , 1_n186 , 1_n187 , 1_n188 , 1_n189 , 1_n191 , 1_n192 , 1_n193 , 1_n194 , 1_n195 , 1_n196 , 1_n197 , 1_n199 , 1_n200 , 1_n201 , 1_n202 , 1_n203 , 1_n205 , 1_n206 , 1_n207 , 1_n208 , 1_n211 , 1_n212 , 1_n213 , 1_n214 , 1_n215 , 1_n216 , 1_n217 , 1_n218 , 1_n219 , 1_n221 , 1_n223 , 1_n224 , 1_n225 , 1_n226 , 1_n227 , 1_n228 , 1_n229 , 1_n234 , 1_n235 , 1_n236 , 1_n237 , 1_n238 , 1_n239 , 1_n241 , 1_n242 , 1_n243 , 1_n244 , 1_n245 , 1_n246 , 1_n247 , 1_n248 , 1_n249 , 1_n250 , 1_n251 , 1_n252 , 1_n254 , 1_n255 , 1_n256 , 1_n257 , 1_n258 , 1_n259 , 1_n260 , 1_n261 , 1_n262 , 1_n263 , 1_n264 , 1_n266 , 1_n267 , 1_n270 , 1_n271 , 1_n272 , 1_n273 , 1_n274 , 1_n275 , 1_n276 , 1_n277 , 1_n278 , 1_n279 , 1_n280 , 1_n281 , 1_n282 , 1_n284 , 1_n285 , 1_n286 , 1_n287 , 1_n288 , 1_n294 , 1_n295 , 1_n297 , 1_n298 , 1_n299 , 1_n300 , 1_n301 , 1_n302 , 1_n303 , 1_n304 , 1_n305 , 1_n306 , 1_n307 , 1_n308 , 1_n309 , 1_n310 , 1_n311 , 1_n312 , 1_n314 , 1_n315 , 1_n316 , 1_n317 , 1_n318 , 1_n319 , 1_n320 , 1_n321 , 1_n322 , 1_n323 , 1_n326 , 1_n327 , 1_n328 , 1_n329 , 1_n331 , 1_n332 , 1_n333 , 1_n334 , 1_n335 , 1_n337 , 1_n338 , 1_n339 , 1_n340 , 1_n341 , 1_n343 , 1_n344 , 1_n345 , 1_n346 , 1_n348 , 1_n349 , 1_n351 , 1_n352 , 1_n353 , 1_n354 , 1_n355 , 1_n357 , 1_n358 , 1_n359 , 1_n360 , 1_n361 , 1_n366 , 1_n367 , 1_n369 , 1_n370 , 1_n371 , 1_n372 , 1_n374 , 1_n375 , 1_n376 , 1_n377 , 1_n378 , 1_n379 , 1_n380 , 1_n381 , 1_n382 , 1_n384 , 1_n385 , 1_n387 , 1_n389 , 1_n390 , 1_n391 , 1_n392 , 1_n393 , 1_n394 , 1_n395 , 1_n396 , 1_n397 , 1_n398 , 1_n399 , 1_n400 , 1_n401 , 1_n402 , 1_n404 , 1_n405 , 1_n406 , 1_n407 , 1_n408 , 1_n409 , 1_n410 , 1_n411 , 1_n412 , 1_n413 , 1_n414 , 1_n416 , 1_n417 , 1_n419 , 1_n420 , 1_n422 , 1_n423 , 1_n424 , 1_n425 , 1_n426 , 1_n428 , 1_n429 , 1_n430 , 1_n431 , 1_n433 , 1_n435 , 1_n436 , 1_n437 , 1_n438 , 1_n439 , 1_n440 , 1_n441 , 1_n442 , 1_n443 , 1_n444 , 1_n445 , 1_n446 , 1_n447 , 1_n448 , 1_n449 , 1_n450 , 1_n451 , 1_n452 , 1_n453 , 1_n454 , 1_n455 , 1_n456 , 1_n457 , 1_n458 , 1_n459 , 1_n460 , 1_n461 , 1_n462 , 1_n463 , 1_n464 , 1_n465 , 1_n466 , 1_n467 , 1_n469 , 1_n470 , 1_n471 , 1_n472 , 1_n473 , 1_n474 , 1_n475 , 1_n477 , 1_n479 , 1_n482 , 1_n483 , 1_n484 , 1_n485 , 1_n486 , 1_n487 , 1_n488 , 1_n491 , 1_n492 , 1_n493 , 1_n494 , 1_n495 , 1_n496 , 1_n497 , 1_n498 , 1_n499 , 1_n500 , 1_n501 , 1_n502 , 1_n503 , 1_n504 , 1_n505 , 1_n508 , 1_n509 , 1_n510 , 1_n511 , 1_n512 , 1_n513 , 1_n515 , 1_n516 , 1_n517 , 1_n518 , 1_n519 , 1_n520 , 1_n521 , 1_n522 , 1_n523 , 1_n525 , 1_n527 , 1_n528 , 1_n529 , 1_n530 , 1_n531 , 1_n533 , 1_n534 , 1_n535 , 1_n536 , 1_n537 , 1_n538 , 1_n539 , 1_n540 , 1_n541 , 1_n542 , 1_n544 , 1_n545 , 1_n546 , 1_n547 , 1_n548 , 1_n549 , 1_n550 , 1_n551 , 1_n552 , 1_n553 , 1_n554 , 1_n555 , 1_n556 , 1_n557 , 1_n558 , 1_n559 , 1_n560 , 1_n561 , 1_n562 , 1_n563 , 1_n564 , 1_n566 , 1_n567 , 1_n568 , 1_n569 , 1_n570 , 1_n571 , 1_n572 , 1_n573 , 1_n575 , 1_n577 , 1_n578 , 1_n580 , 1_n581 , 1_n582 , 1_n583 , 1_n584 , 1_n585 , 1_n586 , 1_n587 , 1_n589 , 1_n590 , 1_n591 , 1_n592 , 1_n593 , 1_n594 , 1_n595 , 1_n597 , 1_n599 , 1_n600 , 1_n601 , 1_n602 , 1_n603 , 1_n604 , 1_n606 , 1_n607 , 1_n609 , 1_n610 , 1_n611 , 1_n612 , 1_n613 , 1_n616 , 1_n617 , 1_n619 , 1_n620 , 1_n621 , 1_n622 , 1_n624 , 1_n625 , 1_n626 , 1_n627 , 1_n628 , 1_n630 , 1_n631 , 1_n632 , 1_n634 , 1_n636 , 1_n637 , 1_n638 , 1_n639 , 1_n641 , 1_n642 , 1_n643 , 1_n644 , 1_n645 , 1_n647 , 1_n648 , 1_n649 , 1_n650 , 1_n651 , 1_n652 , 1_n653 , 1_n655 , 1_n657 , 1_n658 , 1_n659 , 1_n660 , 1_n661 , 1_n662 , 1_n665 , 1_n666 , 1_n667 , 1_n668 , 1_n669 , 1_n670 , 1_n671 , 1_n672 , 1_n673 , 1_n674 , 1_n679 , 1_n680 , 1_n681 , 1_n682 , 1_n683 , 1_n684 , 1_n685 , 1_n686 , 1_n687 , 1_n688 , 1_n689 , 1_n690 , 1_n692 , 1_n694 , 1_n695 , 1_n696 , 1_n697 , 1_n698 , 1_n699 , 1_n700 , 1_n701 , 1_n702 , 1_n703 , 1_n705 , 1_n706 , 1_n707 , 1_n708 , 1_n709 , 1_n711 , 1_n712 , 1_n713 , 1_n714 , 1_n715 , 1_n718 , 1_n719 , 1_n720 , 1_n721 , 1_n723 , 1_n724 , 1_n725 , 1_n728 , 1_n729 , 1_n730 , 1_n731 , 1_n732 , 1_n733 , 1_n734 , 1_n735 , 1_n736 , 1_n738 , 1_n739 , 1_n741 , 1_n742 , 1_n743 , 1_n744 , 1_n745 , 1_n746 , 1_n747 , 1_n748 , 1_n749 , 1_n752 , 1_n753 , 1_n754 , 1_n755 , 1_n756 , 1_n757 , 1_n758 , 1_n759 , 1_n760 , 1_n761 , 1_n762 , 1_n763 , 1_n764 , 1_n766 , 1_n767 , 1_n768 , 1_n770 , 1_n771 , 1_n772 , 1_n773 , 1_n774 , 1_n775 , 1_n776 , 1_n777 , 1_n778 , 1_n779 , 1_n780 , 1_n781 , 1_n782 , 1_n783 , 1_n784 , 1_n787 , 1_n788 , 1_n789 , 1_n791 , 1_n792 , 1_n795 , 1_n796 , 1_n798 , 1_n799 , 1_n801 , 1_n802 , 1_n803 , 1_n804 , 1_n805 , 1_n806 , 1_n807 , 1_n808 , 1_n809 , 1_n810 , 1_n811 , 1_n812 , 1_n813 , 1_n815 , 1_n816 , 1_n817 , 1_n819 , 1_n820 , 1_n822 , 1_n823 , 1_n825 , 1_n826 , 1_n827 , 1_n828 , 1_n830 , 1_n831 , 1_n832 , 1_n833 , 1_n834 , 1_n838 , 1_n839 , 1_n841 , 1_n843 , 1_n844 , 1_n846 , 1_n847 , 1_n849 , 1_n850 , 1_n852 , 1_n853 , 1_n854 , 1_n855 , 1_n856 , 1_n858 , 1_n860 , 1_n861 , 1_n862 , 1_n863 , 1_n864 , 1_n865 , 1_n866 , 1_n867 , 1_n868 , 1_n870 , 1_n871 , 1_n872 , 1_n873 , 1_n874 , 1_n875 , 1_n876 , 1_n878 , 1_n879 , 1_n880 , 1_n881 , 1_n882 , 1_n883 , 1_n884 , 1_n885 , 1_n886 , 1_n888 , 1_n889 , 1_n890 , 1_n891 , 1_n892 , 1_n893 , 1_n895 , 1_n896 , 1_n897 , 1_n898 , 1_n899 , 1_n900 , 1_n902 , 1_n903 , 1_n904 , 1_n905 , 1_n906 , 1_n907 , 1_n908 , 1_n910 , 1_n911 , 1_n912 , 1_n913 , 1_n914 , 1_n915 , 1_n916 , 1_n917 , 1_n918 , 1_n919 , 1_n920 , 1_n921 , 1_n922 , 1_n924 , 1_n925 , 1_n926 , 1_n927 , 1_n929 , 1_n930 , 1_n931 , 1_n932 , 1_n935 , 1_n936 , 1_n937 , 1_n939 , 1_n940 , 1_n941 , 1_n942 , 1_n943 , 1_n944 , 1_n945 , 1_n946 , 1_n947 , 1_n948 , 1_n949 , 1_n951 , 1_n952 , 1_n953 , 1_n954 , 1_n955 , 1_n957 , 1_n958 , 1_n959 , 1_n960 , 1_n961 , 1_n962 , 1_n963 , 1_n965 , 1_n966 , 1_n967 , 1_n968 , 1_n969 , 1_n970 , 1_n971 , 1_n972 , 1_n975 , 1_n976 , 1_n977 , 1_n978 , 1_n979 , 1_n980 , 1_n981 , 1_n982 , 1_n983 , 1_n984 , 1_n985 , 1_n986 , 1_n987 , 1_n988 , 1_n991 , 1_n992 , 1_n993 , 1_n994 , 1_n995 , 1_n996 , 1_n997 , 1_n998 , 1_n999 , 1_n1000 , 1_n1001 , 1_n1002 , 1_n1003 , 1_n1004 , 1_n1005 , 1_n1006 , 1_n1007 , 1_n1008 , 1_n1009 , 1_n1010 , 1_n1011 , 1_n1012 , 1_n1015 , 1_n1016 , 1_n1017 , 1_n1018 , 1_n1020 , 1_n1022 , 1_n1024 , 1_n1027 , 1_n1028 , 1_n1029 , 1_n1031 , 1_n1033 , 1_n1034 , 1_n1035 , 1_n1037 , 1_n1038 , 1_n1040 , 1_n1041 , 1_n1044 , 1_n1045 , 1_n1046 , 1_n1047 , 1_n1048 , 1_n1050 , 1_n1051 , 1_n1053 , 1_n1054 , 1_n1055 , 1_n1056 , 1_n1057 , 1_n1059 , 1_n1060 , 1_n1061 , 1_n1062 , 1_n1063 , 1_n1064 , 1_n1066 , 1_n1067 , 1_n1068 , 1_n1069 , 1_n1071 , 1_n1072 , 1_n1073 , 1_n1074 , 1_n1075 , 1_n1076 , 1_n1077 , 1_n1078 , 1_n1079 , 1_n1080 , 1_n1081 , 1_n1082 , 1_n1083 , 1_n1084 , 1_n1085 , 1_n1086 , 1_n1087 , 1_n1088 , 1_n1089 , 1_n1090 , 1_n1092 , 1_n1094 , 1_n1095 , 1_n1096 , 1_n1097 , 1_n1100 , 1_n1101 , 1_n1102 , 1_n1103 , 1_n1104 , 1_n1105 , 1_n1106 , 1_n1107 , 1_n1109 , 1_n1110 , 1_n1111 , 1_n1112 , 1_n1113 , 1_n1114 , 1_n1115 , 1_n1116 , 1_n1118 , 1_n1119 , 1_n1120 , 1_n1123 , 1_n1124 , 1_n1125 , 1_n1126 , 1_n1127 , 1_n1128 , 1_n1129 , 1_n1130 , 1_n1132 , 1_n1133 , 1_n1135 , 1_n1136 , 1_n1137 , 1_n1139 , 1_n1140 , 1_n1141 , 1_n1142 , 1_n1144 , 1_n1145 , 1_n1147 , 1_n1148 , 1_n1149 , 1_n1152 , 1_n1153 , 1_n1154 , 1_n1155 , 1_n1156 , 1_n1158 , 1_n1159 , 1_n1163 , 1_n1164 , 1_n1166 , 1_n1167 , 1_n1168 , 1_n1169 , 1_n1171 , 1_n1172 , 1_n1173 , 1_n1174 , 1_n1175 , 1_n1176 , 1_n1178 , 1_n1179 , 1_n1180 , 1_n1181 , 1_n1182 , 1_n1183 , 1_n1185 , 1_n1186 , 1_n1188 , 1_n1190 , 1_n1191 , 1_n1193 , 1_n1195 , 1_n1196 , 1_n1197 , 1_n1199 , 1_n1200 , 1_n1201 , 1_n1202 , 1_n1203 , 1_n1204 , 1_n1205 , 1_n1206 , 1_n1207 , 1_n1208 , 1_n1209 , 1_n1210 , 1_n1211 , 1_n1212 , 1_n1213 , 1_n1214 , 1_n1215 , 1_n1216 , 1_n1217 , 1_n1218 , 1_n1219 , 1_n1220 , 1_n1221 , 1_n1222 , 1_n1224 , 1_n1225 , 1_n1226 , 1_n1227 , 1_n1228 , 1_n1229 , 1_n1230 , 1_n1231 , 1_n1232 , 1_n1233 , 1_n1234 , 1_n1235 , 1_n1236 , 1_n1237 , 1_n1238 , 1_n1241 , 1_n1242 , 1_n1244 , 1_n1245 , 1_n1246 , 1_n1247 , 1_n1248 , 1_n1249 , 1_n1250 , 1_n1252 , 1_n1254 , 1_n1256 , 1_n1257 , 1_n1258 , 1_n1259 , 1_n1260 , 1_n1261 , 1_n1262 , 1_n1263 , 1_n1264 , 1_n1265 , 1_n1266 , 1_n1267 , 1_n1268 , 1_n1269 , 1_n1270 , 1_n1271 , 1_n1272 , 1_n1273 , 1_n1274 , 1_n1277 , 1_n1278 , 1_n1279 , 1_n1281 , 1_n1282 , 1_n1283 , 1_n1284 , 1_n1285 , 1_n1286 , 1_n1287 , 1_n1288 , 1_n1289 , 1_n1290 , 1_n1291 , 1_n1292 , 1_n1293 , 1_n1294 , 1_n1295 , 1_n1296 , 1_n1297 , 1_n1298 , 1_n1299 , 1_n1300 , 1_n1301 , 1_n1302 , 1_n1304 , 1_n1305 , 1_n1306 , 1_n1307 , 1_n1308 , 1_n1309 , 1_n1312 , 1_n1313 , 1_n1315 , 1_n1316 , 1_n1317 , 1_n1318 , 1_n1319 , 1_n1320 , 1_n1321 , 1_n1322 , 1_n1323 , 1_n1324 , 1_n1325 , 1_n1326 , 1_n1327 , 1_n1328 , 1_n1329 , 1_n1330 , 1_n1332 , 1_n1333 , 1_n1334 , 1_n1336 , 1_n1337 , 1_n1338 , 1_n1340 , 1_n1341 , 1_n1342 , 1_n1343 , 1_n1344 , 1_n1345 , 1_n1346 , 1_n1347 , 1_n1348 , 1_n1349 , 1_n1350 , 1_n1351 , 1_n1352 , 1_n1353 , 1_n1354 , 1_n1355 , 1_n1356 , 1_n1357 , 1_n1358 , 1_n1359 , 1_n1360 , 1_n1362 , 1_n1363 , 1_n1364 , 1_n1365 , 1_n1367 , 1_n1368 , 1_n1369 , 1_n1370 , 1_n1371 , 1_n1372 , 1_n1374 , 1_n1376 , 1_n1377 , 1_n1379 , 1_n1380 , 1_n1381 , 1_n1382 , 1_n1383 , 1_n1384 , 1_n1385 , 1_n1386 , 1_n1387 , 1_n1388 , 1_n1390 , 1_n1391 , 1_n1393 , 1_n1394 , 1_n1395 , 1_n1397 , 1_n1399 , 1_n1400 , 1_n1401 , 1_n1402 , 1_n1403 , 1_n1404 , 1_n1405 , 1_n1406 , 1_n1408 , 1_n1410 , 1_n1414 , 1_n1415 , 1_n1416 , 1_n1417 , 1_n1419 , 1_n1420 , 1_n1421 , 1_n1423 , 1_n1424 , 1_n1426 , 1_n1427 , 1_n1428 , 1_n1429 , 1_n1430 , 1_n1431 , 1_n1432 , 1_n1433 , 1_n1434 , 1_n1435 , 1_n1436 , 1_n1437 , 1_n1439 , 1_n1440 , 1_n1441 , 1_n1443 , 1_n1444 , 1_n1445 , 1_n1446 , 1_n1447 , 1_n1448 , 1_n1449 , 1_n1450 , 1_n1451 , 1_n1452 , 1_n1453 , 1_n1455 , 1_n1456 , 1_n1457 , 1_n1458 , 1_n1459 , 1_n1460 , 1_n1461 , 1_n1462 , 1_n1463 , 1_n1464 , 1_n1465 , 1_n1466 , 1_n1467 , 1_n1468 , 1_n1469 , 1_n1470 , 1_n1471 , 1_n1472 , 1_n1473 , 1_n1476 , 1_n1477 , 1_n1480 , 1_n1481 , 1_n1482 , 1_n1483 , 1_n1484 , 1_n1486 , 1_n1487 , 1_n1488 , 1_n1489 , 1_n1490 , 1_n1491 , 1_n1492 , 1_n1493 , 1_n1494 , 1_n1495 , 1_n1496 , 1_n1497 , 1_n1498 , 1_n1499 , 1_n1500 , 1_n1501 , 1_n1502 , 1_n1503 , 1_n1504 , 1_n1505 , 1_n1506 , 1_n1507 , 1_n1509 , 1_n1510 , 1_n1513 , 1_n1514 , 1_n1516 , 1_n1517 , 1_n1519 , 1_n1520 , 1_n1521 , 1_n1522 , 1_n1523 , 1_n1524 , 1_n1525 , 1_n1526 , 1_n1527 , 1_n1528 , 1_n1529 , 1_n1532 , 1_n1533 , 1_n1534 , 1_n1535 , 1_n1536 , 1_n1537 , 1_n1538 , 1_n1539 , 1_n1540 , 1_n1541 , 1_n1543 , 1_n1544 , 1_n1546 , 1_n1548 , 1_n1550 , 1_n1553 , 1_n1554 , 1_n1557 , 1_n1558 , 1_n1559 , 1_n1560 , 1_n1561 , 1_n1563 , 1_n1564 , 1_n1565 , 1_n1566 , 1_n1567 , 1_n1568 , 1_n1569 , 1_n1570 , 1_n1571 , 1_n1572 , 1_n1573 , 1_n1576 , 1_n1577 , 1_n1578 , 1_n1579 , 1_n1582 , 1_n1583 , 1_n1584 , 1_n1585 , 1_n1586 , 1_n1587 , 1_n1588 , 1_n1590 , 1_n1591 , 1_n1592 , 1_n1593 , 1_n1595 , 1_n1597 , 1_n1598 , 1_n1599 , 1_n1600 , 1_n1602 , 1_n1603 , 1_n1605 , 1_n1607 , 1_n1608 , 1_n1609 , 1_n1610 , 1_n1611 , 1_n1612 , 1_n1613 , 1_n1614 , 1_n1615 , 1_n1616 , 1_n1617 , 1_n1618 , 1_n1619 , 1_n1621 , 1_n1622 , 1_n1623 , 1_n1624 , 1_n1625 , 1_n1626 , 1_n1627 , 1_n1632 , 1_n1633 , 1_n1634 , 1_n1635 , 1_n1636 , 1_n1637 , 1_n1638 , 1_n1639 , 1_n1640 , 1_n1641 , 1_n1642 , 1_n1643 , 1_n1644 , 1_n1646 , 1_n1647 , 1_n1649 , 1_n1650 , 1_n1651 , 1_n1652 , 1_n1653 , 1_n1654 , 1_n1656 , 1_n1657 , 1_n1658 , 1_n1659 , 1_n1660 , 1_n1661 , 1_n1662 , 1_n1663 , 1_n1664 , 1_n1666 , 1_n1667 , 1_n1668 , 1_n1669 , 1_n1670 , 1_n1672 , 1_n1673 , 1_n1674 , 1_n1675 , 1_n1677 ;
assign 1_n806 = ~(1_n1255 | 1_n1030);
assign 1_n1163 = ~(1_n1422 | 1_n148);
assign 1_n1015 = ~(1_n1041 | 1_n967);
assign 1_n1516 = ~1_n47;
assign 1_n394 = 1_n413 | 1_n513;
assign 1_n1359 = ~(1_n198 | 1_n1053);
assign 1_n360 = ~(1_n1255 | 1_n1251);
assign 1_n1472 = ~1_n1408;
assign 1_n936 = ~1_n51;
assign 1_n1635 = ~(1_n915 ^ 1_n1554);
assign 1_n1447 = ~(1_n1127 ^ 1_n742);
assign 1_n402 = ~(1_n1255 | 1_n209);
assign 1_n1043 = 1_n1629 | 1_n1529;
assign 1_n1294 = ~(1_n605 | 1_n734);
assign 1_n1282 = 1_n1295 ^ 1_n71;
assign 1_n191 = 1_n641 | 1_n539;
assign 1_n1033 = 1_n1348 & 1_n1535;
assign 1_n667 = 1_n1491 & 1_n632;
assign 1_n518 = ~1_n1365;
assign 1_n1007 = 1_n713 | 1_n519;
assign 1_n890 = 1_n1517 | 1_n1139;
assign 1_n1491 = 1_n275 | 1_n277;
assign 1_n71 = 1_n975 & 1_n570;
assign 1_n28 = ~(1_n272 | 1_n1283);
assign 1_n1085 = 1_n944 | 1_n774;
assign 1_n524 = 1_n1629 | 1_n1089;
assign 1_n60 = ~1_n218;
assign 1_n434 = ~1_n1587;
assign 1_n151 = 1_n917 | 1_n783;
assign 1_n822 = ~(1_n1133 | 1_n931);
assign 1_n1496 = 1_n1242 ^ 1_n1265;
assign 1_n1010 = 1_n954 & 1_n938;
assign 1_n610 = 1_n1530 | 1_n245;
assign 1_n1229 = ~1_n729;
assign 1_n720 = 1_n940 | 1_n841;
assign 1_n1384 = ~1_n847;
assign 1_n1320 = ~(1_n1311 | 1_n1030);
assign 1_n1190 = ~1_n770;
assign 1_n1324 = ~1_n825;
assign 1_n79 = 1_n1495 | 1_n1446;
assign 1_n598 = 1_n425 | 1_n177;
assign 1_n1619 = ~(1_n116 ^ 1_n1669);
assign 1_n506 = 1_n1629 | 1_n323;
assign 1_n504 = ~1_n1624;
assign 1_n981 = 1_n1143 & 1_n325;
assign 1_n542 = ~(1_n402 | 1_n1027);
assign 1_n1272 = ~(1_n1274 | 1_n1518);
assign 1_n1609 = 1_n243 | 1_n28;
assign 1_n949 = ~(1_n453 ^ 1_n500);
assign 1_n985 = ~(1_n300 | 1_n1211);
assign 1_n47 = 1_n550 | 1_n320;
assign 1_n287 = 1_n559 | 1_n492;
assign 1_n206 = ~(1_n289 | 1_n62);
assign 1_n163 = ~(1_n1554 ^ 1_n1599);
assign 1_n1344 = ~(1_n10 | 1_n1478);
assign 1_n862 = ~(1_n403 | 1_n789);
assign 1_n1428 = 1_n224 & 1_n514;
assign 1_n1269 = ~1_n397;
assign 1_n427 = 1_n449 | 1_n168;
assign 1_n1593 = ~(1_n960 | 1_n654);
assign 1_n66 = ~1_n1290;
assign 1_n57 = 1_n707 & 1_n877;
assign 1_n1199 = ~1_n1356;
assign 1_n1178 = ~(1_n622 | 1_n677);
assign 1_n140 = ~1_n1378;
assign 1_n339 = ~(1_n1481 ^ 1_n662);
assign 1_n558 = ~1_n532;
assign 1_n400 = ~1_n902;
assign 1_n32 = ~(1_n1629 | 1_n1323);
assign 1_n1181 = ~1_n646;
assign 1_n1368 = 1_n1338 & 1_n1354;
assign 1_n87 = ~(1_n848 | 1_n525);
assign 1_n174 = ~1_n1435;
assign 1_n260 = ~(1_n763 ^ 1_n1058);
assign 1_n725 = 1_n922 | 1_n1420;
assign 1_n550 = ~(1_n1390 ^ 1_n147);
assign 1_n728 = ~(1_n615 | 1_n1199);
assign 1_n2 = ~1_n1108;
assign 1_n761 = ~1_n1147;
assign 1_n83 = 1_n224 & 1_n415;
assign 1_n649 = ~1_n1384;
assign 1_n1100 = 1_n737 & 1_n1243;
assign 1_n927 = ~(1_n483 | 1_n239);
assign 1_n962 = ~1_n1235;
assign 1_n1219 = 1_n584 | 1_n81;
assign 1_n45 = ~(1_n135 | 1_n385);
assign 1_n286 = ~(1_n464 | 1_n248);
assign 1_n746 = ~(1_n121 ^ 1_n600);
assign 1_n540 = 1_n929 & 1_n1339;
assign 1_n41 = 1_n102 | 1_n404;
assign 1_n185 = 1_n242 | 1_n371;
assign 1_n471 = ~(1_n1676 | 1_n1195);
assign 1_n1454 = ~(1_n1099 | 1_n1499);
assign 1_n227 = ~1_n1193;
assign 1_n106 = 1_n969 & 1_n403;
assign 1_n808 = 1_n1180 | 1_n1528;
assign 1_n1647 = 1_n1268 & 1_n726;
assign 1_n895 = ~(1_n950 | 1_n644);
assign 1_n543 = 1_n1629 | 1_n890;
assign 1_n1626 = ~(1_n238 | 1_n1143);
assign 1_n72 = ~1_n956;
assign 1_n534 = 1_n658 | 1_n849;
assign 1_n370 = 1_n1302 & 1_n1379;
assign 1_n754 = ~1_n196;
assign 1_n1275 = 1_n165 | 1_n326;
assign 1_n23 = 1_n1465 & 1_n751;
assign 1_n343 = 1_n1011 & 1_n181;
assign 1_n1371 = ~(1_n527 | 1_n962);
assign 1_n644 = ~(1_n1504 | 1_n1248);
assign 1_n1211 = ~1_n1457;
assign 1_n1244 = ~1_n220;
assign 1_n1246 = ~(1_n6 | 1_n1272);
assign 1_n1258 = ~(1_n120 | 1_n930);
assign 1_n854 = 1_n331 | 1_n104;
assign 1_n517 = ~1_n121;
assign 1_n1179 = ~(1_n42 | 1_n1283);
assign 1_n1417 = 1_n839 | 1_n1371;
assign 1_n1322 = ~(1_n848 | 1_n424);
assign 1_n1060 = ~(1_n960 | 1_n859);
assign 1_n1604 = 1_n1629 | 1_n444;
assign 1_n811 = 1_n319 | 1_n1543;
assign 1_n1547 = ~1_n842;
assign 1_n964 = ~1_n1520;
assign 1_n1477 = ~1_n902;
assign 1_n25 = 1_n647 & 1_n1;
assign 1_n169 = ~(1_n256 | 1_n1645);
assign 1_n954 = 1_n1320 | 1_n1330;
assign 1_n1191 = ~(1_n1524 ^ 1_n1435);
assign 1_n1153 = ~1_n877;
assign 1_n187 = ~1_n297;
assign 1_n695 = 1_n401 & 1_n1108;
assign 1_n7 = 1_n228 | 1_n714;
assign 1_n1419 = ~1_n1038;
assign 1_n463 = ~1_n573;
assign 1_n1476 = 1_n1654 | 1_n736;
assign 1_n1316 = ~(1_n960 | 1_n646);
assign 1_n1617 = ~(1_n112 ^ 1_n125);
assign 1_n398 = ~1_n372;
assign 1_n1250 = ~(1_n561 | 1_n752);
assign 1_n815 = 1_n442 | 1_n7;
assign 1_n961 = ~(1_n454 ^ 1_n594);
assign 1_n1576 = 1_n800 & 1_n507;
assign 1_n682 = 1_n628 & 1_n184;
assign 1_n670 = ~1_n1336;
assign 1_n913 = ~(1_n1255 | 1_n1518);
assign 1_n1046 = 1_n540 | 1_n1203;
assign 1_n529 = ~(1_n1606 | 1_n1181);
assign 1_n1375 = 1_n1629 | 1_n1657;
assign 1_n1416 = 1_n1234 & 1_n93;
assign 1_n589 = 1_n564 & 1_n1378;
assign 1_n270 = ~1_n514;
assign 1_n1531 = 1_n8 | 1_n741;
assign 1_n1657 = 1_n82 | 1_n1079;
assign 1_n438 = ~1_n550;
assign 1_n254 = 1_n4 | 1_n44;
assign 1_n801 = ~1_n863;
assign 1_n1140 = ~(1_n419 ^ 1_n1634);
assign 1_n531 = 1_n135 & 1_n325;
assign 1_n495 = 1_n1046 | 1_n787;
assign 1_n1095 = 1_n943 | 1_n724;
assign 1_n1570 = 1_n1215 | 1_n864;
assign 1_n688 = 1_n1304 ^ 1_n1564;
assign 1_n333 = ~(1_n198 | 1_n72);
assign 1_n1307 = ~1_n393;
assign 1_n1443 = ~(1_n1014 | 1_n166);
assign 1_n1631 = ~1_n523;
assign 1_n1210 = 1_n295 | 1_n1185;
assign 1_n839 = 1_n1524 & 1_n1479;
assign 1_n747 = 1_n1013 & 1_n1606;
assign 1_n836 = 1_n984 | 1_n1559;
assign 1_n789 = ~(1_n772 | 1_n1376);
assign 1_n473 = 1_n1334 | 1_n169;
assign 1_n1493 = ~1_n184;
assign 1_n907 = ~(1_n694 | 1_n590);
assign 1_n880 = 1_n1364 & 1_n765;
assign 1_n1437 = 1_n68 | 1_n1659;
assign 1_n123 = 1_n1140 & 1_n632;
assign 1_n810 = ~(1_n289 | 1_n819);
assign 1_n73 = ~(1_n1410 | 1_n1404);
assign 1_n1301 = ~(1_n198 | 1_n1105);
assign 1_n618 = ~1_n797;
assign 1_n75 = ~1_n932;
assign 1_n849 = 1_n728 | 1_n465;
assign 1_n19 = ~(1_n706 | 1_n1593);
assign 1_n0 = ~1_n997;
assign 1_n1397 = 1_n433 | 1_n1399;
assign 1_n1565 = ~(1_n1367 | 1_n261);
assign 1_n1343 = 1_n1335 | 1_n162;
assign 1_n1497 = ~(1_n1042 | 1_n183);
assign 1_n1018 = ~(1_n735 | 1_n1039);
assign 1_n1076 = ~(1_n870 ^ 1_n1496);
assign 1_n607 = ~(1_n1398 | 1_n1560);
assign 1_n805 = ~(1_n256 | 1_n621);
assign 1_n1129 = ~1_n573;
assign 1_n844 = 1_n118 | 1_n698;
assign 1_n872 = ~(1_n468 | 1_n670);
assign 1_n130 = ~1_n1360;
assign 1_n24 = 1_n1629 | 1_n639;
assign 1_n952 = 1_n1124 | 1_n200;
assign 1_n65 = ~(1_n342 | 1_n757);
assign 1_n1583 = 1_n1243 & 1_n1253;
assign 1_n733 = ~(1_n1 | 1_n1632);
assign 1_n1050 = 1_n856 | 1_n100;
assign 1_n1499 = ~1_n1412;
assign 1_n208 = ~(1_n198 | 1_n1526);
assign 1_n1651 = 1_n1596 & 1_n1606;
assign 1_n1468 = ~(1_n221 | 1_n1302);
assign 1_n416 = ~1_n280;
assign 1_n1214 = 1_n874 | 1_n1449;
assign 1_n1012 = ~1_n517;
assign 1_n500 = ~(1_n620 ^ 1_n241);
assign 1_n1313 = 1_n1221 | 1_n1625;
assign 1_n1109 = ~(1_n1335 ^ 1_n629);
assign 1_n1613 = ~(1_n859 ^ 1_n677);
assign 1_n1394 = ~(1_n283 | 1_n792);
assign 1_n675 = ~1_n196;
assign 1_n515 = ~(1_n1243 | 1_n72);
assign 1_n194 = 1_n103 | 1_n322;
assign 1_n781 = ~1_n1587;
assign 1_n965 = ~(1_n933 | 1_n1156);
assign 1_n112 = ~1_n975;
assign 1_n1578 = ~1_n1405;
assign 1_n1502 = 1_n1140 | 1_n318;
assign 1_n1567 = ~(1_n615 | 1_n1022);
assign 1_n1224 = ~(1_n818 | 1_n544);
assign 1_n1257 = ~(1_n268 ^ 1_n209);
assign 1_n972 = 1_n746 & 1_n632;
assign 1_n219 = 1_n616 & 1_n765;
assign 1_n297 = 1_n747 | 1_n886;
assign 1_n216 = 1_n940 ^ 1_n1329;
assign 1_n1450 = 1_n69 & 1_n1243;
assign 1_n327 = 1_n156 & 1_n145;
assign 1_n81 = ~(1_n1227 | 1_n291);
assign 1_n387 = 1_n1346 | 1_n208;
assign 1_n1273 = ~(1_n1511 | 1_n959);
assign 1_n717 = 1_n1134;
assign 1_n1217 = 1_n579 & 1_n1243;
assign 1_n617 = 1_n956 & 1_n325;
assign 1_n1288 = ~1_n625;
assign 1_n226 = ~(1_n236 | 1_n1251);
assign 1_n930 = ~(1_n1308 ^ 1_n835);
assign 1_n1079 = 1_n1238 | 1_n5;
assign 1_n1402 = ~1_n652;
assign 1_n55 = ~1_n1251;
assign 1_n1039 = ~1_n1440;
assign 1_n846 = 1_n1094 | 1_n983;
assign 1_n911 = ~(1_n361 ^ 1_n1165);
assign 1_n121 = ~(1_n1430 ^ 1_n1389);
assign 1_n1636 = ~1_n931;
assign 1_n1466 = 1_n267 | 1_n1400;
assign 1_n1188 = ~(1_n198 | 1_n884);
assign 1_n1020 = 1_n407 & 1_n632;
assign 1_n1594 = 1_n484 | 1_n475;
assign 1_n1632 = ~(1_n1463 ^ 1_n1434);
assign 1_n1287 = ~(1_n198 | 1_n935);
assign 1_n94 = ~1_n115;
assign 1_n1107 = 1_n1319 ^ 1_n1264;
assign 1_n1399 = ~(1_n735 | 1_n964);
assign 1_n1653 = 1_n490 & 1_n325;
assign 1_n876 = ~(1_n843 | 1_n1177);
assign 1_n1369 = 1_n1413 & 1_n989;
assign 1_n454 = ~(1_n1572 ^ 1_n1591);
assign 1_n887 = ~1_n1247;
assign 1_n1629 = 1_n1090;
assign 1_n1434 = ~(1_n372 ^ 1_n613);
assign 1_n116 = ~(1_n161 ^ 1_n625);
assign 1_n401 = 1_n1600 | 1_n947;
assign 1_n304 = ~1_n982;
assign 1_n1204 = ~1_n306;
assign 1_n464 = ~(1_n1255 | 1_n135);
assign 1_n111 = ~(1_n1398 | 1_n665);
assign 1_n888 = ~(1_n1425 | 1_n999);
assign 1_n1130 = 1_n1481 | 1_n1292;
assign 1_n683 = 1_n140 | 1_n1416;
assign 1_n1154 = 1_n38 | 1_n867;
assign 1_n1483 = ~(1_n1635 ^ 1_n1298);
assign 1_n597 = 1_n149 & 1_n796;
assign 1_n50 = 1_n416 & 1_n570;
assign 1_n199 = 1_n759 | 1_n1359;
assign 1_n1505 = ~(1_n882 | 1_n1256);
assign 1_n1510 = 1_n1293 | 1_n548;
assign 1_n281 = ~(1_n367 | 1_n52);
assign 1_n165 = 1_n1000 | 1_n307;
assign 1_n1427 = ~1_n507;
assign 1_n1633 = ~(1_n1091 | 1_n665);
assign 1_n894 = 1_n1629 | 1_n472;
assign 1_n714 = 1_n1067 & 1_n1520;
assign 1_n1112 = ~(1_n897 | 1_n971);
assign 1_n1644 = 1_n1143 & 1_n230;
assign 1_n1220 = 1_n351 & 1_n869;
assign 1_n443 = ~(1_n738 ^ 1_n1002);
assign 1_n734 = ~1_n908;
assign 1_n259 = ~1_n1615;
assign 1_n486 = ~(1_n1667 | 1_n686);
assign 1_n1247 = ~1_n392;
assign 1_n232 = 1_n480;
assign 1_n702 = ~(1_n1606 | 1_n800);
assign 1_n419 = ~(1_n625 ^ 1_n403);
assign 1_n1062 = ~1_n1432;
assign 1_n580 = ~(1_n355 | 1_n556);
assign 1_n623 = 1_n455 & 1_n521;
assign 1_n320 = ~1_n493;
assign 1_n736 = 1_n1007 | 1_n1437;
assign 1_n1135 = 1_n997 & 1_n1121;
assign 1_n314 = 1_n356 & 1_n1243;
assign 1_n467 = 1_n1471 | 1_n537;
assign 1_n1618 = 1_n481 & 1_n1606;
assign 1_n447 = ~(1_n451 | 1_n316);
assign 1_n1159 = ~1_n731;
assign 1_n1507 = 1_n1492 & 1_n147;
assign 1_n703 = ~(1_n882 | 1_n394);
assign 1_n445 = 1_n176 & 1_n950;
assign 1_n1465 = ~1_n218;
assign 1_n512 = ~1_n1409;
assign 1_n560 = 1_n1331 & 1_n1243;
assign 1_n309 = ~(1_n342 | 1_n649);
assign 1_n730 = 1_n1470 & 1_n1232;
assign 1_n175 = ~(1_n304 | 1_n863);
assign 1_n698 = 1_n681 | 1_n131;
assign 1_n906 = ~(1_n1311 | 1_n135);
assign 1_n1105 = ~1_n135;
assign 1_n347 = 1_n1629 | 1_n1313;
assign 1_n282 = ~(1_n643 ^ 1_n1047);
assign 1_n631 = ~(1_n1108 | 1_n1077);
assign 1_n759 = ~(1_n1311 | 1_n646);
assign 1_n545 = ~1_n1166;
assign 1_n986 = ~(1_n272 | 1_n210);
assign 1_n834 = 1_n416 & 1_n94;
assign 1_n1061 = ~(1_n1184 | 1_n1650);
assign 1_n85 = 1_n1152 & 1_n490;
assign 1_n203 = 1_n23 | 1_n430;
assign 1_n181 = 1_n1357 | 1_n70;
assign 1_n1333 = ~1_n57;
assign 1_n1557 = ~1_n621;
assign 1_n1432 = ~1_n1173;
assign 1_n788 = ~(1_n1047 ^ 1_n1128);
assign 1_n1540 = 1_n1186 | 1_n705;
assign 1_n493 = 1_n274 & 1_n777;
assign 1_n313 = 1_n1629 | 1_n1461;
assign 1_n786 = 1_n478;
assign 1_n1340 = 1_n171 | 1_n764;
assign 1_n1083 = 1_n349 | 1_n1344;
assign 1_n484 = 1_n1607 | 1_n900;
assign 1_n861 = ~1_n1342;
assign 1_n4 = 1_n373 & 1_n1243;
assign 1_n385 = ~1_n365;
assign 1_n902 = ~1_n138;
assign 1_n882 = ~1_n1290;
assign 1_n1084 = ~(1_n1035 ^ 1_n1619);
assign 1_n99 = 1_n1264 | 1_n657;
assign 1_n828 = 1_n1289 | 1_n978;
assign 1_n275 = 1_n968 & 1_n1421;
assign 1_n1292 = ~(1_n1242 | 1_n600);
assign 1_n168 = 1_n1055 | 1_n805;
assign 1_n104 = 1_n186 | 1_n437;
assign 1_n22 = 1_n1382 & 1_n1165;
assign 1_n231 = 1_n284 | 1_n650;
assign 1_n721 = 1_n1226 | 1_n1502;
assign 1_n1654 = 1_n749 | 1_n538;
assign 1_n1215 = ~(1_n1378 | 1_n1527);
assign 1_n966 = 1_n271 | 1_n216;
assign 1_n582 = ~(1_n577 | 1_n643);
assign 1_n125 = ~1_n459;
assign 1_n511 = ~(1_n1311 | 1_n1518);
assign 1_n946 = ~(1_n1146 | 1_n130);
assign 1_n141 = ~(1_n1627 ^ 1_n376);
assign 1_n825 = ~1_n1137;
assign 1_n117 = 1_n811 | 1_n1284;
assign 1_n150 = 1_n1629 | 1_n1154;
assign 1_n706 = 1_n654 & 1_n325;
assign 1_n884 = ~1_n209;
assign 1_n1577 = 1_n375 | 1_n795;
assign 1_n638 = ~(1_n1605 | 1_n824);
assign 1_n43 = ~1_n283;
assign 1_n1185 = ~(1_n1058 | 1_n385);
assign 1_n753 = ~1_n419;
assign 1_n431 = ~(1_n264 ^ 1_n922);
assign 1_n587 = ~(1_n1637 ^ 1_n1045);
assign 1_n93 = 1_n1181 | 1_n700;
assign 1_n34 = ~1_n1436;
assign 1_n1193 = 1_n488 & 1_n1551;
assign 1_n382 = ~(1_n1621 | 1_n860);
assign 1_n1022 = ~1_n1336;
assign 1_n35 = 1_n578 | 1_n571;
assign 1_n183 = ~1_n701;
assign 1_n684 = 1_n965 | 1_n143;
assign 1_n1342 = ~1_n66;
assign 1_n29 = ~(1_n1064 | 1_n124);
assign 1_n1148 = ~1_n1170;
assign 1_n1088 = 1_n1545 & 1_n230;
assign 1_n1519 = 1_n1658 | 1_n1590;
assign 1_n444 = 1_n651 | 1_n976;
assign 1_n1525 = 1_n107 & 1_n1243;
assign 1_n396 = ~(1_n1361 | 1_n1480);
assign 1_n1347 = ~(1_n1309 | 1_n1256);
assign 1_n1453 = ~(1_n909 | 1_n1031);
assign 1_n1055 = ~(1_n1162 | 1_n1480);
assign 1_n1145 = ~(1_n1152 | 1_n1547);
assign 1_n864 = 1_n199 & 1_n1378;
assign 1_n592 = 1_n824 | 1_n385;
assign 1_n685 = 1_n647 & 1_n1555;
assign 1_n100 = 1_n1202 | 1_n555;
assign 1_n900 = ~(1_n1374 | 1_n545);
assign 1_n611 = ~1_n1647;
assign 1_n823 = ~(1_n1430 ^ 1_n361);
assign 1_n1424 = ~(1_n605 | 1_n959);
assign 1_n352 = ~1_n824;
assign 1_n255 = 1_n1494 | 1_n1048;
assign 1_n261 = ~(1_n141 ^ 1_n949);
assign 1_n1658 = 1_n1032 | 1_n523;
assign 1_n466 = ~1_n1592;
assign 1_n91 = 1_n122 & 1_n1005;
assign 1_n621 = 1_n203 | 1_n202;
assign 1_n1283 = 1_n916 | 1_n593;
assign 1_n991 = ~1_n692;
assign 1_n21 = 1_n473 | 1_n1174;
assign 1_n858 = 1_n677 & 1_n325;
assign 1_n1514 = 1_n1278 | 1_n1612;
assign 1_n516 = 1_n1472 & 1_n438;
assign 1_n768 = ~(1_n1002 | 1_n48);
assign 1_n161 = 1_n1381 & 1_n1606;
assign 1_n671 = ~1_n1335;
assign 1_n300 = ~1_n1365;
assign 1_n475 = 1_n567 | 1_n1468;
assign 1_n655 = 1_n448 | 1_n13;
assign 1_n242 = 1_n395 & 1_n1580;
assign 1_n520 = 1_n18 | 1_n1595;
assign 1_n1296 = 1_n956 & 1_n230;
assign 1_n204 = 1_n197 | 1_n712;
assign 1_n657 = 1_n1319 | 1_n854;
assign 1_n1661 = 1_n1489 | 1_n1576;
assign 1_n1356 = ~1_n611;
assign 1_n110 = 1_n1127 | 1_n59;
assign 1_n449 = 1_n745 | 1_n541;
assign 1_n921 = ~(1_n927 ^ 1_n672);
assign 1_n1436 = ~1_n26;
assign 1_n591 = 1_n995 & 1_n753;
assign 1_n739 = ~(1_n1161 | 1_n162);
assign 1_n1386 = ~(1_n1255 | 1_n956);
assign 1_n277 = 1_n577 & 1_n1016;
assign 1_n1524 = 1_n39 | 1_n515;
assign 1_n54 = 1_n1155 | 1_n699;
assign 1_n284 = 1_n1443 | 1_n382;
assign 1_n331 = 1_n1343 & 1_n1315;
assign 1_n496 = ~(1_n933 | 1_n1544);
assign 1_n748 = 1_n467 | 1_n1582;
assign 1_n672 = ~(1_n1158 | 1_n106);
assign 1_n814 = 1_n1214 | 1_n666;
assign 1_n1001 = ~1_n1173;
assign 1_n791 = ~1_n962;
assign 1_n250 = 1_n1126 | 1_n101;
assign 1_n487 = ~(1_n1485 | 1_n1560);
assign 1_n1026 = 1_n740;
assign 1_n774 = ~(1_n861 | 1_n1120);
assign 1_n764 = ~(1_n504 | 1_n1601);
assign 1_n1248 = ~(1_n1605 | 1_n209);
assign 1_n1113 = ~(1_n1427 | 1_n1058);
assign 1_n126 = ~(1_n1146 | 1_n1031);
assign 1_n1408 = ~1_n35;
assign 1_n1435 = 1_n1217 | 1_n108;
assign 1_n1073 = 1_n1369 & 1_n1515;
assign 1_n499 = 1_n511 | 1_n305;
assign 1_n1103 = ~(1_n1024 | 1_n336);
assign 1_n18 = ~(1_n934 | 1_n734);
assign 1_n1350 = 1_n278 | 1_n1266;
assign 1_n1500 = ~(1_n1391 | 1_n682);
assign 1_n298 = 1_n191 | 1_n583;
assign 1_n172 = ~(1_n1629 | 1_n1643);
assign 1_n600 = 1_n685 | 1_n1270;
assign 1_n1256 = 1_n1431 | 1_n547;
assign 1_n1072 = ~(1_n582 ^ 1_n788);
assign 1_n408 = ~(1_n1372 ^ 1_n426);
assign 1_n1584 = ~(1_n956 | 1_n344);
assign 1_n1634 = 1_n77 | 1_n398;
assign 1_n278 = 1_n361 & 1_n1165;
assign 1_n410 = 1_n832 & 1_n654;
assign 1_n1442 = 1_n574;
assign 1_n1364 = 1_n1539 | 1_n45;
assign 1_n1535 = ~1_n1413;
assign 1_n1090 = ~1_n1310;
assign 1_n1537 = ~1_n899;
assign 1_n1149 = ~1_n1243;
assign 1_n461 = ~1_n31;
assign 1_n850 = 1_n1651 | 1_n129;
assign 1_n1387 = 1_n251 & 1_n576;
assign 1_n180 = ~(1_n843 | 1_n566);
assign 1_n953 = ~(1_n152 | 1_n754);
assign 1_n910 = ~1_n1190;
assign 1_n62 = ~1_n1403;
assign 1_n779 = 1_n71 | 1_n50;
assign 1_n146 = 1_n1164 | 1_n828;
assign 1_n1492 = 1_n601 | 1_n508;
assign 1_n873 = ~(1_n1016 | 1_n1159);
assign 1_n1586 = ~(1_n1511 | 1_n1063);
assign 1_n354 = 1_n1368 & 1_n1116;
assign 1_n186 = ~1_n1372;
assign 1_n1662 = ~(1_n1245 | 1_n968);
assign 1_n868 = ~1_n760;
assign 1_n178 = ~(1_n1425 | 1_n352);
assign 1_n1489 = 1_n629 & 1_n325;
assign 1_n1433 = 1_n1647 & 1_n1121;
assign 1_n122 = 1_n637 | 1_n237;
assign 1_n745 = ~(1_n9 | 1_n227);
assign 1_n1202 = ~(1_n1093 | 1_n400);
assign 1_n1169 = 1_n1008 & 1_n283;
assign 1_n10 = ~1_n1033;
assign 1_n636 = 1_n708 | 1_n1010;
assign 1_n328 = ~(1_n557 ^ 1_n1484);
assign 1_n1183 = 1_n1007 & 1_n1005;
assign 1_n115 = ~1_n1663;
assign 1_n1132 = ~(1_n1388 | 1_n566);
assign 1_n578 = 1_n414 & 1_n938;
assign 1_n1484 = ~(1_n554 ^ 1_n1546);
assign 1_n152 = ~1_n536;
assign 1_n1031 = ~1_n1384;
assign 1_n856 = 1_n65 | 1_n436;
assign 1_n170 = 1_n163 | 1_n766;
assign 1_n1319 = 1_n626 | 1_n1501;
assign 1_n1315 = 1_n671 | 1_n832;
assign 1_n1194 = 1_n1629 | 1_n1050;
assign 1_n477 = 1_n2 | 1_n174;
assign 1_n1209 = 1_n1493 | 1_n1419;
assign 1_n1041 = ~(1_n1255 | 1_n859);
assign 1_n154 = 1_n478;
assign 1_n442 = 1_n206 | 1_n88;
assign 1_n915 = ~1_n1548;
assign 1_n963 = ~(1_n851 | 1_n34);
assign 1_n509 = ~1_n1406;
assign 1_n1235 = 1_n1205 | 1_n516;
assign 1_n238 = ~1_n507;
assign 1_n302 = 1_n1497 | 1_n17;
assign 1_n1671 = 1_n423 | 1_n1397;
assign 1_n541 = ~(1_n285 | 1_n1157);
assign 1_n652 = 1_n877 & 1_n182;
assign 1_n1589 = ~1_n889;
assign 1_n1009 = ~(1_n1191 ^ 1_n961);
assign 1_n1558 = ~(1_n1309 | 1_n1003);
assign 1_n249 = 1_n811 & 1_n1005;
assign 1_n1623 = ~(1_n222 | 1_n218);
assign 1_n1338 = 1_n412 & 1_n477;
assign 1_n1411 = ~(1_n1614 ^ 1_n260);
assign 1_n393 = 1_n235 & 1_n84;
assign 1_n809 = ~(1_n1255 | 1_n646);
assign 1_n1133 = 1_n1417 & 1_n1420;
assign 1_n1192 = 1_n1134;
assign 1_n1554 = ~1_n366;
assign 1_n1207 = ~1_n1534;
assign 1_n1122 = 1_n1510 | 1_n1085;
assign 1_n202 = 1_n681 & 1_n632;
assign 1_n1252 = ~(1_n1451 | 1_n1143);
assign 1_n1117 = 1_n110;
assign 1_n1574 = ~(1_n96 & 1_n1150);
assign 1_n994 = ~1_n1033;
assign 1_n755 = ~(1_n1467 | 1_n11);
assign 1_n430 = 1_n1654 & 1_n1005;
assign 1_n1097 = 1_n1503 & 1_n1655;
assign 1_n322 = ~(1_n897 | 1_n640);
assign 1_n735 = ~1_n1097;
assign 1_n494 = ~1_n1624;
assign 1_n879 = ~(1_n482 ^ 1_n1257);
assign 1_n1067 = ~1_n1448;
assign 1_n680 = 1_n327 | 1_n338;
assign 1_n1383 = ~(1_n1350 ^ 1_n1447);
assign 1_n1064 = 1_n1573;
assign 1_n1486 = 1_n1267 | 1_n29;
assign 1_n863 = 1_n1439 | 1_n1325;
assign 1_n1249 = ~(1_n765 | 1_n286);
assign 1_n1048 = ~(1_n329 | 1_n535);
assign 1_n92 = ~(1_n1274 | 1_n135);
assign 1_n892 = 1_n1251 & 1_n325;
assign 1_n246 = ~(1_n1213 | 1_n343);
assign 1_n1317 = ~1_n1377;
assign 1_n1628 = 1_n167 & 1_n794;
assign 1_n1080 = ~(1_n1534 | 1_n1636);
assign 1_n738 = ~(1_n113 ^ 1_n784);
assign 1_n1231 = 1_n1305 | 1_n791;
assign 1_n1119 = 1_n491 & 1_n1005;
assign 1_n1023 = 1_n1630;
assign 1_n661 = 1_n945 | 1_n315;
assign 1_n224 = 1_n421 & 1_n1412;
assign 1_n1295 = 1_n94 & 1_n720;
assign 1_n1225 = ~(1_n1523 | 1_n1395);
assign 1_n228 = ~(1_n1485 | 1_n34);
assign 1_n1314 = 1_n1490 | 1_n357;
assign 1_n265 = 1_n797 | 1_n1244;
assign 1_n1517 = 1_n1273 | 1_n1081;
assign 1_n1008 = ~(1_n1660 ^ 1_n1483);
assign 1_n1541 = ~1_n495;
assign 1_n1490 = 1_n1118 | 1_n1112;
assign 1_n1268 = ~1_n84;
assign 1_n573 = ~1_n1448;
assign 1_n472 = 1_n1212 | 1_n1340;
assign 1_n766 = 1_n431 | 1_n844;
assign 1_n271 = ~(1_n113 ^ 1_n16);
assign 1_n519 = ~(1_n1108 | 1_n1250);
assign 1_n922 = ~1_n857;
assign 1_n1201 = ~(1_n704 | 1_n1269);
assign 1_n458 = ~1_n859;
assign 1_n1380 = ~(1_n870 ^ 1_n339);
assign 1_n1522 = ~(1_n493 | 1_n35);
assign 1_n190 = 1_n761 | 1_n99;
assign 1_n919 = 1_n1677 | 1_n1423;
assign 1_n335 = ~(1_n1098 | 1_n1269);
assign 1_n1068 = ~(1_n147 | 1_n865);
assign 1_n48 = 1_n1338 & 1_n1540;
assign 1_n552 = ~(1_n386 | 1_n130);
assign 1_n1670 = 1_n585 & 1_n683;
assign 1_n1494 = ~(1_n418 | 1_n649);
assign 1_n741 = 1_n335 | 1_n460;
assign 1_n1672 = ~1_n590;
assign 1_n425 = ~(1_n1366 | 1_n218);
assign 1_n58 = ~(1_n435 | 1_n812);
assign 1_n1302 = 1_n912 | 1_n177;
assign 1_n223 = 1_n1251 & 1_n230;
assign 1_n423 = 1_n1322 | 1_n866;
assign 1_n1608 = ~1_n905;
assign 1_n1308 = ~1_n75;
assign 1_n1285 = ~1_n218;
assign 1_n886 = 1_n1675 & 1_n1161;
assign 1_n1334 = ~(1_n526 | 1_n668);
assign 1_n1156 = ~1_n939;
assign 1_n1230 = ~1_n1402;
assign 1_n1245 = ~1_n1351;
assign 1_n1395 = 1_n846 | 1_n86;
assign 1_n1005 = 1_n1445;
assign 1_n1488 = 1_n68 & 1_n1005;
assign 1_n143 = ~(1_n1578 | 1_n466);
assign 1_n1357 = 1_n517 & 1_n30;
assign 1_n109 = ~1_n1417;
assign 1_n348 = 1_n1551 & 1_n1655;
assign 1_n1421 = 1_n1555 | 1_n234;
assign 1_n1546 = 1_n560 | 1_n1429;
assign 1_n80 = ~(1_n1064 | 1_n1652);
assign 1_n762 = ~1_n1350;
assign 1_n1506 = 1_n487 | 1_n266;
assign 1_n1002 = 1_n936 & 1_n841;
assign 1_n980 = ~1_n569;
assign 1_n1242 = ~1_n225;
assign 1_n479 = ~(1_n443 ^ 1_n299);
assign 1_n1649 = 1_n153 | 1_n1018;
assign 1_n1392 = 1_n288 | 1_n337;
assign 1_n390 = ~(1_n1024 | 1_n1532);
assign 1_n993 = 1_n158 | 1_n294;
assign 1_n1173 = ~1_n1445;
assign 1_n663 = 1_n350;
assign 1_n218 = 1_n1362;
assign 1_n1461 = 1_n173 | 1_n687;
assign 1_n1234 = 1_n646 | 1_n1102;
assign 1_n525 = ~1_n57;
assign 1_n406 = ~1_n910;
assign 1_n321 = ~1_n1044;
assign 1_n162 = ~1_n1311;
assign 1_n1600 = ~(1_n1311 | 1_n1143);
assign 1_n105 = ~1_n1406;
assign 1_n366 = ~1_n1564;
assign 1_n674 = ~1_n950;
assign 1_n622 = ~1_n507;
assign 1_n1625 = 1_n1294 | 1_n755;
assign 1_n1139 = 1_n1353 | 1_n1037;
assign 1_n778 = ~1_n1141;
assign 1_n1643 = ~(1_n78 | 1_n813);
assign 1_n1284 = 1_n122 | 1_n748;
assign 1_n1385 = 1_n387 & 1_n1530;
assign 1_n1611 = ~(1_n1394 | 1_n1169);
assign 1_n1337 = ~1_n970;
assign 1_n996 = ~1_n661;
assign 1_n376 = ~(1_n811 ^ 1_n1500);
assign 1_n976 = 1_n1567 | 1_n447;
assign 1_n441 = ~1_n750;
assign 1_n1426 = ~(1_n238 | 1_n956);
assign 1_n947 = ~(1_n198 | 1_n606);
assign 1_n367 = ~(1_n769 | 1_n1246);
assign 1_n1568 = ~1_n138;
assign 1_n258 = ~(1_n67 | 1_n918);
assign 1_n1605 = ~1_n507;
assign 1_n1106 = ~1_n1300;
assign 1_n480 = 1_n132 & 1_n742;
assign 1_n1599 = 1_n609 | 1_n379;
assign 1_n551 = ~(1_n1187 | 1_n400);
assign 1_n1512 = 1_n194 | 1_n257;
assign 1_n1329 = ~(1_n51 | 1_n768);
assign 1_n139 = 1_n1066 | 1_n776;
assign 1_n897 = ~1_n31;
assign 1_n213 = ~(1_n1611 ^ 1_n891);
assign 1_n1665 = ~1_n1610;
assign 1_n1464 = ~(1_n1091 | 1_n406);
assign 1_n1638 = 1_n943 | 1_n420;
assign 1_n1552 = 1_n478;
assign 1_n1274 = ~1_n507;
assign 1_n1429 = ~(1_n1243 | 1_n352);
assign 1_n1236 = ~(1_n631 | 1_n695);
assign 1_n214 = ~(1_n1676 | 1_n1123);
assign 1_n332 = ~(1_n198 | 1_n977);
assign 1_n523 = 1_n512 | 1_n405;
assign 1_n1239 = 1_n984 | 1_n988;
assign 1_n124 = ~(1_n1306 ^ 1_n926);
assign 1_n874 = ~(1_n793 | 1_n311);
assign 1_n565 = 1_n1547;
assign 1_n787 = 1_n431 & 1_n632;
assign 1_n1376 = ~(1_n1425 | 1_n935);
assign 1_n318 = 1_n746 | 1_n312;
assign 1_n306 = ~1_n1498;
assign 1_n606 = ~1_n1143;
assign 1_n319 = ~(1_n1240 | 1_n709);
assign 1_n59 = 1_n932 | 1_n1638;
assign 1_n536 = ~1_n1307;
assign 1_n134 = ~1_n251;
assign 1_n351 = 1_n1258 | 1_n826;
assign 1_n1656 = ~(1_n659 ^ 1_n1616);
assign 1_n630 = ~(1_n1425 | 1_n72);
assign 1_n1138 = 1_n1629 | 1_n1553;
assign 1_n144 = 1_n824 & 1_n325;
assign 1_n1197 = ~(1_n300 | 1_n345);
assign 1_n926 = 1_n14 | 1_n1473;
assign 1_n20 = 1_n661 ^ 1_n1663;
assign 1_n40 = ~(1_n1427 | 1_n490);
assign 1_n1011 = 1_n70 | 1_n600;
assign 1_n1051 = 1_n727 & 1_n1606;
assign 1_n1228 = ~(1_n913 | 1_n888);
assign 1_n1127 = ~1_n1297;
assign 1_n1336 = ~1_n0;
assign 1_n439 = ~(1_n956 ^ 1_n1143);
assign 1_n1374 = ~1_n1405;
assign 1_n77 = 1_n995 & 1_n1555;
assign 1_n1401 = ~(1_n596 | 1_n525);
assign 1_n1615 = ~1_n1333;
assign 1_n1400 = 1_n1656 | 1_n721;
assign 1_n210 = ~1_n212;
assign 1_n33 = 1_n770 & 1_n1515;
assign 1_n807 = ~(1_n1311 | 1_n654);
assign 1_n56 = 1_n163 & 1_n632;
assign 1_n521 = 1_n391 | 1_n193;
assign 1_n98 = ~(1_n1352 ^ 1_n1370);
assign 1_n1118 = ~(1_n1162 | 1_n273);
assign 1_n1452 = ~(1_n568 | 1_n1507);
assign 1_n378 = ~(1_n1621 | 1_n722);
assign 1_n632 = 1_n771;
assign 1_n614 = 1_n991 | 1_n1622;
assign 1_n982 = 1_n1513 | 1_n1034;
assign 1_n1650 = ~1_n939;
assign 1_n1561 = ~(1_n1311 | 1_n677);
assign 1_n522 = 1_n1260 | 1_n333;
assign 1_n1227 = ~1_n1318;
assign 1_n1382 = 1_n1521 | 1_n942;
assign 1_n310 = 1_n609 | 1_n264;
assign 1_n1142 = 1_n852 | 1_n718;
assign 1_n1167 = ~(1_n152 | 1_n1355);
assign 1_n1459 = 1_n1428 & 1_n1549;
assign 1_n640 = ~1_n1059;
assign 1_n200 = ~(1_n1667 | 1_n562);
assign 1_n397 = ~1_n134;
assign 1_n875 = 1_n669 | 1_n1068;
assign 1_n1645 = ~1_n980;
assign 1_n1212 = 1_n817 | 1_n58;
assign 1_n1019 = 1_n1104 | 1_n146;
assign 1_n160 = ~(1_n1042 | 1_n1261);
assign 1_n1028 = ~(1_n1613 ^ 1_n136);
assign 1_n893 = ~1_n536;
assign 1_n1115 = ~(1_n144 | 1_n638);
assign 1_n456 = 1_n1487 | 1_n411;
assign 1_n719 = ~(1_n439 ^ 1_n879);
assign 1_n847 = ~1_n1647;
assign 1_n955 = 1_n27 | 1_n1263;
assign 1_n1205 = 1_n1390 & 1_n147;
assign 1_n1471 = 1_n151 & 1_n950;
assign 1_n1003 = ~1_n980;
assign 1_n782 = 1_n309 | 1_n986;
assign 1_n1328 = ~(1_n596 | 1_n1004);
assign 1_n1346 = ~(1_n1311 | 1_n824);
assign 1_n1669 = ~(1_n1144 ^ 1_n1444);
assign 1_n413 = 1_n572 | 1_n878;
assign 1_n1175 = ~1_n229;
assign 1_n1592 = ~1_n1029;
assign 1_n303 = ~1_n262;
assign 1_n253 = 1_n481;
assign 1_n860 = ~1_n1610;
assign 1_n865 = ~(1_n360 | 1_n830);
assign 1_n173 = 1_n946 | 1_n1132;
assign 1_n625 = 1_n1051 | 1_n831;
assign 1_n240 = 1_n1629 | 1_n723;
assign 1_n613 = ~(1_n659 ^ 1_n1006);
assign 1_n1172 = ~1_n1326;
assign 1_n819 = ~1_n1377;
assign 1_n503 = 1_n610 & 1_n79;
assign 1_n294 = ~(1_n1102 | 1_n1518);
assign 1_n448 = 1_n1455 & 1_n664;
assign 1_n374 = ~1_n652;
assign 1_n470 = ~(1_n1456 | 1_n725);
assign 1_n590 = 1_n655 | 1_n80;
assign 1_n6 = 1_n1518 & 1_n325;
assign 1_n324 = 1_n293;
assign 1_n742 = ~1_n932;
assign 1_n1640 = ~(1_n1441 ^ 1_n1380);
assign 1_n1601 = ~1_n1541;
assign 1_n1372 = 1_n799 | 1_n739;
assign 1_n1040 = 1_n25 | 1_n1270;
assign 1_n37 = 1_n458 | 1_n700;
assign 1_n694 = ~1_n1281;
assign 1_n350 = ~1_n128;
assign 1_n699 = 1_n1491 | 1_n1466;
assign 1_n156 = ~1_n218;
assign 1_n446 = ~1_n624;
assign 1_n889 = ~1_n1355;
assign 1_n1277 = 1_n267 & 1_n632;
assign 1_n639 = 1_n1609 | 1_n520;
assign 1_n1474 = 1_n1629 | 1_n1639;
assign 1_n1610 = ~1_n345;
assign 1_n407 = ~(1_n48 ^ 1_n112);
assign 1_n485 = ~1_n503;
assign 1_n1237 = 1_n673 & 1_n37;
assign 1_n870 = 1_n30 ^ 1_n1012;
assign 1_n1641 = 1_n223 | 1_n226;
assign 1_n650 = 1_n1401 | 1_n1505;
assign 1_n369 = ~(1_n661 | 1_n459);
assign 1_n103 = ~(1_n1581 | 1_n273);
assign 1_n1504 = 1_n209 & 1_n325;
assign 1_n817 = ~(1_n710 | 1_n819);
assign 1_n1571 = 1_n552 | 1_n308;
assign 1_n821 = 1_n1623 | 1_n1486;
assign 1_n1642 = 1_n1453 | 1_n876;
assign 1_n612 = ~(1_n1056 | 1_n1113);
assign 1_n653 = 1_n1526 | 1_n700;
assign 1_n1449 = ~(1_n1374 | 1_n686);
assign 1_n1034 = ~1_n597;
assign 1_n775 = 1_n1264 & 1_n1005;
assign 1_n958 = ~1_n730;
assign 1_n666 = 1_n214 | 1_n937;
assign 1_n420 = ~1_n647;
assign 1_n1195 = ~1_n853;
assign 1_n1668 = 1_n251 & 1_n1648;
assign 1_n708 = ~(1_n938 | 1_n188);
assign 1_n1544 = ~1_n57;
assign 1_n777 = ~1_n1563;
assign 1_n555 = ~(1_n1129 | 1_n392);
assign 1_n1044 = ~1_n1333;
assign 1_n999 = ~1_n1518;
assign 1_n1158 = ~(1_n403 | 1_n612);
assign 1_n678 = 1_n623;
assign 1_n388 = 1_n1013;
assign 1_n392 = 1_n36 | 1_n56;
assign 1_n114 = 1_n807 | 1_n410;
assign 1_n248 = ~(1_n1425 | 1_n1105);
assign 1_n344 = ~1_n365;
assign 1_n453 = ~(1_n1236 ^ 1_n580);
assign 1_n52 = 1_n499 & 1_n769;
assign 1_n452 = 1_n1586 | 1_n1167;
assign 1_n95 = ~(1_n1165 | 1_n1458);
assign 1_n39 = 1_n1407 & 1_n1243;
assign 1_n207 = ~1_n348;
assign 1_n31 = ~1_n1172;
assign 1_n903 = ~(1_n531 | 1_n92);
assign 1_n795 = ~(1_n1324 | 1_n624);
assign 1_n102 = 1_n1030 & 1_n230;
assign 1_n409 = 1_n157 | 1_n966;
assign 1_n559 = 1_n1285 & 1_n1508;
assign 1_n1213 = ~1_n730;
assign 1_n1082 = ~(1_n470 | 1_n1472);
assign 1_n1241 = 1_n407 | 1_n409;
assign 1_n3 = 1_n1328 | 1_n1197;
assign 1_n603 = ~(1_n120 | 1_n1661);
assign 1_n831 = ~(1_n1606 | 1_n935);
assign 1_n562 = 1_n595 | 1_n1486;
assign 1_n608 = 1_n1596;
assign 1_n450 = ~(1_n215 | 1_n1060);
assign 1_n1455 = ~1_n218;
assign 1_n236 = ~1_n365;
assign 1_n1096 = 1_n979 | 1_n1488;
assign 1_n166 = ~1_n1230;
assign 1_n1370 = ~(1_n921 ^ 1_n408);
assign 1_n840 = 1_n1629 | 1_n534;
assign 1_n308 = ~(1_n10 | 1_n345);
assign 1_n428 = ~(1_n1425 | 1_n1053);
assign 1_n508 = ~(1_n198 | 1_n55);
assign 1_n1290 = 1_n1153 & 1_n182;
assign 1_n643 = 1_n589 | 1_n1662;
assign 1_n252 = ~(1_n1435 ^ 1_n1108);
assign 1_n1066 = 1_n1460 & 1_n1049;
assign 1_n358 = ~1_n1001;
assign 1_n983 = 1_n796 & 1_n589;
assign 1_n1354 = 1_n252 | 1_n1171;
assign 1_n1458 = ~(1_n1653 | 1_n40);
assign 1_n987 = 1_n1223 & 1_n1606;
assign 1_n1004 = ~1_n868;
assign 1_n1536 = ~1_n1432;
assign 1_n838 = 1_n1338 & 1_n1663;
assign 1_n1607 = ~(1_n1280 | 1_n311);
assign 1_n1520 = ~1_n394;
assign 1_n604 = ~1_n509;
assign 1_n707 = ~1_n182;
assign 1_n241 = ~(1_n1452 ^ 1_n636);
assign 1_n1664 = ~(1_n1425 | 1_n1545);
assign 1_n855 = ~1_n1545;
assign 1_n1444 = ~(1_n564 ^ 1_n850);
assign 1_n528 = ~(1_n1569 ^ 1_n175);
assign 1_n383 = 1_n1387 | 1_n1222;
assign 1_n433 = ~(1_n1581 | 1_n1123);
assign 1_n148 = ~1_n306;
assign 1_n830 = ~(1_n1425 | 1_n55);
assign 1_n530 = ~1_n229;
assign 1_n790 = ~(1_n1562 & 1_n128);
assign 1_n539 = ~(1_n769 | 1_n1228);
assign 1_n1035 = 1_n1447 ^ 1_n823;
assign 1_n1448 = ~1_n1379;
assign 1_n760 = ~1_n1193;
assign 1_n312 = 1_n1229 | 1_n970;
assign 1_n42 = ~1_n1318;
assign 1_n276 = 1_n646 & 1_n325;
assign 1_n1588 = 1_n452 | 1_n1642;
assign 1_n1174 = 1_n1579 | 1_n907;
assign 1_n712 = 1_n1069 | 1_n377;
assign 1_n1318 = ~1_n994;
assign 1_n263 = ~(1_n622 | 1_n1030);
assign 1_n1196 = 1_n1245 | 1_n982;
assign 1_n372 = 1_n801 & 1_n1196;
assign 1_n457 = ~(1_n346 | 1_n827);
assign 1_n78 = 1_n1433 | 1_n1291;
assign 1_n960 = ~1_n507;
assign 1_n465 = ~(1_n604 | 1_n316);
assign 1_n1616 = 1_n873 | 1_n643;
assign 1_n1456 = ~1_n274;
assign 1_n363 = 1_n808 | 1_n1220;
assign 1_n1286 = ~1_n1190;
assign 1_n76 = 1_n1629 | 1_n1588;
assign 1_n338 = 1_n331 & 1_n1005;
assign 1_n243 = ~(1_n468 | 1_n1317);
assign 1_n359 = 1_n1101 ^ 1_n438;
assign 1_n1591 = 1_n1583 | 1_n599;
assign 1_n336 = ~1_n446;
assign 1_n1332 = ~(1_n1617 ^ 1_n20);
assign 1_n1360 = ~1_n63;
assign 1_n944 = ~(1_n1184 | 1_n1544);
assign 1_n553 = 1_n271 & 1_n632;
assign 1_n391 = ~1_n1240;
assign 1_n1420 = ~(1_n1572 ^ 1_n950);
assign 1_n1391 = ~(1_n184 | 1_n450);
assign 1_n197 = 1_n802 | 1_n1312;
assign 1_n1550 = 1_n160 | 1_n119;
assign 1_n1006 = ~(1_n1159 ^ 1_n234);
assign 1_n1087 = ~1_n293;
assign 1_n951 = ~1_n446;
assign 1_n462 = ~1_n252;
assign 1_n435 = ~1_n105;
assign 1_n1124 = ~(1_n923 | 1_n374);
assign 1_n53 = ~(1_n479 | 1_n1368);
assign 1_n414 = 1_n314 | 1_n211;
assign 1_n1667 = ~1_n1300;
assign 1_n568 = ~(1_n147 | 1_n1136);
assign 1_n1263 = ~(1_n494 | 1_n887);
assign 1_n1152 = ~1_n1606;
assign 1_n866 = ~(1_n285 | 1_n250);
assign 1_n164 = ~(1_n617 | 1_n1426);
assign 1_n482 = ~(1_n1030 ^ 1_n1251);
assign 1_n584 = ~(1_n710 | 1_n1022);
assign 1_n1321 = ~(1_n654 ^ 1_n490);
assign 1_n878 = ~(1_n1062 | 1_n503);
assign 1_n266 = ~(1_n893 | 1_n394);
assign 1_n411 = ~(1_n1106 | 1_n434);
assign 1_n334 = ~(1_n329 | 1_n1665);
assign 1_n90 = ~(1_n1243 | 1_n884);
assign 1_n361 = 1_n987 | 1_n85;
assign 1_n1451 = ~1_n365;
assign 1_n179 = ~1_n705;
assign 1_n280 = ~1_n48;
assign 1_n1379 = 1_n1535 & 1_n989;
assign 1_n1306 = ~(1_n733 | 1_n1674);
assign 1_n802 = ~(1_n362 | 1_n321);
assign 1_n257 = 1_n87 | 1_n703;
assign 1_n74 = 1_n744 | 1_n1519;
assign 1_n1673 = ~(1_n417 | 1_n603);
assign 1_n665 = ~1_n1568;
assign 1_n279 = ~(1_n67 | 1_n1004);
assign 1_n323 = 1_n1571 | 1_n581;
assign 1_n556 = 1_n522 & 1_n1479;
assign 1_n992 = ~1_n149;
assign 1_n269 = 1_n456 | 1_n767;
assign 1_n127 = ~1_n1389;
assign 1_n569 = 1_n89 | 1_n553;
assign 1_n1024 = ~1_n1342;
assign 1_n1585 = 1_n1030 & 1_n325;
assign 1_n498 = ~(1_n290 | 1_n1175);
assign 1_n1513 = ~1_n1271;
assign 1_n239 = ~(1_n198 | 1_n855);
assign 1_n1300 = ~1_n1172;
assign 1_n633 = 1_n3 | 1_n1649;
assign 1_n709 = ~(1_n858 | 1_n1178);
assign 1_n355 = ~(1_n1479 | 1_n164);
assign 1_n1467 = ~1_n393;
assign 1_n833 = 1_n1285 & 1_n1131;
assign 1_n1157 = ~1_n1233;
assign 1_n1111 = ~(1_n1575 ^ 1_n1161);
assign 1_n368 = ~(1_n693 ^ 1_n930);
assign 1_n537 = ~(1_n950 | 1_n542);
assign 1_n679 = 1_n1661 ^ 1_n331;
assign 1_n1222 = 1_n1428 & 1_n1052;
assign 1_n998 = ~1_n1030;
assign 1_n88 = ~(1_n1227 | 1_n250);
assign 1_n1533 = ~(1_n504 | 1_n624);
assign 1_n1089 = 1_n634 | 1_n255;
assign 1_n792 = ~(1_n587 ^ 1_n804);
assign 1_n1029 = 1_n139 | 1_n317;
assign 1_n1566 = 1_n1633 | 1_n1558;
assign 1_n1102 = ~1_n365;
assign 1_n563 = 1_n471 | 1_n486;
assign 1_n1590 = ~1_n1411;
assign 1_n1086 = ~1_n1606;
assign 1_n436 = ~(1_n42 | 1_n1345);
assign 1_n1216 = 1_n1078 | 1_n575;
assign 1_n235 = ~1_n726;
assign 1_n852 = 1_n648 & 1_n635;
assign 1_n1206 = ~(1_n1324 | 1_n495);
assign 1_n307 = ~(1_n1578 | 1_n781);
assign 1_n1144 = ~(1_n743 ^ 1_n234);
assign 1_n155 = 1_n51 ^ 1_n738;
assign 1_n49 = 1_n1025 & 1_n1606;
assign 1_n1639 = 1_n1566 | 1_n1083;
assign 1_n17 = ~(1_n303 | 1_n1355);
assign 1_n225 = 1_n127 | 1_n384;
assign 1_n340 = ~(1_n463 | 1_n495);
assign 1_n1358 = ~1_n403;
assign 1_n1473 = 1_n1040 & 1_n1640;
assign 1_n1092 = ~(1_n1462 | 1_n1385);
assign 1_n326 = 1_n498 | 1_n1666;
assign 1_n1646 = ~1_n770;
assign 1_n757 = ~1_n1360;
assign 1_n1114 = 1_n929 & 1_n1475;
assign 1_n975 = ~(1_n554 ^ 1_n765);
assign 1_n1289 = ~1_n676;
assign 1_n237 = ~(1_n938 | 1_n440);
assign 1_n1603 = ~1_n1351;
assign 1_n14 = ~(1_n1299 | 1_n1040);
assign 1_n984 = ~1_n1150;
assign 1_n1622 = 1_n429 | 1_n1207;
assign 1_n455 = 1_n881 | 1_n1349;
assign 1_n681 = ~(1_n527 ^ 1_n1231);
assign 1_n691 = 1_n619 | 1_n15;
assign 1_n743 = 1_n798 | 1_n1057;
assign 1_n885 = 1_n1460 & 1_n1189;
assign 1_n502 = ~(1_n463 | 1_n951);
assign 1_n732 = 1_n1644 | 1_n1252;
assign 1_n570 = ~1_n996;
assign 1_n11 = ~1_n1440;
assign 1_n693 = ~1_n627;
assign 1_n812 = 1_n871 | 1_n1277;
assign 1_n1390 = 1_n1450 | 1_n1363;
assign 1_n474 = ~(1_n435 | 1_n469);
assign 1_n959 = ~1_n1436;
assign 1_n1462 = ~(1_n1530 | 1_n1115);
assign 1_n548 = ~(1_n461 | 1_n244);
assign 1_n669 = 1_n1641 & 1_n147;
assign 1_n1164 = ~1_n1630;
assign 1_n1293 = ~(1_n1361 | 1_n374);
assign 1_n136 = ~(1_n135 ^ 1_n824);
assign 1_n585 = 1_n1378 | 1_n1415;
assign 1_n1309 = ~1_n1379;
assign 1_n301 = ~1_n113;
assign 1_n626 = ~(1_n1389 | 1_n19);
assign 1_n377 = ~(1_n461 | 1_n590);
assign 1_n1675 = ~1_n1606;
assign 1_n1469 = 1_n419 | 1_n372;
assign 1_n941 = 1_n1455 & 1_n716;
assign 1_n1059 = ~1_n250;
assign 1_n914 = 1_n60 & 1_n1620;
assign 1_n1652 = ~(1_n1308 ^ 1_n246);
assign 1_n723 = 1_n1182 | 1_n1506;
assign 1_n979 = 1_n395 & 1_n233;
assign 1_n1569 = ~(1_n597 | 1_n846);
assign 1_n1457 = ~1_n316;
assign 1_n776 = 1_n191 & 1_n1005;
assign 1_n460 = ~(1_n974 | 1_n1204);
assign 1_n843 = ~1_n509;
assign 1_n1415 = ~(1_n809 | 1_n428);
assign 1_n1171 = 1_n43 | 1_n217;
assign 1_n129 = ~(1_n1606 | 1_n999);
assign 1_n978 = 1_n74 | 1_n1084;
assign 1_n1120 = ~1_n1541;
assign 1_n229 = ~1_n207;
assign 1_n1063 = ~1_n910;
assign 1_n620 = ~(1_n895 | 1_n445);
assign 1_n1057 = 1_n1086 & 1_n1575;
assign 1_n581 = 1_n1424 | 1_n1347;
assign 1_n288 = 1_n258 | 1_n1103;
assign 1_n1081 = ~(1_n346 | 1_n1589);
assign 1_n1659 = 1_n485 | 1_n778;
assign 1_n157 = ~(1_n125 ^ 1_n779);
assign 1_n648 = ~1_n218;
assign 1_n1232 = 1_n1148 | 1_n1675;
assign 1_n341 = ~(1_n1064 | 1_n213);
assign 1_n896 = ~(1_n1101 ^ 1_n924);
assign 1_n1077 = ~(1_n981 | 1_n1626);
assign 1_n705 = 1_n922 | 1_n1207;
assign 1_n113 = ~(1_n254 ^ 1_n1240);
assign 1_n1298 = 1_n1133 | 1_n1080;
assign 1_n554 = 1_n1100 | 1_n12;
assign 1_n827 = 1_n1096 | 1_n1020;
assign 1_n1126 = 1_n833 | 1_n775;
assign 1_n977 = ~1_n859;
assign 1_n1075 = ~(1_n1064 | 1_n1337);
assign 1_n940 = ~1_n1110;
assign 1_n1341 = ~(1_n1070 | 1_n1259);
assign 1_n744 = ~1_n785;
assign 1_n935 = ~1_n1058;
assign 1_n763 = ~(1_n399 ^ 1_n1111);
assign 1_n770 = 1_n726 & 1_n84;
assign 1_n557 = ~(1_n1038 ^ 1_n254);
assign 1_n645 = 1_n216 & 1_n632;
assign 1_n1553 = 1_n782 | 1_n955;
assign 1_n1621 = ~1_n1326;
assign 1_n133 = ~1_n812;
assign 1_n948 = ~1_n198;
assign 1_n1351 = ~1_n187;
assign 1_n908 = ~1_n1646;
assign 1_n1078 = 1_n60 & 1_n1418;
assign 1_n997 = 1_n1348 & 1_n1413;
assign 1_n1094 = 1_n850 & 1_n769;
assign 1_n533 = ~(1_n1608 | 1_n827);
assign 1_n426 = ~(1_n281 ^ 1_n1570);
assign 1_n1218 = ~(1_n1274 | 1_n1251);
assign 1_n1259 = ~1_n397;
assign 1_n832 = ~1_n198;
assign 1_n149 = 1_n564 ^ 1_n1378;
assign 1_n217 = 1_n915 | 1_n47;
assign 1_n957 = 1_n586 | 1_n219;
assign 1_n251 = 1_n1537 & 1_n270;
assign 1_n767 = 1_n1224 | 1_n533;
assign 1_n379 = ~1_n725;
assign 1_n1377 = ~1_n611;
assign 1_n153 = ~(1_n1014 | 1_n668);
assign 1_n594 = ~(1_n414 ^ 1_n1390);
assign 1_n1501 = 1_n114 & 1_n1389;
assign 1_n567 = ~(1_n923 | 1_n530);
assign 1_n5 = ~(1_n1129 | 1_n928);
assign 1_n1587 = ~1_n566;
assign 1_n1233 = ~1_n1283;
assign 1_n159 = ~(1_n1438 | 1_n1204);
assign 1_n1381 = ~1_n574;
assign 1_n63 = ~1_n997;
assign 1_n967 = ~(1_n1425 | 1_n458);
assign 1_n1141 = 1_n389 & 1_n1538;
assign 1_n429 = 1_n881 | 1_n720;
assign 1_n752 = ~(1_n1425 | 1_n606);
assign 1_n1221 = 1_n898 | 1_n334;
assign 1_n697 = ~1_n1572;
assign 1_n1186 = ~1_n692;
assign 1_n799 = 1_n1161 & 1_n198;
assign 1_n920 = ~1_n1302;
assign 1_n311 = ~1_n1193;
assign 1_n12 = ~(1_n1243 | 1_n1105);
assign 1_n1305 = 1_n1516 & 1_n857;
assign 1_n711 = 1_n551 | 1_n340;
assign 1_n205 = 1_n1210 & 1_n403;
assign 1_n46 = ~1_n1670;
assign 1_n883 = ~(1_n1386 | 1_n630);
assign 1_n256 = ~1_n825;
assign 1_n1404 = ~1_n1247;
assign 1_n492 = ~(1_n358 | 1_n1141);
assign 1_n177 = 1_n1565 | 1_n341;
assign 1_n616 = 1_n906 | 1_n1301;
assign 1_n641 = 1_n993 & 1_n769;
assign 1_n690 = 1_n1268 & 1_n235;
assign 1_n1027 = ~(1_n1425 | 1_n884);
assign 1_n912 = 1_n901 & 1_n1065;
assign 1_n1021 = 1_n476 | 1_n1514;
assign 1_n1299 = ~(1_n1383 ^ 1_n1076);
assign 1_n1365 = 1_n488 & 1_n1503;
assign 1_n1074 = ~1_n1034;
assign 1_n167 = ~1_n899;
assign 1_n1254 = 1_n696 & 1_n393;
assign 1_n292 = ~1_n1134;
assign 1_n1539 = 1_n135 & 1_n230;
assign 1_n171 = ~(1_n1187 | 1_n189);
assign 1_n399 = ~(1_n646 ^ 1_n1518);
assign 1_n658 = 1_n501 | 1_n1533;
assign 1_n1125 = 1_n545 & 1_n1033;
assign 1_n601 = ~(1_n1311 | 1_n1251);
assign 1_n1431 = 1_n1168 | 1_n1183;
assign 1_n1367 = ~1_n1001;
assign 1_n1053 = ~1_n646;
assign 1_n1327 = ~(1_n1522 ^ 1_n359);
assign 1_n299 = ~(1_n1617 ^ 1_n1282);
assign 1_n1016 = ~1_n1555;
assign 1_n295 = 1_n1058 & 1_n230;
assign 1_n609 = ~1_n381;
assign 1_n44 = 1_n1149 & 1_n677;
assign 1_n1200 = ~1_n664;
assign 1_n1265 = 1_n762 & 1_n730;
assign 1_n1271 = ~(1_n161 ^ 1_n1545);
assign 1_n881 = ~1_n301;
assign 1_n26 = ~1_n1369;
assign 1_n796 = ~1_n659;
assign 1_n676 = ~(1_n328 ^ 1_n1009);
assign 1_n1423 = ~(1_n1410 | 1_n696);
assign 1_n905 = ~1_n66;
assign 1_n583 = 1_n549 | 1_n46;
assign 1_n212 = ~1_n686;
assign 1_n89 = 1_n1114 | 1_n249;
assign 1_n272 = ~1_n105;
assign 1_n510 = ~(1_n1255 | 1_n824);
assign 1_n898 = ~(1_n386 | 1_n1199);
assign 1_n264 = ~1_n1563;
assign 1_n561 = ~(1_n1255 | 1_n1143);
assign 1_n1470 = 1_n1606 | 1_n671;
assign 1_n662 = ~(1_n958 | 1_n181);
assign 1_n82 = 1_n872 | 1_n1179;
assign 1_n1151 = 1_n1577 | 1_n803;
assign 1_n316 = 1_n680 | 1_n1075;
assign 1_n722 = ~1_n1457;
assign 1_n1393 = ~(1_n1608 | 1_n1262);
assign 1_n195 = 1_n648 & 1_n1303;
assign 1_n1226 = ~(1_n1271 ^ 1_n1225);
assign 1_n1538 = 1_n1493 | 1_n1237;
assign 1_n497 = ~1_n994;
assign 1_n651 = 1_n963 | 1_n502;
assign 1_n929 = ~1_n218;
assign 1_n1278 = ~(1_n330 | 1_n1259);
assign 1_n566 = 1_n185 | 1_n972;
assign 1_n1203 = 1_n467 & 1_n1005;
assign 1_n619 = 1_n1061 | 1_n247;
assign 1_n349 = ~(1_n418 | 1_n62);
assign 1_n1627 = ~(1_n1092 ^ 1_n957);
assign 1_n1267 = ~(1_n1536 | 1_n98);
assign 1_n689 = 1_n1135 | 1_n1125;
assign 1_n101 = ~(1_n1064 | 1_n729);
assign 1_n424 = ~1_n868;
assign 1_n108 = ~(1_n1243 | 1_n606);
assign 1_n729 = ~(1_n911 ^ 1_n1130);
assign 1_n221 = ~1_n262;
assign 1_n1137 = ~1_n1097;
assign 1_n1560 = ~1_n1286;
assign 1_n412 = 1_n1186 | 1_n109;
assign 1_n749 = 1_n353 & 1_n1479;
assign 1_n1660 = ~(1_n1327 ^ 1_n546);
assign 1_n628 = 1_n1176 | 1_n332;
assign 1_n1579 = ~(1_n362 | 1_n227);
assign 1_n871 = 1_n941 | 1_n422;
assign 1_n624 = 1_n287 | 1_n645;
assign 1_n970 = ~(1_n1213 ^ 1_n343);
assign 1_n968 = ~1_n731;
assign 1_n800 = ~1_n629;
assign 1_n1559 = 1_n1201 | 1_n159;
assign 1_n942 = 1_n948 & 1_n490;
assign 1_n27 = ~(1_n1093 | 1_n189);
assign 1_n70 = ~1_n762;
assign 1_n1503 = ~1_n1551;
assign 1_n371 = 1_n1319 & 1_n1005;
assign 1_n1345 = ~1_n212;
assign 1_n451 = ~1_n497;
assign 1_n68 = 1_n880 | 1_n1249;
assign 1_n138 = ~1_n1369;
assign 1_n417 = 1_n1200 & 1_n120;
assign 1_n1478 = ~1_n1672;
assign 1_n1595 = ~(1_n494 | 1_n621);
assign 1_n687 = 1_n111 | 1_n457;
assign 1_n488 = ~1_n1655;
assign 1_n599 = 1_n1149 & 1_n268;
assign 1_n826 = 1_n1652 & 1_n120;
assign 1_n1612 = ~(1_n990 | 1_n148);
assign 1_n1534 = ~1_n217;
assign 1_n1180 = 1_n1276 & 1_n1396;
assign 1_n1353 = ~(1_n909 | 1_n670);
assign 1_n924 = 1_n179 | 1_n1417;
assign 1_n1264 = 1_n95 | 1_n22;
assign 1_n637 = 1_n41 & 1_n938;
assign 1_n274 = 1_n414 ^ 1_n938;
assign 1_n1128 = ~(1_n613 ^ 1_n528);
assign 1_n1564 = ~1_n274;
assign 1_n357 = 1_n1602 | 1_n390;
assign 1_n647 = 1_n591 & 1_n1603;
assign 1_n773 = ~1_n652;
assign 1_n1410 = ~1_n905;
assign 1_n659 = ~(1_n850 ^ 1_n769);
assign 1_n816 = ~(1_n793 | 1_n259);
assign 1_n527 = ~(1_n1524 ^ 1_n1479);
assign 1_n931 = 1_n109 & 1_n777;
assign 1_n1260 = ~(1_n1311 | 1_n956);
assign 1_n1032 = 1_n441 | 1_n1087;
assign 1_n853 = ~1_n1402;
assign 1_n131 = 1_n896 | 1_n1241;
assign 1_n571 = ~(1_n381 | 1_n1456);
assign 1_n1304 = ~1_n550;
assign 1_n1556 = 1_n829;
assign 1_n575 = 1_n875 & 1_n1005;
assign 1_n317 = 1_n1656 & 1_n632;
assign 1_n234 = 1_n297;
assign 1_n1291 = 1_n562 & 1_n690;
assign 1_n188 = ~(1_n1585 | 1_n263);
assign 1_n867 = 1_n607 | 1_n953;
assign 1_n118 = ~(1_n1304 ^ 1_n1082);
assign 1_n1330 = ~(1_n198 | 1_n998);
assign 1_n1038 = 1_n1017 | 1_n602;
assign 1_n1155 = ~1_n1652;
assign 1_n939 = ~1_n760;
assign 1_n1532 = ~1_n1557;
assign 1_n1430 = 1_n49 | 1_n904;
assign 1_n546 = ~(1_n756 ^ 1_n310);
assign 1_n51 = 1_n1414 | 1_n369;
assign 1_n1527 = ~(1_n276 | 1_n1316);
assign 1_n692 = ~1_n252;
assign 1_n64 = 1_n952 | 1_n919;
assign 1_n1463 = ~(1_n282 ^ 1_n1597);
assign 1_n8 = ~1_n1150;
assign 1_n1208 = ~(1_n1311 | 1_n1058);
assign 1_n1674 = 1_n1072 & 1_n1;
assign 1_n1182 = 1_n810 | 1_n474;
assign 1_n285 = ~1_n1281;
assign 1_n440 = ~(1_n806 | 1_n1598);
assign 1_n899 = ~1_n224;
assign 1_n1406 = ~1_n690;
assign 1_n937 = ~(1_n221 | 1_n392);
assign 1_n501 = ~(1_n851 | 1_n406);
assign 1_n1414 = 1_n1546 & 1_n1530;
assign 1_n1348 = ~1_n989;
assign 1_n247 = ~(1_n694 | 1_n812);
assign 1_n820 = 1_n784 | 1_n936;
assign 1_n1323 = ~(1_n689 | 1_n505);
assign 1_n538 = ~(1_n1479 | 1_n883);
assign 1_n627 = ~1_n1155;
assign 1_n1355 = 1_n1216 | 1_n201;
assign 1_n673 = 1_n859 | 1_n1451;
assign 1_n15 = 1_n396 | 1_n1206;
assign 1_n668 = ~1_n348;
assign 1_n1177 = ~1_n1592;
assign 1_n758 = 1_n816 | 1_n73;
assign 1_n346 = ~1_n1067;
assign 1_n1677 = ~(1_n1280 | 1_n259);
assign 1_n1325 = 1_n846 & 1_n1271;
assign 1_n1403 = ~1_n63;
assign 1_n1352 = ~(1_n679 ^ 1_n1107);
assign 1_n61 = 1_n845;
assign 1_n1446 = 1_n592 & 1_n653;
assign 1_n544 = ~1_n1044;
assign 1_n273 = ~1_n853;
assign 1_n564 = 1_n1618 | 1_n529;
assign 1_n602 = ~(1_n1243 | 1_n977);
assign 1_n547 = 1_n896 & 1_n632;
assign 1_n798 = 1_n1606 & 1_n588;
assign 1_n489 = 1_n350;
assign 1_n196 = ~1_n827;
assign 1_n1110 = ~1_n784;
assign 1_n642 = 1_n549 & 1_n1005;
assign 1_n784 = ~(1_n1038 ^ 1_n184);
assign 1_n1045 = ~(1_n381 ^ 1_n1235);
assign 1_n395 = ~1_n218;
assign 1_n813 = 1_n33 | 1_n1254;
assign 1_n1297 = ~1_n958;
assign 1_n1498 = ~1_n1428;
assign 1_n549 = 1_n1088 | 1_n1664;
assign 1_n1526 = ~1_n824;
assign 1_n30 = ~1_n911;
assign 1_n1326 = 1_n707 & 1_n1153;
assign 1_n337 = 1_n1509 | 1_n378;
assign 1_n785 = ~(1_n1028 ^ 1_n719);
assign 1_n505 = 1_n1073 | 1_n370;
assign 1_n211 = ~(1_n1243 | 1_n998);
assign 1_n731 = ~1_n992;
assign 1_n783 = ~(1_n236 | 1_n209);
assign 1_n780 = 1_n1561 | 1_n1279;
assign 1_n1136 = ~(1_n892 | 1_n1218);
assign 1_n928 = ~1_n1557;
assign 1_n595 = 1_n837 & 1_n1065;
assign 1_n1047 = ~(1_n1513 ^ 1_n753);
assign 1_n384 = ~1_n1430;
assign 1_n1168 = 1_n1465 & 1_n432;
assign 1_n841 = 1_n975 | 1_n459;
assign 1_n925 = 1_n991 ^ 1_n1548;
assign 1_n291 = ~1_n133;
assign 1_n353 = 1_n1296 | 1_n1584;
assign 1_n995 = ~1_n982;
assign 1_n1509 = ~(1_n1373 | 1_n773);
assign 1_n513 = 1_n157 & 1_n632;
assign 1_n1521 = ~(1_n1311 | 1_n490);
assign 1_n1460 = ~1_n218;
assign 1_n724 = 1_n1469 & 1_n1054;
assign 1_n686 = 1_n1142 | 1_n667;
assign 1_n158 = 1_n1518 & 1_n230;
assign 1_n1000 = ~(1_n818 | 1_n1650);
assign 1_n1270 = ~1_n724;
assign 1_n16 = ~(1_n1295 | 1_n834);
assign 1_n1597 = ~(1_n1395 ^ 1_n234);
assign 1_n315 = ~1_n554;
assign 1_n1637 = ~(1_n35 ^ 1_n925);
assign 1_n1388 = ~1_n497;
assign 1_n38 = 1_n126 | 1_n180;
assign 1_n1279 = 1_n948 & 1_n677;
assign 1_n215 = 1_n859 & 1_n325;
assign 1_n1495 = ~1_n1530;
assign 1_n459 = ~(1_n1546 ^ 1_n1530);
assign 1_n380 = 1_n496 | 1_n1393;
assign 1_n1054 = 1_n1358 | 1_n1288;
assign 1_n660 = ~(1_n1311 | 1_n209);
assign 1_n1666 = ~(1_n303 | 1_n675);
assign 1_n1104 = ~1_n829;
assign 1_n1363 = ~(1_n1243 | 1_n55);
assign 1_n305 = ~(1_n198 | 1_n999);
assign 1_n1528 = ~(1_n869 | 1_n1673);
assign 1_n1523 = 1_n1074 & 1_n1555;
assign 1_n176 = 1_n660 | 1_n1188;
assign 1_n1101 = ~1_n462;
assign 1_n943 = ~1_n1357;
assign 1_n405 = ~1_n296;
assign 1_n577 = 1_n149 & 1_n1603;
assign 1_n904 = 1_n1086 & 1_n654;
assign 1_n1482 = ~1_n1420;
assign 1_n404 = ~(1_n1030 | 1_n344);
assign 1_n772 = ~(1_n1255 | 1_n1058);
assign 1_n1312 = ~(1_n861 | 1_n569);
assign 1_n1542 = 1_n750;
assign 1_n845 = ~1_n128;
assign 1_n917 = 1_n209 & 1_n230;
assign 1_n945 = ~1_n765;
assign 1_n1543 = 1_n780 & 1_n1240;
assign 1_n1116 = ~(1_n155 ^ 1_n1332);
assign 1_n1563 = ~1_n1482;
assign 1_n1614 = ~(1_n1109 ^ 1_n1321);
assign 1_n535 = ~1_n1672;
assign 1_n192 = ~(1_n1467 | 1_n569);
assign 1_n1056 = 1_n1058 & 1_n325;
assign 1_n1624 = ~1_n1307;
assign 1_n572 = 1_n156 & 1_n973;
assign 1_n142 = 1_n614;
assign 1_n1266 = ~(1_n225 | 1_n911);
assign 1_n696 = ~1_n920;
assign 1_n969 = 1_n1208 | 1_n1287;
assign 1_n193 = ~1_n254;
assign 1_n656 = ~1_n1084;
assign 1_n918 = ~1_n1615;
assign 1_n36 = 1_n195 | 1_n91;
assign 1_n1017 = 1_n137 & 1_n1243;
assign 1_n1598 = ~(1_n1425 | 1_n998);
assign 1_n916 = 1_n642 | 1_n885;
assign 1_n1445 = 1_n1071 & 1_n558;
assign 1_n932 = 1_n1145 | 1_n702;
assign 1_n1176 = ~(1_n1311 | 1_n859);
assign 1_n1166 = ~1_n562;
assign 1_n1573 = 1_n1065 | 1_n558;
assign 1_n1071 = ~1_n1065;
assign 1_n1405 = ~1_n518;
assign 1_n469 = ~1_n1059;
assign 1_n1572 = 1_n1525 | 1_n90;
assign 1_n1238 = ~(1_n934 | 1_n1477);
assign 1_n1349 = 1_n1295 | 1_n838;
assign 1_n1198 = 1_n302 | 1_n684;
assign 1_n345 = 1_n715 | 1_n123;
assign 1_n715 = 1_n914 | 1_n1119;
assign 1_n1481 = 1_n1012 & 1_n225;
assign 1_n1160 = 1_n1629 | 1_n815;
assign 1_n804 = ~(1_n822 ^ 1_n688);
assign 1_n1441 = ~(1_n1447 ^ 1_n181);
assign 1_n756 = ~(1_n1516 | 1_n791);
assign 1_n1069 = ~(1_n526 | 1_n773);
assign 1_n1147 = ~1_n1661;
assign 1_n1362 = 1_n532 | 1_n1071;
assign 1_n329 = ~1_n690;
assign 1_n86 = 1_n597 & 1_n234;
assign 1_n1582 = 1_n875 | 1_n1476;
assign 1_n1602 = ~(1_n9 | 1_n544);
assign 1_n1281 = ~1_n518;
assign 1_n132 = 1_n1095 & 1_n1265;
assign 1_n267 = ~(1_n234 ^ 1_n1555);
assign 1_n593 = 1_n1226 & 1_n632;
assign 1_n771 = ~1_n1573;
assign 1_n1440 = ~1_n1256;
assign 1_n189 = ~1_n908;
assign 1_n262 = ~1_n1137;
assign 1_n740 = 1_n1668 | 1_n1459;
assign 1_n483 = 1_n855 & 1_n325;
assign 1_n491 = 1_n205 | 1_n862;
assign 1_n586 = ~(1_n765 | 1_n903);
assign 1_n1036 = 1_n563 | 1_n758;
assign 1_n1261 = ~1_n1230;
assign 1_n244 = ~1_n133;
assign 1_n97 = 1_n380 | 1_n1550;
assign 1_n375 = ~(1_n1373 | 1_n530);
assign 1_n1663 = 1_n820 & 1_n1209;
assign 1_n364 = 1_n842;
assign 1_n1548 = ~1_n527;
assign 1_n634 = 1_n1464 | 1_n192;
assign 1_n1480 = ~1_n701;
assign 1_n891 = 1_n354 | 1_n53;
assign 1_n13 = 1_n761 & 1_n1005;
assign 1_n713 = 1_n732 & 1_n1108;
assign 1_n422 = ~(1_n1536 | 1_n1372);
assign 1_n119 = ~(1_n1106 | 1_n1029);
assign 1_n1123 = ~1_n348;
assign 1_n389 = 1_n184 | 1_n1015;
assign 1_n803 = 1_n279 | 1_n985;
assign 1_n1529 = 1_n1219 | 1_n711;
assign 1_n476 = ~1_n1150;
assign 1_n971 = ~1_n1233;
assign 1_n1037 = ~(1_n1388 | 1_n1029);
assign 1_n701 = ~1_n207;
assign 1_n1439 = ~(1_n855 | 1_n161);
assign 1_n381 = 1_n674 | 1_n697;
assign 1_n988 = 1_n1341 | 1_n1163;
assign 1_n718 = ~(1_n1367 | 1_n1670);
assign 1_n1262 = ~1_n889;
assign 1_n201 = 1_n118 & 1_n632;
assign 1_n1487 = ~(1_n290 | 1_n166);
assign 1_n700 = ~1_n230;
assign 1_n437 = 1_n491 | 1_n298;
assign 1_n245 = ~(1_n510 | 1_n178);
endmodule
