// Benchmark "top" written by ABC on Sun Jun 11 02:28:37 2023

module top ( 
    \1_n0 , \1_n21 , \1_n36 , \1_n38 , \1_n45 , \1_n49 , \1_n77 , \1_n95 ,
    \1_n98 , \1_n104 , \1_n107 , \1_n108 , \1_n116 , \1_n122 , \1_n127 ,
    \1_n128 , \1_n138 , \1_n153 , \1_n192 , \1_n196 , \1_n200 , \1_n208 ,
    \1_n221 , \1_n231 , \1_n236 , \1_n244 , \1_n245 , \1_n246 , \1_n252 ,
    \1_n258 , \1_n260 , \1_n262 , \1_n267 , \1_n268 , \1_n281 , \1_n284 ,
    \1_n288 , \1_n301 , \1_n305 , \1_n310 , \1_n319 , \1_n323 , \1_n324 ,
    \1_n332 , \1_n336 , \1_n359 , \1_n360 , \1_n364 , \1_n366 , \1_n381 ,
    \1_n384 , \1_n393 , \1_n398 , \1_n421 , \1_n423 , \1_n431 , \1_n433 ,
    \1_n438 , \1_n439 , \1_n441 , \1_n444 , \1_n448 , \1_n449 , \1_n475 ,
    \1_n491 , \1_n500 , \1_n505 , \1_n507 , \1_n510 , \1_n519 , \1_n532 ,
    \1_n536 , \1_n540 , \1_n571 , \1_n577 , \1_n589 , \1_n599 , \1_n610 ,
    \1_n631 , \1_n635 , \1_n640 , \1_n644 , \1_n650 , \1_n657 , \1_n667 ,
    \1_n685 , \1_n688 , \1_n695 , \1_n714 , \1_n716 , \1_n741 , \1_n745 ,
    \1_n749 , \1_n766 , \1_n767 , \1_n771 , \1_n774 , \1_n787 , \1_n802 ,
    \1_n804 , \1_n806 , \1_n818 , \1_n819 , \1_n823 , \1_n825 , \1_n826 ,
    \1_n833 , \1_n839 , \1_n841 , \1_n845 , \1_n851 , \1_n857 , \1_n862 ,
    \1_n863 , \1_n866 , \1_n870 , \1_n879 , \1_n893 , \1_n896 , \1_n901 ,
    \1_n928 , \1_n929 , \1_n936 , \1_n944 , \1_n952 , \1_n955 , \1_n961 ,
    \1_n975 , \1_n976 , \1_n986 , \1_n997 , \1_n1005 , \1_n1022 ,
    \1_n1029 , \1_n1035 , \1_n1036 , \1_n1041 , \1_n1044 , \1_n1045 ,
    \1_n1048 , \1_n1064 , \1_n1067 , \1_n1069 , \1_n1072 , \1_n1073 ,
    \1_n1077 , \1_n1080 , \1_n1081 , \1_n1089 , \1_n1091 , \1_n1097 ,
    \1_n1098 , \1_n1120 , \1_n1131 , \1_n1132 , \1_n1140 , \1_n1141 ,
    \1_n1143 , \1_n1146 , \1_n1151 , \1_n1163 , \1_n1164 , \1_n1180 ,
    \1_n1191 , \1_n1198 , \1_n1219 , \1_n1226 , \1_n1229 , \1_n1231 ,
    \1_n1236 , \1_n1257 , \1_n1269 , \1_n1273 , \1_n1277 , \1_n1279 ,
    \1_n1298 , \1_n1308 , \1_n1311 , \1_n1321 , \1_n1326 , \1_n1342 ,
    \1_n1344 , \1_n1352 ,
    \1_n29 , \1_n34 , \1_n60 , \1_n81 , \1_n82 , \1_n88 , \1_n90 , \1_n91 ,
    \1_n112 , \1_n129 , \1_n130 , \1_n135 , \1_n150 , \1_n159 , \1_n167 ,
    \1_n168 , \1_n175 , \1_n185 , \1_n190 , \1_n193 , \1_n204 , \1_n206 ,
    \1_n207 , \1_n218 , \1_n223 , \1_n227 , \1_n228 , \1_n229 , \1_n240 ,
    \1_n275 , \1_n299 , \1_n307 , \1_n342 , \1_n347 , \1_n374 , \1_n383 ,
    \1_n389 , \1_n408 , \1_n409 , \1_n410 , \1_n415 , \1_n432 , \1_n452 ,
    \1_n456 , \1_n492 , \1_n516 , \1_n554 , \1_n580 , \1_n592 , \1_n598 ,
    \1_n607 , \1_n608 , \1_n613 , \1_n617 , \1_n621 , \1_n623 , \1_n627 ,
    \1_n638 , \1_n651 , \1_n653 , \1_n662 , \1_n679 , \1_n683 , \1_n707 ,
    \1_n710 , \1_n718 , \1_n723 , \1_n733 , \1_n734 , \1_n747 , \1_n779 ,
    \1_n785 , \1_n801 , \1_n807 , \1_n808 , \1_n817 , \1_n835 , \1_n842 ,
    \1_n853 , \1_n854 , \1_n877 , \1_n905 , \1_n908 , \1_n927 , \1_n962 ,
    \1_n966 , \1_n973 , \1_n999 , \1_n1023 , \1_n1027 , \1_n1057 ,
    \1_n1059 , \1_n1061 , \1_n1085 , \1_n1099 , \1_n1150 , \1_n1153 ,
    \1_n1178 , \1_n1184 , \1_n1194 , \1_n1202 , \1_n1206 , \1_n1232 ,
    \1_n1239 , \1_n1259 , \1_n1264 , \1_n1288 , \1_n1301   );
  input  \1_n0 , \1_n21 , \1_n36 , \1_n38 , \1_n45 , \1_n49 , \1_n77 ,
    \1_n95 , \1_n98 , \1_n104 , \1_n107 , \1_n108 , \1_n116 , \1_n122 ,
    \1_n127 , \1_n128 , \1_n138 , \1_n153 , \1_n192 , \1_n196 , \1_n200 ,
    \1_n208 , \1_n221 , \1_n231 , \1_n236 , \1_n244 , \1_n245 , \1_n246 ,
    \1_n252 , \1_n258 , \1_n260 , \1_n262 , \1_n267 , \1_n268 , \1_n281 ,
    \1_n284 , \1_n288 , \1_n301 , \1_n305 , \1_n310 , \1_n319 , \1_n323 ,
    \1_n324 , \1_n332 , \1_n336 , \1_n359 , \1_n360 , \1_n364 , \1_n366 ,
    \1_n381 , \1_n384 , \1_n393 , \1_n398 , \1_n421 , \1_n423 , \1_n431 ,
    \1_n433 , \1_n438 , \1_n439 , \1_n441 , \1_n444 , \1_n448 , \1_n449 ,
    \1_n475 , \1_n491 , \1_n500 , \1_n505 , \1_n507 , \1_n510 , \1_n519 ,
    \1_n532 , \1_n536 , \1_n540 , \1_n571 , \1_n577 , \1_n589 , \1_n599 ,
    \1_n610 , \1_n631 , \1_n635 , \1_n640 , \1_n644 , \1_n650 , \1_