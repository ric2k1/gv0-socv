module top(in1, in2, in3, out1);
  input [18:0] in1, in2, in3;
  output [19:0] out1;
  wire [18:0] in1, in2, in3;
  wire [19:0] out1;
  wire csa_tree_add_6_33_groupi_n_2, csa_tree_add_6_33_groupi_n_3, csa_tree_add_6_33_groupi_n_4, csa_tree_add_6_33_groupi_n_5, csa_tree_add_6_33_groupi_n_6, csa_tree_add_6_33_groupi_n_7, csa_tree_add_6_33_groupi_n_8, csa_tree_add_6_33_groupi_n_9;
  wire csa_tree_add_6_33_groupi_n_10, csa_tree_add_6_33_groupi_n_11, csa_tree_add_6_33_groupi_n_12, csa_tree_add_6_33_groupi_n_13, csa_tree_add_6_33_groupi_n_14, csa_tree_add_6_33_groupi_n_15, csa_tree_add_6_33_groupi_n_16, csa_tree_add_6_33_groupi_n_17;
  wire csa_tree_add_6_33_groupi_n_18, csa_tree_add_6_33_groupi_n_19, csa_tree_add_6_33_groupi_n_20, csa_tree_add_6_33_groupi_n_21, csa_tree_add_6_33_groupi_n_22, csa_tree_add_6_33_groupi_n_23, csa_tree_add_6_33_groupi_n_24, csa_tree_add_6_33_groupi_n_25;
  wire csa_tree_add_6_33_groupi_n_26, csa_tree_add_6_33_groupi_n_27, csa_tree_add_6_33_groupi_n_28, csa_tree_add_6_33_groupi_n_29, csa_tree_add_6_33_groupi_n_30, csa_tree_add_6_33_groupi_n_31, csa_tree_add_6_33_groupi_n_32, csa_tree_add_6_33_groupi_n_33;
  wire csa_tree_add_6_33_groupi_n_34, csa_tree_add_6_33_groupi_n_35, csa_tree_add_6_33_groupi_n_36, csa_tree_add_6_33_groupi_n_37, csa_tree_add_6_33_groupi_n_38, csa_tree_add_6_33_groupi_n_39, csa_tree_add_6_33_groupi_n_40, csa_tree_add_6_33_groupi_n_41;
  wire csa_tree_add_6_33_groupi_n_42, csa_tree_add_6_33_groupi_n_43, csa_tree_add_6_33_groupi_n_44, csa_tree_add_6_33_groupi_n_45, csa_tree_add_6_33_groupi_n_46, csa_tree_add_6_33_groupi_n_47, csa_tree_add_6_33_groupi_n_48, csa_tree_add_6_33_groupi_n_49;
  wire csa_tree_add_6_33_groupi_n_50, csa_tree_add_6_33_groupi_n_51, csa_tree_add_6_33_groupi_n_52, csa_tree_add_6_33_groupi_n_53, csa_tree_add_6_33_groupi_n_54, csa_tree_add_6_33_groupi_n_55, csa_tree_add_6_33_groupi_n_56, csa_tree_add_6_33_groupi_n_57;
  wire csa_tree_add_6_33_groupi_n_58, csa_tree_add_6_33_groupi_n_59, csa_tree_add_6_33_groupi_n_60, csa_tree_add_6_33_groupi_n_61, csa_tree_add_6_33_groupi_n_62, csa_tree_add_6_33_groupi_n_63, csa_tree_add_6_33_groupi_n_64, csa_tree_add_6_33_groupi_n_65;
  wire csa_tree_add_6_33_groupi_n_66, csa_tree_add_6_33_groupi_n_67, csa_tree_add_6_33_groupi_n_68, csa_tree_add_6_33_groupi_n_69, csa_tree_add_6_33_groupi_n_70, csa_tree_add_6_33_groupi_n_71, csa_tree_add_6_33_groupi_n_72, csa_tree_add_6_33_groupi_n_73;
  wire csa_tree_add_6_33_groupi_n_74, csa_tree_add_6_33_groupi_n_75, csa_tree_add_6_33_groupi_n_76, csa_tree_add_6_33_groupi_n_77, csa_tree_add_6_33_groupi_n_78, csa_tree_add_6_33_groupi_n_79, csa_tree_add_6_33_groupi_n_80, csa_tree_add_6_33_groupi_n_81;
  wire csa_tree_add_6_33_groupi_n_82, csa_tree_add_6_33_groupi_n_83, csa_tree_add_6_33_groupi_n_84, csa_tree_add_6_33_groupi_n_85, csa_tree_add_6_33_groupi_n_86, csa_tree_add_6_33_groupi_n_87, csa_tree_add_6_33_groupi_n_88, csa_tree_add_6_33_groupi_n_89;
  wire csa_tree_add_6_33_groupi_n_90, csa_tree_add_6_33_groupi_n_91, csa_tree_add_6_33_groupi_n_92, csa_tree_add_6_33_groupi_n_93, csa_tree_add_6_33_groupi_n_94, csa_tree_add_6_33_groupi_n_95, csa_tree_add_6_33_groupi_n_96, csa_tree_add_6_33_groupi_n_97;
  wire csa_tree_add_6_33_groupi_n_98, csa_tree_add_6_33_groupi_n_99, csa_tree_add_6_33_groupi_n_100, csa_tree_add_6_33_groupi_n_101, csa_tree_add_6_33_groupi_n_102, csa_tree_add_6_33_groupi_n_103, csa_tree_add_6_33_groupi_n_104, csa_tree_add_6_33_groupi_n_105;
  wire csa_tree_add_6_33_groupi_n_106, csa_tree_add_6_33_groupi_n_107, csa_tree_add_6_33_groupi_n_108, csa_tree_add_6_33_groupi_n_109, csa_tree_add_6_33_groupi_n_110, csa_tree_add_6_33_groupi_n_111, csa_tree_add_6_33_groupi_n_112, csa_tree_add_6_33_groupi_n_113;
  wire csa_tree_add_6_33_groupi_n_114, csa_tree_add_6_33_groupi_n_115, csa_tree_add_6_33_groupi_n_116, csa_tree_add_6_33_groupi_n_117, csa_tree_add_6_33_groupi_n_118, csa_tree_add_6_33_groupi_n_119, csa_tree_add_6_33_groupi_n_120, csa_tree_add_6_33_groupi_n_121;
  wire csa_tree_add_6_33_groupi_n_122, csa_tree_add_6_33_groupi_n_123, csa_tree_add_6_33_groupi_n_124, csa_tree_add_6_33_groupi_n_125, csa_tree_add_6_33_groupi_n_126, csa_tree_add_6_33_groupi_n_127, csa_tree_add_6_33_groupi_n_128, csa_tree_add_6_33_groupi_n_129;
  wire csa_tree_add_6_33_groupi_n_130, csa_tree_add_6_33_groupi_n_131, csa_tree_add_6_33_groupi_n_132, csa_tree_add_6_33_groupi_n_133, csa_tree_add_6_33_groupi_n_134, csa_tree_add_6_33_groupi_n_135, csa_tree_add_6_33_groupi_n_136, csa_tree_add_6_33_groupi_n_137;
  wire csa_tree_add_6_33_groupi_n_138, csa_tree_add_6_33_groupi_n_139, csa_tree_add_6_33_groupi_n_140, csa_tree_add_6_33_groupi_n_141, csa_tree_add_6_33_groupi_n_142, csa_tree_add_6_33_groupi_n_143, csa_tree_add_6_33_groupi_n_144, csa_tree_add_6_33_groupi_n_145;
  wire csa_tree_add_6_33_groupi_n_146, csa_tree_add_6_33_groupi_n_147, csa_tree_add_6_33_groupi_n_148, csa_tree_add_6_33_groupi_n_149, csa_tree_add_6_33_groupi_n_150, csa_tree_add_6_33_groupi_n_151, csa_tree_add_6_33_groupi_n_152, csa_tree_add_6_33_groupi_n_153;
  wire csa_tree_add_6_33_groupi_n_154, csa_tree_add_6_33_groupi_n_155, csa_tree_add_6_33_groupi_n_156, csa_tree_add_6_33_groupi_n_157, csa_tree_add_6_33_groupi_n_158, csa_tree_add_6_33_groupi_n_159, csa_tree_add_6_33_groupi_n_160, csa_tree_add_6_33_groupi_n_161;
  wire csa_tree_add_6_33_groupi_n_162, csa_tree_add_6_33_groupi_n_163, csa_tree_add_6_33_groupi_n_165, csa_tree_add_6_33_groupi_n_166, csa_tree_add_6_33_groupi_n_167, csa_tree_add_6_33_groupi_n_168, csa_tree_add_6_33_groupi_n_169, csa_tree_add_6_33_groupi_n_170;
  wire csa_tree_add_6_33_groupi_n_171, csa_tree_add_6_33_groupi_n_172, csa_tree_add_6_33_groupi_n_173, csa_tree_add_6_33_groupi_n_174, csa_tree_add_6_33_groupi_n_175, csa_tree_add_6_33_groupi_n_176, csa_tree_add_6_33_groupi_n_177, csa_tree_add_6_33_groupi_n_178;
  wire csa_tree_add_6_33_groupi_n_179, csa_tree_add_6_33_groupi_n_180, csa_tree_add_6_33_groupi_n_181, csa_tree_add_6_33_groupi_n_182, csa_tree_add_6_33_groupi_n_183, csa_tree_add_6_33_groupi_n_184, csa_tree_add_6_33_groupi_n_185, csa_tree_add_6_33_groupi_n_186;
  wire csa_tree_add_6_33_groupi_n_187, csa_tree_add_6_33_groupi_n_188, csa_tree_add_6_33_groupi_n_189, csa_tree_add_6_33_groupi_n_190, csa_tree_add_6_33_groupi_n_191, csa_tree_add_6_33_groupi_n_192, csa_tree_add_6_33_groupi_n_193, csa_tree_add_6_33_groupi_n_194;
  wire csa_tree_add_6_33_groupi_n_195, csa_tree_add_6_33_groupi_n_196, csa_tree_add_6_33_groupi_n_198, csa_tree_add_6_33_groupi_n_199, csa_tree_add_6_33_groupi_n_200, csa_tree_add_6_33_groupi_n_201, csa_tree_add_6_33_groupi_n_202, csa_tree_add_6_33_groupi_n_203;
  wire csa_tree_add_6_33_groupi_n_204, csa_tree_add_6_33_groupi_n_205, csa_tree_add_6_33_groupi_n_206, csa_tree_add_6_33_groupi_n_207, csa_tree_add_6_33_groupi_n_208, csa_tree_add_6_33_groupi_n_209, csa_tree_add_6_33_groupi_n_210, csa_tree_add_6_33_groupi_n_211;
  wire csa_tree_add_6_33_groupi_n_212, csa_tree_add_6_33_groupi_n_213, csa_tree_add_6_33_groupi_n_214, csa_tree_add_6_33_groupi_n_215, csa_tree_add_6_33_groupi_n_216, csa_tree_add_6_33_groupi_n_217, csa_tree_add_6_33_groupi_n_218, csa_tree_add_6_33_groupi_n_219;
  wire csa_tree_add_6_33_groupi_n_220, csa_tree_add_6_33_groupi_n_221, csa_tree_add_6_33_groupi_n_222, csa_tree_add_6_33_groupi_n_223, csa_tree_add_6_33_groupi_n_224, csa_tree_add_6_33_groupi_n_225, csa_tree_add_6_33_groupi_n_226, csa_tree_add_6_33_groupi_n_227;
  wire csa_tree_add_6_33_groupi_n_228, csa_tree_add_6_33_groupi_n_229, csa_tree_add_6_33_groupi_n_230, csa_tree_add_6_33_groupi_n_231, csa_tree_add_6_33_groupi_n_232, csa_tree_add_6_33_groupi_n_233, csa_tree_add_6_33_groupi_n_234, csa_tree_add_6_33_groupi_n_235;
  wire csa_tree_add_6_33_groupi_n_236, csa_tree_add_6_33_groupi_n_237, csa_tree_add_6_33_groupi_n_238, csa_tree_add_6_33_groupi_n_239, csa_tree_add_6_33_groupi_n_240, csa_tree_add_6_33_groupi_n_241, csa_tree_add_6_33_groupi_n_242, csa_tree_add_6_33_groupi_n_243;
  wire csa_tree_add_6_33_groupi_n_244, csa_tree_add_6_33_groupi_n_245, csa_tree_add_6_33_groupi_n_246, csa_tree_add_6_33_groupi_n_247, csa_tree_add_6_33_groupi_n_248, csa_tree_add_6_33_groupi_n_249, csa_tree_add_6_33_groupi_n_250, csa_tree_add_6_33_groupi_n_251;
  wire csa_tree_add_6_33_groupi_n_252, csa_tree_add_6_33_groupi_n_253, csa_tree_add_6_33_groupi_n_254, csa_tree_add_6_33_groupi_n_255, csa_tree_add_6_33_groupi_n_256, csa_tree_add_6_33_groupi_n_257, csa_tree_add_6_33_groupi_n_258, csa_tree_add_6_33_groupi_n_259;
  wire csa_tree_add_6_33_groupi_n_260, csa_tree_add_6_33_groupi_n_261, csa_tree_add_6_33_groupi_n_262, csa_tree_add_6_33_groupi_n_263, csa_tree_add_6_33_groupi_n_264, csa_tree_add_6_33_groupi_n_265, csa_tree_add_6_33_groupi_n_267, csa_tree_add_6_33_groupi_n_269;
  wire csa_tree_add_6_33_groupi_n_270, csa_tree_add_6_33_groupi_n_271, csa_tree_add_6_33_groupi_n_272, csa_tree_add_6_33_groupi_n_273, csa_tree_add_6_33_groupi_n_275, csa_tree_add_6_33_groupi_n_276, csa_tree_add_6_33_groupi_n_278, csa_tree_add_6_33_groupi_n_279;
  wire csa_tree_add_6_33_groupi_n_281, csa_tree_add_6_33_groupi_n_282, csa_tree_add_6_33_groupi_n_284, csa_tree_add_6_33_groupi_n_285, csa_tree_add_6_33_groupi_n_287, csa_tree_add_6_33_groupi_n_288, csa_tree_add_6_33_groupi_n_290, csa_tree_add_6_33_groupi_n_291;
  wire csa_tree_add_6_33_groupi_n_293, csa_tree_add_6_33_groupi_n_294, csa_tree_add_6_33_groupi_n_296, csa_tree_add_6_33_groupi_n_297, csa_tree_add_6_33_groupi_n_299, csa_tree_add_6_33_groupi_n_300, csa_tree_add_6_33_groupi_n_302, csa_tree_add_6_33_groupi_n_303;
  wire csa_tree_add_6_33_groupi_n_305, csa_tree_add_6_33_groupi_n_306, csa_tree_add_6_33_groupi_n_308, csa_tree_add_6_33_groupi_n_309, csa_tree_add_6_33_groupi_n_311;
  xnor csa_tree_add_6_33_groupi_g862__2398(out1[19] ,csa_tree_add_6_33_groupi_n_219 ,csa_tree_add_6_33_groupi_n_311);
  or csa_tree_add_6_33_groupi_g863__5107(csa_tree_add_6_33_groupi_n_311 ,csa_tree_add_6_33_groupi_n_245 ,csa_tree_add_6_33_groupi_n_309);
  xnor csa_tree_add_6_33_groupi_g864__6260(out1[18] ,csa_tree_add_6_33_groupi_n_308 ,csa_tree_add_6_33_groupi_n_263);
  and csa_tree_add_6_33_groupi_g865__4319(csa_tree_add_6_33_groupi_n_309 ,csa_tree_add_6_33_groupi_n_241 ,csa_tree_add_6_33_groupi_n_308);
  or csa_tree_add_6_33_groupi_g866__8428(csa_tree_add_6_33_groupi_n_308 ,csa_tree_add_6_33_groupi_n_237 ,csa_tree_add_6_33_groupi_n_306);
  xnor csa_tree_add_6_33_groupi_g867__5526(out1[17] ,csa_tree_add_6_33_groupi_n_305 ,csa_tree_add_6_33_groupi_n_264);
  and csa_tree_add_6_33_groupi_g868__6783(csa_tree_add_6_33_groupi_n_306 ,csa_tree_add_6_33_groupi_n_228 ,csa_tree_add_6_33_groupi_n_305);
  or csa_tree_add_6_33_groupi_g869__3680(csa_tree_add_6_33_groupi_n_305 ,csa_tree_add_6_33_groupi_n_227 ,csa_tree_add_6_33_groupi_n_303);
  xnor csa_tree_add_6_33_groupi_g870__1617(out1[16] ,csa_tree_add_6_33_groupi_n_302 ,csa_tree_add_6_33_groupi_n_261);
  and csa_tree_add_6_33_groupi_g871__2802(csa_tree_add_6_33_groupi_n_303 ,csa_tree_add_6_33_groupi_n_244 ,csa_tree_add_6_33_groupi_n_302);
  or csa_tree_add_6_33_groupi_g872__1705(csa_tree_add_6_33_groupi_n_302 ,csa_tree_add_6_33_groupi_n_240 ,csa_tree_add_6_33_groupi_n_300);
  xnor csa_tree_add_6_33_groupi_g873__5122(out1[15] ,csa_tree_add_6_33_groupi_n_299 ,csa_tree_add_6_33_groupi_n_260);
  and csa_tree_add_6_33_groupi_g874__8246(csa_tree_add_6_33_groupi_n_300 ,csa_tree_add_6_33_groupi_n_233 ,csa_tree_add_6_33_groupi_n_299);
  or csa_tree_add_6_33_groupi_g875__7098(csa_tree_add_6_33_groupi_n_299 ,csa_tree_add_6_33_groupi_n_232 ,csa_tree_add_6_33_groupi_n_297);
  xnor csa_tree_add_6_33_groupi_g876__6131(out1[14] ,csa_tree_add_6_33_groupi_n_296 ,csa_tree_add_6_33_groupi_n_259);
  and csa_tree_add_6_33_groupi_g877__1881(csa_tree_add_6_33_groupi_n_297 ,csa_tree_add_6_33_groupi_n_225 ,csa_tree_add_6_33_groupi_n_296);
  or csa_tree_add_6_33_groupi_g878__5115(csa_tree_add_6_33_groupi_n_296 ,csa_tree_add_6_33_groupi_n_224 ,csa_tree_add_6_33_groupi_n_294);
  xnor csa_tree_add_6_33_groupi_g879__7482(out1[13] ,csa_tree_add_6_33_groupi_n_293 ,csa_tree_add_6_33_groupi_n_254);
  and csa_tree_add_6_33_groupi_g880__4733(csa_tree_add_6_33_groupi_n_294 ,csa_tree_add_6_33_groupi_n_248 ,csa_tree_add_6_33_groupi_n_293);
  or csa_tree_add_6_33_groupi_g881__6161(csa_tree_add_6_33_groupi_n_293 ,csa_tree_add_6_33_groupi_n_247 ,csa_tree_add_6_33_groupi_n_291);
  xnor csa_tree_add_6_33_groupi_g882__9315(out1[12] ,csa_tree_add_6_33_groupi_n_290 ,csa_tree_add_6_33_groupi_n_257);
  and csa_tree_add_6_33_groupi_g883__9945(csa_tree_add_6_33_groupi_n_291 ,csa_tree_add_6_33_groupi_n_243 ,csa_tree_add_6_33_groupi_n_290);
  or csa_tree_add_6_33_groupi_g884__2883(csa_tree_add_6_33_groupi_n_290 ,csa_tree_add_6_33_groupi_n_239 ,csa_tree_add_6_33_groupi_n_288);
  xnor csa_tree_add_6_33_groupi_g885__2346(out1[11] ,csa_tree_add_6_33_groupi_n_287 ,csa_tree_add_6_33_groupi_n_256);
  and csa_tree_add_6_33_groupi_g886__1666(csa_tree_add_6_33_groupi_n_288 ,csa_tree_add_6_33_groupi_n_234 ,csa_tree_add_6_33_groupi_n_287);
  or csa_tree_add_6_33_groupi_g887__7410(csa_tree_add_6_33_groupi_n_287 ,csa_tree_add_6_33_groupi_n_222 ,csa_tree_add_6_33_groupi_n_285);
  xnor csa_tree_add_6_33_groupi_g888__6417(out1[10] ,csa_tree_add_6_33_groupi_n_284 ,csa_tree_add_6_33_groupi_n_255);
  and csa_tree_add_6_33_groupi_g889__5477(csa_tree_add_6_33_groupi_n_285 ,csa_tree_add_6_33_groupi_n_231 ,csa_tree_add_6_33_groupi_n_284);
  or csa_tree_add_6_33_groupi_g890__2398(csa_tree_add_6_33_groupi_n_284 ,csa_tree_add_6_33_groupi_n_230 ,csa_tree_add_6_33_groupi_n_282);
  xnor csa_tree_add_6_33_groupi_g891__5107(out1[9] ,csa_tree_add_6_33_groupi_n_281 ,csa_tree_add_6_33_groupi_n_258);
  and csa_tree_add_6_33_groupi_g892__6260(csa_tree_add_6_33_groupi_n_282 ,csa_tree_add_6_33_groupi_n_242 ,csa_tree_add_6_33_groupi_n_281);
  or csa_tree_add_6_33_groupi_g893__4319(csa_tree_add_6_33_groupi_n_281 ,csa_tree_add_6_33_groupi_n_229 ,csa_tree_add_6_33_groupi_n_279);
  xnor csa_tree_add_6_33_groupi_g894__8428(out1[8] ,csa_tree_add_6_33_groupi_n_278 ,csa_tree_add_6_33_groupi_n_253);
  and csa_tree_add_6_33_groupi_g895__5526(csa_tree_add_6_33_groupi_n_279 ,csa_tree_add_6_33_groupi_n_226 ,csa_tree_add_6_33_groupi_n_278);
  or csa_tree_add_6_33_groupi_g896__6783(csa_tree_add_6_33_groupi_n_278 ,csa_tree_add_6_33_groupi_n_223 ,csa_tree_add_6_33_groupi_n_276);
  xnor csa_tree_add_6_33_groupi_g897__3680(out1[7] ,csa_tree_add_6_33_groupi_n_275 ,csa_tree_add_6_33_groupi_n_252);
  and csa_tree_add_6_33_groupi_g898__1617(csa_tree_add_6_33_groupi_n_276 ,csa_tree_add_6_33_groupi_n_235 ,csa_tree_add_6_33_groupi_n_275);
  or csa_tree_add_6_33_groupi_g899__2802(csa_tree_add_6_33_groupi_n_275 ,csa_tree_add_6_33_groupi_n_213 ,csa_tree_add_6_33_groupi_n_273);
  xnor csa_tree_add_6_33_groupi_g900__1705(out1[6] ,csa_tree_add_6_33_groupi_n_272 ,csa_tree_add_6_33_groupi_n_221);
  nor csa_tree_add_6_33_groupi_g901__5122(csa_tree_add_6_33_groupi_n_273 ,csa_tree_add_6_33_groupi_n_212 ,csa_tree_add_6_33_groupi_n_272);
  and csa_tree_add_6_33_groupi_g902__8246(csa_tree_add_6_33_groupi_n_272 ,csa_tree_add_6_33_groupi_n_211 ,csa_tree_add_6_33_groupi_n_271);
  or csa_tree_add_6_33_groupi_g904__7098(csa_tree_add_6_33_groupi_n_271 ,csa_tree_add_6_33_groupi_n_210 ,csa_tree_add_6_33_groupi_n_270);
  and csa_tree_add_6_33_groupi_g906__6131(csa_tree_add_6_33_groupi_n_270 ,csa_tree_add_6_33_groupi_n_246 ,csa_tree_add_6_33_groupi_n_269);
  or csa_tree_add_6_33_groupi_g908__1881(csa_tree_add_6_33_groupi_n_269 ,csa_tree_add_6_33_groupi_n_249 ,csa_tree_add_6_33_groupi_n_267);
  xnor csa_tree_add_6_33_groupi_g909__5115(out1[3] ,csa_tree_add_6_33_groupi_n_250 ,csa_tree_add_6_33_groupi_n_262);
  and csa_tree_add_6_33_groupi_g911__7482(csa_tree_add_6_33_groupi_n_267 ,csa_tree_add_6_33_groupi_n_238 ,csa_tree_add_6_33_groupi_n_265);
  xnor csa_tree_add_6_33_groupi_g912__4733(out1[2] ,csa_tree_add_6_33_groupi_n_191 ,csa_tree_add_6_33_groupi_n_196);
  or csa_tree_add_6_33_groupi_g913__6161(csa_tree_add_6_33_groupi_n_265 ,csa_tree_add_6_33_groupi_n_236 ,csa_tree_add_6_33_groupi_n_250);
  xnor csa_tree_add_6_33_groupi_g914__9315(csa_tree_add_6_33_groupi_n_264 ,csa_tree_add_6_33_groupi_n_182 ,csa_tree_add_6_33_groupi_n_206);
  xnor csa_tree_add_6_33_groupi_g915__9945(csa_tree_add_6_33_groupi_n_263 ,csa_tree_add_6_33_groupi_n_181 ,csa_tree_add_6_33_groupi_n_214);
  xnor csa_tree_add_6_33_groupi_g916__2883(csa_tree_add_6_33_groupi_n_262 ,csa_tree_add_6_33_groupi_n_199 ,csa_tree_add_6_33_groupi_n_148);
  xnor csa_tree_add_6_33_groupi_g917__2346(csa_tree_add_6_33_groupi_n_261 ,csa_tree_add_6_33_groupi_n_180 ,csa_tree_add_6_33_groupi_n_218);
  xnor csa_tree_add_6_33_groupi_g918__1666(csa_tree_add_6_33_groupi_n_260 ,csa_tree_add_6_33_groupi_n_183 ,csa_tree_add_6_33_groupi_n_201);
  xnor csa_tree_add_6_33_groupi_g919__7410(csa_tree_add_6_33_groupi_n_259 ,csa_tree_add_6_33_groupi_n_176 ,csa_tree_add_6_33_groupi_n_202);
  xnor csa_tree_add_6_33_groupi_g920__6417(csa_tree_add_6_33_groupi_n_258 ,csa_tree_add_6_33_groupi_n_189 ,csa_tree_add_6_33_groupi_n_203);
  xnor csa_tree_add_6_33_groupi_g921__5477(csa_tree_add_6_33_groupi_n_257 ,csa_tree_add_6_33_groupi_n_175 ,csa_tree_add_6_33_groupi_n_215);
  xnor csa_tree_add_6_33_groupi_g922__2398(csa_tree_add_6_33_groupi_n_256 ,csa_tree_add_6_33_groupi_n_184 ,csa_tree_add_6_33_groupi_n_208);
  xnor csa_tree_add_6_33_groupi_g923__5107(csa_tree_add_6_33_groupi_n_255 ,csa_tree_add_6_33_groupi_n_190 ,csa_tree_add_6_33_groupi_n_207);
  xnor csa_tree_add_6_33_groupi_g924__6260(csa_tree_add_6_33_groupi_n_254 ,csa_tree_add_6_33_groupi_n_172 ,csa_tree_add_6_33_groupi_n_217);
  xnor csa_tree_add_6_33_groupi_g925__4319(csa_tree_add_6_33_groupi_n_253 ,csa_tree_add_6_33_groupi_n_188 ,csa_tree_add_6_33_groupi_n_200);
  xnor csa_tree_add_6_33_groupi_g926__8428(csa_tree_add_6_33_groupi_n_252 ,csa_tree_add_6_33_groupi_n_187 ,csa_tree_add_6_33_groupi_n_216);
  xnor csa_tree_add_6_33_groupi_g927__5526(csa_tree_add_6_33_groupi_n_251 ,csa_tree_add_6_33_groupi_n_174 ,csa_tree_add_6_33_groupi_n_205);
  nor csa_tree_add_6_33_groupi_g928__6783(csa_tree_add_6_33_groupi_n_249 ,csa_tree_add_6_33_groupi_n_174 ,csa_tree_add_6_33_groupi_n_205);
  or csa_tree_add_6_33_groupi_g929__3680(csa_tree_add_6_33_groupi_n_248 ,csa_tree_add_6_33_groupi_n_172 ,csa_tree_add_6_33_groupi_n_217);
  and csa_tree_add_6_33_groupi_g930__1617(csa_tree_add_6_33_groupi_n_247 ,csa_tree_add_6_33_groupi_n_175 ,csa_tree_add_6_33_groupi_n_215);
  or csa_tree_add_6_33_groupi_g931__2802(csa_tree_add_6_33_groupi_n_246 ,csa_tree_add_6_33_groupi_n_173 ,csa_tree_add_6_33_groupi_n_204);
  and csa_tree_add_6_33_groupi_g932__1705(csa_tree_add_6_33_groupi_n_245 ,csa_tree_add_6_33_groupi_n_181 ,csa_tree_add_6_33_groupi_n_214);
  or csa_tree_add_6_33_groupi_g933__5122(csa_tree_add_6_33_groupi_n_244 ,csa_tree_add_6_33_groupi_n_180 ,csa_tree_add_6_33_groupi_n_218);
  or csa_tree_add_6_33_groupi_g934__8246(csa_tree_add_6_33_groupi_n_243 ,csa_tree_add_6_33_groupi_n_175 ,csa_tree_add_6_33_groupi_n_215);
  or csa_tree_add_6_33_groupi_g935__7098(csa_tree_add_6_33_groupi_n_242 ,csa_tree_add_6_33_groupi_n_189 ,csa_tree_add_6_33_groupi_n_203);
  or csa_tree_add_6_33_groupi_g936__6131(csa_tree_add_6_33_groupi_n_241 ,csa_tree_add_6_33_groupi_n_181 ,csa_tree_add_6_33_groupi_n_214);
  and csa_tree_add_6_33_groupi_g937__1881(csa_tree_add_6_33_groupi_n_240 ,csa_tree_add_6_33_groupi_n_183 ,csa_tree_add_6_33_groupi_n_201);
  and csa_tree_add_6_33_groupi_g938__5115(csa_tree_add_6_33_groupi_n_239 ,csa_tree_add_6_33_groupi_n_184 ,csa_tree_add_6_33_groupi_n_208);
  or csa_tree_add_6_33_groupi_g939__7482(csa_tree_add_6_33_groupi_n_238 ,csa_tree_add_6_33_groupi_n_148 ,csa_tree_add_6_33_groupi_n_198);
  and csa_tree_add_6_33_groupi_g940__4733(csa_tree_add_6_33_groupi_n_237 ,csa_tree_add_6_33_groupi_n_182 ,csa_tree_add_6_33_groupi_n_206);
  nor csa_tree_add_6_33_groupi_g941__6161(csa_tree_add_6_33_groupi_n_236 ,csa_tree_add_6_33_groupi_n_147 ,csa_tree_add_6_33_groupi_n_199);
  or csa_tree_add_6_33_groupi_g942__9315(csa_tree_add_6_33_groupi_n_235 ,csa_tree_add_6_33_groupi_n_187 ,csa_tree_add_6_33_groupi_n_216);
  and csa_tree_add_6_33_groupi_g943__9945(csa_tree_add_6_33_groupi_n_250 ,csa_tree_add_6_33_groupi_n_194 ,csa_tree_add_6_33_groupi_n_209);
  or csa_tree_add_6_33_groupi_g944__2883(csa_tree_add_6_33_groupi_n_234 ,csa_tree_add_6_33_groupi_n_184 ,csa_tree_add_6_33_groupi_n_208);
  or csa_tree_add_6_33_groupi_g945__2346(csa_tree_add_6_33_groupi_n_233 ,csa_tree_add_6_33_groupi_n_183 ,csa_tree_add_6_33_groupi_n_201);
  and csa_tree_add_6_33_groupi_g946__1666(csa_tree_add_6_33_groupi_n_232 ,csa_tree_add_6_33_groupi_n_176 ,csa_tree_add_6_33_groupi_n_202);
  or csa_tree_add_6_33_groupi_g947__7410(csa_tree_add_6_33_groupi_n_231 ,csa_tree_add_6_33_groupi_n_190 ,csa_tree_add_6_33_groupi_n_207);
  and csa_tree_add_6_33_groupi_g948__6417(csa_tree_add_6_33_groupi_n_230 ,csa_tree_add_6_33_groupi_n_189 ,csa_tree_add_6_33_groupi_n_203);
  and csa_tree_add_6_33_groupi_g949__5477(csa_tree_add_6_33_groupi_n_229 ,csa_tree_add_6_33_groupi_n_188 ,csa_tree_add_6_33_groupi_n_200);
  or csa_tree_add_6_33_groupi_g950__2398(csa_tree_add_6_33_groupi_n_228 ,csa_tree_add_6_33_groupi_n_182 ,csa_tree_add_6_33_groupi_n_206);
  and csa_tree_add_6_33_groupi_g951__5107(csa_tree_add_6_33_groupi_n_227 ,csa_tree_add_6_33_groupi_n_180 ,csa_tree_add_6_33_groupi_n_218);
  or csa_tree_add_6_33_groupi_g952__6260(csa_tree_add_6_33_groupi_n_226 ,csa_tree_add_6_33_groupi_n_188 ,csa_tree_add_6_33_groupi_n_200);
  or csa_tree_add_6_33_groupi_g953__4319(csa_tree_add_6_33_groupi_n_225 ,csa_tree_add_6_33_groupi_n_176 ,csa_tree_add_6_33_groupi_n_202);
  and csa_tree_add_6_33_groupi_g954__8428(csa_tree_add_6_33_groupi_n_224 ,csa_tree_add_6_33_groupi_n_172 ,csa_tree_add_6_33_groupi_n_217);
  and csa_tree_add_6_33_groupi_g955__5526(csa_tree_add_6_33_groupi_n_223 ,csa_tree_add_6_33_groupi_n_187 ,csa_tree_add_6_33_groupi_n_216);
  and csa_tree_add_6_33_groupi_g956__6783(csa_tree_add_6_33_groupi_n_222 ,csa_tree_add_6_33_groupi_n_190 ,csa_tree_add_6_33_groupi_n_207);
  xnor csa_tree_add_6_33_groupi_g957__3680(csa_tree_add_6_33_groupi_n_221 ,csa_tree_add_6_33_groupi_n_178 ,csa_tree_add_6_33_groupi_n_186);
  xnor csa_tree_add_6_33_groupi_g958__1617(csa_tree_add_6_33_groupi_n_220 ,csa_tree_add_6_33_groupi_n_185 ,csa_tree_add_6_33_groupi_n_177);
  xnor csa_tree_add_6_33_groupi_g959__2802(csa_tree_add_6_33_groupi_n_219 ,csa_tree_add_6_33_groupi_n_65 ,csa_tree_add_6_33_groupi_n_195);
  nor csa_tree_add_6_33_groupi_g960__1705(csa_tree_add_6_33_groupi_n_213 ,csa_tree_add_6_33_groupi_n_179 ,csa_tree_add_6_33_groupi_n_186);
  and csa_tree_add_6_33_groupi_g961__5122(csa_tree_add_6_33_groupi_n_212 ,csa_tree_add_6_33_groupi_n_179 ,csa_tree_add_6_33_groupi_n_186);
  or csa_tree_add_6_33_groupi_g962__8246(csa_tree_add_6_33_groupi_n_211 ,csa_tree_add_6_33_groupi_n_177 ,csa_tree_add_6_33_groupi_n_185);
  and csa_tree_add_6_33_groupi_g963__7098(csa_tree_add_6_33_groupi_n_210 ,csa_tree_add_6_33_groupi_n_177 ,csa_tree_add_6_33_groupi_n_185);
  or csa_tree_add_6_33_groupi_g964__6131(csa_tree_add_6_33_groupi_n_209 ,csa_tree_add_6_33_groupi_n_193 ,csa_tree_add_6_33_groupi_n_192);
  xnor csa_tree_add_6_33_groupi_g965__1881(csa_tree_add_6_33_groupi_n_218 ,csa_tree_add_6_33_groupi_n_69 ,csa_tree_add_6_33_groupi_n_161);
  xnor csa_tree_add_6_33_groupi_g966__5115(csa_tree_add_6_33_groupi_n_217 ,csa_tree_add_6_33_groupi_n_58 ,csa_tree_add_6_33_groupi_n_163);
  xnor csa_tree_add_6_33_groupi_g967__7482(csa_tree_add_6_33_groupi_n_216 ,csa_tree_add_6_33_groupi_n_64 ,csa_tree_add_6_33_groupi_n_149);
  xnor csa_tree_add_6_33_groupi_g968__4733(csa_tree_add_6_33_groupi_n_215 ,csa_tree_add_6_33_groupi_n_57 ,csa_tree_add_6_33_groupi_n_160);
  xnor csa_tree_add_6_33_groupi_g969__6161(csa_tree_add_6_33_groupi_n_214 ,csa_tree_add_6_33_groupi_n_63 ,csa_tree_add_6_33_groupi_n_162);
  not csa_tree_add_6_33_groupi_g970(csa_tree_add_6_33_groupi_n_204 ,csa_tree_add_6_33_groupi_n_205);
  not csa_tree_add_6_33_groupi_g971(csa_tree_add_6_33_groupi_n_198 ,csa_tree_add_6_33_groupi_n_199);
  xnor csa_tree_add_6_33_groupi_g972__9315(out1[1] ,csa_tree_add_6_33_groupi_n_133 ,csa_tree_add_6_33_groupi_n_152);
  xnor csa_tree_add_6_33_groupi_g973__9945(csa_tree_add_6_33_groupi_n_196 ,csa_tree_add_6_33_groupi_n_165 ,csa_tree_add_6_33_groupi_n_56);
  xnor csa_tree_add_6_33_groupi_g974__2883(csa_tree_add_6_33_groupi_n_208 ,csa_tree_add_6_33_groupi_n_67 ,csa_tree_add_6_33_groupi_n_157);
  xnor csa_tree_add_6_33_groupi_g975__2346(csa_tree_add_6_33_groupi_n_207 ,csa_tree_add_6_33_groupi_n_68 ,csa_tree_add_6_33_groupi_n_154);
  xnor csa_tree_add_6_33_groupi_g976__1666(csa_tree_add_6_33_groupi_n_206 ,csa_tree_add_6_33_groupi_n_59 ,csa_tree_add_6_33_groupi_n_150);
  xnor csa_tree_add_6_33_groupi_g977__7410(csa_tree_add_6_33_groupi_n_205 ,csa_tree_add_6_33_groupi_n_71 ,csa_tree_add_6_33_groupi_n_159);
  xnor csa_tree_add_6_33_groupi_g978__6417(csa_tree_add_6_33_groupi_n_203 ,csa_tree_add_6_33_groupi_n_62 ,csa_tree_add_6_33_groupi_n_155);
  xnor csa_tree_add_6_33_groupi_g979__5477(csa_tree_add_6_33_groupi_n_202 ,csa_tree_add_6_33_groupi_n_60 ,csa_tree_add_6_33_groupi_n_156);
  xnor csa_tree_add_6_33_groupi_g980__2398(csa_tree_add_6_33_groupi_n_201 ,csa_tree_add_6_33_groupi_n_74 ,csa_tree_add_6_33_groupi_n_153);
  xnor csa_tree_add_6_33_groupi_g981__5107(csa_tree_add_6_33_groupi_n_200 ,csa_tree_add_6_33_groupi_n_76 ,csa_tree_add_6_33_groupi_n_151);
  xnor csa_tree_add_6_33_groupi_g982__6260(csa_tree_add_6_33_groupi_n_199 ,csa_tree_add_6_33_groupi_n_61 ,csa_tree_add_6_33_groupi_n_158);
  nor csa_tree_add_6_33_groupi_g983__4319(csa_tree_add_6_33_groupi_n_195 ,csa_tree_add_6_33_groupi_n_143 ,csa_tree_add_6_33_groupi_n_167);
  or csa_tree_add_6_33_groupi_g984__8428(csa_tree_add_6_33_groupi_n_194 ,csa_tree_add_6_33_groupi_n_3 ,csa_tree_add_6_33_groupi_n_165);
  and csa_tree_add_6_33_groupi_g985__5526(csa_tree_add_6_33_groupi_n_193 ,csa_tree_add_6_33_groupi_n_56 ,csa_tree_add_6_33_groupi_n_165);
  not csa_tree_add_6_33_groupi_g986(csa_tree_add_6_33_groupi_n_192 ,csa_tree_add_6_33_groupi_n_191);
  or csa_tree_add_6_33_groupi_g987__6783(csa_tree_add_6_33_groupi_n_191 ,csa_tree_add_6_33_groupi_n_132 ,csa_tree_add_6_33_groupi_n_170);
  or csa_tree_add_6_33_groupi_g988__3680(csa_tree_add_6_33_groupi_n_190 ,csa_tree_add_6_33_groupi_n_140 ,csa_tree_add_6_33_groupi_n_169);
  or csa_tree_add_6_33_groupi_g989__1617(csa_tree_add_6_33_groupi_n_189 ,csa_tree_add_6_33_groupi_n_139 ,csa_tree_add_6_33_groupi_n_168);
  or csa_tree_add_6_33_groupi_g990__2802(csa_tree_add_6_33_groupi_n_188 ,csa_tree_add_6_33_groupi_n_145 ,csa_tree_add_6_33_groupi_n_166);
  or csa_tree_add_6_33_groupi_g991__1705(csa_tree_add_6_33_groupi_n_187 ,csa_tree_add_6_33_groupi_n_122 ,csa_tree_add_6_33_groupi_n_171);
  xnor csa_tree_add_6_33_groupi_g992__5122(csa_tree_add_6_33_groupi_n_186 ,csa_tree_add_6_33_groupi_n_86 ,csa_tree_add_6_33_groupi_n_120);
  xnor csa_tree_add_6_33_groupi_g993__8246(csa_tree_add_6_33_groupi_n_185 ,csa_tree_add_6_33_groupi_n_87 ,csa_tree_add_6_33_groupi_n_121);
  not csa_tree_add_6_33_groupi_g994(csa_tree_add_6_33_groupi_n_179 ,csa_tree_add_6_33_groupi_n_178);
  not csa_tree_add_6_33_groupi_g995(csa_tree_add_6_33_groupi_n_173 ,csa_tree_add_6_33_groupi_n_174);
  nor csa_tree_add_6_33_groupi_g996__7098(csa_tree_add_6_33_groupi_n_171 ,csa_tree_add_6_33_groupi_n_75 ,csa_tree_add_6_33_groupi_n_136);
  and csa_tree_add_6_33_groupi_g997__6131(csa_tree_add_6_33_groupi_n_170 ,csa_tree_add_6_33_groupi_n_133 ,csa_tree_add_6_33_groupi_n_126);
  nor csa_tree_add_6_33_groupi_g998__1881(csa_tree_add_6_33_groupi_n_169 ,csa_tree_add_6_33_groupi_n_62 ,csa_tree_add_6_33_groupi_n_138);
  nor csa_tree_add_6_33_groupi_g999__5115(csa_tree_add_6_33_groupi_n_168 ,csa_tree_add_6_33_groupi_n_76 ,csa_tree_add_6_33_groupi_n_142);
  nor csa_tree_add_6_33_groupi_g1000__7482(csa_tree_add_6_33_groupi_n_167 ,csa_tree_add_6_33_groupi_n_63 ,csa_tree_add_6_33_groupi_n_144);
  nor csa_tree_add_6_33_groupi_g1001__4733(csa_tree_add_6_33_groupi_n_166 ,csa_tree_add_6_33_groupi_n_64 ,csa_tree_add_6_33_groupi_n_137);
  or csa_tree_add_6_33_groupi_g1002__6161(csa_tree_add_6_33_groupi_n_184 ,csa_tree_add_6_33_groupi_n_108 ,csa_tree_add_6_33_groupi_n_129);
  or csa_tree_add_6_33_groupi_g1003__9315(csa_tree_add_6_33_groupi_n_183 ,csa_tree_add_6_33_groupi_n_101 ,csa_tree_add_6_33_groupi_n_128);
  or csa_tree_add_6_33_groupi_g1004__9945(csa_tree_add_6_33_groupi_n_182 ,csa_tree_add_6_33_groupi_n_106 ,csa_tree_add_6_33_groupi_n_123);
  or csa_tree_add_6_33_groupi_g1005__2883(csa_tree_add_6_33_groupi_n_181 ,csa_tree_add_6_33_groupi_n_103 ,csa_tree_add_6_33_groupi_n_127);
  or csa_tree_add_6_33_groupi_g1006__2346(csa_tree_add_6_33_groupi_n_180 ,csa_tree_add_6_33_groupi_n_117 ,csa_tree_add_6_33_groupi_n_134);
  or csa_tree_add_6_33_groupi_g1007__1666(csa_tree_add_6_33_groupi_n_178 ,csa_tree_add_6_33_groupi_n_116 ,csa_tree_add_6_33_groupi_n_125);
  and csa_tree_add_6_33_groupi_g1008__7410(csa_tree_add_6_33_groupi_n_177 ,csa_tree_add_6_33_groupi_n_112 ,csa_tree_add_6_33_groupi_n_146);
  or csa_tree_add_6_33_groupi_g1009__6417(csa_tree_add_6_33_groupi_n_176 ,csa_tree_add_6_33_groupi_n_119 ,csa_tree_add_6_33_groupi_n_130);
  or csa_tree_add_6_33_groupi_g1010__5477(csa_tree_add_6_33_groupi_n_175 ,csa_tree_add_6_33_groupi_n_111 ,csa_tree_add_6_33_groupi_n_124);
  or csa_tree_add_6_33_groupi_g1011__2398(csa_tree_add_6_33_groupi_n_174 ,csa_tree_add_6_33_groupi_n_78 ,csa_tree_add_6_33_groupi_n_131);
  or csa_tree_add_6_33_groupi_g1012__5107(csa_tree_add_6_33_groupi_n_172 ,csa_tree_add_6_33_groupi_n_118 ,csa_tree_add_6_33_groupi_n_135);
  xnor csa_tree_add_6_33_groupi_g1013__6260(out1[0] ,csa_tree_add_6_33_groupi_n_77 ,in3[0]);
  xnor csa_tree_add_6_33_groupi_g1014__4319(csa_tree_add_6_33_groupi_n_163 ,csa_tree_add_6_33_groupi_n_94 ,in2[13]);
  xnor csa_tree_add_6_33_groupi_g1015__8428(csa_tree_add_6_33_groupi_n_162 ,csa_tree_add_6_33_groupi_n_85 ,in2[18]);
  xnor csa_tree_add_6_33_groupi_g1016__5526(csa_tree_add_6_33_groupi_n_161 ,csa_tree_add_6_33_groupi_n_88 ,in2[16]);
  xnor csa_tree_add_6_33_groupi_g1017__6783(csa_tree_add_6_33_groupi_n_160 ,csa_tree_add_6_33_groupi_n_95 ,in2[12]);
  xnor csa_tree_add_6_33_groupi_g1018__3680(csa_tree_add_6_33_groupi_n_159 ,csa_tree_add_6_33_groupi_n_91 ,in2[4]);
  xnor csa_tree_add_6_33_groupi_g1019__1617(csa_tree_add_6_33_groupi_n_158 ,csa_tree_add_6_33_groupi_n_92 ,in2[3]);
  xnor csa_tree_add_6_33_groupi_g1020__2802(csa_tree_add_6_33_groupi_n_157 ,csa_tree_add_6_33_groupi_n_97 ,in2[11]);
  xnor csa_tree_add_6_33_groupi_g1021__1705(csa_tree_add_6_33_groupi_n_156 ,csa_tree_add_6_33_groupi_n_89 ,in2[14]);
  xnor csa_tree_add_6_33_groupi_g1022__5122(csa_tree_add_6_33_groupi_n_155 ,csa_tree_add_6_33_groupi_n_81 ,in2[9]);
  xnor csa_tree_add_6_33_groupi_g1023__8246(csa_tree_add_6_33_groupi_n_154 ,csa_tree_add_6_33_groupi_n_93 ,in2[10]);
  xnor csa_tree_add_6_33_groupi_g1024__7098(csa_tree_add_6_33_groupi_n_153 ,csa_tree_add_6_33_groupi_n_96 ,in2[15]);
  xnor csa_tree_add_6_33_groupi_g1025__6131(csa_tree_add_6_33_groupi_n_152 ,csa_tree_add_6_33_groupi_n_80 ,in1[1]);
  xnor csa_tree_add_6_33_groupi_g1026__1881(csa_tree_add_6_33_groupi_n_151 ,csa_tree_add_6_33_groupi_n_83 ,in2[8]);
  xnor csa_tree_add_6_33_groupi_g1027__5115(csa_tree_add_6_33_groupi_n_150 ,csa_tree_add_6_33_groupi_n_90 ,in2[17]);
  xnor csa_tree_add_6_33_groupi_g1028__7482(csa_tree_add_6_33_groupi_n_149 ,csa_tree_add_6_33_groupi_n_82 ,in2[7]);
  and csa_tree_add_6_33_groupi_g1029__4733(csa_tree_add_6_33_groupi_n_165 ,csa_tree_add_6_33_groupi_n_141 ,csa_tree_add_6_33_groupi_n_147);
  not csa_tree_add_6_33_groupi_g1030(csa_tree_add_6_33_groupi_n_147 ,csa_tree_add_6_33_groupi_n_148);
  or csa_tree_add_6_33_groupi_g1031__6161(csa_tree_add_6_33_groupi_n_146 ,csa_tree_add_6_33_groupi_n_110 ,csa_tree_add_6_33_groupi_n_91);
  nor csa_tree_add_6_33_groupi_g1032__9315(csa_tree_add_6_33_groupi_n_145 ,csa_tree_add_6_33_groupi_n_32 ,csa_tree_add_6_33_groupi_n_82);
  and csa_tree_add_6_33_groupi_g1033__9945(csa_tree_add_6_33_groupi_n_144 ,csa_tree_add_6_33_groupi_n_7 ,csa_tree_add_6_33_groupi_n_85);
  and csa_tree_add_6_33_groupi_g1034__2883(csa_tree_add_6_33_groupi_n_143 ,in2[18] ,csa_tree_add_6_33_groupi_n_84);
  and csa_tree_add_6_33_groupi_g1035__2346(csa_tree_add_6_33_groupi_n_142 ,csa_tree_add_6_33_groupi_n_37 ,csa_tree_add_6_33_groupi_n_83);
  or csa_tree_add_6_33_groupi_g1036__1666(csa_tree_add_6_33_groupi_n_141 ,csa_tree_add_6_33_groupi_n_28 ,csa_tree_add_6_33_groupi_n_98);
  nor csa_tree_add_6_33_groupi_g1037__7410(csa_tree_add_6_33_groupi_n_140 ,csa_tree_add_6_33_groupi_n_8 ,csa_tree_add_6_33_groupi_n_81);
  nor csa_tree_add_6_33_groupi_g1038__6417(csa_tree_add_6_33_groupi_n_139 ,csa_tree_add_6_33_groupi_n_37 ,csa_tree_add_6_33_groupi_n_83);
  and csa_tree_add_6_33_groupi_g1039__5477(csa_tree_add_6_33_groupi_n_138 ,csa_tree_add_6_33_groupi_n_8 ,csa_tree_add_6_33_groupi_n_81);
  and csa_tree_add_6_33_groupi_g1040__2398(csa_tree_add_6_33_groupi_n_137 ,csa_tree_add_6_33_groupi_n_32 ,csa_tree_add_6_33_groupi_n_82);
  nor csa_tree_add_6_33_groupi_g1041__5107(csa_tree_add_6_33_groupi_n_136 ,in2[6] ,csa_tree_add_6_33_groupi_n_86);
  nor csa_tree_add_6_33_groupi_g1042__6260(csa_tree_add_6_33_groupi_n_135 ,csa_tree_add_6_33_groupi_n_79 ,csa_tree_add_6_33_groupi_n_95);
  nor csa_tree_add_6_33_groupi_g1043__4319(csa_tree_add_6_33_groupi_n_134 ,csa_tree_add_6_33_groupi_n_115 ,csa_tree_add_6_33_groupi_n_96);
  and csa_tree_add_6_33_groupi_g1044__8428(csa_tree_add_6_33_groupi_n_148 ,csa_tree_add_6_33_groupi_n_28 ,csa_tree_add_6_33_groupi_n_98);
  and csa_tree_add_6_33_groupi_g1045__5526(csa_tree_add_6_33_groupi_n_132 ,in1[1] ,csa_tree_add_6_33_groupi_n_80);
  nor csa_tree_add_6_33_groupi_g1046__6783(csa_tree_add_6_33_groupi_n_131 ,csa_tree_add_6_33_groupi_n_109 ,csa_tree_add_6_33_groupi_n_92);
  nor csa_tree_add_6_33_groupi_g1047__3680(csa_tree_add_6_33_groupi_n_130 ,csa_tree_add_6_33_groupi_n_113 ,csa_tree_add_6_33_groupi_n_94);
  nor csa_tree_add_6_33_groupi_g1048__1617(csa_tree_add_6_33_groupi_n_129 ,csa_tree_add_6_33_groupi_n_107 ,csa_tree_add_6_33_groupi_n_93);
  nor csa_tree_add_6_33_groupi_g1049__2802(csa_tree_add_6_33_groupi_n_128 ,csa_tree_add_6_33_groupi_n_104 ,csa_tree_add_6_33_groupi_n_89);
  nor csa_tree_add_6_33_groupi_g1050__1705(csa_tree_add_6_33_groupi_n_127 ,csa_tree_add_6_33_groupi_n_100 ,csa_tree_add_6_33_groupi_n_90);
  or csa_tree_add_6_33_groupi_g1051__5122(csa_tree_add_6_33_groupi_n_126 ,in1[1] ,csa_tree_add_6_33_groupi_n_80);
  and csa_tree_add_6_33_groupi_g1052__8246(csa_tree_add_6_33_groupi_n_125 ,csa_tree_add_6_33_groupi_n_114 ,csa_tree_add_6_33_groupi_n_87);
  nor csa_tree_add_6_33_groupi_g1053__7098(csa_tree_add_6_33_groupi_n_124 ,csa_tree_add_6_33_groupi_n_99 ,csa_tree_add_6_33_groupi_n_97);
  nor csa_tree_add_6_33_groupi_g1054__6131(csa_tree_add_6_33_groupi_n_123 ,csa_tree_add_6_33_groupi_n_102 ,csa_tree_add_6_33_groupi_n_88);
  and csa_tree_add_6_33_groupi_g1055__1881(csa_tree_add_6_33_groupi_n_122 ,in2[6] ,csa_tree_add_6_33_groupi_n_86);
  xnor csa_tree_add_6_33_groupi_g1056__5115(csa_tree_add_6_33_groupi_n_121 ,csa_tree_add_6_33_groupi_n_73 ,in2[5]);
  xnor csa_tree_add_6_33_groupi_g1057__7482(csa_tree_add_6_33_groupi_n_120 ,csa_tree_add_6_33_groupi_n_75 ,in2[6]);
  or csa_tree_add_6_33_groupi_g1058__4733(csa_tree_add_6_33_groupi_n_133 ,csa_tree_add_6_33_groupi_n_55 ,csa_tree_add_6_33_groupi_n_105);
  nor csa_tree_add_6_33_groupi_g1059__6161(csa_tree_add_6_33_groupi_n_119 ,csa_tree_add_6_33_groupi_n_33 ,csa_tree_add_6_33_groupi_n_58);
  nor csa_tree_add_6_33_groupi_g1060__9315(csa_tree_add_6_33_groupi_n_118 ,csa_tree_add_6_33_groupi_n_30 ,csa_tree_add_6_33_groupi_n_57);
  nor csa_tree_add_6_33_groupi_g1061__9945(csa_tree_add_6_33_groupi_n_117 ,csa_tree_add_6_33_groupi_n_4 ,csa_tree_add_6_33_groupi_n_74);
  nor csa_tree_add_6_33_groupi_g1062__2883(csa_tree_add_6_33_groupi_n_116 ,csa_tree_add_6_33_groupi_n_34 ,csa_tree_add_6_33_groupi_n_73);
  and csa_tree_add_6_33_groupi_g1063__2346(csa_tree_add_6_33_groupi_n_115 ,csa_tree_add_6_33_groupi_n_4 ,csa_tree_add_6_33_groupi_n_74);
  or csa_tree_add_6_33_groupi_g1064__1666(csa_tree_add_6_33_groupi_n_114 ,in2[5] ,csa_tree_add_6_33_groupi_n_72);
  and csa_tree_add_6_33_groupi_g1065__7410(csa_tree_add_6_33_groupi_n_113 ,csa_tree_add_6_33_groupi_n_33 ,csa_tree_add_6_33_groupi_n_58);
  or csa_tree_add_6_33_groupi_g1066__6417(csa_tree_add_6_33_groupi_n_112 ,csa_tree_add_6_33_groupi_n_10 ,csa_tree_add_6_33_groupi_n_71);
  nor csa_tree_add_6_33_groupi_g1067__5477(csa_tree_add_6_33_groupi_n_111 ,csa_tree_add_6_33_groupi_n_9 ,csa_tree_add_6_33_groupi_n_67);
  nor csa_tree_add_6_33_groupi_g1068__2398(csa_tree_add_6_33_groupi_n_110 ,in2[4] ,csa_tree_add_6_33_groupi_n_70);
  and csa_tree_add_6_33_groupi_g1069__5107(csa_tree_add_6_33_groupi_n_109 ,csa_tree_add_6_33_groupi_n_6 ,csa_tree_add_6_33_groupi_n_61);
  nor csa_tree_add_6_33_groupi_g1070__6260(csa_tree_add_6_33_groupi_n_108 ,csa_tree_add_6_33_groupi_n_31 ,csa_tree_add_6_33_groupi_n_68);
  and csa_tree_add_6_33_groupi_g1071__4319(csa_tree_add_6_33_groupi_n_107 ,csa_tree_add_6_33_groupi_n_31 ,csa_tree_add_6_33_groupi_n_68);
  nor csa_tree_add_6_33_groupi_g1072__8428(csa_tree_add_6_33_groupi_n_106 ,csa_tree_add_6_33_groupi_n_36 ,csa_tree_add_6_33_groupi_n_69);
  and csa_tree_add_6_33_groupi_g1073__5526(csa_tree_add_6_33_groupi_n_105 ,in3[0] ,csa_tree_add_6_33_groupi_n_54);
  and csa_tree_add_6_33_groupi_g1074__6783(csa_tree_add_6_33_groupi_n_104 ,csa_tree_add_6_33_groupi_n_5 ,csa_tree_add_6_33_groupi_n_60);
  nor csa_tree_add_6_33_groupi_g1075__3680(csa_tree_add_6_33_groupi_n_103 ,csa_tree_add_6_33_groupi_n_35 ,csa_tree_add_6_33_groupi_n_59);
  and csa_tree_add_6_33_groupi_g1076__1617(csa_tree_add_6_33_groupi_n_102 ,csa_tree_add_6_33_groupi_n_36 ,csa_tree_add_6_33_groupi_n_69);
  nor csa_tree_add_6_33_groupi_g1077__2802(csa_tree_add_6_33_groupi_n_101 ,csa_tree_add_6_33_groupi_n_5 ,csa_tree_add_6_33_groupi_n_60);
  and csa_tree_add_6_33_groupi_g1078__1705(csa_tree_add_6_33_groupi_n_100 ,csa_tree_add_6_33_groupi_n_35 ,csa_tree_add_6_33_groupi_n_59);
  and csa_tree_add_6_33_groupi_g1079__5122(csa_tree_add_6_33_groupi_n_99 ,csa_tree_add_6_33_groupi_n_9 ,csa_tree_add_6_33_groupi_n_67);
  not csa_tree_add_6_33_groupi_g1080(csa_tree_add_6_33_groupi_n_84 ,csa_tree_add_6_33_groupi_n_85);
  and csa_tree_add_6_33_groupi_g1081__8246(csa_tree_add_6_33_groupi_n_79 ,csa_tree_add_6_33_groupi_n_30 ,csa_tree_add_6_33_groupi_n_57);
  nor csa_tree_add_6_33_groupi_g1082__7098(csa_tree_add_6_33_groupi_n_78 ,csa_tree_add_6_33_groupi_n_6 ,csa_tree_add_6_33_groupi_n_61);
  xnor csa_tree_add_6_33_groupi_g1083__6131(csa_tree_add_6_33_groupi_n_77 ,in1[0] ,in2[0]);
  xnor csa_tree_add_6_33_groupi_g1084__1881(csa_tree_add_6_33_groupi_n_98 ,in3[2] ,in1[2]);
  xnor csa_tree_add_6_33_groupi_g1085__5115(csa_tree_add_6_33_groupi_n_97 ,in3[11] ,in1[11]);
  xnor csa_tree_add_6_33_groupi_g1086__7482(csa_tree_add_6_33_groupi_n_96 ,in3[15] ,in1[15]);
  xnor csa_tree_add_6_33_groupi_g1087__4733(csa_tree_add_6_33_groupi_n_95 ,in3[12] ,in1[12]);
  xnor csa_tree_add_6_33_groupi_g1088__6161(csa_tree_add_6_33_groupi_n_94 ,in3[13] ,in1[13]);
  xnor csa_tree_add_6_33_groupi_g1089__9315(csa_tree_add_6_33_groupi_n_93 ,in3[10] ,in1[10]);
  xnor csa_tree_add_6_33_groupi_g1090__9945(csa_tree_add_6_33_groupi_n_92 ,in3[3] ,in1[3]);
  xnor csa_tree_add_6_33_groupi_g1091__2883(csa_tree_add_6_33_groupi_n_91 ,in3[4] ,in1[4]);
  xnor csa_tree_add_6_33_groupi_g1092__2346(csa_tree_add_6_33_groupi_n_90 ,in3[17] ,in1[17]);
  xnor csa_tree_add_6_33_groupi_g1093__1666(csa_tree_add_6_33_groupi_n_89 ,in3[14] ,in1[14]);
  xnor csa_tree_add_6_33_groupi_g1094__7410(csa_tree_add_6_33_groupi_n_88 ,in3[16] ,in1[16]);
  xnor csa_tree_add_6_33_groupi_g1095__6417(csa_tree_add_6_33_groupi_n_87 ,in3[5] ,in1[5]);
  xnor csa_tree_add_6_33_groupi_g1096__5477(csa_tree_add_6_33_groupi_n_86 ,in3[6] ,in1[6]);
  xnor csa_tree_add_6_33_groupi_g1097__2398(csa_tree_add_6_33_groupi_n_85 ,in3[18] ,in1[18]);
  xnor csa_tree_add_6_33_groupi_g1098__5107(csa_tree_add_6_33_groupi_n_83 ,in3[8] ,in1[8]);
  xnor csa_tree_add_6_33_groupi_g1099__6260(csa_tree_add_6_33_groupi_n_82 ,in3[7] ,in1[7]);
  xnor csa_tree_add_6_33_groupi_g1100__4319(csa_tree_add_6_33_groupi_n_81 ,in3[9] ,in1[9]);
  or csa_tree_add_6_33_groupi_g1101__8428(csa_tree_add_6_33_groupi_n_80 ,csa_tree_add_6_33_groupi_n_66 ,csa_tree_add_6_33_groupi_n_3);
  not csa_tree_add_6_33_groupi_g1102(csa_tree_add_6_33_groupi_n_72 ,csa_tree_add_6_33_groupi_n_73);
  not csa_tree_add_6_33_groupi_g1103(csa_tree_add_6_33_groupi_n_70 ,csa_tree_add_6_33_groupi_n_71);
  and csa_tree_add_6_33_groupi_g1104__5526(csa_tree_add_6_33_groupi_n_66 ,in3[1] ,in2[1]);
  nand csa_tree_add_6_33_groupi_g1105__6783(csa_tree_add_6_33_groupi_n_65 ,in3[18] ,in1[18]);
  or csa_tree_add_6_33_groupi_g1106__3680(csa_tree_add_6_33_groupi_n_76 ,csa_tree_add_6_33_groupi_n_52 ,csa_tree_add_6_33_groupi_n_15);
  and csa_tree_add_6_33_groupi_g1107__1617(csa_tree_add_6_33_groupi_n_75 ,csa_tree_add_6_33_groupi_n_41 ,csa_tree_add_6_33_groupi_n_39);
  or csa_tree_add_6_33_groupi_g1108__2802(csa_tree_add_6_33_groupi_n_74 ,csa_tree_add_6_33_groupi_n_40 ,csa_tree_add_6_33_groupi_n_48);
  or csa_tree_add_6_33_groupi_g1109__1705(csa_tree_add_6_33_groupi_n_73 ,csa_tree_add_6_33_groupi_n_46 ,csa_tree_add_6_33_groupi_n_18);
  or csa_tree_add_6_33_groupi_g1110__5122(csa_tree_add_6_33_groupi_n_71 ,csa_tree_add_6_33_groupi_n_22 ,csa_tree_add_6_33_groupi_n_27);
  or csa_tree_add_6_33_groupi_g1111__8246(csa_tree_add_6_33_groupi_n_69 ,csa_tree_add_6_33_groupi_n_16 ,csa_tree_add_6_33_groupi_n_13);
  or csa_tree_add_6_33_groupi_g1112__7098(csa_tree_add_6_33_groupi_n_68 ,csa_tree_add_6_33_groupi_n_47 ,csa_tree_add_6_33_groupi_n_43);
  or csa_tree_add_6_33_groupi_g1113__6131(csa_tree_add_6_33_groupi_n_67 ,csa_tree_add_6_33_groupi_n_11 ,csa_tree_add_6_33_groupi_n_42);
  and csa_tree_add_6_33_groupi_g1114__1881(csa_tree_add_6_33_groupi_n_55 ,in1[0] ,in2[0]);
  or csa_tree_add_6_33_groupi_g1115__5115(csa_tree_add_6_33_groupi_n_54 ,in1[0] ,in2[0]);
  and csa_tree_add_6_33_groupi_g1116__7482(csa_tree_add_6_33_groupi_n_64 ,csa_tree_add_6_33_groupi_n_50 ,csa_tree_add_6_33_groupi_n_14);
  or csa_tree_add_6_33_groupi_g1117__4733(csa_tree_add_6_33_groupi_n_63 ,csa_tree_add_6_33_groupi_n_23 ,csa_tree_add_6_33_groupi_n_45);
  or csa_tree_add_6_33_groupi_g1118__6161(csa_tree_add_6_33_groupi_n_62 ,csa_tree_add_6_33_groupi_n_24 ,csa_tree_add_6_33_groupi_n_12);
  or csa_tree_add_6_33_groupi_g1119__9315(csa_tree_add_6_33_groupi_n_61 ,csa_tree_add_6_33_groupi_n_21 ,csa_tree_add_6_33_groupi_n_20);
  or csa_tree_add_6_33_groupi_g1120__9945(csa_tree_add_6_33_groupi_n_60 ,csa_tree_add_6_33_groupi_n_38 ,csa_tree_add_6_33_groupi_n_19);
  or csa_tree_add_6_33_groupi_g1121__2883(csa_tree_add_6_33_groupi_n_59 ,csa_tree_add_6_33_groupi_n_17 ,csa_tree_add_6_33_groupi_n_51);
  or csa_tree_add_6_33_groupi_g1122__2346(csa_tree_add_6_33_groupi_n_58 ,csa_tree_add_6_33_groupi_n_25 ,csa_tree_add_6_33_groupi_n_26);
  or csa_tree_add_6_33_groupi_g1123__1666(csa_tree_add_6_33_groupi_n_57 ,csa_tree_add_6_33_groupi_n_49 ,csa_tree_add_6_33_groupi_n_44);
  and csa_tree_add_6_33_groupi_g1124__7410(csa_tree_add_6_33_groupi_n_56 ,csa_tree_add_6_33_groupi_n_29 ,csa_tree_add_6_33_groupi_n_53);
  not csa_tree_add_6_33_groupi_g1125(csa_tree_add_6_33_groupi_n_53 ,in2[1]);
  not csa_tree_add_6_33_groupi_g1126(csa_tree_add_6_33_groupi_n_52 ,in3[7]);
  not csa_tree_add_6_33_groupi_g1127(csa_tree_add_6_33_groupi_n_51 ,in1[16]);
  not csa_tree_add_6_33_groupi_g1128(csa_tree_add_6_33_groupi_n_50 ,in3[6]);
  not csa_tree_add_6_33_groupi_g1129(csa_tree_add_6_33_groupi_n_49 ,in3[11]);
  not csa_tree_add_6_33_groupi_g1130(csa_tree_add_6_33_groupi_n_48 ,in1[14]);
  not csa_tree_add_6_33_groupi_g1131(csa_tree_add_6_33_groupi_n_47 ,in3[9]);
  not csa_tree_add_6_33_groupi_g1132(csa_tree_add_6_33_groupi_n_46 ,in3[4]);
  not csa_tree_add_6_33_groupi_g1133(csa_tree_add_6_33_groupi_n_45 ,in1[17]);
  not csa_tree_add_6_33_groupi_g1134(csa_tree_add_6_33_groupi_n_44 ,in1[11]);
  not csa_tree_add_6_33_groupi_g1135(csa_tree_add_6_33_groupi_n_43 ,in1[9]);
  not csa_tree_add_6_33_groupi_g1136(csa_tree_add_6_33_groupi_n_42 ,in1[10]);
  not csa_tree_add_6_33_groupi_g1137(csa_tree_add_6_33_groupi_n_41 ,in3[5]);
  not csa_tree_add_6_33_groupi_g1138(csa_tree_add_6_33_groupi_n_40 ,in3[14]);
  not csa_tree_add_6_33_groupi_g1139(csa_tree_add_6_33_groupi_n_39 ,in1[5]);
  not csa_tree_add_6_33_groupi_g1140(csa_tree_add_6_33_groupi_n_38 ,in3[13]);
  not csa_tree_add_6_33_groupi_g1141(csa_tree_add_6_33_groupi_n_37 ,in2[8]);
  not csa_tree_add_6_33_groupi_g1142(csa_tree_add_6_33_groupi_n_36 ,in2[16]);
  not csa_tree_add_6_33_groupi_g1143(csa_tree_add_6_33_groupi_n_35 ,in2[17]);
  not csa_tree_add_6_33_groupi_g1144(csa_tree_add_6_33_groupi_n_34 ,in2[5]);
  not csa_tree_add_6_33_groupi_g1145(csa_tree_add_6_33_groupi_n_33 ,in2[13]);
  not csa_tree_add_6_33_groupi_g1146(csa_tree_add_6_33_groupi_n_32 ,in2[7]);
  not csa_tree_add_6_33_groupi_g1147(csa_tree_add_6_33_groupi_n_31 ,in2[10]);
  not csa_tree_add_6_33_groupi_g1148(csa_tree_add_6_33_groupi_n_30 ,in2[12]);
  not csa_tree_add_6_33_groupi_g1149(csa_tree_add_6_33_groupi_n_29 ,in3[1]);
  not csa_tree_add_6_33_groupi_g1150(csa_tree_add_6_33_groupi_n_28 ,in2[2]);
  not csa_tree_add_6_33_groupi_g1151(csa_tree_add_6_33_groupi_n_27 ,in1[3]);
  not csa_tree_add_6_33_groupi_g1152(csa_tree_add_6_33_groupi_n_26 ,in1[12]);
  not csa_tree_add_6_33_groupi_g1153(csa_tree_add_6_33_groupi_n_25 ,in3[12]);
  not csa_tree_add_6_33_groupi_g1154(csa_tree_add_6_33_groupi_n_24 ,in3[8]);
  not csa_tree_add_6_33_groupi_g1155(csa_tree_add_6_33_groupi_n_23 ,in3[17]);
  not csa_tree_add_6_33_groupi_g1156(csa_tree_add_6_33_groupi_n_22 ,in3[3]);
  not csa_tree_add_6_33_groupi_g1157(csa_tree_add_6_33_groupi_n_21 ,in3[2]);
  not csa_tree_add_6_33_groupi_g1158(csa_tree_add_6_33_groupi_n_20 ,in1[2]);
  not csa_tree_add_6_33_groupi_g1159(csa_tree_add_6_33_groupi_n_19 ,in1[13]);
  not csa_tree_add_6_33_groupi_g1160(csa_tree_add_6_33_groupi_n_18 ,in1[4]);
  not csa_tree_add_6_33_groupi_g1161(csa_tree_add_6_33_groupi_n_17 ,in3[16]);
  not csa_tree_add_6_33_groupi_g1162(csa_tree_add_6_33_groupi_n_16 ,in3[15]);
  not csa_tree_add_6_33_groupi_g1163(csa_tree_add_6_33_groupi_n_15 ,in1[7]);
  not csa_tree_add_6_33_groupi_g1164(csa_tree_add_6_33_groupi_n_14 ,in1[6]);
  not csa_tree_add_6_33_groupi_g1165(csa_tree_add_6_33_groupi_n_13 ,in1[15]);
  not csa_tree_add_6_33_groupi_g1166(csa_tree_add_6_33_groupi_n_12 ,in1[8]);
  not csa_tree_add_6_33_groupi_g1167(csa_tree_add_6_33_groupi_n_11 ,in3[10]);
  not csa_tree_add_6_33_groupi_g1168(csa_tree_add_6_33_groupi_n_10 ,in2[4]);
  not csa_tree_add_6_33_groupi_g1169(csa_tree_add_6_33_groupi_n_9 ,in2[11]);
  not csa_tree_add_6_33_groupi_g1170(csa_tree_add_6_33_groupi_n_8 ,in2[9]);
  not csa_tree_add_6_33_groupi_g1171(csa_tree_add_6_33_groupi_n_7 ,in2[18]);
  not csa_tree_add_6_33_groupi_g1172(csa_tree_add_6_33_groupi_n_6 ,in2[3]);
  not csa_tree_add_6_33_groupi_g1173(csa_tree_add_6_33_groupi_n_5 ,in2[14]);
  not csa_tree_add_6_33_groupi_g1174(csa_tree_add_6_33_groupi_n_4 ,in2[15]);
  not csa_tree_add_6_33_groupi_drc_bufs1175(csa_tree_add_6_33_groupi_n_3 ,csa_tree_add_6_33_groupi_n_2);
  not csa_tree_add_6_33_groupi_drc_bufs1176(csa_tree_add_6_33_groupi_n_2 ,csa_tree_add_6_33_groupi_n_56);
  xor csa_tree_add_6_33_groupi_g2__6417(out1[5] ,csa_tree_add_6_33_groupi_n_270 ,csa_tree_add_6_33_groupi_n_220);
  xor csa_tree_add_6_33_groupi_g1179__5477(out1[4] ,csa_tree_add_6_33_groupi_n_267 ,csa_tree_add_6_33_groupi_n_251);
endmodule
