module top( n5 , n16 , n23 , n24 , n31 , n38 , n41 , n44 , n46 , n53 , n55 , n57 , n62 , n63 , n68 , n71 , n72 , n78 , n79 , n84 , n92 , n96 , n98 , n101 , n106 , n107 , n120 , n123 , n126 , n136 , n142 , n144 , n145 , n153 , n165 , n177 , n182 , n216 , n220 );
    input n16 , n23 , n24 , n31 , n38 , n41 , n44 , n46 , n53 , n55 , n57 , n62 , n68 , n71 , n72 , n79 , n84 , n92 , n96 , n98 , n101 , n106 , n107 , n120 , n123 , n136 , n145 , n165 , n177 , n182 , n216 , n220 ;
    output n5 , n63 , n78 , n126 , n142 , n144 , n153 ;
    wire n0 , n1 , n2 , n3 , n4 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n17 , n18 , n19 , n20 , n21 , n22 , n25 , n26 , n27 , n28 , n29 , n30 , n32 , n33 , n34 , n35 , n36 , n37 , n39 , n40 , n42 , n43 , n45 , n47 , n48 , n49 , n50 , n51 , n52 , n54 , n56 , n58 , n59 , n60 , n61 , n64 , n65 , n66 , n67 , n69 , n70 , n73 , n74 , n75 , n76 , n77 , n80 , n81 , n82 , n83 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n93 , n94 , n95 , n97 , n99 , n100 , n102 , n103 , n104 , n105 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n121 , n122 , n124 , n125 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n137 , n138 , n139 , n140 , n141 , n143 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n178 , n179 , n180 , n181 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n217 , n218 , n219 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 ;
assign n17 = ~n38;
assign n211 = n18 & n116;
assign n193 = ~n195;
assign n81 = n118 & n84;
assign n75 = n173 | n113;
assign n180 = n132 & n55;
assign n89 = n125 & n136;
assign n103 = n164 | n131;
assign n127 = n226 & n176;
assign n155 = ~(n198 | n179);
assign n18 = ~n195;
assign n21 = n180 & n59;
assign n42 = n121 & n170;
assign n209 = n159 & n98;
assign n28 = ~(n107 | n70);
assign n135 = n139 & n96;
assign n100 = n209 | n1;
assign n172 = n8 | n230;
assign n78 = n97 | n115;
assign n186 = n229 | n86;
assign n111 = n28 & n68;
assign n88 = ~n37;
assign n95 = ~n129;
assign n199 = n193 & n71;
assign n2 = ~(n190 | n118);
assign n47 = ~n61;
assign n179 = n199 | n81;
assign n200 = ~(n58 | n194);
assign n205 = n155 & n38;
assign n26 = ~(n75 | n115);
assign n105 = ~n170;
assign n152 = n153 & n120;
assign n131 = n88 & n31;
assign n201 = ~n212;
assign n80 = n227 & n53;
assign n217 = ~n67;
assign n51 = n41 | n7;
assign n109 = n218 & n10;
assign n11 = ~(n33 | n64);
assign n215 = n80 & n50;
assign n52 = ~n106;
assign n159 = ~n47;
assign n114 = ~(n157 | n125);
assign n110 = ~(n79 | n82);
assign n83 = n95 & n79;
assign n133 = n171 | n2;
assign n162 = n66 & n9;
assign n112 = ~n182;
assign n138 = ~(n89 | n102);
assign n174 = ~n217;
assign n39 = n50 | n204;
assign n99 = n0 & n35;
assign n116 = n71 | n17;
assign n50 = n25 & n53;
assign n70 = n5 & n206;
assign n194 = n138 & n53;
assign n160 = n6 & n11;
assign n82 = n159 & n163;
assign n212 = n223 & n51;
assign n161 = n193 & n165;
assign n183 = n171 & n162;
assign n6 = ~(n181 | n196);
assign n158 = n80 | n137;
assign n91 = n29 & n48;
assign n29 = n210 & n38;
assign n204 = n29 | n221;
assign n102 = n166 | n60;
assign n35 = n169 | n180;
assign n169 = n168 & n182;
assign n32 = n147 | n191;
assign n25 = ~(n136 | n54);
assign n33 = n119 | n85;
assign n154 = n141 & n51;
assign n73 = n46 | n112;
assign n139 = ~(n62 | n186);
assign n227 = ~(n177 | n54);
assign n143 = n172 | n78;
assign n184 = ~(n31 | n128);
assign n141 = n44 | n77;
assign n59 = n110 & n55;
assign n27 = n213 & n230;
assign n178 = n137 & n111;
assign n124 = ~n145;
assign n22 = n111 | n108;
assign n148 = n52 | n76;
assign n86 = n153 & n32;
assign n45 = ~n195;
assign n153 = ~n49;
assign n214 = ~n75;
assign n173 = ~n68;
assign n66 = ~n190;
assign n74 = n169 & n189;
assign n9 = ~n92;
assign n134 = n83 | n222;
assign n208 = n34 & n36;
assign n7 = ~n84;
assign n163 = n165 | n56;
assign n170 = n147 | n104;
assign n30 = ~(n182 | n143);
assign n54 = n45 & n141;
assign n128 = n90 & n10;
assign n130 = ~n103;
assign n157 = ~(n48 | n34);
assign n225 = ~n13;
assign n5 = ~n192;
assign n15 = ~(n185 | n140);
assign n34 = n184 & n84;
assign n12 = ~n101;
assign n48 = n228 & n7;
assign n10 = ~n185;
assign n140 = n195 & n84;
assign n171 = n66 & n24;
assign n206 = n57 | n173;
assign n226 = n20 & n116;
assign n4 = n87 & n73;
assign n122 = ~n211;
assign n63 = n149 & n103;
assign n13 = ~n40;
assign n20 = n154 & n73;
assign n207 = n91 | n208;
assign n164 = n15 | n152;
assign n166 = n45 & n44;
assign n228 = n122 & n38;
assign n67 = ~n203;
assign n121 = ~(n200 | n26);
assign n0 = n203;
assign n65 = ~(n189 | n39);
assign n40 = ~n76;
assign n189 = n175 & n182;
assign n132 = ~(n16 | n82);
assign n168 = ~(n220 | n4);
assign n175 = ~(n123 | n4);
assign n156 = ~(n216 | n70);
assign n119 = n215 | n178;
assign n94 = n127 & n163;
assign n56 = ~n55;
assign n60 = n225 & n177;
assign n187 = n201 & n52;
assign n149 = n3 | n42;
assign n76 = n160 & n219;
assign n142 = ~n13;
assign n198 = n146 & n23;
assign n19 = n146 & n72;
assign n3 = n148 & n201;
assign n185 = n12 & n84;
assign n144 = ~(n205 | n30);
assign n167 = n74 | n21;
assign n117 = n18 & n57;
assign n181 = n167 | n99;
assign n190 = n124 | n87;
assign n230 = n194 | n214;
assign n210 = ~(n23 | n211);
assign n191 = n72 | n229;
assign n150 = n88 & n216;
assign n8 = ~n58;
assign n113 = n224 | n93;
assign n126 = ~(n97 | n27);
assign n36 = n43 & n84;
assign n64 = n207 | n114;
assign n176 = n98 | n147;
assign n196 = n183 | n135;
assign n129 = ~n67;
assign n43 = ~(n120 | n128);
assign n218 = n94 & n206;
assign n213 = ~n115;
assign n137 = n156 & n68;
assign n104 = n19 | n100;
assign n146 = ~n129;
assign n61 = ~n109;
assign n49 = ~n174;
assign n97 = n130 | n3;
assign n188 = ~n32;
assign n203 = n65 & n212;
assign n197 = n59 | n22;
assign n223 = ~n140;
assign n202 = n133 & n151;
assign n221 = n36 | n197;
assign n90 = ~n47;
assign n195 = n109;
assign n229 = n90 & n176;
assign n85 = n0 & n158;
assign n147 = ~n96;
assign n69 = n225 & n16;
assign n87 = ~n192;
assign n224 = n95 & n107;
assign n151 = n9 | n0;
assign n125 = ~n217;
assign n108 = n188 | n162;
assign n93 = n117 | n150;
assign n115 = n202 | n105;
assign n77 = ~n53;
assign n1 = n142 & n62;
assign n58 = n56 | n134;
assign n192 = ~n61;
assign n37 = ~n40;
assign n222 = n161 | n69;
assign n219 = ~(n187 | n14);
assign n118 = ~n37;
assign n14 = n0 & n171;
endmodule
