module top( n1 , n8 , n9 , n21 , n24 , n32 , n54 , n61 , n64 , n67 , n69 , n76 , n83 , n84 , n96 , n97 , n107 , n110 , n117 , n120 , n128 , n135 , n137 , n142 , n145 , n147 , n150 , n154 , n167 , n170 , n172 , n182 , n184 , n190 , n198 , n204 , n209 , n210 , n220 , n222 , n230 , n231 , n232 , n233 , n240 , n253 , n265 , n268 , n269 , n283 , n289 , n290 , n291 , n292 , n293 , n296 , n313 , n324 , n325 , n330 , n336 , n342 , n347 , n350 , n356 , n362 , n363 , n364 , n365 , n368 , n373 , n383 , n386 , n388 , n403 , n415 , n418 , n421 , n427 , n432 , n434 , n468 , n476 , n478 , n480 , n481 , n489 , n490 , n506 , n507 , n514 , n524 , n526 , n532 , n543 , n565 , n574 , n576 , n579 , n588 , n596 , n598 , n605 , n608 , n614 , n615 , n618 , n623 , n629 , n633 , n635 , n640 , n646 , n654 , n656 , n663 , n664 , n675 , n676 , n677 , n678 , n691 , n693 , n704 , n710 , n716 , n717 , n722 , n726 , n727 , n737 , n740 , n750 , n751 , n765 , n769 , n785 , n786 , n790 , n793 , n794 , n797 , n800 , n814 , n818 , n821 , n824 , n829 , n835 , n836 , n837 , n840 , n842 , n845 , n848 , n851 , n857 , n859 , n869 , n877 , n887 , n894 , n901 , n909 , n923 , n928 , n933 , n934 , n938 , n950 , n956 , n964 , n973 , n974 , n989 , n990 , n1013 , n1014 , n1019 , n1021 , n1023 , n1025 , n1026 , n1030 , n1032 , n1036 , n1039 , n1042 , n1043 , n1049 , n1052 , n1058 , n1065 , n1070 , n1091 , n1093 , n1098 , n1099 , n1108 , n1117 , n1121 , n1122 , n1131 , n1134 , n1138 , n1143 , n1146 , n1150 , n1151 , n1157 , n1160 , n1161 , n1162 , n1165 , n1170 , n1177 , n1184 , n1187 , n1189 , n1192 , n1194 , n1198 , n1223 , n1239 , n1240 , n1243 , n1251 , n1253 , n1255 , n1275 , n1276 , n1280 , n1303 , n1310 , n1311 , n1314 , n1331 , n1335 , n1339 , n1361 , n1366 , n1373 , n1375 , n1378 , n1389 , n1392 , n1396 , n1398 , n1407 , n1409 , n1411 , n1412 , n1413 , n1418 , n1422 , n1425 , n1438 , n1442 , n1454 , n1474 , n1475 , n1478 , n1479 , n1485 , n1508 , n1511 , n1512 , n1515 , n1518 , n1530 , n1531 , n1542 , n1545 , n1547 , n1549 , n1551 , n1552 , n1555 , n1556 , n1562 , n1574 , n1575 , n1580 , n1581 , n1589 , n1594 , n1596 , n1601 , n1604 , n1606 , n1620 , n1628 , n1629 , n1630 , n1631 , n1645 , n1648 , n1655 , n1665 , n1671 , n1676 );
    input n1 , n9 , n67 , n69 , n84 , n96 , n107 , n120 , n128 , n135 , n137 , n145 , n147 , n182 , n184 , n198 , n209 , n220 , n222 , n230 , n233 , n268 , n283 , n289 , n290 , n293 , n296 , n325 , n330 , n342 , n356 , n362 , n365 , n373 , n386 , n403 , n415 , n418 , n421 , n432 , n468 , n478 , n481 , n490 , n507 , n514 , n526 , n532 , n574 , n576 , n579 , n588 , n596 , n605 , n615 , n629 , n635 , n646 , n654 , n664 , n677 , n704 , n710 , n716 , n726 , n727 , n737 , n750 , n751 , n765 , n769 , n793 , n794 , n797 , n818 , n824 , n829 , n835 , n837 , n842 , n848 , n851 , n857 , n859 , n869 , n877 , n901 , n909 , n923 , n933 , n934 , n938 , n950 , n956 , n973 , n974 , n989 , n990 , n1013 , n1014 , n1025 , n1030 , n1042 , n1049 , n1052 , n1058 , n1065 , n1070 , n1091 , n1093 , n1098 , n1099 , n1108 , n1121 , n1131 , n1134 , n1143 , n1146 , n1150 , n1161 , n1162 , n1165 , n1170 , n1184 , n1187 , n1189 , n1223 , n1240 , n1243 , n1251 , n1253 , n1255 , n1276 , n1280 , n1303 , n1310 , n1311 , n1331 , n1335 , n1339 , n1361 , n1366 , n1373 , n1378 , n1389 , n1396 , n1398 , n1407 , n1409 , n1412 , n1413 , n1418 , n1422 , n1425 , n1438 , n1475 , n1479 , n1485 , n1508 , n1511 , n1515 , n1518 , n1530 , n1545 , n1549 , n1551 , n1555 , n1562 , n1575 , n1580 , n1581 , n1596 , n1606 , n1620 , n1630 , n1648 , n1655 , n1676 ;
    output n8 , n21 , n24 , n32 , n54 , n61 , n64 , n76 , n83 , n97 , n110 , n117 , n142 , n150 , n154 , n167 , n170 , n172 , n190 , n204 , n210 , n231 , n232 , n240 , n253 , n265 , n269 , n291 , n292 , n313 , n324 , n336 , n347 , n350 , n363 , n364 , n368 , n383 , n388 , n427 , n434 , n476 , n480 , n489 , n506 , n524 , n543 , n565 , n598 , n608 , n614 , n618 , n623 , n633 , n640 , n656 , n663 , n675 , n676 , n678 , n691 , n693 , n717 , n722 , n740 , n785 , n786 , n790 , n800 , n814 , n821 , n836 , n840 , n845 , n887 , n894 , n928 , n964 , n1019 , n1021 , n1023 , n1026 , n1032 , n1036 , n1039 , n1043 , n1117 , n1122 , n1138 , n1151 , n1157 , n1160 , n1177 , n1192 , n1194 , n1198 , n1239 , n1275 , n1314 , n1375 , n1392 , n1411 , n1442 , n1454 , n1474 , n1478 , n1512 , n1531 , n1542 , n1547 , n1552 , n1556 , n1574 , n1589 , n1594 , n1601 , n1604 , n1628 , n1629 , n1631 , n1645 , n1665 , n1671 ;
    wire n0 , n2 , n3 , n4 , n5 , n6 , n7 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n22 , n23 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n55 , n56 , n57 , n58 , n59 , n60 , n62 , n63 , n65 , n66 , n68 , n70 , n71 , n72 , n73 , n74 , n75 , n77 , n78 , n79 , n80 , n81 , n82 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n108 , n109 , n111 , n112 , n113 , n114 , n115 , n116 , n118 , n119 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n129 , n130 , n131 , n132 , n133 , n134 , n136 , n138 , n139 , n140 , n141 , n143 , n144 , n146 , n148 , n149 , n151 , n152 , n153 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n168 , n169 , n171 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n183 , n185 , n186 , n187 , n188 , n189 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n199 , n200 , n201 , n202 , n203 , n205 , n206 , n207 , n208 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n221 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n234 , n235 , n236 , n237 , n238 , n239 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n266 , n267 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n284 , n285 , n286 , n287 , n288 , n294 , n295 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n326 , n327 , n328 , n329 , n331 , n332 , n333 , n334 , n335 , n337 , n338 , n339 , n340 , n341 , n343 , n344 , n345 , n346 , n348 , n349 , n351 , n352 , n353 , n354 , n355 , n357 , n358 , n359 , n360 , n361 , n366 , n367 , n369 , n370 , n371 , n372 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n384 , n385 , n387 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n416 , n417 , n419 , n420 , n422 , n423 , n424 , n425 , n426 , n428 , n429 , n430 , n431 , n433 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n477 , n479 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n508 , n509 , n510 , n511 , n512 , n513 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n525 , n527 , n528 , n529 , n530 , n531 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n575 , n577 , n578 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n597 , n599 , n600 , n601 , n602 , n603 , n604 , n606 , n607 , n609 , n610 , n611 , n612 , n613 , n616 , n617 , n619 , n620 , n621 , n622 , n624 , n625 , n626 , n627 , n628 , n630 , n631 , n632 , n634 , n636 , n637 , n638 , n639 , n641 , n642 , n643 , n644 , n645 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n655 , n657 , n658 , n659 , n660 , n661 , n662 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n692 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n705 , n706 , n707 , n708 , n709 , n711 , n712 , n713 , n714 , n715 , n718 , n719 , n720 , n721 , n723 , n724 , n725 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n738 , n739 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n766 , n767 , n768 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n787 , n788 , n789 , n791 , n792 , n795 , n796 , n798 , n799 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n815 , n816 , n817 , n819 , n820 , n822 , n823 , n825 , n826 , n827 , n828 , n830 , n831 , n832 , n833 , n834 , n838 , n839 , n841 , n843 , n844 , n846 , n847 , n849 , n850 , n852 , n853 , n854 , n855 , n856 , n858 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n888 , n889 , n890 , n891 , n892 , n893 , n895 , n896 , n897 , n898 , n899 , n900 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n924 , n925 , n926 , n927 , n929 , n930 , n931 , n932 , n935 , n936 , n937 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n951 , n952 , n953 , n954 , n955 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1015 , n1016 , n1017 , n1018 , n1020 , n1022 , n1024 , n1027 , n1028 , n1029 , n1031 , n1033 , n1034 , n1035 , n1037 , n1038 , n1040 , n1041 , n1044 , n1045 , n1046 , n1047 , n1048 , n1050 , n1051 , n1053 , n1054 , n1055 , n1056 , n1057 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1066 , n1067 , n1068 , n1069 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1092 , n1094 , n1095 , n1096 , n1097 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1118 , n1119 , n1120 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1132 , n1133 , n1135 , n1136 , n1137 , n1139 , n1140 , n1141 , n1142 , n1144 , n1145 , n1147 , n1148 , n1149 , n1152 , n1153 , n1154 , n1155 , n1156 , n1158 , n1159 , n1163 , n1164 , n1166 , n1167 , n1168 , n1169 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1185 , n1186 , n1188 , n1190 , n1191 , n1193 , n1195 , n1196 , n1197 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1241 , n1242 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1252 , n1254 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1277 , n1278 , n1279 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1312 , n1313 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1332 , n1333 , n1334 , n1336 , n1337 , n1338 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1362 , n1363 , n1364 , n1365 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1374 , n1376 , n1377 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1390 , n1391 , n1393 , n1394 , n1395 , n1397 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1408 , n1410 , n1414 , n1415 , n1416 , n1417 , n1419 , n1420 , n1421 , n1423 , n1424 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1439 , n1440 , n1441 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1476 , n1477 , n1480 , n1481 , n1482 , n1483 , n1484 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1509 , n1510 , n1513 , n1514 , n1516 , n1517 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1543 , n1544 , n1546 , n1548 , n1550 , n1553 , n1554 , n1557 , n1558 , n1559 , n1560 , n1561 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1576 , n1577 , n1578 , n1579 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1590 , n1591 , n1592 , n1593 , n1595 , n1597 , n1598 , n1599 , n1600 , n1602 , n1603 , n1605 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1646 , n1647 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1666 , n1667 , n1668 , n1669 , n1670 , n1672 , n1673 , n1674 , n1675 , n1677 ;
assign n806 = ~(n1255 | n1030);
assign n1163 = ~(n1422 | n148);
assign n1015 = ~(n1041 | n967);
assign n1516 = ~n47;
assign n394 = n413 | n513;
assign n1359 = ~(n198 | n1053);
assign n360 = ~(n1255 | n1251);
assign n1472 = ~n1408;
assign n936 = ~n51;
assign n1635 = ~(n915 ^ n1554);
assign n1447 = ~(n1127 ^ n742);
assign n402 = ~(n1255 | n209);
assign n1043 = n1629 | n1529;
assign n1294 = ~(n605 | n734);
assign n1282 = n1295 ^ n71;
assign n191 = n641 | n539;
assign n1033 = n1348 & n1535;
assign n667 = n1491 & n632;
assign n518 = ~n1365;
assign n1007 = n713 | n519;
assign n890 = n1517 | n1139;
assign n1491 = n275 | n277;
assign n71 = n975 & n570;
assign n28 = ~(n272 | n1283);
assign n1085 = n944 | n774;
assign n524 = n1629 | n1089;
assign n60 = ~n218;
assign n434 = ~n1587;
assign n151 = n917 | n783;
assign n822 = ~(n1133 | n931);
assign n1496 = n1242 ^ n1265;
assign n1010 = n954 & n938;
assign n610 = n1530 | n245;
assign n1229 = ~n729;
assign n720 = n940 | n841;
assign n1384 = ~n847;
assign n1320 = ~(n1311 | n1030);
assign n1190 = ~n770;
assign n1324 = ~n825;
assign n79 = n1495 | n1446;
assign n598 = n425 | n177;
assign n1619 = ~(n116 ^ n1669);
assign n506 = n1629 | n323;
assign n504 = ~n1624;
assign n981 = n1143 & n325;
assign n542 = ~(n402 | n1027);
assign n1272 = ~(n1274 | n1518);
assign n1609 = n243 | n28;
assign n949 = ~(n453 ^ n500);
assign n985 = ~(n300 | n1211);
assign n47 = n550 | n320;
assign n287 = n559 | n492;
assign n206 = ~(n289 | n62);
assign n163 = ~(n1554 ^ n1599);
assign n1344 = ~(n10 | n1478);
assign n862 = ~(n403 | n789);
assign n1428 = n224 & n514;
assign n1269 = ~n397;
assign n427 = n449 | n168;
assign n1593 = ~(n960 | n654);
assign n66 = ~n1290;
assign n57 = n707 & n877;
assign n1199 = ~n1356;
assign n1178 = ~(n622 | n677);
assign n140 = ~n1378;
assign n339 = ~(n1481 ^ n662);
assign n558 = ~n532;
assign n400 = ~n902;
assign n32 = ~(n1629 | n1323);
assign n1181 = ~n646;
assign n1368 = n1338 & n1354;
assign n87 = ~(n848 | n525);
assign n174 = ~n1435;
assign n260 = ~(n763 ^ n1058);
assign n725 = n922 | n1420;
assign n550 = ~(n1390 ^ n147);
assign n728 = ~(n615 | n1199);
assign n2 = ~n1108;
assign n761 = ~n1147;
assign n83 = n224 & n415;
assign n649 = ~n1384;
assign n1100 = n737 & n1243;
assign n927 = ~(n483 | n239);
assign n962 = ~n1235;
assign n1219 = n584 | n81;
assign n45 = ~(n135 | n385);
assign n286 = ~(n464 | n248);
assign n746 = ~(n121 ^ n600);
assign n540 = n929 & n1339;
assign n41 = n102 | n404;
assign n185 = n242 | n371;
assign n471 = ~(n1676 | n1195);
assign n1454 = ~(n1099 | n1499);
assign n227 = ~n1193;
assign n106 = n969 & n403;
assign n808 = n1180 | n1528;
assign n1647 = n1268 & n726;
assign n895 = ~(n950 | n644);
assign n543 = n1629 | n890;
assign n1626 = ~(n238 | n1143);
assign n72 = ~n956;
assign n534 = n658 | n849;
assign n370 = n1302 & n1379;
assign n754 = ~n196;
assign n1275 = n165 | n326;
assign n23 = n1465 & n751;
assign n343 = n1011 & n181;
assign n1371 = ~(n527 | n962);
assign n644 = ~(n1504 | n1248);
assign n1211 = ~n1457;
assign n1244 = ~n220;
assign n1246 = ~(n6 | n1272);
assign n1258 = ~(n120 | n930);
assign n854 = n331 | n104;
assign n517 = ~n121;
assign n1179 = ~(n42 | n1283);
assign n1417 = n839 | n1371;
assign n1322 = ~(n848 | n424);
assign n1060 = ~(n960 | n859);
assign n1604 = n1629 | n444;
assign n811 = n319 | n1543;
assign n1547 = ~n842;
assign n964 = ~n1520;
assign n1477 = ~n902;
assign n25 = n647 & n1;
assign n169 = ~(n256 | n1645);
assign n954 = n1320 | n1330;
assign n1191 = ~(n1524 ^ n1435);
assign n1153 = ~n877;
assign n187 = ~n297;
assign n695 = n401 & n1108;
assign n7 = n228 | n714;
assign n1419 = ~n1038;
assign n463 = ~n573;
assign n1476 = n1654 | n736;
assign n1316 = ~(n960 | n646);
assign n1617 = ~(n112 ^ n125);
assign n398 = ~n372;
assign n1250 = ~(n561 | n752);
assign n815 = n442 | n7;
assign n961 = ~(n454 ^ n594);
assign n1576 = n800 & n507;
assign n682 = n628 & n184;
assign n670 = ~n1336;
assign n913 = ~(n1255 | n1518);
assign n1046 = n540 | n1203;
assign n529 = ~(n1606 | n1181);
assign n1375 = n1629 | n1657;
assign n1416 = n1234 & n93;
assign n589 = n564 & n1378;
assign n270 = ~n514;
assign n1531 = n8 | n741;
assign n1657 = n82 | n1079;
assign n438 = ~n550;
assign n254 = n4 | n44;
assign n801 = ~n863;
assign n1140 = ~(n419 ^ n1634);
assign n531 = n135 & n325;
assign n495 = n1046 | n787;
assign n1095 = n943 | n724;
assign n1570 = n1215 | n864;
assign n688 = n1304 ^ n1564;
assign n333 = ~(n198 | n72);
assign n1307 = ~n393;
assign n1443 = ~(n1014 | n166);
assign n1631 = ~n523;
assign n1210 = n295 | n1185;
assign n839 = n1524 & n1479;
assign n747 = n1013 & n1606;
assign n836 = n984 | n1559;
assign n789 = ~(n772 | n1376);
assign n473 = n1334 | n169;
assign n1493 = ~n184;
assign n907 = ~(n694 | n590);
assign n880 = n1364 & n765;
assign n1437 = n68 | n1659;
assign n123 = n1140 & n632;
assign n810 = ~(n289 | n819);
assign n73 = ~(n1410 | n1404);
assign n1301 = ~(n198 | n1105);
assign n618 = ~n797;
assign n75 = ~n932;
assign n849 = n728 | n465;
assign n19 = ~(n706 | n1593);
assign n0 = ~n997;
assign n1397 = n433 | n1399;
assign n1565 = ~(n1367 | n261);
assign n1343 = n1335 | n162;
assign n1497 = ~(n1042 | n183);
assign n1018 = ~(n735 | n1039);
assign n1076 = ~(n870 ^ n1496);
assign n607 = ~(n1398 | n1560);
assign n805 = ~(n256 | n621);
assign n1129 = ~n573;
assign n844 = n118 | n698;
assign n872 = ~(n468 | n670);
assign n130 = ~n1360;
assign n24 = n1629 | n639;
assign n952 = n1124 | n200;
assign n65 = ~(n342 | n757);
assign n1583 = n1243 & n1253;
assign n733 = ~(n1 | n1632);
assign n1050 = n856 | n100;
assign n1499 = ~n1412;
assign n208 = ~(n198 | n1526);
assign n1651 = n1596 & n1606;
assign n1468 = ~(n221 | n1302);
assign n416 = ~n280;
assign n1214 = n874 | n1449;
assign n1012 = ~n517;
assign n500 = ~(n620 ^ n241);
assign n1313 = n1221 | n1625;
assign n1109 = ~(n1335 ^ n629);
assign n1613 = ~(n859 ^ n677);
assign n1394 = ~(n283 | n792);
assign n675 = ~n196;
assign n515 = ~(n1243 | n72);
assign n194 = n103 | n322;
assign n781 = ~n1587;
assign n965 = ~(n933 | n1156);
assign n112 = ~n975;
assign n1578 = ~n1405;
assign n1502 = n1140 | n318;
assign n1567 = ~(n615 | n1022);
assign n1224 = ~(n818 | n544);
assign n1257 = ~(n268 ^ n209);
assign n972 = n746 & n632;
assign n219 = n616 & n765;
assign n297 = n747 | n886;
assign n216 = n940 ^ n1329;
assign n1450 = n69 & n1243;
assign n327 = n156 & n145;
assign n81 = ~(n1227 | n291);
assign n387 = n1346 | n208;
assign n1273 = ~(n1511 | n959);
assign n717 = n1134;
assign n1217 = n579 & n1243;
assign n617 = n956 & n325;
assign n1288 = ~n625;
assign n226 = ~(n236 | n1251);
assign n930 = ~(n1308 ^ n835);
assign n1079 = n1238 | n5;
assign n1402 = ~n652;
assign n55 = ~n1251;
assign n1039 = ~n1440;
assign n846 = n1094 | n983;
assign n911 = ~(n361 ^ n1165);
assign n121 = ~(n1430 ^ n1389);
assign n1636 = ~n931;
assign n1466 = n267 | n1400;
assign n1188 = ~(n198 | n884);
assign n1020 = n407 & n632;
assign n1594 = n484 | n475;
assign n1632 = ~(n1463 ^ n1434);
assign n1287 = ~(n198 | n935);
assign n94 = ~n115;
assign n1107 = n1319 ^ n1264;
assign n1399 = ~(n735 | n964);
assign n1653 = n490 & n325;
assign n876 = ~(n843 | n1177);
assign n1369 = n1413 & n989;
assign n454 = ~(n1572 ^ n1591);
assign n887 = ~n1247;
assign n1629 = n1090;
assign n1434 = ~(n372 ^ n613);
assign n116 = ~(n161 ^ n625);
assign n401 = n1600 | n947;
assign n304 = ~n982;
assign n1204 = ~n306;
assign n464 = ~(n1255 | n135);
assign n111 = ~(n1398 | n665);
assign n888 = ~(n1425 | n999);
assign n1130 = n1481 | n1292;
assign n683 = n140 | n1416;
assign n1154 = n38 | n867;
assign n1483 = ~(n1635 ^ n1298);
assign n597 = n149 & n796;
assign n50 = n416 & n570;
assign n199 = n759 | n1359;
assign n1505 = ~(n882 | n1256);
assign n1510 = n1293 | n548;
assign n281 = ~(n367 | n52);
assign n165 = n1000 | n307;
assign n1427 = ~n507;
assign n1633 = ~(n1091 | n665);
assign n894 = n1629 | n472;
assign n714 = n1067 & n1520;
assign n1112 = ~(n897 | n971);
assign n1644 = n1143 & n230;
assign n1220 = n351 & n869;
assign n443 = ~(n738 ^ n1002);
assign n734 = ~n908;
assign n259 = ~n1615;
assign n486 = ~(n1667 | n686);
assign n1247 = ~n392;
assign n232 = n480;
assign n702 = ~(n1606 | n800);
assign n419 = ~(n625 ^ n403);
assign n1062 = ~n1432;
assign n580 = ~(n355 | n556);
assign n623 = n455 & n521;
assign n320 = ~n493;
assign n736 = n1007 | n1437;
assign n1135 = n997 & n1121;
assign n314 = n356 & n1243;
assign n467 = n1471 | n537;
assign n1618 = n481 & n1606;
assign n447 = ~(n451 | n316);
assign n1159 = ~n731;
assign n1507 = n1492 & n147;
assign n703 = ~(n882 | n394);
assign n445 = n176 & n950;
assign n1465 = ~n218;
assign n512 = ~n1409;
assign n560 = n1331 & n1243;
assign n309 = ~(n342 | n649);
assign n730 = n1470 & n1232;
assign n175 = ~(n304 | n863);
assign n698 = n681 | n131;
assign n906 = ~(n1311 | n135);
assign n1105 = ~n135;
assign n347 = n1629 | n1313;
assign n282 = ~(n643 ^ n1047);
assign n631 = ~(n1108 | n1077);
assign n759 = ~(n1311 | n646);
assign n545 = ~n1166;
assign n986 = ~(n272 | n210);
assign n834 = n416 & n94;
assign n1061 = ~(n1184 | n1650);
assign n85 = n1152 & n490;
assign n203 = n23 | n430;
assign n181 = n1357 | n70;
assign n1333 = ~n57;
assign n1557 = ~n621;
assign n1432 = ~n1173;
assign n788 = ~(n1047 ^ n1128);
assign n1540 = n1186 | n705;
assign n493 = n274 & n777;
assign n313 = n1629 | n1461;
assign n786 = n478;
assign n1340 = n171 | n764;
assign n1083 = n349 | n1344;
assign n484 = n1607 | n900;
assign n861 = ~n1342;
assign n4 = n373 & n1243;
assign n385 = ~n365;
assign n902 = ~n138;
assign n882 = ~n1290;
assign n1084 = ~(n1035 ^ n1619);
assign n99 = n1264 | n657;
assign n828 = n1289 | n978;
assign n275 = n968 & n1421;
assign n1292 = ~(n1242 | n600);
assign n168 = n1055 | n805;
assign n104 = n186 | n437;
assign n22 = n1382 & n1165;
assign n231 = n284 | n650;
assign n721 = n1226 | n1502;
assign n1654 = n749 | n538;
assign n1215 = ~(n1378 | n1527);
assign n966 = n271 | n216;
assign n582 = ~(n577 | n643);
assign n125 = ~n459;
assign n511 = ~(n1311 | n1518);
assign n946 = ~(n1146 | n130);
assign n141 = ~(n1627 ^ n376);
assign n825 = ~n1137;
assign n117 = n811 | n1284;
assign n150 = n1629 | n1154;
assign n706 = n654 & n325;
assign n884 = ~n209;
assign n1577 = n375 | n795;
assign n638 = ~(n1605 | n824);
assign n43 = ~n283;
assign n1185 = ~(n1058 | n385);
assign n753 = ~n419;
assign n431 = ~(n264 ^ n922);
assign n587 = ~(n1637 ^ n1045);
assign n93 = n1181 | n700;
assign n34 = ~n1436;
assign n1193 = n488 & n1551;
assign n382 = ~(n1621 | n860);
assign n1022 = ~n1336;
assign n35 = n578 | n571;
assign n183 = ~n701;
assign n684 = n965 | n143;
assign n1342 = ~n66;
assign n29 = ~(n1064 | n124);
assign n1148 = ~n1170;
assign n1088 = n1545 & n230;
assign n1519 = n1658 | n1590;
assign n444 = n651 | n976;
assign n1525 = n107 & n1243;
assign n396 = ~(n1361 | n1480);
assign n1347 = ~(n1309 | n1256);
assign n1453 = ~(n909 | n1031);
assign n1055 = ~(n1162 | n1480);
assign n1145 = ~(n1152 | n1547);
assign n864 = n199 & n1378;
assign n592 = n824 | n385;
assign n685 = n647 & n1555;
assign n100 = n1202 | n555;
assign n900 = ~(n1374 | n545);
assign n611 = ~n1647;
assign n823 = ~(n1430 ^ n361);
assign n1424 = ~(n605 | n959);
assign n352 = ~n824;
assign n255 = n1494 | n1048;
assign n261 = ~(n141 ^ n949);
assign n1658 = n1032 | n523;
assign n466 = ~n1592;
assign n91 = n122 & n1005;
assign n621 = n203 | n202;
assign n1283 = n916 | n593;
assign n991 = ~n692;
assign n21 = n473 | n1174;
assign n858 = n677 & n325;
assign n1514 = n1278 | n1612;
assign n516 = n1472 & n438;
assign n768 = ~(n1002 | n48);
assign n161 = n1381 & n1606;
assign n671 = ~n1335;
assign n300 = ~n1365;
assign n475 = n567 | n1468;
assign n655 = n448 | n13;
assign n242 = n395 & n1580;
assign n520 = n18 | n1595;
assign n1296 = n956 & n230;
assign n204 = n197 | n712;
assign n657 = n1319 | n854;
assign n1661 = n1489 | n1576;
assign n1356 = ~n611;
assign n110 = n1127 | n59;
assign n449 = n745 | n541;
assign n921 = ~(n927 ^ n672);
assign n1436 = ~n26;
assign n591 = n995 & n753;
assign n739 = ~(n1161 | n162);
assign n1386 = ~(n1255 | n956);
assign n277 = n577 & n1016;
assign n1524 = n39 | n515;
assign n54 = n1155 | n699;
assign n284 = n1443 | n382;
assign n331 = n1343 & n1315;
assign n496 = ~(n933 | n1544);
assign n748 = n467 | n1582;
assign n672 = ~(n1158 | n106);
assign n814 = n1214 | n666;
assign n1001 = ~n1173;
assign n791 = ~n962;
assign n250 = n1126 | n101;
assign n487 = ~(n1485 | n1560);
assign n1026 = n740;
assign n774 = ~(n861 | n1120);
assign n764 = ~(n504 | n1601);
assign n1248 = ~(n1605 | n209);
assign n1113 = ~(n1427 | n1058);
assign n126 = ~(n1146 | n1031);
assign n1408 = ~n35;
assign n1435 = n1217 | n108;
assign n1073 = n1369 & n1515;
assign n499 = n511 | n305;
assign n1103 = ~(n1024 | n336);
assign n18 = ~(n934 | n734);
assign n1350 = n278 | n1266;
assign n1500 = ~(n1391 | n682);
assign n298 = n191 | n583;
assign n172 = ~(n1629 | n1643);
assign n600 = n685 | n1270;
assign n1256 = n1431 | n547;
assign n1072 = ~(n582 ^ n788);
assign n408 = ~(n1372 ^ n426);
assign n1584 = ~(n956 | n344);
assign n1634 = n77 | n398;
assign n278 = n361 & n1165;
assign n410 = n832 & n654;
assign n1442 = n574;
assign n1364 = n1539 | n45;
assign n1535 = ~n1413;
assign n1090 = ~n1310;
assign n1537 = ~n899;
assign n1149 = ~n1243;
assign n461 = ~n31;
assign n850 = n1651 | n129;
assign n1387 = n251 & n576;
assign n180 = ~(n843 | n566);
assign n953 = ~(n152 | n754);
assign n910 = ~n1190;
assign n62 = ~n1403;
assign n779 = n71 | n50;
assign n146 = n1164 | n828;
assign n1492 = n601 | n508;
assign n873 = ~(n1016 | n1159);
assign n1586 = ~(n1511 | n1063);
assign n354 = n1368 & n1116;
assign n186 = ~n1372;
assign n1662 = ~(n1245 | n968);
assign n868 = ~n760;
assign n178 = ~(n1425 | n352);
assign n1489 = n629 & n325;
assign n1433 = n1647 & n1121;
assign n122 = n637 | n237;
assign n745 = ~(n9 | n227);
assign n1202 = ~(n1093 | n400);
assign n1169 = n1008 & n283;
assign n10 = ~n1033;
assign n636 = n708 | n1010;
assign n328 = ~(n557 ^ n1484);
assign n1183 = n1007 & n1005;
assign n115 = ~n1663;
assign n1132 = ~(n1388 | n566);
assign n578 = n414 & n938;
assign n1484 = ~(n554 ^ n1546);
assign n152 = ~n536;
assign n1031 = ~n1384;
assign n856 = n65 | n436;
assign n170 = n163 | n766;
assign n1319 = n626 | n1501;
assign n1315 = n671 | n832;
assign n1194 = n1629 | n1050;
assign n477 = n2 | n174;
assign n1209 = n1493 | n1419;
assign n1041 = ~(n1255 | n859);
assign n154 = n478;
assign n442 = n206 | n88;
assign n915 = ~n1548;
assign n963 = ~(n851 | n34);
assign n509 = ~n1406;
assign n1235 = n1205 | n516;
assign n238 = ~n507;
assign n302 = n1497 | n17;
assign n1671 = n423 | n1397;
assign n541 = ~(n285 | n1157);
assign n652 = n877 & n182;
assign n1589 = ~n889;
assign n1009 = ~(n1191 ^ n961);
assign n1558 = ~(n1309 | n1003);
assign n249 = n811 & n1005;
assign n1623 = ~(n222 | n218);
assign n1338 = n412 & n477;
assign n1411 = ~(n1614 ^ n260);
assign n393 = n235 & n84;
assign n809 = ~(n1255 | n646);
assign n1133 = n1417 & n1420;
assign n1192 = n1134;
assign n1554 = ~n366;
assign n1207 = ~n1534;
assign n1122 = n1510 | n1085;
assign n202 = n681 & n632;
assign n1252 = ~(n1451 | n1143);
assign n1117 = n110;
assign n1574 = ~(n96 & n1150);
assign n994 = ~n1033;
assign n755 = ~(n1467 | n11);
assign n430 = n1654 & n1005;
assign n1097 = n1503 & n1655;
assign n322 = ~(n897 | n640);
assign n735 = ~n1097;
assign n494 = ~n1624;
assign n879 = ~(n482 ^ n1257);
assign n1067 = ~n1448;
assign n680 = n327 | n338;
assign n1383 = ~(n1350 ^ n1447);
assign n1064 = n1573;
assign n1486 = n1267 | n29;
assign n863 = n1439 | n1325;
assign n1249 = ~(n765 | n286);
assign n1048 = ~(n329 | n535);
assign n92 = ~(n1274 | n135);
assign n892 = n1251 & n325;
assign n246 = ~(n1213 | n343);
assign n1317 = ~n1377;
assign n1628 = n167 & n794;
assign n1080 = ~(n1534 | n1636);
assign n738 = ~(n113 ^ n784);
assign n1231 = n1305 | n791;
assign n1119 = n491 & n1005;
assign n1023 = n1630;
assign n661 = n945 | n315;
assign n224 = n421 & n1412;
assign n1295 = n94 & n720;
assign n1225 = ~(n1523 | n1395);
assign n228 = ~(n1485 | n34);
assign n1314 = n1490 | n357;
assign n265 = n797 | n1244;
assign n1517 = n1273 | n1081;
assign n1008 = ~(n1660 ^ n1483);
assign n1541 = ~n495;
assign n1490 = n1118 | n1112;
assign n1268 = ~n84;
assign n573 = ~n1448;
assign n472 = n1212 | n1340;
assign n766 = n431 | n844;
assign n271 = ~(n113 ^ n16);
assign n519 = ~(n1108 | n1250);
assign n922 = ~n857;
assign n1201 = ~(n704 | n1269);
assign n458 = ~n859;
assign n1380 = ~(n870 ^ n339);
assign n1522 = ~(n493 | n35);
assign n190 = n761 | n99;
assign n919 = n1677 | n1423;
assign n335 = ~(n1098 | n1269);
assign n1068 = ~(n147 | n865);
assign n48 = n1338 & n1540;
assign n552 = ~(n386 | n130);
assign n1670 = n585 & n683;
assign n1494 = ~(n418 | n649);
assign n741 = n335 | n460;
assign n1672 = ~n590;
assign n425 = ~(n1366 | n218);
assign n58 = ~(n435 | n812);
assign n1302 = n912 | n177;
assign n223 = n1251 & n230;
assign n423 = n1322 | n866;
assign n1608 = ~n905;
assign n1308 = ~n75;
assign n1285 = ~n218;
assign n886 = n1675 & n1161;
assign n1334 = ~(n526 | n668);
assign n1156 = ~n939;
assign n1230 = ~n1402;
assign n1245 = ~n1351;
assign n1395 = n846 | n86;
assign n1005 = n1445;
assign n1488 = n68 & n1005;
assign n143 = ~(n1578 | n466);
assign n1357 = n517 & n30;
assign n109 = ~n1417;
assign n348 = n1551 & n1655;
assign n1421 = n1555 | n234;
assign n1546 = n560 | n1429;
assign n80 = ~(n1064 | n1652);
assign n762 = ~n1350;
assign n1506 = n487 | n266;
assign n1002 = n936 & n841;
assign n980 = ~n569;
assign n1242 = ~n225;
assign n479 = ~(n443 ^ n299);
assign n1649 = n153 | n1018;
assign n1392 = n288 | n337;
assign n390 = ~(n1024 | n1532);
assign n993 = n158 | n294;
assign n1173 = ~n1445;
assign n663 = n350;
assign n218 = n1362;
assign n1461 = n173 | n687;
assign n1234 = n646 | n1102;
assign n525 = ~n57;
assign n406 = ~n910;
assign n321 = ~n1044;
assign n162 = ~n1311;
assign n1600 = ~(n1311 | n1143);
assign n105 = ~n1406;
assign n366 = ~n1564;
assign n674 = ~n950;
assign n622 = ~n507;
assign n1625 = n1294 | n755;
assign n1139 = n1353 | n1037;
assign n778 = ~n1141;
assign n1643 = ~(n78 | n813);
assign n1284 = n122 | n748;
assign n1385 = n387 & n1530;
assign n1611 = ~(n1394 | n1169);
assign n1337 = ~n970;
assign n996 = ~n661;
assign n376 = ~(n811 ^ n1500);
assign n976 = n1567 | n447;
assign n441 = ~n750;
assign n1426 = ~(n238 | n956);
assign n947 = ~(n198 | n606);
assign n367 = ~(n769 | n1246);
assign n1568 = ~n138;
assign n258 = ~(n67 | n918);
assign n1605 = ~n507;
assign n1106 = ~n1300;
assign n480 = n132 & n742;
assign n1599 = n609 | n379;
assign n551 = ~(n1187 | n400);
assign n1512 = n194 | n257;
assign n1329 = ~(n51 | n768);
assign n139 = n1066 | n776;
assign n897 = ~n31;
assign n213 = ~(n1611 ^ n891);
assign n1665 = ~n1610;
assign n1464 = ~(n1091 | n406);
assign n1638 = n943 | n420;
assign n1552 = n478;
assign n1274 = ~n507;
assign n1429 = ~(n1243 | n352);
assign n1236 = ~(n631 | n695);
assign n214 = ~(n1676 | n1123);
assign n332 = ~(n198 | n977);
assign n523 = n512 | n405;
assign n1239 = n984 | n988;
assign n124 = ~(n1306 ^ n926);
assign n874 = ~(n793 | n311);
assign n565 = n1547;
assign n787 = n431 & n632;
assign n1376 = ~(n1425 | n935);
assign n318 = n746 | n312;
assign n306 = ~n1498;
assign n606 = ~n1143;
assign n319 = ~(n1240 | n709);
assign n59 = n932 | n1638;
assign n536 = ~n1307;
assign n134 = ~n251;
assign n351 = n1258 | n826;
assign n1656 = ~(n659 ^ n1616);
assign n630 = ~(n1425 | n72);
assign n1138 = n1629 | n1553;
assign n144 = n824 & n325;
assign n1197 = ~(n300 | n345);
assign n926 = n14 | n1473;
assign n20 = n661 ^ n1663;
assign n40 = ~(n1427 | n490);
assign n1011 = n70 | n600;
assign n1051 = n727 & n1606;
assign n1228 = ~(n913 | n888);
assign n1127 = ~n1297;
assign n1336 = ~n0;
assign n439 = ~(n956 ^ n1143);
assign n1374 = ~n1405;
assign n77 = n995 & n1555;
assign n1401 = ~(n596 | n525);
assign n1615 = ~n1333;
assign n1400 = n1656 | n721;
assign n210 = ~n212;
assign n33 = n770 & n1515;
assign n807 = ~(n1311 | n654);
assign n56 = n163 & n632;
assign n521 = n391 | n193;
assign n98 = ~(n1352 ^ n1370);
assign n1118 = ~(n1162 | n273);
assign n1452 = ~(n568 | n1507);
assign n378 = ~(n1621 | n722);
assign n632 = n771;
assign n614 = n991 | n1622;
assign n982 = n1513 | n1034;
assign n1650 = ~n939;
assign n1561 = ~(n1311 | n677);
assign n522 = n1260 | n333;
assign n1227 = ~n1318;
assign n1382 = n1521 | n942;
assign n310 = n609 | n264;
assign n1142 = n852 | n718;
assign n1167 = ~(n152 | n1355);
assign n1459 = n1428 & n1549;
assign n640 = ~n1059;
assign n200 = ~(n1667 | n562);
assign n397 = ~n134;
assign n875 = n669 | n1068;
assign n1645 = ~n980;
assign n1212 = n817 | n58;
assign n1019 = n1104 | n146;
assign n160 = ~(n1042 | n1261);
assign n1028 = ~(n1613 ^ n136);
assign n893 = ~n536;
assign n1115 = ~(n144 | n638);
assign n456 = n1487 | n411;
assign n719 = ~(n439 ^ n879);
assign n847 = ~n1647;
assign n955 = n27 | n1263;
assign n1205 = n1390 & n147;
assign n1471 = n151 & n950;
assign n1003 = ~n980;
assign n782 = n309 | n986;
assign n1328 = ~(n596 | n1004);
assign n1346 = ~(n1311 | n824);
assign n1669 = ~(n1144 ^ n1444);
assign n413 = n572 | n878;
assign n1175 = ~n229;
assign n1592 = ~n1029;
assign n303 = ~n262;
assign n253 = n481;
assign n860 = ~n1610;
assign n865 = ~(n360 | n830);
assign n173 = n946 | n1132;
assign n625 = n1051 | n831;
assign n240 = n1629 | n723;
assign n613 = ~(n659 ^ n1006);
assign n1172 = ~n1326;
assign n819 = ~n1377;
assign n503 = n610 & n79;
assign n294 = ~(n1102 | n1518);
assign n448 = n1455 & n664;
assign n374 = ~n652;
assign n470 = ~(n1456 | n725);
assign n590 = n655 | n80;
assign n6 = n1518 & n325;
assign n324 = n293;
assign n742 = ~n932;
assign n1640 = ~(n1441 ^ n1380);
assign n1601 = ~n1541;
assign n1372 = n799 | n739;
assign n1040 = n25 | n1270;
assign n37 = n458 | n700;
assign n694 = ~n1281;
assign n350 = ~n128;
assign n699 = n1491 | n1466;
assign n156 = ~n218;
assign n446 = ~n624;
assign n889 = ~n1355;
assign n1277 = n267 & n632;
assign n639 = n1609 | n520;
assign n1474 = n1629 | n1639;
assign n1610 = ~n345;
assign n407 = ~(n48 ^ n112);
assign n485 = ~n503;
assign n1237 = n673 & n37;
assign n870 = n30 ^ n1012;
assign n1641 = n223 | n226;
assign n650 = n1401 | n1505;
assign n369 = ~(n661 | n459);
assign n103 = ~(n1581 | n273);
assign n1504 = n209 & n325;
assign n817 = ~(n710 | n819);
assign n1571 = n552 | n308;
assign n821 = n1623 | n1486;
assign n1642 = n1453 | n876;
assign n612 = ~(n1056 | n1113);
assign n653 = n1526 | n700;
assign n1449 = ~(n1374 | n686);
assign n1034 = ~n597;
assign n775 = n1264 & n1005;
assign n958 = ~n730;
assign n666 = n214 | n937;
assign n420 = ~n647;
assign n1195 = ~n853;
assign n1668 = n251 & n1648;
assign n708 = ~(n938 | n188);
assign n1544 = ~n57;
assign n777 = ~n1563;
assign n555 = ~(n1129 | n392);
assign n1044 = ~n1333;
assign n999 = ~n1518;
assign n1158 = ~(n403 | n612);
assign n678 = n623;
assign n388 = n1013;
assign n392 = n36 | n56;
assign n114 = n807 | n410;
assign n248 = ~(n1425 | n1105);
assign n344 = ~n365;
assign n453 = ~(n1236 ^ n580);
assign n52 = n499 & n769;
assign n452 = n1586 | n1167;
assign n95 = ~(n1165 | n1458);
assign n39 = n1407 & n1243;
assign n207 = ~n348;
assign n31 = ~n1172;
assign n903 = ~(n531 | n92);
assign n795 = ~(n1324 | n624);
assign n102 = n1030 & n230;
assign n409 = n157 | n966;
assign n559 = n1285 & n1508;
assign n1213 = ~n730;
assign n1082 = ~(n470 | n1472);
assign n1241 = n407 | n409;
assign n3 = n1328 | n1197;
assign n603 = ~(n120 | n1661);
assign n831 = ~(n1606 | n935);
assign n562 = n595 | n1486;
assign n608 = n1596;
assign n450 = ~(n215 | n1060);
assign n1455 = ~n218;
assign n236 = ~n365;
assign n1096 = n979 | n1488;
assign n166 = ~n1230;
assign n1370 = ~(n921 ^ n408);
assign n840 = n1629 | n534;
assign n308 = ~(n10 | n345);
assign n428 = ~(n1425 | n1053);
assign n508 = ~(n198 | n55);
assign n1290 = n1153 & n182;
assign n643 = n589 | n1662;
assign n252 = ~(n1435 ^ n1108);
assign n1066 = n1460 & n1049;
assign n358 = ~n1001;
assign n983 = n796 & n589;
assign n1354 = n252 | n1171;
assign n1458 = ~(n1653 | n40);
assign n987 = n1223 & n1606;
assign n1004 = ~n868;
assign n1536 = ~n1432;
assign n838 = n1338 & n1663;
assign n1607 = ~(n1280 | n311);
assign n1520 = ~n394;
assign n604 = ~n509;
assign n707 = ~n182;
assign n241 = ~(n1452 ^ n636);
assign n1664 = ~(n1425 | n1545);
assign n855 = ~n1545;
assign n1444 = ~(n564 ^ n850);
assign n528 = ~(n1569 ^ n175);
assign n383 = n1387 | n1222;
assign n433 = ~(n1581 | n1123);
assign n148 = ~n306;
assign n830 = ~(n1425 | n55);
assign n530 = ~n229;
assign n790 = ~(n1562 & n128);
assign n539 = ~(n769 | n1228);
assign n1035 = n1447 ^ n823;
assign n1448 = ~n1379;
assign n760 = ~n1193;
assign n312 = n1229 | n970;
assign n42 = ~n1318;
assign n276 = n646 & n325;
assign n1588 = n452 | n1642;
assign n1174 = n1579 | n907;
assign n712 = n1069 | n377;
assign n1318 = ~n994;
assign n263 = ~(n622 | n1030);
assign n1196 = n1245 | n982;
assign n372 = n801 & n1196;
assign n457 = ~(n346 | n827);
assign n78 = n1433 | n1291;
assign n960 = ~n507;
assign n465 = ~(n604 | n316);
assign n1616 = n873 | n643;
assign n1456 = ~n274;
assign n363 = n808 | n1220;
assign n1286 = ~n1190;
assign n76 = n1629 | n1588;
assign n338 = n331 & n1005;
assign n243 = ~(n468 | n1317);
assign n359 = n1101 ^ n438;
assign n1591 = n1583 | n599;
assign n336 = ~n446;
assign n1332 = ~(n1617 ^ n20);
assign n1360 = ~n63;
assign n944 = ~(n1184 | n1544);
assign n553 = n271 & n632;
assign n391 = ~n1240;
assign n1420 = ~(n1572 ^ n950);
assign n1391 = ~(n184 | n450);
assign n197 = n802 | n1312;
assign n1550 = n160 | n119;
assign n1006 = ~(n1159 ^ n234);
assign n1087 = ~n293;
assign n951 = ~n446;
assign n462 = ~n252;
assign n435 = ~n105;
assign n1124 = ~(n923 | n374);
assign n53 = ~(n479 | n1368);
assign n414 = n314 | n211;
assign n1667 = ~n1300;
assign n568 = ~(n147 | n1136);
assign n1263 = ~(n494 | n887);
assign n1152 = ~n1606;
assign n866 = ~(n285 | n250);
assign n164 = ~(n617 | n1426);
assign n482 = ~(n1030 ^ n1251);
assign n584 = ~(n710 | n1022);
assign n1321 = ~(n654 ^ n490);
assign n878 = ~(n1062 | n503);
assign n266 = ~(n893 | n394);
assign n411 = ~(n1106 | n434);
assign n334 = ~(n329 | n1665);
assign n90 = ~(n1243 | n884);
assign n361 = n987 | n85;
assign n1451 = ~n365;
assign n179 = ~n705;
assign n280 = ~n48;
assign n1379 = n1535 & n989;
assign n1306 = ~(n733 | n1674);
assign n802 = ~(n362 | n321);
assign n257 = n87 | n703;
assign n74 = n744 | n1519;
assign n1673 = ~(n417 | n603);
assign n665 = ~n1568;
assign n279 = ~(n67 | n1004);
assign n323 = n1571 | n581;
assign n556 = n522 & n1479;
assign n992 = ~n149;
assign n269 = n456 | n767;
assign n127 = ~n1389;
assign n569 = n89 | n553;
assign n1024 = ~n1342;
assign n1585 = n1030 & n325;
assign n498 = ~(n290 | n1175);
assign n1513 = ~n1271;
assign n239 = ~(n198 | n855);
assign n1300 = ~n1172;
assign n633 = n3 | n1649;
assign n709 = ~(n858 | n1178);
assign n355 = ~(n1479 | n164);
assign n1467 = ~n393;
assign n833 = n1285 & n1131;
assign n1157 = ~n1233;
assign n1111 = ~(n1575 ^ n1161);
assign n368 = ~(n693 ^ n930);
assign n537 = ~(n950 | n542);
assign n679 = n1661 ^ n331;
assign n1222 = n1428 & n1052;
assign n998 = ~n1030;
assign n88 = ~(n1227 | n250);
assign n1533 = ~(n504 | n624);
assign n1089 = n634 | n255;
assign n792 = ~(n587 ^ n804);
assign n1029 = n139 | n317;
assign n1566 = n1633 | n1558;
assign n1102 = ~n365;
assign n563 = n471 | n486;
assign n1590 = ~n1411;
assign n1086 = ~n1606;
assign n436 = ~(n42 | n1345);
assign n1216 = n1078 | n575;
assign n235 = ~n726;
assign n852 = n648 & n635;
assign n1206 = ~(n1324 | n495);
assign n307 = ~(n1578 | n781);
assign n1144 = ~(n743 ^ n234);
assign n155 = n51 ^ n738;
assign n49 = n1025 & n1606;
assign n1639 = n1566 | n1083;
assign n17 = ~(n303 | n1355);
assign n225 = n127 | n384;
assign n340 = ~(n463 | n495);
assign n1358 = ~n403;
assign n1473 = n1040 & n1640;
assign n1092 = ~(n1462 | n1385);
assign n326 = n498 | n1666;
assign n1646 = ~n770;
assign n757 = ~n1360;
assign n1114 = n929 & n1475;
assign n975 = ~(n554 ^ n765);
assign n1289 = ~n676;
assign n237 = ~(n938 | n440);
assign n1603 = ~n1351;
assign n14 = ~(n1299 | n1040);
assign n984 = ~n1150;
assign n1622 = n429 | n1207;
assign n455 = n881 | n1349;
assign n681 = ~(n527 ^ n1231);
assign n691 = n619 | n15;
assign n743 = n798 | n1057;
assign n885 = n1460 & n1189;
assign n502 = ~(n463 | n951);
assign n732 = n1644 | n1252;
assign n570 = ~n996;
assign n11 = ~n1440;
assign n693 = ~n627;
assign n812 = n871 | n1277;
assign n1390 = n1450 | n1363;
assign n474 = ~(n435 | n469);
assign n959 = ~n1436;
assign n1462 = ~(n1530 | n1115);
assign n548 = ~(n461 | n244);
assign n669 = n1641 & n147;
assign n1164 = ~n1630;
assign n1293 = ~(n1361 | n374);
assign n136 = ~(n135 ^ n824);
assign n585 = n1378 | n1415;
assign n1309 = ~n1379;
assign n301 = ~n113;
assign n626 = ~(n1389 | n19);
assign n377 = ~(n461 | n590);
assign n1675 = ~n1606;
assign n1469 = n419 | n372;
assign n941 = n1455 & n716;
assign n1059 = ~n250;
assign n914 = n60 & n1620;
assign n1652 = ~(n1308 ^ n246);
assign n723 = n1182 | n1506;
assign n979 = n395 & n233;
assign n1569 = ~(n597 | n846);
assign n1457 = ~n316;
assign n776 = n191 & n1005;
assign n460 = ~(n974 | n1204);
assign n843 = ~n509;
assign n1415 = ~(n809 | n428);
assign n1171 = n43 | n217;
assign n129 = ~(n1606 | n999);
assign n978 = n74 | n1084;
assign n1120 = ~n1541;
assign n229 = ~n207;
assign n1063 = ~n910;
assign n620 = ~(n895 | n445);
assign n1057 = n1086 & n1575;
assign n581 = n1424 | n1347;
assign n288 = n258 | n1103;
assign n1081 = ~(n346 | n1589);
assign n1659 = n485 | n778;
assign n157 = ~(n125 ^ n779);
assign n648 = ~n218;
assign n1232 = n1148 | n1675;
assign n341 = ~(n1064 | n213);
assign n896 = ~(n1101 ^ n924);
assign n1077 = ~(n981 | n1626);
assign n705 = n922 | n1207;
assign n113 = ~(n254 ^ n1240);
assign n1298 = n1133 | n1080;
assign n554 = n1100 | n12;
assign n827 = n1096 | n1020;
assign n1126 = n833 | n775;
assign n977 = ~n859;
assign n1075 = ~(n1064 | n1337);
assign n940 = ~n1110;
assign n1341 = ~(n1070 | n1259);
assign n744 = ~n785;
assign n935 = ~n1058;
assign n763 = ~(n399 ^ n1111);
assign n770 = n726 & n84;
assign n557 = ~(n1038 ^ n254);
assign n645 = n216 & n632;
assign n1553 = n782 | n955;
assign n1621 = ~n1326;
assign n133 = ~n812;
assign n948 = ~n198;
assign n1351 = ~n187;
assign n908 = ~n1646;
assign n1078 = n60 & n1418;
assign n997 = n1348 & n1413;
assign n1094 = n850 & n769;
assign n533 = ~(n1608 | n827);
assign n426 = ~(n281 ^ n1570);
assign n1218 = ~(n1274 | n1251);
assign n1259 = ~n397;
assign n832 = ~n198;
assign n149 = n564 ^ n1378;
assign n217 = n915 | n47;
assign n957 = n586 | n219;
assign n251 = n1537 & n270;
assign n767 = n1224 | n533;
assign n379 = ~n725;
assign n1377 = ~n611;
assign n153 = ~(n1014 | n668);
assign n594 = ~(n414 ^ n1390);
assign n1501 = n114 & n1389;
assign n567 = ~(n923 | n530);
assign n5 = ~(n1129 | n928);
assign n1587 = ~n566;
assign n1233 = ~n1283;
assign n159 = ~(n1438 | n1204);
assign n1381 = ~n574;
assign n63 = ~n997;
assign n967 = ~(n1425 | n458);
assign n1141 = n389 & n1538;
assign n429 = n881 | n720;
assign n752 = ~(n1425 | n606);
assign n1221 = n898 | n334;
assign n697 = ~n1572;
assign n1186 = ~n692;
assign n799 = n1161 & n198;
assign n920 = ~n1302;
assign n311 = ~n1193;
assign n12 = ~(n1243 | n1105);
assign n1305 = n1516 & n857;
assign n711 = n551 | n340;
assign n205 = n1210 & n403;
assign n46 = ~n1670;
assign n883 = ~(n1386 | n630);
assign n256 = ~n825;
assign n1404 = ~n1247;
assign n492 = ~(n358 | n1141);
assign n177 = n1565 | n341;
assign n616 = n906 | n1301;
assign n641 = n993 & n769;
assign n690 = n1268 & n235;
assign n1027 = ~(n1425 | n884);
assign n912 = n901 & n1065;
assign n1021 = n476 | n1514;
assign n1299 = ~(n1383 ^ n1076);
assign n1365 = n488 & n1503;
assign n1074 = ~n1034;
assign n167 = ~n899;
assign n1254 = n696 & n393;
assign n292 = ~n1134;
assign n1539 = n135 & n230;
assign n171 = ~(n1187 | n189);
assign n399 = ~(n646 ^ n1518);
assign n658 = n501 | n1533;
assign n1125 = n545 & n1033;
assign n601 = ~(n1311 | n1251);
assign n1431 = n1168 | n1183;
assign n1367 = ~n1001;
assign n1053 = ~n646;
assign n1327 = ~(n1522 ^ n359);
assign n299 = ~(n1617 ^ n1282);
assign n1016 = ~n1555;
assign n295 = n1058 & n230;
assign n609 = ~n381;
assign n44 = n1149 & n677;
assign n1200 = ~n664;
assign n1265 = n762 & n730;
assign n1271 = ~(n161 ^ n1545);
assign n881 = ~n301;
assign n26 = ~n1369;
assign n796 = ~n659;
assign n676 = ~(n328 ^ n1009);
assign n1423 = ~(n1410 | n696);
assign n905 = ~n66;
assign n583 = n549 | n46;
assign n212 = ~n686;
assign n89 = n1114 | n249;
assign n272 = ~n105;
assign n510 = ~(n1255 | n824);
assign n898 = ~(n386 | n1199);
assign n264 = ~n1563;
assign n561 = ~(n1255 | n1143);
assign n1470 = n1606 | n671;
assign n662 = ~(n958 | n181);
assign n82 = n872 | n1179;
assign n1151 = n1577 | n803;
assign n316 = n680 | n1075;
assign n722 = ~n1457;
assign n1393 = ~(n1608 | n1262);
assign n195 = n648 & n1303;
assign n1226 = ~(n1271 ^ n1225);
assign n1538 = n1493 | n1237;
assign n497 = ~n994;
assign n651 = n963 | n502;
assign n929 = ~n218;
assign n1278 = ~(n330 | n1259);
assign n566 = n185 | n972;
assign n1203 = n467 & n1005;
assign n619 = n1061 | n247;
assign n349 = ~(n418 | n62);
assign n1627 = ~(n1092 ^ n957);
assign n1267 = ~(n1536 | n98);
assign n689 = n1135 | n1125;
assign n101 = ~(n1064 | n729);
assign n424 = ~n868;
assign n108 = ~(n1243 | n606);
assign n729 = ~(n911 ^ n1130);
assign n221 = ~n262;
assign n1137 = ~n1097;
assign n1560 = ~n1286;
assign n412 = n1186 | n109;
assign n749 = n353 & n1479;
assign n1660 = ~(n1327 ^ n546);
assign n628 = n1176 | n332;
assign n1579 = ~(n362 | n227);
assign n871 = n941 | n422;
assign n624 = n287 | n645;
assign n970 = ~(n1213 ^ n343);
assign n968 = ~n731;
assign n800 = ~n629;
assign n1559 = n1201 | n159;
assign n942 = n948 & n490;
assign n27 = ~(n1093 | n189);
assign n70 = ~n762;
assign n1503 = ~n1551;
assign n371 = n1319 & n1005;
assign n1345 = ~n212;
assign n451 = ~n497;
assign n68 = n880 | n1249;
assign n138 = ~n1369;
assign n417 = n1200 & n120;
assign n1478 = ~n1672;
assign n1595 = ~(n494 | n621);
assign n687 = n111 | n457;
assign n488 = ~n1655;
assign n599 = n1149 & n268;
assign n826 = n1652 & n120;
assign n1612 = ~(n990 | n148);
assign n1534 = ~n217;
assign n1180 = n1276 & n1396;
assign n1353 = ~(n909 | n670);
assign n924 = n179 | n1417;
assign n1264 = n95 | n22;
assign n637 = n41 & n938;
assign n274 = n414 ^ n938;
assign n1128 = ~(n613 ^ n528);
assign n1564 = ~n274;
assign n357 = n1602 | n390;
assign n647 = n591 & n1603;
assign n773 = ~n652;
assign n1410 = ~n905;
assign n659 = ~(n850 ^ n769);
assign n816 = ~(n793 | n259);
assign n527 = ~(n1524 ^ n1479);
assign n931 = n109 & n777;
assign n1260 = ~(n1311 | n956);
assign n1032 = n441 | n1087;
assign n853 = ~n1402;
assign n131 = n896 | n1241;
assign n571 = ~(n381 | n1456);
assign n1304 = ~n550;
assign n1556 = n829;
assign n575 = n875 & n1005;
assign n317 = n1656 & n632;
assign n234 = n297;
assign n1291 = n562 & n690;
assign n188 = ~(n1585 | n263);
assign n867 = n607 | n953;
assign n118 = ~(n1304 ^ n1082);
assign n1330 = ~(n198 | n998);
assign n1038 = n1017 | n602;
assign n1155 = ~n1652;
assign n939 = ~n760;
assign n1532 = ~n1557;
assign n1430 = n49 | n904;
assign n546 = ~(n756 ^ n310);
assign n51 = n1414 | n369;
assign n1527 = ~(n276 | n1316);
assign n692 = ~n252;
assign n64 = n952 | n919;
assign n1463 = ~(n282 ^ n1597);
assign n8 = ~n1150;
assign n1208 = ~(n1311 | n1058);
assign n1674 = n1072 & n1;
assign n1182 = n810 | n474;
assign n285 = ~n1281;
assign n440 = ~(n806 | n1598);
assign n899 = ~n224;
assign n1406 = ~n690;
assign n937 = ~(n221 | n392);
assign n501 = ~(n851 | n406);
assign n1414 = n1546 & n1530;
assign n1348 = ~n989;
assign n247 = ~(n694 | n812);
assign n820 = n784 | n936;
assign n1323 = ~(n689 | n505);
assign n538 = ~(n1479 | n883);
assign n627 = ~n1155;
assign n1355 = n1216 | n201;
assign n673 = n859 | n1451;
assign n15 = n396 | n1206;
assign n668 = ~n348;
assign n1177 = ~n1592;
assign n758 = n816 | n73;
assign n346 = ~n1067;
assign n1677 = ~(n1280 | n259);
assign n1325 = n846 & n1271;
assign n1403 = ~n63;
assign n1352 = ~(n679 ^ n1107);
assign n61 = n845;
assign n1446 = n592 & n653;
assign n544 = ~n1044;
assign n273 = ~n853;
assign n564 = n1618 | n529;
assign n602 = ~(n1243 | n977);
assign n547 = n896 & n632;
assign n798 = n1606 & n588;
assign n489 = n350;
assign n196 = ~n827;
assign n1110 = ~n784;
assign n642 = n549 & n1005;
assign n784 = ~(n1038 ^ n184);
assign n1045 = ~(n381 ^ n1235);
assign n395 = ~n218;
assign n813 = n33 | n1254;
assign n1297 = ~n958;
assign n1498 = ~n1428;
assign n549 = n1088 | n1664;
assign n1526 = ~n824;
assign n30 = ~n911;
assign n1326 = n707 & n1153;
assign n337 = n1509 | n378;
assign n785 = ~(n1028 ^ n719);
assign n505 = n1073 | n370;
assign n211 = ~(n1243 | n998);
assign n731 = ~n992;
assign n783 = ~(n236 | n209);
assign n780 = n1561 | n1279;
assign n1136 = ~(n892 | n1218);
assign n928 = ~n1557;
assign n595 = n837 & n1065;
assign n1047 = ~(n1513 ^ n753);
assign n384 = ~n1430;
assign n1168 = n1465 & n432;
assign n841 = n975 | n459;
assign n925 = n991 ^ n1548;
assign n291 = ~n133;
assign n353 = n1296 | n1584;
assign n995 = ~n982;
assign n1509 = ~(n1373 | n773);
assign n513 = n157 & n632;
assign n1521 = ~(n1311 | n490);
assign n1460 = ~n218;
assign n724 = n1469 & n1054;
assign n686 = n1142 | n667;
assign n158 = n1518 & n230;
assign n1000 = ~(n818 | n1650);
assign n1270 = ~n724;
assign n16 = ~(n1295 | n834);
assign n1597 = ~(n1395 ^ n234);
assign n315 = ~n554;
assign n1637 = ~(n35 ^ n925);
assign n1388 = ~n497;
assign n38 = n126 | n180;
assign n1279 = n948 & n677;
assign n215 = n859 & n325;
assign n1495 = ~n1530;
assign n459 = ~(n1546 ^ n1530);
assign n380 = n496 | n1393;
assign n1054 = n1358 | n1288;
assign n660 = ~(n1311 | n209);
assign n1666 = ~(n303 | n675);
assign n1104 = ~n829;
assign n1363 = ~(n1243 | n55);
assign n305 = ~(n198 | n999);
assign n1528 = ~(n869 | n1673);
assign n1523 = n1074 & n1555;
assign n176 = n660 | n1188;
assign n1101 = ~n462;
assign n943 = ~n1357;
assign n405 = ~n296;
assign n577 = n149 & n1603;
assign n904 = n1086 & n654;
assign n1482 = ~n1420;
assign n404 = ~(n1030 | n344);
assign n772 = ~(n1255 | n1058);
assign n1312 = ~(n861 | n569);
assign n1542 = n750;
assign n845 = ~n128;
assign n917 = n209 & n230;
assign n945 = ~n765;
assign n1543 = n780 & n1240;
assign n1116 = ~(n155 ^ n1332);
assign n1563 = ~n1482;
assign n1614 = ~(n1109 ^ n1321);
assign n535 = ~n1672;
assign n192 = ~(n1467 | n569);
assign n1056 = n1058 & n325;
assign n1624 = ~n1307;
assign n572 = n156 & n973;
assign n142 = n614;
assign n1266 = ~(n225 | n911);
assign n696 = ~n920;
assign n969 = n1208 | n1287;
assign n193 = ~n254;
assign n656 = ~n1084;
assign n918 = ~n1615;
assign n36 = n195 | n91;
assign n1017 = n137 & n1243;
assign n1598 = ~(n1425 | n998);
assign n916 = n642 | n885;
assign n1445 = n1071 & n558;
assign n932 = n1145 | n702;
assign n1176 = ~(n1311 | n859);
assign n1166 = ~n562;
assign n1573 = n1065 | n558;
assign n1071 = ~n1065;
assign n1405 = ~n518;
assign n469 = ~n1059;
assign n1572 = n1525 | n90;
assign n1238 = ~(n934 | n1477);
assign n1349 = n1295 | n838;
assign n1198 = n302 | n684;
assign n345 = n715 | n123;
assign n715 = n914 | n1119;
assign n1481 = n1012 & n225;
assign n1160 = n1629 | n815;
assign n804 = ~(n822 ^ n688);
assign n1441 = ~(n1447 ^ n181);
assign n756 = ~(n1516 | n791);
assign n1069 = ~(n526 | n773);
assign n1147 = ~n1661;
assign n1362 = n532 | n1071;
assign n329 = ~n690;
assign n86 = n597 & n234;
assign n1582 = n875 | n1476;
assign n1602 = ~(n9 | n544);
assign n1281 = ~n518;
assign n132 = n1095 & n1265;
assign n267 = ~(n234 ^ n1555);
assign n593 = n1226 & n632;
assign n771 = ~n1573;
assign n1440 = ~n1256;
assign n189 = ~n908;
assign n262 = ~n1137;
assign n740 = n1668 | n1459;
assign n483 = n855 & n325;
assign n491 = n205 | n862;
assign n586 = ~(n765 | n903);
assign n1036 = n563 | n758;
assign n1261 = ~n1230;
assign n244 = ~n133;
assign n97 = n380 | n1550;
assign n375 = ~(n1373 | n530);
assign n1663 = n820 & n1209;
assign n364 = n842;
assign n1548 = ~n527;
assign n634 = n1464 | n192;
assign n1480 = ~n701;
assign n891 = n354 | n53;
assign n13 = n761 & n1005;
assign n713 = n732 & n1108;
assign n422 = ~(n1536 | n1372);
assign n119 = ~(n1106 | n1029);
assign n1123 = ~n348;
assign n389 = n184 | n1015;
assign n803 = n279 | n985;
assign n1529 = n1219 | n711;
assign n476 = ~n1150;
assign n971 = ~n1233;
assign n1037 = ~(n1388 | n1029);
assign n701 = ~n207;
assign n1439 = ~(n855 | n161);
assign n381 = n674 | n697;
assign n988 = n1341 | n1163;
assign n718 = ~(n1367 | n1670);
assign n1262 = ~n889;
assign n201 = n118 & n632;
assign n1487 = ~(n290 | n166);
assign n700 = ~n230;
assign n437 = n491 | n298;
assign n245 = ~(n510 | n178);
endmodule
