module top( 1_n1 , 1_n3 , 1_n4 , 1_n15 , 1_n21 , 1_n23 , 1_n28 , 1_n32 , 1_n37 , 1_n38 , 1_n40 , 1_n45 , 1_n47 , 1_n50 , 1_n52 , 1_n53 , 1_n54 , 1_n60 , 1_n72 , 1_n75 , 1_n79 , 1_n81 , 1_n83 , 1_n86 , 1_n87 , 1_n91 , 1_n95 , 1_n97 , 1_n99 , 1_n105 , 1_n111 , 1_n114 , 1_n117 , 1_n122 , 1_n139 , 1_n152 , 1_n154 , 1_n155 , 1_n160 , 1_n162 , 1_n168 , 1_n176 , 1_n183 , 1_n185 , 1_n187 , 1_n191 , 1_n194 , 1_n197 , 1_n198 , 1_n200 , 1_n205 , 1_n206 , 1_n208 , 1_n211 , 1_n214 , 1_n215 , 1_n218 , 1_n220 , 1_n227 , 1_n228 , 1_n231 , 1_n242 , 1_n243 , 1_n248 , 1_n254 , 1_n262 , 1_n265 , 1_n269 , 1_n273 , 1_n276 , 1_n278 , 1_n280 , 1_n283 );
    input 1_n1 , 1_n4 , 1_n15 , 1_n21 , 1_n23 , 1_n28 , 1_n37 , 1_n38 , 1_n45 , 1_n52 , 1_n53 , 1_n60 , 1_n75 , 1_n79 , 1_n83 , 1_n87 , 1_n95 , 1_n105 , 1_n114 , 1_n117 , 1_n122 , 1_n152 , 1_n155 , 1_n160 , 1_n162 , 1_n168 , 1_n183 , 1_n187 , 1_n194 , 1_n198 , 1_n206 , 1_n215 , 1_n218 , 1_n227 , 1_n228 , 1_n231 , 1_n242 , 1_n269 , 1_n276 , 1_n278 , 1_n280 ;
    output 1_n3 , 1_n32 , 1_n40 , 1_n47 , 1_n50 , 1_n54 , 1_n72 , 1_n81 , 1_n86 , 1_n91 , 1_n97 , 1_n99 , 1_n111 , 1_n139 , 1_n154 , 1_n176 , 1_n185 , 1_n191 , 1_n197 , 1_n200 , 1_n205 , 1_n208 , 1_n211 , 1_n214 , 1_n220 , 1_n243 , 1_n248 , 1_n254 , 1_n262 , 1_n265 , 1_n273 , 1_n283 ;
    wire 1_n0 , 1_n2 , 1_n5 , 1_n6 , 1_n7 , 1_n8 , 1_n9 , 1_n10 , 1_n11 , 1_n12 , 1_n13 , 1_n14 , 1_n16 , 1_n17 , 1_n18 , 1_n19 , 1_n20 , 1_n22 , 1_n24 , 1_n25 , 1_n26 , 1_n27 , 1_n29 , 1_n30 , 1_n31 , 1_n33 , 1_n34 , 1_n35 , 1_n36 , 1_n39 , 1_n41 , 1_n42 , 1_n43 , 1_n44 , 1_n46 , 1_n48 , 1_n49 , 1_n51 , 1_n55 , 1_n56 , 1_n57 , 1_n58 , 1_n59 , 1_n61 , 1_n62 , 1_n63 , 1_n64 , 1_n65 , 1_n66 , 1_n67 , 1_n68 , 1_n69 , 1_n70 , 1_n71 , 1_n73 , 1_n74 , 1_n76 , 1_n77 , 1_n78 , 1_n80 , 1_n82 , 1_n84 , 1_n85 , 1_n88 , 1_n89 , 1_n90 , 1_n92 , 1_n93 , 1_n94 , 1_n96 , 1_n98 , 1_n100 , 1_n101 , 1_n102 , 1_n103 , 1_n104 , 1_n106 , 1_n107 , 1_n108 , 1_n109 , 1_n110 , 1_n112 , 1_n113 , 1_n115 , 1_n116 , 1_n118 , 1_n119 , 1_n120 , 1_n121 , 1_n123 , 1_n124 , 1_n125 , 1_n126 , 1_n127 , 1_n128 , 1_n129 , 1_n130 , 1_n131 , 1_n132 , 1_n133 , 1_n134 , 1_n135 , 1_n136 , 1_n137 , 1_n138 , 1_n140 , 1_n141 , 1_n142 , 1_n143 , 1_n144 , 1_n145 , 1_n146 , 1_n147 , 1_n148 , 1_n149 , 1_n150 , 1_n151 , 1_n153 , 1_n156 , 1_n157 , 1_n158 , 1_n159 , 1_n161 , 1_n163 , 1_n164 , 1_n165 , 1_n166 , 1_n167 , 1_n169 , 1_n170 , 1_n171 , 1_n172 , 1_n173 , 1_n174 , 1_n175 , 1_n177 , 1_n178 , 1_n179 , 1_n180 , 1_n181 , 1_n182 , 1_n184 , 1_n186 , 1_n188 , 1_n189 , 1_n190 , 1_n192 , 1_n193 , 1_n195 , 1_n196 , 1_n199 , 1_n201 , 1_n202 , 1_n203 , 1_n204 , 1_n207 , 1_n209 , 1_n210 , 1_n212 , 1_n213 , 1_n216 , 1_n217 , 1_n219 , 1_n221 , 1_n222 , 1_n223 , 1_n224 , 1_n225 , 1_n226 , 1_n229 , 1_n230 , 1_n232 , 1_n233 , 1_n234 , 1_n235 , 1_n236 , 1_n237 , 1_n238 , 1_n239 , 1_n240 , 1_n241 , 1_n244 , 1_n245 , 1_n246 , 1_n247 , 1_n249 , 1_n250 , 1_n251 , 1_n252 , 1_n253 , 1_n255 , 1_n256 , 1_n257 , 1_n258 , 1_n259 , 1_n260 , 1_n261 , 1_n263 , 1_n264 , 1_n266 , 1_n267 , 1_n268 , 1_n270 , 1_n271 , 1_n272 , 1_n274 , 1_n275 , 1_n277 , 1_n279 , 1_n281 , 1_n282 , 1_n284 , 1_n285 ;
assign 1_n140 = 1_n247 & 1_n201;
assign 1_n72 = ~(1_n126 ^ 1_n162);
assign 1_n244 = 1_n173 | 1_n230;
assign 1_n18 = 1_n141 | 1_n136;
assign 1_n43 = ~1_n4;
assign 1_n177 = ~1_n198;
assign 1_n16 = ~(1_n215 ^ 1_n206);
assign 1_n80 = 1_n237 | 1_n252;
assign 1_n81 = ~(1_n216 ^ 1_n194);
assign 1_n261 = ~1_n193;
assign 1_n55 = ~1_n172;
assign 1_n148 = ~1_n168;
assign 1_n136 = ~(1_n209 ^ 1_n77);
assign 1_n263 = ~(1_n206 ^ 1_n183);
assign 1_n257 = ~(1_n280 ^ 1_n21);
assign 1_n159 = ~(1_n285 ^ 1_n24);
assign 1_n254 = 1_n0 ^ 1_n28;
assign 1_n33 = 1_n115 | 1_n256;
assign 1_n110 = 1_n55 | 1_n18;
assign 1_n68 = ~(1_n227 ^ 1_n21);
assign 1_n181 = ~(1_n187 ^ 1_n45);
assign 1_n49 = ~1_n26;
assign 1_n126 = 1_n90 | 1_n235;
assign 1_n225 = ~1_n12;
assign 1_n202 = 1_n103 | 1_n235;
assign 1_n200 = ~(1_n186 ^ 1_n23);
assign 1_n30 = 1_n78 | 1_n101;
assign 1_n123 = ~1_n137;
assign 1_n281 = 1_n193 | 1_n169;
assign 1_n50 = ~(1_n179 ^ 1_n87);
assign 1_n164 = ~(1_n28 ^ 1_n15);
assign 1_n47 = 1_n272 ^ 1_n38;
assign 1_n137 = ~1_n35;
assign 1_n27 = 1_n142 | 1_n5;
assign 1_n175 = ~1_n128;
assign 1_n277 = 1_n223 | 1_n108;
assign 1_n149 = 1_n2 & 1_n240;
assign 1_n213 = ~(1_n89 ^ 1_n165);
assign 1_n66 = ~1_n275;
assign 1_n103 = ~1_n224;
assign 1_n190 = 1_n226 | 1_n281;
assign 1_n115 = ~1_n224;
assign 1_n42 = 1_n137 | 1_n222;
assign 1_n56 = ~1_n114;
assign 1_n283 = ~(1_n48 ^ 1_n105);
assign 1_n259 = 1_n59 | 1_n43;
assign 1_n48 = 1_n195 | 1_n157;
assign 1_n11 = ~1_n199;
assign 1_n104 = 1_n7 | 1_n232;
assign 1_n209 = ~(1_n170 ^ 1_n188);
assign 1_n78 = ~1_n250;
assign 1_n174 = 1_n55 | 1_n150;
assign 1_n239 = ~1_n2;
assign 1_n176 = ~(1_n33 ^ 1_n95);
assign 1_n17 = 1_n173 | 1_n235;
assign 1_n219 = ~(1_n112 ^ 1_n16);
assign 1_n249 = ~1_n60;
assign 1_n40 = ~(1_n147 ^ 1_n183);
assign 1_n134 = 1_n203 | 1_n43;
assign 1_n274 = 1_n65 & 1_n239;
assign 1_n41 = 1_n107 | 1_n266;
assign 1_n236 = ~(1_n228 ^ 1_n95);
assign 1_n77 = ~(1_n279 ^ 1_n258);
assign 1_n119 = 1_n49 | 1_n88;
assign 1_n74 = ~(1_n278 ^ 1_n52);
assign 1_n270 = 1_n161 & 1_n7;
assign 1_n163 = 1_n78 | 1_n19;
assign 1_n100 = ~(1_n82 ^ 1_n74);
assign 1_n284 = ~(1_n271 ^ 1_n20);
assign 1_n241 = ~(1_n75 ^ 1_n45);
assign 1_n131 = 1_n249 | 1_n127;
assign 1_n97 = ~(1_n27 ^ 1_n53);
assign 1_n94 = ~(1_n138 ^ 1_n212);
assign 1_n54 = ~(1_n124 ^ 1_n160);
assign 1_n224 = ~1_n104;
assign 1_n237 = ~1_n149;
assign 1_n31 = ~(1_n152 ^ 1_n280);
assign 1_n203 = ~1_n218;
assign 1_n165 = ~(1_n152 ^ 1_n227);
assign 1_n129 = ~(1_n237 | 1_n190);
assign 1_n193 = ~(1_n71 ^ 1_n62);
assign 1_n166 = ~1_n26;
assign 1_n256 = ~1_n247;
assign 1_n107 = ~1_n136;
assign 1_n144 = 1_n166 | 1_n163;
assign 1_n2 = ~(1_n245 ^ 1_n217);
assign 1_n240 = ~1_n65;
assign 1_n153 = ~(1_n276 ^ 1_n95);
assign 1_n111 = ~(1_n264 ^ 1_n83);
assign 1_n268 = 1_n173 | 1_n36;
assign 1_n29 = ~(1_n28 ^ 1_n1);
assign 1_n125 = ~(1_n8 ^ 1_n31);
assign 1_n51 = 1_n180 | 1_n196;
assign 1_n272 = ~(1_n182 | 1_n190);
assign 1_n19 = 1_n121 | 1_n260;
assign 1_n141 = ~1_n266;
assign 1_n118 = ~1_n210;
assign 1_n5 = 1_n252 | 1_n275;
assign 1_n212 = ~(1_n23 ^ 1_n83);
assign 1_n179 = 1_n115 | 1_n230;
assign 1_n88 = 1_n174 | 1_n196;
assign 1_n245 = ~(1_n9 ^ 1_n68);
assign 1_n91 = ~(1_n119 ^ 1_n152);
assign 1_n92 = 1_n26 & 1_n46;
assign 1_n71 = ~(1_n8 ^ 1_n178);
assign 1_n26 = 1_n6 & 1_n35;
assign 1_n82 = ~(1_n242 ^ 1_n87);
assign 1_n143 = 1_n226 | 1_n36;
assign 1_n20 = ~(1_n219 ^ 1_n134);
assign 1_n170 = ~(1_n167 ^ 1_n257);
assign 1_n196 = 1_n261 | 1_n96;
assign 1_n169 = 1_n192 | 1_n123;
assign 1_n7 = ~1_n225;
assign 1_n172 = ~1_n58;
assign 1_n204 = ~(1_n135 ^ 1_n73);
assign 1_n246 = 1_n169 | 1_n19;
assign 1_n161 = ~1_n41;
assign 1_n147 = 1_n260 | 1_n143;
assign 1_n69 = ~1_n210;
assign 1_n138 = ~(1_n53 ^ 1_n155);
assign 1_n130 = 1_n103 | 1_n282;
assign 1_n265 = 1_n238 ^ 1_n79;
assign 1_n262 = 1_n129 ^ 1_n1;
assign 1_n90 = ~1_n270;
assign 1_n3 = ~(1_n130 ^ 1_n278);
assign 1_n22 = ~(1_n100 ^ 1_n263);
assign 1_n234 = ~(1_n83 ^ 1_n52);
assign 1_n145 = 1_n275 | 1_n19;
assign 1_n208 = ~(1_n63 ^ 1_n52);
assign 1_n184 = 1_n177 | 1_n108;
assign 1_n73 = 1_n148 | 1_n127;
assign 1_n207 = ~(1_n105 ^ 1_n194);
assign 1_n98 = ~(1_n1 ^ 1_n38);
assign 1_n135 = ~(1_n153 ^ 1_n102);
assign 1_n217 = ~(1_n234 ^ 1_n76);
assign 1_n85 = ~(1_n162 ^ 1_n183);
assign 1_n93 = 1_n180 | 1_n101;
assign 1_n112 = ~(1_n122 ^ 1_n187);
assign 1_n267 = 1_n69 | 1_n80;
assign 1_n157 = 1_n128 | 1_n174;
assign 1_n106 = 1_n56 | 1_n221;
assign 1_n271 = ~(1_n23 ^ 1_n278);
assign 1_n199 = 1_n92 & 1_n149;
assign 1_n84 = 1_n173 | 1_n80;
assign 1_n142 = ~1_n158;
assign 1_n61 = 1_n222 | 1_n123;
assign 1_n191 = ~(1_n133 ^ 1_n215);
assign 1_n101 = ~1_n92;
assign 1_n158 = ~1_n233;
assign 1_n243 = ~(1_n202 ^ 1_n45);
assign 1_n222 = ~1_n192;
assign 1_n235 = 1_n182 | 1_n128;
assign 1_n279 = ~(1_n79 ^ 1_n276);
assign 1_n230 = 1_n142 | 1_n281;
assign 1_n201 = ~1_n110;
assign 1_n12 = ~(1_n116 ^ 1_n151);
assign 1_n156 = ~1_n231;
assign 1_n260 = ~1_n274;
assign 1_n180 = ~1_n66;
assign 1_n24 = ~(1_n9 ^ 1_n277);
assign 1_n197 = ~(1_n44 ^ 1_n242);
assign 1_n39 = ~(1_n170 ^ 1_n259);
assign 1_n57 = ~(1_n98 ^ 1_n39);
assign 1_n109 = ~(1_n213 ^ 1_n184);
assign 1_n133 = 1_n90 | 1_n80;
assign 1_n25 = 1_n156 | 1_n221;
assign 1_n238 = 1_n199 & 1_n201;
assign 1_n250 = ~1_n174;
assign 1_n8 = ~(1_n13 ^ 1_n29);
assign 1_n89 = ~(1_n105 ^ 1_n160);
assign 1_n275 = 1_n12 | 1_n41;
assign 1_n96 = ~1_n149;
assign 1_n178 = ~(1_n160 ^ 1_n37);
assign 1_n285 = ~(1_n53 ^ 1_n242);
assign 1_n233 = 1_n240 | 1_n239;
assign 1_n9 = ~(1_n241 ^ 1_n85);
assign 1_n210 = ~1_n104;
assign 1_n70 = ~1_n233;
assign 1_n221 = ~1_n4;
assign 1_n132 = 1_n118 | 1_n11;
assign 1_n226 = 1_n58 | 1_n232;
assign 1_n58 = ~1_n12;
assign 1_n151 = ~(1_n236 ^ 1_n10);
assign 1_n128 = 1_n121 | 1_n42;
assign 1_n186 = 1_n166 | 1_n51;
assign 1_n59 = ~1_n269;
assign 1_n86 = ~(1_n244 ^ 1_n37);
assign 1_n171 = ~(1_n155 ^ 1_n87);
assign 1_n62 = ~(1_n171 ^ 1_n204);
assign 1_n6 = ~(1_n146 ^ 1_n159);
assign 1_n223 = ~1_n117;
assign 1_n264 = 1_n49 | 1_n145;
assign 1_n113 = ~(1_n215 ^ 1_n162);
assign 1_n167 = ~(1_n194 ^ 1_n37);
assign 1_n127 = ~1_n4;
assign 1_n258 = ~(1_n213 ^ 1_n131);
assign 1_n13 = ~(1_n79 ^ 1_n228);
assign 1_n108 = ~1_n4;
assign 1_n139 = 1_n189 ^ 1_n155;
assign 1_n220 = ~(1_n144 ^ 1_n227);
assign 1_n44 = 1_n195 | 1_n251;
assign 1_n65 = ~(1_n125 ^ 1_n284);
assign 1_n247 = 1_n92 & 1_n274;
assign 1_n102 = ~(1_n15 ^ 1_n38);
assign 1_n252 = ~1_n175;
assign 1_n255 = ~(1_n94 ^ 1_n113);
assign 1_n150 = 1_n136 | 1_n266;
assign 1_n229 = ~1_n70;
assign 1_n0 = 1_n199 & 1_n270;
assign 1_n182 = ~1_n274;
assign 1_n67 = ~(1_n164 ^ 1_n109);
assign 1_n173 = 1_n110;
assign 1_n214 = ~(1_n267 ^ 1_n187);
assign 1_n121 = ~1_n34;
assign 1_n188 = ~(1_n122 ^ 1_n75);
assign 1_n116 = ~(1_n100 ^ 1_n181);
assign 1_n216 = 1_n229 | 1_n268;
assign 1_n14 = 1_n173 | 1_n282;
assign 1_n192 = ~1_n6;
assign 1_n146 = ~(1_n219 ^ 1_n207);
assign 1_n36 = 1_n261 | 1_n61;
assign 1_n154 = ~(1_n64 ^ 1_n206);
assign 1_n120 = 1_n247 & 1_n270;
assign 1_n32 = ~(1_n132 ^ 1_n228);
assign 1_n189 = ~(1_n233 | 1_n93);
assign 1_n205 = ~(1_n253 ^ 1_n21);
assign 1_n266 = ~(1_n255 ^ 1_n67);
assign 1_n35 = ~(1_n22 ^ 1_n57);
assign 1_n185 = 1_n140 ^ 1_n276;
assign 1_n211 = ~(1_n84 ^ 1_n122);
assign 1_n46 = ~1_n193;
assign 1_n64 = 1_n96 | 1_n143;
assign 1_n253 = 1_n173 | 1_n246;
assign 1_n195 = ~1_n158;
assign 1_n34 = ~1_n46;
assign 1_n124 = 1_n229 | 1_n30;
assign 1_n232 = 1_n107 | 1_n141;
assign 1_n10 = ~(1_n94 ^ 1_n106);
assign 1_n63 = 1_n69 | 1_n246;
assign 1_n273 = ~(1_n17 ^ 1_n75);
assign 1_n251 = 1_n36 | 1_n118;
assign 1_n248 = 1_n120 ^ 1_n15;
assign 1_n76 = ~(1_n135 ^ 1_n25);
assign 1_n282 = 1_n169 | 1_n196;
assign 1_n99 = ~(1_n14 ^ 1_n280);
endmodule
