module top(in1, in2, in3, in4, in5, in6, in7, in8, in9, in10, in11, in12, in13, in14, in15, out1, out2, out3, out4, out5);
  input [11:0] in1, in2, in7;
  input in3, in4, in5, in6, in8, in9, in10, in11, in12, in13, in14, in15;
  output out1, out2, out3, out4, out5;
  wire [11:0] in1, in2, in7;
  wire in3, in4, in5, in6, in8, in9, in10, in11, in12, in13, in14, in15;
  wire out1, out2, out3, out4, out5;
  wire lt_42_22_n_0, lt_42_22_n_1, lt_42_22_n_2, lt_42_22_n_3, lt_42_22_n_4, lt_42_22_n_5, lt_42_22_n_6, lt_42_22_n_7;
  wire lt_42_22_n_8, lt_42_22_n_9, lt_42_22_n_10, lt_42_22_n_11, lt_42_22_n_12, lt_42_22_n_13, lt_42_22_n_14, lt_42_22_n_15;
  wire lt_42_22_n_16, lt_42_22_n_17, lt_42_22_n_18, lt_42_22_n_19, lt_42_22_n_20, lt_42_22_n_21, lt_42_22_n_22, lt_42_22_n_23;
  wire lt_42_22_n_24, lt_42_22_n_25, lt_42_22_n_26, lt_42_22_n_27, lt_42_22_n_28, lt_42_22_n_29, lt_42_22_n_30, lt_42_22_n_31;
  wire lt_42_22_n_32, lt_42_22_n_33, lt_42_22_n_34, lt_42_22_n_35, lt_42_22_n_36, lt_42_22_n_37, lt_42_22_n_38, lt_42_22_n_39;
  wire lt_42_22_n_40, lt_42_22_n_41, lt_42_22_n_42, lt_42_22_n_43, lt_42_22_n_44, lt_42_22_n_45, lt_42_22_n_46, lt_42_22_n_47;
  wire lt_42_22_n_48, lt_42_22_n_49, lt_42_22_n_50, lt_42_22_n_51, lt_42_22_n_52, lt_42_22_n_53, lt_42_22_n_54, lt_42_22_n_55;
  wire lt_42_22_n_56, lt_42_22_n_57, lt_42_22_n_58, lt_42_22_n_59, lt_42_22_n_60, lt_42_22_n_61, lt_42_22_n_62, lt_42_22_n_63;
  wire lt_42_22_n_64, lt_42_22_n_65, lt_42_22_n_66, lt_42_22_n_67, lt_42_22_n_68, lt_42_22_n_69, lt_42_22_n_70, lt_42_22_n_71;
  wire lt_42_22_n_72, lt_42_22_n_73, lt_43_22_n_0, lt_43_22_n_1, lt_43_22_n_2, lt_43_22_n_3, lt_43_22_n_4, lt_43_22_n_5;
  wire lt_43_22_n_6, lt_43_22_n_7, lt_43_22_n_8, lt_43_22_n_9, lt_43_22_n_10, lt_43_22_n_11, lt_43_22_n_12, lt_43_22_n_13;
  wire lt_43_22_n_14, lt_43_22_n_15, lt_43_22_n_16, lt_43_22_n_17, lt_43_22_n_18, lt_43_22_n_19, lt_43_22_n_20, lt_43_22_n_21;
  wire lt_43_22_n_22, lt_43_22_n_23, lt_43_22_n_24, lt_43_22_n_25, lt_43_22_n_26, lt_43_22_n_27, lt_43_22_n_28, lt_43_22_n_29;
  wire lt_43_22_n_30, lt_43_22_n_31, lt_43_22_n_32, lt_43_22_n_33, lt_43_22_n_34, lt_43_22_n_35, lt_43_22_n_36, lt_43_22_n_37;
  wire lt_43_22_n_38, lt_43_22_n_39, lt_43_22_n_40, lt_43_22_n_41, lt_43_22_n_42, lt_43_22_n_43, lt_43_22_n_44, lt_43_22_n_45;
  wire lt_43_22_n_46, lt_43_22_n_47, lt_43_22_n_48, lt_43_22_n_49, lt_43_22_n_50, lt_43_22_n_51, lt_43_22_n_52, lt_43_22_n_53;
  wire lt_43_22_n_54, lt_43_22_n_55, lt_43_22_n_56, lt_43_22_n_57, lt_43_22_n_58, lt_43_22_n_59, lt_43_22_n_60, lt_43_22_n_61;
  wire lt_43_22_n_62, lt_43_22_n_63, lt_43_22_n_64, lt_43_22_n_65, lt_43_22_n_66, lt_43_22_n_67, lt_43_22_n_68, lt_43_22_n_69;
  wire lt_43_22_n_70, lt_43_22_n_71, lt_43_22_n_72, lt_43_22_n_73, lt_44_22_n_0, lt_44_22_n_1, lt_44_22_n_2, lt_44_22_n_3;
  wire lt_44_22_n_4, lt_44_22_n_5, lt_44_22_n_6, lt_44_22_n_7, lt_44_22_n_8, lt_44_22_n_9, lt_44_22_n_10, lt_44_22_n_11;
  wire lt_44_22_n_12, lt_44_22_n_13, lt_44_22_n_14, lt_44_22_n_15, lt_44_22_n_16, lt_44_22_n_17, lt_44_22_n_18, lt_44_22_n_19;
  wire lt_44_22_n_20, lt_44_22_n_21, lt_44_22_n_22, lt_44_22_n_23, lt_44_22_n_24, lt_44_22_n_25, lt_44_22_n_26, lt_44_22_n_27;
  wire lt_44_22_n_28, lt_44_22_n_29, lt_44_22_n_30, lt_44_22_n_31, lt_44_22_n_32, lt_44_22_n_33, lt_44_22_n_34, lt_44_22_n_35;
  wire lt_44_22_n_36, lt_44_22_n_37, lt_44_22_n_38, lt_44_22_n_39, lt_44_22_n_40, lt_44_22_n_41, lt_44_22_n_42, lt_44_22_n_43;
  wire lt_44_22_n_44, lt_44_22_n_45, lt_44_22_n_46, lt_44_22_n_47, lt_44_22_n_48, lt_44_22_n_49, lt_44_22_n_50, lt_44_22_n_51;
  wire lt_44_22_n_52, lt_44_22_n_53, lt_44_22_n_54, lt_44_22_n_55, lt_44_22_n_56, lt_44_22_n_57, lt_44_22_n_58, lt_44_22_n_59;
  wire lt_44_22_n_60, lt_44_22_n_61, lt_44_22_n_62, lt_44_22_n_63, lt_44_22_n_64, lt_44_22_n_65, lt_44_22_n_66, lt_44_22_n_67;
  wire lt_44_22_n_68, lt_44_22_n_69, lt_44_22_n_70, lt_44_22_n_71, lt_44_22_n_72, lt_44_22_n_73, n_0, n_1;
  wire n_2, n_3, n_4, n_5, n_6, n_7, n_8, n_9;
  wire n_10, n_11, n_12, n_13, n_14, n_15, n_16, n_17;
  wire n_18, n_19, n_20, n_21, n_22, n_23, n_24, n_25;
  wire n_26, n_27, n_28, n_29, n_30, n_31, n_32, n_33;
  wire n_34, n_35, n_36, n_37, n_38, n_39, n_40, n_41;
  wire n_42, n_43, n_44, n_45, n_46, n_47, n_48, n_49;
  wire n_50, n_51, n_52, n_53, n_54, n_55, n_56, n_57;
  wire n_58, n_59, n_60, n_61, n_62, n_63, n_64, n_65;
  wire n_66, n_67, n_68, n_69, n_70, n_71, n_72, n_73;
  wire n_74, n_75, n_76, n_77, n_78, n_79, n_80, n_81;
  wire n_82, n_83, n_84, n_85, n_86, n_87, n_88, n_89;
  wire n_90, n_91, n_92, n_93, n_94, n_95, n_96, n_97;
  wire n_98, n_99, n_100, n_101, n_102, n_103, n_104, n_105;
  wire n_106, n_107, n_108, n_109, n_110, n_111, n_112, n_113;
  wire n_114, n_115, n_116, n_117, n_118, n_119, n_120, n_121;
  wire n_122, n_123, n_124, n_125, n_126, n_127, n_128, n_129;
  wire n_130, n_131, n_132, n_133, n_134, n_135, n_136, n_137;
  wire n_138, n_139, n_140, n_141, n_142, n_143, n_144, n_145;
  wire n_146, n_147, n_148, n_149, n_150, n_151, n_152, n_153;
  wire n_154, n_155, n_156, n_157, n_158, n_159, n_160, n_161;
  wire n_162, n_163, n_164, n_165, n_166, n_167, n_168, n_169;
  wire n_170, n_171, n_172, n_173, n_174, n_175, n_176, n_177;
  wire n_178, n_179, n_180, n_181, n_182, n_183, n_184, n_185;
  wire n_186, n_187, n_188, n_189, n_190, n_191, n_192, n_193;
  wire n_194, n_195, n_196, n_197, n_198, n_199, n_200, n_201;
  wire n_202, n_203, n_204, n_205, n_206, n_207, n_208, n_209;
  wire n_210, n_211, n_212, n_213, n_214, n_215, n_216, n_217;
  wire n_218, n_219, n_220, n_221, n_222, n_223, n_224, n_225;
  wire n_226, n_227, n_228, n_229, n_230, n_231, n_232, n_233;
  wire n_234, n_235, n_236, n_237, n_238, n_239, n_240, n_241;
  wire n_242, n_243, n_244, n_245, n_246, n_247, n_248, n_249;
  wire n_250, n_251, n_252, n_253, n_254, n_255, n_256, n_257;
  wire n_258, n_259, n_260, n_261, n_262, n_263, n_264, n_265;
  wire n_266, n_267, n_268, n_269, n_270, n_271, n_272, n_273;
  wire n_274, n_275, n_276, n_277, n_278, n_279, n_280, n_281;
  wire n_282, n_283, n_284, n_285, n_286, n_287, n_288, n_289;
  wire n_290, n_291, n_292, n_293, n_294, n_295, n_296, n_297;
  wire n_298, n_299, n_300, n_301, n_302, n_303, n_304, n_305;
  wire n_306, n_307, n_308, n_309, n_310, n_311, n_312, n_313;
  wire n_314, n_315, n_316, n_317, n_318, n_319, n_320, n_321;
  wire n_322, n_323, n_324, n_325, n_326, n_327, n_328, n_329;
  wire n_330, n_331, n_332, n_333, n_334, n_335, n_336, n_337;
  wire n_338, n_339, n_340, n_341, n_343, n_344, n_345, n_346;
  wire n_347, n_348, n_349, n_350, n_351, n_352, n_353, n_354;
  wire n_355, n_356, n_357, n_358, n_359, n_360, n_361, n_362;
  wire n_363, n_364, n_365, n_366, n_367, n_368, n_369, n_370;
  wire n_371, n_372, n_373, n_374, n_375, n_376, n_377, n_378;
  wire n_379, n_380, n_381, n_382, n_383, n_384, n_385, n_386;
  wire n_387, n_388, n_389, n_390, n_391, n_392, n_393, n_394;
  wire n_395, n_396, n_397, n_398, n_399, n_400, n_401, n_402;
  wire n_403, n_404, n_405, n_406, n_407, n_408, n_409, n_410;
  wire n_411, n_412, n_413, n_414, n_415, n_416, n_417, n_418;
  wire n_419, n_420, n_421, n_422, n_423, n_424, n_425, n_426;
  wire n_427, n_428, n_429, n_430, n_431, n_432, n_434, n_435;
  wire n_436, n_437, n_438, n_439, n_440, n_441, n_442, n_443;
  wire n_444, n_445, n_446, n_447, n_448, n_449, n_450, n_451;
  wire n_452, n_453, n_454, n_455, n_456, n_457, n_458, n_459;
  wire n_460, n_461, n_462, n_463, n_464, n_465, n_466, n_467;
  wire n_468, n_469, n_470, n_471, sub_32_21_n_2, sub_32_21_n_3, sub_32_21_n_4, sub_32_21_n_5;
  wire sub_32_21_n_6, sub_32_21_n_7, sub_32_21_n_8, sub_32_21_n_9, sub_32_21_n_10, sub_32_21_n_11, sub_32_21_n_12, sub_32_21_n_13;
  wire sub_32_21_n_14, sub_32_21_n_15, sub_32_21_n_16, sub_32_21_n_17, sub_32_21_n_18, sub_32_21_n_19, sub_32_21_n_20, sub_32_21_n_21;
  wire sub_32_21_n_22, sub_32_21_n_23, sub_32_21_n_24, sub_32_21_n_25, sub_32_21_n_26, sub_32_21_n_27, sub_32_21_n_28, sub_32_21_n_29;
  wire sub_32_21_n_30, sub_32_21_n_31, sub_32_21_n_32, sub_32_21_n_33, sub_32_21_n_34, sub_32_21_n_35, sub_32_21_n_36, sub_32_21_n_37;
  wire sub_32_21_n_38, sub_32_21_n_39, sub_32_21_n_40, sub_32_21_n_41, sub_32_21_n_42, sub_32_21_n_43, sub_32_21_n_44, sub_32_21_n_45;
  wire sub_32_21_n_46, sub_32_21_n_47, sub_32_21_n_48, sub_32_21_n_49, sub_32_21_n_50, sub_32_21_n_51, sub_32_21_n_52, sub_32_21_n_53;
  wire sub_32_21_n_54, sub_32_21_n_55, sub_32_21_n_56, sub_32_21_n_57, sub_32_21_n_58, sub_32_21_n_59, sub_32_21_n_61, sub_32_21_n_63;
  wire sub_32_21_n_64, sub_32_21_n_66, sub_32_21_n_67, sub_32_21_n_69, sub_32_21_n_70, sub_32_21_n_72, sub_32_21_n_73, sub_32_21_n_75;
  wire sub_32_21_n_76, sub_32_21_n_78, sub_32_21_n_79, sub_32_21_n_81, sub_32_21_n_82, sub_32_21_n_84, sub_32_21_n_85, sub_32_21_n_87;
  wire sub_32_21_n_88, sub_32_21_n_90, sub_33_31_n_0, sub_33_31_n_1, sub_33_31_n_2, sub_33_31_n_3, sub_33_31_n_4, sub_33_31_n_5;
  wire sub_33_31_n_6, sub_33_31_n_7, sub_33_31_n_8, sub_33_31_n_9, sub_33_31_n_10, sub_33_31_n_24, sub_33_31_n_25, sub_33_31_n_26;
  wire sub_33_31_n_27, sub_33_31_n_28, sub_33_31_n_29, sub_33_31_n_30, sub_33_31_n_31, sub_33_31_n_32, sub_33_31_n_33, sub_33_31_n_34;
  wire sub_33_31_n_35, sub_33_31_n_36, sub_33_31_n_37, sub_33_31_n_38, sub_33_31_n_39, sub_33_31_n_40, sub_33_31_n_41, sub_33_31_n_42;
  wire sub_33_31_n_43, sub_33_31_n_44, sub_33_31_n_45, sub_33_31_n_46, sub_33_31_n_47, sub_33_31_n_48, sub_33_31_n_49, sub_33_31_n_50;
  wire sub_33_31_n_51, sub_35_21_n_2, sub_35_21_n_3, sub_35_21_n_4, sub_35_21_n_5, sub_35_21_n_6, sub_35_21_n_7, sub_35_21_n_8;
  wire sub_35_21_n_9, sub_35_21_n_10, sub_35_21_n_11, sub_35_21_n_12, sub_35_21_n_13, sub_35_21_n_14, sub_35_21_n_15, sub_35_21_n_16;
  wire sub_35_21_n_17, sub_35_21_n_18, sub_35_21_n_19, sub_35_21_n_20, sub_35_21_n_21, sub_35_21_n_22, sub_35_21_n_23, sub_35_21_n_24;
  wire sub_35_21_n_25, sub_35_21_n_26, sub_35_21_n_27, sub_35_21_n_28, sub_35_21_n_29, sub_35_21_n_30, sub_35_21_n_31, sub_35_21_n_32;
  wire sub_35_21_n_33, sub_35_21_n_34, sub_35_21_n_35, sub_35_21_n_36, sub_35_21_n_37, sub_35_21_n_38, sub_35_21_n_39, sub_35_21_n_40;
  wire sub_35_21_n_41, sub_35_21_n_42, sub_35_21_n_43, sub_35_21_n_44, sub_35_21_n_45, sub_35_21_n_46, sub_35_21_n_47, sub_35_21_n_48;
  wire sub_35_21_n_49, sub_35_21_n_50, sub_35_21_n_51, sub_35_21_n_52, sub_35_21_n_53, sub_35_21_n_54, sub_35_21_n_55, sub_35_21_n_56;
  wire sub_35_21_n_57, sub_35_21_n_58, sub_35_21_n_59, sub_35_21_n_61, sub_35_21_n_63, sub_35_21_n_64, sub_35_21_n_66, sub_35_21_n_67;
  wire sub_35_21_n_69, sub_35_21_n_70, sub_35_21_n_72, sub_35_21_n_73, sub_35_21_n_75, sub_35_21_n_76, sub_35_21_n_78, sub_35_21_n_79;
  wire sub_35_21_n_81, sub_35_21_n_82, sub_35_21_n_84, sub_35_21_n_85, sub_35_21_n_87, sub_35_21_n_88, sub_35_21_n_90, sub_36_31_n_0;
  wire sub_36_31_n_1, sub_36_31_n_2, sub_36_31_n_3, sub_36_31_n_4, sub_36_31_n_5, sub_36_31_n_6, sub_36_31_n_7, sub_36_31_n_8;
  wire sub_36_31_n_9, sub_36_31_n_10, sub_36_31_n_24, sub_36_31_n_25, sub_36_31_n_26, sub_36_31_n_27, sub_36_31_n_28, sub_36_31_n_29;
  wire sub_36_31_n_30, sub_36_31_n_31, sub_36_31_n_32, sub_36_31_n_33, sub_36_31_n_34, sub_36_31_n_35, sub_36_31_n_36, sub_36_31_n_37;
  wire sub_36_31_n_38, sub_36_31_n_39, sub_36_31_n_40, sub_36_31_n_41, sub_36_31_n_42, sub_36_31_n_43, sub_36_31_n_44, sub_36_31_n_45;
  wire sub_36_31_n_46, sub_36_31_n_47, sub_36_31_n_48, sub_36_31_n_49, sub_36_31_n_50, sub_36_31_n_51;
  or g777__2398(n_392 ,n_294 ,n_329);
  or g778__5107(n_366 ,n_278 ,n_315);
  or g779__6260(n_361 ,n_295 ,n_330);
  or g780__4319(n_394 ,n_298 ,n_339);
  or g781__8428(n_438 ,n_301 ,n_337);
  or g782__5526(n_437 ,n_299 ,n_336);
  or g783__6783(n_436 ,n_290 ,n_334);
  or g784__3680(n_393 ,n_303 ,n_339);
  or g785__1617(n_435 ,n_277 ,n_332);
  or g786__2802(n_368 ,n_287 ,n_340);
  or g787__1705(n_434 ,n_300 ,n_331);
  or g788__5122(n_391 ,n_293 ,n_328);
  or g789__8246(n_390 ,n_289 ,n_327);
  or g790__7098(n_364 ,n_281 ,n_321);
  or g791__6131(n_360 ,n_285 ,n_323);
  or g792__1881(n_389 ,n_286 ,n_325);
  or g793__5115(n_388 ,n_282 ,n_324);
  or g794__7482(n_387 ,n_280 ,n_320);
  or g795__4733(n_359 ,n_288 ,n_316);
  or g796__6161(n_386 ,n_279 ,n_319);
  or g797__9315(n_385 ,n_284 ,n_318);
  or g798__9945(n_384 ,n_292 ,n_317);
  or g799__2883(n_367 ,n_269 ,n_340);
  or g800__2346(n_363 ,n_272 ,n_309);
  or g801__1666(n_358 ,n_270 ,n_310);
  or g802__7410(n_383 ,n_274 ,n_314);
  or g803__6417(n_382 ,n_296 ,n_313);
  or g804__5477(n_357 ,n_268 ,n_306);
  or g805__2398(n_446 ,n_297 ,n_341);
  or g806__5107(n_445 ,n_267 ,n_341);
  or g807__6260(n_444 ,n_291 ,n_308);
  or g808__4319(n_365 ,n_302 ,n_333);
  or g809__8428(n_443 ,n_276 ,n_307);
  or g810__5526(n_442 ,n_271 ,n_312);
  or g811__6783(n_441 ,n_273 ,n_305);
  or g812__3680(n_362 ,n_338 ,n_335);
  or g813__1617(n_356 ,n_275 ,n_311);
  or g814__2802(n_440 ,n_304 ,n_322);
  or g815__1705(n_439 ,n_283 ,n_326);
  and g816__5122(n_338 ,n_210 ,n_453);
  and g817__8246(n_337 ,n_239 ,n_181);
  and g818__7098(n_336 ,n_236 ,n_182);
  and g819__6131(n_335 ,n_221 ,n_175);
  and g820__1881(n_334 ,n_233 ,n_200);
  and g821__5115(n_333 ,n_227 ,n_176);
  and g822__7482(n_332 ,n_242 ,n_182);
  and g823__4733(n_331 ,n_224 ,n_181);
  and g824__6161(n_330 ,n_218 ,n_198);
  and g825__9315(n_329 ,n_203 ,n_187);
  and g826__9945(n_328 ,n_226 ,n_188);
  and g827__2883(n_327 ,n_245 ,n_196);
  and g828__2346(n_326 ,n_217 ,n_184);
  and g829__1666(n_325 ,n_230 ,n_188);
  and g830__7410(n_324 ,n_220 ,n_187);
  and g831__6417(n_323 ,n_238 ,n_176);
  and g832__5477(n_322 ,n_221 ,n_184);
  and g833__2398(n_321 ,n_244 ,n_175);
  and g834__5107(n_320 ,n_218 ,n_172);
  and g835__6260(n_319 ,n_239 ,n_172);
  and g836__4319(n_318 ,n_235 ,n_263);
  and g837__8428(n_317 ,n_232 ,n_263);
  and g838__5526(n_316 ,n_236 ,n_178);
  and g839__6783(n_315 ,n_202 ,n_178);
  and g840__3680(n_314 ,n_241 ,n_196);
  and g841__1617(n_313 ,n_223 ,n_173);
  and g842__2802(n_312 ,n_245 ,n_251);
  and g843__1705(n_311 ,n_224 ,n_257);
  and g844__5122(n_310 ,n_233 ,n_257);
  and g845__8246(n_309 ,n_229 ,n_198);
  and g846__7098(n_308 ,n_203 ,n_251);
  and g847__6131(n_307 ,n_227 ,n_200);
  and g848__1881(n_306 ,n_242 ,n_179);
  and g849__5115(n_305 ,n_230 ,n_185);
  and g850__7482(n_341 ,n_248 ,n_185);
  and g851__4733(n_340 ,n_247 ,n_179);
  and g852__6161(n_339 ,n_248 ,n_173);
  and g853__9315(n_304 ,n_206 ,n_453);
  and g854__9945(n_303 ,n_204 ,n_458);
  and g855__2883(n_302 ,n_211 ,n_456);
  and g856__2346(n_301 ,n_207 ,n_451);
  and g857__1666(n_300 ,n_253 ,n_447);
  and g858__7410(n_299 ,n_192 ,n_450);
  and g859__6417(n_298 ,n_205 ,n_459);
  and g860__5477(n_297 ,n_207 ,n_459);
  and g861__2398(n_296 ,n_265 ,n_447);
  and g862__5107(n_295 ,n_259 ,n_452);
  and g863__6260(n_294 ,n_194 ,n_457);
  and g864__4319(n_293 ,n_205 ,n_456);
  and g865__8428(n_292 ,n_262 ,n_449);
  and g866__5526(n_291 ,n_250 ,n_457);
  and g867__6783(n_290 ,n_192 ,n_449);
  and g868__3680(n_289 ,n_194 ,n_455);
  and g869__1617(n_288 ,n_190 ,n_450);
  and g870__2802(n_287 ,n_211 ,n_459);
  and g871__1705(n_286 ,n_212 ,n_454);
  and g872__5122(n_285 ,n_256 ,n_451);
  and g873__8246(n_284 ,n_204 ,n_450);
  and g874__7098(n_283 ,n_208 ,n_452);
  and g875__6131(n_282 ,n_262 ,n_453);
  and g876__1881(n_281 ,n_190 ,n_455);
  and g877__5115(n_280 ,n_213 ,n_452);
  and g878__7482(n_279 ,n_213 ,n_451);
  and g879__4733(n_278 ,n_214 ,n_457);
  and g880__6161(n_277 ,n_206 ,n_448);
  and g881__9315(n_276 ,n_250 ,n_456);
  and g882__9945(n_275 ,n_210 ,n_447);
  and g883__2883(n_274 ,n_212 ,n_448);
  and g884__2346(n_273 ,n_209 ,n_454);
  and g885__1666(n_272 ,n_256 ,n_454);
  and g886__7410(n_271 ,n_209 ,n_455);
  and g887__6417(n_270 ,n_215 ,n_449);
  and g888__5477(n_269 ,n_215 ,n_458);
  and g889__2398(n_268 ,n_214 ,n_448);
  and g890__5107(n_267 ,n_208 ,n_458);
  not g891(n_266 ,in10);
  not g892(n_265 ,n_264);
  not g894(n_264 ,in10);
  not g895(n_263 ,in10);
  not g896(n_262 ,n_261);
  not g898(n_261 ,in10);
  not g899(n_260 ,in14);
  not g900(n_259 ,n_258);
  not g902(n_258 ,in14);
  not g903(n_257 ,in14);
  not g904(n_256 ,n_255);
  not g906(n_255 ,in14);
  not g907(n_254 ,in3);
  not g908(n_253 ,n_252);
  not g910(n_252 ,in3);
  not g911(n_251 ,in3);
  not g912(n_250 ,n_249);
  not g914(n_249 ,in3);
  not drc_bufs929(n_248 ,n_246);
  not drc_bufs930(n_247 ,n_246);
  not drc_bufs931(n_246 ,out5);
  not drc_bufs933(n_245 ,n_243);
  not drc_bufs934(n_244 ,n_243);
  not drc_bufs935(n_243 ,n_469);
  not drc_bufs937(n_242 ,n_240);
  not drc_bufs938(n_241 ,n_240);
  not drc_bufs939(n_240 ,n_462);
  not drc_bufs941(n_239 ,n_237);
  not drc_bufs942(n_238 ,n_237);
  not drc_bufs943(n_237 ,n_465);
  not drc_bufs945(n_236 ,n_234);
  not drc_bufs946(n_235 ,n_234);
  not drc_bufs947(n_234 ,n_464);
  not drc_bufs949(n_233 ,n_231);
  not drc_bufs950(n_232 ,n_231);
  not drc_bufs951(n_231 ,n_463);
  not drc_bufs953(n_230 ,n_228);
  not drc_bufs954(n_229 ,n_228);
  not drc_bufs955(n_228 ,n_468);
  not drc_bufs957(n_227 ,n_225);
  not drc_bufs958(n_226 ,n_225);
  not drc_bufs959(n_225 ,n_470);
  not drc_bufs961(n_224 ,n_222);
  not drc_bufs962(n_223 ,n_222);
  not drc_bufs963(n_222 ,n_461);
  not drc_bufs965(n_221 ,n_219);
  not drc_bufs966(n_220 ,n_219);
  not drc_bufs967(n_219 ,n_467);
  not drc_bufs969(n_218 ,n_216);
  not drc_bufs970(n_217 ,n_216);
  not drc_bufs971(n_216 ,n_466);
  not drc_bufs973(n_215 ,n_255);
  not drc_bufs974(n_214 ,n_255);
  not drc_bufs977(n_213 ,n_261);
  not drc_bufs978(n_212 ,n_261);
  not drc_bufs981(n_211 ,n_258);
  not drc_bufs982(n_210 ,n_258);
  not drc_bufs985(n_209 ,n_249);
  not drc_bufs986(n_208 ,n_249);
  not drc_bufs989(n_207 ,n_252);
  not drc_bufs990(n_206 ,n_252);
  not drc_bufs993(n_205 ,n_264);
  not drc_bufs994(n_204 ,n_264);
  not drc_bufs997(n_203 ,n_201);
  not drc_bufs998(n_202 ,n_201);
  not drc_bufs999(n_201 ,n_471);
  not drc_bufs1002(n_200 ,n_199);
  not drc_bufs1003(n_199 ,n_251);
  not drc_bufs1006(n_198 ,n_197);
  not drc_bufs1007(n_197 ,n_257);
  not drc_bufs1010(n_196 ,n_195);
  not drc_bufs1011(n_195 ,n_263);
  not drc_bufs1013(n_194 ,n_193);
  not drc_bufs1015(n_193 ,n_265);
  not drc_bufs1017(n_192 ,n_191);
  not drc_bufs1019(n_191 ,n_253);
  not drc_bufs1021(n_190 ,n_189);
  not drc_bufs1023(n_189 ,n_259);
  not drc_bufs1025(n_188 ,n_186);
  not drc_bufs1026(n_187 ,n_186);
  not drc_bufs1027(n_186 ,n_266);
  not drc_bufs1029(n_185 ,n_183);
  not drc_bufs1030(n_184 ,n_183);
  not drc_bufs1031(n_183 ,n_254);
  not drc_bufs1033(n_182 ,n_180);
  not drc_bufs1034(n_181 ,n_180);
  not drc_bufs1035(n_180 ,n_254);
  not drc_bufs1037(n_179 ,n_177);
  not drc_bufs1038(n_178 ,n_177);
  not drc_bufs1039(n_177 ,n_260);
  not drc_bufs1041(n_176 ,n_174);
  not drc_bufs1042(n_175 ,n_174);
  not drc_bufs1043(n_174 ,n_260);
  not drc_bufs1045(n_173 ,n_171);
  not drc_bufs1046(n_172 ,n_171);
  not drc_bufs1047(n_171 ,n_266);
  or g1050__6260(n_379 ,n_123 ,n_158);
  or g1051__4319(n_353 ,n_107 ,n_144);
  or g1052__8428(n_348 ,n_124 ,n_159);
  or g1053__5526(n_381 ,n_127 ,n_168);
  or g1054__6783(n_399 ,n_130 ,n_166);
  or g1055__3680(n_398 ,n_128 ,n_165);
  or g1056__1617(n_397 ,n_119 ,n_163);
  or g1057__2802(n_380 ,n_132 ,n_168);
  or g1058__1705(n_396 ,n_106 ,n_161);
  or g1059__5122(n_355 ,n_116 ,n_169);
  or g1060__8246(n_395 ,n_129 ,n_160);
  or g1061__7098(n_378 ,n_122 ,n_157);
  or g1062__6131(n_377 ,n_118 ,n_156);
  or g1063__1881(n_351 ,n_110 ,n_150);
  or g1064__5115(n_347 ,n_114 ,n_152);
  or g1065__7482(n_376 ,n_115 ,n_154);
  or g1066__4733(n_375 ,n_111 ,n_153);
  or g1067__6161(n_374 ,n_109 ,n_149);
  or g1068__9315(n_346 ,n_117 ,n_145);
  or g1069__9945(n_373 ,n_108 ,n_148);
  or g1070__2883(n_372 ,n_113 ,n_147);
  or g1071__2346(n_371 ,n_121 ,n_146);
  or g1072__1666(n_354 ,n_98 ,n_169);
  or g1073__7410(n_350 ,n_101 ,n_138);
  or g1074__6417(n_345 ,n_99 ,n_139);
  or g1075__5477(n_370 ,n_103 ,n_143);
  or g1076__2398(n_369 ,n_125 ,n_142);
  or g1077__5107(n_344 ,n_97 ,n_135);
  or g1078__6260(n_407 ,n_126 ,n_170);
  or g1079__4319(n_406 ,n_96 ,n_170);
  or g1080__8428(n_405 ,n_120 ,n_137);
  or g1081__5526(n_352 ,n_131 ,n_162);
  or g1082__6783(n_404 ,n_105 ,n_136);
  or g1083__3680(n_403 ,n_100 ,n_141);
  or g1084__1617(n_402 ,n_102 ,n_134);
  or g1085__2802(n_349 ,n_167 ,n_164);
  or g1086__1705(n_343 ,n_104 ,n_140);
  or g1087__5122(n_401 ,n_133 ,n_151);
  or g1088__8246(n_400 ,n_112 ,n_155);
  and g1089__7098(n_167 ,n_39 ,n_414);
  and g1090__6131(n_166 ,n_68 ,n_10);
  and g1091__1881(n_165 ,n_65 ,n_11);
  and g1092__5115(n_164 ,n_50 ,n_4);
  and g1093__7482(n_163 ,n_62 ,n_29);
  and g1094__4733(n_162 ,n_56 ,n_5);
  and g1095__6161(n_161 ,n_71 ,n_11);
  and g1096__9315(n_160 ,n_53 ,n_10);
  and g1097__9945(n_159 ,n_47 ,n_27);
  and g1098__2883(n_158 ,n_32 ,n_16);
  and g1099__2346(n_157 ,n_55 ,n_17);
  and g1100__1666(n_156 ,n_74 ,n_25);
  and g1101__7410(n_155 ,n_46 ,n_13);
  and g1102__6417(n_154 ,n_59 ,n_17);
  and g1103__5477(n_153 ,n_49 ,n_16);
  and g1104__2398(n_152 ,n_67 ,n_5);
  and g1105__5107(n_151 ,n_50 ,n_13);
  and g1106__6260(n_150 ,n_73 ,n_4);
  and g1107__4319(n_149 ,n_47 ,n_1);
  and g1108__8428(n_148 ,n_68 ,n_1);
  and g1109__5526(n_147 ,n_64 ,n_92);
  and g1110__6783(n_146 ,n_61 ,n_92);
  and g1111__3680(n_145 ,n_65 ,n_7);
  and g1112__1617(n_144 ,n_31 ,n_7);
  and g1113__2802(n_143 ,n_70 ,n_25);
  and g1114__1705(n_142 ,n_52 ,n_2);
  and g1115__5122(n_141 ,n_74 ,n_80);
  and g1116__8246(n_140 ,n_53 ,n_86);
  and g1117__7098(n_139 ,n_62 ,n_86);
  and g1118__6131(n_138 ,n_58 ,n_27);
  and g1119__1881(n_137 ,n_32 ,n_80);
  and g1120__5115(n_136 ,n_56 ,n_29);
  and g1121__7482(n_135 ,n_71 ,n_8);
  and g1122__4733(n_134 ,n_59 ,n_14);
  and g1123__6161(n_170 ,n_77 ,n_14);
  and g1124__9315(n_169 ,n_76 ,n_8);
  and g1125__9945(n_168 ,n_77 ,n_2);
  and g1126__2883(n_133 ,n_35 ,n_414);
  and g1127__2346(n_132 ,n_33 ,n_419);
  and g1128__1666(n_131 ,n_40 ,n_417);
  and g1129__7410(n_130 ,n_36 ,n_412);
  and g1130__6417(n_129 ,n_82 ,n_408);
  and g1131__5477(n_128 ,n_21 ,n_411);
  and g1132__2398(n_127 ,n_34 ,n_420);
  and g1133__5107(n_126 ,n_36 ,n_420);
  and g1134__6260(n_125 ,n_94 ,n_408);
  and g1135__4319(n_124 ,n_88 ,n_413);
  and g1136__8428(n_123 ,n_23 ,n_418);
  and g1137__5526(n_122 ,n_34 ,n_417);
  and g1138__6783(n_121 ,n_91 ,n_410);
  and g1139__3680(n_120 ,n_79 ,n_418);
  and g1140__1617(n_119 ,n_21 ,n_410);
  and g1141__2802(n_118 ,n_23 ,n_416);
  and g1142__1705(n_117 ,n_19 ,n_411);
  and g1143__5122(n_116 ,n_40 ,n_420);
  and g1144__8246(n_115 ,n_41 ,n_415);
  and g1145__7098(n_114 ,n_85 ,n_412);
  and g1146__6131(n_113 ,n_33 ,n_411);
  and g1147__1881(n_112 ,n_37 ,n_413);
  and g1148__5115(n_111 ,n_91 ,n_414);
  and g1149__7482(n_110 ,n_19 ,n_416);
  and g1150__4733(n_109 ,n_42 ,n_413);
  and g1151__6161(n_108 ,n_42 ,n_412);
  and g1152__9315(n_107 ,n_43 ,n_418);
  and g1153__9945(n_106 ,n_35 ,n_409);
  and g1154__2883(n_105 ,n_79 ,n_417);
  and g1155__2346(n_104 ,n_39 ,n_408);
  and g1156__1666(n_103 ,n_41 ,n_409);
  and g1157__7410(n_102 ,n_38 ,n_415);
  and g1158__6417(n_101 ,n_85 ,n_415);
  and g1159__5477(n_100 ,n_38 ,n_416);
  and g1160__2398(n_99 ,n_44 ,n_410);
  and g1161__5107(n_98 ,n_44 ,n_419);
  and g1162__6260(n_97 ,n_43 ,n_409);
  and g1163__4319(n_96 ,n_37 ,n_419);
  not g1164(n_95 ,in8);
  not g1165(n_94 ,n_93);
  not g1166(n_93 ,in8);
  not g1167(n_92 ,in8);
  not g1168(n_91 ,n_90);
  not g1169(n_90 ,in8);
  not g1170(n_89 ,in12);
  not g1171(n_88 ,n_87);
  not g1172(n_87 ,in12);
  not g1173(n_86 ,in12);
  not g1174(n_85 ,n_84);
  not g1175(n_84 ,in12);
  not g1176(n_83 ,in5);
  not g1177(n_82 ,n_81);
  not g1178(n_81 ,in5);
  not g1179(n_80 ,in5);
  not g1180(n_79 ,n_78);
  not g1181(n_78 ,in5);
  not drc_bufs1182(n_77 ,n_75);
  not drc_bufs1183(n_76 ,n_75);
  not drc_bufs1184(n_75 ,out4);
  not drc_bufs1185(n_74 ,n_72);
  not drc_bufs1186(n_73 ,n_72);
  not drc_bufs1187(n_72 ,n_430);
  not drc_bufs1188(n_71 ,n_69);
  not drc_bufs1189(n_70 ,n_69);
  not drc_bufs1190(n_69 ,n_423);
  not drc_bufs1191(n_68 ,n_66);
  not drc_bufs1192(n_67 ,n_66);
  not drc_bufs1193(n_66 ,n_426);
  not drc_bufs1194(n_65 ,n_63);
  not drc_bufs1195(n_64 ,n_63);
  not drc_bufs1196(n_63 ,n_425);
  not drc_bufs1197(n_62 ,n_60);
  not drc_bufs1198(n_61 ,n_60);
  not drc_bufs1199(n_60 ,n_424);
  not drc_bufs1200(n_59 ,n_57);
  not drc_bufs1201(n_58 ,n_57);
  not drc_bufs1202(n_57 ,n_429);
  not drc_bufs1203(n_56 ,n_54);
  not drc_bufs1204(n_55 ,n_54);
  not drc_bufs1205(n_54 ,n_431);
  not drc_bufs1206(n_53 ,n_51);
  not drc_bufs1207(n_52 ,n_51);
  not drc_bufs1208(n_51 ,n_422);
  not drc_bufs1209(n_50 ,n_48);
  not drc_bufs1210(n_49 ,n_48);
  not drc_bufs1211(n_48 ,n_428);
  not drc_bufs1212(n_47 ,n_45);
  not drc_bufs1213(n_46 ,n_45);
  not drc_bufs1214(n_45 ,n_427);
  not drc_bufs1215(n_44 ,n_84);
  not drc_bufs1216(n_43 ,n_84);
  not drc_bufs1217(n_42 ,n_90);
  not drc_bufs1218(n_41 ,n_90);
  not drc_bufs1219(n_40 ,n_87);
  not drc_bufs1220(n_39 ,n_87);
  not drc_bufs1221(n_38 ,n_78);
  not drc_bufs1222(n_37 ,n_78);
  not drc_bufs1223(n_36 ,n_81);
  not drc_bufs1224(n_35 ,n_81);
  not drc_bufs1225(n_34 ,n_93);
  not drc_bufs1226(n_33 ,n_93);
  not drc_bufs1227(n_32 ,n_30);
  not drc_bufs1228(n_31 ,n_30);
  not drc_bufs1229(n_30 ,n_432);
  not drc_bufs1230(n_29 ,n_28);
  not drc_bufs1231(n_28 ,n_80);
  not drc_bufs1232(n_27 ,n_26);
  not drc_bufs1233(n_26 ,n_86);
  not drc_bufs1234(n_25 ,n_24);
  not drc_bufs1235(n_24 ,n_92);
  not drc_bufs1236(n_23 ,n_22);
  not drc_bufs1237(n_22 ,n_94);
  not drc_bufs1238(n_21 ,n_20);
  not drc_bufs1239(n_20 ,n_82);
  not drc_bufs1240(n_19 ,n_18);
  not drc_bufs1241(n_18 ,n_88);
  not drc_bufs1242(n_17 ,n_15);
  not drc_bufs1243(n_16 ,n_15);
  not drc_bufs1244(n_15 ,n_95);
  not drc_bufs1245(n_14 ,n_12);
  not drc_bufs1246(n_13 ,n_12);
  not drc_bufs1247(n_12 ,n_83);
  not drc_bufs1248(n_11 ,n_9);
  not drc_bufs1249(n_10 ,n_9);
  not drc_bufs1250(n_9 ,n_83);
  not drc_bufs1251(n_8 ,n_6);
  not drc_bufs1252(n_7 ,n_6);
  not drc_bufs1253(n_6 ,n_89);
  not drc_bufs1254(n_5 ,n_3);
  not drc_bufs1255(n_4 ,n_3);
  not drc_bufs1256(n_3 ,n_89);
  not drc_bufs1257(n_2 ,n_0);
  not drc_bufs1258(n_1 ,n_0);
  not drc_bufs1259(n_0 ,n_95);
  or lt_42_22_g242__8428(out1 ,lt_42_22_n_33 ,lt_42_22_n_73);
  nor lt_42_22_g243__5526(lt_42_22_n_73 ,lt_42_22_n_24 ,lt_42_22_n_72);
  or lt_42_22_g244__6783(lt_42_22_n_72 ,lt_42_22_n_41 ,lt_42_22_n_71);
  nor lt_42_22_g245__3680(lt_42_22_n_71 ,lt_42_22_n_29 ,lt_42_22_n_70);
  nor lt_42_22_g246__1617(lt_42_22_n_70 ,lt_42_22_n_40 ,lt_42_22_n_69);
  nor lt_42_22_g247__2802(lt_42_22_n_69 ,lt_42_22_n_36 ,lt_42_22_n_68);
  nor lt_42_22_g248__1705(lt_42_22_n_68 ,lt_42_22_n_35 ,lt_42_22_n_67);
  nor lt_42_22_g249__5122(lt_42_22_n_67 ,lt_42_22_n_31 ,lt_42_22_n_66);
  nor lt_42_22_g250__8246(lt_42_22_n_66 ,lt_42_22_n_28 ,lt_42_22_n_65);
  nor lt_42_22_g251__7098(lt_42_22_n_65 ,lt_42_22_n_22 ,lt_42_22_n_64);
  nor lt_42_22_g252__6131(lt_42_22_n_64 ,lt_42_22_n_44 ,lt_42_22_n_63);
  nor lt_42_22_g253__1881(lt_42_22_n_63 ,lt_42_22_n_26 ,lt_42_22_n_62);
  nor lt_42_22_g254__5115(lt_42_22_n_62 ,lt_42_22_n_37 ,lt_42_22_n_61);
  nor lt_42_22_g255__7482(lt_42_22_n_61 ,lt_42_22_n_38 ,lt_42_22_n_60);
  nor lt_42_22_g256__4733(lt_42_22_n_60 ,lt_42_22_n_34 ,lt_42_22_n_59);
  nor lt_42_22_g257__6161(lt_42_22_n_59 ,lt_42_22_n_32 ,lt_42_22_n_58);
  nor lt_42_22_g258__9315(lt_42_22_n_58 ,lt_42_22_n_30 ,lt_42_22_n_57);
  nor lt_42_22_g259__9945(lt_42_22_n_57 ,lt_42_22_n_27 ,lt_42_22_n_56);
  nor lt_42_22_g260__2883(lt_42_22_n_56 ,lt_42_22_n_25 ,lt_42_22_n_55);
  nor lt_42_22_g261__2346(lt_42_22_n_55 ,lt_42_22_n_23 ,lt_42_22_n_54);
  nor lt_42_22_g262__1666(lt_42_22_n_54 ,lt_42_22_n_39 ,lt_42_22_n_53);
  nor lt_42_22_g263__7410(lt_42_22_n_53 ,lt_42_22_n_43 ,lt_42_22_n_52);
  nor lt_42_22_g264__6417(lt_42_22_n_52 ,lt_42_22_n_42 ,lt_42_22_n_51);
  nor lt_42_22_g265__5477(lt_42_22_n_51 ,lt_42_22_n_45 ,lt_42_22_n_50);
  nor lt_42_22_g266__2398(lt_42_22_n_50 ,lt_42_22_n_48 ,lt_42_22_n_49);
  nor lt_42_22_g267__5107(lt_42_22_n_49 ,n_395 ,lt_42_22_n_47);
  and lt_42_22_g268__6260(lt_42_22_n_48 ,n_434 ,lt_42_22_n_46);
  nor lt_42_22_g269__4319(lt_42_22_n_47 ,n_434 ,lt_42_22_n_46);
  nor lt_42_22_g270__8428(lt_42_22_n_45 ,lt_42_22_n_13 ,n_435);
  nor lt_42_22_g271__5526(lt_42_22_n_44 ,lt_42_22_n_18 ,n_402);
  nor lt_42_22_g272__6783(lt_42_22_n_43 ,lt_42_22_n_19 ,n_436);
  nor lt_42_22_g273__3680(lt_42_22_n_42 ,lt_42_22_n_11 ,n_396);
  nor lt_42_22_g274__1617(lt_42_22_n_41 ,lt_42_22_n_3 ,n_406);
  nor lt_42_22_g275__2802(lt_42_22_n_40 ,lt_42_22_n_20 ,n_405);
  nor lt_42_22_g276__1705(lt_42_22_n_39 ,lt_42_22_n_16 ,n_397);
  nor lt_42_22_g277__5122(lt_42_22_n_38 ,lt_42_22_n_10 ,n_440);
  nor lt_42_22_g278__8246(lt_42_22_n_37 ,lt_42_22_n_15 ,n_401);
  nor lt_42_22_g279__7098(lt_42_22_n_36 ,lt_42_22_n_8 ,n_444);
  nor lt_42_22_g280__6131(lt_42_22_n_35 ,lt_42_22_n_1 ,n_404);
  or lt_42_22_g281__1881(lt_42_22_n_46 ,lt_42_22_n_7 ,n_460);
  nor lt_42_22_g282__5115(lt_42_22_n_34 ,lt_42_22_n_14 ,n_400);
  nor lt_42_22_g283__7482(lt_42_22_n_33 ,lt_42_22_n_5 ,n_407);
  nor lt_42_22_g284__4733(lt_42_22_n_32 ,lt_42_22_n_6 ,n_439);
  and lt_42_22_g285__6161(lt_42_22_n_31 ,n_404 ,lt_42_22_n_1);
  nor lt_42_22_g286__9315(lt_42_22_n_30 ,lt_42_22_n_9 ,n_399);
  and lt_42_22_g287__9945(lt_42_22_n_29 ,n_406 ,lt_42_22_n_3);
  nor lt_42_22_g288__2883(lt_42_22_n_28 ,lt_42_22_n_21 ,n_403);
  nor lt_42_22_g289__2346(lt_42_22_n_27 ,lt_42_22_n_2 ,n_438);
  and lt_42_22_g290__1666(lt_42_22_n_26 ,n_402 ,lt_42_22_n_18);
  nor lt_42_22_g291__7410(lt_42_22_n_25 ,lt_42_22_n_12 ,n_398);
  nor lt_42_22_g292__6417(lt_42_22_n_24 ,lt_42_22_n_17 ,n_446);
  nor lt_42_22_g293__5477(lt_42_22_n_23 ,lt_42_22_n_4 ,n_437);
  nor lt_42_22_g294__2398(lt_42_22_n_22 ,lt_42_22_n_0 ,n_442);
  not lt_42_22_g295(lt_42_22_n_21 ,n_442);
  not lt_42_22_g296(lt_42_22_n_20 ,n_444);
  not lt_42_22_g297(lt_42_22_n_19 ,n_397);
  not lt_42_22_g298(lt_42_22_n_18 ,n_441);
  not lt_42_22_g299(lt_42_22_n_17 ,n_407);
  not lt_42_22_g300(lt_42_22_n_16 ,n_436);
  not lt_42_22_g301(lt_42_22_n_15 ,n_440);
  not lt_42_22_g302(lt_42_22_n_14 ,n_439);
  not lt_42_22_g303(lt_42_22_n_13 ,n_396);
  not lt_42_22_g304(lt_42_22_n_12 ,n_437);
  not lt_42_22_g305(lt_42_22_n_11 ,n_435);
  not lt_42_22_g306(lt_42_22_n_10 ,n_401);
  not lt_42_22_g307(lt_42_22_n_9 ,n_438);
  not lt_42_22_g308(lt_42_22_n_8 ,n_405);
  not lt_42_22_g309(lt_42_22_n_7 ,n_421);
  not lt_42_22_g310(lt_42_22_n_6 ,n_400);
  not lt_42_22_g311(lt_42_22_n_5 ,n_446);
  not lt_42_22_g312(lt_42_22_n_4 ,n_398);
  not lt_42_22_g313(lt_42_22_n_3 ,n_445);
  not lt_42_22_g314(lt_42_22_n_2 ,n_399);
  not lt_42_22_g315(lt_42_22_n_1 ,n_443);
  not lt_42_22_g316(lt_42_22_n_0 ,n_403);
  or lt_43_22_g242__5107(out2 ,lt_43_22_n_33 ,lt_43_22_n_73);
  nor lt_43_22_g243__6260(lt_43_22_n_73 ,lt_43_22_n_24 ,lt_43_22_n_72);
  or lt_43_22_g244__4319(lt_43_22_n_72 ,lt_43_22_n_41 ,lt_43_22_n_71);
  nor lt_43_22_g245__8428(lt_43_22_n_71 ,lt_43_22_n_29 ,lt_43_22_n_70);
  nor lt_43_22_g246__5526(lt_43_22_n_70 ,lt_43_22_n_40 ,lt_43_22_n_69);
  nor lt_43_22_g247__6783(lt_43_22_n_69 ,lt_43_22_n_36 ,lt_43_22_n_68);
  nor lt_43_22_g248__3680(lt_43_22_n_68 ,lt_43_22_n_35 ,lt_43_22_n_67);
  nor lt_43_22_g249__1617(lt_43_22_n_67 ,lt_43_22_n_31 ,lt_43_22_n_66);
  nor lt_43_22_g250__2802(lt_43_22_n_66 ,lt_43_22_n_28 ,lt_43_22_n_65);
  nor lt_43_22_g251__1705(lt_43_22_n_65 ,lt_43_22_n_22 ,lt_43_22_n_64);
  nor lt_43_22_g252__5122(lt_43_22_n_64 ,lt_43_22_n_44 ,lt_43_22_n_63);
  nor lt_43_22_g253__8246(lt_43_22_n_63 ,lt_43_22_n_26 ,lt_43_22_n_62);
  nor lt_43_22_g254__7098(lt_43_22_n_62 ,lt_43_22_n_37 ,lt_43_22_n_61);
  nor lt_43_22_g255__6131(lt_43_22_n_61 ,lt_43_22_n_38 ,lt_43_22_n_60);
  nor lt_43_22_g256__1881(lt_43_22_n_60 ,lt_43_22_n_34 ,lt_43_22_n_59);
  nor lt_43_22_g257__5115(lt_43_22_n_59 ,lt_43_22_n_32 ,lt_43_22_n_58);
  nor lt_43_22_g258__7482(lt_43_22_n_58 ,lt_43_22_n_30 ,lt_43_22_n_57);
  nor lt_43_22_g259__4733(lt_43_22_n_57 ,lt_43_22_n_27 ,lt_43_22_n_56);
  nor lt_43_22_g260__6161(lt_43_22_n_56 ,lt_43_22_n_25 ,lt_43_22_n_55);
  nor lt_43_22_g261__9315(lt_43_22_n_55 ,lt_43_22_n_23 ,lt_43_22_n_54);
  nor lt_43_22_g262__9945(lt_43_22_n_54 ,lt_43_22_n_39 ,lt_43_22_n_53);
  nor lt_43_22_g263__2883(lt_43_22_n_53 ,lt_43_22_n_43 ,lt_43_22_n_52);
  nor lt_43_22_g264__2346(lt_43_22_n_52 ,lt_43_22_n_42 ,lt_43_22_n_51);
  nor lt_43_22_g265__1666(lt_43_22_n_51 ,lt_43_22_n_45 ,lt_43_22_n_50);
  nor lt_43_22_g266__7410(lt_43_22_n_50 ,lt_43_22_n_48 ,lt_43_22_n_49);
  nor lt_43_22_g267__6417(lt_43_22_n_49 ,n_369 ,lt_43_22_n_47);
  and lt_43_22_g268__5477(lt_43_22_n_48 ,n_382 ,lt_43_22_n_46);
  nor lt_43_22_g269__2398(lt_43_22_n_47 ,n_382 ,lt_43_22_n_46);
  nor lt_43_22_g270__5107(lt_43_22_n_45 ,lt_43_22_n_13 ,n_383);
  nor lt_43_22_g271__6260(lt_43_22_n_44 ,lt_43_22_n_18 ,n_376);
  nor lt_43_22_g272__4319(lt_43_22_n_43 ,lt_43_22_n_19 ,n_384);
  nor lt_43_22_g273__8428(lt_43_22_n_42 ,lt_43_22_n_11 ,n_370);
  nor lt_43_22_g274__5526(lt_43_22_n_41 ,lt_43_22_n_3 ,n_380);
  nor lt_43_22_g275__6783(lt_43_22_n_40 ,lt_43_22_n_20 ,n_379);
  nor lt_43_22_g276__3680(lt_43_22_n_39 ,lt_43_22_n_16 ,n_371);
  nor lt_43_22_g277__1617(lt_43_22_n_38 ,lt_43_22_n_10 ,n_388);
  nor lt_43_22_g278__2802(lt_43_22_n_37 ,lt_43_22_n_15 ,n_375);
  nor lt_43_22_g279__1705(lt_43_22_n_36 ,lt_43_22_n_8 ,n_392);
  nor lt_43_22_g280__5122(lt_43_22_n_35 ,lt_43_22_n_1 ,n_378);
  or lt_43_22_g281__8246(lt_43_22_n_46 ,lt_43_22_n_7 ,n_460);
  nor lt_43_22_g282__7098(lt_43_22_n_34 ,lt_43_22_n_14 ,n_374);
  nor lt_43_22_g283__6131(lt_43_22_n_33 ,lt_43_22_n_5 ,n_381);
  nor lt_43_22_g284__1881(lt_43_22_n_32 ,lt_43_22_n_6 ,n_387);
  and lt_43_22_g285__5115(lt_43_22_n_31 ,n_378 ,lt_43_22_n_1);
  nor lt_43_22_g286__7482(lt_43_22_n_30 ,lt_43_22_n_9 ,n_373);
  and lt_43_22_g287__4733(lt_43_22_n_29 ,n_380 ,lt_43_22_n_3);
  nor lt_43_22_g288__6161(lt_43_22_n_28 ,lt_43_22_n_21 ,n_377);
  nor lt_43_22_g289__9315(lt_43_22_n_27 ,lt_43_22_n_2 ,n_386);
  and lt_43_22_g290__9945(lt_43_22_n_26 ,n_376 ,lt_43_22_n_18);
  nor lt_43_22_g291__2883(lt_43_22_n_25 ,lt_43_22_n_12 ,n_372);
  nor lt_43_22_g292__2346(lt_43_22_n_24 ,lt_43_22_n_17 ,n_394);
  nor lt_43_22_g293__1666(lt_43_22_n_23 ,lt_43_22_n_4 ,n_385);
  nor lt_43_22_g294__7410(lt_43_22_n_22 ,lt_43_22_n_0 ,n_390);
  not lt_43_22_g295(lt_43_22_n_21 ,n_390);
  not lt_43_22_g296(lt_43_22_n_20 ,n_392);
  not lt_43_22_g297(lt_43_22_n_19 ,n_371);
  not lt_43_22_g298(lt_43_22_n_18 ,n_389);
  not lt_43_22_g299(lt_43_22_n_17 ,n_381);
  not lt_43_22_g300(lt_43_22_n_16 ,n_384);
  not lt_43_22_g301(lt_43_22_n_15 ,n_388);
  not lt_43_22_g302(lt_43_22_n_14 ,n_387);
  not lt_43_22_g303(lt_43_22_n_13 ,n_370);
  not lt_43_22_g304(lt_43_22_n_12 ,n_385);
  not lt_43_22_g305(lt_43_22_n_11 ,n_383);
  not lt_43_22_g306(lt_43_22_n_10 ,n_375);
  not lt_43_22_g307(lt_43_22_n_9 ,n_386);
  not lt_43_22_g308(lt_43_22_n_8 ,n_379);
  not lt_43_22_g309(lt_43_22_n_7 ,n_421);
  not lt_43_22_g310(lt_43_22_n_6 ,n_374);
  not lt_43_22_g311(lt_43_22_n_5 ,n_394);
  not lt_43_22_g312(lt_43_22_n_4 ,n_372);
  not lt_43_22_g313(lt_43_22_n_3 ,n_393);
  not lt_43_22_g314(lt_43_22_n_2 ,n_373);
  not lt_43_22_g315(lt_43_22_n_1 ,n_391);
  not lt_43_22_g316(lt_43_22_n_0 ,n_377);
  or lt_44_22_g242__6417(out3 ,lt_44_22_n_33 ,lt_44_22_n_73);
  nor lt_44_22_g243__5477(lt_44_22_n_73 ,lt_44_22_n_24 ,lt_44_22_n_72);
  or lt_44_22_g244__2398(lt_44_22_n_72 ,lt_44_22_n_41 ,lt_44_22_n_71);
  nor lt_44_22_g245__5107(lt_44_22_n_71 ,lt_44_22_n_29 ,lt_44_22_n_70);
  nor lt_44_22_g246__6260(lt_44_22_n_70 ,lt_44_22_n_40 ,lt_44_22_n_69);
  nor lt_44_22_g247__4319(lt_44_22_n_69 ,lt_44_22_n_36 ,lt_44_22_n_68);
  nor lt_44_22_g248__8428(lt_44_22_n_68 ,lt_44_22_n_35 ,lt_44_22_n_67);
  nor lt_44_22_g249__5526(lt_44_22_n_67 ,lt_44_22_n_31 ,lt_44_22_n_66);
  nor lt_44_22_g250__6783(lt_44_22_n_66 ,lt_44_22_n_28 ,lt_44_22_n_65);
  nor lt_44_22_g251__3680(lt_44_22_n_65 ,lt_44_22_n_22 ,lt_44_22_n_64);
  nor lt_44_22_g252__1617(lt_44_22_n_64 ,lt_44_22_n_44 ,lt_44_22_n_63);
  nor lt_44_22_g253__2802(lt_44_22_n_63 ,lt_44_22_n_26 ,lt_44_22_n_62);
  nor lt_44_22_g254__1705(lt_44_22_n_62 ,lt_44_22_n_37 ,lt_44_22_n_61);
  nor lt_44_22_g255__5122(lt_44_22_n_61 ,lt_44_22_n_38 ,lt_44_22_n_60);
  nor lt_44_22_g256__8246(lt_44_22_n_60 ,lt_44_22_n_34 ,lt_44_22_n_59);
  nor lt_44_22_g257__7098(lt_44_22_n_59 ,lt_44_22_n_32 ,lt_44_22_n_58);
  nor lt_44_22_g258__6131(lt_44_22_n_58 ,lt_44_22_n_30 ,lt_44_22_n_57);
  nor lt_44_22_g259__1881(lt_44_22_n_57 ,lt_44_22_n_27 ,lt_44_22_n_56);
  nor lt_44_22_g260__5115(lt_44_22_n_56 ,lt_44_22_n_25 ,lt_44_22_n_55);
  nor lt_44_22_g261__7482(lt_44_22_n_55 ,lt_44_22_n_23 ,lt_44_22_n_54);
  nor lt_44_22_g262__4733(lt_44_22_n_54 ,lt_44_22_n_39 ,lt_44_22_n_53);
  nor lt_44_22_g263__6161(lt_44_22_n_53 ,lt_44_22_n_43 ,lt_44_22_n_52);
  nor lt_44_22_g264__9315(lt_44_22_n_52 ,lt_44_22_n_42 ,lt_44_22_n_51);
  nor lt_44_22_g265__9945(lt_44_22_n_51 ,lt_44_22_n_45 ,lt_44_22_n_50);
  nor lt_44_22_g266__2883(lt_44_22_n_50 ,lt_44_22_n_48 ,lt_44_22_n_49);
  nor lt_44_22_g267__2346(lt_44_22_n_49 ,n_343 ,lt_44_22_n_47);
  and lt_44_22_g268__1666(lt_44_22_n_48 ,n_356 ,lt_44_22_n_46);
  nor lt_44_22_g269__7410(lt_44_22_n_47 ,n_356 ,lt_44_22_n_46);
  nor lt_44_22_g270__6417(lt_44_22_n_45 ,lt_44_22_n_13 ,n_357);
  nor lt_44_22_g271__5477(lt_44_22_n_44 ,lt_44_22_n_18 ,n_350);
  nor lt_44_22_g272__2398(lt_44_22_n_43 ,lt_44_22_n_19 ,n_358);
  nor lt_44_22_g273__5107(lt_44_22_n_42 ,lt_44_22_n_11 ,n_344);
  nor lt_44_22_g274__6260(lt_44_22_n_41 ,lt_44_22_n_3 ,n_354);
  nor lt_44_22_g275__4319(lt_44_22_n_40 ,lt_44_22_n_20 ,n_353);
  nor lt_44_22_g276__8428(lt_44_22_n_39 ,lt_44_22_n_16 ,n_345);
  nor lt_44_22_g277__5526(lt_44_22_n_38 ,lt_44_22_n_10 ,n_362);
  nor lt_44_22_g278__6783(lt_44_22_n_37 ,lt_44_22_n_15 ,n_349);
  nor lt_44_22_g279__3680(lt_44_22_n_36 ,lt_44_22_n_8 ,n_366);
  nor lt_44_22_g280__1617(lt_44_22_n_35 ,lt_44_22_n_1 ,n_352);
  or lt_44_22_g281__2802(lt_44_22_n_46 ,lt_44_22_n_7 ,n_460);
  nor lt_44_22_g282__1705(lt_44_22_n_34 ,lt_44_22_n_14 ,n_348);
  nor lt_44_22_g283__5122(lt_44_22_n_33 ,lt_44_22_n_5 ,n_355);
  nor lt_44_22_g284__8246(lt_44_22_n_32 ,lt_44_22_n_6 ,n_361);
  and lt_44_22_g285__7098(lt_44_22_n_31 ,n_352 ,lt_44_22_n_1);
  nor lt_44_22_g286__6131(lt_44_22_n_30 ,lt_44_22_n_9 ,n_347);
  and lt_44_22_g287__1881(lt_44_22_n_29 ,n_354 ,lt_44_22_n_3);
  nor lt_44_22_g288__5115(lt_44_22_n_28 ,lt_44_22_n_21 ,n_351);
  nor lt_44_22_g289__7482(lt_44_22_n_27 ,lt_44_22_n_2 ,n_360);
  and lt_44_22_g290__4733(lt_44_22_n_26 ,n_350 ,lt_44_22_n_18);
  nor lt_44_22_g291__6161(lt_44_22_n_25 ,lt_44_22_n_12 ,n_346);
  nor lt_44_22_g292__9315(lt_44_22_n_24 ,lt_44_22_n_17 ,n_368);
  nor lt_44_22_g293__9945(lt_44_22_n_23 ,lt_44_22_n_4 ,n_359);
  nor lt_44_22_g294__2883(lt_44_22_n_22 ,lt_44_22_n_0 ,n_364);
  not lt_44_22_g295(lt_44_22_n_21 ,n_364);
  not lt_44_22_g296(lt_44_22_n_20 ,n_366);
  not lt_44_22_g297(lt_44_22_n_19 ,n_345);
  not lt_44_22_g298(lt_44_22_n_18 ,n_363);
  not lt_44_22_g299(lt_44_22_n_17 ,n_355);
  not lt_44_22_g300(lt_44_22_n_16 ,n_358);
  not lt_44_22_g301(lt_44_22_n_15 ,n_362);
  not lt_44_22_g302(lt_44_22_n_14 ,n_361);
  not lt_44_22_g303(lt_44_22_n_13 ,n_344);
  not lt_44_22_g304(lt_44_22_n_12 ,n_359);
  not lt_44_22_g305(lt_44_22_n_11 ,n_357);
  not lt_44_22_g306(lt_44_22_n_10 ,n_349);
  not lt_44_22_g307(lt_44_22_n_9 ,n_360);
  not lt_44_22_g308(lt_44_22_n_8 ,n_353);
  not lt_44_22_g309(lt_44_22_n_7 ,n_421);
  not lt_44_22_g310(lt_44_22_n_6 ,n_348);
  not lt_44_22_g311(lt_44_22_n_5 ,n_368);
  not lt_44_22_g312(lt_44_22_n_4 ,n_346);
  not lt_44_22_g313(lt_44_22_n_3 ,n_367);
  not lt_44_22_g314(lt_44_22_n_2 ,n_347);
  not lt_44_22_g315(lt_44_22_n_1 ,n_365);
  not lt_44_22_g316(lt_44_22_n_0 ,n_351);
  or sub_32_21_g297__2346(sub_32_21_n_90 ,sub_32_21_n_32 ,sub_32_21_n_88);
  xnor sub_32_21_g298__1666(n_471 ,sub_32_21_n_87 ,sub_32_21_n_54);
  and sub_32_21_g299__7410(sub_32_21_n_88 ,sub_32_21_n_23 ,sub_32_21_n_87);
  and sub_32_21_g300__6417(sub_32_21_n_87 ,sub_32_21_n_41 ,sub_32_21_n_85);
  xnor sub_32_21_g301__5477(n_470 ,sub_32_21_n_84 ,sub_32_21_n_55);
  or sub_32_21_g302__2398(sub_32_21_n_85 ,sub_32_21_n_27 ,sub_32_21_n_84);
  and sub_32_21_g303__5107(sub_32_21_n_84 ,sub_32_21_n_35 ,sub_32_21_n_82);
  xnor sub_32_21_g304__6260(n_469 ,sub_32_21_n_81 ,sub_32_21_n_56);
  or sub_32_21_g305__4319(sub_32_21_n_82 ,sub_32_21_n_37 ,sub_32_21_n_81);
  and sub_32_21_g306__8428(sub_32_21_n_81 ,sub_32_21_n_36 ,sub_32_21_n_79);
  xnor sub_32_21_g307__5526(n_468 ,sub_32_21_n_78 ,sub_32_21_n_46);
  or sub_32_21_g308__6783(sub_32_21_n_79 ,sub_32_21_n_30 ,sub_32_21_n_78);
  and sub_32_21_g309__3680(sub_32_21_n_78 ,sub_32_21_n_26 ,sub_32_21_n_76);
  xnor sub_32_21_g310__1617(n_467 ,sub_32_21_n_75 ,sub_32_21_n_51);
  or sub_32_21_g311__2802(sub_32_21_n_76 ,sub_32_21_n_43 ,sub_32_21_n_75);
  and sub_32_21_g312__1705(sub_32_21_n_75 ,sub_32_21_n_39 ,sub_32_21_n_73);
  xnor sub_32_21_g313__5122(n_466 ,sub_32_21_n_72 ,sub_32_21_n_50);
  or sub_32_21_g314__8246(sub_32_21_n_73 ,sub_32_21_n_44 ,sub_32_21_n_72);
  and sub_32_21_g315__7098(sub_32_21_n_72 ,sub_32_21_n_38 ,sub_32_21_n_70);
  xnor sub_32_21_g316__6131(n_465 ,sub_32_21_n_69 ,sub_32_21_n_49);
  or sub_32_21_g317__1881(sub_32_21_n_70 ,sub_32_21_n_40 ,sub_32_21_n_69);
  and sub_32_21_g318__5115(sub_32_21_n_69 ,sub_32_21_n_28 ,sub_32_21_n_67);
  xnor sub_32_21_g319__7482(n_464 ,sub_32_21_n_66 ,sub_32_21_n_48);
  or sub_32_21_g320__4733(sub_32_21_n_67 ,sub_32_21_n_29 ,sub_32_21_n_66);
  and sub_32_21_g321__6161(sub_32_21_n_66 ,sub_32_21_n_34 ,sub_32_21_n_64);
  xnor sub_32_21_g322__9315(n_463 ,sub_32_21_n_63 ,sub_32_21_n_47);
  or sub_32_21_g323__9945(sub_32_21_n_64 ,sub_32_21_n_25 ,sub_32_21_n_63);
  and sub_32_21_g324__2883(sub_32_21_n_63 ,sub_32_21_n_24 ,sub_32_21_n_61);
  xnor sub_32_21_g325__2346(n_462 ,sub_32_21_n_59 ,sub_32_21_n_52);
  or sub_32_21_g326__1666(sub_32_21_n_61 ,sub_32_21_n_33 ,sub_32_21_n_59);
  xnor sub_32_21_g327__7410(n_461 ,sub_32_21_n_45 ,sub_32_21_n_53);
  and sub_32_21_g328__6417(sub_32_21_n_59 ,sub_32_21_n_31 ,sub_32_21_n_58);
  or sub_32_21_g329__5477(sub_32_21_n_58 ,sub_32_21_n_42 ,sub_32_21_n_45);
  xor sub_32_21_g330__2398(sub_32_21_n_57 ,in1[0] ,in2[0]);
  xnor sub_32_21_g331__5107(sub_32_21_n_56 ,in1[9] ,in2[9]);
  xnor sub_32_21_g332__6260(sub_32_21_n_55 ,in1[10] ,in2[10]);
  xnor sub_32_21_g333__4319(sub_32_21_n_54 ,in1[11] ,in2[11]);
  xnor sub_32_21_g334__8428(sub_32_21_n_53 ,in1[1] ,in2[1]);
  xnor sub_32_21_g335__5526(sub_32_21_n_52 ,in1[2] ,in2[2]);
  xnor sub_32_21_g336__6783(sub_32_21_n_51 ,in1[7] ,in2[7]);
  xnor sub_32_21_g337__3680(sub_32_21_n_50 ,in1[6] ,in2[6]);
  xnor sub_32_21_g338__1617(sub_32_21_n_49 ,in1[5] ,in2[5]);
  xnor sub_32_21_g339__2802(sub_32_21_n_48 ,in1[4] ,in2[4]);
  xnor sub_32_21_g340__1705(sub_32_21_n_47 ,in1[3] ,in2[3]);
  xnor sub_32_21_g341__5122(sub_32_21_n_46 ,in1[8] ,in2[8]);
  nor sub_32_21_g342__8246(sub_32_21_n_44 ,sub_32_21_n_7 ,in1[6]);
  nor sub_32_21_g343__7098(sub_32_21_n_43 ,sub_32_21_n_18 ,in1[7]);
  nor sub_32_21_g344__6131(sub_32_21_n_42 ,sub_32_21_n_9 ,in1[1]);
  or sub_32_21_g345__1881(sub_32_21_n_41 ,sub_32_21_n_3 ,in2[10]);
  nor sub_32_21_g346__5115(sub_32_21_n_40 ,sub_32_21_n_4 ,in1[5]);
  or sub_32_21_g347__7482(sub_32_21_n_39 ,sub_32_21_n_22 ,in2[6]);
  or sub_32_21_g348__4733(sub_32_21_n_38 ,sub_32_21_n_16 ,in2[5]);
  nor sub_32_21_g349__6161(sub_32_21_n_37 ,sub_32_21_n_15 ,in1[9]);
  or sub_32_21_g350__9315(sub_32_21_n_36 ,sub_32_21_n_8 ,in2[8]);
  or sub_32_21_g351__9945(sub_32_21_n_35 ,sub_32_21_n_12 ,in2[9]);
  and sub_32_21_g352__2883(sub_32_21_n_45 ,in2[0] ,sub_32_21_n_11);
  or sub_32_21_g353__2346(sub_32_21_n_34 ,sub_32_21_n_13 ,in2[3]);
  nor sub_32_21_g354__1666(sub_32_21_n_33 ,sub_32_21_n_14 ,in1[2]);
  nor sub_32_21_g355__7410(sub_32_21_n_32 ,sub_32_21_n_20 ,in2[11]);
  or sub_32_21_g356__6417(sub_32_21_n_31 ,sub_32_21_n_10 ,in2[1]);
  and sub_32_21_g357__5477(sub_32_21_n_30 ,in2[8] ,sub_32_21_n_8);
  nor sub_32_21_g358__2398(sub_32_21_n_29 ,sub_32_21_n_2 ,in1[4]);
  or sub_32_21_g359__5107(sub_32_21_n_28 ,sub_32_21_n_21 ,in2[4]);
  and sub_32_21_g360__6260(sub_32_21_n_27 ,in2[10] ,sub_32_21_n_3);
  or sub_32_21_g361__4319(sub_32_21_n_26 ,sub_32_21_n_5 ,in2[7]);
  nor sub_32_21_g362__8428(sub_32_21_n_25 ,sub_32_21_n_17 ,in1[3]);
  or sub_32_21_g363__5526(sub_32_21_n_24 ,sub_32_21_n_19 ,in2[2]);
  or sub_32_21_g364__6783(sub_32_21_n_23 ,sub_32_21_n_6 ,in1[11]);
  not sub_32_21_g365(sub_32_21_n_22 ,in1[6]);
  not sub_32_21_g366(sub_32_21_n_21 ,in1[4]);
  not sub_32_21_g367(sub_32_21_n_20 ,in1[11]);
  not sub_32_21_g368(sub_32_21_n_19 ,in1[2]);
  not sub_32_21_g369(sub_32_21_n_18 ,in2[7]);
  not sub_32_21_g370(sub_32_21_n_17 ,in2[3]);
  not sub_32_21_g371(sub_32_21_n_16 ,in1[5]);
  not sub_32_21_g372(sub_32_21_n_15 ,in2[9]);
  not sub_32_21_g373(sub_32_21_n_14 ,in2[2]);
  not sub_32_21_g374(sub_32_21_n_13 ,in1[3]);
  not sub_32_21_g375(sub_32_21_n_12 ,in1[9]);
  not sub_32_21_g376(sub_32_21_n_11 ,in1[0]);
  not sub_32_21_g377(sub_32_21_n_10 ,in1[1]);
  not sub_32_21_g378(sub_32_21_n_9 ,in2[1]);
  not sub_32_21_g379(sub_32_21_n_8 ,in1[8]);
  not sub_32_21_g380(sub_32_21_n_7 ,in2[6]);
  not sub_32_21_g381(sub_32_21_n_6 ,in2[11]);
  not sub_32_21_g382(sub_32_21_n_5 ,in1[7]);
  not sub_32_21_g383(sub_32_21_n_4 ,in2[5]);
  not sub_32_21_g384(sub_32_21_n_3 ,in1[10]);
  not sub_32_21_g385(sub_32_21_n_2 ,in2[4]);
  buf sub_32_21_drc_bufs(n_460 ,sub_32_21_n_57);
  buf sub_32_21_drc_bufs386(out5 ,sub_32_21_n_90);
  and sub_33_31_g204__3680(sub_33_31_n_51 ,sub_33_31_n_31 ,sub_33_31_n_49);
  and sub_33_31_g205__1617(sub_33_31_n_50 ,sub_33_31_n_47 ,sub_33_31_n_49);
  not sub_33_31_g206(sub_33_31_n_49 ,sub_33_31_n_48);
  and sub_33_31_g207__2802(sub_33_31_n_48 ,sub_33_31_n_36 ,sub_33_31_n_46);
  or sub_33_31_g208__1705(sub_33_31_n_47 ,sub_33_31_n_36 ,sub_33_31_n_46);
  and sub_33_31_g210__5122(sub_33_31_n_46 ,sub_33_31_n_32 ,sub_33_31_n_45);
  and sub_33_31_g212__8246(sub_33_31_n_45 ,sub_33_31_n_25 ,sub_33_31_n_44);
  and sub_33_31_g214__7098(sub_33_31_n_44 ,sub_33_31_n_29 ,sub_33_31_n_43);
  and sub_33_31_g216__6131(sub_33_31_n_43 ,sub_33_31_n_27 ,sub_33_31_n_42);
  and sub_33_31_g218__1881(sub_33_31_n_42 ,sub_33_31_n_35 ,sub_33_31_n_41);
  and sub_33_31_g220__5115(sub_33_31_n_41 ,sub_33_31_n_26 ,sub_33_31_n_40);
  and sub_33_31_g222__7482(sub_33_31_n_40 ,sub_33_31_n_28 ,sub_33_31_n_39);
  and sub_33_31_g224__4733(sub_33_31_n_39 ,sub_33_31_n_24 ,sub_33_31_n_38);
  and sub_33_31_g226__6161(sub_33_31_n_38 ,sub_33_31_n_30 ,sub_33_31_n_37);
  and sub_33_31_g228__9315(sub_33_31_n_37 ,sub_33_31_n_33 ,sub_33_31_n_34);
  not sub_33_31_g232(sub_33_31_n_36 ,n_471);
  not sub_33_31_drc_bufs243(sub_33_31_n_31 ,out5);
  not sub_33_31_drc_bufs247(sub_33_31_n_24 ,n_463);
  not sub_33_31_drc_bufs251(sub_33_31_n_27 ,n_467);
  not sub_33_31_drc_bufs255(sub_33_31_n_29 ,n_468);
  not sub_33_31_drc_bufs259(sub_33_31_n_28 ,n_464);
  not sub_33_31_drc_bufs263(sub_33_31_n_25 ,n_469);
  not sub_33_31_drc_bufs267(sub_33_31_n_32 ,n_470);
  not sub_33_31_drc_bufs271(sub_33_31_n_33 ,n_461);
  not sub_33_31_drc_bufs275(sub_33_31_n_30 ,n_462);
  not sub_33_31_drc_bufs279(sub_33_31_n_26 ,n_465);
  not sub_33_31_drc_bufs283(sub_33_31_n_35 ,n_466);
  not sub_33_31_drc_bufs287(sub_33_31_n_34 ,n_460);
  buf sub_33_31_drc_bufs290(n_458 ,sub_33_31_n_10);
  buf sub_33_31_drc_bufs291(n_453 ,sub_33_31_n_8);
  buf sub_33_31_drc_bufs292(n_452 ,sub_33_31_n_0);
  buf sub_33_31_drc_bufs293(n_450 ,sub_33_31_n_6);
  buf sub_33_31_drc_bufs294(n_449 ,sub_33_31_n_9);
  buf sub_33_31_drc_bufs295(n_448 ,sub_33_31_n_2);
  buf sub_33_31_drc_bufs296(n_455 ,sub_33_31_n_5);
  buf sub_33_31_drc_bufs297(n_451 ,sub_33_31_n_1);
  buf sub_33_31_drc_bufs298(n_454 ,sub_33_31_n_7);
  buf sub_33_31_drc_bufs299(n_456 ,sub_33_31_n_4);
  buf sub_33_31_drc_bufs300(n_447 ,sub_33_31_n_3);
  buf sub_33_31_drc_bufs301(n_457 ,sub_33_31_n_50);
  buf sub_33_31_drc_bufs302(n_459 ,sub_33_31_n_51);
  xor sub_33_31_g2__9945(sub_33_31_n_10 ,sub_33_31_n_48 ,sub_33_31_n_31);
  xor sub_33_31_g315__2883(sub_33_31_n_9 ,sub_33_31_n_38 ,sub_33_31_n_24);
  xor sub_33_31_g316__2346(sub_33_31_n_8 ,sub_33_31_n_42 ,sub_33_31_n_27);
  xor sub_33_31_g317__1666(sub_33_31_n_7 ,sub_33_31_n_43 ,sub_33_31_n_29);
  xor sub_33_31_g318__7410(sub_33_31_n_6 ,sub_33_31_n_39 ,sub_33_31_n_28);
  xor sub_33_31_g319__6417(sub_33_31_n_5 ,sub_33_31_n_44 ,sub_33_31_n_25);
  xor sub_33_31_g320__5477(sub_33_31_n_4 ,sub_33_31_n_45 ,sub_33_31_n_32);
  xor sub_33_31_g321__2398(sub_33_31_n_3 ,sub_33_31_n_34 ,sub_33_31_n_33);
  xor sub_33_31_g322__5107(sub_33_31_n_2 ,sub_33_31_n_37 ,sub_33_31_n_30);
  xor sub_33_31_g323__6260(sub_33_31_n_1 ,sub_33_31_n_40 ,sub_33_31_n_26);
  xor sub_33_31_g324__4319(sub_33_31_n_0 ,sub_33_31_n_41 ,sub_33_31_n_35);
  or sub_35_21_g297__8428(sub_35_21_n_90 ,sub_35_21_n_32 ,sub_35_21_n_88);
  xnor sub_35_21_g298__5526(n_432 ,sub_35_21_n_87 ,sub_35_21_n_54);
  and sub_35_21_g299__6783(sub_35_21_n_88 ,sub_35_21_n_23 ,sub_35_21_n_87);
  and sub_35_21_g300__3680(sub_35_21_n_87 ,sub_35_21_n_41 ,sub_35_21_n_85);
  xnor sub_35_21_g301__1617(n_431 ,sub_35_21_n_84 ,sub_35_21_n_55);
  or sub_35_21_g302__2802(sub_35_21_n_85 ,sub_35_21_n_27 ,sub_35_21_n_84);
  and sub_35_21_g303__1705(sub_35_21_n_84 ,sub_35_21_n_35 ,sub_35_21_n_82);
  xnor sub_35_21_g304__5122(n_430 ,sub_35_21_n_81 ,sub_35_21_n_56);
  or sub_35_21_g305__8246(sub_35_21_n_82 ,sub_35_21_n_37 ,sub_35_21_n_81);
  and sub_35_21_g306__7098(sub_35_21_n_81 ,sub_35_21_n_36 ,sub_35_21_n_79);
  xnor sub_35_21_g307__6131(n_429 ,sub_35_21_n_78 ,sub_35_21_n_46);
  or sub_35_21_g308__1881(sub_35_21_n_79 ,sub_35_21_n_30 ,sub_35_21_n_78);
  and sub_35_21_g309__5115(sub_35_21_n_78 ,sub_35_21_n_26 ,sub_35_21_n_76);
  xnor sub_35_21_g310__7482(n_428 ,sub_35_21_n_75 ,sub_35_21_n_51);
  or sub_35_21_g311__4733(sub_35_21_n_76 ,sub_35_21_n_43 ,sub_35_21_n_75);
  and sub_35_21_g312__6161(sub_35_21_n_75 ,sub_35_21_n_39 ,sub_35_21_n_73);
  xnor sub_35_21_g313__9315(n_427 ,sub_35_21_n_72 ,sub_35_21_n_50);
  or sub_35_21_g314__9945(sub_35_21_n_73 ,sub_35_21_n_44 ,sub_35_21_n_72);
  and sub_35_21_g315__2883(sub_35_21_n_72 ,sub_35_21_n_38 ,sub_35_21_n_70);
  xnor sub_35_21_g316__2346(n_426 ,sub_35_21_n_69 ,sub_35_21_n_49);
  or sub_35_21_g317__1666(sub_35_21_n_70 ,sub_35_21_n_40 ,sub_35_21_n_69);
  and sub_35_21_g318__7410(sub_35_21_n_69 ,sub_35_21_n_28 ,sub_35_21_n_67);
  xnor sub_35_21_g319__6417(n_425 ,sub_35_21_n_66 ,sub_35_21_n_48);
  or sub_35_21_g320__5477(sub_35_21_n_67 ,sub_35_21_n_29 ,sub_35_21_n_66);
  and sub_35_21_g321__2398(sub_35_21_n_66 ,sub_35_21_n_34 ,sub_35_21_n_64);
  xnor sub_35_21_g322__5107(n_424 ,sub_35_21_n_63 ,sub_35_21_n_47);
  or sub_35_21_g323__6260(sub_35_21_n_64 ,sub_35_21_n_25 ,sub_35_21_n_63);
  and sub_35_21_g324__4319(sub_35_21_n_63 ,sub_35_21_n_24 ,sub_35_21_n_61);
  xnor sub_35_21_g325__8428(n_423 ,sub_35_21_n_59 ,sub_35_21_n_52);
  or sub_35_21_g326__5526(sub_35_21_n_61 ,sub_35_21_n_33 ,sub_35_21_n_59);
  xnor sub_35_21_g327__6783(n_422 ,sub_35_21_n_45 ,sub_35_21_n_53);
  and sub_35_21_g328__3680(sub_35_21_n_59 ,sub_35_21_n_31 ,sub_35_21_n_58);
  or sub_35_21_g329__1617(sub_35_21_n_58 ,sub_35_21_n_42 ,sub_35_21_n_45);
  xor sub_35_21_g330__2802(sub_35_21_n_57 ,in2[0] ,in7[0]);
  xnor sub_35_21_g331__1705(sub_35_21_n_56 ,in2[9] ,in7[9]);
  xnor sub_35_21_g332__5122(sub_35_21_n_55 ,in2[10] ,in7[10]);
  xnor sub_35_21_g333__8246(sub_35_21_n_54 ,in2[11] ,in7[11]);
  xnor sub_35_21_g334__7098(sub_35_21_n_53 ,in2[1] ,in7[1]);
  xnor sub_35_21_g335__6131(sub_35_21_n_52 ,in2[2] ,in7[2]);
  xnor sub_35_21_g336__1881(sub_35_21_n_51 ,in2[7] ,in7[7]);
  xnor sub_35_21_g337__5115(sub_35_21_n_50 ,in2[6] ,in7[6]);
  xnor sub_35_21_g338__7482(sub_35_21_n_49 ,in2[5] ,in7[5]);
  xnor sub_35_21_g339__4733(sub_35_21_n_48 ,in2[4] ,in7[4]);
  xnor sub_35_21_g340__6161(sub_35_21_n_47 ,in2[3] ,in7[3]);
  xnor sub_35_21_g341__9315(sub_35_21_n_46 ,in2[8] ,in7[8]);
  nor sub_35_21_g342__9945(sub_35_21_n_44 ,sub_35_21_n_7 ,in2[6]);
  nor sub_35_21_g343__2883(sub_35_21_n_43 ,sub_35_21_n_18 ,in2[7]);
  nor sub_35_21_g344__2346(sub_35_21_n_42 ,sub_35_21_n_9 ,in2[1]);
  or sub_35_21_g345__1666(sub_35_21_n_41 ,sub_35_21_n_3 ,in7[10]);
  nor sub_35_21_g346__7410(sub_35_21_n_40 ,sub_35_21_n_4 ,in2[5]);
  or sub_35_21_g347__6417(sub_35_21_n_39 ,sub_35_21_n_22 ,in7[6]);
  or sub_35_21_g348__5477(sub_35_21_n_38 ,sub_35_21_n_16 ,in7[5]);
  nor sub_35_21_g349__2398(sub_35_21_n_37 ,sub_35_21_n_15 ,in2[9]);
  or sub_35_21_g350__5107(sub_35_21_n_36 ,sub_35_21_n_8 ,in7[8]);
  or sub_35_21_g351__6260(sub_35_21_n_35 ,sub_35_21_n_12 ,in7[9]);
  and sub_35_21_g352__4319(sub_35_21_n_45 ,in7[0] ,sub_35_21_n_11);
  or sub_35_21_g353__8428(sub_35_21_n_34 ,sub_35_21_n_13 ,in7[3]);
  nor sub_35_21_g354__5526(sub_35_21_n_33 ,sub_35_21_n_14 ,in2[2]);
  nor sub_35_21_g355__6783(sub_35_21_n_32 ,sub_35_21_n_20 ,in7[11]);
  or sub_35_21_g356__3680(sub_35_21_n_31 ,sub_35_21_n_10 ,in7[1]);
  and sub_35_21_g357__1617(sub_35_21_n_30 ,in7[8] ,sub_35_21_n_8);
  nor sub_35_21_g358__2802(sub_35_21_n_29 ,sub_35_21_n_2 ,in2[4]);
  or sub_35_21_g359__1705(sub_35_21_n_28 ,sub_35_21_n_21 ,in7[4]);
  and sub_35_21_g360__5122(sub_35_21_n_27 ,in7[10] ,sub_35_21_n_3);
  or sub_35_21_g361__8246(sub_35_21_n_26 ,sub_35_21_n_5 ,in7[7]);
  nor sub_35_21_g362__7098(sub_35_21_n_25 ,sub_35_21_n_17 ,in2[3]);
  or sub_35_21_g363__6131(sub_35_21_n_24 ,sub_35_21_n_19 ,in7[2]);
  or sub_35_21_g364__1881(sub_35_21_n_23 ,sub_35_21_n_6 ,in2[11]);
  not sub_35_21_g365(sub_35_21_n_22 ,in2[6]);
  not sub_35_21_g366(sub_35_21_n_21 ,in2[4]);
  not sub_35_21_g367(sub_35_21_n_20 ,in2[11]);
  not sub_35_21_g368(sub_35_21_n_19 ,in2[2]);
  not sub_35_21_g369(sub_35_21_n_18 ,in7[7]);
  not sub_35_21_g370(sub_35_21_n_17 ,in7[3]);
  not sub_35_21_g371(sub_35_21_n_16 ,in2[5]);
  not sub_35_21_g372(sub_35_21_n_15 ,in7[9]);
  not sub_35_21_g373(sub_35_21_n_14 ,in7[2]);
  not sub_35_21_g374(sub_35_21_n_13 ,in2[3]);
  not sub_35_21_g375(sub_35_21_n_12 ,in2[9]);
  not sub_35_21_g376(sub_35_21_n_11 ,in2[0]);
  not sub_35_21_g377(sub_35_21_n_10 ,in2[1]);
  not sub_35_21_g378(sub_35_21_n_9 ,in7[1]);
  not sub_35_21_g379(sub_35_21_n_8 ,in2[8]);
  not sub_35_21_g380(sub_35_21_n_7 ,in7[6]);
  not sub_35_21_g381(sub_35_21_n_6 ,in7[11]);
  not sub_35_21_g382(sub_35_21_n_5 ,in2[7]);
  not sub_35_21_g383(sub_35_21_n_4 ,in7[5]);
  not sub_35_21_g384(sub_35_21_n_3 ,in2[10]);
  not sub_35_21_g385(sub_35_21_n_2 ,in7[4]);
  buf sub_35_21_drc_bufs(n_421 ,sub_35_21_n_57);
  buf sub_35_21_drc_bufs386(out4 ,sub_35_21_n_90);
  and sub_36_31_g204__5115(sub_36_31_n_51 ,sub_36_31_n_31 ,sub_36_31_n_49);
  and sub_36_31_g205__7482(sub_36_31_n_50 ,sub_36_31_n_47 ,sub_36_31_n_49);
  not sub_36_31_g206(sub_36_31_n_49 ,sub_36_31_n_48);
  and sub_36_31_g207__4733(sub_36_31_n_48 ,sub_36_31_n_36 ,sub_36_31_n_46);
  or sub_36_31_g208__6161(sub_36_31_n_47 ,sub_36_31_n_36 ,sub_36_31_n_46);
  and sub_36_31_g210__9315(sub_36_31_n_46 ,sub_36_31_n_32 ,sub_36_31_n_45);
  and sub_36_31_g212__9945(sub_36_31_n_45 ,sub_36_31_n_25 ,sub_36_31_n_44);
  and sub_36_31_g214__2883(sub_36_31_n_44 ,sub_36_31_n_29 ,sub_36_31_n_43);
  and sub_36_31_g216__2346(sub_36_31_n_43 ,sub_36_31_n_27 ,sub_36_31_n_42);
  and sub_36_31_g218__1666(sub_36_31_n_42 ,sub_36_31_n_35 ,sub_36_31_n_41);
  and sub_36_31_g220__7410(sub_36_31_n_41 ,sub_36_31_n_26 ,sub_36_31_n_40);
  and sub_36_31_g222__6417(sub_36_31_n_40 ,sub_36_31_n_28 ,sub_36_31_n_39);
  and sub_36_31_g224__5477(sub_36_31_n_39 ,sub_36_31_n_24 ,sub_36_31_n_38);
  and sub_36_31_g226__2398(sub_36_31_n_38 ,sub_36_31_n_30 ,sub_36_31_n_37);
  and sub_36_31_g228__5107(sub_36_31_n_37 ,sub_36_31_n_33 ,sub_36_31_n_34);
  not sub_36_31_g232(sub_36_31_n_36 ,n_432);
  not sub_36_31_drc_bufs243(sub_36_31_n_31 ,out4);
  not sub_36_31_drc_bufs247(sub_36_31_n_24 ,n_424);
  not sub_36_31_drc_bufs251(sub_36_31_n_27 ,n_428);
  not sub_36_31_drc_bufs255(sub_36_31_n_29 ,n_429);
  not sub_36_31_drc_bufs259(sub_36_31_n_28 ,n_425);
  not sub_36_31_drc_bufs263(sub_36_31_n_25 ,n_430);
  not sub_36_31_drc_bufs267(sub_36_31_n_32 ,n_431);
  not sub_36_31_drc_bufs271(sub_36_31_n_33 ,n_422);
  not sub_36_31_drc_bufs275(sub_36_31_n_30 ,n_423);
  not sub_36_31_drc_bufs279(sub_36_31_n_26 ,n_426);
  not sub_36_31_drc_bufs283(sub_36_31_n_35 ,n_427);
  not sub_36_31_drc_bufs287(sub_36_31_n_34 ,n_421);
  buf sub_36_31_drc_bufs290(n_419 ,sub_36_31_n_10);
  buf sub_36_31_drc_bufs291(n_414 ,sub_36_31_n_8);
  buf sub_36_31_drc_bufs292(n_413 ,sub_36_31_n_0);
  buf sub_36_31_drc_bufs293(n_411 ,sub_36_31_n_6);
  buf sub_36_31_drc_bufs294(n_410 ,sub_36_31_n_9);
  buf sub_36_31_drc_bufs295(n_409 ,sub_36_31_n_2);
  buf sub_36_31_drc_bufs296(n_416 ,sub_36_31_n_5);
  buf sub_36_31_drc_bufs297(n_412 ,sub_36_31_n_1);
  buf sub_36_31_drc_bufs298(n_415 ,sub_36_31_n_7);
  buf sub_36_31_drc_bufs299(n_417 ,sub_36_31_n_4);
  buf sub_36_31_drc_bufs300(n_408 ,sub_36_31_n_3);
  buf sub_36_31_drc_bufs301(n_418 ,sub_36_31_n_50);
  buf sub_36_31_drc_bufs302(n_420 ,sub_36_31_n_51);
  xor sub_36_31_g2__6260(sub_36_31_n_10 ,sub_36_31_n_48 ,sub_36_31_n_31);
  xor sub_36_31_g315__4319(sub_36_31_n_9 ,sub_36_31_n_38 ,sub_36_31_n_24);
  xor sub_36_31_g316__8428(sub_36_31_n_8 ,sub_36_31_n_42 ,sub_36_31_n_27);
  xor sub_36_31_g317__5526(sub_36_31_n_7 ,sub_36_31_n_43 ,sub_36_31_n_29);
  xor sub_36_31_g318__6783(sub_36_31_n_6 ,sub_36_31_n_39 ,sub_36_31_n_28);
  xor sub_36_31_g319__3680(sub_36_31_n_5 ,sub_36_31_n_44 ,sub_36_31_n_25);
  xor sub_36_31_g320__1617(sub_36_31_n_4 ,sub_36_31_n_45 ,sub_36_31_n_32);
  xor sub_36_31_g321__2802(sub_36_31_n_3 ,sub_36_31_n_34 ,sub_36_31_n_33);
  xor sub_36_31_g322__1705(sub_36_31_n_2 ,sub_36_31_n_37 ,sub_36_31_n_30);
  xor sub_36_31_g323__5122(sub_36_31_n_1 ,sub_36_31_n_40 ,sub_36_31_n_26);
  xor sub_36_31_g324__8246(sub_36_31_n_0 ,sub_36_31_n_41 ,sub_36_31_n_35);
endmodule
