/* This is a
  Multi line comment
  example */
module addbit (
a,
b,
ci,
sum,
co);

// Input Ports  Single line comment
input           a;
input           b;
input           ci;
// Output ports
output         sum;
output         co;
// Data Types      
wire            a;
wire            b;
wire            ci;
wire            sum;
wire            co; 

endmodule
