module top( 2_n4 , 2_n14 , 2_n23 , 2_n25 , 2_n28 , 2_n32 , 2_n34 , 2_n38 , 2_n40 , 2_n50 , 2_n55 , 2_n58 , 2_n59 , 2_n60 , 2_n63 , 2_n65 );
    input 2_n4 , 2_n23 , 2_n25 , 2_n28 , 2_n32 , 2_n38 , 2_n50 , 2_n55 , 2_n58 , 2_n60 , 2_n63 , 2_n65 ;
    output 2_n14 , 2_n34 , 2_n40 , 2_n59 ;
    wire 2_n0 , 2_n1 , 2_n2 , 2_n3 , 2_n5 , 2_n6 , 2_n7 , 2_n8 , 2_n9 , 2_n10 , 2_n11 , 2_n12 , 2_n13 , 2_n15 , 2_n16 , 2_n17 , 2_n18 , 2_n19 , 2_n20 , 2_n21 , 2_n22 , 2_n24 , 2_n26 , 2_n27 , 2_n29 , 2_n30 , 2_n31 , 2_n33 , 2_n35 , 2_n36 , 2_n37 , 2_n39 , 2_n41 , 2_n42 , 2_n43 , 2_n44 , 2_n45 , 2_n46 , 2_n47 , 2_n48 , 2_n49 , 2_n51 , 2_n52 , 2_n53 , 2_n54 , 2_n56 , 2_n57 , 2_n61 , 2_n62 , 2_n64 , 2_n66 , 2_n67 , 2_n68 ;
assign 2_n49 = ~(2_n47 | 2_n13);
assign 2_n12 = ~(2_n1 ^ 2_n47);
assign 2_n57 = ~(2_n8 ^ 2_n23);
assign 2_n62 = ~(2_n0 | 2_n45);
assign 2_n56 = 2_n37 | 2_n44;
assign 2_n22 = ~(2_n32 & 2_n60);
assign 2_n44 = ~2_n25;
assign 2_n47 = 2_n3 | 2_n19;
assign 2_n46 = 2_n65 | 2_n61;
assign 2_n33 = 2_n53 | 2_n31;
assign 2_n31 = 2_n3 | 2_n44;
assign 2_n66 = 2_n37 | 2_n36;
assign 2_n2 = ~2_n58;
assign 2_n11 = ~2_n7;
assign 2_n51 = ~2_n32;
assign 2_n9 = ~2_n5;
assign 2_n68 = ~(2_n26 ^ 2_n21);
assign 2_n7 = 2_n51 | 2_n44;
assign 2_n42 = ~(2_n23 | 2_n52);
assign 2_n43 = 2_n27 | 2_n64;
assign 2_n64 = ~(2_n42 | 2_n8);
assign 2_n35 = ~(2_n41 ^ 2_n68);
assign 2_n52 = ~2_n33;
assign 2_n29 = 2_n9 | 2_n24;
assign 2_n21 = 2_n15 | 2_n44;
assign 2_n40 = ~(2_n30 | 2_n52);
assign 2_n16 = 2_n10 & 2_n7;
assign 2_n53 = ~2_n4;
assign 2_n45 = 2_n43 & 2_n46;
assign 2_n24 = ~(2_n56 ^ 2_n12);
assign 2_n15 = ~2_n55;
assign 2_n26 = 2_n3 | 2_n2;
assign 2_n19 = ~2_n60;
assign 2_n27 = 2_n23 & 2_n52;
assign 2_n30 = ~(2_n4 | 2_n39);
assign 2_n37 = ~2_n63;
assign 2_n48 = ~(2_n62 ^ 2_n28);
assign 2_n36 = ~2_n38;
assign 2_n13 = 2_n1 & 2_n56;
assign 2_n39 = ~2_n31;
assign 2_n18 = ~(2_n6 ^ 2_n48);
assign 2_n8 = 2_n16 | 2_n5;
assign 2_n67 = ~(2_n17 | 2_n49);
assign 2_n17 = ~(2_n1 | 2_n56);
assign 2_n20 = ~(2_n61 ^ 2_n65);
assign 2_n5 = 2_n54 & 2_n11;
assign 2_n0 = 2_n65 & 2_n61;
assign 2_n14 = ~(2_n43 ^ 2_n20);
assign 2_n41 = ~(2_n22 ^ 2_n66);
assign 2_n10 = ~2_n54;
assign 2_n61 = ~(2_n5 ^ 2_n24);
assign 2_n1 = 2_n51 | 2_n36;
assign 2_n54 = 2_n50 & 2_n38;
assign 2_n59 = ~(2_n35 ^ 2_n18);
assign 2_n6 = ~(2_n67 ^ 2_n29);
assign 2_n3 = ~2_n50;
assign 2_n34 = ~(2_n33 ^ 2_n57);
endmodule
