module top( n45 , n112 , n137 , n159 , n217 , n226 , n381 , n397 , n405 , n447 , n503 , n521 , n533 , n615 , n658 , n671 , n753 , n783 , n806 , n837 , n844 , n911 , n992 , n996 , n1020 , n1067 , n1094 , n1097 , n1136 , n1138 , n1198 , n1199 , n1209 , n1269 , n1333 , n1353 , n1357 , n1471 , n1478 , n1510 , n1512 , n1523 , n1564 , n1576 , n1658 , n1798 , n1835 , n1847 , n1906 , n1980 , n2024 , n2087 , n2096 , n2131 , n2226 , n2253 , n2278 , n2301 , n2316 , n2347 , n2383 , n2393 , n2425 , n2431 , n2433 , n2434 , n2464 , n2498 , n2507 , n2508 , n2509 , n2512 , n2515 , n2522 , n2530 , n2551 , n2558 , n2564 , n2577 , n2581 , n2585 , n2624 , n2679 , n2708 , n2749 , n2802 , n2818 , n2879 , n2902 , n3022 , n3071 , n3124 , n3146 , n3172 , n3214 , n3230 , n3272 , n3287 , n3339 , n3342 , n3456 , n3602 , n3616 , n3627 , n3654 , n3661 , n3677 , n3719 , n3754 , n3842 , n3849 , n3865 , n3932 , n3986 , n3992 , n4005 , n4086 , n4088 , n4094 , n4141 , n4155 , n4159 , n4187 , n4189 , n4190 , n4203 , n4226 , n4230 , n4300 , n4312 , n4326 , n4333 , n4370 , n4378 , n4397 , n4436 , n4499 , n4516 , n4553 , n4634 , n4686 , n4689 , n4722 , n4733 , n4757 , n4805 , n4817 , n4826 , n4828 , n4903 , n4921 , n4928 , n4938 , n4970 , n4971 , n5030 , n5034 , n5069 , n5094 , n5105 , n5132 , n5153 , n5191 , n5198 , n5212 , n5240 , n5257 , n5283 , n5305 , n5314 , n5319 , n5320 , n5331 , n5411 , n5435 , n5579 , n5641 , n5645 , n5670 , n5693 , n5694 , n5760 , n5767 , n5798 , n5814 , n5857 , n5860 , n5934 , n5964 , n6016 , n6038 , n6089 , n6126 , n6192 , n6254 , n6273 , n6294 , n6358 , n6359 , n6429 , n6431 , n6441 , n6445 , n6578 , n6604 , n6611 , n6645 , n6687 , n6689 , n6703 , n6742 , n6770 , n6776 , n6797 , n6806 , n6809 , n6822 , n6826 , n6860 , n6877 , n6986 , n7159 , n7160 , n7193 , n7236 , n7265 , n7270 , n7294 , n7320 , n7354 , n7388 , n7436 , n7456 , n7500 , n7523 , n7546 , n7568 , n7610 , n7646 , n7676 , n7690 , n7730 , n7733 , n7823 , n7862 , n7891 , n7946 , n7965 , n7966 , n7981 , n8028 , n8065 , n8100 , n8138 , n8202 , n8236 , n8276 , n8303 , n8336 , n8384 , n8398 , n8433 , n8476 , n8595 , n8665 , n8717 , n8759 , n8819 , n9080 , n9111 , n9137 , n9189 , n9195 , n9241 , n9387 , n9400 , n9457 , n9571 , n9578 , n9583 , n9637 , n9640 , n9706 , n9725 , n9756 , n9763 , n9767 , n9820 , n9920 , n9938 , n9956 , n10022 , n10174 , n10217 , n10223 , n10278 , n10327 , n10391 , n10439 , n10451 , n10476 , n10510 , n10545 , n10547 , n10589 , n10644 , n10678 , n10685 , n10695 , n10789 , n10848 , n10851 , n10898 , n10913 , n10928 , n10949 , n10965 , n10990 , n11023 , n11153 , n11216 , n11222 , n11257 , n11296 , n11311 , n11326 , n11407 , n11423 , n11478 , n11536 , n11662 , n11707 , n11728 , n11755 , n11757 , n11780 , n11791 , n11821 , n11876 , n11877 , n11892 , n11917 , n11919 , n11922 , n11967 , n11999 , n12000 , n12005 , n12014 , n12020 , n12025 , n12044 , n12069 , n12076 , n12111 , n12145 , n12221 , n12247 , n12299 , n12391 , n12444 , n12489 , n12511 , n12591 , n12648 , n12704 , n12705 , n12706 , n12709 , n12720 , n12753 , n12777 , n12807 , n12826 , n12925 , n12947 );
    input n45 , n137 , n159 , n217 , n405 , n447 , n503 , n521 , n533 , n615 , n753 , n783 , n806 , n996 , n1067 , n1094 , n1097 , n1198 , n1199 , n1209 , n1333 , n1353 , n1357 , n1471 , n1478 , n1510 , n1512 , n1564 , n1576 , n1798 , n1835 , n1906 , n1980 , n2024 , n2087 , n2226 , n2253 , n2278 , n2347 , n2393 , n2433 , n2464 , n2498 , n2507 , n2508 , n2509 , n2512 , n2515 , n2522 , n2530 , n2551 , n2558 , n2564 , n2577 , n2585 , n2749 , n2802 , n2879 , n3022 , n3146 , n3172 , n3342 , n3602 , n3616 , n3627 , n3719 , n3754 , n3842 , n3865 , n3932 , n3986 , n3992 , n4005 , n4086 , n4094 , n4141 , n4187 , n4189 , n4190 , n4203 , n4312 , n4370 , n4436 , n4499 , n4516 , n4634 , n4722 , n4805 , n4817 , n4826 , n4828 , n4903 , n4921 , n4928 , n4938 , n4970 , n5069 , n5105 , n5153 , n5198 , n5212 , n5240 , n5283 , n5305 , n5314 , n5319 , n5320 , n5331 , n5579 , n5645 , n5694 , n5760 , n5767 , n5798 , n5814 , n5857 , n5860 , n5964 , n6016 , n6038 , n6126 , n6254 , n6294 , n6358 , n6359 , n6429 , n6431 , n6441 , n6578 , n6604 , n6611 , n6687 , n6703 , n6770 , n6776 , n6797 , n6806 , n6826 , n6877 , n6986 , n7159 , n7160 , n7236 , n7265 , n7270 , n7294 , n7320 , n7354 , n7388 , n7436 , n7456 , n7500 , n7523 , n7546 , n7610 , n7646 , n7690 , n7730 , n7733 , n7823 , n7862 , n7891 , n7946 , n7965 , n8028 , n8065 , n8236 , n8276 , n8336 , n8384 , n8433 , n8476 , n8595 , n8665 , n8717 , n8759 , n8819 , n9080 , n9111 , n9189 , n9195 , n9241 , n9400 , n9457 , n9583 , n9637 , n9640 , n9725 , n9763 , n9920 , n9956 , n10022 , n10174 , n10217 , n10223 , n10278 , n10327 , n10391 , n10439 , n10451 , n10510 , n10545 , n10547 , n10644 , n10678 , n10685 , n10848 , n10898 , n10928 , n10965 , n10990 , n11023 , n11153 , n11222 , n11257 , n11296 , n11311 , n11407 , n11423 , n11478 , n11536 , n11662 , n11728 , n11757 , n11791 , n11821 , n11876 , n11877 , n11892 , n11917 , n11922 , n11967 , n11999 , n12000 , n12025 , n12044 , n12069 , n12145 , n12221 , n12247 , n12299 , n12391 , n12489 , n12511 , n12591 , n12648 , n12704 , n12705 , n12706 , n12709 , n12720 , n12753 , n12777 , n12826 , n12925 , n12947 ;
    output n112 , n226 , n381 , n397 , n658 , n671 , n837 , n844 , n911 , n992 , n1020 , n1136 , n1138 , n1269 , n1523 , n1658 , n1847 , n2096 , n2131 , n2301 , n2316 , n2383 , n2425 , n2431 , n2434 , n2581 , n2624 , n2679 , n2708 , n2818 , n2902 , n3071 , n3124 , n3214 , n3230 , n3272 , n3287 , n3339 , n3456 , n3654 , n3661 , n3677 , n3849 , n4088 , n4155 , n4159 , n4226 , n4230 , n4300 , n4326 , n4333 , n4378 , n4397 , n4553 , n4686 , n4689 , n4733 , n4757 , n4971 , n5030 , n5034 , n5094 , n5132 , n5191 , n5257 , n5411 , n5435 , n5641 , n5670 , n5693 , n5934 , n6089 , n6192 , n6273 , n6445 , n6645 , n6689 , n6742 , n6809 , n6822 , n6860 , n7193 , n7568 , n7676 , n7966 , n7981 , n8100 , n8138 , n8202 , n8303 , n8398 , n9137 , n9387 , n9571 , n9578 , n9706 , n9756 , n9767 , n9820 , n9938 , n10476 , n10589 , n10695 , n10789 , n10851 , n10913 , n10949 , n11216 , n11326 , n11707 , n11755 , n11780 , n11919 , n12005 , n12014 , n12020 , n12076 , n12111 , n12444 , n12807 ;
    wire n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n838 , n839 , n840 , n841 , n842 , n843 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n993 , n994 , n995 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1095 , n1096 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1137 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1354 , n1355 , n1356 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1511 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2426 , n2427 , n2428 , n2429 , n2430 , n2432 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2510 , n2511 , n2513 , n2514 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2559 , n2560 , n2561 , n2562 , n2563 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2578 , n2579 , n2580 , n2582 , n2583 , n2584 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3340 , n3341 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3987 , n3988 , n3989 , n3990 , n3991 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4087 , n4089 , n4090 , n4091 , n4092 , n4093 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4156 , n4157 , n4158 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4188 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4227 , n4228 , n4229 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4687 , n4688 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4827 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5031 , n5032 , n5033 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5315 , n5316 , n5317 , n5318 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5642 , n5643 , n5644 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5858 , n5859 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6430 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6442 , n6443 , n6444 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6688 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6771 , n6772 , n6773 , n6774 , n6775 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6807 , n6808 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6823 , n6824 , n6825 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7266 , n7267 , n7268 , n7269 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7731 , n7732 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9190 , n9191 , n9192 , n9193 , n9194 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9579 , n9580 , n9581 , n9582 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9638 , n9639 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9764 , n9765 , n9766 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10218 , n10219 , n10220 , n10221 , n10222 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10546 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10849 , n10850 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11217 , n11218 , n11219 , n11220 , n11221 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11756 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11918 , n11920 , n11921 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n12001 , n12002 , n12003 , n12004 , n12006 , n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12015 , n12016 , n12017 , n12018 , n12019 , n12021 , n12022 , n12023 , n12024 , n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , n12701 , n12702 , n12703 , n12707 , n12708 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , n12750 , n12751 , n12752 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12808 , n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12827 , n12828 , n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , n12926 , n12927 , n12928 , n12929 , n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , n12948 , n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , n12960 ;
assign n2141 = n2530 & n521;
assign n206 = ~(n491 ^ n5906);
assign n3102 = n4112 & n2282;
assign n2523 = n12144 | n5251;
assign n2468 = n491 | n9006;
assign n5935 = ~(n5205 | n1662);
assign n12452 = n3831 & n6309;
assign n3584 = n9389 | n6402;
assign n12769 = ~(n12488 ^ n2077);
assign n9132 = ~(n8037 ^ n4937);
assign n8628 = ~(n8093 ^ n65);
assign n7698 = ~(n8387 ^ n966);
assign n490 = ~n5531;
assign n999 = n9750 | n4371;
assign n5811 = ~(n7893 | n291);
assign n4271 = ~(n3168 | n10348);
assign n12068 = n636 | n12735;
assign n2076 = ~n12706;
assign n10627 = ~(n9510 ^ n851);
assign n8741 = ~(n5885 ^ n10164);
assign n6963 = n9723 | n12736;
assign n5770 = n10925 | n11911;
assign n2237 = ~(n6664 ^ n8627);
assign n7708 = ~n10979;
assign n8228 = n6073 & n8947;
assign n8420 = ~(n6208 ^ n6269);
assign n1335 = ~n12713;
assign n6572 = ~(n1342 | n7497);
assign n12308 = ~(n5629 ^ n8716);
assign n3369 = n12792 & n2220;
assign n3113 = ~(n9048 ^ n5993);
assign n5819 = ~(n10889 ^ n7455);
assign n5150 = ~(n7321 ^ n2104);
assign n6886 = n9202 & n7379;
assign n6118 = ~(n10013 ^ n9298);
assign n171 = ~n8009;
assign n10492 = n638 & n7227;
assign n9668 = ~(n2213 ^ n1443);
assign n10042 = n7236 & n11876;
assign n12212 = n1392 & n2337;
assign n3581 = n11073 | n5965;
assign n6875 = n246 & n5633;
assign n12285 = ~(n1762 | n5238);
assign n2936 = n8903 | n5834;
assign n8724 = ~(n11543 ^ n924);
assign n11838 = n989 | n1546;
assign n4629 = ~(n11708 ^ n11243);
assign n4319 = n7130 | n2371;
assign n8111 = n12237 | n12535;
assign n6562 = ~(n11596 ^ n5864);
assign n2487 = n1989 & n3600;
assign n6692 = ~(n10970 ^ n11448);
assign n3458 = ~(n2834 ^ n2017);
assign n10494 = ~(n638 ^ n1446);
assign n2545 = ~(n9828 ^ n952);
assign n9965 = ~(n5371 ^ n1780);
assign n8178 = ~(n5532 | n2604);
assign n11147 = n11923 | n4527;
assign n1622 = ~(n4430 ^ n2054);
assign n1082 = n11026 | n10916;
assign n8348 = n2099 | n1163;
assign n8486 = n3207 & n10957;
assign n1757 = n7749 | n8602;
assign n10124 = n4250 | n7101;
assign n2478 = ~(n3943 | n7708);
assign n1228 = ~(n9428 ^ n9981);
assign n4157 = ~(n8423 ^ n7315);
assign n8463 = ~(n3767 ^ n8601);
assign n9317 = ~(n2340 ^ n6152);
assign n8303 = n5732 ^ n5336;
assign n10085 = n9122 & n4460;
assign n8631 = n242 | n12250;
assign n10958 = ~(n3380 | n4252);
assign n1579 = n1699 | n6071;
assign n5316 = n4358 & n10165;
assign n10473 = ~(n9382 ^ n3001);
assign n2321 = n8428 | n2815;
assign n4965 = n9271 & n1866;
assign n3103 = n7916 & n2642;
assign n8152 = ~n5213;
assign n3034 = ~(n8018 ^ n744);
assign n10839 = n9370 | n12328;
assign n10454 = ~(n1661 ^ n6545);
assign n10310 = n4175 | n457;
assign n6142 = n1653 | n10896;
assign n4910 = ~(n6400 ^ n2360);
assign n8690 = ~n7121;
assign n10461 = n6718 | n12120;
assign n11803 = ~n6866;
assign n372 = n5350 & n3540;
assign n9377 = ~n6787;
assign n4958 = n9561 | n11702;
assign n6911 = n1937 | n12816;
assign n8730 = n6510 | n49;
assign n2061 = ~(n5956 ^ n2369);
assign n11117 = ~(n1930 ^ n9047);
assign n2307 = n3655 & n4653;
assign n12594 = ~(n7659 | n9923);
assign n8651 = ~(n6335 ^ n5728);
assign n7187 = n8623 & n7113;
assign n2050 = ~n8938;
assign n3442 = n3127 | n10419;
assign n5257 = ~(n10357 ^ n5568);
assign n5834 = n5489 & n10173;
assign n2462 = ~(n4717 ^ n12433);
assign n7483 = ~(n3418 ^ n2490);
assign n7076 = n3218 | n3846;
assign n4520 = ~(n1033 ^ n617);
assign n5455 = ~n11016;
assign n9277 = n12138 | n7132;
assign n12377 = ~(n11098 | n2315);
assign n11028 = ~(n1179 | n7664);
assign n1103 = ~(n12125 ^ n1204);
assign n12342 = n11892 & n217;
assign n6480 = ~(n2246 ^ n9569);
assign n9422 = ~n8937;
assign n4639 = ~(n3509 | n727);
assign n221 = ~(n5107 | n258);
assign n9126 = n2956 | n6653;
assign n11397 = ~(n842 ^ n10764);
assign n1049 = n12442 | n10382;
assign n3740 = ~n6165;
assign n1169 = n4760 & n10105;
assign n12150 = n8181 & n8485;
assign n4048 = ~n11265;
assign n2984 = n10904 | n126;
assign n8290 = n1183 | n10854;
assign n8158 = ~n5745;
assign n6389 = ~n2879;
assign n7837 = n295 | n8415;
assign n9153 = ~(n9388 ^ n6619);
assign n5683 = ~n4809;
assign n3724 = n12398 | n4655;
assign n1355 = n9512 & n5173;
assign n8260 = n3127 | n8524;
assign n12831 = n2099 | n12441;
assign n8029 = ~(n6075 ^ n12581);
assign n7347 = n2671 | n9678;
assign n8443 = ~(n4210 | n5871);
assign n8006 = n1146 | n8593;
assign n12126 = ~(n7468 ^ n271);
assign n7882 = ~(n8058 ^ n6323);
assign n4258 = ~(n8581 ^ n4231);
assign n8100 = ~(n750 ^ n863);
assign n2201 = n6577 | n8414;
assign n1179 = ~n7009;
assign n9690 = n8042 | n1905;
assign n9775 = n7843 & n3005;
assign n8929 = ~n2945;
assign n8182 = ~(n2474 | n6830);
assign n1955 = n4456 | n10442;
assign n11129 = n5659 | n366;
assign n7119 = n12862 & n5595;
assign n661 = n6349 | n8350;
assign n3565 = n4744 & n171;
assign n3098 = ~n9572;
assign n7791 = n11923 | n9078;
assign n8763 = n11892 & n2749;
assign n9184 = ~(n9621 ^ n1490);
assign n1142 = ~(n2600 | n12332);
assign n10231 = n9878 | n10854;
assign n6119 = n7046 & n11778;
assign n3993 = n1998 & n6081;
assign n9684 = ~(n10144 ^ n10484);
assign n7261 = n10546 | n1307;
assign n5800 = n3757 | n10363;
assign n12481 = n5559 & n496;
assign n2007 = ~(n2086 ^ n7547);
assign n6659 = ~(n7359 ^ n8616);
assign n11289 = n4498 | n5497;
assign n10195 = ~(n2608 | n4615);
assign n1467 = ~n670;
assign n12265 = ~(n11377 ^ n4052);
assign n9114 = n3096 | n6197;
assign n12106 = ~(n887 ^ n8942);
assign n12785 = ~(n9065 ^ n141);
assign n11886 = ~(n4999 ^ n4897);
assign n2345 = ~(n3978 ^ n3515);
assign n11694 = n7391 | n1851;
assign n1064 = n118 & n5957;
assign n11474 = ~n7519;
assign n6846 = n2125 & n9796;
assign n12160 = ~(n5177 ^ n4626);
assign n9081 = n11026 | n9568;
assign n9402 = ~n5697;
assign n5261 = ~n9539;
assign n4451 = n1941 | n11820;
assign n12075 = ~(n747 ^ n4069);
assign n1443 = n5436 & n6471;
assign n676 = ~n9677;
assign n7897 = n12406 & n5121;
assign n9592 = n6030 & n3866;
assign n6858 = ~(n5377 ^ n10765);
assign n1968 = ~(n1557 | n7030);
assign n10924 = ~(n176 ^ n6873);
assign n10008 = ~(n1689 ^ n9950);
assign n1682 = n7449 | n6922;
assign n4784 = n9978 | n2489;
assign n2632 = n3992 & n8433;
assign n5703 = n8535 | n2410;
assign n9494 = ~(n4980 | n8875);
assign n9082 = n7391 | n7881;
assign n4696 = n7116 | n12816;
assign n7725 = ~n716;
assign n11913 = n1161 & n134;
assign n12192 = n11434 | n10153;
assign n3185 = ~(n12347 | n9480);
assign n1397 = n10545 & n7159;
assign n3564 = ~(n10959 ^ n3879);
assign n8596 = n10142 | n2076;
assign n500 = n10657 | n11861;
assign n9942 = n7363 & n10684;
assign n3555 = n9004 | n3164;
assign n8213 = ~(n10527 ^ n4227);
assign n2670 = n994 | n1162;
assign n1528 = ~(n1139 ^ n5098);
assign n5190 = n11969 & n5585;
assign n5526 = n12391 & n2558;
assign n6193 = ~n1185;
assign n12583 = n5395 & n1952;
assign n10722 = ~(n8066 ^ n9294);
assign n8639 = ~(n4777 ^ n7475);
assign n10497 = ~(n6177 ^ n10713);
assign n141 = ~(n9073 ^ n4641);
assign n7553 = ~n270;
assign n3900 = n3562 | n10796;
assign n7127 = n6601 & n7223;
assign n5167 = n11736 & n569;
assign n7230 = n12675 & n11381;
assign n10258 = n11204 & n243;
assign n6464 = ~(n12351 ^ n5804);
assign n4032 = n3967 | n8057;
assign n6740 = n3746 | n11820;
assign n9773 = n4966 & n5161;
assign n442 = ~(n690 | n11084);
assign n1693 = ~(n12004 ^ n5033);
assign n9719 = ~(n4012 ^ n1971);
assign n5673 = n9199 & n2302;
assign n2623 = ~(n8863 ^ n7766);
assign n839 = n6590 | n11930;
assign n11893 = ~n9547;
assign n7577 = n4787 & n1889;
assign n3734 = n7810 | n4538;
assign n9652 = n6718 | n9144;
assign n9954 = n2995 & n10800;
assign n1130 = ~n1584;
assign n6681 = n5530 | n5326;
assign n7139 = n12803 & n11117;
assign n12032 = ~(n11324 ^ n12756);
assign n639 = ~(n2381 ^ n8506);
assign n1461 = n2456 | n6071;
assign n3623 = n10435 & n4895;
assign n11001 = ~(n8123 ^ n6774);
assign n10036 = ~(n9152 ^ n9509);
assign n5449 = n7906 | n9794;
assign n2236 = n12930 | n6947;
assign n886 = ~(n2837 | n5360);
assign n8020 = n4960 | n4945;
assign n5473 = n9373 | n12771;
assign n1311 = ~n1594;
assign n186 = n12705 & n3932;
assign n10142 = ~n6687;
assign n9203 = n11923 | n2020;
assign n9070 = n2056 | n10008;
assign n10747 = ~(n5294 ^ n4748);
assign n2654 = n4579 | n1167;
assign n11602 = n8216 | n10480;
assign n9159 = n5160 | n9283;
assign n1496 = ~(n6993 ^ n8633);
assign n5652 = n4628 | n530;
assign n1005 = ~(n11813 | n8922);
assign n64 = n2842 & n6424;
assign n10675 = n6032 | n3801;
assign n8405 = ~n6578;
assign n11788 = ~(n11610 ^ n2547);
assign n4774 = n4972 & n2542;
assign n11068 = n5945 | n2232;
assign n8169 = n2382 | n948;
assign n4396 = ~(n5092 | n3074);
assign n1714 = n12610 | n7794;
assign n11266 = n11923 | n4875;
assign n11608 = n3127 | n11827;
assign n8210 = ~n8772;
assign n9482 = n12273 & n9256;
assign n6458 = n5788 | n7673;
assign n7728 = ~(n2009 ^ n12921);
assign n5978 = n4481 & n10634;
assign n4176 = ~n6751;
assign n6028 = n11941 | n4793;
assign n12190 = ~(n9490 | n767);
assign n1730 = ~(n5559 | n496);
assign n11371 = ~(n6067 | n8182);
assign n1151 = n4275 & n9813;
assign n7449 = ~n7388;
assign n3704 = ~(n6984 ^ n2543);
assign n1366 = ~(n4714 ^ n1118);
assign n5735 = ~n10425;
assign n8668 = ~(n10743 ^ n8721);
assign n8135 = n288 | n11386;
assign n10134 = n3829 | n10384;
assign n12158 = ~(n1091 ^ n10497);
assign n7652 = ~(n4794 ^ n7799);
assign n3389 = n4247 | n554;
assign n4228 = n10196 | n8643;
assign n1547 = n10824 | n6501;
assign n2262 = ~n10831;
assign n2825 = ~(n5454 ^ n9125);
assign n1686 = n1261 & n2366;
assign n12867 = n7683 & n12954;
assign n10831 = n2093 | n6102;
assign n3359 = n9829 & n5541;
assign n4421 = ~n5207;
assign n11610 = ~(n5784 ^ n10591);
assign n9902 = ~(n8484 ^ n4363);
assign n5983 = ~(n11624 ^ n3484);
assign n2045 = n8428 | n6197;
assign n5276 = n3627 & n6038;
assign n8357 = ~(n6135 ^ n12459);
assign n4122 = ~(n12931 | n9495);
assign n8649 = n27 | n1050;
assign n8783 = ~(n6467 ^ n11860);
assign n3278 = n11923 | n4864;
assign n7199 = ~(n4512 | n11170);
assign n10118 = n5765 | n9144;
assign n2353 = ~(n2549 | n1680);
assign n2093 = ~(n7115 | n310);
assign n5045 = ~n7464;
assign n8328 = ~(n5647 | n10263);
assign n2589 = ~n2278;
assign n4046 = n6072 | n891;
assign n12401 = n3251 & n1274;
assign n3705 = ~(n2906 ^ n6699);
assign n1292 = n12722 | n1763;
assign n12759 = n3491 & n8543;
assign n12122 = n2099 | n9188;
assign n10981 = ~(n5109 ^ n12295);
assign n2187 = n8229 | n1276;
assign n416 = ~(n7504 ^ n224);
assign n12307 = ~n12664;
assign n2949 = ~(n1760 ^ n12766);
assign n7022 = ~n4386;
assign n8096 = n11552 | n8830;
assign n2795 = n9379 & n1356;
assign n2663 = n7116 | n8768;
assign n9745 = ~(n2314 ^ n268);
assign n2765 = ~(n2644 ^ n12810);
assign n6843 = n7283 | n9589;
assign n1239 = n7243 | n2460;
assign n6803 = ~(n8118 ^ n11933);
assign n10530 = n8583 | n9144;
assign n1494 = n4347 & n6375;
assign n1602 = n4369 & n467;
assign n8141 = ~(n4717 | n12302);
assign n2705 = n11328 & n6043;
assign n11482 = ~(n7551 ^ n9867);
assign n5091 = ~(n8163 | n3914);
assign n12323 = ~(n11550 ^ n5176);
assign n6479 = ~(n1654 ^ n8571);
assign n2455 = n6574 | n8331;
assign n7550 = n10843 | n11295;
assign n2352 = ~(n11617 ^ n8400);
assign n8505 = ~n2500;
assign n2119 = ~(n10456 ^ n32);
assign n3216 = ~n9437;
assign n2113 = n4059 | n561;
assign n307 = n4492 | n11901;
assign n11355 = n9905 & n10792;
assign n10096 = n2687 & n7153;
assign n10752 = n2159 & n12822;
assign n12184 = ~(n1637 | n11325);
assign n163 = ~(n10497 | n1091);
assign n1819 = ~(n7763 ^ n185);
assign n2988 = n12727 | n8005;
assign n6836 = n2217 | n1476;
assign n12416 = n12853 | n8109;
assign n7622 = ~(n4137 ^ n4640);
assign n11950 = n12699 & n4113;
assign n10182 = n7116 | n11122;
assign n4842 = n9136 | n7642;
assign n3749 = ~(n2674 ^ n11847);
assign n4558 = ~(n3769 ^ n3070);
assign n7215 = ~(n5887 ^ n11904);
assign n11812 = ~n255;
assign n3757 = n5765 | n1047;
assign n11320 = ~(n9000 ^ n11598);
assign n12746 = n5355 | n4400;
assign n9672 = ~(n11646 ^ n1203);
assign n826 = ~n5645;
assign n2185 = ~(n10639 | n6479);
assign n9950 = ~n4967;
assign n42 = ~(n12508 ^ n2994);
assign n409 = ~(n715 ^ n4000);
assign n6489 = n1985 & n4186;
assign n7796 = ~(n2307 ^ n12902);
assign n12480 = ~(n3541 ^ n11067);
assign n11720 = ~(n817 ^ n9361);
assign n6409 = n6642 & n1893;
assign n7063 = ~n10556;
assign n10319 = ~(n6580 ^ n5304);
assign n11105 = ~(n11280 ^ n8825);
assign n2679 = ~(n68 ^ n1876);
assign n8406 = ~(n11983 ^ n1036);
assign n4978 = ~(n4669 ^ n9650);
assign n2004 = ~(n3148 ^ n6821);
assign n7775 = ~(n5983 ^ n9347);
assign n260 = n10208 | n11932;
assign n1400 = ~(n7686 ^ n10079);
assign n10621 = n41 & n1255;
assign n10953 = n9529 & n7950;
assign n8567 = ~(n2432 ^ n213);
assign n9812 = n5108 & n9198;
assign n878 = n756 | n12428;
assign n3433 = ~n4270;
assign n12098 = n6373 | n4875;
assign n12419 = n6001 | n1152;
assign n584 = n4994 | n2980;
assign n534 = ~(n6889 ^ n6179);
assign n8356 = n3627 & n11407;
assign n4467 = ~(n7684 | n12162);
assign n7743 = ~(n2717 ^ n5282);
assign n8151 = ~(n8055 ^ n8344);
assign n727 = ~n7528;
assign n724 = n3275 | n9293;
assign n9475 = n8753 & n5752;
assign n3448 = ~(n3068 ^ n12058);
assign n7346 = n4716 & n7;
assign n1120 = ~(n633 ^ n1221);
assign n1220 = n5960 & n10664;
assign n12316 = n994 | n9589;
assign n5113 = ~(n9903 ^ n7362);
assign n5603 = ~(n6964 ^ n2143);
assign n11455 = n5589 & n11291;
assign n906 = n4453 | n4706;
assign n9658 = n11535 & n11767;
assign n4061 = n10750 | n6071;
assign n8378 = ~(n9863 ^ n12860);
assign n7033 = n921 | n8298;
assign n6069 = n2838 & n6164;
assign n1019 = n9389 | n11746;
assign n3815 = n10640 & n5223;
assign n7778 = n6358 & n217;
assign n545 = n333 | n487;
assign n8987 = n8490 & n5321;
assign n7813 = n8945 & n1859;
assign n3337 = n8158 & n5616;
assign n11399 = ~(n6515 ^ n11471);
assign n4013 = n2045 | n11274;
assign n3333 = n0 & n9322;
assign n7378 = n4911 | n1455;
assign n425 = ~(n75 ^ n1823);
assign n8933 = n8363 & n5806;
assign n8407 = ~n2695;
assign n8451 = n12924 | n1124;
assign n4891 = n10843 & n11295;
assign n11833 = ~(n408 ^ n11082);
assign n813 = n7306 & n10584;
assign n10366 = ~(n2457 ^ n2517);
assign n2667 = n2266 | n11618;
assign n5722 = ~(n11021 ^ n9660);
assign n6945 = n8583 | n8830;
assign n2085 = n12299 & n8819;
assign n3413 = ~(n9709 | n2015);
assign n10485 = n11108 | n11637;
assign n779 = n10642 | n9973;
assign n12774 = ~(n11137 | n470);
assign n10176 = n8758 & n12630;
assign n523 = n2367 | n4474;
assign n2252 = ~n8447;
assign n3269 = ~(n12210 ^ n12536);
assign n9535 = ~(n1062 ^ n12811);
assign n11902 = n5466 | n4578;
assign n5663 = n1808 | n2210;
assign n11496 = ~(n4742 ^ n8621);
assign n6113 = ~(n9298 | n10013);
assign n9436 = ~(n6161 ^ n12599);
assign n938 = n10354 | n1502;
assign n6696 = ~n9391;
assign n4526 = ~(n9493 ^ n10069);
assign n428 = n4121 | n11975;
assign n6093 = n2013 | n8542;
assign n4749 = ~(n9079 ^ n6695);
assign n7024 = ~(n1242 ^ n6378);
assign n12728 = ~(n3225 ^ n7099);
assign n2814 = n11358 | n6201;
assign n7169 = n11416 | n2535;
assign n9803 = n11832 & n9681;
assign n12148 = ~(n4703 ^ n11570);
assign n9925 = n9802 | n9220;
assign n12850 = ~(n9368 ^ n809);
assign n2695 = n12503 | n2020;
assign n10909 = ~(n7441 | n3009);
assign n8765 = ~(n11563 ^ n5192);
assign n8034 = ~(n7579 | n10073);
assign n3538 = ~n733;
assign n3101 = ~(n5016 ^ n12202);
assign n3434 = ~n3443;
assign n4231 = ~(n771 ^ n1829);
assign n12242 = n10835 | n9160;
assign n3793 = n3837 | n9096;
assign n9797 = n10835 | n10916;
assign n4610 = ~n4784;
assign n8264 = n5847 | n136;
assign n6933 = ~(n645 | n4043);
assign n1184 = ~n6474;
assign n6893 = n10874 | n1300;
assign n2764 = ~(n11538 ^ n8798);
assign n12610 = ~(n12118 ^ n3721);
assign n2369 = ~(n522 ^ n8401);
assign n3050 = n10835 | n1047;
assign n9670 = n5384 & n12652;
assign n5592 = n8115 | n1106;
assign n2351 = n8467 | n8231;
assign n7266 = n11271 | n8239;
assign n9060 = n9119 & n1182;
assign n1542 = n10326 & n9618;
assign n10619 = n11719 | n10066;
assign n5902 = ~n6826;
assign n9345 = n9236 & n1559;
assign n1538 = ~(n11605 ^ n3278);
assign n9235 = ~n3460;
assign n1976 = ~(n10746 | n10577);
assign n11124 = n3381 & n10811;
assign n5218 = ~(n11548 | n4523);
assign n11467 = ~(n6907 ^ n3610);
assign n8434 = ~(n3840 ^ n4151);
assign n4333 = ~(n8792 ^ n6372);
assign n9794 = n9878 | n12535;
assign n8962 = ~n8732;
assign n2012 = ~n8790;
assign n3522 = ~n1027;
assign n1661 = ~(n2063 ^ n7466);
assign n1445 = n8959 | n6197;
assign n10573 = n12237 | n3224;
assign n5617 = ~(n12195 ^ n4622);
assign n10225 = n10336 & n11677;
assign n11469 = ~(n1248 ^ n8440);
assign n11350 = ~n10914;
assign n10641 = ~n9738;
assign n6556 = ~(n3085 ^ n2554);
assign n947 = n8152 | n11942;
assign n9432 = n5355 | n7703;
assign n1168 = ~(n6413 ^ n12778);
assign n8107 = ~(n9358 ^ n547);
assign n8956 = ~(n7092 ^ n4030);
assign n1871 = ~n3978;
assign n10673 = n5384 | n12652;
assign n2221 = ~n1611;
assign n837 = ~(n5483 ^ n5072);
assign n1043 = n6577 | n9741;
assign n7768 = n2097 | n3792;
assign n1406 = ~(n6889 | n9422);
assign n12290 = n9368 & n809;
assign n12928 = ~(n11234 ^ n2359);
assign n4284 = ~(n2069 ^ n10458);
assign n5851 = ~n3865;
assign n5772 = ~(n8287 ^ n10188);
assign n2600 = n12119 | n12446;
assign n9689 = ~(n7070 | n10571);
assign n3765 = n9933 & n8729;
assign n8705 = n3771 & n3302;
assign n11299 = n2497 | n9001;
assign n566 = n6934 & n1377;
assign n6799 = ~(n4926 ^ n2745);
assign n1038 = ~(n7285 ^ n6498);
assign n11093 = n3766 & n11974;
assign n1917 = n849 | n4575;
assign n3814 = n3581 & n6230;
assign n2441 = n3236 & n3067;
assign n7696 = ~(n3517 ^ n823);
assign n3751 = ~(n1252 | n9565);
assign n8854 = n196 & n11477;
assign n5829 = ~(n6794 | n3545);
assign n3652 = n6550 | n5792;
assign n10418 = n8071 | n7595;
assign n8137 = n5850 | n1347;
assign n4264 = n6977 | n5012;
assign n11031 = ~n11501;
assign n3405 = n1051 | n12816;
assign n11775 = ~n3602;
assign n5594 = ~n6087;
assign n1520 = ~(n11112 ^ n5123);
assign n12843 = ~n4921;
assign n7279 = ~(n9194 ^ n2480);
assign n1911 = n7735 & n1324;
assign n4801 = ~(n7817 | n9118);
assign n7096 = n10742 & n12001;
assign n10101 = ~n1515;
assign n3739 = n6766 | n395;
assign n3214 = ~(n4583 ^ n4276);
assign n7326 = ~n12710;
assign n3301 = ~(n7746 ^ n4743);
assign n1317 = n2217 | n9160;
assign n270 = n12531 | n5565;
assign n2395 = n5915 | n3224;
assign n3166 = n10142 | n4400;
assign n5192 = n7449 | n9521;
assign n6287 = n9570 & n12050;
assign n4849 = n4059 | n1455;
assign n11369 = ~n12632;
assign n6942 = ~(n3985 ^ n5112);
assign n4369 = n10551 | n7988;
assign n8282 = n6977 | n8414;
assign n8459 = n9896 & n9815;
assign n3151 = ~(n11343 ^ n6106);
assign n10632 = n9262 | n4474;
assign n6602 = ~(n10525 | n9466);
assign n8684 = ~n7143;
assign n9783 = ~(n12142 ^ n12061);
assign n11232 = n3746 | n7395;
assign n6985 = ~n4079;
assign n10472 = n4202 & n9496;
assign n11794 = n3324 | n1509;
assign n1348 = ~(n9063 | n9580);
assign n1201 = ~(n3584 ^ n4037);
assign n5606 = n11950 & n5127;
assign n3465 = n4187 & n3602;
assign n2277 = ~(n221 | n3529);
assign n1448 = ~n10904;
assign n12409 = ~(n2912 ^ n4192);
assign n9882 = n11152 & n10482;
assign n469 = ~(n6220 ^ n59);
assign n12589 = ~(n10983 ^ n91);
assign n11505 = n10108 | n11827;
assign n12407 = ~(n5424 | n9337);
assign n9433 = n7221 | n6453;
assign n10312 = n2593 | n8497;
assign n12268 = ~(n7386 ^ n8651);
assign n8606 = ~(n3077 ^ n2627);
assign n3272 = ~(n5354 ^ n6014);
assign n10562 = ~(n1785 ^ n12143);
assign n2387 = ~(n2637 ^ n8950);
assign n4771 = ~(n6090 ^ n1698);
assign n2982 = n5089 | n10823;
assign n3589 = n7905 | n12431;
assign n10384 = ~(n721 | n9327);
assign n12094 = ~(n7483 ^ n5297);
assign n10980 = ~(n4541 | n7995);
assign n10128 = n3324 | n4474;
assign n3541 = n10508 | n10930;
assign n10636 = n10199 | n7637;
assign n6597 = ~(n9446 | n9051);
assign n11384 = n1705 | n12251;
assign n11501 = n12815 & n10109;
assign n6127 = ~(n10744 ^ n5913);
assign n9874 = ~(n9145 ^ n12649);
assign n4887 = ~(n9499 ^ n11096);
assign n4414 = n12069 & n1564;
assign n4668 = n3265 & n1454;
assign n323 = n12879 & n7792;
assign n7512 = ~n2640;
assign n9278 = ~(n2011 | n4899);
assign n10087 = n6087 ^ n3134;
assign n5106 = ~(n6168 ^ n4418);
assign n10741 = n5289 & n6166;
assign n12363 = ~n11842;
assign n9112 = n4013 & n9800;
assign n382 = ~(n8140 ^ n10253);
assign n11508 = n6776 & n6703;
assign n3426 = n3693 | n12795;
assign n9989 = ~(n4930 | n12448);
assign n5098 = ~n6683;
assign n10704 = ~(n9278 | n12352);
assign n10681 = ~(n10815 ^ n9254);
assign n5217 = ~(n7244 ^ n2890);
assign n5541 = ~n11256;
assign n7287 = n11425 | n6025;
assign n11768 = ~(n5846 ^ n12628);
assign n9796 = n12283 | n8333;
assign n691 = ~(n7496 ^ n3436);
assign n10843 = ~(n11533 ^ n12068);
assign n3367 = ~(n2488 ^ n6203);
assign n9806 = n5809 | n12080;
assign n8191 = n7283 | n2076;
assign n4803 = n5231 & n5217;
assign n12449 = ~(n8313 ^ n879);
assign n4238 = n10735 | n4091;
assign n3285 = ~(n3884 ^ n734);
assign n8084 = ~(n12203 ^ n10593);
assign n4034 = n3274 & n3755;
assign n350 = ~(n1065 | n4039);
assign n8900 = n7236 & n5760;
assign n8782 = n7271 | n11263;
assign n2639 = ~(n10918 | n12900);
assign n1561 = n5020 & n3916;
assign n5721 = ~(n12873 ^ n10513);
assign n6384 = n8176 & n2388;
assign n8789 = n5575 | n11896;
assign n7437 = n4428 | n8797;
assign n1745 = n1507 | n9168;
assign n134 = n10521 | n1828;
assign n699 = n8903 & n5834;
assign n10822 = n3666 | n7068;
assign n12100 = ~(n10091 ^ n3560);
assign n12091 = ~(n6195 ^ n7571);
assign n1551 = ~(n5284 ^ n12676);
assign n12443 = n994 | n1079;
assign n4052 = ~n10042;
assign n2188 = n9797 | n2900;
assign n8293 = ~n10741;
assign n1361 = ~(n8027 ^ n228);
assign n5325 = ~(n1408 ^ n11875);
assign n7395 = ~n10278;
assign n10075 = n11462 | n11148;
assign n976 = n2651 | n4394;
assign n9636 = ~n10080;
assign n3536 = ~(n11568 ^ n8846);
assign n3729 = n3746 | n10919;
assign n4453 = ~(n6485 | n1187);
assign n368 = ~(n1571 ^ n9891);
assign n10633 = n4522 | n4656;
assign n10774 = n5204 | n283;
assign n7705 = ~n5432;
assign n7653 = ~(n5795 ^ n6118);
assign n7846 = n7283 | n1738;
assign n5846 = ~(n10393 ^ n2540);
assign n5932 = ~(n1989 | n3600);
assign n10024 = ~(n10457 ^ n7820);
assign n893 = n5026 & n9139;
assign n4466 = n8941 | n1418;
assign n7776 = n12658 & n6327;
assign n1931 = ~n7312;
assign n4811 = ~n10517;
assign n3546 = ~(n11267 ^ n4751);
assign n4952 = ~n6203;
assign n11358 = n7168 | n3047;
assign n10742 = n9920 & n4921;
assign n2145 = n991 & n354;
assign n5376 = n1215 & n5055;
assign n8744 = ~(n7146 ^ n9552);
assign n11377 = ~n2824;
assign n4841 = ~n8773;
assign n9471 = ~(n2739 | n1033);
assign n5651 = ~(n6857 ^ n4544);
assign n3017 = n11892 & n11791;
assign n9534 = ~n11468;
assign n11200 = n10332 | n12934;
assign n6539 = n3746 | n11122;
assign n11394 = n5493 | n5019;
assign n2849 = ~n4;
assign n7674 = n9075 | n4840;
assign n512 = ~(n4233 ^ n11553);
assign n7820 = n7453 & n2059;
assign n7040 = ~(n3651 | n3183);
assign n8535 = ~(n4655 ^ n4825);
assign n8528 = n2427 & n1157;
assign n7636 = ~(n1050 ^ n2544);
assign n10907 = ~(n10297 ^ n2983);
assign n3618 = n12474 | n881;
assign n5317 = ~(n7844 ^ n12378);
assign n6499 = ~(n5501 ^ n4792);
assign n6588 = ~(n5848 ^ n3913);
assign n4864 = ~n1510;
assign n454 = ~(n10904 ^ n5789);
assign n8255 = n817 | n9817;
assign n6110 = ~(n12867 ^ n3443);
assign n4128 = ~(n8189 ^ n5797);
assign n1750 = ~(n11564 ^ n5015);
assign n2388 = ~(n5009 ^ n821);
assign n4105 = n3992 & n8028;
assign n8172 = ~(n2272 ^ n10258);
assign n6332 = ~(n2625 | n4874);
assign n5522 = n11887 | n9188;
assign n5625 = n4780 | n10436;
assign n2227 = n12680 & n3783;
assign n3758 = ~(n775 ^ n11071);
assign n516 = ~(n11417 ^ n1314);
assign n195 = ~(n9999 ^ n7478);
assign n4998 = ~(n5942 ^ n11064);
assign n6444 = n3964 & n1334;
assign n80 = n6801 & n6011;
assign n11212 = n4628 | n5781;
assign n3944 = n1699 | n1932;
assign n9192 = n213 | n2432;
assign n8540 = n11422 & n10028;
assign n3019 = ~(n10441 ^ n12904);
assign n10424 = n2901 & n2938;
assign n4689 = ~(n595 ^ n10785);
assign n2590 = n12723 & n1130;
assign n4678 = ~(n669 ^ n10559);
assign n5457 = n7284 & n10144;
assign n7803 = ~n12162;
assign n11708 = ~(n3592 ^ n12383);
assign n1001 = ~(n2979 ^ n9476);
assign n8296 = ~(n7608 ^ n10632);
assign n6633 = ~(n3600 ^ n8107);
assign n10263 = ~(n610 | n469);
assign n6176 = ~(n6098 ^ n1845);
assign n5840 = ~n6824;
assign n7358 = ~n10947;
assign n9595 = ~(n4886 ^ n5135);
assign n7150 = ~(n12875 | n6875);
assign n8060 = ~(n11036 ^ n5252);
assign n12612 = ~(n9244 | n4025);
assign n11850 = n6738 | n11179;
assign n2738 = n11259 & n6119;
assign n5561 = n4184 & n3169;
assign n5704 = ~n5236;
assign n11412 = ~(n6945 ^ n7023);
assign n5016 = n8026 | n10903;
assign n10730 = n7839 | n2815;
assign n4524 = ~(n1366 ^ n8351);
assign n3303 = n7161 | n8765;
assign n10888 = ~(n901 | n11252);
assign n4459 = n11593 | n4584;
assign n2659 = n5915 | n826;
assign n9889 = n2832 | n6389;
assign n12810 = ~(n4413 ^ n10803);
assign n10254 = ~(n9649 ^ n12726);
assign n8804 = ~(n2611 ^ n286);
assign n5956 = ~(n3523 ^ n9682);
assign n9228 = n1051 | n2815;
assign n9858 = n4828 & n2498;
assign n3064 = n12299 & n2522;
assign n12737 = n7668 & n9130;
assign n1342 = n5765 | n8285;
assign n367 = n9795 | n9719;
assign n3320 = ~(n8092 ^ n8358);
assign n2409 = n6590 & n11930;
assign n9914 = ~(n12294 | n6665);
assign n586 = n10838 | n3060;
assign n8757 = n10157 | n3606;
assign n5970 = ~n5192;
assign n10658 = ~(n8790 ^ n4089);
assign n1857 = ~n1949;
assign n8108 = n6931 | n4506;
assign n9638 = n11028 | n8;
assign n7632 = ~(n2874 ^ n9587);
assign n5774 = n222 & n9742;
assign n1286 = ~n12159;
assign n10462 = n6373 | n609;
assign n7428 = ~(n7794 ^ n11888);
assign n2916 = n8011 & n4866;
assign n6285 = ~(n2629 ^ n8062);
assign n2417 = ~n7043;
assign n4848 = ~n11878;
assign n1672 = ~(n8712 ^ n10344);
assign n809 = n5765 | n9160;
assign n92 = n7407 | n10662;
assign n12034 = ~n6520;
assign n6760 = ~(n10580 ^ n9095);
assign n11182 = n8428 | n7425;
assign n9972 = n8428 | n8414;
assign n12682 = ~(n11694 ^ n4377);
assign n5165 = ~(n12772 ^ n9264);
assign n6974 = n7826 & n12034;
assign n10306 = n12797 | n7876;
assign n268 = ~(n3006 ^ n2446);
assign n2620 = ~n5327;
assign n5346 = n8844 & n302;
assign n3457 = n7449 | n4654;
assign n1360 = n9331 | n1592;
assign n5715 = ~n7024;
assign n4416 = ~(n11995 ^ n8168);
assign n9497 = n8738 | n12771;
assign n12849 = n12260 | n1501;
assign n5214 = n4059 | n7881;
assign n9545 = ~(n9749 ^ n7513);
assign n6817 = n4498 | n1915;
assign n2945 = n12237 | n8109;
assign n9619 = n12731 & n2110;
assign n8610 = n4815 | n5729;
assign n1281 = ~(n12736 ^ n2764);
assign n3885 = n1051 | n10903;
assign n4730 = ~(n3704 ^ n9396);
assign n5513 = ~(n11259 ^ n6119);
assign n2092 = ~(n4469 ^ n1428);
assign n8119 = n5809 | n5326;
assign n5026 = ~(n11750 ^ n10935);
assign n2909 = ~(n12911 ^ n2198);
assign n11734 = n7082 & n10579;
assign n5215 = n1675 | n344;
assign n6684 = n3241 | n6236;
assign n9234 = ~(n5542 ^ n11232);
assign n3 = ~(n1451 ^ n9676);
assign n6668 = ~(n7035 ^ n11168);
assign n7975 = ~(n12490 ^ n6916);
assign n9573 = n11172 | n6019;
assign n10643 = n3746 | n6169;
assign n7623 = ~(n7526 ^ n4988);
assign n6166 = n7001 | n6401;
assign n3295 = n10565 | n10570;
assign n10926 = n4059 | n1851;
assign n138 = n6589 & n4049;
assign n6601 = n9108 | n3983;
assign n2882 = ~(n5931 ^ n4617);
assign n8319 = n7832 & n11869;
assign n4897 = n4201 & n11762;
assign n4731 = n113 | n10259;
assign n9602 = ~(n6368 ^ n12416);
assign n1270 = n2367 | n2020;
assign n7282 = n5064 | n8974;
assign n9448 = ~n7779;
assign n216 = ~(n8035 ^ n6322);
assign n5068 = ~n12319;
assign n4170 = ~(n9794 ^ n4954);
assign n10017 = n4531 & n4885;
assign n1394 = ~n6904;
assign n3738 = ~(n459 ^ n8609);
assign n3327 = n8555 & n11568;
assign n11771 = ~(n4366 ^ n10752);
assign n7677 = ~(n10160 ^ n12201);
assign n5913 = n2289 & n12192;
assign n5697 = n9472 & n9462;
assign n6307 = ~n1706;
assign n761 = ~(n6244 ^ n4042);
assign n1245 = ~(n11246 ^ n7814);
assign n9154 = ~(n808 ^ n5849);
assign n6011 = n8026 | n10919;
assign n12241 = n8759 & n3719;
assign n11428 = ~n11882;
assign n11465 = n3455 & n5392;
assign n6781 = n7626 & n7913;
assign n12893 = ~(n745 ^ n10583);
assign n2215 = n2099 | n12686;
assign n9944 = ~(n4860 ^ n1497);
assign n4489 = ~(n5022 ^ n2864);
assign n7772 = ~(n4790 ^ n3029);
assign n5548 = ~(n7710 | n3531);
assign n4606 = ~(n7874 ^ n4992);
assign n4478 = n2269 | n6987;
assign n5318 = n3337 & n10736;
assign n181 = ~(n808 | n9934);
assign n1623 = n2003 | n12762;
assign n6866 = n7891 & n7610;
assign n3984 = n10142 | n10419;
assign n2348 = n11694 & n4377;
assign n5740 = n3570 & n9972;
assign n5194 = n3219 & n1956;
assign n3743 = ~n7236;
assign n10365 = n8187 | n1851;
assign n5383 = ~n6367;
assign n11512 = ~(n12006 ^ n5953);
assign n3971 = ~(n2791 ^ n278);
assign n10968 = ~(n7154 ^ n7994);
assign n3622 = ~n7684;
assign n4194 = ~(n4263 ^ n8131);
assign n9667 = n499 | n819;
assign n12205 = n1417 | n12331;
assign n7136 = ~n10965;
assign n7032 = n4778 | n8740;
assign n7853 = n5945 | n5012;
assign n10811 = n994 | n6389;
assign n1358 = n7391 | n8524;
assign n12827 = ~(n7958 ^ n9537);
assign n10528 = n4189 & n7456;
assign n4394 = ~(n7511 | n12711);
assign n6794 = n6425 & n10409;
assign n6233 = ~(n103 ^ n1273);
assign n5302 = ~(n706 ^ n12314);
assign n12441 = ~n7546;
assign n2973 = n11742 | n11342;
assign n2147 = n11680 & n5625;
assign n4098 = n8687 | n795;
assign n5654 = n2127 | n3333;
assign n7411 = ~(n10999 ^ n1976);
assign n9712 = ~(n7925 ^ n5545);
assign n4403 = n6583 | n10700;
assign n2914 = ~(n12053 ^ n4464);
assign n12809 = ~n290;
assign n10317 = ~(n12189 ^ n4476);
assign n12837 = n1044 | n6668;
assign n3832 = n7640 | n1489;
assign n1652 = ~(n7484 ^ n10495);
assign n6361 = n3171 & n8421;
assign n6223 = ~(n8913 ^ n4605);
assign n10964 = n10692 & n1210;
assign n10714 = n6044 & n12521;
assign n1958 = ~(n10012 ^ n5837);
assign n12213 = n9878 | n12735;
assign n5696 = n6287 | n10666;
assign n9040 = ~(n7217 | n11996);
assign n5329 = n1675 & n344;
assign n8617 = n3743 | n9280;
assign n3014 = n3115 | n8324;
assign n12216 = ~(n7166 ^ n7878);
assign n9525 = ~n2346;
assign n1732 = ~(n7024 ^ n1942);
assign n3436 = ~(n703 ^ n9491);
assign n11554 = n11272 & n9192;
assign n10961 = ~n6010;
assign n4043 = ~(n4475 | n7910);
assign n6052 = ~(n8122 ^ n1466);
assign n3304 = n12461 | n8212;
assign n11748 = ~n3831;
assign n12844 = n6901 & n12638;
assign n9446 = ~(n7693 | n3330);
assign n2575 = n4001 | n592;
assign n6225 = ~(n7969 | n3357);
assign n6143 = n11799 & n8502;
assign n2336 = n7236 & n10898;
assign n12274 = ~n7823;
assign n7627 = ~(n10837 ^ n10968);
assign n6589 = ~n11554;
assign n6954 = n9875 & n7674;
assign n12611 = n4104 & n8504;
assign n411 = n5925 | n4882;
assign n11543 = n2357 | n12434;
assign n7466 = n10622 | n4876;
assign n4986 = n8187 | n10066;
assign n7794 = ~(n10140 ^ n11763);
assign n2276 = ~(n4358 ^ n10715);
assign n224 = n6977 | n2232;
assign n12392 = ~(n7929 | n732);
assign n11631 = ~n3006;
assign n3911 = ~n1798;
assign n1852 = n686 | n1413;
assign n11364 = n9319 | n5751;
assign n4186 = n1057 | n2441;
assign n5550 = n9584 | n795;
assign n7753 = ~(n9976 ^ n11224);
assign n10985 = ~(n9701 | n2799);
assign n4055 = ~n7171;
assign n3111 = ~(n1515 ^ n6366);
assign n8653 = n6461 & n3148;
assign n3774 = n144 & n7137;
assign n9368 = n2217 | n9144;
assign n9532 = ~n492;
assign n12660 = n5918 | n11409;
assign n3688 = n2069 | n10458;
assign n10653 = ~n4727;
assign n8373 = n9218 | n10559;
assign n12545 = n8583 | n7506;
assign n2631 = n8794 | n2257;
assign n5748 = n12935 & n9808;
assign n4714 = ~(n11179 ^ n10232);
assign n2071 = n12361 | n11820;
assign n10568 = n8127 | n7881;
assign n10049 = n7504 | n224;
assign n6904 = ~(n10537 ^ n9412);
assign n8906 = n7967 & n7261;
assign n12755 = ~(n11029 | n11685);
assign n12064 = ~(n9829 ^ n11256);
assign n8857 = ~(n7980 ^ n6183);
assign n10465 = ~n7209;
assign n9054 = n10270 & n6999;
assign n6283 = n2217 | n12120;
assign n1227 = ~(n10555 ^ n2162);
assign n11190 = ~(n3375 ^ n1986);
assign n4243 = n12071 | n9046;
assign n7377 = n11047 & n7479;
assign n4363 = ~(n6985 ^ n11077);
assign n10860 = n9878 | n12686;
assign n9862 = n6767 & n6250;
assign n10646 = n8354 | n12535;
assign n11589 = n8583 | n12120;
assign n11847 = ~(n590 | n9762);
assign n6144 = ~n11414;
assign n9450 = n8583 | n4642;
assign n4299 = n5690 | n1607;
assign n281 = n8374 | n7235;
assign n3379 = n11154 | n9405;
assign n484 = n7587 & n2343;
assign n1926 = n9997 | n12576;
assign n7971 = n9176 & n12409;
assign n4534 = ~n7664;
assign n7243 = n3743 | n12120;
assign n6538 = n12147 | n85;
assign n12169 = ~(n4676 ^ n8590);
assign n9312 = ~n12404;
assign n9177 = ~(n6564 ^ n2896);
assign n11131 = n11674 & n2726;
assign n4939 = n4674 | n6513;
assign n1059 = ~(n8899 ^ n8565);
assign n1165 = ~(n4461 | n10766);
assign n9921 = n1423 & n5471;
assign n10533 = n5423 & n1528;
assign n4902 = ~(n9205 | n8089);
assign n1670 = n7661 & n8724;
assign n12017 = ~(n1874 | n8233);
assign n6642 = n4782 | n4554;
assign n2621 = n2448 & n3799;
assign n3797 = n8025 & n3280;
assign n3267 = ~n6548;
assign n5883 = n807 | n11775;
assign n4770 = n896 | n10155;
assign n4659 = n12404 & n6493;
assign n5177 = ~(n2752 ^ n9236);
assign n9949 = n3569 | n2707;
assign n5850 = n5915 | n8655;
assign n11002 = n2406 & n8073;
assign n2644 = ~(n5147 ^ n8691);
assign n4991 = ~(n789 ^ n1056);
assign n9937 = n8127 | n7341;
assign n9688 = n9373 | n4875;
assign n5359 = ~n10608;
assign n8266 = ~(n9683 ^ n6559);
assign n12176 = ~(n2192 | n11761);
assign n180 = n7209 | n6807;
assign n6951 = ~n2385;
assign n10579 = ~(n10416 ^ n4569);
assign n11303 = ~(n9196 ^ n4996);
assign n1866 = ~(n12473 ^ n10784);
assign n12644 = ~(n8526 ^ n12250);
assign n12327 = n9370 | n1079;
assign n7808 = ~(n1121 | n11510);
assign n3708 = ~(n4045 | n1635);
assign n12791 = ~(n5959 ^ n10748);
assign n3595 = ~(n7939 ^ n11065);
assign n12369 = n962 | n12771;
assign n3706 = n3743 | n5914;
assign n2300 = n9148 | n4417;
assign n9138 = ~n1338;
assign n2154 = ~(n11834 | n12355);
assign n370 = n12119 | n2259;
assign n5116 = ~(n11233 | n5078);
assign n8058 = ~(n11928 ^ n11308);
assign n19 = n8990 | n1720;
assign n4274 = ~(n6944 | n8783);
assign n4124 = n2217 | n6138;
assign n6623 = ~(n8139 ^ n1473);
assign n5060 = n11927 | n8157;
assign n5429 = n9308 | n9562;
assign n129 = n636 | n10422;
assign n2870 = n2541 | n10427;
assign n11356 = n191 | n8735;
assign n1331 = ~(n9854 ^ n10430);
assign n11959 = n7283 | n5851;
assign n7787 = ~(n4304 ^ n3074);
assign n8292 = ~(n11372 ^ n6918);
assign n5379 = n3659 & n4993;
assign n6690 = ~(n6579 ^ n9997);
assign n8011 = n10157 | n9144;
assign n6334 = ~(n2600 ^ n12332);
assign n9421 = n6174 | n157;
assign n4693 = n3625 | n9031;
assign n3237 = ~(n6636 ^ n6991);
assign n6735 = ~(n10779 ^ n1902);
assign n7110 = ~(n9924 | n2185);
assign n3899 = n11874 & n6793;
assign n7902 = n3078 | n6895;
assign n7080 = ~(n3171 ^ n2831);
assign n10638 = ~(n10362 ^ n1251);
assign n6092 = n8946 & n1593;
assign n9844 = ~n3546;
assign n10977 = ~(n2064 ^ n2267);
assign n3082 = n1574 & n7706;
assign n1487 = ~(n6519 ^ n5549);
assign n3357 = ~(n9657 | n1807);
assign n6881 = n752 | n6197;
assign n212 = ~(n1759 | n11817);
assign n892 = ~n11166;
assign n6483 = ~(n4010 ^ n6300);
assign n8920 = n3127 | n1079;
assign n4630 = n807 | n7876;
assign n4615 = n7449 | n4864;
assign n7893 = n2832 | n3911;
assign n7030 = n5027 & n10477;
assign n10083 = ~(n11613 ^ n5928);
assign n4044 = ~(n12844 | n9183);
assign n355 = ~(n4492 ^ n6521);
assign n5159 = n8631 | n1453;
assign n7452 = ~(n12956 ^ n11030);
assign n11660 = ~(n11959 ^ n8659);
assign n11114 = ~(n5216 ^ n8306);
assign n2972 = ~(n9141 | n5149);
assign n11633 = n6247 & n6973;
assign n7719 = ~(n8897 ^ n9213);
assign n5943 = n7037 & n3232;
assign n599 = n7057 | n3489;
assign n2703 = ~(n7267 | n8470);
assign n8864 = n2047 & n12130;
assign n244 = n9754 | n4491;
assign n8352 = ~(n330 | n2628);
assign n10435 = n191 | n1915;
assign n8893 = ~(n7133 ^ n9918);
assign n41 = n1937 | n995;
assign n7681 = n9240 & n11264;
assign n9752 = n962 | n4875;
assign n11136 = ~(n939 ^ n12824);
assign n5334 = ~n9739;
assign n6168 = n2872 | n6169;
assign n8419 = ~(n3619 | n7592);
assign n1302 = n10668 | n2397;
assign n6281 = ~(n10352 | n8815);
assign n5168 = n8120 & n4248;
assign n9297 = n9807 & n6295;
assign n466 = ~n11800;
assign n7391 = ~n4312;
assign n2784 = n11311 & n8819;
assign n6715 = ~(n2626 ^ n4041);
assign n6297 = n301 & n3154;
assign n2785 = ~(n12759 | n7915);
assign n2656 = ~(n11784 | n9281);
assign n3415 = ~n773;
assign n6823 = n1978 & n5237;
assign n6568 = ~(n4859 ^ n8618);
assign n687 = n8793 | n7736;
assign n6396 = ~n5174;
assign n5229 = ~(n2337 ^ n9930);
assign n8464 = ~(n7992 ^ n8569);
assign n4074 = n8173 & n3834;
assign n3118 = n4510 & n6410;
assign n11663 = ~(n12659 ^ n6846);
assign n1441 = n12647 & n11313;
assign n2128 = n12069 & n1067;
assign n7757 = n11347 | n6405;
assign n11521 = n11443 | n11237;
assign n597 = n870 & n1257;
assign n12595 = ~(n3954 ^ n8955);
assign n6720 = n5455 | n7785;
assign n7130 = n5915 | n9188;
assign n445 = ~(n12491 ^ n6657);
assign n11282 = ~n9438;
assign n4914 = ~(n5582 ^ n1691);
assign n8952 = n5314 & n806;
assign n10020 = n1031 & n8378;
assign n1629 = ~(n3216 ^ n3120);
assign n6976 = ~(n4057 | n176);
assign n1708 = n4628 | n8655;
assign n6304 = n1298 | n11303;
assign n8412 = ~(n1850 ^ n12356);
assign n1469 = n1890 & n3343;
assign n6595 = ~n3000;
assign n11340 = ~(n9836 ^ n249);
assign n9620 = ~(n7867 ^ n2545);
assign n8801 = ~n4337;
assign n7844 = ~(n10884 ^ n3143);
assign n7116 = ~n2226;
assign n11385 = ~(n7871 ^ n6817);
assign n10253 = ~(n2533 ^ n3099);
assign n5362 = ~n8670;
assign n5558 = n5236 & n10301;
assign n9938 = ~(n7323 ^ n7518);
assign n11525 = n1432 | n4923;
assign n4798 = n7774 & n7127;
assign n4461 = ~(n3196 | n2274);
assign n7309 = n5355 | n12843;
assign n435 = ~(n2234 ^ n12414);
assign n7189 = ~(n10980 ^ n4614);
assign n12895 = n2476 & n9102;
assign n7481 = ~(n9383 | n8195);
assign n1995 = n686 | n5540;
assign n2787 = n7550 & n12390;
assign n2655 = ~(n8603 | n6969);
assign n4103 = n11905 | n11186;
assign n1293 = ~(n12914 | n10920);
assign n5374 = n11292 | n9517;
assign n10291 = n2784 & n12315;
assign n10746 = ~(n11613 | n10710);
assign n8397 = n11966 | n5091;
assign n6354 = ~n6318;
assign n2082 = ~n7699;
assign n2533 = n1825 & n3229;
assign n10331 = ~n9130;
assign n11873 = n4057 & n176;
assign n5994 = ~n2610;
assign n4816 = n9487 | n3897;
assign n12009 = n10993 | n8928;
assign n12177 = n3746 | n7952;
assign n1939 = ~(n3646 ^ n1201);
assign n4993 = n6577 | n11122;
assign n7951 = n10139 & n3615;
assign n5588 = ~(n4908 ^ n12345);
assign n7591 = n10535 | n1457;
assign n3302 = n4018 & n9159;
assign n4513 = ~(n5241 ^ n245);
assign n2712 = n8034 | n5868;
assign n9442 = ~(n9337 ^ n5587);
assign n1876 = ~(n11760 ^ n1301);
assign n3537 = ~(n2684 | n9962);
assign n61 = n5765 | n6138;
assign n6903 = n11843 & n6440;
assign n9420 = ~n6899;
assign n144 = n12119 | n12883;
assign n1329 = ~(n7563 ^ n6609);
assign n9948 = n9918 | n7575;
assign n9717 = ~(n2885 | n11989);
assign n6929 = n10835 | n5086;
assign n7672 = n4911 | n12843;
assign n5370 = n11887 | n1932;
assign n10753 = n2606 & n11485;
assign n5454 = ~(n452 ^ n12646);
assign n2199 = ~(n8180 ^ n761);
assign n8500 = ~(n9974 ^ n3392);
assign n479 = ~(n679 ^ n9045);
assign n8511 = n7944 | n2594;
assign n7750 = n10729 | n8018;
assign n5803 = ~n12081;
assign n4879 = ~(n9538 ^ n10503);
assign n9479 = n8354 | n3224;
assign n2808 = n3018 & n6810;
assign n8159 = ~(n2043 ^ n7717);
assign n3822 = n6560 | n3741;
assign n4491 = ~(n4815 ^ n10041);
assign n11926 = ~n7984;
assign n10550 = ~(n3131 ^ n10813);
assign n4250 = n8428 | n3903;
assign n5129 = ~(n1123 | n396);
assign n1144 = ~n7200;
assign n3511 = n11613 & n10710;
assign n6582 = n319 | n1234;
assign n10590 = n2217 | n9280;
assign n5560 = n7380 | n1634;
assign n10251 = ~(n11280 | n6141);
assign n8302 = ~n1213;
assign n4898 = ~(n6248 ^ n3497);
assign n4472 = n2424 & n12846;
assign n9770 = n2217 | n3451;
assign n4818 = ~n2802;
assign n4682 = n2176 ^ n4779;
assign n7451 = ~(n1598 ^ n8724);
assign n5865 = n1272 & n8761;
assign n2854 = n12853 | n3924;
assign n175 = n1659 | n4714;
assign n6199 = n5365 | n479;
assign n2691 = ~(n11499 ^ n1216);
assign n5782 = ~n4233;
assign n11984 = n191 | n1546;
assign n12465 = ~n6723;
assign n8194 = n9170 | n1851;
assign n2616 = n7391 | n5497;
assign n5185 = ~n1339;
assign n3816 = n5828 | n5186;
assign n1340 = ~(n8052 | n7989);
assign n9881 = n4002 | n6061;
assign n9330 = ~(n3386 ^ n9746);
assign n6375 = n9459 | n2193;
assign n4772 = n2931 & n4376;
assign n5059 = n12541 & n12031;
assign n11479 = ~(n4918 ^ n1268);
assign n10935 = ~n11201;
assign n3085 = ~(n6892 ^ n12469);
assign n7910 = ~(n12522 ^ n12928);
assign n7107 = n9836 | n8081;
assign n2734 = ~n8702;
assign n5281 = n2872 | n6455;
assign n1057 = n3746 | n11775;
assign n8555 = n5895 & n11374;
assign n91 = n3127 | n1162;
assign n3888 = ~(n1590 ^ n1954);
assign n1549 = ~n8562;
assign n6557 = ~(n7481 | n9494);
assign n8570 = ~n3219;
assign n11982 = ~(n8159 ^ n2238);
assign n12512 = n2534 | n4747;
assign n1295 = ~(n9266 ^ n8711);
assign n560 = n2140 | n12656;
assign n4475 = n9450 & n8067;
assign n2758 = ~(n3943 ^ n4262);
assign n10202 = n10157 | n4875;
assign n8754 = ~(n5604 ^ n8837);
assign n5446 = ~(n6697 ^ n12225);
assign n7349 = ~(n610 ^ n5647);
assign n8926 = n9670 | n10048;
assign n10389 = n8674 & n5642;
assign n11499 = ~(n9153 ^ n8379);
assign n3209 = ~(n4730 ^ n12060);
assign n859 = ~(n12355 ^ n10125);
assign n2372 = ~(n5267 ^ n9406);
assign n1666 = ~(n2359 | n3212);
assign n12182 = n7116 | n1413;
assign n6527 = n191 | n11827;
assign n12558 = n11134 & n401;
assign n1000 = ~n8631;
assign n11609 = ~(n4905 ^ n620);
assign n5527 = ~n8816;
assign n1768 = ~(n3689 | n9332);
assign n11447 = ~(n4961 ^ n231);
assign n10845 = n7862 & n1798;
assign n7974 = ~n1241;
assign n11343 = ~n6626;
assign n10288 = n9373 | n12120;
assign n3193 = n10040 | n7990;
assign n1138 = ~(n12461 ^ n12672);
assign n9023 = ~n1648;
assign n3319 = ~(n10585 ^ n8728);
assign n11936 = n7160 & n11922;
assign n12272 = ~(n6929 ^ n275);
assign n11398 = ~(n6836 ^ n332);
assign n8571 = ~(n2618 ^ n4564);
assign n2342 = ~(n2721 ^ n11628);
assign n3268 = ~(n12306 ^ n9351);
assign n8183 = ~n3689;
assign n5406 = ~n7096;
assign n5682 = n8175 | n11003;
assign n12021 = ~n11275;
assign n3154 = n4603 | n10468;
assign n8437 = ~(n2677 ^ n9579);
assign n7982 = n9301 | n2028;
assign n1660 = n3127 | n6389;
assign n2056 = n8870 | n3924;
assign n989 = ~n2564;
assign n2709 = n6625 & n12959;
assign n6390 = n11278 & n441;
assign n1690 = ~(n10202 ^ n6271);
assign n8427 = ~(n3538 | n682);
assign n2952 = n10879 | n5497;
assign n11918 = ~(n3689 ^ n206);
assign n11378 = n4314 & n9089;
assign n5463 = ~n8990;
assign n1187 = n1337 & n4054;
assign n2014 = n3252 | n12542;
assign n8148 = n337 & n12329;
assign n463 = ~n1872;
assign n3274 = n8737 | n5874;
assign n625 = n3648 & n9664;
assign n8365 = ~n4771;
assign n9512 = n6294 & n2498;
assign n5433 = ~(n2599 ^ n1083);
assign n3577 = n10463 & n5119;
assign n12582 = ~(n3062 ^ n2242);
assign n6619 = ~(n3007 ^ n8561);
assign n322 = ~(n5169 ^ n42);
assign n313 = n5765 | n2020;
assign n4697 = n3127 | n4242;
assign n6465 = n4085 & n6000;
assign n7933 = ~n7716;
assign n2489 = ~(n11530 ^ n8625);
assign n7906 = n1699 | n8655;
assign n4296 = ~(n8732 ^ n1280);
assign n12029 = ~n4742;
assign n10749 = n7370 | n3125;
assign n1674 = ~(n1953 ^ n10276);
assign n7307 = n10555 & n7791;
assign n10706 = n5107 & n258;
assign n10810 = n994 | n8859;
assign n104 = ~(n1687 ^ n3785);
assign n10470 = n1461 & n3374;
assign n937 = n10847 & n12626;
assign n11345 = n1102 & n468;
assign n7390 = n12518 & n10688;
assign n7432 = n9834 | n7467;
assign n10873 = ~(n3857 ^ n9008);
assign n2172 = ~(n5144 ^ n5705);
assign n9910 = ~(n2250 ^ n1977);
assign n3937 = n7978 | n9566;
assign n3063 = ~(n969 ^ n5046);
assign n3170 = n11290 & n497;
assign n4550 = n8416 & n2933;
assign n8308 = n5809 | n7382;
assign n12786 = n10378 | n2620;
assign n908 = n279 & n2876;
assign n7100 = n5575 | n7952;
assign n1743 = n12881 & n10884;
assign n10737 = n8354 | n5468;
assign n2880 = ~(n4846 ^ n11562);
assign n6228 = ~(n1029 ^ n8639);
assign n9208 = n1746 | n2404;
assign n9174 = n6078 & n2672;
assign n1557 = ~n6834;
assign n1101 = n4290 | n10113;
assign n4553 = n253 ^ n11227;
assign n6628 = n12757 & n5057;
assign n7863 = ~(n7407 ^ n10662);
assign n2950 = n5735 & n1058;
assign n5166 = n2217 | n795;
assign n5291 = n8276 & n9640;
assign n1758 = ~(n908 | n6976);
assign n8769 = ~(n12033 ^ n6781);
assign n10776 = ~(n5333 ^ n257);
assign n9826 = ~n9662;
assign n2332 = n5765 | n10916;
assign n7782 = n10169 & n1411;
assign n10014 = ~(n6486 ^ n1464);
assign n198 = ~n5608;
assign n79 = ~(n8295 ^ n2862);
assign n8197 = ~(n352 ^ n8973);
assign n6714 = n4635 & n12369;
assign n4149 = ~n3775;
assign n2454 = ~n3710;
assign n12935 = n2217 | n8830;
assign n11966 = n2822 & n5265;
assign n1737 = n7864 | n8099;
assign n2048 = ~(n5108 | n9198);
assign n12642 = n10620 & n11302;
assign n12571 = n4145 & n11459;
assign n7318 = n3820 | n2020;
assign n670 = n3465 & n9147;
assign n10666 = ~(n1899 ^ n9575);
assign n7514 = ~(n2424 ^ n8822);
assign n7643 = n11958 | n6114;
assign n2568 = ~(n2130 ^ n2037);
assign n1116 = ~n10423;
assign n12479 = ~n10255;
assign n9265 = n8384 & n806;
assign n3131 = n2099 | n530;
assign n5260 = ~(n3030 ^ n8394);
assign n8453 = n9674 | n2691;
assign n9604 = ~(n5229 | n12653);
assign n2233 = ~(n8591 ^ n3731);
assign n1477 = ~(n8960 | n12466);
assign n8232 = n8026 | n3468;
assign n1085 = n4943 | n3189;
assign n49 = n3674 & n1636;
assign n6655 = ~(n9638 ^ n3555);
assign n4988 = ~(n4554 ^ n3935);
assign n1429 = ~(n11641 ^ n6333);
assign n3598 = ~(n11353 | n10000);
assign n6871 = n11285 | n6537;
assign n3290 = n78 | n1934;
assign n12703 = n7495 | n7424;
assign n6909 = n3591 | n8082;
assign n6360 = ~n3330;
assign n7940 = n12172 & n7096;
assign n967 = ~n2717;
assign n3364 = n5171 | n4317;
assign n5196 = n10103 & n411;
assign n1967 = ~n12087;
assign n6914 = n3746 | n7425;
assign n3853 = n11335 & n6518;
assign n6983 = ~(n1206 ^ n5300);
assign n9776 = n11433 | n2232;
assign n1779 = ~(n2557 | n10923);
assign n9032 = ~(n128 ^ n5460);
assign n2120 = ~n157;
assign n9246 = n7388 & n12947;
assign n5842 = ~(n11745 ^ n4969);
assign n6786 = n12391 & n6806;
assign n7527 = n8583 | n8643;
assign n5595 = ~(n8568 ^ n9116);
assign n7980 = ~(n12901 | n8105);
assign n8691 = n11719 | n11746;
assign n2801 = n4445 | n11105;
assign n1769 = ~(n6500 ^ n6593);
assign n9886 = ~n8284;
assign n5793 = n12119 | n6071;
assign n1785 = ~(n5310 | n5912);
assign n3419 = ~(n6669 ^ n3568);
assign n4079 = n11222 & n9111;
assign n983 = ~(n12795 ^ n9407);
assign n11103 = ~n3296;
assign n2809 = ~(n6292 | n9824);
assign n3535 = ~(n5273 ^ n108);
assign n3351 = n1726 & n3718;
assign n2791 = n3743 | n7921;
assign n11389 = ~n5048;
assign n290 = n10006 | n10659;
assign n123 = ~(n3509 ^ n1188);
assign n2669 = n2447 & n9150;
assign n8827 = ~(n787 ^ n12944);
assign n4002 = n10142 | n561;
assign n9105 = n6777 | n2908;
assign n52 = ~(n11856 ^ n11998);
assign n7217 = n9172 & n11949;
assign n7174 = ~(n2285 ^ n7801);
assign n3194 = n8127 | n11827;
assign n8382 = n7123 | n10074;
assign n1161 = n4956 | n5000;
assign n3662 = ~(n8810 ^ n318);
assign n2727 = n1599 | n11816;
assign n8035 = n3939 & n1368;
assign n2132 = ~(n12457 ^ n3366);
assign n5096 = n9000 & n5391;
assign n4555 = n7760 | n11617;
assign n10402 = n12237 | n10854;
assign n6859 = n2808 | n11903;
assign n905 = n4498 | n1079;
assign n8874 = ~(n99 ^ n11008);
assign n8812 = n9900 & n5063;
assign n306 = n9373 | n1509;
assign n7143 = n686 | n12816;
assign n6065 = n4824 | n11273;
assign n6531 = n3746 | n1413;
assign n9370 = ~n3172;
assign n10324 = ~(n12165 ^ n2720);
assign n10421 = ~(n3189 ^ n6176);
assign n8784 = n10572 & n2741;
assign n4929 = n5739 | n10241;
assign n3428 = n3096 | n2232;
assign n5520 = ~(n6449 | n4626);
assign n3031 = ~(n856 ^ n7324);
assign n2379 = n12797 | n6169;
assign n1795 = ~(n9925 ^ n8658);
assign n12798 = ~(n3018 | n6810);
assign n7234 = n12361 | n11410;
assign n12958 = ~n8912;
assign n4782 = ~n9967;
assign n4713 = n6718 | n609;
assign n12848 = ~(n4741 | n4384);
assign n811 = n5224 | n3851;
assign n4197 = n9801 | n8528;
assign n5480 = ~(n12691 ^ n306);
assign n9576 = n11552 | n8643;
assign n6649 = ~(n6129 | n4700);
assign n5687 = n8498 | n7279;
assign n6000 = ~n10245;
assign n4823 = ~(n1730 | n1772);
assign n7816 = ~n3204;
assign n8329 = n9690 & n5546;
assign n9263 = n2107 & n5239;
assign n2484 = ~(n9296 ^ n2712);
assign n8538 = n12231 & n3958;
assign n2696 = n7912 | n4136;
assign n12504 = n4668 | n5572;
assign n5928 = n962 | n1509;
assign n4868 = ~(n3513 ^ n10491);
assign n106 = ~(n5947 ^ n5261);
assign n8346 = ~(n6379 | n9484);
assign n8133 = ~(n10613 ^ n12740);
assign n8208 = n11958 | n2754;
assign n7873 = ~(n219 ^ n10523);
assign n12794 = n10770 & n4048;
assign n8506 = n11747 | n4058;
assign n8279 = n37 | n11316;
assign n11016 = ~(n4512 ^ n9986);
assign n8015 = ~(n847 ^ n11950);
assign n8446 = n9758 & n9408;
assign n8306 = n931 | n1735;
assign n10635 = n9420 & n5665;
assign n11882 = n11433 | n6169;
assign n6212 = ~n10778;
assign n11418 = ~n1776;
assign n10189 = ~(n8677 ^ n1369);
assign n2389 = ~(n4462 ^ n11363);
assign n10286 = n4678 | n10234;
assign n1583 = n1670 | n8700;
assign n2586 = ~(n9865 ^ n8654);
assign n7342 = ~(n7566 ^ n2932);
assign n3182 = ~(n5998 ^ n9577);
assign n11276 = ~(n9205 ^ n1069);
assign n4192 = ~(n8310 ^ n8450);
assign n4847 = ~(n10926 ^ n5600);
assign n12740 = n9584 | n4474;
assign n6371 = n855 & n10699;
assign n8289 = ~(n4484 ^ n1777);
assign n6445 = ~(n9566 ^ n336);
assign n3844 = ~(n9937 ^ n6224);
assign n2810 = n3746 | n184;
assign n9220 = ~(n4649 | n8075);
assign n4963 = ~(n8536 ^ n1656);
assign n4584 = n8189 & n5797;
assign n590 = n4434 & n1584;
assign n6798 = n8757 & n3021;
assign n4807 = ~(n2948 ^ n11083);
assign n683 = n12853 | n12080;
assign n9171 = n7501 & n1628;
assign n496 = n5915 | n530;
assign n802 = n9887 & n9226;
assign n5206 = n7258 & n2988;
assign n5021 = ~(n1552 ^ n2091);
assign n11874 = n12691 | n6543;
assign n3040 = ~(n1563 | n7062);
assign n286 = ~(n4070 ^ n4017);
assign n4937 = ~(n7118 | n4093);
assign n146 = ~(n10243 ^ n9707);
assign n1399 = ~n4581;
assign n10218 = ~(n1439 ^ n4412);
assign n12902 = ~(n4497 ^ n731);
assign n3872 = n12180 | n4558;
assign n5017 = ~n6328;
assign n11871 = ~(n6652 | n6046);
assign n6939 = n10142 | n4775;
assign n8964 = n9389 | n1455;
assign n6059 = n4843 | n11314;
assign n10243 = ~(n7640 ^ n2396);
assign n6625 = n5530 | n8648;
assign n3250 = n6797 & n12489;
assign n4119 = n8656 & n3144;
assign n2249 = n2703 | n850;
assign n1816 = ~(n7501 | n1628);
assign n7232 = n11400 & n7590;
assign n341 = ~n8754;
assign n408 = ~(n2228 ^ n5286);
assign n968 = ~(n10795 | n12909);
assign n12557 = n10835 | n8745;
assign n12765 = ~(n11140 ^ n7163);
assign n7173 = n11445 & n247;
assign n755 = ~(n9674 ^ n2691);
assign n12502 = n9341 & n8154;
assign n12688 = n2693 & n11525;
assign n1784 = n6373 | n4474;
assign n5707 = ~(n8372 ^ n1480);
assign n5841 = n6977 | n7425;
assign n5807 = ~(n1088 ^ n1479);
assign n2360 = ~(n1398 ^ n2338);
assign n5598 = n4022 & n9318;
assign n3093 = n9389 | n4400;
assign n10183 = ~n8743;
assign n8272 = n5179 & n8417;
assign n6994 = ~(n3368 ^ n1326);
assign n12555 = ~n10493;
assign n9821 = n12910 | n5296;
assign n1285 = n928 & n6381;
assign n85 = n7895 & n89;
assign n6764 = ~n9872;
assign n5092 = ~n4304;
assign n3683 = ~(n589 ^ n12321);
assign n8711 = n5915 | n5468;
assign n5138 = ~(n10070 | n7997);
assign n10412 = n8894 | n10256;
assign n4023 = ~(n11429 ^ n9761);
assign n12770 = n3970 & n1364;
assign n650 = ~(n12601 ^ n4149);
assign n7091 = n1305 & n1928;
assign n885 = n2099 | n12124;
assign n12451 = ~n10448;
assign n6173 = n2711 & n2807;
assign n6192 = ~(n7079 ^ n9911);
assign n8001 = ~(n11741 | n1447);
assign n12613 = ~n9419;
assign n12942 = ~n2828;
assign n10941 = n6618 & n12588;
assign n2710 = ~(n392 | n9940);
assign n1216 = n12197 & n8637;
assign n10397 = n8896 & n4710;
assign n6349 = n10338 & n6123;
assign n8542 = ~(n4268 ^ n5586);
assign n5950 = n9074 & n972;
assign n11606 = ~(n3336 | n3752);
assign n11706 = n12694 & n7386;
assign n11865 = ~(n7146 | n7691);
assign n5539 = ~(n9034 ^ n11359);
assign n12016 = ~(n7819 | n7339);
assign n12814 = n8118 | n9965;
assign n11438 = n111 | n4618;
assign n12546 = ~n6556;
assign n12295 = ~(n6746 ^ n3119);
assign n5960 = ~n11345;
assign n4763 = n10339 | n8740;
assign n11376 = ~n6262;
assign n11086 = ~(n9016 ^ n10026);
assign n9162 = ~(n8268 ^ n10669);
assign n7257 = ~(n11415 ^ n12606);
assign n5862 = ~n9380;
assign n5877 = ~(n7620 | n1724);
assign n8625 = ~(n2400 ^ n2705);
assign n8007 = ~(n10403 | n6870);
assign n10374 = n5355 | n11430;
assign n4876 = ~(n6406 | n3542);
assign n312 = n2762 & n5782;
assign n3543 = ~(n6187 ^ n7403);
assign n12833 = ~(n6390 | n8238);
assign n8507 = n1396 & n10946;
assign n7223 = n10147 | n12838;
assign n6006 = n9079 & n6414;
assign n8917 = ~(n2957 ^ n3671);
assign n5058 = n11043 | n9721;
assign n6878 = ~n11749;
assign n6998 = n678 & n1703;
assign n3423 = ~(n4346 ^ n1308);
assign n8681 = ~(n10036 ^ n3526);
assign n11172 = ~(n7229 ^ n10749);
assign n5426 = ~n1373;
assign n12400 = n249 | n11480;
assign n12008 = ~(n6081 ^ n12609);
assign n7463 = ~(n9581 ^ n10924);
assign n887 = ~(n12258 ^ n4705);
assign n5348 = n9373 | n28;
assign n12623 = n5303 & n3393;
assign n4075 = n807 | n2815;
assign n12397 = ~n3895;
assign n5220 = ~(n229 ^ n11915);
assign n1433 = n1941 | n11896;
assign n10045 = n2459 | n4594;
assign n7081 = n5677 & n11125;
assign n3863 = ~(n6237 ^ n12917);
assign n3315 = ~(n12308 ^ n227);
assign n11515 = ~(n8999 ^ n11371);
assign n9553 = ~(n11724 ^ n9919);
assign n3510 = n2602 & n4014;
assign n11979 = ~(n5277 | n7517);
assign n5613 = ~(n4700 ^ n6129);
assign n10404 = n3326 & n2364;
assign n11337 = ~(n7401 ^ n6412);
assign n5135 = ~(n4247 ^ n554);
assign n2599 = n5575 | n11410;
assign n3752 = ~(n1859 ^ n12339);
assign n6748 = ~(n1878 ^ n10861);
assign n12873 = n7449 | n6138;
assign n2708 = ~(n7749 ^ n3281);
assign n12056 = n4602 & n2676;
assign n11801 = n11026 | n4875;
assign n2532 = ~(n1722 ^ n1055);
assign n773 = n11389 | n1159;
assign n9302 = ~n7177;
assign n460 = ~(n1339 ^ n6299);
assign n4025 = ~(n6569 | n12796);
assign n4 = n270 | n11231;
assign n8966 = n6031 | n3787;
assign n6438 = ~(n7564 ^ n8019);
assign n7544 = n1966 | n7784;
assign n7262 = ~(n1672 ^ n2553);
assign n3942 = ~(n2345 ^ n8444);
assign n3173 = ~(n2555 ^ n12042);
assign n204 = n4777 | n7475;
assign n7367 = ~n3604;
assign n2597 = n7688 | n11465;
assign n10582 = ~n1151;
assign n1099 = n763 | n5976;
assign n5057 = ~n12118;
assign n4692 = ~n1687;
assign n1891 = ~(n3048 | n5978);
assign n6791 = ~(n2854 ^ n7701);
assign n7821 = ~(n292 ^ n2428);
assign n11381 = n8438 | n12190;
assign n11011 = ~n6209;
assign n6497 = ~(n1348 ^ n10372);
assign n4599 = ~n8963;
assign n784 = n8481 & n1048;
assign n9579 = n8572 & n11579;
assign n11534 = n3558 | n1927;
assign n3260 = n989 | n1162;
assign n12888 = ~n39;
assign n378 = ~n10155;
assign n9168 = ~(n10061 | n10316);
assign n9417 = ~n10362;
assign n9994 = ~(n3620 ^ n5718);
assign n4733 = ~(n12019 ^ n8661);
assign n10605 = ~(n12464 ^ n2122);
assign n1582 = n1871 & n3515;
assign n5504 = ~(n495 ^ n1189);
assign n2840 = n5414 | n10759;
assign n109 = ~n5517;
assign n4523 = ~(n4514 ^ n7677);
assign n2770 = ~(n2842 | n6424);
assign n9045 = ~(n5328 ^ n2683);
assign n695 = n2217 | n4864;
assign n9389 = ~n4189;
assign n12022 = n12960 & n10487;
assign n542 = n725 & n8146;
assign n3569 = n5765 | n28;
assign n4341 = ~(n10180 ^ n4234);
assign n5046 = n7439 & n5891;
assign n12600 = ~(n10226 ^ n9680);
assign n6861 = n607 & n419;
assign n5435 = ~(n1385 ^ n4009);
assign n4213 = ~(n588 ^ n156);
assign n3048 = ~n37;
assign n314 = ~(n8789 ^ n1733);
assign n11468 = n6718 | n4642;
assign n9147 = ~n7131;
assign n11611 = ~n1865;
assign n7786 = ~n1264;
assign n179 = ~(n5023 ^ n10401);
assign n7920 = n11220 & n7829;
assign n11786 = ~(n3879 | n10499);
assign n9014 = n2479 & n2317;
assign n4587 = ~n7642;
assign n11884 = n4565 | n1281;
assign n11191 = ~n2861;
assign n5757 = n9370 | n510;
assign n9817 = n24 & n7334;
assign n9769 = ~(n8232 | n7679);
assign n6326 = ~(n6233 ^ n11513);
assign n2273 = ~(n5423 ^ n9921);
assign n11930 = n9370 | n11746;
assign n10966 = ~n2311;
assign n5339 = ~n7775;
assign n1650 = ~(n7864 ^ n8099);
assign n3310 = n7116 | n11775;
assign n7393 = n5530 | n12883;
assign n8863 = ~(n6694 ^ n11733);
assign n11639 = ~(n10876 | n10982);
assign n5884 = n5679 & n2963;
assign n4164 = ~n4920;
assign n12779 = ~(n2903 ^ n10734);
assign n6534 = n8026 | n3903;
assign n6392 = ~(n10341 ^ n6357);
assign n4422 = ~(n5090 ^ n1993);
assign n9453 = ~(n12658 ^ n8392);
assign n10453 = n2832 | n1455;
assign n3645 = ~(n4580 | n7561);
assign n9348 = n7028 & n898;
assign n9911 = ~(n3811 ^ n7135);
assign n6114 = ~n7730;
assign n6474 = n9052 & n2716;
assign n2163 = n4343 | n6513;
assign n2429 = n4605 & n1678;
assign n6900 = n8428 | n7395;
assign n2205 = ~(n1341 ^ n3362);
assign n2778 = ~(n2045 ^ n11274);
assign n7284 = n2456 | n8655;
assign n7767 = ~n4529;
assign n12783 = ~(n12091 ^ n12682);
assign n6322 = ~(n5149 ^ n6035);
assign n4875 = ~n4086;
assign n6430 = n7834 & n8364;
assign n5235 = ~(n7121 ^ n8944);
assign n2036 = n5915 | n3924;
assign n688 = n1051 | n995;
assign n6485 = ~n9054;
assign n4068 = n9027 & n1588;
assign n1726 = n10142 | n1851;
assign n3238 = ~(n12563 ^ n9703);
assign n4429 = ~(n1411 ^ n1925);
assign n12042 = ~(n12035 ^ n6063);
assign n6551 = n8690 & n3904;
assign n4942 = ~(n8219 ^ n6815);
assign n12513 = n7449 | n609;
assign n909 = ~(n4525 ^ n11382);
assign n11353 = n1025 & n4933;
assign n9216 = n15 | n5218;
assign n11298 = ~(n3665 ^ n9355);
assign n5870 = ~(n12571 ^ n619);
assign n9020 = ~(n1583 ^ n4473);
assign n2305 = n752 | n5540;
assign n5624 = ~(n940 ^ n9984);
assign n11680 = n1043 | n11532;
assign n1530 = ~(n1754 | n2291);
assign n7656 = n11576 & n1712;
assign n9711 = ~(n8331 ^ n5351);
assign n5459 = n12497 & n7033;
assign n4984 = ~(n2610 ^ n9541);
assign n7303 = n2456 | n4913;
assign n7964 = n2136 | n10652;
assign n11718 = ~(n7448 | n3231);
assign n8257 = ~n12571;
assign n5308 = ~(n2447 ^ n2313);
assign n9996 = n5680 & n4883;
assign n9868 = ~(n7487 ^ n8251);
assign n6298 = n9564 & n706;
assign n4980 = n10339 | n6513;
assign n10708 = ~(n9245 ^ n8383);
assign n12231 = n3989 & n5970;
assign n10934 = n5765 | n9280;
assign n7599 = n8738 | n4654;
assign n7271 = n3743 | n9078;
assign n10900 = n12142 & n4458;
assign n6814 = n5355 | n1738;
assign n1539 = ~n2087;
assign n11709 = n6863 | n4427;
assign n6219 = n2376 | n3679;
assign n2630 = n12748 | n1336;
assign n4992 = n9389 | n5497;
assign n267 = ~(n956 ^ n8680);
assign n3176 = n5738 & n9642;
assign n1821 = n7562 & n12889;
assign n8776 = ~(n8975 ^ n1619);
assign n12425 = n7713 & n4012;
assign n6506 = n5689 & n10134;
assign n11380 = ~(n7920 ^ n8715);
assign n4411 = ~n1723;
assign n266 = n2865 | n1942;
assign n3041 = ~(n4446 | n1491);
assign n5011 = n4559 | n10651;
assign n493 = n6395 | n2806;
assign n643 = ~(n5087 | n5357);
assign n558 = n11069 & n10056;
assign n7113 = n7624 | n3139;
assign n8424 = ~(n5673 ^ n8784);
assign n4519 = n22 | n5261;
assign n12303 = n8211 & n12745;
assign n11278 = n526 | n12480;
assign n2241 = ~(n122 ^ n11504);
assign n3276 = n1886 & n4382;
assign n8586 = ~(n3749 ^ n8995);
assign n3263 = ~(n140 ^ n7811);
assign n7442 = ~(n3807 ^ n1967);
assign n7947 = n9231 | n6051;
assign n1134 = ~n634;
assign n6857 = n6373 | n3606;
assign n9597 = ~(n694 | n1527);
assign n11052 = ~(n4122 ^ n4225);
assign n634 = n556 & n9483;
assign n3846 = n5850 & n1347;
assign n9603 = n11478 & n12489;
assign n8301 = ~n1242;
assign n613 = n10142 | n12843;
assign n406 = ~n8914;
assign n11544 = n10157 | n6922;
assign n8064 = n5542 & n7234;
assign n11081 = ~(n11276 ^ n5298);
assign n9795 = n10199 & n7637;
assign n12617 = ~n9519;
assign n10875 = ~(n2781 ^ n2132);
assign n2544 = ~(n11679 ^ n1702);
assign n12538 = ~(n3065 | n577);
assign n10105 = n5999 | n7753;
assign n4276 = ~(n12788 ^ n1120);
assign n969 = n7391 | n1079;
assign n7103 = ~(n9887 ^ n9226);
assign n6377 = n1881 | n3482;
assign n5488 = n3051 | n2323;
assign n12227 = n4628 | n3924;
assign n12186 = ~n10644;
assign n5946 = ~n935;
assign n353 = ~(n8242 ^ n6266);
assign n8440 = ~(n3138 ^ n5747);
assign n4087 = ~(n9228 ^ n776);
assign n3966 = ~(n8534 ^ n12791);
assign n1425 = n6571 | n11787;
assign n417 = ~(n7501 ^ n5037);
assign n4540 = ~n8163;
assign n10917 = n8097 & n3621;
assign n11522 = ~(n331 ^ n9121);
assign n10146 = n9431 & n421;
assign n6351 = n6635 & n9863;
assign n10995 = n12797 | n2815;
assign n881 = n12933 & n4152;
assign n1847 = ~(n3521 ^ n6605);
assign n11327 = n10251 | n7741;
assign n9507 = n10551 & n7988;
assign n1262 = ~(n9784 ^ n945);
assign n4727 = n8336 & n12709;
assign n6824 = n12141 & n11811;
assign n2223 = n5809 | n12735;
assign n8519 = ~n4650;
assign n9485 = n11821 & n1798;
assign n12174 = ~(n1808 ^ n2210);
assign n1846 = ~(n3474 | n5126);
assign n6512 = ~(n4017 | n4070);
assign n338 = n11782 & n5114;
assign n12270 = ~(n5791 ^ n3300);
assign n9104 = ~n6988;
assign n158 = n4911 | n7881;
assign n11858 = n3196 ^ n10766;
assign n8903 = n5575 | n10903;
assign n1717 = ~n5948;
assign n11678 = n4961 & n231;
assign n11627 = ~n9395;
assign n10642 = n8921 | n1555;
assign n1072 = n5355 | n6402;
assign n6501 = n4243 & n8520;
assign n921 = ~(n7936 | n1021);
assign n5642 = n3756 & n2970;
assign n9530 = n10196 | n4474;
assign n5771 = n1462 | n10617;
assign n9572 = n6376 & n7343;
assign n12499 = ~n9896;
assign n6448 = ~(n8675 | n9295);
assign n8392 = n6888 & n11121;
assign n8794 = n7058 & n6484;
assign n9647 = ~(n11392 ^ n10994);
assign n6405 = ~(n2303 ^ n6676);
assign n7277 = n11126 & n687;
assign n8969 = ~n4756;
assign n9786 = n2595 | n920;
assign n11109 = n6977 | n3421;
assign n3218 = n8552 | n10854;
assign n9646 = ~(n11094 ^ n7005);
assign n11258 = ~(n9176 ^ n11849);
assign n3575 = ~(n7527 ^ n5344);
assign n899 = n10157 | n5759;
assign n2378 = n1663 & n4964;
assign n1490 = ~(n3403 ^ n3675);
assign n4347 = n12841 | n6563;
assign n7912 = n7283 | n7881;
assign n8048 = n659 | n2151;
assign n2110 = ~(n5358 ^ n764);
assign n9872 = n7177 & n8407;
assign n11561 = ~(n9894 ^ n5047);
assign n12863 = ~(n10377 ^ n11);
assign n4827 = n6931 & n4506;
assign n2209 = n5355 | n11827;
assign n4908 = n2538 & n2861;
assign n8585 = n12119 | n10854;
assign n12576 = n6579 & n3093;
assign n5340 = n8371 | n4073;
assign n6178 = ~(n8579 ^ n1647);
assign n1439 = n6743 & n4503;
assign n9875 = n9653 | n3928;
assign n9356 = ~(n4949 ^ n3083);
assign n4096 = ~n5380;
assign n8483 = ~(n9799 ^ n12802);
assign n3087 = n10750 | n826;
assign n3954 = n12237 | n1932;
assign n9139 = ~(n2028 ^ n3245);
assign n8930 = ~(n7587 ^ n10511);
assign n12072 = ~(n5523 ^ n12349);
assign n11238 = ~n8660;
assign n9151 = n9835 | n11151;
assign n254 = ~n4135;
assign n10570 = n7899 & n5485;
assign n12580 = ~n3945;
assign n11887 = ~n6797;
assign n1194 = ~(n12155 ^ n10506);
assign n7916 = n10142 | n9589;
assign n7797 = n9849 & n8268;
assign n8444 = ~(n4110 ^ n11565);
assign n1856 = n6277 & n8368;
assign n6505 = ~n5869;
assign n6116 = ~(n4360 ^ n702);
assign n7247 = ~(n11899 ^ n477);
assign n11074 = n4932 | n12548;
assign n11388 = n9454 & n6302;
assign n3794 = ~(n5877 | n653);
assign n2807 = n11608 | n6029;
assign n2816 = n8617 | n2375;
assign n10290 = n11521 & n7438;
assign n5351 = ~n6574;
assign n11711 = n3197 & n6057;
assign n10639 = n12178 & n5402;
assign n11653 = n2579 | n4751;
assign n3275 = ~n4664;
assign n3636 = ~n12068;
assign n7718 = n11923 | n4474;
assign n12665 = n854 | n1710;
assign n9590 = n12299 & n11023;
assign n6132 = n8738 | n28;
assign n798 = ~(n1853 ^ n1577);
assign n710 = ~(n2777 ^ n10319);
assign n8892 = ~(n4998 ^ n6646);
assign n10214 = ~(n82 ^ n3917);
assign n7895 = n1629 | n11103;
assign n4974 = n3461 | n8923;
assign n11781 = ~(n3471 ^ n355);
assign n9320 = ~(n504 ^ n8915);
assign n9824 = ~n2869;
assign n4687 = ~(n7144 ^ n4713);
assign n3053 = ~n3396;
assign n7424 = ~n12720;
assign n5778 = n264 | n3350;
assign n11647 = ~(n5882 | n786);
assign n11864 = n12853 | n9188;
assign n7731 = ~n7401;
assign n3716 = n12501 & n7631;
assign n4648 = ~n10167;
assign n6741 = n5466 & n4578;
assign n2220 = n876 | n11561;
assign n5330 = n375 | n11346;
assign n9251 = ~(n12632 ^ n2990);
assign n8870 = ~n7160;
assign n2261 = n4488 | n11502;
assign n1164 = ~n7252;
assign n11227 = ~(n6239 ^ n8808);
assign n5554 = n3587 | n2295;
assign n12219 = n1333 & n6038;
assign n10299 = ~(n7916 ^ n2642);
assign n12860 = ~(n6635 ^ n9193);
assign n12055 = ~(n11303 ^ n1614);
assign n3821 = n6849 | n10786;
assign n7198 = n8002 & n8934;
assign n9472 = n8390 | n2744;
assign n1069 = ~(n7756 ^ n4681);
assign n9230 = ~(n1260 ^ n1053);
assign n11383 = ~(n2073 ^ n8420);
assign n1154 = n2217 | n5086;
assign n11140 = ~(n5801 ^ n4160);
assign n10535 = n10938 | n5356;
assign n7252 = ~(n12268 ^ n4486);
assign n113 = n2033 & n8014;
assign n11839 = ~(n9324 | n12805);
assign n11454 = ~(n7083 ^ n12586);
assign n4089 = n3746 | n12816;
assign n3159 = ~(n8143 ^ n976);
assign n903 = n5940 & n6495;
assign n3437 = ~(n12387 ^ n4258);
assign n11642 = n12886 & n4117;
assign n8904 = ~(n5428 ^ n2647);
assign n2492 = ~(n8193 ^ n4752);
assign n7351 = ~n9059;
assign n7415 = ~(n2704 ^ n6163);
assign n5313 = ~(n11080 ^ n3441);
assign n11041 = n8377 & n5770;
assign n5750 = ~(n8736 ^ n6643);
assign n6678 = ~n3910;
assign n1214 = n5650 & n11675;
assign n9459 = n12841 & n6563;
assign n1259 = n4633 & n6062;
assign n2835 = ~(n2779 | n8001);
assign n10566 = ~(n2869 ^ n6292);
assign n8168 = ~(n10320 | n2747);
assign n5479 = ~n2100;
assign n2980 = n9370 | n12843;
assign n8771 = ~(n5023 | n4063);
assign n6756 = n2906 | n6213;
assign n2693 = ~(n9778 ^ n4240);
assign n10333 = n4469 & n1428;
assign n12938 = n9563 | n3881;
assign n340 = ~(n8795 ^ n12151);
assign n5277 = n9389 | n12328;
assign n1804 = ~(n5122 ^ n10977);
assign n4734 = n6770 & n2508;
assign n936 = n5177 & n10438;
assign n5534 = ~(n7684 ^ n12162);
assign n9560 = n673 & n7022;
assign n2310 = ~(n2502 ^ n11123);
assign n9680 = ~n6768;
assign n1625 = n10612 & n12938;
assign n4781 = n4212 & n4350;
assign n11868 = ~n4991;
assign n8578 = ~(n2945 ^ n5725);
assign n7046 = n9043 | n10840;
assign n5581 = ~(n2897 ^ n12421);
assign n11816 = n8583 | n12771;
assign n1241 = n994 | n10419;
assign n6385 = n9616 & n5262;
assign n8670 = n1239 & n5737;
assign n5510 = ~(n7563 | n9272);
assign n472 = ~(n2761 ^ n1190);
assign n220 = ~n3264;
assign n9641 = ~(n10728 ^ n8985);
assign n5297 = ~(n12717 ^ n10156);
assign n3923 = ~(n7310 ^ n11202);
assign n2405 = n10339 | n9188;
assign n12173 = n11259 | n6119;
assign n2531 = ~n12276;
assign n7777 = n752 | n10919;
assign n4379 = ~(n11957 ^ n7460);
assign n6071 = ~n503;
assign n992 = ~(n4977 ^ n104);
assign n7446 = ~(n11555 ^ n11609);
assign n3585 = n7839 | n6169;
assign n7041 = ~n7566;
assign n10040 = ~(n1810 | n10778);
assign n7913 = n4992 | n875;
assign n10788 = ~(n7215 ^ n4269);
assign n2027 = ~(n6567 ^ n11161);
assign n3394 = n4675 & n5818;
assign n5940 = n12467 | n918;
assign n3987 = ~(n9366 ^ n3063);
assign n4654 = ~n405;
assign n3090 = ~(n11221 ^ n3260);
assign n12666 = n4180 & n4990;
assign n8530 = ~n2342;
assign n12691 = n6718 | n1047;
assign n2339 = n12479 & n8174;
assign n11904 = ~(n10118 ^ n5601);
assign n10188 = ~n12637;
assign n11780 = ~(n11241 ^ n2062);
assign n8274 = n3127 | n11746;
assign n626 = ~(n12271 ^ n12707);
assign n4748 = ~(n1872 ^ n625);
assign n8710 = ~(n4239 | n5998);
assign n12366 = n7071 & n8338;
assign n10367 = n8870 | n10422;
assign n6944 = ~n9487;
assign n1747 = n349 | n3520;
assign n4180 = ~n9869;
assign n5178 = n4294 | n1120;
assign n10674 = n4263 | n8131;
assign n4447 = n5145 & n1247;
assign n10219 = ~(n9445 | n651);
assign n10925 = n6577 | n5012;
assign n1621 = n5038 & n2570;
assign n1117 = ~n3074;
assign n10341 = ~(n10380 ^ n4609);
assign n6033 = n11887 | n8740;
assign n9958 = ~n6039;
assign n10509 = n3322 | n9842;
assign n8695 = ~n8808;
assign n3004 = ~(n223 ^ n4172);
assign n4450 = n1599 & n11816;
assign n9340 = ~(n6952 ^ n4592);
assign n1731 = n3747 | n12249;
assign n7278 = ~(n7467 ^ n1063);
assign n11834 = ~(n812 ^ n11007);
assign n1388 = ~(n9261 | n9726);
assign n10092 = ~(n11234 | n12522);
assign n8016 = ~(n6612 ^ n3069);
assign n2957 = n11887 | n8655;
assign n4595 = n11980 & n3142;
assign n1851 = ~n12591;
assign n11498 = n5765 | n795;
assign n9701 = n11796 & n5093;
assign n1004 = ~n11208;
assign n7612 = n8026 | n3421;
assign n7566 = n6474 & n10755;
assign n10477 = n12 | n3805;
assign n7501 = ~(n5742 ^ n10360);
assign n10411 = n9365 | n3307;
assign n12114 = n8552 | n12535;
assign n3640 = n7038 & n6907;
assign n7373 = ~(n4576 | n7365);
assign n6730 = n4504 | n12036;
assign n4997 = ~(n3577 ^ n4372);
assign n12132 = n288 & n11386;
assign n11008 = n9693 | n8708;
assign n1807 = ~(n3626 ^ n5062);
assign n1256 = n1542 & n9639;
assign n2546 = ~(n9677 ^ n4331);
assign n8576 = n9370 | n11430;
assign n3117 = n6407 & n2208;
assign n506 = n6325 & n12504;
assign n11417 = n3746 | n10903;
assign n9500 = n321 & n3426;
assign n7468 = n989 | n7341;
assign n3610 = ~(n12047 ^ n4004);
assign n9392 = ~(n1959 ^ n5349);
assign n8561 = n10832 & n7421;
assign n8541 = ~n8712;
assign n1421 = n236 | n3770;
assign n6289 = ~(n3208 ^ n6757);
assign n3803 = ~n4004;
assign n5173 = ~n5522;
assign n7570 = ~(n2318 | n9475);
assign n1141 = ~(n2598 | n7576);
assign n8896 = n5530 | n5781;
assign n3684 = n8187 | n6402;
assign n6993 = n7449 | n9280;
assign n11091 = ~(n835 ^ n7979);
assign n7163 = ~(n4723 ^ n8905);
assign n7822 = n3467 | n11304;
assign n1243 = ~n833;
assign n1975 = n6306 & n12452;
assign n11475 = ~n1973;
assign n7416 = n3137 | n1711;
assign n4793 = ~n12286;
assign n832 = n3920 & n4934;
assign n4612 = n8738 | n4474;
assign n3696 = ~(n11971 ^ n10228);
assign n4822 = ~n3779;
assign n12202 = n10721 & n8976;
assign n5353 = n9560 & n12439;
assign n8742 = ~(n716 ^ n8670);
assign n7694 = n1941 | n995;
assign n11379 = ~n9851;
assign n21 = n12363 & n9142;
assign n3527 = n7801 | n6651;
assign n12117 = n10879 | n12843;
assign n3006 = n6364 & n8599;
assign n6710 = n9785 & n574;
assign n1456 = n8428 | n5538;
assign n12758 = n337 | n12329;
assign n10135 = n8583 | n3606;
assign n11646 = ~(n12054 ^ n2173);
assign n11166 = n3172 & n7456;
assign n4021 = ~(n11700 ^ n11456);
assign n8886 = ~(n5466 ^ n4578);
assign n956 = ~(n12918 ^ n4606);
assign n191 = ~n7862;
assign n2355 = ~(n12200 | n6975);
assign n12180 = n752 | n6084;
assign n1981 = n8506 | n2381;
assign n143 = n9250 & n10453;
assign n10876 = n12955 & n873;
assign n6369 = n5305 & n6038;
assign n7567 = n962 | n1047;
assign n10082 = ~n1187;
assign n12051 = n8055 | n3802;
assign n6439 = n2612 | n10166;
assign n2376 = ~(n9993 ^ n1281);
assign n12338 = ~(n2263 ^ n6568);
assign n10828 = ~(n2333 ^ n9209);
assign n7536 = n6560 & n3741;
assign n1970 = ~(n8663 | n5056);
assign n10544 = ~(n12544 ^ n9334);
assign n11568 = ~(n6708 ^ n7781);
assign n6758 = n6347 & n9890;
assign n5274 = n7982 & n7184;
assign n2780 = n4343 | n3224;
assign n8894 = n7391 | n4400;
assign n2652 = ~(n11120 ^ n280);
assign n3868 = ~n1520;
assign n9523 = n3746 | n9971;
assign n8887 = n10992 | n12749;
assign n1841 = ~n1511;
assign n10185 = n11671 | n7681;
assign n9205 = n10108 | n3911;
assign n4556 = n5374 & n3182;
assign n7012 = n3127 | n7703;
assign n2769 = ~n1156;
assign n760 = ~(n5000 ^ n3649);
assign n3205 = n989 | n10419;
assign n9879 = ~(n9909 | n5227);
assign n3239 = ~(n12023 ^ n7734);
assign n5208 = n619 & n8257;
assign n1224 = n6836 | n2004;
assign n8985 = ~(n899 ^ n4424);
assign n8478 = ~n479;
assign n10456 = ~(n363 ^ n7411);
assign n438 = n8428 | n6455;
assign n9294 = ~(n1695 ^ n276);
assign n7504 = n8026 | n9741;
assign n11211 = n3188 | n689;
assign n10361 = n10196 | n9144;
assign n3026 = n726 & n3800;
assign n1922 = n7449 | n4474;
assign n1598 = ~(n6201 ^ n1957);
assign n12149 = n6069 | n2586;
assign n1044 = n8583 | n1047;
assign n10450 = ~(n6361 ^ n4163);
assign n9985 = ~(n6598 ^ n10704);
assign n6917 = ~(n689 ^ n12152);
assign n8023 = ~(n841 ^ n7242);
assign n51 = n8127 | n1079;
assign n10358 = ~(n5646 | n3134);
assign n2280 = ~(n11142 ^ n10187);
assign n117 = ~n9923;
assign n6694 = ~(n5769 ^ n7239);
assign n8093 = n629 & n8432;
assign n4237 = n12237 | n9188;
assign n2294 = ~(n9390 ^ n9482);
assign n1518 = n834 & n5431;
assign n2447 = n5575 | n9741;
assign n5821 = ~(n9103 ^ n11114);
assign n12492 = ~(n8666 ^ n10557);
assign n2719 = ~n1624;
assign n5999 = n4366 & n10752;
assign n12283 = n6697 & n12225;
assign n1380 = n8183 | n4720;
assign n10065 = ~n774;
assign n9351 = n5945 | n6169;
assign n3181 = n1183 | n8109;
assign n5365 = n6570 & n11756;
assign n9295 = ~(n8243 | n2510);
assign n440 = n3796 & n5592;
assign n8683 = ~n4307;
assign n6308 = ~(n10056 ^ n9809);
assign n255 = n7116 | n10903;
assign n1507 = n9622 & n2782;
assign n9227 = ~(n3116 | n9931);
assign n11102 = n7116 | n11410;
assign n12918 = n8187 | n4400;
assign n11815 = ~(n2019 | n11218);
assign n4756 = ~(n38 ^ n6317);
assign n275 = n2367 | n4527;
assign n11413 = n4059 | n11827;
assign n5552 = ~(n10846 ^ n11890);
assign n5357 = n989 | n4775;
assign n1724 = n10108 | n4400;
assign n9206 = ~(n9442 ^ n12158);
assign n11254 = n4961 | n231;
assign n11637 = ~n4684;
assign n4136 = n4059 | n5497;
assign n10801 = n3632 | n2416;
assign n4457 = n8428 | n7558;
assign n6975 = ~(n1586 ^ n4236);
assign n745 = ~(n845 ^ n5325);
assign n11825 = n824 | n261;
assign n7977 = n10751 | n4114;
assign n10821 = ~(n4124 ^ n1342);
assign n11021 = ~(n6004 ^ n7204);
assign n1389 = ~(n7194 ^ n3514);
assign n10383 = n813 | n9865;
assign n1029 = ~(n3021 ^ n7548);
assign n698 = ~n5337;
assign n884 = n5501 & n4792;
assign n1385 = n8279 & n3861;
assign n2827 = n8336 & n6703;
assign n10436 = n1043 & n11532;
assign n2947 = n9878 | n3924;
assign n3002 = n1795 | n1748;
assign n1091 = n8269 & n5528;
assign n12251 = n7283 | n1162;
assign n4070 = n9441 & n7837;
assign n7596 = ~(n3829 ^ n8150);
assign n6167 = n10075 & n4837;
assign n8975 = ~(n6414 ^ n4749);
assign n1200 = ~n6535;
assign n9309 = n12429 | n6135;
assign n2873 = n11641 & n12379;
assign n12258 = ~(n7143 ^ n1997);
assign n6340 = ~n8564;
assign n8976 = n3215 | n2682;
assign n2812 = n6859 & n8559;
assign n1786 = ~(n1724 ^ n3122);
assign n1289 = ~(n2292 ^ n9276);
assign n4651 = n1421 & n1254;
assign n12469 = ~(n4167 ^ n5007);
assign n9430 = n3405 | n9833;
assign n2820 = ~(n10238 ^ n3850);
assign n1191 = ~(n10771 ^ n9904);
assign n6263 = ~(n10745 ^ n3082);
assign n161 = n5575 | n12899;
assign n12321 = n614 & n4443;
assign n4512 = n12361 | n11122;
assign n8484 = ~(n10 ^ n11277);
assign n10842 = n636 | n3924;
assign n9738 = n4324 & n1085;
assign n8226 = n7606 | n9822;
assign n1626 = ~(n12483 | n3830);
assign n8200 = ~(n8806 | n110);
assign n9975 = ~(n5709 | n886);
assign n8752 = n1937 | n6455;
assign n7676 = ~(n4439 ^ n9375);
assign n11213 = ~(n3762 ^ n9060);
assign n12634 = ~(n9648 ^ n5802);
assign n2863 = ~(n5607 | n7712);
assign n10401 = n6616 & n10578;
assign n8697 = n6265 | n8041;
assign n8186 = n11588 & n5476;
assign n4131 = ~(n2233 ^ n1184);
assign n8299 = n12853 | n530;
assign n3670 = ~n6948;
assign n1287 = n12237 | n4818;
assign n7926 = ~(n3116 ^ n4061);
assign n4249 = ~n1576;
assign n3772 = n6530 | n3167;
assign n3338 = n7994 | n7450;
assign n10079 = n8187 | n5497;
assign n4754 = n9510 | n11586;
assign n12352 = ~(n6268 | n2420);
assign n9716 = n8406 & n2607;
assign n11924 = ~n7097;
assign n6278 = n6066 & n5292;
assign n11206 = ~(n1012 ^ n5547);
assign n4400 = ~n11407;
assign n1703 = n11310 | n6964;
assign n12095 = ~(n5621 | n4075);
assign n10016 = ~(n8908 ^ n3736);
assign n9748 = n994 | n4242;
assign n3766 = n9748 | n10395;
assign n8277 = ~n9319;
assign n10335 = n10975 & n2152;
assign n9634 = n5279 | n12258;
assign n464 = n7396 & n5885;
assign n8071 = n2215 & n6729;
assign n12236 = ~n11545;
assign n3121 = ~(n11177 ^ n7836);
assign n505 = n12853 | n8655;
assign n5465 = n12742 | n11768;
assign n6663 = n5355 | n9397;
assign n6915 = ~(n4510 ^ n6410);
assign n6579 = n10142 | n7881;
assign n6302 = ~n12055;
assign n6064 = n11211 & n3438;
assign n1320 = n7083 & n672;
assign n10329 = n5279 & n12258;
assign n11807 = ~(n1542 ^ n5317);
assign n7944 = n5923 & n412;
assign n8785 = n10374 | n3898;
assign n12005 = ~(n9737 ^ n3263);
assign n6420 = ~(n1628 ^ n417);
assign n3061 = ~(n1312 ^ n2518);
assign n9103 = ~(n317 ^ n4065);
assign n4330 = ~(n3362 | n2178);
assign n10373 = ~n6086;
assign n6241 = n7133 | n2395;
assign n12650 = ~(n5899 ^ n3201);
assign n9621 = ~(n12865 ^ n6627);
assign n11084 = ~(n1371 | n6392);
assign n7392 = n1908 & n315;
assign n9519 = n3127 | n1546;
assign n8297 = ~n10535;
assign n2946 = n3603 | n2715;
assign n880 = ~n8719;
assign n11667 = ~(n8474 | n3774);
assign n3030 = n11026 | n12120;
assign n5483 = ~(n8668 ^ n2206);
assign n11641 = ~(n9405 ^ n1794);
assign n3079 = ~n7074;
assign n5916 = n1777 & n304;
assign n9478 = ~(n2535 ^ n11416);
assign n10697 = ~(n7612 ^ n10080);
assign n3681 = n11550 & n7051;
assign n1818 = ~(n1774 ^ n3777);
assign n4885 = n10656 | n7948;
assign n10164 = ~(n7396 ^ n1995);
assign n12310 = n3105 | n358;
assign n310 = ~n1979;
assign n7798 = n3742 & n390;
assign n12506 = n8049 & n12510;
assign n6919 = ~(n11879 | n11392);
assign n6148 = ~(n1608 ^ n9668);
assign n9086 = n8169 & n6633;
assign n1767 = ~(n1457 ^ n8297);
assign n4505 = ~(n4210 ^ n12769);
assign n7968 = ~n6289;
assign n3975 = ~(n8454 ^ n5734);
assign n2283 = ~(n12612 ^ n5537);
assign n12763 = ~(n7630 | n5736);
assign n9839 = ~(n6234 ^ n11982);
assign n1643 = ~n7454;
assign n10857 = n10902 & n1393;
assign n4144 = n9370 | n1738;
assign n9155 = n11026 | n7506;
assign n10855 = n11076 | n7067;
assign n5018 = ~n5976;
assign n3867 = ~n3858;
assign n7834 = ~n11289;
assign n6426 = n10835 | n8830;
assign n5033 = ~(n9054 ^ n1187);
assign n489 = ~(n5542 | n7234);
assign n7353 = ~(n3510 | n7366);
assign n5909 = n4134 & n1943;
assign n3882 = ~(n9429 | n7092);
assign n11143 = ~(n6246 ^ n10345);
assign n1719 = n12853 | n4913;
assign n8797 = n5730 & n10407;
assign n1511 = n11474 | n9371;
assign n1028 = ~(n11335 | n6518);
assign n9269 = n12867 & n3434;
assign n9011 = ~(n8682 | n1525);
assign n4107 = n1183 | n1932;
assign n4557 = ~n3776;
assign n10121 = n11682 | n12092;
assign n4663 = ~(n4716 ^ n7053);
assign n10572 = n5066 | n3226;
assign n9864 = ~(n1074 | n5426);
assign n11978 = ~n3877;
assign n10967 = ~(n5491 ^ n3664);
assign n7054 = n10108 | n10066;
assign n11443 = n5530 | n8259;
assign n3717 = ~n3565;
assign n8948 = ~(n6122 ^ n189);
assign n504 = n11958 | n3356;
assign n11055 = n7862 & n2879;
assign n4159 = ~(n4766 ^ n3635);
assign n5295 = ~(n7251 ^ n4264);
assign n1552 = ~(n10046 ^ n6927);
assign n7228 = n10104 | n10498;
assign n5287 = n10269 | n3308;
assign n12832 = ~(n905 | n11505);
assign n6372 = ~(n9708 ^ n4822);
assign n9352 = ~n4948;
assign n11651 = ~(n1611 ^ n11337);
assign n6885 = ~n11373;
assign n2370 = ~(n2244 ^ n5697);
assign n1897 = n11890 | n4291;
assign n7400 = n12361 | n3468;
assign n5585 = n5889 | n802;
assign n3895 = n752 | n1413;
assign n8734 = ~(n8124 ^ n3270);
assign n5747 = n12565 | n903;
assign n12358 = ~(n3988 ^ n11105);
assign n11265 = n8738 | n795;
assign n5835 = ~(n1017 | n4853);
assign n3257 = n8336 & n7500;
assign n2267 = n11254 & n7847;
assign n12140 = ~(n11462 ^ n5398);
assign n5577 = n10641 & n3867;
assign n6079 = ~(n11451 ^ n6853);
assign n4564 = n7495 | n12843;
assign n455 = n8752 | n1918;
assign n10350 = ~n2365;
assign n5419 = ~n7304;
assign n4029 = n4380 | n5245;
assign n5795 = ~(n12671 ^ n1615);
assign n12151 = n12136 | n9779;
assign n12374 = ~(n9745 ^ n3112);
assign n12456 = n12503 | n4875;
assign n11551 = n12774 | n2423;
assign n9936 = ~(n6367 | n987);
assign n2779 = ~(n4301 | n2204);
assign n12652 = n12839 & n1279;
assign n12731 = n11754 | n3073;
assign n10513 = n6373 | n8285;
assign n8089 = n7756 & n4681;
assign n11552 = ~n5767;
assign n7616 = ~(n9035 ^ n4616);
assign n11395 = ~(n11720 ^ n11089);
assign n9863 = ~(n9247 ^ n9033);
assign n2967 = ~(n1612 | n4673);
assign n2772 = n12245 | n300;
assign n2293 = n11928 | n11308;
assign n11294 = ~n7658;
assign n6780 = n8854 | n1035;
assign n6046 = n12739 & n3108;
assign n4951 = ~(n5463 | n12693);
assign n718 = n7074 & n4105;
assign n1842 = n6625 | n12959;
assign n12429 = n7176 & n506;
assign n5438 = n3127 | n1851;
assign n8371 = ~n391;
assign n11312 = ~(n3416 ^ n4687);
assign n6036 = ~n7796;
assign n1720 = ~n12693;
assign n12933 = n7173 | n8125;
assign n8824 = ~(n3405 ^ n10106);
assign n11494 = ~n6338;
assign n2438 = ~(n1124 ^ n8110);
assign n5959 = n5355 | n510;
assign n2579 = ~n11267;
assign n1614 = ~(n10735 ^ n4091);
assign n5309 = ~(n3628 ^ n894);
assign n8989 = ~(n862 ^ n2668);
assign n5366 = n1941 | n2815;
assign n10718 = n12214 & n4423;
assign n11624 = n6718 | n9521;
assign n8620 = n12009 | n788;
assign n12162 = ~(n5749 ^ n8809);
assign n11492 = n8294 & n6316;
assign n5403 = ~(n1412 ^ n12957);
assign n4462 = ~(n11824 ^ n1545);
assign n10094 = n754 | n624;
assign n3931 = ~(n10215 ^ n4848);
assign n6137 = n191 | n9589;
assign n6319 = n6003 & n11614;
assign n4619 = ~(n5758 ^ n8210);
assign n8995 = ~(n8972 ^ n2667);
assign n9410 = n11879 & n11392;
assign n2965 = ~(n11532 ^ n1195);
assign n8327 = n343 | n7278;
assign n3568 = ~(n11053 ^ n5745);
assign n8022 = ~(n1803 ^ n6421);
assign n9358 = ~(n11723 ^ n8487);
assign n1229 = n10545 & n7733;
assign n9218 = ~n669;
assign n3811 = ~(n1707 ^ n700);
assign n8624 = ~n1132;
assign n4071 = n10698 & n7208;
assign n11934 = n12814 & n8431;
assign n12621 = ~n1410;
assign n10109 = n10714 | n43;
assign n2898 = ~n860;
assign n3015 = n5575 | n6084;
assign n7062 = ~(n1569 ^ n7211);
assign n3969 = ~(n11042 | n6350);
assign n3033 = n9286 | n2889;
assign n12370 = n12393 | n1463;
assign n11835 = ~(n6097 ^ n4496);
assign n4446 = n11923 | n1476;
assign n649 = n191 | n10066;
assign n11065 = n1699 | n12754;
assign n3829 = n9003 & n7006;
assign n8123 = n2099 | n2259;
assign n11259 = n8870 | n12080;
assign n4723 = n8870 | n9586;
assign n4407 = n6720 & n7516;
assign n9095 = ~(n656 ^ n3516);
assign n3400 = ~(n2183 | n5920);
assign n7901 = n1230 & n811;
assign n388 = ~n3646;
assign n173 = n11222 & n10848;
assign n1438 = n3127 | n3911;
assign n7866 = ~(n3055 ^ n10950);
assign n11260 = ~(n5632 ^ n6483);
assign n3884 = ~n9858;
assign n10863 = ~(n6543 ^ n5480);
assign n2853 = n8552 | n8740;
assign n9315 = ~n11499;
assign n5535 = ~(n9748 ^ n10395);
assign n1010 = ~(n11088 ^ n9952);
assign n11629 = ~(n10658 ^ n10946);
assign n4776 = ~(n6423 ^ n1125);
assign n8938 = ~(n4446 ^ n6647);
assign n1848 = n7564 | n1363;
assign n5020 = n6470 | n7392;
assign n6548 = n11691 & n8511;
assign n2570 = n4831 & n426;
assign n10447 = ~(n7762 | n8302);
assign n1451 = n3926 & n10474;
assign n11883 = n3088 | n8080;
assign n4334 = ~(n2111 ^ n7631);
assign n5087 = n10142 | n5851;
assign n1532 = n9652 & n9798;
assign n1349 = n9621 & n1490;
assign n3199 = ~n10191;
assign n10379 = n8738 | n9144;
assign n916 = ~n12553;
assign n2139 = ~n1451;
assign n6883 = n6741 | n3136;
assign n6739 = n6426 & n11009;
assign n8909 = ~n4883;
assign n3080 = ~n7977;
assign n66 = ~(n12263 ^ n3569);
assign n6888 = n7322 | n256;
assign n12035 = ~(n9117 ^ n3266);
assign n7710 = ~n3804;
assign n10177 = ~(n1923 | n6640);
assign n2122 = ~n8356;
assign n2788 = n5413 & n10170;
assign n1186 = n7151 | n7714;
assign n601 = ~(n7488 ^ n8876);
assign n5390 = ~(n6686 ^ n7599);
assign n3755 = n6644 | n2461;
assign n4244 = n8026 | n184;
assign n6382 = ~n1324;
assign n9236 = n12614 & n1022;
assign n8736 = n5575 | n9971;
assign n4920 = n10835 | n9521;
assign n6961 = ~(n4076 ^ n10213);
assign n9543 = n6868 | n793;
assign n12385 = ~n2350;
assign n7225 = ~(n9336 | n11463);
assign n6680 = n12223 & n7114;
assign n12019 = n12183 | n10177;
assign n6850 = ~(n2664 | n7797);
assign n6147 = n4387 | n4162;
assign n5720 = ~(n6110 ^ n4199);
assign n11480 = n9836 & n8081;
assign n5371 = n7495 | n10066;
assign n3283 = ~(n4322 ^ n512);
assign n6386 = n10744 | n2240;
assign n5378 = n1003 | n6517;
assign n1499 = ~(n9752 ^ n7238);
assign n9 = ~(n12538 | n10690);
assign n544 = ~(n2249 ^ n9983);
assign n4353 = ~(n11356 ^ n5342);
assign n12686 = ~n7610;
assign n3736 = n8959 | n3421;
assign n9021 = n10018 & n10021;
assign n11430 = ~n12000;
assign n1263 = n1679 & n10359;
assign n6979 = n289 | n11772;
assign n805 = n9335 & n11031;
assign n9823 = ~(n10195 | n3161);
assign n235 = ~(n4121 ^ n11975);
assign n11386 = n8583 | n1509;
assign n4701 = ~(n8030 ^ n8060);
assign n8727 = n9504 | n11910;
assign n7293 = ~n5898;
assign n9347 = n12218 & n2632;
assign n3228 = ~(n6624 | n10834);
assign n3515 = ~(n5577 ^ n3204);
assign n4576 = n5530 | n12124;
assign n2183 = n10004 ^ n6289;
assign n6821 = ~(n6461 ^ n3211);
assign n12584 = n81 & n12343;
assign n1898 = n2003 & n12762;
assign n7748 = n4059 | n2358;
assign n12761 = n989 | n5851;
assign n3105 = n12361 | n9741;
assign n7595 = ~(n12114 ^ n944);
assign n11470 = n4120 | n2805;
assign n4270 = ~(n9757 ^ n5806);
assign n4129 = n7941 | n9113;
assign n7164 = ~(n5981 ^ n282);
assign n6164 = n1073 & n6790;
assign n10770 = n5860 & n10848;
assign n3808 = ~n7405;
assign n12567 = n2286 | n7581;
assign n5736 = n7544 & n7228;
assign n11944 = ~n12811;
assign n8959 = ~n7436;
assign n1466 = ~(n1486 ^ n4221);
assign n7178 = n6698 & n2158;
assign n4172 = ~(n1330 ^ n106);
assign n486 = ~n10023;
assign n4161 = n10750 | n12883;
assign n1959 = ~(n12887 | n539);
assign n9555 = ~(n11284 ^ n5626);
assign n8482 = ~(n3065 ^ n7032);
assign n7175 = ~(n8776 ^ n123);
assign n8404 = n3096 | n11896;
assign n10354 = n12119 | n7928;
assign n12054 = ~(n10809 ^ n11107);
assign n11162 = n6681 | n10894;
assign n11219 = ~(n815 ^ n11075);
assign n1372 = n5066 & n3226;
assign n9318 = n3664 | n6712;
assign n4709 = ~(n2215 ^ n6729);
assign n3058 = ~n4838;
assign n12014 = ~(n2805 ^ n5521);
assign n10991 = ~(n1361 | n8577);
assign n6654 = n8870 | n7382;
assign n2689 = ~n1479;
assign n8165 = n23 & n7844;
assign n825 = ~(n11745 | n2578);
assign n3229 = ~n5819;
assign n3391 = ~(n9281 ^ n8563);
assign n1971 = ~(n7713 ^ n9343);
assign n4964 = n10975 | n2152;
assign n4674 = ~n4499;
assign n7818 = ~(n705 ^ n8192);
assign n10480 = n12361 | n6169;
assign n3354 = ~(n933 ^ n12666);
assign n9932 = ~(n6222 ^ n9902);
assign n4802 = ~n1880;
assign n2565 = ~(n396 ^ n8802);
assign n8408 = ~(n11489 ^ n1403);
assign n7943 = ~n12700;
assign n9169 = n1128 & n6110;
assign n7482 = ~(n2382 ^ n6633);
assign n8090 = ~n8799;
assign n7887 = ~(n3804 ^ n3531);
assign n4676 = n8738 | n3606;
assign n11721 = ~(n3327 | n11046);
assign n10982 = ~n12003;
assign n243 = n6146 | n6749;
assign n12856 = n9370 | n1455;
assign n11547 = n10157 | n8643;
assign n2790 = ~n5888;
assign n2922 = n7012 & n2026;
assign n10957 = n9193 | n6351;
assign n12097 = ~(n3209 ^ n8681);
assign n78 = n5530 | n12080;
assign n12733 = n11222 & n405;
assign n770 = n6348 | n10175;
assign n1053 = n11719 | n12843;
assign n9536 = ~n10734;
assign n3689 = ~(n3966 ^ n11977);
assign n1266 = n6577 | n2815;
assign n12693 = n508 & n8530;
assign n1712 = ~(n4542 ^ n5403);
assign n8569 = n12127 & n3081;
assign n10773 = ~n8900;
assign n7766 = ~(n1787 ^ n7591);
assign n11249 = n1539 | n1455;
assign n4206 = n7283 | n7424;
assign n2296 = ~(n8353 ^ n1922);
assign n7108 = n6650 | n5386;
assign n10359 = ~(n3182 ^ n4082);
assign n8098 = n6111 | n212;
assign n1485 = ~(n10313 ^ n6603);
assign n10910 = ~n82;
assign n7465 = n8026 | n11775;
assign n1736 = n646 & n494;
assign n7370 = n4204 | n5028;
assign n6023 = ~(n12884 ^ n4139);
assign n8847 = n12119 | n2964;
assign n5462 = ~n3284;
assign n6291 = n4811 & n8090;
assign n8138 = ~(n8460 ^ n5610);
assign n5533 = ~(n11935 ^ n10821);
assign n8659 = n4059 | n4775;
assign n9510 = n4498 | n11827;
assign n11292 = ~n3206;
assign n9335 = ~n11188;
assign n5831 = ~(n8704 ^ n11689);
assign n10808 = n12853 | n7928;
assign n3682 = ~n5284;
assign n5880 = n8587 & n10206;
assign n6702 = ~(n8320 ^ n6588);
assign n2804 = ~n742;
assign n9947 = ~(n9620 ^ n9238);
assign n2932 = ~(n1356 ^ n10540);
assign n6533 = ~(n11997 ^ n930);
assign n8680 = ~(n6073 ^ n8947);
assign n5350 = n11841 & n3002;
assign n10974 = n4628 | n12535;
assign n8945 = n1051 | n9741;
assign n4686 = n1027 ^ n3950;
assign n10157 = ~n3992;
assign n7029 = ~(n10878 | n5623);
assign n10559 = ~(n2397 ^ n12403);
assign n10587 = n8552 | n7382;
assign n6701 = n11445 | n247;
assign n985 = ~(n1266 ^ n6324);
assign n2672 = n8552 | n8109;
assign n7426 = ~(n5263 ^ n3657);
assign n365 = n1699 | n10854;
assign n10403 = n1594 & n10964;
assign n5486 = n8583 | n9521;
assign n4445 = ~(n3988 | n5039);
assign n8237 = n10118 & n5887;
assign n1854 = n11226 | n2658;
assign n3356 = ~n8236;
assign n1319 = ~(n4718 | n3634);
assign n4278 = ~(n7643 | n913);
assign n7275 = n637 & n5996;
assign n8878 = n10434 & n9894;
assign n6024 = n197 & n8330;
assign n6398 = n3713 | n3227;
assign n1323 = ~(n6865 | n9059);
assign n11119 = ~n6353;
assign n6117 = n1856 | n3748;
assign n6581 = n8354 | n6513;
assign n1177 = ~(n12471 ^ n535);
assign n11035 = ~(n12524 | n8898);
assign n7067 = n762 & n6312;
assign n7301 = n2251 & n4277;
assign n2196 = ~(n7897 | n4918);
assign n3124 = ~(n12267 ^ n7399);
assign n9753 = n9279 & n10331;
assign n5844 = n11182 | n4200;
assign n600 = ~(n3906 ^ n11203);
assign n7222 = ~(n1536 ^ n12651);
assign n11284 = ~(n1347 ^ n7216);
assign n5517 = ~(n9467 ^ n9312);
assign n4856 = n5575 | n8768;
assign n1639 = n8428 | n12816;
assign n4348 = ~n707;
assign n8844 = n2226 & n2522;
assign n9586 = ~n11967;
assign n10711 = ~(n10724 ^ n10581);
assign n9887 = n6977 | n9741;
assign n4919 = n2930 & n4901;
assign n5251 = n636 | n3224;
assign n2707 = n12263 & n9203;
assign n10705 = ~(n582 ^ n11014);
assign n2796 = ~(n3976 ^ n10429);
assign n8211 = ~n7277;
assign n6182 = ~n1082;
assign n2320 = ~(n4191 ^ n6555);
assign n10693 = ~(n3396 ^ n12700);
assign n10606 = ~n10171;
assign n12088 = ~(n6894 | n7105);
assign n12628 = n1842 & n10943;
assign n12058 = ~(n6514 ^ n5373);
assign n11246 = ~(n4597 ^ n394);
assign n458 = ~(n1873 ^ n11223);
assign n8751 = n10835 | n1739;
assign n1428 = ~(n2274 ^ n11858);
assign n6226 = n7243 & n2460;
assign n3869 = ~(n8097 ^ n4520);
assign n10192 = ~(n3888 ^ n10029);
assign n12689 = n116 & n5826;
assign n7540 = n9656 & n12411;
assign n10259 = n1951 & n11244;
assign n5099 = ~(n9461 | n6363);
assign n9962 = ~(n5963 | n4102);
assign n112 = n9321 ^ n3824;
assign n12943 = ~(n8545 ^ n4824);
assign n11973 = n9389 | n11430;
assign n4469 = ~(n1949 ^ n12487);
assign n9405 = ~(n8949 ^ n6724);
assign n11263 = n8322 & n6737;
assign n12887 = ~(n6751 | n3519);
assign n1112 = n1051 | n7425;
assign n4675 = n2613 | n3826;
assign n1118 = ~(n4001 ^ n592);
assign n2398 = n4628 | n6513;
assign n5304 = ~(n6728 ^ n3827);
assign n6938 = ~(n2991 ^ n8769);
assign n540 = ~(n2561 | n6572);
assign n3100 = ~(n9230 ^ n8689);
assign n6834 = ~(n4437 ^ n5220);
assign n1379 = ~(n1127 | n11848);
assign n482 = n10697 & n4968;
assign n9613 = ~(n3792 ^ n1244);
assign n5555 = ~(n7009 ^ n7664);
assign n12912 = n11887 | n12080;
assign n6520 = ~(n5334 ^ n4884);
assign n11804 = ~(n5335 | n9207);
assign n3046 = ~(n11960 ^ n3273);
assign n2414 = n3145 | n1267;
assign n2584 = ~(n7983 ^ n2334);
assign n5109 = ~(n4315 ^ n8832);
assign n6037 = ~(n10203 | n7219);
assign n8840 = ~(n5988 ^ n6856);
assign n6341 = ~(n6874 | n10455);
assign n2146 = ~(n8635 ^ n2698);
assign n8942 = ~(n35 ^ n9110);
assign n9502 = ~(n9432 ^ n7226);
assign n7781 = ~(n8319 ^ n8044);
assign n2445 = ~n5371;
assign n11216 = ~(n7230 ^ n9154);
assign n10247 = ~(n8092 | n5459);
assign n12111 = ~(n7708 ^ n2758);
assign n4384 = n1288 | n2868;
assign n10486 = n2854 & n1961;
assign n9210 = ~n292;
assign n9622 = n11228 | n8573;
assign n6560 = n5765 | n4642;
assign n4024 = ~(n3928 ^ n9075);
assign n5859 = ~(n8254 ^ n6490);
assign n4058 = ~(n2975 ^ n10901);
assign n1468 = ~(n3329 | n9053);
assign n2861 = n7965 & n9763;
assign n4538 = ~(n10048 ^ n9129);
assign n9643 = ~(n3954 | n8955);
assign n10727 = n346 | n7721;
assign n11905 = n1937 | n7876;
assign n8946 = n60 | n11213;
assign n1267 = n8428 | n5012;
assign n2893 = n5355 | n7341;
assign n5986 = ~(n12870 | n10107);
assign n3617 = ~n1199;
assign n4994 = n994 | n7341;
assign n2874 = n5575 | n8414;
assign n2134 = ~n6946;
assign n1566 = n10010 | n10815;
assign n2436 = n8900 & n5531;
assign n5639 = ~(n3653 ^ n2021);
assign n7552 = n11317 & n1265;
assign n8102 = n10464 & n4164;
assign n1305 = n2064 | n5122;
assign n11133 = n2619 | n4978;
assign n3785 = ~(n4256 ^ n5534);
assign n5006 = ~n8765;
assign n1024 = n12119 | n1163;
assign n6455 = ~n3719;
assign n2716 = ~n8275;
assign n5589 = n10835 | n4642;
assign n12090 = n3715 | n9788;
assign n1695 = n9370 | n7881;
assign n8981 = n5059 | n11994;
assign n7008 = ~(n110 ^ n2882);
assign n269 = ~n9581;
assign n8991 = n2850 | n9469;
assign n11732 = n2408 & n1931;
assign n10210 = n4778 | n7382;
assign n12857 = ~(n9907 | n9927);
assign n8621 = ~(n6085 ^ n4762);
assign n5997 = ~(n7037 ^ n8613);
assign n9196 = n8187 | n3911;
assign n7417 = ~(n6165 | n8787);
assign n7039 = ~(n10877 ^ n4406);
assign n1531 = n7195 & n7793;
assign n230 = ~(n7457 ^ n9017);
assign n10724 = ~(n11537 ^ n11206);
assign n8883 = ~(n8750 | n10537);
assign n4941 = n7503 | n11066;
assign n5121 = ~n5590;
assign n5117 = ~(n5969 ^ n11591);
assign n7509 = n6577 | n6455;
assign n7121 = n5765 | n1476;
assign n5732 = n191 | n1455;
assign n12508 = ~(n12059 ^ n2796);
assign n1900 = n6131 & n2060;
assign n12680 = n8406 | n2607;
assign n2060 = n3486 & n7825;
assign n8953 = ~(n12761 ^ n50);
assign n3731 = ~(n10435 ^ n4895);
assign n9412 = ~(n8750 ^ n6167);
assign n5156 = ~n8289;
assign n11777 = n9138 & n2135;
assign n265 = ~n7576;
assign n2162 = n5765 | n7921;
assign n2732 = n7149 | n9026;
assign n8050 = n12385 & n12353;
assign n12326 = n4500 & n1483;
assign n3763 = ~(n9814 | n9609);
assign n3321 = n6650 & n5386;
assign n11169 = n1899 | n5376;
assign n101 = n1197 | n4827;
assign n12238 = ~(n2227 | n9716);
assign n10542 = n8496 | n4583;
assign n1047 = ~n1980;
assign n1102 = n2363 | n229;
assign n12491 = ~(n10346 | n7372);
assign n8603 = n5077 & n12350;
assign n10382 = ~n5029;
assign n3597 = ~n11953;
assign n7634 = ~n3881;
assign n4254 = n11958 | n5311;
assign n10654 = ~(n5569 ^ n1877);
assign n3450 = ~(n9108 ^ n3983);
assign n1175 = ~n11198;
assign n830 = n6090 | n2811;
assign n2806 = n9231 & n6051;
assign n12603 = ~n11685;
assign n1575 = ~n4492;
assign n5453 = n2217 | n3599;
assign n9739 = n4805 & n1564;
assign n5948 = n8026 | n11410;
assign n8470 = ~n9842;
assign n1146 = n9797 & n2900;
assign n3898 = ~(n1037 ^ n2402);
assign n10806 = n11239 | n5980;
assign n6128 = ~n5673;
assign n9792 = ~(n7827 ^ n711);
assign n4289 = n752 | n3468;
assign n3678 = n11923 | n609;
assign n10081 = n5995 & n769;
assign n3630 = ~(n8817 | n4099);
assign n7259 = ~(n9655 ^ n865);
assign n2326 = n7449 | n3606;
assign n170 = ~(n12492 ^ n425);
assign n4305 = ~n3257;
assign n4973 = ~n3428;
assign n3676 = ~(n12104 ^ n11215);
assign n7334 = n4059 | n6389;
assign n9726 = ~n2440;
assign n7114 = n9389 | n8524;
assign n1941 = ~n4187;
assign n3619 = n12052 & n9818;
assign n1218 = ~(n2268 ^ n7047);
assign n11234 = n11552 | n9144;
assign n7560 = ~n131;
assign n11998 = n6577 | n2232;
assign n8979 = ~(n10730 ^ n4507);
assign n8375 = ~n267;
assign n628 = n3097 | n7281;
assign n2375 = ~(n6326 ^ n6631);
assign n4900 = n1814 & n739;
assign n3280 = ~n5405;
assign n8729 = n9976 | n1638;
assign n9000 = n10835 | n3606;
assign n4010 = n2562 & n5484;
assign n48 = ~(n11025 ^ n6958);
assign n9908 = n2213 | n1443;
assign n8256 = n973 | n12170;
assign n12048 = ~(n12879 ^ n10887);
assign n5911 = ~(n54 ^ n11751);
assign n7680 = n250 ^ n11151;
assign n10599 = ~(n10018 ^ n10021);
assign n7205 = n1471 & n8028;
assign n9367 = n7268 & n1767;
assign n11252 = n9141 & n5149;
assign n10827 = ~n7233;
assign n449 = n10532 & n7374;
assign n1232 = n8538 & n1504;
assign n6244 = n11552 | n3606;
assign n8919 = n5577 & n7816;
assign n8971 = ~(n4561 ^ n10280);
assign n12239 = ~(n12775 ^ n12157);
assign n5133 = ~(n7605 ^ n3031);
assign n6631 = n9182 & n6245;
assign n10309 = n3743 | n8830;
assign n12435 = n1708 & n12114;
assign n11621 = n6413 | n166;
assign n6742 = n3166 ^ n3894;
assign n6600 = ~(n12129 | n12573);
assign n3038 = n9370 | n11827;
assign n10567 = ~(n3543 ^ n4861);
assign n1166 = n11433 | n12816;
assign n9283 = ~(n2817 ^ n12589);
assign n6436 = ~(n12370 ^ n10650);
assign n1943 = n2118 | n1155;
assign n169 = ~(n11073 ^ n10424);
assign n3075 = ~(n8054 ^ n9338);
assign n385 = n5038 | n2570;
assign n1996 = ~n7035;
assign n1137 = n1233 | n6330;
assign n10220 = n2536 & n12112;
assign n5505 = n2067 | n12568;
assign n10481 = ~(n7332 ^ n6932);
assign n9308 = n10142 | n2358;
assign n12350 = n3874 | n6060;
assign n7128 = n6055 | n6997;
assign n11293 = n705 | n1310;
assign n6868 = ~(n9692 | n4439);
assign n2046 = ~n1104;
assign n2243 = n10390 | n10883;
assign n10364 = ~n12949;
assign n10417 = ~(n267 ^ n3548);
assign n9388 = ~(n1630 ^ n2046);
assign n305 = n6977 | n7952;
assign n12607 = ~(n6993 | n9915);
assign n4235 = ~(n8945 | n1859);
assign n11382 = n6080 | n2953;
assign n10005 = ~(n6872 ^ n7751);
assign n11441 = ~(n4728 ^ n12275);
assign n11879 = n3743 | n6922;
assign n11531 = n2593 & n8497;
assign n3998 = ~n2209;
assign n8828 = ~(n978 ^ n977);
assign n4118 = ~(n3372 ^ n5322);
assign n4367 = n8521 ^ n10445;
assign n3572 = ~(n3302 ^ n3771);
assign n7376 = n11958 | n3903;
assign n11897 = ~(n6722 ^ n8318);
assign n5988 = n3617 | n826;
assign n5328 = ~n9606;
assign n9793 = n215 | n939;
assign n7779 = ~(n2788 ^ n12627);
assign n2556 = n9584 | n9521;
assign n4627 = n12091 | n2348;
assign n3871 = ~(n11444 ^ n439);
assign n6469 = ~(n1646 ^ n11022);
assign n3164 = ~(n12421 | n10063);
assign n11888 = ~(n12610 ^ n10283);
assign n9326 = n2099 | n12535;
assign n12183 = ~(n10100 | n9839);
assign n351 = ~n400;
assign n11860 = ~n3797;
assign n5537 = n3746 | n12899;
assign n2603 = n6027 & n2250;
assign n9077 = ~n12952;
assign n3702 = ~(n7491 | n10470);
assign n3271 = n10663 | n8937;
assign n11290 = n6939 | n208;
assign n11974 = n8203 | n10722;
assign n9750 = ~(n7667 | n9348);
assign n7162 = ~(n3404 ^ n12828);
assign n3374 = n1699 | n530;
assign n8353 = n10835 | n12771;
assign n3032 = n9048 | n5993;
assign n12854 = ~(n2729 ^ n647);
assign n6053 = n5530 | n7928;
assign n11373 = ~(n9084 ^ n9478);
assign n4303 = n4059 | n1162;
assign n2341 = ~(n3376 | n12134);
assign n3135 = ~(n7542 | n12896);
assign n4498 = ~n5240;
assign n4894 = n5779 & n10102;
assign n473 = n5674 & n11330;
assign n12230 = ~(n7493 ^ n8075);
assign n10939 = ~n3424;
assign n10269 = n7116 | n2815;
assign n9306 = n2292 | n662;
assign n4395 = ~(n5364 ^ n12595);
assign n588 = n6718 | n8643;
assign n12859 = ~n4325;
assign n10830 = n5967 & n3028;
assign n9444 = n994 | n1455;
assign n4474 = ~n9763;
assign n7948 = n5441 & n1862;
assign n6017 = ~(n3577 | n46);
assign n7654 = n12310 & n9430;
assign n1121 = n3133 & n10313;
assign n10561 = ~n3769;
assign n6964 = ~(n8547 ^ n4020);
assign n6401 = ~(n7779 | n10248);
assign n3903 = ~n6126;
assign n10303 = ~(n12436 ^ n12389);
assign n12635 = ~(n7170 | n9038);
assign n9935 = ~(n1537 | n8188);
assign n2037 = n7313 | n3640;
assign n10651 = ~(n10423 ^ n4517);
assign n8441 = n2686 | n10618;
assign n11273 = n8545 & n12783;
assign n3924 = ~n8665;
assign n819 = n11744 & n2222;
assign n1472 = n10761 & n3234;
assign n7629 = n3984 | n3902;
assign n4014 = ~n2106;
assign n3220 = n5116 | n11361;
assign n3470 = n4299 & n5698;
assign n3122 = ~(n7620 ^ n1181);
assign n3658 = ~n6631;
assign n8826 = ~(n3221 | n3314);
assign n11957 = ~(n9162 ^ n7106);
assign n2733 = n12818 | n541;
assign n10266 = n5138 | n8471;
assign n6084 = ~n8065;
assign n9607 = ~n4659;
assign n2316 = ~(n11439 ^ n1609);
assign n3471 = ~(n7335 ^ n8466);
assign n12944 = ~(n4246 ^ n4265);
assign n6165 = n8451 & n5430;
assign n1264 = n12079 & n1704;
assign n8225 = n5515 & n6683;
assign n9286 = ~(n10560 | n5029);
assign n11 = n4628 | n8259;
assign n10785 = ~(n9844 ^ n9225);
assign n357 = n7283 | n7341;
assign n592 = n9990 & n2840;
assign n495 = ~(n602 ^ n10024);
assign n2458 = ~(n10289 ^ n6679);
assign n633 = n9554 | n8507;
assign n3049 = ~(n12008 ^ n5555);
assign n209 = ~n7936;
assign n833 = ~(n3220 ^ n5675);
assign n10442 = ~n2826;
assign n1986 = ~(n5571 ^ n537);
assign n57 = ~(n2950 ^ n7252);
assign n3673 = n1623 & n7323;
assign n9541 = n9370 | n1546;
assign n5416 = n6256 | n7489;
assign n5815 = n9107 & n2986;
assign n10729 = ~n4468;
assign n18 = ~(n4514 | n9659);
assign n11832 = n10945 | n7318;
assign n3563 = ~(n5101 | n9206);
assign n7210 = ~(n8273 ^ n4909);
assign n2319 = n2217 | n6922;
assign n7088 = n8870 | n6513;
assign n10012 = n9170 | n6389;
assign n11769 = n1075 | n8013;
assign n4151 = ~(n6050 ^ n3424);
assign n5368 = n309 & n8529;
assign n7042 = ~(n11443 ^ n11237);
assign n5031 = n6718 | n28;
assign n3760 = ~n3001;
assign n12527 = n636 | n8109;
assign n10699 = ~(n3428 ^ n1166);
assign n1794 = ~n11154;
assign n6190 = ~(n832 | n3178);
assign n2684 = n4332 & n9232;
assign n10199 = n5530 | n4818;
assign n12866 = ~(n8045 ^ n7557);
assign n929 = n8127 | n12843;
assign n8658 = ~(n5415 ^ n4248);
assign n2179 = ~(n9064 | n3185);
assign n1581 = n3976 | n12059;
assign n6711 = ~(n5733 ^ n1237);
assign n4636 = ~n313;
assign n8280 = ~n8281;
assign n2921 = n6948 | n8357;
assign n10805 = n11061 | n9759;
assign n1527 = ~(n6151 | n11219);
assign n6141 = ~n6330;
assign n5424 = n7273 & n5985;
assign n11792 = n6072 & n891;
assign n5938 = n3042 | n2965;
assign n6646 = ~(n5865 ^ n8480);
assign n276 = n3127 | n5497;
assign n9575 = ~(n1215 ^ n5055);
assign n9456 = ~(n6516 ^ n9533);
assign n2491 = n582 | n11014;
assign n715 = ~(n12912 ^ n8916);
assign n4372 = ~(n10776 ^ n4809);
assign n3078 = n989 | n2358;
assign n6660 = n8187 | n1546;
assign n5358 = ~(n4917 ^ n5870);
assign n12851 = ~(n11397 ^ n5821);
assign n11208 = ~(n2395 ^ n8893);
assign n3786 = n5989 & n6704;
assign n10315 = n11026 | n1509;
assign n11985 = n3324 | n12771;
assign n845 = ~(n5244 ^ n5443);
assign n7865 = n6457 | n12627;
assign n12448 = n8748 & n4814;
assign n9287 = n8054 | n3524;
assign n876 = n11527 & n8072;
assign n2913 = n4862 & n5230;
assign n1087 = n9212 & n9932;
assign n12171 = n5473 | n11792;
assign n11164 = ~(n9910 ^ n4795);
assign n3507 = n1695 & n8066;
assign n1825 = ~n1697;
assign n309 = ~n12348;
assign n4912 = ~n9026;
assign n11764 = n9432 | n7226;
assign n3088 = n8649 & n9624;
assign n7614 = ~(n5485 ^ n5083);
assign n898 = n7701 | n10486;
assign n1662 = ~(n5161 ^ n4915);
assign n6293 = n9389 | n11827;
assign n9598 = n9698 & n665;
assign n11994 = ~n4099;
assign n8193 = n8554 & n10561;
assign n10862 = n8326 | n10044;
assign n5213 = ~(n438 ^ n12631);
assign n5963 = ~(n9819 ^ n10795);
assign n381 = ~(n3941 ^ n11054);
assign n12836 = ~(n5247 ^ n9020);
assign n11301 = ~(n4034 ^ n400);
assign n4657 = n7687 | n2352;
assign n8884 = ~(n8544 ^ n5051);
assign n10433 = ~(n4500 | n1483);
assign n3880 = ~(n346 ^ n7721);
assign n2078 = n1909 & n1773;
assign n9249 = ~(n2444 | n1176);
assign n1442 = ~n7909;
assign n9253 = ~(n2918 ^ n10425);
assign n8097 = n2082 & n7007;
assign n205 = ~(n6966 | n11981);
assign n7336 = ~n10751;
assign n637 = n10601 | n3576;
assign n12877 = n10196 | n8830;
assign n5430 = n8110 | n2767;
assign n5912 = n7715 & n3883;
assign n8564 = n11457 | n4240;
assign n11122 = ~n2433;
assign n12543 = ~n10998;
assign n4819 = n4778 | n10854;
assign n6130 = n8305 | n1667;
assign n6096 = n9170 | n1162;
assign n9437 = n6687 & n2879;
assign n3951 = n3609 | n11286;
assign n7037 = n3127 | n7424;
assign n9605 = ~(n3474 ^ n8780);
assign n7000 = ~(n11233 ^ n3489);
assign n7070 = ~(n9179 | n9479);
assign n9847 = ~(n8163 ^ n4448);
assign n4640 = ~(n9846 ^ n5409);
assign n9301 = n7391 | n7341;
assign n12845 = n11547 | n6832;
assign n2281 = ~(n11390 ^ n3431);
assign n167 = n8345 | n2635;
assign n1987 = ~n7505;
assign n5124 = ~(n3864 ^ n10234);
assign n5765 = ~n11153;
assign n4662 = ~(n4135 | n5339);
assign n1872 = n2924 & n2141;
assign n3701 = ~(n10332 ^ n9484);
assign n3580 = ~n9194;
assign n2115 = ~(n4480 ^ n7123);
assign n4199 = n1972 & n3977;
assign n860 = ~(n469 ^ n7349);
assign n12540 = n2537 & n151;
assign n5616 = ~n11053;
assign n12495 = n8792 | n7972;
assign n6421 = ~(n11155 ^ n3574);
assign n5545 = ~(n10359 ^ n8424);
assign n1111 = n3743 | n3606;
assign n5562 = n12853 | n8740;
assign n10170 = ~n10034;
assign n3043 = ~(n2060 ^ n6131);
assign n2612 = ~n12619;
assign n4625 = n7977 | n755;
assign n6373 = ~n11892;
assign n1246 = n8221 | n11268;
assign n4833 = n12683 & n6552;
assign n8354 = ~n3616;
assign n2219 = n5708 & n12892;
assign n2908 = ~(n5819 ^ n1697);
assign n7227 = ~(n4170 ^ n10599);
assign n709 = n6628 & n11372;
assign n6222 = n12087 & n4267;
assign n4857 = ~(n3885 ^ n11729);
assign n2202 = ~n9275;
assign n7193 = ~(n1505 ^ n4118);
assign n11156 = ~(n4021 ^ n10654);
assign n9044 = ~(n7295 | n2785);
assign n9244 = ~(n7316 | n9090);
assign n8429 = ~n7824;
assign n2993 = n12186 | n2815;
assign n2593 = ~(n10028 ^ n4651);
assign n2557 = ~n9982;
assign n4568 = n10852 & n12019;
assign n3672 = n24 | n7334;
assign n5292 = n6718 | n795;
assign n7352 = n4100 | n9385;
assign n5042 = ~n9307;
assign n1326 = n11552 | n4642;
assign n5706 = n3820 | n8643;
assign n1190 = n7788 & n11654;
assign n4065 = n5858 | n1455;
assign n6552 = n2478 | n2387;
assign n93 = ~(n6767 ^ n1508);
assign n4360 = n4498 | n1455;
assign n6273 = ~(n10382 ^ n11167);
assign n5081 = n5964 & n11662;
assign n9982 = n7124 & n4307;
assign n7408 = ~(n12272 ^ n6950);
assign n11730 = n1757 & n303;
assign n6805 = ~(n8532 | n442);
assign n10090 = ~(n6995 ^ n9305);
assign n12273 = n4856 | n10610;
assign n6356 = ~(n913 ^ n8493);
assign n4442 = n10647 ^ n10009;
assign n2428 = n1224 & n8422;
assign n11463 = n10078 & n8652;
assign n3711 = ~(n6962 ^ n7049);
assign n8204 = n6776 & n12145;
assign n4859 = n2099 | n9586;
assign n11753 = ~n3541;
assign n10667 = n2217 | n8745;
assign n10665 = ~(n8197 ^ n1098);
assign n380 = ~n9698;
assign n8321 = n10879 | n7424;
assign n4405 = ~n4070;
assign n6802 = n9806 & n8579;
assign n10420 = ~(n3365 | n5811);
assign n9799 = ~(n9669 | n12196);
assign n9145 = ~(n1622 ^ n10189);
assign n1813 = n2102 & n517;
assign n1787 = ~(n7663 ^ n11886);
assign n11666 = n6244 & n8180;
assign n7028 = n2854 | n1961;
assign n397 = n649 ^ n8270;
assign n12220 = ~n6553;
assign n3378 = n4272 | n11833;
assign n88 = ~n1795;
assign n9094 = ~(n7254 ^ n11190);
assign n4418 = n9528 | n10054;
assign n3665 = n3819 & n2966;
assign n11113 = ~(n4060 | n2225);
assign n9083 = ~n4463;
assign n10553 = ~n987;
assign n12795 = ~(n1560 ^ n12697);
assign n12275 = n2414 & n1920;
assign n10089 = n8959 | n11122;
assign n11076 = n12853 | n3224;
assign n12062 = ~(n4273 | n11934);
assign n3361 = ~n9627;
assign n2021 = ~(n3757 ^ n10363);
assign n4976 = n632 & n4881;
assign n12685 = ~(n2230 | n7302);
assign n7984 = ~(n5332 ^ n12952);
assign n6889 = ~(n5380 ^ n4305);
assign n3074 = n6509 & n2657;
assign n4146 = n2872 | n2815;
assign n5179 = n752 | n11122;
assign n5137 = ~(n7418 ^ n3061);
assign n9736 = ~n5931;
assign n4202 = n10196 | n9568;
assign n11928 = n752 | n7395;
assign n5144 = ~(n9 ^ n12486);
assign n7129 = ~n11307;
assign n5702 = ~(n9340 ^ n263);
assign n4503 = n9945 | n11486;
assign n9097 = ~(n4074 | n5104);
assign n3750 = n10741 | n10149;
assign n6364 = n5860 & n10898;
assign n9695 = ~(n3508 ^ n12096);
assign n9260 = n11719 | n4400;
assign n815 = ~(n7062 ^ n145);
assign n2636 = ~(n2098 ^ n6959);
assign n12762 = ~(n1458 ^ n3942);
assign n6229 = ~(n3228 | n2603);
assign n12563 = ~(n6620 ^ n11660);
assign n418 = n5809 | n9188;
assign n11686 = ~(n9905 ^ n10792);
assign n9537 = ~(n861 ^ n9545);
assign n2928 = n2559 & n502;
assign n15 = n10615 & n4699;
assign n2480 = ~(n4349 ^ n4927);
assign n6043 = n5061 | n11720;
assign n6325 = n3265 | n1454;
assign n2022 = n8137 & n7076;
assign n8525 = n2833 & n553;
assign n44 = ~(n12223 ^ n4389);
assign n9986 = ~(n3464 ^ n8805);
assign n2255 = ~(n7984 ^ n6362);
assign n10137 = ~(n3233 | n4402);
assign n10141 = n8552 | n9586;
assign n1889 = n5084 & n562;
assign n10954 = ~(n9872 ^ n6941);
assign n376 = n959 | n5155;
assign n12344 = n2969 | n11072;
assign n1009 = n5575 | n2232;
assign n3491 = n7391 | n4242;
assign n5641 = n1548 ^ n6838;
assign n6345 = n4178 | n1751;
assign n10377 = n2099 | n12446;
assign n5542 = n752 | n184;
assign n2866 = ~n6085;
assign n9390 = ~(n5476 ^ n8360);
assign n1993 = n11749 | n4165;
assign n6160 = n11181 & n4268;
assign n8212 = ~(n12537 | n11978);
assign n4178 = n239 | n8788;
assign n10720 = ~(n1059 ^ n10875);
assign n11953 = n5032 | n760;
assign n11684 = ~(n489 | n10184);
assign n12059 = ~(n366 ^ n2035);
assign n8560 = n7539 | n1328;
assign n2003 = ~(n11173 ^ n8603);
assign n9743 = ~n1853;
assign n3486 = n12033 | n6781;
assign n11947 = n584 & n8887;
assign n12687 = ~n1166;
assign n4565 = ~n9993;
assign n12402 = ~(n6125 ^ n2867);
assign n4337 = n12837 & n12554;
assign n396 = n12361 | n3421;
assign n164 = n11856 | n6911;
assign n1290 = ~(n12859 | n2412);
assign n3070 = n6147 & n9876;
assign n2510 = ~(n6551 | n2086);
assign n7020 = ~(n8553 ^ n5073);
assign n5228 = n10833 | n7761;
assign n1568 = ~(n1424 | n8707);
assign n4971 = ~(n12818 ^ n11461);
assign n7528 = ~(n11414 ^ n11375);
assign n12312 = ~n7390;
assign n5013 = ~n1688;
assign n6177 = n1699 | n7928;
assign n6997 = n6795 & n11424;
assign n8961 = n11421 | n6212;
assign n10108 = ~n9080;
assign n5559 = n2099 | n7136;
assign n2650 = n5198 & n9111;
assign n3983 = n839 & n69;
assign n9188 = ~n2558;
assign n8481 = n8026 | n6197;
assign n7831 = ~(n8022 ^ n724);
assign n2516 = ~(n8449 ^ n4758);
assign n11824 = ~(n1038 ^ n3466);
assign n3762 = ~(n11559 ^ n6978);
assign n7669 = n5902 | n3911;
assign n7333 = ~(n7021 ^ n10726);
assign n4688 = ~(n8557 ^ n7275);
assign n6175 = n6977 | n7876;
assign n7269 = ~(n4963 ^ n9362);
assign n491 = n11200 & n9393;
assign n1642 = n11958 | n7425;
assign n5864 = n8354 | n8740;
assign n514 = n11013 & n1346;
assign n1780 = ~n8600;
assign n6777 = n5355 | n7246;
assign n10710 = n3324 | n795;
assign n10637 = ~(n9395 ^ n10386);
assign n11644 = ~(n5438 ^ n1856);
assign n3190 = n10882 | n9665;
assign n12789 = n9433 & n11196;
assign n8269 = n683 | n12834;
assign n5335 = n676 & n4331;
assign n1534 = n8387 | n12856;
assign n653 = ~(n1181 | n12808);
assign n12869 = ~n4331;
assign n3112 = ~(n987 ^ n6367);
assign n6335 = n2505 & n8388;
assign n9777 = n7176 | n506;
assign n1126 = n7391 | n10066;
assign n8589 = n11584 | n4156;
assign n11634 = n4311 | n2572;
assign n8307 = n10522 & n2943;
assign n7295 = n1387 & n2954;
assign n6775 = ~n8966;
assign n6808 = ~n10658;
assign n1213 = ~(n2519 ^ n4673);
assign n12234 = ~(n53 ^ n7541);
assign n2675 = n5190 | n6371;
assign n11562 = ~(n9381 ^ n7277);
assign n8821 = n298 & n8746;
assign n7603 = ~(n12730 ^ n3123);
assign n9759 = ~(n9615 | n5253);
assign n4739 = ~(n4451 | n1852);
assign n6491 = ~n2721;
assign n8579 = n8354 | n9188;
assign n4015 = n11266 | n8286;
assign n9554 = ~(n10658 | n2513);
assign n6565 = ~(n4049 ^ n11554);
assign n73 = n7884 & n1930;
assign n4702 = n7470 | n1286;
assign n6800 = n1311 & n799;
assign n6250 = ~(n6285 ^ n7515);
assign n7457 = n2099 | n12883;
assign n1701 = n7154 | n10837;
assign n2211 = n8727 & n6756;
assign n9106 = ~n253;
assign n6004 = n5575 | n2754;
assign n7260 = ~n5500;
assign n928 = n10750 | n8740;
assign n7135 = ~(n5137 ^ n7340);
assign n4476 = n7709 | n12771;
assign n2064 = ~(n3284 ^ n5841);
assign n8395 = n5915 | n6513;
assign n935 = n4727 & n4140;
assign n6155 = ~(n10843 ^ n1169);
assign n5310 = ~(n1479 | n1088);
assign n8227 = n3743 | n4864;
assign n7663 = n2099 | n8259;
assign n415 = n3776 | n7665;
assign n7989 = n4576 & n7365;
assign n2180 = n1684 & n3408;
assign n3656 = ~(n11556 ^ n6173);
assign n3158 = n6654 & n8578;
assign n11760 = ~(n12037 ^ n8968);
assign n2364 = n8476 & n5645;
assign n9645 = n5179 | n8417;
assign n8873 = ~(n548 | n2184);
assign n574 = n7709 | n9521;
assign n3206 = ~(n6518 ^ n9790);
assign n663 = ~(n9678 ^ n9384);
assign n3927 = n8443 | n12769;
assign n4142 = ~(n11400 | n7590);
assign n402 = ~(n1299 ^ n11634);
assign n8466 = ~(n6548 ^ n3910);
assign n11987 = n8441 & n10645;
assign n1611 = ~(n3213 ^ n9694);
assign n11051 = n11764 & n7533;
assign n757 = n7902 & n10675;
assign n2090 = n3145 & n1267;
assign n10067 = ~(n8827 ^ n364);
assign n1365 = ~(n8652 ^ n5293);
assign n11795 = ~(n9755 ^ n10274);
assign n5246 = ~(n9227 | n11615);
assign n10307 = ~(n1142 | n5933);
assign n5700 = n12659 & n6846;
assign n5571 = n6577 | n3468;
assign n2427 = n6577 | n3903;
assign n5620 = ~(n4719 | n5723);
assign n10066 = ~n6038;
assign n12914 = n989 | n561;
assign n1863 = n9465 & n3003;
assign n8242 = ~(n5118 ^ n4081);
assign n1593 = n257 | n5333;
assign n10490 = ~(n11400 ^ n4691);
assign n4509 = n12177 | n12386;
assign n5418 = n2564 & n9956;
assign n1573 = ~(n49 ^ n8775);
assign n7183 = ~(n4699 ^ n7565);
assign n3349 = n5470 | n4672;
assign n5037 = ~(n4799 ^ n4607);
assign n11773 = n6857 | n4544;
assign n6094 = ~(n9615 ^ n10981);
assign n1288 = n9376 & n11160;
assign n3466 = ~(n10530 ^ n3470);
assign n10086 = n2832 | n12843;
assign n9369 = n9170 | n7881;
assign n10617 = ~(n623 ^ n5157);
assign n11546 = n9492 | n4420;
assign n2519 = n10534 & n12546;
assign n1687 = ~(n11231 ^ n7553);
assign n6895 = ~(n7752 ^ n9868);
assign n3476 = ~(n5242 ^ n79);
assign n6712 = n5491 & n7743;
assign n7142 = ~(n762 ^ n6312);
assign n8340 = ~n203;
assign n10378 = ~(n8912 ^ n7830);
assign n3420 = n9895 & n1832;
assign n3533 = ~(n3880 ^ n9498);
assign n1840 = ~n5820;
assign n1076 = n3291 & n8686;
assign n8240 = ~n2680;
assign n11908 = ~(n3038 ^ n1030);
assign n6145 = n8959 | n12816;
assign n2955 = ~(n12939 ^ n6858);
assign n6759 = ~n8850;
assign n2074 = n7822 & n5165;
assign n4530 = ~(n11248 | n7525);
assign n5791 = n5530 | n4249;
assign n3224 = ~n1564;
assign n11943 = n8387 & n12856;
assign n12245 = ~(n12367 | n11600);
assign n12926 = ~(n5564 ^ n7451);
assign n10560 = ~(n4058 ^ n1554);
assign n7057 = ~(n3016 ^ n5356);
assign n1949 = ~(n312 ^ n11600);
assign n2989 = n10922 | n8021;
assign n8091 = n10928 & n4141;
assign n3626 = ~(n1786 ^ n10971);
assign n4279 = ~(n7603 ^ n11951);
assign n1435 = ~(n5346 | n9704);
assign n3485 = n3765 | n3158;
assign n2774 = ~(n7186 | n11809);
assign n9355 = n8679 & n1360;
assign n997 = ~(n8646 | n7314);
assign n7213 = n11569 | n4115;
assign n5254 = n618 | n7139;
assign n6355 = ~(n6625 ^ n7625);
assign n7525 = n4442 & n4110;
assign n8222 = n3024 & n7596;
assign n12909 = ~n9819;
assign n572 = ~(n12661 ^ n1211);
assign n1113 = n12643 & n4537;
assign n8720 = ~n11987;
assign n6477 = ~(n9657 ^ n7969);
assign n12010 = n8127 | n1851;
assign n1373 = ~(n2150 ^ n5723);
assign n2617 = ~(n9825 ^ n9776);
assign n8988 = n1151 | n4573;
assign n7335 = ~(n7915 ^ n11435);
assign n8214 = ~n9810;
assign n4959 = ~(n7001 ^ n12897);
assign n494 = n6718 | n7506;
assign n12683 = n7831 | n10979;
assign n10064 = n10018 | n10021;
assign n10563 = ~(n12460 ^ n360);
assign n2062 = ~(n12930 ^ n9350);
assign n11127 = n3131 & n10813;
assign n10161 = ~(n1975 | n11606);
assign n4604 = ~n4437;
assign n6204 = n191 | n7703;
assign n10796 = ~(n10004 | n7968);
assign n3024 = n868 | n8323;
assign n6060 = ~(n3791 ^ n11806);
assign n10526 = ~(n1681 ^ n7048);
assign n9057 = ~(n4063 ^ n179);
assign n297 = ~(n1830 | n3860);
assign n1983 = ~n9567;
assign n8079 = ~(n9928 ^ n2501);
assign n5661 = n8187 | n11827;
assign n6784 = n1315 | n2211;
assign n10446 = ~(n1439 | n9427);
assign n5195 = n3367 | n3056;
assign n6054 = ~n6335;
assign n10104 = ~(n8198 ^ n4403);
assign n11697 = ~(n5574 | n9133);
assign n11695 = n3617 | n4913;
assign n10363 = n11923 | n1509;
assign n11669 = ~(n7280 ^ n11909);
assign n6032 = n12413 & n8866;
assign n4154 = ~n12702;
assign n5597 = n2638 & n8358;
assign n9952 = ~n11459;
assign n6707 = n4560 & n11334;
assign n5998 = ~(n10710 ^ n10083);
assign n696 = ~(n8174 ^ n12937);
assign n1223 = ~(n1354 ^ n9167);
assign n5495 = ~(n5048 ^ n1159);
assign n707 = ~(n11931 ^ n4008);
assign n557 = n12346 & n12083;
assign n11309 = ~(n1352 ^ n7851);
assign n5501 = n10142 | n8524;
assign n10988 = ~n588;
assign n2781 = ~(n11279 ^ n11020);
assign n8856 = ~n5665;
assign n2938 = n10132 | n3476;
assign n843 = n3608 & n3488;
assign n4465 = n6977 | n2815;
assign n8298 = ~(n4135 ^ n8076);
assign n10400 = n3470 | n9175;
assign n2371 = n5089 & n10823;
assign n3534 = n3614 & n8539;
assign n7684 = ~(n272 ^ n3095);
assign n4198 = ~(n74 | n7776);
assign n940 = n10339 | n826;
assign n6487 = ~(n3106 ^ n1759);
assign n8838 = n11838 & n7344;
assign n9395 = n3820 | n1509;
assign n8761 = n7196 | n4087;
assign n10622 = n8831 & n3918;
assign n3328 = n6814 | n2929;
assign n904 = n10750 | n10422;
assign n7904 = n4674 | n9188;
assign n1778 = ~(n10839 | n5248);
assign n9632 = ~n2428;
assign n4589 = ~(n1632 | n11730);
assign n1907 = n8217 & n10941;
assign n12934 = ~(n11327 ^ n7000);
assign n10936 = n12119 | n8957;
assign n816 = n2099 | n3224;
assign n12228 = ~(n4435 ^ n10033);
assign n9046 = ~n11230;
assign n3592 = ~(n6282 ^ n12279);
assign n6667 = ~n7563;
assign n7958 = ~(n7873 ^ n9771);
assign n5489 = n7998 | n4153;
assign n5660 = n5886 & n770;
assign n8487 = n6275 & n3907;
assign n2690 = ~(n8429 ^ n7326);
assign n242 = ~n8526;
assign n10234 = ~n3246;
assign n10110 = n11490 & n1919;
assign n6344 = ~(n8194 ^ n4035);
assign n8477 = n11153 & n7270;
assign n7551 = n6577 | n6169;
assign n4134 = n6053 | n5830;
assign n9805 = ~(n12496 ^ n5124);
assign n8669 = n11005 | n11297;
assign n5219 = n2099 | n8655;
assign n12386 = n8959 | n6169;
assign n5633 = ~(n6350 ^ n11412);
assign n7717 = ~n1882;
assign n10034 = ~(n8395 ^ n7863);
assign n4535 = n10157 | n4642;
assign n6955 = n5054 & n6300;
assign n3294 = ~(n8520 ^ n7815);
assign n3212 = n11234 & n12522;
assign n10166 = ~(n2688 ^ n5315);
assign n291 = n8194 & n4035;
assign n6779 = ~(n5975 | n2362);
assign n2254 = n1799 | n8544;
assign n2005 = ~(n9304 ^ n549);
assign n9329 = n6544 | n6422;
assign n7176 = n12119 | n9586;
assign n9047 = ~(n11934 ^ n4273);
assign n12760 = n6941 & n6764;
assign n7249 = ~(n10153 ^ n8437);
assign n918 = ~n9270;
assign n5516 = n603 | n12688;
assign n1145 = n1696 | n3102;
assign n8414 = ~n4928;
assign n10340 = n10732 | n476;
assign n8499 = n9373 | n5502;
assign n2962 = n6408 & n5787;
assign n6959 = ~(n8141 | n12804);
assign n5993 = n7108 & n12164;
assign n5547 = n8411 & n4596;
assign n4837 = n5398 | n3248;
assign n2618 = n4911 | n7341;
assign n11437 = ~(n2138 ^ n723);
assign n11220 = n585 & n4670;
assign n8795 = ~(n9514 | n3751);
assign n154 = ~(n9017 | n8199);
assign n2943 = n6709 & n8356;
assign n8587 = n11556 | n6173;
assign n11247 = n3155 & n7213;
assign n10594 = n4116 | n7188;
assign n8431 = n11933 | n11322;
assign n8270 = ~(n6520 ^ n5991);
assign n5756 = ~(n6517 ^ n10246);
assign n9215 = n8221 & n11268;
assign n10754 = n3617 | n5468;
assign n6227 = n11060 | n11247;
assign n8814 = n10157 | n1509;
assign n11243 = n9777 & n9309;
assign n10471 = ~(n8518 | n5697);
assign n9375 = ~(n7758 ^ n793);
assign n7182 = ~(n4395 ^ n7923);
assign n9808 = n6142 & n830;
assign n3988 = ~(n9197 ^ n12110);
assign n12776 = n2564 & n2585;
assign n2292 = ~n3817;
assign n877 = ~(n12178 ^ n1481);
assign n5384 = n5355 | n1546;
assign n461 = ~(n2885 ^ n9715);
assign n8250 = ~(n359 ^ n9357);
assign n130 = ~n2512;
assign n1713 = ~(n2365 ^ n932);
assign n39 = ~(n10152 ^ n1693);
assign n3775 = n3992 & n11876;
assign n536 = ~(n5206 ^ n2311);
assign n2443 = ~(n2481 ^ n3504);
assign n480 = ~(n6039 ^ n10488);
assign n11409 = ~(n11076 ^ n7142);
assign n11852 = ~n4990;
assign n3092 = ~(n10844 ^ n8471);
assign n10891 = ~n9385;
assign n5675 = ~(n7268 ^ n1767);
assign n5783 = n8336 & n9640;
assign n3722 = ~(n11352 ^ n12265);
assign n3152 = ~n187;
assign n2065 = ~(n3665 | n2452);
assign n654 = ~(n8282 ^ n12298);
assign n3737 = ~(n11405 | n9285);
assign n8061 = ~(n1031 ^ n9297);
assign n2526 = ~(n10414 ^ n10369);
assign n7311 = n10339 | n12535;
assign n10537 = ~(n4829 ^ n11301);
assign n7327 = n2217 | n4527;
assign n2692 = ~(n7835 | n8885);
assign n6830 = ~(n3108 ^ n6610);
assign n354 = n636 | n6513;
assign n836 = ~n5418;
assign n4080 = ~n5841;
assign n10386 = ~n7205;
assign n8243 = n2792 & n5060;
assign n2830 = ~n4017;
assign n2750 = n6475 | n10867;
assign n7852 = ~(n3826 ^ n2613);
assign n4072 = ~(n6556 ^ n6007);
assign n7724 = ~(n11128 | n558);
assign n10614 = n6914 | n4447;
assign n26 = ~n7922;
assign n4577 = ~(n985 ^ n5558);
assign n11405 = n3324 | n9521;
assign n6901 = n9792 | n7554;
assign n2407 = ~(n1844 | n6094);
assign n4824 = n11567 & n4209;
assign n4594 = ~(n5001 ^ n6787);
assign n9866 = ~(n2329 ^ n8000);
assign n9758 = n12155 | n6473;
assign n5989 = n10835 | n4875;
assign n9687 = n9529 | n7950;
assign n7601 = ~n1905;
assign n1274 = ~(n10790 ^ n11235);
assign n12244 = n982 & n8230;
assign n1749 = n10129 | n11946;
assign n10308 = n4238 & n6304;
assign n11583 = ~(n1459 ^ n1984);
assign n1771 = ~(n961 ^ n1359);
assign n2023 = ~n8410;
assign n12547 = n8309 & n10441;
assign n6605 = ~(n8412 ^ n3429);
assign n2649 = n10874 & n1300;
assign n5551 = n8229 & n1276;
assign n2911 = ~(n4442 | n4110);
assign n7668 = n137 & n7610;
assign n3621 = ~n4520;
assign n8447 = ~(n4357 ^ n10299);
assign n4109 = ~(n240 ^ n1076);
assign n10140 = ~(n5044 ^ n7639);
assign n6310 = n10750 | n12446;
assign n12509 = ~(n7599 | n8910);
assign n4272 = ~(n2304 ^ n4839);
assign n8201 = ~n11363;
assign n6570 = ~(n12055 ^ n8246);
assign n2486 = ~(n2838 ^ n6164);
assign n72 = ~(n10015 ^ n12517);
assign n316 = ~n985;
assign n2715 = ~n10443;
assign n11218 = ~(n9453 | n9646);
assign n888 = n610 & n469;
assign n12585 = ~n11784;
assign n9440 = n399 & n7949;
assign n8349 = n1960 & n1019;
assign n4376 = ~n10974;
assign n4417 = ~(n12432 ^ n6162);
assign n712 = ~(n644 ^ n9966);
assign n8185 = ~n6935;
assign n6083 = ~(n8481 ^ n1048);
assign n2006 = n10893 & n9121;
assign n6237 = n9373 | n4474;
assign n10487 = n2456 | n12754;
assign n6559 = n4079 & n150;
assign n1788 = ~(n6607 | n10753);
assign n7027 = n10750 | n12535;
assign n2613 = ~(n685 ^ n12191);
assign n5638 = ~n1637;
assign n9229 = ~(n11171 ^ n5712);
assign n9916 = n5794 & n4340;
assign n5400 = n10057 & n5822;
assign n11036 = n11958 | n11122;
assign n12129 = ~n3467;
assign n4313 = n7301 | n10158;
assign n3110 = n9616 | n5262;
assign n1156 = n2973 | n9613;
assign n6201 = ~(n12180 ^ n4558);
assign n3819 = ~n10414;
assign n1910 = n5404 | n6823;
assign n6672 = n11801 | n10413;
assign n5836 = n4628 | n2964;
assign n11553 = n10899 & n7532;
assign n11591 = n11887 | n4913;
assign n10923 = n6481 & n7437;
assign n7231 = n2012 & n11497;
assign n11972 = ~(n3067 ^ n1793);
assign n11042 = n6945 & n423;
assign n6220 = ~(n6585 ^ n12534);
assign n11573 = ~n3027;
assign n2330 = ~(n10498 ^ n7857);
assign n11328 = n5780 | n960;
assign n6108 = n1621 | n1331;
assign n8977 = n9784 | n6920;
assign n7477 = n4567 & n9960;
assign n12622 = n6577 | n11820;
assign n5070 = ~(n3716 | n3586);
assign n6908 = n7167 & n2477;
assign n4605 = ~(n12231 ^ n5041);
assign n7431 = ~n12166;
assign n6097 = ~(n7073 ^ n9628);
assign n4945 = ~n4851;
assign n5115 = ~(n6497 ^ n10554);
assign n4927 = ~(n5368 ^ n11651);
assign n11906 = ~(n4388 ^ n4898);
assign n7679 = n7643 & n913;
assign n7840 = n1854 & n4620;
assign n11400 = ~(n3089 ^ n3692);
assign n6314 = ~n9444;
assign n6063 = ~(n8902 ^ n12784);
assign n1408 = n9394 & n6789;
assign n10117 = n12833 | n984;
assign n6810 = n4724 | n7896;
assign n8393 = n11923 | n8285;
assign n11964 = n10740 & n5703;
assign n10849 = n3930 | n4483;
assign n11099 = n1911 & n1004;
assign n3197 = ~n9131;
assign n7543 = ~(n7127 ^ n7774);
assign n786 = ~(n95 | n6792);
assign n392 = n9170 | n7424;
assign n12874 = n9005 | n1608;
assign n3709 = n969 & n5046;
assign n4866 = n9373 | n4527;
assign n10692 = n5860 & n5760;
assign n11951 = ~(n7502 ^ n12213);
assign n1368 = n566 | n5656;
assign n6669 = n5355 | n4775;
assign n4362 = ~(n2458 ^ n12238);
assign n9009 = n9343 | n12425;
assign n2101 = n2448 | n3799;
assign n10068 = ~n11653;
assign n6504 = n3625 & n9031;
assign n11128 = n11433 | n5540;
assign n7 = ~(n3476 ^ n1193);
assign n12087 = n12069 & n2558;
assign n12240 = ~(n12318 ^ n6900);
assign n1596 = ~(n10374 ^ n3898);
assign n5899 = n2913 ^ n368;
assign n11336 = n7043 & n7190;
assign n3162 = n10983 & n2817;
assign n3309 = n11036 & n8030;
assign n1140 = ~(n11692 | n12484);
assign n8693 = ~(n9348 ^ n7667);
assign n1946 = n10196 | n4642;
assign n8766 = n9389 | n1738;
assign n4718 = n1041 & n11364;
assign n4569 = ~(n7726 ^ n5533);
assign n7626 = n7874 | n12918;
assign n8890 = ~n3163;
assign n5162 = ~(n10960 ^ n10315);
assign n1619 = n8743 & n9505;
assign n4018 = n9884 | n3411;
assign n682 = n8785 & n6021;
assign n10123 = ~n6001;
assign n3106 = n11070 & n4599;
assign n5027 = n8412 | n3521;
assign n10874 = n5530 | n1163;
assign n11702 = ~(n3397 ^ n6382);
assign n5341 = n994 | n1546;
assign n2740 = ~n9298;
assign n1722 = n11900 & n8871;
assign n2426 = ~(n7376 ^ n7465);
assign n7306 = n8428 | n11896;
assign n9515 = ~(n7585 ^ n8283);
assign n9401 = n2917 | n2465;
assign n6008 = ~(n6051 ^ n9635);
assign n12485 = ~(n3712 | n9805);
assign n6210 = ~(n1884 ^ n3312);
assign n12735 = ~n6254;
assign n8075 = ~(n6506 ^ n12372);
assign n8737 = n11026 | n1047;
assign n10949 = ~(n948 ^ n7482);
assign n6159 = n8418 & n11472;
assign n10734 = n5215 & n8095;
assign n11802 = n9970 & n2224;
assign n6303 = n4604 | n5220;
assign n6205 = n6995 & n2405;
assign n3721 = ~n12757;
assign n6013 = n8192 | n10193;
assign n6807 = ~(n10610 ^ n1855);
assign n4479 = ~(n2109 | n6274);
assign n4342 = ~n11491;
assign n3265 = n12119 | n12735;
assign n12549 = n4674 | n826;
assign n12816 = ~n12709;
assign n2298 = n5573 & n7618;
assign n2951 = ~(n7732 | n11246);
assign n2302 = ~n6015;
assign n9705 = n10396 | n11491;
assign n2789 = ~(n9515 ^ n2825);
assign n12920 = n7283 | n7389;
assign n1990 = n3743 | n1476;
assign n9814 = n395 ^ n8479;
assign n7322 = n2217 | n8285;
assign n5917 = n1446 | n10492;
assign n8077 = ~(n574 ^ n6427);
assign n6656 = ~n4273;
assign n580 = ~n6242;
assign n11054 = ~(n8836 ^ n11376);
assign n4502 = n2272 & n10258;
assign n3284 = n8026 | n11122;
assign n987 = n7617 & n9667;
assign n2753 = n12644 | n265;
assign n1247 = n6145 | n3647;
assign n6195 = n7495 | n3911;
assign n4613 = n10196 | n1047;
assign n8614 = ~(n11984 ^ n6460);
assign n6949 = ~(n10155 ^ n2140);
assign n6855 = n3627 & n7265;
assign n8241 = n7965 & n10848;
assign n8490 = ~(n478 ^ n12475);
assign n1308 = n686 | n3903;
assign n7191 = ~(n11343 | n3499);
assign n10851 = n11557 ^ n12360;
assign n12195 = n3746 | n995;
assign n11683 = ~(n9987 | n2361);
assign n6664 = ~(n8786 ^ n2419);
assign n3741 = n5151 & n11670;
assign n6172 = n4666 | n10863;
assign n10522 = n6770 & n4370;
assign n8438 = ~n12123;
assign n9314 = n880 | n11758;
assign n6940 = ~(n1448 | n5789);
assign n9381 = ~(n11148 ^ n12140);
assign n7120 = n2017 | n2883;
assign n8273 = n2456 | n12735;
assign n3505 = n10091 & n100;
assign n12870 = n1717 & n3813;
assign n9878 = ~n6294;
assign n1129 = ~n1689;
assign n9859 = n636 | n2964;
assign n7788 = n2584 | n9258;
assign n6047 = ~(n6033 | n214);
assign n2843 = ~n9465;
assign n7224 = n7236 & n8028;
assign n8 = n3156 & n12008;
assign n2902 = ~(n11187 ^ n7671);
assign n1515 = n12007 | n2328;
assign n9764 = n8552 | n8648;
assign n2268 = n9389 | n3911;
assign n10585 = n1051 | n7876;
assign n4869 = ~n10399;
assign n11620 = ~(n7898 ^ n2622);
assign n4855 = ~(n7911 | n5323);
assign n12900 = ~n85;
assign n5456 = n5575 | n6197;
assign n3532 = ~(n1409 ^ n12780);
assign n2327 = n418 | n7924;
assign n2306 = ~(n4781 | n138);
assign n2970 = n6237 | n9526;
assign n7092 = ~(n11405 ^ n11665);
assign n1865 = n12361 | n11896;
assign n7888 = n5838 | n10892;
assign n7645 = n1890 | n3343;
assign n4591 = n5765 | n609;
assign n5804 = ~(n8191 ^ n11176);
assign n166 = ~n12778;
assign n8965 = ~(n10467 ^ n12288);
assign n11975 = n11668 & n7538;
assign n12203 = n191 | n4775;
assign n228 = ~(n3075 ^ n314);
assign n11648 = n11856 & n6911;
assign n2521 = n3026 | n3896;
assign n3976 = n5355 | n8524;
assign n1002 = n6894 & n7105;
assign n3516 = n7044 & n10185;
assign n2008 = n12361 | n2232;
assign n6416 = ~n10466;
assign n12749 = n4994 & n2980;
assign n6261 = n8214 | n10857;
assign n5984 = n6718 | n7921;
assign n546 = ~(n10019 | n11667);
assign n5753 = n3153 | n6982;
assign n4233 = ~(n8378 ^ n8061);
assign n5482 = n2067 & n12568;
assign n1855 = ~(n4856 ^ n3348);
assign n6755 = ~n2903;
assign n3960 = ~(n8934 ^ n10460);
assign n3410 = n444 & n12829;
assign n9506 = n3620 & n5718;
assign n3449 = n3820 | n5258;
assign n2121 = n11080 & n12597;
assign n9316 = ~(n10059 ^ n10827);
assign n10265 = n2226 & n8819;
assign n7385 = ~(n12827 ^ n1674);
assign n14 = ~(n4994 ^ n2980);
assign n1436 = n4644 & n11624;
assign n12371 = ~n1322;
assign n6863 = ~n3354;
assign n3905 = n10347 | n12182;
assign n6391 = n5016 | n12202;
assign n5441 = n2456 | n3924;
assign n9625 = ~n8370;
assign n11530 = ~(n11286 ^ n12320);
assign n3388 = n5404 & n6823;
assign n9588 = n3050 | n11524;
assign n4821 = ~(n7247 ^ n199);
assign n9207 = ~(n1350 | n1912);
assign n1071 = n7536 | n1191;
assign n1754 = ~(n646 | n494);
assign n858 = ~(n1746 ^ n2404);
assign n10320 = ~(n11490 | n1919);
assign n3233 = ~(n5969 | n1313);
assign n10139 = n2217 | n4642;
assign n11391 = ~(n6801 ^ n6011);
assign n177 = ~n9289;
assign n133 = n10108 | n5497;
assign n11763 = ~(n10587 ^ n12727);
assign n7298 = n602 | n10024;
assign n6333 = ~(n8445 ^ n9766);
assign n871 = ~(n11712 ^ n9574);
assign n6129 = ~(n3335 ^ n9062);
assign n8645 = n2244 | n9402;
assign n62 = n12324 & n2736;
assign n3143 = ~(n12653 ^ n5229);
assign n11244 = n2033 | n8014;
assign n4432 = n989 | n4400;
assign n10838 = n10157 | n8830;
assign n644 = ~(n8116 ^ n9576);
assign n7002 = n2652 & n3518;
assign n12084 = ~(n2899 ^ n4182);
assign n2098 = ~(n1907 | n12566);
assign n5576 = ~(n5584 ^ n5672);
assign n4173 = n2874 | n9587;
assign n8575 = n12698 | n2298;
assign n446 = ~(n9363 ^ n4807);
assign n11012 = ~(n10810 ^ n4144);
assign n7532 = n884 | n3639;
assign n11891 = ~n6439;
assign n9895 = n3344 | n11086;
assign n3382 = n10343 | n9535;
assign n10940 = n9170 | n2358;
assign n5367 = ~(n5720 | n6565);
assign n10501 = n9908 & n12874;
assign n1947 = n7417 | n2149;
assign n4452 = ~n623;
assign n9373 = ~n6358;
assign n2759 = ~(n1154 ^ n10804);
assign n10997 = n8187 | n12328;
assign n9665 = n432 & n9549;
assign n12739 = n3096 | n3903;
assign n6753 = ~(n8580 ^ n6223);
assign n9293 = ~(n6938 ^ n5481);
assign n8950 = ~(n880 ^ n5131);
assign n5528 = n12953 | n4878;
assign n1483 = n11719 | n3911;
assign n12102 = ~n5901;
assign n11161 = n6320 | n2821;
assign n1727 = n2539 | n5910;
assign n6184 = n9101 | n9516;
assign n11853 = ~(n12200 ^ n12789);
assign n10132 = n515 & n5941;
assign n6217 = ~(n4791 ^ n5925);
assign n1269 = ~(n10631 ^ n2095);
assign n55 = n4984 & n9153;
assign n2070 = ~(n646 ^ n11540);
assign n6782 = n4498 | n7424;
assign n9819 = ~(n10648 ^ n8179);
assign n2611 = ~(n1680 ^ n31);
assign n335 = n4948 & n12021;
assign n8462 = n3262 | n4072;
assign n11916 = ~(n2713 | n6937);
assign n5136 = n3617 | n8740;
assign n7268 = ~(n9460 ^ n6159);
assign n12690 = n9274 & n10814;
assign n4352 = ~(n10279 | n9855);
assign n11977 = ~n8051;
assign n10313 = ~(n7650 ^ n3);
assign n524 = ~n2481;
assign n3107 = n1898 | n3673;
assign n9807 = n11838 | n7344;
assign n11722 = n2976 | n11495;
assign n4248 = ~(n10255 ^ n696);
assign n8700 = n1598 & n5564;
assign n1885 = ~(n11535 ^ n8403);
assign n1048 = n3933 & n3406;
assign n3648 = n9176 | n12409;
assign n4285 = ~n4414;
assign n11368 = n7709 | n9160;
assign n4349 = ~(n2321 ^ n5704);
assign n6473 = n3820 | n9521;
assign n6752 = ~(n2319 | n10252);
assign n2574 = ~n2761;
assign n199 = ~(n11517 ^ n5883);
assign n5749 = n4274 | n11810;
assign n6107 = ~(n3533 ^ n1284);
assign n11681 = n4957 & n7771;
assign n10084 = ~(n4747 ^ n2534);
assign n4544 = n11026 | n28;
assign n591 = n11142 & n10187;
assign n2894 = n10738 & n3150;
assign n12718 = ~(n9853 ^ n1831);
assign n2493 = n4657 | n3971;
assign n4884 = ~n7224;
assign n3427 = ~(n1007 | n10410);
assign n4350 = ~n1485;
assign n6841 = ~(n9518 ^ n5197);
assign n8326 = ~n9591;
assign n8565 = ~(n3915 ^ n11558);
assign n10237 = n7906 & n9794;
assign n8911 = ~(n457 ^ n8086);
assign n6074 = n9170 | n4400;
assign n5739 = n191 | n2358;
assign n585 = n6877 & n3602;
assign n7157 = ~(n2352 ^ n2643);
assign n10970 = ~(n1433 ^ n5853);
assign n4716 = n2099 | n8648;
assign n6498 = n12503 | n4527;
assign n12260 = ~(n8608 | n8160);
assign n11542 = n11641 | n12379;
assign n6793 = n306 | n40;
assign n10252 = n11923 | n5502;
assign n3165 = n4352 | n1388;
assign n4001 = n989 | n7703;
assign n1691 = ~n972;
assign n2792 = n5235 | n433;
assign n12155 = n6718 | n4875;
assign n12289 = n2099 | n6071;
assign n4311 = ~(n4224 | n7290);
assign n7941 = n11324 & n12756;
assign n9379 = n191 | n510;
assign n2333 = ~(n8499 ^ n7574);
assign n2095 = ~(n3184 ^ n11333);
assign n7707 = n4183 | n3886;
assign n12885 = ~(n6174 ^ n1885);
assign n6066 = n3743 | n1047;
assign n11703 = ~(n11713 ^ n4695);
assign n3945 = n10845 & n8426;
assign n4825 = ~n12398;
assign n9659 = ~n10160;
assign n5447 = ~(n11835 ^ n2891);
assign n8666 = ~(n8439 ^ n8953);
assign n8845 = ~n12455;
assign n10978 = ~(n5739 ^ n10241);
assign n4409 = ~(n7509 ^ n9998);
assign n8180 = n7709 | n2020;
assign n2217 = ~n11222;
assign n10279 = ~n2569;
assign n5047 = ~(n10434 ^ n1362);
assign n8188 = ~(n8290 | n5095);
assign n12332 = n2456 | n8259;
assign n10295 = n5209 & n10312;
assign n8635 = ~(n6393 | n1343);
assign n3950 = ~n6369;
assign n9970 = n8002 | n8934;
assign n9660 = ~(n4726 ^ n8098);
assign n2257 = n2097 & n3792;
assign n5665 = n9400 & n7354;
assign n12721 = n320 | n8869;
assign n11433 = ~n10678;
assign n5420 = ~(n9980 | n1587);
assign n5355 = ~n5305;
assign n7711 = ~(n9701 ^ n6861);
assign n2828 = ~(n12336 ^ n3572);
assign n12662 = ~n3513;
assign n9762 = ~(n2590 | n1544);
assign n5204 = n7449 | n1047;
assign n7869 = n5765 | n7506;
assign n4413 = n7391 | n510;
assign n4078 = n597 | n5896;
assign n6827 = n3383 | n2297;
assign n3746 = ~n6776;
assign n6723 = n11893 & n9885;
assign n11772 = ~(n8374 ^ n3113);
assign n11268 = ~(n2100 ^ n4650);
assign n10866 = ~(n8847 ^ n9356);
assign n5500 = ~(n12856 ^ n7698);
assign n1437 = ~n10753;
assign n10355 = n4535 & n501;
assign n9310 = ~(n1435 ^ n9040);
assign n5734 = ~(n8954 ^ n6852);
assign n9026 = ~(n5405 ^ n8025);
assign n9934 = ~n5849;
assign n2017 = n10614 & n7859;
assign n3809 = ~(n3968 ^ n11016);
assign n4695 = ~(n11419 | n12685);
assign n246 = n3240 | n8801;
assign n11593 = n3127 | n10066;
assign n8047 = ~(n2308 ^ n10415);
assign n3418 = n12119 | n4249;
assign n4027 = ~(n8102 | n5006);
assign n11366 = n1791 & n5344;
assign n11422 = ~n4651;
assign n2291 = ~(n11540 | n1736);
assign n7331 = n3746 | n5538;
assign n2213 = n10835 | n5258;
assign n10349 = ~(n5567 | n7187);
assign n4510 = n5765 | n5258;
assign n4795 = ~(n9982 ^ n10923);
assign n11144 = ~n9676;
assign n8851 = n5331 & n5645;
assign n7810 = ~n8672;
assign n10423 = n3838 | n5529;
assign n8249 = ~(n6331 ^ n1383);
assign n10850 = n804 & n3714;
assign n11179 = n9170 | n10066;
assign n4390 = n7283 | n12328;
assign n11575 = n1114 & n12030;
assign n2404 = ~(n5475 ^ n1395);
assign n6811 = ~n3821;
assign n12294 = ~n12248;
assign n4820 = ~(n810 | n2058);
assign n4719 = ~n2150;
assign n4152 = n6910 | n2668;
assign n7274 = ~n3601;
assign n4038 = n12340 | n1385;
assign n1061 = n1699 | n9586;
assign n3893 = ~(n4119 ^ n6949);
assign n2367 = ~n45;
assign n6481 = n5730 | n10407;
assign n10715 = n1402 & n5866;
assign n7123 = n6784 & n2103;
assign n127 = n5832 | n6531;
assign n2077 = ~(n5269 ^ n1535);
assign n2138 = ~(n1694 ^ n3727);
assign n11159 = ~n7954;
assign n4003 = ~(n8799 ^ n4811);
assign n8703 = ~n3588;
assign n9466 = n7732 & n11246;
assign n4653 = ~n6342;
assign n3395 = n10196 | n5258;
assign n759 = ~(n4036 ^ n9503);
assign n10044 = ~(n9610 ^ n8172);
assign n1560 = n11552 | n795;
assign n12817 = n3747 & n12249;
assign n2680 = n12705 & n2879;
assign n608 = ~n7039;
assign n5601 = n11923 | n9160;
assign n1565 = n4750 | n4652;
assign n6726 = ~n8130;
assign n1577 = n949 & n5917;
assign n2899 = n5355 | n130;
assign n5990 = n910 | n9852;
assign n12475 = ~(n4460 ^ n5272);
assign n4232 = n2099 | n8957;
assign n70 = ~(n3758 ^ n7031);
assign n168 = n11305 | n10501;
assign n1377 = n6451 | n2894;
assign n8265 = ~n1922;
assign n1254 = n8094 | n12865;
assign n5395 = n4469 | n1428;
assign n2506 = ~n6092;
assign n6268 = n2099 | n5781;
assign n7021 = n8552 | n530;
assign n3184 = ~(n5221 ^ n8032);
assign n4735 = ~n8049;
assign n1823 = ~(n7942 ^ n2484);
assign n12340 = ~n6813;
assign n12043 = n11093 | n9211;
assign n10600 = ~n3705;
assign n6266 = ~(n6779 ^ n4801);
assign n1601 = n5397 | n9174;
assign n9582 = ~n3350;
assign n4671 = ~(n3579 | n4342);
assign n12542 = n2660 & n10205;
assign n8367 = ~n1201;
assign n86 = ~(n10964 ^ n1311);
assign n7785 = ~n3968;
assign n6965 = ~(n12502 | n11276);
assign n519 = n1539 | n11827;
assign n2133 = n2400 & n2705;
assign n3512 = n4997 & n3937;
assign n7348 = n752 | n12274;
assign n1196 = ~(n2858 | n10188);
assign n6792 = ~(n2373 ^ n3696);
assign n9360 = n9826 & n3979;
assign n6076 = ~n42;
assign n9394 = n7037 | n3232;
assign n12157 = n7391 | n1162;
assign n9458 = ~n11086;
assign n3979 = ~n6771;
assign n5519 = n8197 & n1098;
assign n2979 = n9170 | n1079;
assign n8685 = ~n2632;
assign n9165 = n1277 & n4946;
assign n10152 = n9377 & n6523;
assign n5897 = ~n10558;
assign n3925 = ~(n8447 | n203);
assign n9200 = ~(n5231 ^ n7537);
assign n10387 = ~(n12064 ^ n11987);
assign n1545 = ~(n5859 ^ n12038);
assign n6317 = n3257 & n4096;
assign n6887 = ~n3894;
assign n8313 = n10835 | n8643;
assign n2256 = ~n2007;
assign n995 = ~n9189;
assign n3360 = ~(n8260 ^ n12065);
assign n245 = ~(n8362 ^ n12232);
assign n1359 = n2524 & n11431;
assign n3189 = ~(n538 ^ n8465);
assign n11253 = n11509 | n6804;
assign n4890 = ~(n2176 | n8516);
assign n12601 = ~n2336;
assign n11774 = ~(n7912 ^ n4136);
assign n4620 = ~(n6479 ^ n877);
assign n12292 = ~(n6370 ^ n5408);
assign n10175 = ~(n5746 ^ n7472);
assign n6183 = ~(n7330 | n11630);
assign n8998 = ~(n4823 ^ n7140);
assign n1633 = ~n10138;
assign n823 = ~(n9438 ^ n8744);
assign n9135 = ~(n1249 ^ n7963);
assign n12667 = ~(n4392 ^ n11710);
assign n5242 = n5809 | n3224;
assign n1080 = ~(n4732 ^ n8773);
assign n4297 = n8567 | n10536;
assign n5127 = ~n847;
assign n9974 = n8187 | n8524;
assign n5614 = n12648 & n521;
assign n320 = n6577 | n7952;
assign n12168 = n3271 & n6179;
assign n7324 = n7116 | n3421;
assign n7233 = n2226 & n8595;
assign n9600 = n10180 | n4234;
assign n6719 = n2605 | n11921;
assign n730 = ~(n2032 ^ n1939);
assign n1387 = ~n3491;
assign n2435 = ~(n888 | n8328);
assign n4168 = n6687 & n7265;
assign n7801 = n3746 | n2232;
assign n12930 = ~n84;
assign n9662 = n9645 & n12301;
assign n75 = ~(n5100 ^ n6264);
assign n3531 = n3870 & n7120;
assign n7288 = n5494 | n5401;
assign n11341 = ~n6222;
assign n9648 = n12361 | n3903;
assign n7957 = ~(n4968 ^ n6992);
assign n5746 = n9306 & n4078;
assign n8551 = n11466 | n8222;
assign n1540 = ~(n12823 ^ n1143);
assign n1849 = ~(n6759 ^ n11160);
assign n10767 = ~n11325;
assign n5611 = n11723 & n12821;
assign n3412 = n3020 & n1355;
assign n10114 = n4589 | n9128;
assign n140 = ~n7452;
assign n6839 = ~n1702;
assign n11080 = n752 | n12899;
assign n6865 = ~(n9915 ^ n1496);
assign n8496 = ~n12788;
assign n8762 = ~(n6686 | n5407);
assign n5817 = n12248 | n7723;
assign n2373 = ~(n6308 ^ n5352);
assign n264 = ~n11997;
assign n12423 = n12119 | n1932;
assign n10205 = n6095 | n781;
assign n5164 = n3658 & n10207;
assign n12110 = n12397 & n11508;
assign n2862 = n8552 | n4913;
assign n5472 = ~(n8406 ^ n3783);
assign n10238 = ~(n11312 ^ n8586);
assign n9158 = n2516 | n11559;
assign n4226 = n6527 ^ n10214;
assign n12606 = n3279 & n6871;
assign n4836 = ~(n12552 ^ n8115);
assign n7894 = ~n10152;
assign n782 = n11476 | n1125;
assign n8498 = ~(n7861 | n5327);
assign n1953 = ~(n12224 ^ n5268);
assign n4165 = ~(n8081 ^ n11340);
assign n4628 = ~n8476;
assign n11236 = n1937 | n5012;
assign n9323 = n4784 | n3419;
assign n3273 = n10108 | n1162;
assign n11198 = ~(n7627 ^ n12128);
assign n10696 = n9389 | n561;
assign n1181 = n8127 | n5497;
assign n781 = ~(n10567 ^ n2771);
assign n911 = ~(n11756 ^ n10459);
assign n3021 = n9373 | n2020;
assign n890 = n1811 | n829;
assign n11347 = ~n7440;
assign n6763 = n7901 | n5701;
assign n7430 = ~(n9146 ^ n2453);
assign n10592 = ~(n9565 ^ n6469);
assign n6639 = ~(n251 ^ n8980);
assign n11828 = ~(n9310 ^ n10043);
assign n11819 = ~(n6442 ^ n3462);
assign n3999 = ~(n10887 | n323);
assign n5061 = n5780 & n960;
assign n8743 = n8759 & n2024;
assign n5344 = n2813 & n7613;
assign n2259 = ~n5694;
assign n4511 = n9367 | n7471;
assign n1729 = ~n11508;
assign n457 = ~(n10656 ^ n12903);
assign n6245 = n8207 | n8650;
assign n8925 = n3845 & n10733;
assign n5830 = ~(n8468 ^ n8278);
assign n9616 = n10750 | n5326;
assign n3848 = n5219 | n4926;
assign n11595 = n8026 | n9971;
assign n2686 = n2099 | n8644;
assign n1964 = ~(n5404 ^ n6823);
assign n5646 = n5594 & n11095;
assign n8199 = n7457 & n872;
assign n7606 = ~(n463 | n625);
assign n12468 = n488 | n10691;
assign n8852 = n6718 | n8285;
assign n2971 = ~n8656;
assign n7147 = ~n8266;
assign n8324 = ~(n2467 ^ n311);
assign n10656 = n12853 | n826;
assign n247 = ~(n4429 ^ n4659);
assign n6412 = ~n3472;
assign n11894 = n9837 | n6529;
assign n10515 = n5681 & n10646;
assign n7134 = n9688 & n8446;
assign n7101 = n6577 | n11775;
assign n2704 = n3743 | n3451;
assign n11017 = n8127 | n10066;
assign n7839 = ~n10510;
assign n10615 = ~(n8009 ^ n4744);
assign n10179 = n12800 | n9418;
assign n12185 = ~(n9391 | n5302);
assign n680 = n1557 & n7030;
assign n11089 = ~(n5780 ^ n960);
assign n1321 = n1051 | n6197;
assign n6068 = n11822 & n8382;
assign n7745 = n10745 | n12072;
assign n11751 = n8959 | n8768;
assign n2111 = n8959 | n7558;
assign n8118 = n7391 | n7424;
assign n2477 = ~(n9360 ^ n4260);
assign n1491 = n8550 & n10934;
assign n6475 = n8187 | n12843;
assign n4373 = n2217 | n609;
assign n4789 = n8395 | n10588;
assign n7950 = n11110 & n10794;
assign n7812 = ~(n7429 ^ n4344);
assign n6923 = ~(n10128 | n6714);
assign n7625 = n10636 & n367;
assign n2157 = n7992 & n8569;
assign n8310 = n8552 | n12080;
assign n11053 = ~(n3987 ^ n11636);
assign n6896 = n10466 & n2678;
assign n8283 = ~(n12046 ^ n1287);
assign n11829 = n8778 | n12718;
assign n8550 = n2217 | n5759;
assign n11287 = ~n9720;
assign n11657 = n4205 | n10817;
assign n8513 = ~n917;
assign n12092 = n9661 & n5130;
assign n4658 = n4788 & n9620;
assign n12187 = ~n5622;
assign n4035 = n10879 | n11746;
assign n517 = n4179 | n8266;
assign n548 = n9370 | n8524;
assign n4030 = ~(n7276 ^ n5974);
assign n9319 = ~(n285 ^ n180);
assign n5755 = n1070 & n4306;
assign n5868 = ~(n3433 | n1722);
assign n10078 = n3836 | n12371;
assign n9129 = ~(n5384 ^ n12652);
assign n11043 = n1382 & n11657;
assign n4145 = n10545 & n1512;
assign n6414 = n12361 | n2815;
assign n6395 = n10212 & n907;
assign n4704 = ~(n1760 | n2859);
assign n6336 = ~(n12579 | n6506);
assign n4747 = n10224 & n11452;
assign n11004 = ~(n805 | n7656);
assign n3579 = ~(n3753 ^ n2941);
assign n6156 = ~(n12870 ^ n440);
assign n9861 = ~(n2947 | n940);
assign n5269 = ~(n10608 ^ n5950);
assign n9481 = n4628 | n12446;
assign n5088 = ~n11533;
assign n12052 = n8187 | n1915;
assign n11665 = ~(n10148 ^ n7996);
assign n5731 = ~(n9626 ^ n1597);
assign n3459 = ~(n867 ^ n4731);
assign n334 = n9878 | n3224;
assign n7692 = ~(n7151 ^ n1501);
assign n6039 = n12673 & n10440;
assign n5125 = n9688 | n8446;
assign n5439 = ~n3130;
assign n9686 = ~(n12123 ^ n9490);
assign n1741 = ~n7920;
assign n11274 = n10124 & n455;
assign n9113 = ~(n4420 ^ n1603);
assign n492 = n9370 | n4242;
assign n3920 = n2845 & n4177;
assign n5556 = ~(n10667 ^ n8317);
assign n8251 = n8187 | n6389;
assign n89 = n3363 | n5509;
assign n7814 = ~(n4524 ^ n10068);
assign n6734 = n8193 & n5002;
assign n9876 = n4894 | n36;
assign n1608 = ~(n9787 ^ n1904);
assign n10539 = ~(n1705 ^ n12251);
assign n8577 = ~n9550;
assign n5259 = ~(n1112 ^ n8588);
assign n10057 = n8870 | n8655;
assign n2897 = ~(n7505 ^ n3049);
assign n3128 = ~(n9339 ^ n4763);
assign n10184 = ~(n11232 | n8064);
assign n10041 = ~(n349 ^ n3520);
assign n6812 = ~(n8522 | n3882);
assign n6370 = n12119 | n12535;
assign n9820 = ~(n1264 ^ n4776);
assign n4785 = n9379 | n1356;
assign n851 = ~(n12327 ^ n1660);
assign n5231 = n8583 | n4875;
assign n812 = ~(n6175 ^ n11006);
assign n1562 = ~n3928;
assign n2285 = n752 | n9741;
assign n11245 = n11026 | n3606;
assign n11010 = ~(n7243 ^ n2460);
assign n7095 = ~(n8904 ^ n12193);
assign n9651 = n4911 | n5497;
assign n11948 = n9029 & n2615;
assign n6450 = n1016 | n1979;
assign n3375 = ~(n12532 ^ n1620);
assign n11896 = ~n5105;
assign n7657 = ~n1216;
assign n9028 = ~n9655;
assign n2073 = ~(n4224 ^ n7155);
assign n8830 = ~n7294;
assign n689 = ~(n1255 ^ n10444);
assign n3948 = ~n3519;
assign n12748 = ~n11050;
assign n9732 = n3795 | n10294;
assign n4810 = ~(n1475 ^ n5414);
assign n6124 = ~n1505;
assign n1450 = ~(n9089 ^ n11980);
assign n7402 = ~(n5832 ^ n6531);
assign n10813 = n681 & n10418;
assign n373 = ~n3921;
assign n10115 = ~(n1721 ^ n10114);
assign n12649 = ~(n7375 ^ n5256);
assign n917 = n7588 & n9543;
assign n6234 = ~n5299;
assign n7075 = ~(n3337 ^ n3294);
assign n8042 = n3642 & n10963;
assign n5336 = ~(n5432 ^ n12292);
assign n11126 = n8835 | n9595;
assign n8958 = n7218 & n4313;
assign n8839 = n11958 | n11410;
assign n3207 = n6635 | n9863;
assign n5393 = n11958 | n3468;
assign n6747 = ~n11038;
assign n8972 = ~(n9988 | n6332);
assign n6105 = n11953 | n11242;
assign n4741 = ~(n3869 ^ n6209);
assign n11419 = ~(n6374 | n5757);
assign n6153 = n3096 | n7558;
assign n11822 = n4480 | n7866;
assign n603 = ~(n9499 | n17);
assign n1013 = ~(n4142 | n4691);
assign n10945 = n6718 | n3606;
assign n2842 = n6786 & n10373;
assign n12261 = n432 | n9549;
assign n3787 = ~(n2193 ^ n4708);
assign n3393 = n5547 | n5810;
assign n8520 = ~(n3883 ^ n5807);
assign n10769 = ~(n1390 ^ n1292);
assign n6021 = n6772 | n1596;
assign n7701 = n5285 & n6902;
assign n3991 = n7657 & n9315;
assign n2225 = ~(n9164 | n6802);
assign n5784 = ~(n12799 ^ n12253);
assign n1956 = n11627 & n7205;
assign n575 = ~(n102 | n5875);
assign n873 = n12090 | n4871;
assign n12588 = n5319 & n9763;
assign n12790 = n12115 & n1761;
assign n11740 = n1419 | n9216;
assign n214 = n2947 & n940;
assign n841 = ~(n5370 ^ n339);
assign n5967 = n11026 | n8643;
assign n6657 = ~(n3412 | n12407);
assign n9212 = n12941 | n1624;
assign n1663 = n10219 | n7477;
assign n5475 = ~(n11264 ^ n3744);
assign n11466 = ~(n3198 | n12772);
assign n6851 = n1900 | n9556;
assign n12698 = n5247 & n9020;
assign n7993 = n7236 & n9111;
assign n9851 = ~(n6313 ^ n498);
assign n3045 = ~(n12950 | n1381);
assign n2072 = n97 | n2129;
assign n4975 = ~(n4138 ^ n9929);
assign n4724 = n9101 & n9516;
assign n1654 = n11719 | n1455;
assign n2948 = ~(n2075 | n6972);
assign n100 = ~(n11184 ^ n11018);
assign n10449 = ~n6997;
assign n5856 = ~(n5324 ^ n518);
assign n4108 = n2069 & n10458;
assign n2766 = ~n5627;
assign n10751 = n1200 | n1482;
assign n9822 = n3700 & n5294;
assign n10904 = n6867 & n187;
assign n1694 = ~(n11929 ^ n6253);
assign n4966 = n11319 | n4310;
assign n3492 = ~(n5605 ^ n3745);
assign n9765 = n8645 & n9594;
assign n3404 = ~(n6576 ^ n5150);
assign n4177 = ~n6705;
assign n1646 = n8959 | n11896;
assign n12954 = ~n11708;
assign n9090 = n5945 | n11775;
assign n11060 = n7283 | n1546;
assign n8916 = n10339 | n5468;
assign n10136 = n7409 | n1868;
assign n419 = n12038 | n1913;
assign n5888 = ~(n6070 ^ n56);
assign n12771 = ~n9111;
assign n11676 = ~(n6190 ^ n11658);
assign n6476 = ~(n4647 ^ n11236);
assign n3840 = n12750 & n376;
assign n7440 = n5916 & n6785;
assign n5885 = n114 | n6169;
assign n12343 = n4189 & n4370;
assign n8501 = ~(n737 ^ n6132);
assign n8445 = n1316 | n6898;
assign n2805 = n12135 & n1380;
assign n9366 = ~(n1275 ^ n8240);
assign n4437 = n8823 & n2049;
assign n10913 = ~(n10857 ^ n8385);
assign n8073 = ~n6498;
assign n278 = ~(n458 ^ n2992);
assign n8068 = ~(n3340 ^ n4228);
assign n10392 = n8839 | n10927;
assign n11283 = ~(n5213 | n12602);
assign n5512 = n807 | n2232;
assign n2315 = ~(n1359 | n6658);
assign n9197 = ~(n3076 ^ n7402);
assign n6080 = n2541 & n10427;
assign n1457 = ~(n663 ^ n9039);
assign n11899 = ~(n8165 | n297);
assign n3571 = ~n1426;
assign n1484 = n2967 | n10447;
assign n2408 = n8759 & n3602;
assign n3406 = n9538 | n4064;
assign n7209 = n1741 | n8715;
assign n9049 = n12388 & n2492;
assign n10634 = ~n5336;
assign n11851 = n7283 | n2358;
assign n11723 = ~(n1518 ^ n3536);
assign n8940 = n10247 | n5597;
assign n9067 = n4255 & n10411;
assign n5853 = n686 | n7952;
assign n1195 = ~(n1043 ^ n4780);
assign n9469 = ~(n8752 ^ n9850);
assign n9029 = n4639 | n6140;
assign n7697 = ~(n10039 ^ n5591);
assign n7991 = ~(n12859 ^ n2652);
assign n4607 = ~(n8266 ^ n2102);
assign n6042 = ~n5533;
assign n3266 = n3573 | n10624;
assign n2867 = n11059 | n12300;
assign n6134 = n10626 & n12317;
assign n2344 = n621 & n6844;
assign n6362 = ~n1541;
assign n10593 = ~(n5603 ^ n11345);
assign n10677 = n2534 & n4747;
assign n8430 = n1465 | n6272;
assign n7406 = n8136 | n4879;
assign n9449 = ~(n3546 | n9225);
assign n1634 = n5685 & n5658;
assign n12466 = n11717 & n9120;
assign n9657 = n7974 & n9532;
assign n11248 = n11460 ^ n39;
assign n5923 = n5214 | n2616;
assign n3587 = ~(n8334 | n6234);
assign n9431 = n10799 | n917;
assign n6296 = n10142 | n8735;
assign n2668 = ~n8121;
assign n11487 = n422 | n12482;
assign n10716 = ~n146;
assign n1454 = n1627 & n5813;
assign n5656 = n2700 & n3268;
assign n10709 = ~n9708;
assign n5126 = n4451 & n1852;
assign n7059 = ~(n1477 | n11049);
assign n5605 = n5530 | n2964;
assign n7729 = n11305 & n10501;
assign n1031 = ~(n11687 ^ n6599);
assign n7738 = ~(n12107 ^ n6632);
assign n12651 = ~(n9985 ^ n5777);
assign n7908 = n2564 & n7265;
assign n4425 = ~n2973;
assign n8618 = n3887 & n3583;
assign n5737 = n6226 | n7666;
assign n47 = ~n2085;
assign n6943 = n7015 | n9959;
assign n12654 = ~(n8510 ^ n8274);
assign n9273 = n5341 | n11947;
assign n1233 = ~n11280;
assign n8403 = ~(n7299 ^ n2239);
assign n12253 = n5945 | n7952;
assign n10332 = ~n6379;
assign n5413 = n9233 & n8244;
assign n12710 = ~(n2014 ^ n12259);
assign n2465 = n7376 & n7465;
assign n12823 = n8738 | n9568;
assign n5777 = n9507 | n1602;
assign n8861 = ~(n431 ^ n8546);
assign n11237 = ~(n531 ^ n1338);
assign n5895 = n9400 & n12145;
assign n711 = ~n12776;
assign n5572 = ~(n4458 ^ n9783);
assign n74 = n6465 & n4645;
assign n4281 = n2699 & n1618;
assign n7635 = ~(n11932 ^ n8841);
assign n7851 = n7839 | n2232;
assign n5399 = n3878 & n1565;
assign n5591 = ~(n10291 | n11261);
assign n5122 = ~(n10699 ^ n5490);
assign n2726 = n11026 | n9521;
assign n5848 = n12237 | n12080;
assign n8527 = ~(n8149 | n5517);
assign n3483 = ~(n121 ^ n1389);
assign n668 = n6339 | n3157;
assign n1679 = n5673 | n8756;
assign n4240 = ~(n9322 ^ n3475);
assign n11796 = n11153 & n159;
assign n5761 = n3127 | n4400;
assign n3653 = n8583 | n795;
assign n2860 = n5340 & n11957;
assign n756 = n8273 & n4909;
assign n9237 = ~n4105;
assign n1957 = ~n11358;
assign n4444 = ~(n8535 ^ n2410);
assign n12165 = n4778 | n8655;
assign n2535 = n9880 & n10801;
assign n116 = n12195 | n4622;
assign n9073 = n12186 | n7876;
assign n7479 = n10748 | n2039;
assign n7702 = n8046 | n4497;
assign n6970 = ~(n4206 ^ n4303);
assign n3322 = ~n7267;
assign n8973 = n6482 & n4586;
assign n399 = n5754 & n1983;
assign n11306 = ~(n11718 ^ n350);
assign n5301 = n8342 & n4051;
assign n5930 = n4812 & n2573;
assign n4906 = n1220 & n12621;
assign n7363 = n4289 | n3035;
assign n7397 = ~n5003;
assign n2959 = ~n12178;
assign n2038 = ~(n583 ^ n6202);
assign n3877 = ~(n7416 ^ n950);
assign n4174 = ~(n1916 ^ n655);
assign n8448 = ~(n4158 | n4407);
assign n9268 = ~(n5728 | n6335);
assign n4761 = ~(n10361 ^ n12246);
assign n12474 = ~(n862 | n8121);
assign n12031 = n2464 & n8595;
assign n1434 = ~(n4577 | n10423);
assign n2776 = ~(n9832 ^ n8657);
assign n8238 = n6076 & n5169;
assign n7281 = ~(n12871 | n5649);
assign n5253 = ~(n5109 | n12295);
assign n3217 = ~(n12639 ^ n9823);
assign n11805 = n3931 | n9720;
assign n12438 = n4624 & n8281;
assign n12641 = ~(n1867 ^ n8734);
assign n2105 = n92 & n4789;
assign n6103 = n10842 | n5823;
assign n7005 = n3382 & n8620;
assign n203 = n1910 & n3114;
assign n8080 = ~(n6773 | n9419);
assign n535 = n5771 & n415;
assign n7196 = n4562 & n12689;
assign n12807 = ~(n310 ^ n3008);
assign n5929 = ~n6136;
assign n4439 = n1345 & n6887;
assign n10598 = n12280 & n2937;
assign n10938 = ~n3016;
assign n6795 = n4023 | n1870;
assign n3851 = ~(n8894 ^ n11774);
assign n12639 = ~(n9936 | n2634);
assign n12486 = ~(n7798 | n2194);
assign n9498 = n10862 | n10421;
assign n1268 = ~(n5590 ^ n12406);
assign n4251 = ~(n8229 ^ n1276);
assign n6529 = n7468 & n271;
assign n11510 = ~(n6541 | n1219);
assign n5232 = ~(n925 ^ n10714);
assign n7650 = ~(n10000 ^ n6912);
assign n11197 = n12775 & n12913;
assign n10062 = ~(n2602 ^ n2106);
assign n7433 = n2483 & n4040;
assign n11675 = n7449 | n8285;
assign n7549 = n8583 | n9078;
assign n6236 = ~(n10438 ^ n12160);
assign n12518 = n12659 | n6846;
assign n1684 = n3767 | n7600;
assign n2460 = n4693 & n5182;
assign n2009 = ~(n7102 ^ n7017);
assign n10262 = ~(n12747 ^ n8685);
assign n9187 = ~(n9770 ^ n2556);
assign n5531 = n3992 & n10990;
assign n977 = ~(n10367 ^ n2164);
assign n190 = n8929 & n11141;
assign n7671 = ~(n10711 ^ n6094);
assign n2362 = ~(n6886 | n8213);
assign n5161 = ~(n9629 ^ n11870);
assign n5995 = n10157 | n9280;
assign n10835 = ~n7965;
assign n7240 = n6442 & n10619;
assign n9924 = n2959 & n1481;
assign n2200 = ~(n5026 ^ n4539);
assign n641 = ~n12071;
assign n6518 = n6718 | n9078;
assign n10695 = ~(n6665 ^ n8726);
assign n2782 = n3402 | n3391;
assign n12804 = ~(n12433 | n5417);
assign n8122 = ~(n12242 ^ n8909);
assign n7369 = n6022 | n8427;
assign n10983 = n9370 | n7424;
assign n12939 = ~(n10700 ^ n7435);
assign n7145 = n4498 | n7703;
assign n6041 = ~(n4635 | n12369);
assign n777 = ~(n3726 | n8031);
assign n12719 = n307 & n3471;
assign n5407 = n8687 | n9521;
assign n788 = ~(n10343 ^ n9535);
assign n925 = n8187 | n1079;
assign n5826 = n1205 | n4282;
assign n7842 = ~(n12945 ^ n9859);
assign n8370 = n7780 & n8901;
assign n2317 = ~n8144;
assign n10858 = ~(n10365 ^ n8512);
assign n9574 = ~(n8130 ^ n9284);
assign n7921 = ~n5814;
assign n4440 = ~(n7188 ^ n10807);
assign n2168 = n2326 | n10869;
assign n7911 = ~(n11972 ^ n11732);
assign n197 = ~(n12012 ^ n3054);
assign n7077 = n9900 | n5063;
assign n5249 = n9844 | n7976;
assign n10163 = n5372 | n4163;
assign n12152 = ~(n3188 ^ n5561);
assign n10270 = ~n1354;
assign n12936 = n4126 | n12608;
assign n8637 = n10715 | n5316;
assign n4133 = ~(n578 ^ n8938);
assign n10911 = n5774 | n10011;
assign n12531 = ~n1837;
assign n1495 = n1941 | n7558;
assign n10498 = n5141 & n545;
assign n587 = n505 | n12592;
assign n8411 = n6204 | n11735;
assign n7494 = n5981 & n5661;
assign n5327 = n7476 & n10942;
assign n4059 = ~n1097;
assign n12047 = n12297 & n11611;
assign n3417 = ~(n8733 | n5632);
assign n12764 = n8476 & n6806;
assign n9492 = n6977 | n995;
assign n81 = ~n3205;
assign n4562 = n3746 | n7558;
assign n8275 = ~(n8369 ^ n4284);
assign n8629 = ~n10231;
assign n2560 = n3352 & n1765;
assign n8418 = n9996 & n6634;
assign n5908 = n7709 | n1509;
assign n6005 = ~(n10335 | n2378);
assign n7152 = ~(n6003 ^ n2919);
assign n11460 = n10045 & n6345;
assign n1760 = n12067 & n9214;
assign n4944 = ~(n7300 | n9252);
assign n10647 = n5465 & n6783;
assign n11067 = ~(n2877 ^ n7973);
assign n23 = n1519 & n564;
assign n801 = ~(n1207 ^ n10696);
assign n842 = ~(n8998 ^ n8575);
assign n10028 = ~(n1516 ^ n2181);
assign n10546 = n12023 & n7734;
assign n5356 = ~(n12282 ^ n4631);
assign n2547 = ~(n12728 ^ n340);
assign n1276 = n636 | n10854;
assign n4033 = ~(n10921 | n7522);
assign n240 = n2217 | n9078;
assign n3397 = ~n7735;
assign n12626 = n7283 | n6389;
assign n1605 = n8228 | n956;
assign n5053 = n8336 & n7946;
assign n8017 = ~(n5280 | n1801);
assign n10009 = ~(n3313 ^ n11809);
assign n5209 = n1349 | n8258;
assign n6614 = ~(n451 ^ n9502);
assign n8223 = ~(n5148 | n6675);
assign n5934 = ~(n917 ^ n7262);
assign n12359 = n8074 & n735;
assign n1327 = n6674 & n7075;
assign n5052 = ~(n12667 ^ n11737);
assign n2662 = ~(n1792 ^ n8636);
assign n7035 = n12503 | n795;
assign n7153 = n8764 | n8918;
assign n9581 = n11473 & n6925;
assign n7201 = ~(n4863 ^ n7145);
assign n11269 = ~(n9746 | n6586);
assign n2540 = ~(n9791 ^ n7905);
assign n3791 = n10142 | n7246;
assign n12421 = n77 & n8056;
assign n5955 = n3605 & n9888;
assign n4315 = ~(n2586 ^ n2486);
assign n9219 = n1076 | n3439;
assign n3982 = ~(n6597 ^ n6845);
assign n10883 = n2031 & n650;
assign n10950 = ~(n9656 ^ n12411);
assign n10282 = n5769 | n7239;
assign n1555 = ~(n7838 ^ n9135);
assign n9100 = n11697 | n2985;
assign n6718 = ~n8384;
assign n6829 = ~(n9508 | n146);
assign n183 = n11958 | n7395;
assign n8825 = ~(n6330 ^ n6996);
assign n8813 = n7376 | n7465;
assign n6544 = n9373 | n795;
assign n3798 = ~(n12789 | n2355);
assign n1879 = n11433 | n5012;
assign n8687 = ~n5857;
assign n9156 = ~(n3944 ^ n1719);
assign n3052 = ~(n11079 | n3847);
assign n3501 = ~n927;
assign n5708 = ~(n290 ^ n4551);
assign n8522 = n7778 & n7276;
assign n8837 = ~n2921;
assign n7015 = ~n6891;
assign n7195 = n10966 | n7447;
assign n9015 = ~n5846;
assign n8113 = ~n8556;
assign n7799 = ~(n10912 ^ n6143);
assign n10555 = n2217 | n11698;
assign n10820 = n4778 | n12080;
assign n9724 = ~n6343;
assign n4077 = ~(n852 | n8335);
assign n563 = ~n8927;
assign n1648 = n3478 & n1104;
assign n10700 = ~(n1307 ^ n3239);
assign n9209 = ~(n11544 ^ n5944);
assign n855 = n7116 | n9741;
assign n3072 = n636 | n8655;
assign n12387 = ~(n4416 ^ n4253);
assign n6197 = ~n8595;
assign n7344 = n9066 & n11894;
assign n7365 = n636 | n7928;
assign n9427 = ~(n3222 | n12228);
assign n749 = ~(n7253 | n12848);
assign n11645 = ~n5808;
assign n9374 = n11433 | n995;
assign n10226 = ~n8851;
assign n8467 = n8410 | n6101;
assign n10233 = ~(n4759 | n1569);
assign n7364 = n6559 & n2977;
assign n785 = n3665 & n2452;
assign n4402 = ~(n11591 | n9841);
assign n2987 = n10847 | n12626;
assign n2702 = ~(n8381 | n3163);
assign n4273 = ~(n10529 ^ n626);
assign n12210 = n5081 & n3953;
assign n10257 = ~n3795;
assign n1407 = n4247 & n554;
assign n8082 = ~n1408;
assign n10921 = n10947 & n11800;
assign n7618 = n8209 | n160;
assign n9969 = ~(n5129 | n11770);
assign n4062 = n6115 & n1566;
assign n11737 = ~(n10306 ^ n1042);
assign n5514 = n4296 | n11865;
assign n4494 = ~(n5567 ^ n4959);
assign n7156 = n338 | n11885;
assign n8935 = ~(n333 ^ n2955);
assign n12001 = n3627 & n9956;
assign n7047 = ~(n1726 ^ n3718);
assign n6109 = n7487 & n7752;
assign n8014 = ~(n8628 ^ n12625);
assign n12537 = ~(n1837 ^ n5565);
assign n12846 = n1699 | n6513;
assign n4999 = ~(n1588 ^ n12677);
assign n1853 = ~(n3576 ^ n6403);
assign n12196 = ~(n3516 | n11845);
assign n889 = ~n4697;
assign n7588 = n7758 | n1861;
assign n1721 = ~(n6229 ^ n3473);
assign n1723 = n3445 & n10261;
assign n11489 = n10661 & n5276;
assign n12109 = ~(n9989 | n10408);
assign n4950 = n7071 | n8338;
assign n8131 = ~(n11242 ^ n3597);
assign n2057 = ~(n5987 ^ n8723);
assign n10181 = n12335 & n9743;
assign n10804 = n9584 | n4527;
assign n2361 = ~(n4564 | n4487);
assign n6931 = n5765 | n3606;
assign n12154 = ~(n11219 ^ n4800);
assign n6459 = ~(n7267 ^ n11797);
assign n8664 = ~(n2855 ^ n8874);
assign n9509 = ~(n8208 ^ n5512);
assign n9486 = ~n6423;
assign n8630 = n2600 & n12332;
assign n8799 = n9838 & n11645;
assign n11027 = n8489 & n5696;
assign n4287 = n7638 | n7419;
assign n2158 = ~(n6896 ^ n7636);
assign n412 = n8584 | n12605;
assign n10165 = ~(n6116 ^ n4188);
assign n9010 = n3992 & n6611;
assign n2711 = n12443 | n1734;
assign n12632 = n7397 & n11166;
assign n3823 = n7577 | n5796;
assign n7117 = n6373 | n12771;
assign n4404 = ~(n928 ^ n3650);
assign n4135 = n5778 & n1591;
assign n10037 = ~(n12057 ^ n654);
assign n404 = n373 | n10191;
assign n11945 = ~(n12854 ^ n7589);
assign n8558 = n5951 | n5678;
assign n9272 = ~n604;
assign n12357 = ~n4190;
assign n3132 = ~(n10864 ^ n4198);
assign n4283 = n8428 | n995;
assign n11250 = n8428 | n3468;
assign n8374 = ~(n12692 ^ n11882);
assign n2397 = ~(n6561 ^ n10705);
assign n3685 = n7393 & n12362;
assign n1728 = n9792 & n7554;
assign n12012 = n740 & n406;
assign n2978 = n5809 | n8740;
assign n972 = n10928 & n3719;
assign n12159 = ~(n6405 ^ n7440);
assign n5170 = n3544 & n4715;
assign n10652 = n6718 | n1509;
assign n10896 = n5765 | n1509;
assign n10432 = ~(n7457 | n872);
assign n2482 = n12119 | n10311;
assign n1845 = n713 & n96;
assign n8667 = ~(n650 ^ n2031);
assign n10376 = ~n12880;
assign n11529 = ~(n10199 ^ n7637);
assign n3202 = n10750 | n7928;
assign n4931 = n8189 | n5797;
assign n11359 = ~(n9697 | n1778);
assign n2745 = ~(n5219 ^ n3461);
assign n11135 = ~n8467;
assign n6284 = n2659 | n3186;
assign n7023 = n3401 & n1996;
assign n9845 = ~(n12760 | n2199);
assign n6447 = ~(n7866 ^ n2115);
assign n9966 = ~(n9068 ^ n9871);
assign n5936 = n12584 & n5733;
assign n12341 = n8789 & n1733;
assign n10131 = ~(n2172 ^ n11897);
assign n11910 = n10750 | n10854;
assign n8986 = ~(n8896 | n4710);
assign n5111 = n697 | n1109;
assign n5110 = n12380 & n4985;
assign n931 = ~(n269 | n10924);
assign n4104 = ~n5652;
assign n5921 = ~(n8469 ^ n2617);
assign n8677 = ~(n11578 ^ n975);
assign n4399 = ~(n12266 ^ n2438);
assign n10771 = n11552 | n4527;
assign n2896 = n9262 | n2020;
assign n5183 = n1339 | n8940;
assign n3213 = ~n7993;
assign n10336 = n6358 & n11791;
assign n9778 = n7993 & n5845;
assign n12788 = ~(n1520 ^ n8247);
assign n7074 = n7236 & n10848;
assign n6922 = ~n12247;
assign n9836 = n5575 | n3421;
assign n1770 = ~(n8079 ^ n741);
assign n1453 = ~(n9555 ^ n10550);
assign n4791 = n7283 | n7703;
assign n12676 = ~(n11287 ^ n11954);
assign n10565 = n6373 | n9160;
assign n6051 = ~(n12718 ^ n234);
assign n11072 = ~n11783;
assign n11406 = n12361 | n11775;
assign n2682 = n3141 & n4721;
assign n1206 = ~(n902 ^ n5829);
assign n8672 = n2941 & n1567;
assign n10765 = ~(n11445 ^ n247);
assign n3936 = n11026 | n5502;
assign n6700 = n11607 | n10719;
assign n6423 = ~(n7206 ^ n11655);
assign n6918 = ~(n6628 ^ n1424);
assign n5197 = ~(n8996 ^ n4053);
assign n10103 = n4791 | n5762;
assign n9382 = n4411 & n10007;
assign n3850 = ~(n409 ^ n12094);
assign n9031 = n12842 & n5654;
assign n8652 = ~(n8979 ^ n4334);
assign n3081 = n6695 | n6006;
assign n1559 = ~n2752;
assign n8012 = ~(n11366 | n7237);
assign n5672 = ~(n12024 | n8821);
assign n8602 = ~(n4385 ^ n7266);
assign n1773 = n7540 | n3055;
assign n12730 = n11887 | n7382;
assign n612 = ~(n11369 | n2990);
assign n1171 = ~n10788;
assign n7624 = ~(n5898 | n633);
assign n10396 = ~n3579;
assign n7141 = n1784 | n11355;
assign n3570 = n5575 | n3356;
assign n532 = ~(n1912 ^ n2546);
assign n5044 = ~n1397;
assign n960 = n2987 & n6214;
assign n4924 = ~n2180;
assign n12796 = n7316 & n9090;
assign n17 = ~n4923;
assign n7332 = ~(n225 ^ n8039);
assign n12903 = ~(n5441 ^ n1862);
assign n4536 = n2456 | n4818;
assign n1632 = n2532 & n4802;
assign n12884 = ~(n5799 ^ n801);
assign n5202 = n6577 | n11410;
assign n12144 = n5530 | n1932;
assign n4815 = n9878 | n9188;
assign n10004 = n10282 & n3409;
assign n12657 = ~(n9029 ^ n3500);
assign n2746 = ~(n7516 ^ n3809);
assign n11040 = n9241 & n6703;
assign n6981 = n5765 | n11698;
assign n3631 = n4343 | n826;
assign n4911 = ~n12705;
assign n3443 = ~(n11348 ^ n472);
assign n3286 = n10365 & n10723;
assign n2677 = n5575 | n7425;
assign n9737 = n3325 & n1386;
assign n432 = n2217 | n4875;
assign n8882 = n5915 | n10854;
assign n4316 = ~(n1256 | n3254);
assign n12551 = n1403 & n765;
assign n12319 = ~(n5965 ^ n169);
assign n12501 = ~n2111;
assign n10438 = n7197 | n8069;
assign n12640 = ~n3732;
assign n69 = n1438 | n2409;
assign n7961 = n4716 | n7;
assign n9423 = ~(n11838 ^ n7344);
assign n3810 = n12237 | n7382;
assign n7945 = n7807 & n1412;
assign n1612 = ~n2519;
assign n10356 = n595 | n9449;
assign n12053 = n4059 | n7341;
assign n8452 = n6373 | n9568;
assign n11325 = ~(n4771 ^ n5082);
assign n4765 = ~(n11961 | n1090);
assign n3967 = n8552 | n826;
assign n1595 = n10180 & n4234;
assign n12130 = ~n6725;
assign n964 = n8687 | n9160;
assign n12825 = n11282 | n3517;
assign n6541 = n1018 & n6093;
assign n12713 = ~(n9115 ^ n11924);
assign n1202 = ~(n8857 ^ n7842);
assign n7660 = ~(n4819 | n10515);
assign n9264 = ~(n3198 ^ n7596);
assign n9142 = ~n7027;
assign n7859 = n5971 | n8824;
assign n3149 = ~(n4535 ^ n501);
assign n1609 = ~(n2109 ^ n859);
assign n9327 = ~n3990;
assign n3231 = n6130 & n6708;
assign n10429 = n10673 & n8926;
assign n12950 = n12210 & n601;
assign n1874 = n5765 | n4864;
assign n3148 = ~(n10798 ^ n10707);
assign n616 = n7284 | n10144;
assign n671 = ~(n10853 ^ n11300);
assign n2086 = ~(n553 ^ n4133);
assign n5024 = n11026 | n4474;
assign n11107 = ~(n202 | n9086);
assign n6869 = n5110 | n2795;
assign n7584 = n9304 | n8148;
assign n315 = n5664 | n2145;
assign n1401 = n2154 | n6459;
assign n9243 = ~n11225;
assign n3861 = n1891 | n11920;
assign n1212 = n1960 | n1019;
assign n3297 = n9370 | n6402;
assign n3300 = n8405 | n9188;
assign n12046 = n8870 | n8648;
assign n9496 = n8687 | n4474;
assign n6471 = n11598 | n5096;
assign n9681 = n5348 | n581;
assign n4006 = ~(n2937 ^ n1297);
assign n9338 = ~(n11968 ^ n6);
assign n5893 = n6221 | n9851;
assign n3578 = ~n3003;
assign n12745 = ~n9381;
assign n10475 = ~n10394;
assign n856 = n6977 | n10919;
assign n12524 = n3617 | n6513;
assign n3777 = n11032 | n12830;
assign n9834 = n1937 | n11820;
assign n6502 = ~(n11937 ^ n1547);
assign n6989 = ~(n100 ^ n12100);
assign n4632 = n3494 & n2646;
assign n8749 = ~n1304;
assign n11275 = n9858 & n10972;
assign n12554 = n5602 | n2463;
assign n4247 = n7449 | n8830;
assign n5965 = ~(n1010 ^ n5187);
assign n8509 = ~n2533;
assign n10224 = n4535 | n501;
assign n9119 = n12324 | n2736;
assign n8402 = ~(n730 ^ n4345);
assign n499 = n9093 & n5682;
assign n7520 = n9886 & n3370;
assign n155 = ~(n2826 ^ n758);
assign n7515 = ~(n6365 ^ n9702);
assign n9034 = ~(n6512 | n12681);
assign n4643 = ~n8580;
assign n9096 = ~(n946 ^ n3258);
assign n6187 = ~(n8339 ^ n9540);
assign n225 = ~(n8448 ^ n10161);
assign n1700 = ~n3531;
assign n2099 = ~n5331;
assign n4100 = ~n12582;
assign n4853 = ~n8324;
assign n4009 = ~(n6813 ^ n4156);
assign n10504 = n5575 | n7395;
assign n2525 = n12361 | n12816;
assign n9048 = n7116 | n7952;
assign n9907 = n8750 & n10537;
assign n3115 = ~n1017;
assign n5151 = n10118 | n5887;
assign n7448 = ~(n8044 | n8319);
assign n6453 = ~(n10008 ^ n8494);
assign n3989 = ~n11563;
assign n7642 = n2407 | n12137;
assign n5270 = ~(n7953 ^ n12148);
assign n5078 = ~(n7531 ^ n9259);
assign n7414 = n10677 | n5079;
assign n12390 = n1169 | n4891;
assign n6062 = n7984 | n1541;
assign n1414 = ~(n5260 ^ n1108);
assign n2996 = ~(n2120 ^ n12885);
assign n5538 = ~n4141;
assign n11698 = ~n4903;
assign n6460 = n1534 & n8112;
assign n8951 = ~n1646;
assign n4434 = ~n12723;
assign n4728 = n5575 | n7558;
assign n5354 = n4568 | n12558;
assign n11527 = ~(n1456 ^ n8842);
assign n3938 = n12633 | n6508;
assign n326 = n5989 | n6704;
assign n6828 = ~(n12430 | n6281);
assign n8698 = n4422 | n12809;
assign n11688 = n5619 & n7308;
assign n7048 = ~(n7474 ^ n7654);
assign n12364 = ~(n2536 ^ n2670);
assign n2420 = n2011 & n4899;
assign n11659 = n8304 & n10469;
assign n6239 = n11958 | n6455;
assign n6399 = ~(n8781 | n4330);
assign n3254 = n2506 & n11807;
assign n3583 = n7384 | n2005;
assign n11976 = ~n6303;
assign n105 = n11037 & n10573;
assign n7795 = n8510 & n8274;
assign n11420 = n10202 & n9729;
assign n3834 = n5419 & n11619;
assign n11656 = n3176 & n8167;
assign n6357 = ~(n9414 ^ n2038);
assign n7319 = n9081 | n6258;
assign n12450 = ~(n8304 ^ n190);
assign n7780 = n10761 | n3234;
assign n4585 = n4725 | n12396;
assign n6924 = n10750 | n7382;
assign n1344 = ~n165;
assign n10221 = ~(n8436 ^ n86);
assign n4150 = n11694 | n4377;
assign n12927 = ~(n6566 | n4542);
assign n483 = n9621 | n1490;
assign n652 = ~(n4962 ^ n10016);
assign n642 = ~(n296 ^ n6837);
assign n952 = ~(n9134 ^ n5775);
assign n7066 = ~(n6659 ^ n7524);
assign n10687 = ~(n9445 ^ n4567);
assign n6400 = ~(n474 ^ n1556);
assign n3230 = ~(n12359 ^ n94);
assign n2231 = n8730 & n5588;
assign n7988 = ~(n5881 ^ n9979);
assign n4169 = ~n11628;
assign n6295 = n8838 | n8029;
assign n7770 = n5600 | n2793;
assign n984 = ~(n6076 | n5169);
assign n3712 = ~n5495;
assign n4571 = n955 | n5442;
assign n1828 = n4956 & n5000;
assign n6352 = n6290 | n11439;
assign n3454 = ~(n12422 | n8568);
assign n9128 = ~(n2532 | n4802);
assign n10895 = n3065 & n577;
assign n2137 = n11417 | n1314;
assign n11597 = n10101 | n2218;
assign n1858 = ~(n9969 ^ n7604);
assign n2815 = ~n7946;
assign n5332 = ~(n3608 ^ n11467);
assign n10626 = n11037 | n10573;
assign n4548 = n10564 | n9733;
assign n4560 = n11390 | n3431;
assign n9409 = ~(n4536 ^ n4220);
assign n7329 = n7404 & n11438;
assign n3841 = n5913 | n2751;
assign n11393 = ~(n9942 ^ n2477);
assign n3788 = ~(n8557 | n7653);
assign n5763 = ~n12115;
assign n1122 = ~n2413;
assign n1862 = n1699 | n8740;
assign n2768 = n11621 & n11956;
assign n1739 = ~n6431;
assign n4996 = ~(n1960 ^ n1019);
assign n3355 = ~(n11992 | n1293);
assign n2410 = ~(n195 ^ n12049);
assign n12878 = ~n2038;
assign n131 = n11601 | n10724;
assign n4482 = n7474 & n1681;
assign n4398 = n3549 & n98;
assign n6733 = ~(n1804 ^ n1105);
assign n8381 = ~(n5202 ^ n12240);
assign n4423 = ~n302;
assign n3714 = ~n1716;
assign n4126 = n11958 | n10919;
assign n5410 = ~n8940;
assign n12702 = ~(n8864 ^ n8788);
assign n3908 = n3891 | n8409;
assign n11517 = n11958 | n12357;
assign n2762 = ~n11553;
assign n10149 = ~(n7248 | n12159);
assign n77 = n8227 | n10209;
assign n4282 = n12195 & n4622;
assign n1430 = ~(n4910 ^ n4361);
assign n2182 = n994 | n2076;
assign n12015 = n686 | n5012;
assign n4532 = n2078 | n10596;
assign n7843 = n12632 | n10244;
assign n7202 = n2626 | n4041;
assign n6034 = n2288 & n1145;
assign n10859 = ~(n9744 ^ n3963);
assign n8203 = n9748 & n10395;
assign n4563 = ~(n3463 | n8178);
assign n7756 = n4498 | n1851;
assign n10277 = ~(n8277 | n12370);
assign n7168 = n6595 | n6639;
assign n364 = ~(n3551 ^ n12205);
assign n4227 = ~(n3210 ^ n11192);
assign n5123 = ~(n2155 ^ n5786);
assign n8311 = n4768 | n9619;
assign n2206 = ~(n5618 ^ n1430);
assign n5762 = ~(n12913 ^ n12239);
assign n11817 = ~(n3106 | n11945);
assign n8807 = ~n3465;
assign n5023 = n674 & n10606;
assign n401 = n10852 | n12019;
assign n10162 = n2756 | n327;
assign n11990 = n8984 & n12268;
assign n4216 = ~n4275;
assign n2041 = n12157 | n11197;
assign n10514 = ~n10711;
assign n7764 = n12503 | n4654;
assign n7305 = n6242 & n8791;
assign n8679 = n2526 | n8491;
assign n10193 = n705 & n1310;
assign n10558 = ~(n12880 ^ n2690);
assign n7848 = ~(n8713 | n6850);
assign n5792 = n4932 & n12548;
assign n2567 = ~(n2686 ^ n10618);
assign n8252 = ~(n8011 ^ n10518);
assign n1488 = ~n11227;
assign n8435 = n4637 & n11288;
assign n2748 = ~n5916;
assign n6449 = ~(n5177 | n10438);
assign n10775 = n677 & n7811;
assign n8491 = ~(n6258 ^ n12412);
assign n9787 = n11026 | n2020;
assign n2235 = ~(n9109 ^ n6207);
assign n9084 = ~(n1961 ^ n6791);
assign n8796 = ~n3179;
assign n1920 = n1266 | n2090;
assign n8261 = n3126 & n188;
assign n12905 = n7998 & n4153;
assign n8722 = ~n9541;
assign n8593 = ~(n5024 ^ n5255);
assign n1489 = n3050 & n11524;
assign n11566 = ~(n7572 ^ n7394);
assign n5954 = ~n5967;
assign n11030 = ~(n7761 ^ n3259);
assign n2011 = n4628 | n12754;
assign n5685 = n3743 | n9144;
assign n8083 = n1471 & n8433;
assign n638 = n12119 | n530;
assign n991 = n5530 | n7382;
assign n4829 = ~(n7148 ^ n8106);
assign n12781 = n5575 | n12274;
assign n4380 = n10142 | n7703;
assign n913 = n6977 | n11122;
assign n9121 = ~(n597 ^ n1289);
assign n12879 = n1051 | n11820;
assign n4064 = n6534 & n10826;
assign n11024 = n8127 | n4400;
assign n12561 = n12669 | n6360;
assign n12946 = ~n8353;
assign n12712 = n996 & n11791;
assign n10033 = n1727 & n12514;
assign n796 = n5341 & n11947;
assign n3550 = n1153 | n55;
assign n869 = ~(n3440 | n5755);
assign n2998 = ~(n436 | n3299);
assign n6342 = ~(n6293 ^ n9157);
assign n1655 = n12110 & n1133;
assign n2497 = n7864 & n8099;
assign n5487 = ~(n8299 ^ n10860);
assign n5028 = ~(n9719 ^ n11529);
assign n1382 = n12622 | n3919;
assign n11584 = ~(n6813 | n10871);
assign n2309 = n12200 & n6975;
assign n10029 = ~(n12765 ^ n8664);
assign n12674 = ~(n205 ^ n11965);
assign n10869 = n6373 | n28;
assign n8536 = n191 | n8970;
assign n8136 = n8423 & n7315;
assign n5890 = n9222 | n342;
assign n5009 = ~(n9480 ^ n6956);
assign n4650 = n11887 | n3224;
assign n7491 = n12119 | n7136;
assign n12636 = n4266 & n3626;
assign n3462 = n7495 | n1162;
assign n9426 = n1808 & n2210;
assign n7404 = n8348 | n12282;
assign n543 = ~n7530;
assign n3620 = n4059 | n1079;
assign n11869 = n383 | n10621;
assign n3671 = n10339 | n10854;
assign n10915 = n6461 | n3148;
assign n6221 = ~n4868;
assign n5223 = ~n2629;
assign n10058 = ~(n1061 | n12022);
assign n1296 = ~(n4986 ^ n4810);
assign n12138 = ~n6816;
assign n6716 = ~(n6894 ^ n1616);
assign n11859 = ~(n4389 | n6680);
assign n7521 = ~(n5644 | n7220);
assign n1782 = ~n12764;
assign n1405 = n3285 | n2738;
assign n9298 = ~(n3374 ^ n11789);
assign n8247 = n4953 & n8301;
assign n2925 = n11689 | n11058;
assign n12747 = n3743 | n4654;
assign n2475 = n7504 & n224;
assign n5822 = ~(n10402 ^ n3249);
assign n12616 = n11556 & n6173;
assign n963 = ~(n2893 ^ n1014);
assign n8619 = n3804 | n1700;
assign n10886 = n5945 | n3903;
assign n4017 = ~(n10839 ^ n600);
assign n10893 = n6717 | n5867;
assign n8059 = ~n4700;
assign n3188 = ~(n12734 ^ n1283);
assign n8489 = n9570 | n12050;
assign n2148 = ~(n688 | n7853);
assign n11557 = n5355 | n1455;
assign n6198 = ~(n5234 | n9597);
assign n2380 = ~n3083;
assign n6612 = ~(n7312 ^ n8718);
assign n1606 = n636 | n8259;
assign n3728 = n1511 | n7602;
assign n6980 = ~(n3005 ^ n9251);
assign n2114 = ~(n3201 | n10782);
assign n8246 = ~n9454;
assign n12433 = n12503 | n12771;
assign n4570 = ~(n10481 ^ n6480);
assign n11006 = ~(n5064 ^ n8974);
assign n3482 = ~n2871;
assign n3076 = n12361 | n7876;
assign n4757 = ~(n8573 ^ n9691);
assign n10076 = ~(n5364 | n9781);
assign n12586 = n2597 & n934;
assign n11270 = ~(n6242 ^ n2469);
assign n149 = ~n2913;
assign n160 = n5710 & n12926;
assign n576 = ~n7726;
assign n9706 = ~(n4427 ^ n1110);
assign n7932 = n8545 | n12783;
assign n9585 = n7662 & n1800;
assign n330 = n7919 & n5872;
assign n9976 = n12237 | n6513;
assign n2714 = n6977 | n11896;
assign n4618 = n8348 & n12282;
assign n11782 = n7449 | n5258;
assign n4518 = ~n11623;
assign n7754 = n3746 | n6114;
assign n12410 = ~(n10401 | n8771);
assign n90 = ~(n5995 | n769);
assign n4872 = n2089 | n7962;
assign n3264 = n12025 & n9956;
assign n4345 = ~(n5503 ^ n12844);
assign n5596 = n4958 & n5514;
assign n7112 = n4498 | n3911;
assign n1803 = n10142 | n11430;
assign n2250 = ~(n6702 ^ n9901);
assign n3203 = ~(n6582 ^ n10121);
assign n9288 = n11294 & n7507;
assign n8125 = n5377 & n6701;
assign n1431 = ~(n6994 ^ n1538);
assign n7742 = ~n2094;
assign n11261 = ~(n9165 | n2729);
assign n11581 = n11433 | n3903;
assign n11738 = ~(n9699 ^ n2084);
assign n9679 = ~(n6137 ^ n3901);
assign n11000 = ~(n1177 | n5354);
assign n2752 = ~(n10480 ^ n1173);
assign n12198 = n7685 & n3179;
assign n7007 = ~n4241;
assign n3221 = n5355 | n8859;
assign n3234 = n348 & n5667;
assign n4925 = ~n9390;
assign n3330 = n9070 & n9786;
assign n4488 = n8291 & n3104;
assign n453 = n8674 | n5642;
assign n769 = n6718 | n1476;
assign n8876 = ~(n10443 ^ n5544);
assign n4905 = ~(n10568 ^ n133);
assign n10736 = ~n3294;
assign n6135 = ~(n12428 ^ n7210);
assign n11558 = ~(n3684 ^ n12333);
assign n8109 = ~n7159;
assign n6179 = ~(n4468 ^ n3034);
assign n6378 = ~n4953;
assign n6256 = n4628 | n1163;
assign n6773 = ~(n6688 ^ n6255);
assign n3693 = n8692 & n2421;
assign n2210 = n2786 & n9009;
assign n9140 = n2584 & n9258;
assign n6262 = ~(n5018 ^ n12593);
assign n11649 = n9825 & n8469;
assign n10766 = n5209 ^ n7241;
assign n1167 = ~(n11864 ^ n11458);
assign n9615 = n857 & n6691;
assign n11176 = n4059 | n7246;
assign n2469 = n1397 & n8359;
assign n11483 = ~n9351;
assign n6801 = n11958 | n9971;
assign n5086 = ~n12511;
assign n9292 = n3567 | n11440;
assign n4954 = ~(n7906 ^ n4338);
assign n4183 = n3746 | n5540;
assign n5466 = n2099 | n4818;
assign n7573 = ~n9838;
assign n9361 = ~(n24 ^ n7334);
assign n2864 = n5743 | n7840;
assign n6837 = n7709 | n28;
assign n2683 = ~n544;
assign n3826 = n2137 & n4335;
assign n3475 = ~(n0 ^ n2127);
assign n12050 = n1212 & n3039;
assign n10782 = n5899 & n2928;
assign n10116 = ~(n6935 ^ n12438);
assign n5062 = ~(n11642 ^ n8562);
assign n289 = ~(n2714 ^ n7125);
assign n8818 = n7084 | n9091;
assign n2673 = ~(n6301 ^ n2823);
assign n539 = n4769 & n8956;
assign n2058 = n3014 & n9939;
assign n5975 = n9036 & n8225;
assign n5728 = ~(n496 ^ n2939);
assign n56 = ~(n8342 ^ n5900);
assign n11183 = n1054 | n12657;
assign n324 = n5378 & n8697;
assign n10323 = n8959 | n1413;
assign n2912 = ~(n12478 ^ n7759);
assign n5250 = n8847 | n9356;
assign n5931 = n5291 & n11040;
assign n12306 = n1051 | n5540;
assign n9761 = ~n2742;
assign n6666 = n5456 | n87;
assign n12597 = n12361 | n8768;
assign n8574 = n969 | n5046;
assign n251 = ~(n11285 ^ n33);
assign n1620 = n686 | n9741;
assign n11691 = n9082 | n10865;
assign n6496 = ~(n12318 | n6900);
assign n11088 = ~n4145;
assign n1251 = n10392 & n10911;
assign n9870 = n1642 & n12325;
assign n5828 = n5355 | n1915;
assign n12824 = ~(n1418 ^ n8941);
assign n7883 = n9370 | n4400;
assign n11635 = ~(n12479 | n8174);
assign n994 = ~n1333;
assign n11092 = ~(n5368 | n2221);
assign n8943 = n5394 & n5152;
assign n5904 = ~(n6149 | n3454);
assign n6419 = ~(n3930 ^ n4483);
assign n4116 = n6977 | n3903;
assign n10352 = n8738 | n1509;
assign n3461 = n4628 | n10854;
assign n9628 = ~(n4857 ^ n2310);
assign n6820 = n636 | n12754;
assign n5055 = n8187 | n11746;
assign n11986 = ~(n1657 ^ n9030);
assign n6598 = ~(n2783 | n1531);
assign n7412 = ~(n7221 ^ n10500);
assign n5296 = ~n6188;
assign n11344 = n10953 | n9999;
assign n9275 = n7431 & n1175;
assign n1063 = ~(n9834 ^ n11043);
assign n5188 = n12053 & n4464;
assign n7789 = ~n9311;
assign n3644 = ~n11908;
assign n8030 = ~(n5805 ^ n11447);
assign n1814 = ~(n8084 ^ n11976);
assign n924 = ~(n4272 ^ n11833);
assign n8132 = n2472 | n11952;
assign n3956 = n504 & n3873;
assign n6270 = ~n12537;
assign n10871 = ~n1385;
assign n562 = n5982 | n9166;
assign n6206 = ~n6748;
assign n10680 = ~(n9134 | n10397);
assign n10912 = n2217 | n10916;
assign n4091 = n3552 & n7061;
assign n8474 = n1699 | n8648;
assign n5043 = ~(n8917 ^ n5487);
assign n12082 = ~(n10432 | n154);
assign n10052 = n7050 & n2106;
assign n3677 = ~(n4720 ^ n11918);
assign n7712 = n8308 & n6581;
assign n2944 = ~(n384 | n5972);
assign n9802 = n7493 & n8551;
assign n5768 = ~(n5972 ^ n384);
assign n4753 = ~n4960;
assign n4979 = ~(n6951 | n12081);
assign n7857 = ~(n10104 ^ n4835);
assign n12113 = ~(n12456 ^ n12743);
assign n11039 = ~(n11351 ^ n6023);
assign n1225 = n7551 | n10825;
assign n640 = n12177 & n12386;
assign n9727 = n4628 | n9188;
assign n9122 = n12119 | n8655;
assign n4755 = n5530 | n10311;
assign n5530 = ~n12069;
assign n497 = n7266 | n4385;
assign n12282 = ~(n3967 ^ n5927);
assign n2717 = n3096 | n5012;
assign n7361 = ~(n107 ^ n11005);
assign n7368 = ~(n9274 ^ n12513);
assign n5546 = n3642 | n10963;
assign n12813 = ~n3258;
assign n3629 = n276 | n3507;
assign n6746 = n7191 | n942;
assign n3613 = ~(n3747 ^ n1561);
assign n8190 = ~(n5202 | n9513);
assign n6972 = ~(n6788 | n1214);
assign n1398 = n8738 | n4875;
assign n12487 = n507 & n2797;
assign n3707 = n8390 & n2744;
assign n6547 = ~n10531;
assign n12945 = n10750 | n12124;
assign n7389 = ~n9583;
assign n7140 = n9268 | n11706;
assign n4336 = n686 | n11820;
assign n5627 = n4529 & n8749;
assign n3392 = n9170 | n1546;
assign n11855 = n11390 & n3431;
assign n1999 = ~(n9931 ^ n7926);
assign n1937 = ~n11311;
assign n5678 = ~(n6208 | n5878);
assign n8494 = ~(n2056 ^ n2595);
assign n8235 = ~(n10421 ^ n11367);
assign n5008 = ~n555;
assign n700 = ~(n1202 ^ n10115);
assign n1006 = ~(n6442 | n10619);
assign n2088 = ~(n3810 ^ n3181);
assign n11449 = n4304 | n1117;
assign n5640 = ~(n8296 ^ n1427);
assign n7928 = ~n6016;
assign n8504 = n2530 & n7610;
assign n4309 = ~(n11039 ^ n6641);
assign n8000 = n1699 | n2964;
assign n6977 = ~n6986;
assign n6535 = n393 & n7260;
assign n10388 = ~(n7890 | n9162);
assign n12864 = n5016 & n12202;
assign n8040 = ~n308;
assign n6960 = n5505 & n5009;
assign n10655 = ~n8538;
assign n5681 = n5809 | n8655;
assign n1919 = n6373 | n9078;
assign n2609 = ~(n4415 ^ n8175);
assign n2488 = n7283 | n10419;
assign n2474 = n10827 & n10944;
assign n6550 = n453 & n9013;
assign n5549 = n4911 | n7703;
assign n12049 = ~n12256;
assign n1716 = n6354 & n10952;
assign n12575 = ~(n7850 ^ n3394);
assign n9033 = ~n12001;
assign n7518 = ~(n2003 ^ n12762);
assign n10586 = ~(n10701 | n7148);
assign n10897 = ~n4657;
assign n2658 = ~n5274;
assign n2016 = ~n3064;
assign n10394 = n3992 & n7270;
assign n726 = n8452 | n8978;
assign n2833 = n2050 | n4736;
assign n1734 = n9370 | n6389;
assign n2423 = ~(n10290 | n12640);
assign n4318 = ~(n432 ^ n10882);
assign n4322 = n10142 | n1738;
assign n12133 = n12391 & n4970;
assign n12124 = ~n2347;
assign n4099 = n3912 & n10030;
assign n11142 = n7449 | n4642;
assign n2331 = ~(n10272 ^ n3390);
assign n660 = ~n6624;
assign n6574 = n12596 | n3288;
assign n182 = n5809 | n826;
assign n1979 = n10298 | n9596;
assign n12658 = ~(n6465 ^ n8843);
assign n10534 = ~n6007;
assign n6608 = n12454 | n1029;
assign n9547 = n4498 | n6389;
assign n7502 = n12853 | n9586;
assign n12444 = ~(n6913 ^ n11383);
assign n622 = ~(n5366 ^ n6476);
assign n2161 = n7319 & n2521;
assign n8889 = ~n8373;
assign n529 = n2887 & n6963;
assign n10588 = n7407 & n10662;
assign n5690 = n11923 | n9144;
assign n5602 = n8135 & n2229;
assign n8184 = ~(n7072 ^ n12449);
assign n4656 = ~(n6814 ^ n2929);
assign n2594 = n9082 & n10865;
assign n10180 = n191 | n7881;
assign n1410 = ~(n8804 ^ n8391);
assign n12373 = ~(n12713 | n10027);
assign n2985 = ~(n2550 | n2422);
assign n11223 = ~(n3226 ^ n5066);
assign n2440 = ~(n2569 ^ n9855);
assign n10010 = n12262 & n8253;
assign n9387 = ~(n739 ^ n1318);
assign n6585 = ~(n4075 ^ n3385);
assign n2415 = n2363 & n229;
assign n5007 = n10351 & n3629;
assign n8994 = ~(n8550 | n10934);
assign n6953 = n1466 | n7055;
assign n2403 = n9190 | n8079;
assign n2513 = ~n9124;
assign n6026 = ~(n11037 ^ n1883);
assign n10887 = n5945 | n1413;
assign n5511 = n9297 | n10020;
assign n1718 = n8428 | n3356;
assign n10399 = ~(n2744 ^ n1553);
assign n3339 = ~(n2412 ^ n7991);
assign n6576 = ~(n1544 ^ n9558);
assign n6402 = ~n2585;
assign n4893 = n9389 | n510;
assign n7638 = ~(n7882 | n8454);
assign n8267 = n636 | n7382;
assign n5401 = n9732 & n3404;
assign n12096 = n114 | n1413;
assign n398 = n928 | n6381;
assign n3169 = n11041 | n7423;
assign n3713 = ~n10497;
assign n6191 = n11415 | n12606;
assign n8582 = n11425 & n6025;
assign n8860 = n8582 | n772;
assign n9571 = ~(n767 ^ n9686);
assign n7830 = ~n11055;
assign n4846 = n10835 | n7921;
assign n4588 = ~(n5681 | n10646);
assign n4525 = ~(n546 ^ n7011);
assign n1315 = n5530 | n12686;
assign n3018 = ~(n7740 ^ n12724);
assign n7461 = n3131 | n10813;
assign n3421 = ~n12145;
assign n3748 = n5438 & n11986;
assign n9828 = n5543 & n3485;
assign n6905 = n7690 & n12925;
assign n8563 = ~(n11784 ^ n5536);
assign n12276 = ~(n858 ^ n7757);
assign n9926 = ~(n5982 ^ n3923);
assign n993 = n11887 | n12535;
assign n12477 = n6407 | n2208;
assign n3227 = ~n1091;
assign n5004 = n4647 & n11236;
assign n12027 = n7283 | n11430;
assign n6899 = n5575 | n5540;
assign n10743 = ~(n11620 ^ n3100);
assign n2002 = ~n11541;
assign n6594 = ~(n400 | n4034);
assign n5861 = n4911 | n11827;
assign n8806 = n4617 & n9736;
assign n3838 = ~(n4349 | n3580);
assign n4529 = n8247 & n3868;
assign n6879 = n5666 & n8134;
assign n10300 = ~(n1990 ^ n8207);
assign n9526 = n10502 & n6189;
assign n6967 = n2633 | n11339;
assign n6615 = ~n5282;
assign n4579 = n4561 & n10280;
assign n7892 = n11127 | n9555;
assign n810 = ~n8537;
assign n3343 = n5312 | n2886;
assign n3472 = n11478 & n2558;
assign n9125 = ~(n34 ^ n11214);
assign n12346 = n2599 | n10681;
assign n9549 = n11923 | n9521;
assign n8650 = n1990 & n7635;
assign n7896 = n4508 & n6184;
assign n11541 = n7449 | n1476;
assign n9612 = ~n7081;
assign n12529 = ~(n12582 ^ n3893);
assign n7992 = n752 | n7558;
assign n9708 = ~(n9293 ^ n4664);
assign n8139 = n8187 | n10419;
assign n10890 = ~(n6228 ^ n9525);
assign n1680 = ~(n11505 ^ n520);
assign n12464 = ~n6709;
assign n5953 = n11719 | n6389;
assign n552 = n5361 & n6282;
assign n2026 = ~n3834;
assign n10589 = ~(n6997 ^ n5692);
assign n3939 = n2700 | n3268;
assign n4768 = ~(n2504 | n3814);
assign n7272 = ~(n6914 ^ n4447);
assign n1250 = n2147 | n10329;
assign n2150 = n8505 & n11731;
assign n5586 = ~(n11181 ^ n9803);
assign n11110 = n4644 | n11624;
assign n12320 = ~(n11851 ^ n9255);
assign n1989 = ~n9358;
assign n10267 = ~n3953;
assign n11334 = n2197 | n11855;
assign n4907 = n989 | n8859;
assign n9173 = ~(n7812 ^ n559);
assign n7137 = n2456 | n8644;
assign n12249 = ~(n7753 ^ n11771);
assign n4531 = n5441 | n1862;
assign n7762 = n8462 & n736;
assign n7924 = n1811 & n829;
assign n2184 = n9744 & n3963;
assign n7068 = ~(n1310 ^ n7818);
assign n3200 = ~(n3056 ^ n3367);
assign n4392 = n11958 | n2589;
assign n973 = ~n10228;
assign n1590 = ~(n7700 ^ n9132);
assign n10051 = n6687 & n2509;
assign n1271 = n2605 & n11921;
assign n5926 = n807 | n5540;
assign n2391 = ~(n387 | n11859);
assign n2175 = n11317 | n1265;
assign n1546 = ~n3842;
assign n5719 = ~(n10973 ^ n4399);
assign n2399 = ~(n11711 | n4833);
assign n5148 = ~(n1392 | n2337);
assign n656 = n9246 & n3017;
assign n8493 = ~(n7643 ^ n8232);
assign n5875 = ~(n12551 | n8647);
assign n252 = n8187 | n1162;
assign n11149 = ~(n5075 ^ n9434);
assign n8062 = ~n10640;
assign n9332 = n2494 | n10775;
assign n3594 = n11782 | n5114;
assign n5382 = ~(n12375 | n7444);
assign n6650 = n7116 | n5540;
assign n7563 = ~(n3027 ^ n8459);
assign n12917 = ~(n10502 ^ n6189);
assign n10809 = ~(n10260 ^ n9975);
assign n2872 = ~n10174;
assign n8638 = ~(n11744 ^ n499);
assign n10784 = ~(n3126 ^ n188);
assign n12553 = ~(n3679 ^ n4494);
assign n10274 = n1259 | n3778;
assign n7832 = n41 | n1255;
assign n5288 = n12617 & n1648;
assign n895 = ~n4422;
assign n11104 = n688 & n7853;
assign n2340 = n5530 | n8957;
assign n12889 = n2919 | n6319;
assign n1808 = n10750 | n4818;
assign n11719 = ~n11257;
assign n4601 = ~(n8352 ^ n9879);
assign n9565 = ~(n3585 ^ n3554);
assign n1062 = ~(n11295 ^ n6155);
assign n3917 = ~n6621;
assign n4200 = n164 & n10881;
assign n9304 = n8552 | n6513;
assign n9056 = ~n12031;
assign n9981 = ~(n2828 ^ n12623);
assign n11507 = n10750 | n8644;
assign n1895 = n1827 & n11479;
assign n9152 = ~(n1892 ^ n481);
assign n4302 = n1384 | n9194;
assign n12136 = ~(n6322 | n8035);
assign n12915 = n10928 & n6703;
assign n5584 = ~(n4767 | n4987);
assign n11661 = ~(n8329 | n11063);
assign n10768 = n994 | n7389;
assign n3806 = ~(n9163 ^ n402);
assign n7208 = n3561 | n8312;
assign n9439 = ~(n12084 ^ n6502);
assign n5925 = n12330 & n3980;
assign n3916 = n4796 | n9493;
assign n565 = ~(n10842 ^ n2123);
assign n5036 = n12033 & n6781;
assign n1092 = ~n3988;
assign n11535 = n1271 | n12528;
assign n6209 = n4173 & n7858;
assign n7664 = n12512 & n7414;
assign n8792 = n6252 & n7089;
assign n4582 = n8313 | n879;
assign n11277 = ~n5526;
assign n7056 = ~(n10776 | n5683);
assign n9754 = n4121 & n11975;
assign n11007 = n5783 & n12915;
assign n3398 = ~(n11332 ^ n2772);
assign n742 = ~(n8927 ^ n9071);
assign n12454 = n4777 & n7475;
assign n1616 = n12503 | n1509;
assign n3964 = n5355 | n7389;
assign n10292 = n12503 | n9144;
assign n6279 = ~(n4207 | n3371);
assign n6950 = ~(n10379 ^ n964);
assign n1339 = ~(n6807 ^ n10465);
assign n6968 = ~n6430;
assign n1683 = n5739 & n10241;
assign n4831 = n4510 | n6410;
assign n12036 = ~(n7766 | n12898);
assign n1809 = n12237 | n8655;
assign n1702 = n10750 | n6513;
assign n8502 = n7718 | n5884;
assign n8422 = n332 | n3703;
assign n822 = n5362 & n7725;
assign n9091 = n11602 & n7707;
assign n3191 = ~(n1755 | n6913);
assign n4720 = ~n9332;
assign n5101 = n10797 & n7954;
assign n8516 = n1141 | n1192;
assign n9495 = ~(n7317 | n11492);
assign n2303 = ~(n11885 ^ n9804);
assign n8389 = n11150 & n6726;
assign n2356 = ~n6786;
assign n5392 = n8882 | n12435;
assign n280 = ~(n1335 ^ n10027);
assign n2392 = n149 & n368;
assign n6309 = ~n7458;
assign n3817 = ~(n3247 ^ n5028);
assign n2091 = ~(n5904 ^ n1379);
assign n2964 = ~n5798;
assign n12714 = ~(n2312 ^ n3899);
assign n10672 = n3638 | n7528;
assign n2534 = ~(n11468 ^ n7789);
assign n4364 = ~n8544;
assign n8147 = ~(n12277 ^ n1769);
assign n5610 = ~(n7405 ^ n11066);
assign n6249 = n6881 & n6489;
assign n9051 = n12561 & n1586;
assign n9728 = n1471 & n9763;
assign n4522 = n3734 | n12508;
assign n12890 = ~(n4292 | n3690);
assign n763 = ~n5128;
assign n194 = ~(n5281 ^ n8777);
assign n4780 = n1937 | n2232;
assign n6637 = ~(n8719 | n2637);
assign n3352 = ~n9341;
assign n9252 = n708 & n2032;
assign n4241 = ~(n11561 ^ n4067);
assign n595 = n9248 & n6592;
assign n10018 = n2456 | n12686;
assign n7317 = n8026 | n7395;
assign n10951 = n5554 & n11625;
assign n3259 = ~(n5828 ^ n5186);
assign n11502 = n9943 & n9035;
assign n6282 = ~(n10604 ^ n7356);
assign n3831 = n8276 & n11728;
assign n9930 = ~(n1392 ^ n1992);
assign n2193 = ~(n5345 ^ n2614);
assign n6264 = ~(n5922 ^ n9614);
assign n7343 = ~n11155;
assign n2335 = n9370 | n4775;
assign n8458 = n9370 | n7341;
assign n6825 = ~(n9861 | n6047);
assign n2968 = n1963 & n11769;
assign n8041 = n1003 & n6517;
assign n5529 = n4302 & n4927;
assign n1133 = ~n9197;
assign n5396 = ~n3208;
assign n2001 = n1170 | n6748;
assign n1870 = ~n6745;
assign n8745 = ~n10022;
assign n741 = ~(n9190 ^ n7901);
assign n4752 = ~(n7350 ^ n454);
assign n4328 = n8405 | n12535;
assign n8263 = ~(n9676 | n1451);
assign n4685 = n7641 & n9910;
assign n10865 = ~(n9651 ^ n12543);
assign n8508 = n5486 | n3557;
assign n6328 = n962 | n2020;
assign n8461 = n12284 & n663;
assign n6020 = n3211 | n8653;
assign n4290 = n1051 | n6455;
assign n12847 = n4363 | n6321;
assign n10080 = n6977 | n7558;
assign n10250 = n1123 & n396;
assign n7085 = ~(n11905 ^ n6715);
assign n7759 = ~n9102;
assign n3922 = ~n4462;
assign n9718 = ~(n11306 ^ n5381);
assign n6467 = ~(n8350 ^ n4455);
assign n8032 = ~(n6754 ^ n6573);
assign n10281 = n10912 | n6143;
assign n11914 = ~n11679;
assign n226 = ~(n5350 ^ n5175);
assign n5119 = n4256 | n4467;
assign n2563 = n2108 & n5590;
assign n6651 = n2285 & n2525;
assign n12670 = n1445 & n5727;
assign n6363 = n4356 & n6210;
assign n9064 = n2413 & n10802;
assign n10311 = ~n4436;
assign n747 = ~(n7772 ^ n5421);
assign n10133 = n11266 & n8286;
assign n9945 = ~(n12951 ^ n12840);
assign n9035 = ~(n10413 ^ n12254);
assign n11459 = n7690 & n1564;
assign n1282 = n6696 | n1938;
assign n9042 = ~(n9328 ^ n11826);
assign n11057 = n1903 | n3332;
assign n12839 = n2893 | n1014;
assign n4677 = ~n1500;
assign n6788 = n6373 | n7506;
assign n1330 = n10349 | n7328;
assign n721 = ~(n11099 ^ n3288);
assign n11622 = ~(n12088 | n3490);
assign n6946 = n2456 | n530;
assign n2151 = ~(n4365 | n4323);
assign n9606 = ~(n6816 ^ n7132);
assign n4355 = n5445 | n9215;
assign n7597 = ~(n9250 ^ n12117);
assign n201 = ~n6239;
assign n444 = n9122 | n4460;
assign n8654 = ~(n7306 ^ n10584);
assign n10791 = n8810 | n318;
assign n8688 = n5101 & n9206;
assign n1978 = n7686 | n6074;
assign n10825 = n7100 & n9714;
assign n2606 = n7083 | n672;
assign n1375 = n2285 | n2525;
assign n3236 = n752 | n3903;
assign n10609 = n724 | n8022;
assign n8788 = ~(n983 ^ n4109);
assign n12365 = n3746 | n3903;
assign n8907 = n2613 & n3826;
assign n2123 = n8870 | n8740;
assign n6693 = n9364 & n1458;
assign n1473 = n9170 | n4242;
assign n3604 = n7862 & n3932;
assign n10007 = ~n7616;
assign n2504 = ~n11754;
assign n5666 = ~n11184;
assign n1354 = n5765 | n9078;
assign n6367 = ~(n7019 ^ n9666);
assign n791 = n3618 ^ n11585;
assign n988 = n11531 | n10295;
assign n10905 = n9021 | n4170;
assign n7587 = n7283 | n1915;
assign n4391 = ~n6905;
assign n1733 = n4426 & n1225;
assign n12515 = ~(n9179 ^ n4217);
assign n6339 = n4059 | n10066;
assign n8607 = ~n8634;
assign n12243 = n10169 | n1411;
assign n2018 = n7306 | n10584;
assign n2248 = ~(n161 | n550);
assign n12892 = n1814 | n739;
assign n7547 = ~(n6551 ^ n8243);
assign n5553 = ~(n7569 ^ n12207);
assign n2554 = ~(n8262 ^ n11093);
assign n704 = ~(n9201 ^ n5911);
assign n1345 = ~n3166;
assign n4592 = n1539 | n4400;
assign n1522 = ~(n10417 ^ n3660);
assign n6936 = ~(n5181 ^ n3410);
assign n3097 = ~(n8983 | n4172);
assign n1584 = n2650 & n9728;
assign n10427 = ~(n4384 ^ n6587);
assign n974 = n7221 & n6453;
assign n3913 = n1183 | n5468;
assign n2934 = n1936 & n6723;
assign n5858 = ~n10547;
assign n12360 = ~(n3460 ^ n12229);
assign n3380 = ~(n5533 | n7726);
assign n799 = ~n10964;
assign n7651 = n7391 | n12328;
assign n1172 = n7992 | n8569;
assign n6151 = n5994 & n8722;
assign n8322 = n10309 | n11180;
assign n11015 = n11674 | n2726;
assign n1529 = n4071 | n5612;
assign n537 = n1937 | n11122;
assign n9631 = n7564 & n1363;
assign n7006 = n5596 | n6829;
assign n10829 = n9791 | n10393;
assign n5380 = n8026 | n6169;
assign n5692 = ~(n4806 ^ n6236);
assign n8800 = n8020 & n1644;
assign n12200 = n5507 & n5045;
assign n10099 = ~(n12423 ^ n7303);
assign n8960 = ~(n12597 ^ n5313);
assign n8869 = n1941 | n6169;
assign n629 = ~n11913;
assign n10884 = ~(n6830 ^ n9316);
assign n3222 = ~(n12353 ^ n2350);
assign n11177 = n6718 | n2020;
assign n10362 = ~(n6989 ^ n4836);
assign n8515 = n7678 & n1526;
assign n12415 = ~(n12466 ^ n8960);
assign n1832 = n5120 | n174;
assign n12328 = ~n9195;
assign n5637 = n3453 | n2809;
assign n3995 = n998 & n4129;
assign n11330 = n5031 | n6798;
assign n11682 = ~(n3058 | n5901);
assign n11615 = ~(n4061 | n10437);
assign n8816 = n1937 | n11896;
assign n3699 = n4131 | n10190;
assign n6452 = ~(n605 | n9288);
assign n9490 = ~n9544;
assign n2051 = ~(n8839 ^ n5774);
assign n3318 = n855 | n10699;
assign n12503 = ~n5319;
assign n5444 = ~(n8315 ^ n2789);
assign n7118 = ~(n6244 | n8180);
assign n1777 = n5013 & n3588;
assign n8787 = ~n10116;
assign n9618 = ~n3762;
assign n729 = ~(n11409 ^ n9032);
assign n1681 = ~(n7458 ^ n11748);
assign n7181 = n1249 | n7963;
assign n547 = ~(n2684 ^ n5103);
assign n3695 = n4798 | n4368;
assign n2572 = n4286 & n8472;
assign n7379 = ~n8225;
assign n7576 = ~(n8184 ^ n10655);
assign n9296 = ~(n5338 | n8933);
assign n10119 = n4911 | n2358;
assign n12899 = ~n10391;
assign n1294 = ~(n6392 ^ n4090);
assign n10601 = ~(n6946 ^ n9104);
assign n2550 = n12819 & n3379;
assign n7098 = ~(n5097 | n9773);
assign n7291 = ~(n2148 | n5275);
assign n9501 = ~(n9365 ^ n3307);
assign n2900 = n7802 & n7141;
assign n3756 = n10502 | n6189;
assign n11938 = ~(n11545 ^ n5067);
assign n4067 = ~(n8072 ^ n11527);
assign n8400 = ~(n7271 ^ n11263);
assign n1020 = n2177 ^ n1150;
assign n9226 = n7116 | n2232;
assign n2222 = ~(n7286 ^ n7443);
assign n8718 = ~n2408;
assign n448 = n11543 & n3378;
assign n2052 = ~n1105;
assign n11322 = n8118 & n9965;
assign n8351 = ~(n7071 ^ n8338);
assign n162 = ~(n8835 ^ n8793);
assign n4590 = ~(n2448 ^ n12070);
assign n3077 = ~(n11828 ^ n5133);
assign n9161 = ~n9416;
assign n7575 = n7133 & n2395;
assign n5991 = ~n7826;
assign n11756 = n6352 & n1533;
assign n7177 = n5767 & n5760;
assign n10285 = ~(n8714 ^ n10468);
assign n12453 = ~n458;
assign n9185 = ~n10604;
assign n8723 = ~(n6933 ^ n3994);
assign n12772 = ~n8323;
assign n6112 = ~(n2180 ^ n927);
assign n6971 = ~(n6121 | n5946);
assign n3862 = ~n9099;
assign n2094 = ~(n10922 ^ n11650);
assign n3376 = n580 & n2469;
assign n8116 = n8583 | n1476;
assign n6393 = ~(n4892 | n583);
assign n6433 = ~n535;
assign n7819 = ~(n11875 | n1408);
assign n6561 = n8870 | n9188;
assign n4246 = n4628 | n12883;
assign n11528 = n4561 | n10280;
assign n2960 = ~(n2909 ^ n6280);
assign n6948 = n2630 | n5324;
assign n9337 = ~(n2405 ^ n10090);
assign n719 = n7862 & n4921;
assign n11062 = ~(n5166 ^ n4285);
assign n9489 = n2653 & n12359;
assign n872 = n5915 | n8648;
assign n10689 = n2293 & n10956;
assign n706 = n12594 | n5469;
assign n2142 = ~(n8473 | n2442);
assign n8823 = n7578 & n3644;
assign n9344 = ~n2047;
assign n456 = ~(n3262 ^ n4072);
assign n5307 = ~n9443;
assign n528 = ~(n4379 ^ n11693);
assign n4426 = n7100 | n9714;
assign n3480 = n2830 | n4405;
assign n6709 = n9920 & n5212;
assign n4415 = n11026 | n9160;
assign n7192 = ~(n5695 | n6745);
assign n11059 = ~(n10996 | n8292);
assign n3910 = ~(n12630 ^ n5074);
assign n6670 = n4393 & n4829;
assign n3825 = n1581 & n437;
assign n349 = n1699 | n12080;
assign n3943 = ~n7831;
assign n7362 = ~(n4019 ^ n2027);
assign n12949 = ~(n10034 ^ n5413);
assign n430 = n2456 | n10854;
assign n1424 = n1714 & n2592;
assign n7099 = n3746 | n3356;
assign n8271 = ~(n8166 ^ n3253);
assign n5980 = ~(n2416 ^ n9088);
assign n7078 = n6577 | n7876;
assign n6044 = n7487 | n7752;
assign n7043 = n5860 & n9111;
assign n2624 = ~(n651 ^ n10687);
assign n4280 = ~n10178;
assign n11532 = n1941 | n12816;
assign n3596 = ~(n10228 | n11971);
assign n6677 = n10057 | n5822;
assign n2963 = n5765 | n12771;
assign n8773 = n12243 & n11331;
assign n11523 = ~(n3000 ^ n6639);
assign n5876 = ~n7377;
assign n1781 = ~n4522;
assign n94 = ~(n10686 ^ n8935);
assign n369 = ~(n6066 ^ n8814);
assign n7585 = ~(n4107 ^ n11695);
assign n10305 = n2670 | n10220;
assign n7985 = ~(n2216 ^ n2810);
assign n10073 = n3433 & n1722;
assign n508 = n7862 & n11407;
assign n7359 = ~(n10210 ^ n8366);
assign n4047 = n10926 | n11396;
assign n12123 = ~(n12379 ^ n1429);
assign n9676 = ~(n494 ^ n2070);
assign n12775 = n4059 | n7424;
assign n475 = ~(n9413 ^ n9022);
assign n9546 = ~(n11788 ^ n3641);
assign n8004 = n744 | n11432;
assign n2890 = n12503 | n9521;
assign n7658 = n648 & n6769;
assign n5102 = n10530 | n1038;
assign n2104 = ~(n10461 ^ n12523);
assign n7554 = n2575 & n175;
assign n423 = ~n7023;
assign n9781 = n3954 & n8955;
assign n4930 = ~(n4893 ^ n5085);
assign n6787 = n3961 & n9219;
assign n2995 = n8129 | n12603;
assign n8202 = ~(n3296 ^ n5557);
assign n2794 = ~(n3297 | n12424);
assign n6288 = ~n1190;
assign n12556 = ~(n2702 | n449);
assign n8362 = ~(n3128 ^ n12381);
assign n1637 = ~(n10023 ^ n11085);
assign n3545 = ~(n8142 | n6308);
assign n2578 = ~n9216;
assign n11983 = ~(n3991 ^ n12154);
assign n7036 = ~(n4904 ^ n5493);
assign n1591 = n10262 | n5630;
assign n12287 = ~(n6544 ^ n6435);
assign n1370 = n7839 | n1413;
assign n3559 = ~(n4114 ^ n7336);
assign n10348 = n905 & n11505;
assign n1316 = n2619 & n4978;
assign n1073 = n8789 | n1733;
assign n2977 = ~n9683;
assign n2582 = ~n8763;
assign n10370 = n2911 | n4530;
assign n4809 = ~(n11534 ^ n9184);
assign n10385 = n8814 | n6278;
assign n3847 = ~(n7157 | n6746);
assign n5112 = ~(n5578 ^ n780);
assign n8284 = n6386 & n3841;
assign n1015 = ~(n4566 ^ n10370);
assign n5175 = ~(n382 ^ n1060);
assign n8163 = ~(n8239 ^ n11857);
assign n12572 = ~(n6650 ^ n305);
assign n2583 = ~(n10269 ^ n5295);
assign n7441 = n1051 | n7952;
assign n3994 = ~(n10092 | n1666);
assign n3796 = n12552 | n6989;
assign n6635 = n8187 | n7341;
assign n1299 = ~(n3244 | n6024);
assign n3409 = n5450 | n6694;
assign n3720 = ~(n10761 ^ n3234);
assign n12505 = ~(n9572 ^ n6711);
assign n7824 = ~(n4259 ^ n10003);
assign n5434 = ~n8347;
assign n10459 = ~(n6570 ^ n8478);
assign n3554 = ~(n7441 ^ n3009);
assign n1350 = n9677 & n12869;
assign n9238 = ~(n4788 ^ n2787);
assign n10529 = n4059 | n6402;
assign n4684 = n9299 & n11158;
assign n7850 = n6002 & n9590;
assign n1948 = ~(n816 ^ n7530);
assign n579 = ~(n2856 ^ n3165);
assign n6894 = n11552 | n1047;
assign n9967 = ~(n3895 ^ n1729);
assign n6641 = ~(n6488 ^ n5731);
assign n5469 = n2249 & n1676;
assign n8897 = ~(n12399 | n4889);
assign n8312 = n12098 & n5499;
assign n11497 = ~n4089;
assign n34 = ~(n64 | n5143);
assign n11185 = ~(n10575 ^ n3187);
assign n8613 = n11616 & n3023;
assign n2400 = n5355 | n12328;
assign n5451 = ~(n4562 ^ n12689);
assign n8468 = ~(n4237 ^ n12852);
assign n7721 = ~(n3858 ^ n9738);
assign n6323 = ~n525;
assign n4265 = n5915 | n8644;
assign n9816 = n8206 | n3195;
assign n5067 = n2816 & n9378;
assign n5321 = n254 | n7775;
assign n5484 = n180 | n285;
assign n655 = ~(n6045 ^ n6432);
assign n4593 = ~n2485;
assign n7736 = n8835 & n9595;
assign n6898 = n2308 & n11133;
assign n176 = ~(n4620 ^ n9912);
assign n9594 = ~(n1712 ^ n11632);
assign n1667 = ~n8319;
assign n12578 = n7111 | n11131;
assign n8836 = ~(n11395 ^ n4735);
assign n11690 = n1051 | n7558;
assign n9407 = ~(n8692 ^ n2421);
assign n1255 = ~(n5808 ^ n7573);
assign n11342 = ~(n6018 ^ n5892);
assign n9900 = ~(n2492 ^ n12099);
assign n2844 = ~n10013;
assign n7403 = ~(n2332 ^ n6034);
assign n7050 = ~n2602;
assign n8539 = ~n1420;
assign n7703 = ~n2508;
assign n4245 = ~(n10838 ^ n3060);
assign n5670 = ~(n5649 ^ n3004);
assign n6819 = ~(n2073 | n12028);
assign n4881 = n8705 | n12336;
assign n1300 = n398 & n2322;
assign n10344 = n1442 & n3668;
assign n12514 = n12840 | n12951;
assign n1764 = ~(n6612 | n4896);
assign n4477 = ~(n2943 ^ n11097);
assign n1014 = n7283 | n12843;
assign n2591 = n5786 | n9464;
assign n6337 = ~(n4438 ^ n12498);
assign n3837 = ~(n7507 ^ n7658);
assign n7938 = ~n11526;
assign n5186 = n10739 & n3938;
assign n3551 = ~(n10249 ^ n12082);
assign n1419 = ~(n3565 ^ n1894);
assign n12379 = n9696 | n6394;
assign n1516 = n9953 & n6396;
assign n3060 = n7964 & n9329;
assign n2573 = n6251 | n3403;
assign n11766 = ~(n2531 ^ n9945);
assign n1314 = n2511 & n926;
assign n9943 = ~(n11541 ^ n4936);
assign n2503 = n12503 | n1047;
assign n7949 = ~n2467;
assign n9460 = ~(n5 ^ n3720);
assign n6768 = n7965 & n11876;
assign n3804 = n2437 & n2085;
assign n11809 = ~(n6424 ^ n1332);
assign n7867 = ~(n11408 ^ n12450);
assign n2605 = ~(n7956 ^ n11251);
assign n4645 = ~n8843;
assign n1638 = n8267 & n11939;
assign n9714 = n8428 | n5540;
assign n9983 = ~(n7659 ^ n117);
assign n1928 = n2267 | n1096;
assign n10381 = n2456 | n2964;
assign n2470 = n5305 & n3932;
assign n570 = ~(n10071 | n1604);
assign n12724 = ~n3728;
assign n3253 = n8026 | n12899;
assign n3054 = ~(n11715 ^ n12575);
assign n10552 = ~(n4739 | n1846);
assign n59 = ~(n5598 ^ n11672);
assign n11034 = n7914 & n4351;
assign n4408 = ~(n12513 | n12690);
assign n10948 = ~(n9250 | n10453);
assign n2831 = ~(n6381 ^ n4404);
assign n4401 = n6660 & n5406;
assign n10347 = n6977 | n11820;
assign n10172 = n8552 | n7928;
assign n646 = n3743 | n6138;
assign n7060 = n12155 & n6473;
assign n11196 = n10500 | n974;
assign n2265 = ~(n1006 | n9217);
assign n3639 = ~(n8029 ^ n9423);
assign n9052 = n3604 & n4421;
assign n3503 = ~(n5936 | n2998);
assign n3311 = n4092 | n5907;
assign n10780 = ~n12623;
assign n3771 = ~(n1776 ^ n9452);
assign n12281 = n2099 | n10311;
assign n5467 = ~(n9860 ^ n9100);
assign n1594 = n2393 & n11791;
assign n11993 = n6303 | n8084;
assign n2638 = n11380 | n11115;
assign n7493 = ~(n4171 ^ n10077);
assign n7720 = n5961 & n2804;
assign n9428 = n191 | n7246;
assign n7929 = ~(n1240 ^ n10183);
assign n11137 = ~n11777;
assign n8417 = ~(n8824 ^ n7272);
assign n3783 = ~(n4718 ^ n11260);
assign n6925 = ~n3633;
assign n3883 = ~(n12291 ^ n923);
assign n8355 = n10222 & n3828;
assign n6003 = n1937 | n3903;
assign n9987 = ~(n2618 | n1654);
assign n2757 = ~(n10057 ^ n5399);
assign n156 = ~n9010;
assign n12250 = ~(n7595 ^ n4709);
assign n2308 = n2548 | n8435;
assign n3003 = n186 & n3435;
assign n12381 = ~(n2852 ^ n1789);
assign n4106 = ~(n11684 ^ n10731);
assign n2581 = ~(n3945 ^ n7259);
assign n4708 = ~(n12841 ^ n6563);
assign n7800 = ~n8779;
assign n10261 = n4185 | n4965;
assign n5237 = n10079 | n10538;
assign n743 = ~(n4211 | n6259);
assign n7732 = ~n7814;
assign n9905 = n10835 | n9568;
assign n9918 = n4628 | n4913;
assign n3001 = ~(n5872 ^ n9018);
assign n10275 = ~n4034;
assign n1337 = n1223 | n2892;
assign n2311 = ~(n4899 ^ n4329);
assign n2499 = ~n613;
assign n3035 = ~(n6771 ^ n9662);
assign n3114 = n10605 | n3388;
assign n8721 = ~(n70 ^ n11210);
assign n10726 = n5809 | n12686;
assign n5813 = n8822 | n4472;
assign n2634 = n12708 & n9745;
assign n12767 = n196 | n11477;
assign n6246 = ~(n12074 ^ n1540);
assign n11087 = ~(n9810 | n11696);
assign n5604 = ~(n11281 ^ n4629);
assign n12066 = ~(n8919 | n1582);
assign n828 = ~(n7400 ^ n10089);
assign n7557 = n114 | n11775;
assign n11946 = ~(n3420 ^ n594);
assign n10187 = n10088 & n3295;
assign n3249 = ~n6884;
assign n7484 = ~(n4630 ^ n7722);
assign n11735 = n2042 & n10305;
assign n96 = n4502 | n9610;
assign n1627 = n2424 | n12846;
assign n11452 = n10355 | n5863;
assign n11130 = ~(n8017 ^ n3364);
assign n2666 = ~(n5756 ^ n11913);
assign n9548 = ~n11934;
assign n10448 = n10879 | n3911;
assign n12797 = ~n7523;
assign n7263 = ~(n6812 ^ n12018);
assign n3624 = ~n933;
assign n11758 = n8961 & n3193;
assign n10499 = n2262 & n2066;
assign n6892 = ~(n11289 ^ n11024);
assign n2042 = n2536 | n12112;
assign n8503 = ~(n7393 | n12362);
assign n9650 = ~n1;
assign n1913 = n5859 & n11824;
assign n8130 = ~(n12409 ^ n11258);
assign n5969 = n9878 | n1932;
assign n733 = ~(n5167 ^ n11781);
assign n768 = ~(n5852 ^ n4095);
assign n9992 = ~(n683 ^ n12953);
assign n3892 = ~(n5594 | n11095);
assign n4501 = n1699 | n10422;
assign n5725 = ~n11141;
assign n8196 = ~(n3115 ^ n4853);
assign n7204 = n114 | n2232;
assign n299 = ~n3874;
assign n11078 = n10194 | n9928;
assign n2576 = ~(n1995 | n464);
assign n4084 = ~n6174;
assign n12548 = ~(n6272 ^ n2126);
assign n12347 = n1122 & n12427;
assign n10304 = ~n2924;
assign n7589 = ~(n2871 ^ n6415);
assign n10002 = n962 | n3606;
assign n11668 = n5394 | n5152;
assign n5225 = ~(n3420 | n7634);
assign n669 = n6462 & n7742;
assign n5871 = ~n3479;
assign n12829 = n430 | n10085;
assign n2671 = n6256 & n7489;
assign n2730 = ~n10061;
assign n311 = ~n399;
assign n6962 = ~(n7594 | n4902);
assign n12801 = ~n3087;
assign n10971 = ~(n4697 ^ n6430);
assign n10296 = n11449 & n1365;
assign n5095 = n1809 & n882;
assign n165 = n10142 | n3911;
assign n11594 = n12662 | n10491;
assign n7212 = ~n5758;
assign n2354 = n9787 | n7619;
assign n2068 = n1561 | n12817;
assign n1671 = ~(n8227 ^ n10209);
assign n38 = ~(n12426 ^ n12085);
assign n8114 = ~n2307;
assign n7094 = n3413 | n4877;
assign n11157 = ~(n10541 ^ n8852);
assign n5961 = ~n12746;
assign n10431 = ~(n9570 ^ n12050);
assign n1418 = n7593 & n3377;
assign n10719 = n9929 & n4842;
assign n3985 = ~(n6727 ^ n9439);
assign n5788 = ~n7667;
assign n853 = ~(n6773 ^ n9419);
assign n9984 = ~(n2947 ^ n6033);
assign n122 = ~(n6825 ^ n6100);
assign n10800 = ~(n4637 ^ n4454);
assign n1404 = n7749 & n8602;
assign n8622 = ~n7820;
assign n5437 = ~(n10433 | n4485);
assign n3178 = n8678 & n10154;
assign n12602 = ~n11942;
assign n12476 = n4698 & n3815;
assign n12784 = n1319 | n3417;
assign n7459 = ~(n6788 ^ n4495);
assign n9477 = ~(n6896 | n9856);
assign n374 = n1111 | n11177;
assign n12723 = n9373 | n10916;
assign n10437 = n3116 & n9931;
assign n6832 = n5816 & n6522;
assign n7722 = ~(n1415 ^ n4431);
assign n9521 = ~n8433;
assign n110 = ~(n7792 ^ n12048);
assign n2152 = ~(n8329 ^ n6434);
assign n5775 = ~(n8896 ^ n4710);
assign n7611 = n4380 & n5245;
assign n4669 = ~(n9898 ^ n1513);
assign n2425 = ~(n85 ^ n2884);
assign n6567 = ~(n3784 | n3317);
assign n7339 = n6909 & n845;
assign n6022 = ~(n11752 | n11781);
assign n3562 = ~(n5396 | n6757);
assign n8968 = ~(n356 ^ n3398);
assign n4389 = n989 | n1738;
assign n7900 = n3820 | n10916;
assign n8268 = n114 | n6455;
assign n8368 = n7112 | n7795;
assign n9350 = ~n6947;
assign n9741 = ~n6429;
assign n9591 = n6317 & n12929;
assign n5306 = n4059 | n12843;
assign n5612 = n11801 & n10413;
assign n6329 = n8598 | n5581;
assign n1226 = n11867 | n6075;
assign n6120 = ~(n2541 ^ n10427);
assign n7864 = n4628 | n5326;
assign n11165 = ~n8973;
assign n10795 = n5250 & n2214;
assign n3854 = ~(n8765 ^ n29);
assign n3958 = ~n5041;
assign n1045 = ~(n2700 ^ n566);
assign n7109 = n11652 | n5939;
assign n8401 = n8687 | n1509;
assign n5787 = ~n528;
assign n1236 = n6294 & n1067;
assign n9832 = ~(n5576 ^ n4353);
assign n510 = ~n11662;
assign n10755 = ~n2233;
assign n11603 = n2123 | n11101;
assign n1742 = ~(n9753 | n12671);
assign n1237 = ~(n12584 ^ n436);
assign n3242 = ~n11936;
assign n6838 = ~(n8475 ^ n12600);
assign n5298 = ~(n9341 ^ n1765);
assign n5544 = ~(n1334 ^ n5566);
assign n9995 = n1183 | n12080;
assign n3800 = n9530 | n7879;
assign n3591 = ~n11875;
assign n2191 = n4984 | n9153;
assign n11770 = ~(n3729 | n10250);
assign n3084 = n1092 | n3175;
assign n7649 = ~n3089;
assign n2155 = n5355 | n7881;
assign n9222 = n10196 | n795;
assign n12156 = n4059 | n11430;
assign n3770 = ~(n5174 ^ n6068);
assign n1381 = ~(n12536 | n883);
assign n3174 = n8262 | n3085;
assign n5432 = n5575 | n6455;
assign n3518 = n4325 | n628;
assign n4314 = n137 & n11922;
assign n12226 = ~(n3863 ^ n3293);
assign n7517 = n5087 & n5357;
assign n6528 = ~(n6662 ^ n8311);
assign n8153 = n10844 | n5699;
assign n10271 = ~(n6834 ^ n2996);
assign n9556 = ~(n10605 ^ n1964);
assign n2476 = n10545 & n2498;
assign n915 = ~(n3221 ^ n7846);
assign n5372 = ~n6361;
assign n7758 = ~(n7909 ^ n4432);
assign n11861 = ~(n10666 ^ n10431);
assign n6640 = n3699 & n2733;
assign n2271 = n9131 & n12463;
assign n2286 = ~(n12235 | n12154);
assign n6873 = ~(n4057 ^ n908);
assign n10059 = n3053 & n7943;
assign n6590 = n994 | n1851;
assign n11436 = ~(n952 | n9828);
assign n9818 = ~n6440;
assign n12471 = ~(n4602 ^ n6980);
assign n11650 = ~(n78 ^ n1934);
assign n5766 = ~n173;
assign n12883 = ~n12044;
assign n7004 = n11417 & n1314;
assign n3341 = ~(n11523 | n7973);
assign n10701 = n8113 & n8626;
assign n9877 = ~n10253;
assign n10870 = n800 & n2468;
assign n7286 = n8738 | n4527;
assign n462 = ~(n9453 ^ n9646);
assign n9267 = ~(n5958 | n4765);
assign n4597 = n5271 | n2006;
assign n1180 = n11552 | n5258;
assign n8712 = ~(n3093 ^ n6690);
assign n7861 = ~n10378;
assign n12074 = ~(n8751 ^ n523);
assign n7973 = ~n572;
assign n9224 = ~(n7084 ^ n9091);
assign n5474 = ~n3931;
assign n12530 = n3743 | n8285;
assign n4638 = n4546 | n7545;
assign n4691 = ~(n3088 ^ n853);
assign n6890 = n9878 | n4818;
assign n12388 = ~n12099;
assign n5839 = n573 & n11044;
assign n2751 = n10744 & n2240;
assign n6415 = ~(n4993 ^ n6099);
assign n6864 = n9432 & n7226;
assign n7105 = n7709 | n795;
assign n12736 = ~(n6145 ^ n12101);
assign n8259 = ~n12826;
assign n4393 = n351 | n10275;
assign n3161 = ~(n7019 | n3782);
assign n3150 = n1051 | n6169;
assign n4514 = n4858 & n2243;
assign n3246 = ~(n7652 ^ n4830);
assign n2457 = ~(n9935 ^ n9488);
assign n9101 = ~(n8911 ^ n2734);
assign n4473 = ~(n9900 ^ n5063);
assign n12135 = n1768 | n206;
assign n5324 = ~(n5572 ^ n12908);
assign n4063 = ~(n6210 ^ n6112);
assign n5074 = ~(n8758 ^ n12027);
assign n1793 = ~(n3236 ^ n1057);
assign n10255 = n6336 | n4077;
assign n8009 = ~(n7078 ^ n838);
assign n3904 = n5314 & n217;
assign n5143 = ~(n6260 | n2770);
assign n6831 = n8981 & n4379;
assign n3768 = ~n5368;
assign n279 = n5026 | n9139;
assign n9693 = ~(n12555 | n9947);
assign n2197 = n6977 | n12816;
assign n7997 = n8855 & n10760;
assign n6101 = ~(n5980 ^ n3532);
assign n4300 = ~(n9734 ^ n2857);
assign n10204 = ~(n8633 | n5713);
assign n219 = ~(n12832 | n4271);
assign n12414 = n274 | n11815;
assign n9464 = n2155 & n11112;
assign n9376 = n8850 | n10805;
assign n7937 = ~(n8492 | n6188);
assign n3972 = ~(n8682 ^ n6736);
assign n807 = ~n7320;
assign n7170 = ~n7526;
assign n607 = n5859 | n11824;
assign n6688 = ~(n354 ^ n12793);
assign n11329 = n5204 & n283;
assign n7825 = n5036 | n2991;
assign n3244 = n12012 & n11889;
assign n2856 = ~(n8101 | n10885);
assign n11416 = ~(n866 ^ n1580);
assign n2502 = n12361 | n7395;
assign n10787 = n1867 & n7371;
assign n9349 = n4465 | n12916;
assign n8868 = n11074 & n3652;
assign n12904 = n3256 & n1081;
assign n1901 = n3210 & n10527;
assign n9473 = ~(n10927 ^ n2051);
assign n5710 = n10117 | n5140;
assign n10748 = n3816 & n5228;
assign n10469 = ~n190;
assign n8217 = ~n2699;
assign n6085 = ~(n1009 ^ n1639);
assign n215 = n8941 & n1418;
assign n12820 = ~(n8308 ^ n5607);
assign n273 = n7480 | n1080;
assign n9977 = ~(n4914 | n4364);
assign n4449 = ~n1229;
assign n11677 = n6185 & n5017;
assign n1537 = ~(n1809 | n882);
assign n5780 = n5355 | n2358;
assign n740 = ~n11802;
assign n5573 = n5247 | n9020;
assign n10922 = n636 | n9188;
assign n9685 = n6579 | n3093;
assign n1446 = n3698 & n2394;
assign n12581 = ~(n11867 ^ n6475);
assign n7847 = n11678 | n5805;
assign n288 = n11923 | n1047;
assign n4751 = ~(n1296 ^ n12948);
assign n6257 = ~n7869;
assign n12380 = n10435 | n4895;
assign n4223 = ~n11955;
assign n12937 = ~(n2880 ^ n792);
assign n3348 = n6666 & n8991;
assign n2039 = n5959 & n8534;
assign n7631 = n11577 & n8053;
assign n4621 = ~(n2275 ^ n4543);
assign n1508 = n6191 & n8895;
assign n6211 = ~(n7396 | n5885);
assign n185 = ~(n6204 ^ n11735);
assign n2126 = ~(n1465 ^ n848);
assign n11077 = ~n150;
assign n1890 = ~(n755 ^ n3080);
assign n8820 = ~(n8087 ^ n10371);
assign n11538 = n752 | n7425;
assign n1961 = ~(n6454 ^ n177);
assign n3383 = ~n7459;
assign n6662 = ~(n3359 | n10047);
assign n12361 = ~n12299;
assign n6676 = ~(n11305 ^ n10501);
assign n9217 = ~(n3462 | n7240);
assign n5299 = n825 | n10284;
assign n5580 = n11221 & n3260;
assign n384 = ~(n10252 ^ n8932);
assign n748 = ~n9265;
assign n12291 = ~(n2204 ^ n751);
assign n9953 = ~n6068;
assign n1763 = ~(n1645 | n11000);
assign n262 = ~(n3723 ^ n712);
assign n6673 = n5915 | n10422;
assign n1965 = ~(n929 | n11453);
assign n5040 = n945 | n4521;
assign n2566 = ~(n804 ^ n1716);
assign n1230 = n835 | n7979;
assign n4957 = n8181 | n8485;
assign n7396 = n1941 | n7952;
assign n33 = ~(n12365 ^ n11406);
assign n6577 = ~n2464;
assign n2975 = ~(n5762 ^ n6217);
assign n5716 = ~(n11138 | n10218);
assign n864 = n3996 | n1046;
assign n708 = n8367 | n388;
assign n12286 = n9843 & n1066;
assign n868 = ~(n9345 ^ n3167);
assign n1217 = n2384 & n3852;
assign n3612 = n3682 & n8958;
assign n5322 = ~(n6010 ^ n2117);
assign n12368 = ~(n9785 | n574);
assign n3109 = ~(n9187 ^ n12113);
assign n8594 = n3743 | n5759;
assign n12071 = n4773 & n403;
assign n3083 = n938 & n3311;
assign n238 = ~(n4799 | n7147);
assign n11154 = n11878 | n10215;
assign n12901 = ~(n5848 | n3913);
assign n12656 = ~(n4119 | n378);
assign n5635 = ~(n3667 ^ n3090);
assign n7826 = n6877 & n7354;
assign n8770 = ~(n12271 | n12707);
assign n5077 = n3791 | n11806;
assign n3386 = n5530 | n12446;
assign n2580 = n10682 | n4011;
assign n6383 = n7441 & n3009;
assign n5745 = n10239 & n9325;
assign n11189 = n6877 & n9640;
assign n10879 = ~n3627;
assign n10268 = ~(n6554 ^ n5201);
assign n6274 = ~n11439;
assign n949 = n638 | n7227;
assign n2724 = n10955 | n6744;
assign n1838 = n4683 & n2732;
assign n11205 = ~(n9123 | n3969);
assign n7628 = ~(n12520 ^ n12664);
assign n10019 = ~(n144 | n7137);
assign n8244 = ~n2398;
assign n12298 = n7116 | n5538;
assign n3235 = n1297 & n1391;
assign n5873 = ~(n5553 ^ n2765);
assign n12679 = n3076 | n10868;
assign n8149 = ~n874;
assign n394 = ~(n8235 ^ n10175);
assign n11958 = ~n8336;
assign n2562 = n3015 | n2294;
assign n3133 = n12093 & n10939;
assign n1969 = ~(n10874 ^ n1300);
assign n12672 = ~(n6270 ^ n11978);
assign n5264 = ~n12133;
assign n11520 = ~n11983;
assign n1272 = n4562 | n12689;
assign n5241 = ~(n353 ^ n10828);
assign n775 = n752 | n12357;
assign n5071 = n3533 | n5660;
assign n8566 = ~(n6399 ^ n1740);
assign n1610 = ~(n12129 ^ n5165);
assign n11049 = n10340 & n1460;
assign n3005 = ~(n11081 ^ n3086);
assign n6077 = n7850 | n3566;
assign n6259 = ~(n4357 | n3103);
assign n8124 = n12940 & n4297;
assign n4506 = n8583 | n2020;
assign n2742 = n5964 & n6038;
assign n7667 = ~(n4501 ^ n6334);
assign n7806 = n10142 | n130;
assign n907 = n4528 | n6187;
assign n3718 = n989 | n11746;
assign n866 = n2456 | n10422;
assign n6163 = n9262 | n9521;
assign n3255 = n2099 | n8109;
assign n4031 = ~(n7316 ^ n9090);
assign n6403 = ~(n10601 ^ n1802);
assign n10833 = n5828 & n5186;
assign n5879 = ~(n1688 ^ n8703);
assign n5852 = ~(n6663 ^ n8456);
assign n2918 = ~(n672 ^ n11454);
assign n4185 = n4582 & n3955;
assign n3633 = ~(n9139 ^ n2200);
assign n10186 = n6293 | n11194;
assign n4922 = n8831 ^ n6406;
assign n6365 = n8959 | n3903;
assign n5015 = ~(n11027 ^ n3611);
assign n12085 = ~(n58 ^ n6146);
assign n8798 = n1375 & n3527;
assign n10892 = n6283 & n3543;
assign n8559 = n6554 | n5201;
assign n9514 = n8951 & n11022;
assign n10732 = ~n8960;
assign n2169 = ~n5635;
assign n6921 = n1583 & n7077;
assign n4351 = n4101 & n9349;
assign n10207 = ~n6326;
assign n12256 = n1078 | n5983;
assign n9852 = n2696 & n10412;
assign n3637 = ~(n1044 ^ n5602);
assign n5022 = ~(n8826 | n631);
assign n9170 = ~n9920;
assign n11241 = n4038 & n8589;
assign n5436 = n9000 | n5391;
assign n9979 = ~(n10218 ^ n11393);
assign n12520 = n1185 & n7755;
assign n9065 = ~(n3452 ^ n1370);
assign n7031 = ~(n4195 ^ n12121);
assign n8309 = ~n12904;
assign n2381 = ~(n6777 ^ n2908);
assign n4504 = n4511 & n8863;
assign n7522 = ~(n3593 | n12291);
assign n8552 = ~n12648;
assign n7340 = ~(n6337 ^ n9447);
assign n6425 = ~n12539;
assign n11940 = n5915 | n8740;
assign n5644 = ~(n1415 | n4630);
assign n8099 = n10725 & n5111;
assign n2066 = ~n10959;
assign n7617 = n11744 | n2222;
assign n3293 = ~(n3625 ^ n9031);
assign n10781 = n7405 | n1148;
assign n12956 = n7427 & n11868;
assign n6884 = n2515 & n12925;
assign n6050 = n10157 | n7506;
assign n12348 = n12119 | n9188;
assign n6523 = ~n5001;
assign n7555 = ~n8083;
assign n9005 = n2213 & n1443;
assign n5284 = ~(n9973 ^ n7180);
assign n5695 = ~n4023;
assign n9894 = ~(n6661 ^ n4493);
assign n7267 = n4770 & n560;
assign n8822 = n2456 | n8109;
assign n253 = n10142 | n1455;
assign n9837 = n8187 | n1455;
assign n7833 = ~(n10975 ^ n2152);
assign n4485 = ~(n3469 | n12326);
assign n2592 = n10283 | n4947;
assign n3875 = n11552 | n2020;
assign n4672 = ~(n12625 | n9963);
assign n2109 = ~(n1218 ^ n4600);
assign n5901 = n8967 & n1673;
assign n2295 = n10216 & n2238;
assign n2797 = n4 | n3283;
assign n1523 = ~(n2262 ^ n3564);
assign n1050 = ~(n1706 ^ n313);
assign n10671 = n2228 | n5286;
assign n12941 = ~n4619;
assign n3401 = n5767 & n10848;
assign n3000 = n11732 & n5506;
assign n7854 = ~n2488;
assign n6822 = ~(n7030 ^ n10271);
assign n5758 = n11958 | n5012;
assign n2081 = n5416 & n7347;
assign n3248 = n11462 & n11148;
assign n9798 = n3820 | n4527;
assign n5222 = ~(n7082 | n10579);
assign n5405 = ~(n9549 ^ n4318);
assign n8671 = n5240 & n3932;
assign n8936 = ~(n2731 ^ n5702);
assign n5157 = n4785 & n6869;
assign n8398 = ~(n7997 ^ n3092);
assign n4758 = ~n564;
assign n12738 = n9388 | n10302;
assign n11229 = n12569 | n9067;
assign n610 = n4983 & n9636;
assign n12953 = n1747 & n8610;
assign n8315 = ~(n6961 ^ n9019);
assign n9202 = ~n9036;
assign n12802 = ~(n9527 | n8050);
assign n8005 = n10587 & n10140;
assign n12865 = ~(n236 ^ n3770);
assign n11003 = n4415 & n325;
assign n9696 = ~(n5474 | n11287);
assign n6727 = ~(n2372 ^ n1032);
assign n12697 = ~(n288 ^ n11386);
assign n3292 = ~n9277;
assign n8150 = ~(n5518 ^ n9327);
assign n7221 = ~(n904 ^ n7464);
assign n7572 = n7449 | n5759;
assign n5818 = n8907 | n10483;
assign n4960 = n6353 & n3601;
assign n9346 = ~n5140;
assign n4307 = n7891 & n521;
assign n7064 = n686 | n7876;
assign n8682 = n2832 | n4400;
assign n4012 = n8870 | n3224;
assign n3305 = n12853 | n8648;
assign n8701 = n5025 & n56;
assign n5869 = ~(n2525 ^ n7174);
assign n9160 = ~n10898;
assign n477 = n12797 | n6455;
assign n3710 = n8738 | n9521;
assign n835 = n5355 | n4242;
assign n8662 = ~(n9564 | n706);
assign n12815 = n925 | n1958;
assign n9017 = n4628 | n8644;
assign n1384 = ~n4349;
assign n10836 = ~(n2048 | n8939);
assign n10408 = n4222 & n11724;
assign n9774 = ~(n2820 ^ n9672);
assign n6411 = n3251 | n1274;
assign n11125 = n12635 | n4988;
assign n111 = n10849 & n6284;
assign n1833 = n5181 & n3410;
assign n5945 = ~n9241;
assign n12455 = n11923 | n5258;
assign n900 = ~(n7796 | n4348);
assign n3047 = ~(n4162 ^ n10406);
assign n11448 = ~(n2201 ^ n12725);
assign n6381 = n636 | n826;
assign n8678 = ~n5955;
assign n6269 = ~(n2055 ^ n9941);
assign n3977 = n2921 | n5604;
assign n8521 = n3797 & n10816;
assign n11664 = ~(n6835 ^ n11469);
assign n5201 = ~(n1671 ^ n5862);
assign n10662 = n4628 | n8109;
assign n2773 = ~(n6211 | n2576);
assign n7407 = n2099 | n7382;
assign n3935 = ~(n9967 ^ n1893);
assign n5524 = n1937 | n2815;
assign n848 = n4046 & n12171;
assign n3820 = ~n5198;
assign n1498 = ~n993;
assign n2192 = ~(n10555 | n7791);
assign n9892 = n11552 | n10916;
assign n7537 = n4015 & n4740;
assign n6407 = n5575 | n3903;
assign n2450 = ~n6772;
assign n6202 = ~(n4892 ^ n4591);
assign n6542 = n5793 | n798;
assign n2756 = ~n2885;
assign n814 = ~(n6496 | n8190);
assign n1888 = ~(n7082 ^ n7845);
assign n8442 = n2300 & n4130;
assign n10048 = ~(n11569 ^ n7880);
assign n4366 = n10750 | n12735;
assign n9675 = ~(n3934 ^ n8888);
assign n3566 = ~n3394;
assign n1896 = n4536 & n4220;
assign n8780 = ~(n4451 ^ n1852);
assign n5805 = ~(n5889 ^ n7103);
assign n6368 = n1699 | n7382;
assign n6840 = ~(n7207 ^ n12674);
assign n12296 = n11026 | n9078;
assign n6231 = n752 | n5538;
assign n1699 = ~n5283;
assign n9529 = n3743 | n8643;
assign n5866 = n1982 | n7621;
assign n202 = n2382 & n948;
assign n3745 = ~(n6705 ^ n5909);
assign n3603 = ~n5544;
assign n11988 = n10879 | n7881;
assign n3331 = ~(n7462 ^ n2105);
assign n2817 = n4498 | n10066;
assign n1089 = n1024 | n7498;
assign n3836 = ~n2565;
assign n4622 = n12361 | n5012;
assign n7429 = ~(n5453 ^ n5550);
assign n9245 = n2872 | n7876;
assign n1193 = ~(n515 ^ n5941);
assign n429 = ~(n6629 ^ n8667);
assign n2030 = n7961 & n10969;
assign n10761 = n10835 | n5502;
assign n11066 = ~(n8937 ^ n534);
assign n9733 = ~(n422 ^ n12482);
assign n11844 = ~(n2760 ^ n1555);
assign n4406 = ~(n12122 ^ n11191);
assign n5933 = ~(n4501 | n8630);
assign n1569 = n10108 | n1455;
assign n12004 = ~(n5633 ^ n9424);
assign n7829 = ~n4409;
assign n9063 = ~(n621 | n6844);
assign n3675 = ~n6251;
assign n1836 = ~n10783;
assign n1356 = ~(n12838 ^ n3450);
assign n10844 = ~(n7309 ^ n9083);
assign n5349 = ~(n90 | n12732);
assign n2232 = ~n11728;
assign n1007 = n989 | n7246;
assign n8573 = n1944 & n782;
assign n1279 = n4849 | n1935;
assign n300 = ~(n12487 | n1857);
assign n8732 = n7449 | n795;
assign n11885 = ~(n8848 ^ n5651);
assign n53 = ~(n7227 ^ n10494);
assign n1023 = ~(n1034 ^ n5722);
assign n4578 = n6241 & n9948;
assign n6461 = n5765 | n8643;
assign n8997 = ~(n5415 | n389);
assign n5039 = n10679 | n6409;
assign n7126 = n5575 | n5311;
assign n1328 = ~(n5822 ^ n2757);
assign n12741 = ~n9246;
assign n11901 = ~n6521;
assign n10663 = ~n6889;
assign n681 = n2215 | n6729;
assign n7034 = ~(n12960 | n10487);
assign n6563 = n127 & n12679;
assign n1570 = ~(n10720 ^ n8088);
assign n10690 = ~(n7032 | n10895);
assign n2956 = n9607 | n4429;
assign n227 = ~(n8205 ^ n6820);
assign n1035 = ~(n5397 ^ n6346);
assign n3479 = n4441 & n4854;
assign n12533 = ~(n12701 ^ n5309);
assign n470 = ~(n6975 ^ n11853);
assign n8088 = ~(n5643 ^ n9173);
assign n1556 = n2367 | n9521;
assign n11616 = n10983 | n2817;
assign n8421 = ~n2831;
assign n474 = n10835 | n3451;
assign n10444 = ~(n41 ^ n383);
assign n2156 = n10518 | n2916;
assign n874 = ~(n2571 ^ n11342);
assign n7765 = ~n10096;
assign n2010 = n9943 | n9035;
assign n9771 = ~(n8612 ^ n2335);
assign n3407 = ~(n4619 | n2719);
assign n3918 = n7937 | n11145;
assign n6804 = ~(n8003 | n11638);
assign n7648 = ~(n3645 ^ n3493);
assign n6926 = ~n508;
assign n6571 = n5915 | n4913;
assign n1352 = n752 | n2754;
assign n10816 = ~n6467;
assign n12193 = ~(n7045 ^ n10937);
assign n8492 = ~n12910;
assign n3952 = n4514 & n9659;
assign n7455 = ~(n1665 ^ n5196);
assign n522 = n8738 | n1047;
assign n7087 = ~(n6801 | n6011);
assign n11079 = n760 ^ n12835;
assign n1155 = n6053 & n5830;
assign n1899 = n9170 | n3911;
assign n7207 = ~(n7288 ^ n4845);
assign n9055 = n7527 & n9772;
assign n10744 = n5575 | n11122;
assign n11866 = ~n11022;
assign n1903 = ~(n5544 | n10443);
assign n4298 = n2832 | n11827;
assign n1982 = n11984 & n6460;
assign n4167 = n3127 | n7881;
assign n1086 = ~(n8776 | n11526);
assign n9447 = ~(n12270 ^ n11676);
assign n12139 = ~(n7549 ^ n8096);
assign n10906 = ~n9414;
assign n3574 = n7629 & n2112;
assign n2832 = ~n4516;
assign n7381 = ~(n9028 | n3945);
assign n9860 = ~(n3276 | n10787);
assign n6025 = n10818 & n9949;
assign n541 = n4131 & n10190;
assign n4878 = n683 & n12834;
assign n2883 = n2834 & n10526;
assign n8855 = ~n11557;
assign n46 = n10776 & n5683;
assign n5837 = ~n6855;
assign n9186 = n12878 & n10906;
assign n1280 = ~n8241;
assign n5114 = n2168 & n2354;
assign n9281 = n379 | n5193;
assign n1132 = ~(n2659 ^ n6419);
assign n6136 = n124 & n11883;
assign n7899 = n7449 | n9144;
assign n10597 = ~(n37 ^ n11920);
assign n7578 = n11055 & n12958;
assign n6874 = ~(n10488 | n6039);
assign n12633 = n7283 | n11746;
assign n2635 = ~(n1866 ^ n10603);
assign n6566 = n12957 & n71;
assign n5107 = n12237 | n3924;
assign n10603 = ~(n9271 ^ n4185);
assign n8154 = ~n1765;
assign n9959 = ~n8455;
assign n2216 = ~(n8288 | n3999);
assign n4410 = ~(n420 ^ n10308);
assign n11970 = ~n8122;
assign n11969 = n9887 | n9226;
assign n1656 = n5902 | n1455;
assign n8345 = ~n1232;
assign n3270 = ~(n5720 ^ n6565);
assign n8359 = n7690 & n12489;
assign n4022 = n5491 | n7743;
assign n5855 = n1072 | n2975;
assign n7608 = n3743 | n1739;
assign n9364 = ~n2345;
assign n1649 = n1231 | n10446;
assign n7316 = n1051 | n3903;
assign n4358 = n191 | n8524;
assign n7427 = n2470 & n1994;
assign n9596 = ~(n2653 | n12359);
assign n12891 = ~(n7894 | n1693);
assign n3586 = ~(n8829 | n8979);
assign n7881 = ~n11877;
assign n4268 = ~(n10929 ^ n6328);
assign n118 = n8481 | n1048;
assign n2598 = ~n12644;
assign n2170 = n10846 | n5525;
assign n7942 = ~(n10405 ^ n11004);
assign n2877 = ~n11523;
assign n8912 = n994 | n11827;
assign n1640 = n3196 & n2274;
assign n10097 = n4929 & n6833;
assign n4056 = n10051 & n1836;
assign n3946 = ~(n11069 | n10056);
assign n8999 = ~(n9604 | n1743);
assign n5874 = ~(n11265 ^ n957);
assign n7716 = n7731 & n3472;
assign n11132 = n4973 & n12687;
assign n3251 = n8870 | n1932;
assign n2876 = n4539 | n893;
assign n10541 = n10157 | n6138;
assign n12057 = ~(n8404 ^ n11739);
assign n6437 = n11341 | n8484;
assign n4294 = ~(n12788 | n11907);
assign n9517 = ~n1820;
assign n2793 = n10926 & n11396;
assign n10159 = n10377 & n6673;
assign n11537 = ~(n9283 ^ n9623);
assign n128 = n12119 | n4818;
assign n12288 = n5915 | n2964;
assign n11235 = ~n2537;
assign n1231 = n3222 & n12228;
assign n4661 = ~n7720;
assign n10702 = n7965 & n10990;
assign n7827 = n9389 | n7703;
assign n498 = ~(n6944 ^ n3897);
assign n5759 = ~n11296;
assign n978 = ~(n8386 ^ n5136);
assign n9656 = n10750 | n12686;
assign n12955 = n12858 | n8742;
assign n5373 = n3324 | n9160;
assign n4967 = n2515 & n5645;
assign n9036 = n6358 & n2749;
assign n9024 = ~(n2979 | n4298);
assign n6292 = n2287 & n12313;
assign n2238 = ~(n6810 ^ n635);
assign n3703 = n6836 & n2004;
assign n3878 = n3072 | n8111;
assign n3744 = ~(n9240 ^ n11671);
assign n9623 = ~(n9884 ^ n3411);
assign n4852 = ~(n370 ^ n2780);
assign n4711 = ~(n7322 ^ n256);
assign n8604 = ~(n11526 ^ n7175);
assign n9339 = n11887 | n3924;
assign n3856 = ~n1994;
assign n9363 = ~(n4563 ^ n8007);
assign n12896 = ~(n2981 | n6444);
assign n71 = ~n1412;
assign n4191 = ~(n7848 ^ n10574);
assign n3460 = ~(n9326 ^ n4920);
assign n4608 = n1896 | n1135;
assign n3219 = n6358 & n7294;
assign n24 = n7283 | n1079;
assign n8815 = n4613 & n4098;
assign n11820 = ~n3022;
assign n970 = n8295 | n5242;
assign n5919 = n10417 & n10146;
assign n11685 = n12468 & n1749;
assign n6440 = n11038 & n12451;
assign n9043 = n636 | n12080;
assign n2272 = n11958 | n11896;
assign n6935 = ~(n7409 ^ n10099);
assign n11432 = ~(n4468 | n7508);
assign n10001 = n1407 | n4886;
assign n3020 = n137 & n521;
assign n7488 = ~(n6937 ^ n12257);
assign n6757 = ~(n12374 ^ n7179);
assign n7444 = ~(n9776 | n11649);
assign n12447 = n1937 | n5540;
assign n9829 = n5631 & n5068;
assign n12262 = n8428 | n10903;
assign n4481 = ~n5732;
assign n961 = n953 & n10528;
assign n1504 = ~n8184;
assign n9359 = ~(n7539 ^ n2078);
assign n11403 = ~n7168;
assign n189 = n1937 | n8768;
assign n7001 = n1470 & n1917;
assign n3296 = n4168 & n4572;
assign n7214 = n6924 & n12527;
assign n11201 = n1097 & n3842;
assign n10919 = ~n12221;
assign n5268 = ~(n12781 ^ n3843);
assign n1460 = ~(n8341 ^ n8747);
assign n7665 = ~(n1462 ^ n10617);
assign n1312 = ~(n11589 ^ n9892);
assign n3635 = ~(n9346 ^ n12926);
assign n3897 = ~n8783;
assign n468 = n10097 | n2415;
assign n7641 = n9982 | n2386;
assign n9398 = ~(n2449 ^ n5721);
assign n12105 = n8164 & n4762;
assign n8394 = n10196 | n10916;
assign n8085 = n114 | n2815;
assign n5838 = n10281 & n9087;
assign n3142 = ~n9089;
assign n1883 = n636 | n1932;
assign n10783 = n989 | n10066;
assign n8115 = n6391 & n5824;
assign n8106 = ~(n12794 ^ n8113);
assign n1310 = ~(n2203 ^ n6915);
assign n9749 = n3127 | n12328;
assign n589 = n10142 | n1546;
assign n9968 = ~(n5043 ^ n2237);
assign n12013 = ~n5742;
assign n8915 = n8026 | n8414;
assign n1188 = ~(n7528 ^ n12216);
assign n5729 = n349 & n3520;
assign n2054 = ~(n6843 ^ n12156);
assign n5789 = n2324 & n3730;
assign n11488 = ~n11577;
assign n9085 = n5172 | n3111;
assign n8369 = n9370 | n3911;
assign n6638 = ~(n12098 ^ n3561);
assign n11590 = ~(n1157 ^ n12418);
assign n8967 = n4213 | n6233;
assign n7093 = ~(n10060 ^ n11229);
assign n366 = ~(n7378 ^ n2914);
assign n9087 = n3607 | n4794;
assign n3725 = n6561 | n8008;
assign n11797 = ~(n9842 ^ n7080);
assign n2167 = n10091 | n100;
assign n11207 = ~n6990;
assign n6286 = ~n12516;
assign n387 = ~(n12223 | n7114);
assign n2108 = n7160 & n7610;
assign n1624 = n5053 & n12655;
assign n3481 = ~(n2710 | n4982);
assign n9734 = n6538 & n10035;
assign n11493 = ~n9342;
assign n11549 = ~(n2036 ^ n2853);
assign n6207 = ~(n6426 ^ n11009);
assign n7297 = ~(n12857 ^ n2212);
assign n2731 = ~(n10544 ^ n3315);
assign n148 = n10569 | n3479;
assign n8304 = n8870 | n12735;
assign n4179 = ~n4799;
assign n2080 = n284 & n10693;
assign n12696 = n7757 | n858;
assign n11123 = n8959 | n11410;
assign n7620 = n4498 | n7881;
assign n12330 = n4206 | n4303;
assign n10932 = ~(n7415 ^ n1499);
assign n2895 = ~(n11373 ^ n9883);
assign n9922 = n191 | n9397;
assign n5582 = n11958 | n11775;
assign n3016 = n10404 & n8624;
assign n9117 = ~(n6930 | n8873);
assign n4224 = n4287 & n12376;
assign n10240 = ~(n1783 ^ n906);
assign n4895 = n3688 & n12045;
assign n4559 = ~(n12309 | n4593);
assign n11204 = n58 | n12426;
assign n11314 = ~(n11861 ^ n4410);
assign n5799 = ~(n10420 ^ n1875);
assign n8387 = n191 | n7341;
assign n7741 = n6996 & n1137;
assign n4969 = ~(n4508 ^ n8495);
assign n8663 = n380 & n12540;
assign n7300 = n8367 & n388;
assign n10203 = ~(n6137 | n9404);
assign n11349 = n11433 | n11820;
assign n3521 = n1824 & n5011;
assign n11305 = n10835 | n7506;
assign n10460 = ~(n8002 ^ n1494);
assign n9891 = ~(n2799 ^ n7711);
assign n8581 = ~(n12296 ^ n12877);
assign n10148 = n3820 | n4875;
assign n119 = ~(n5563 | n5749);
assign n2479 = n1222 & n9417;
assign n3990 = ~(n2235 ^ n5763);
assign n11061 = n5109 & n12295;
assign n6213 = n9504 & n11910;
assign n3657 = ~(n12642 ^ n1589);
assign n3287 = ~(n6443 ^ n8820);
assign n1500 = n3743 | n2020;
assign n9633 = n6827 & n10221;
assign n7592 = ~(n7893 ^ n6344);
assign n7828 = ~(n11068 | n7813);
assign n3204 = ~(n6792 ^ n6315);
assign n10649 = ~n1088;
assign n12871 = ~n223;
assign n5536 = ~(n6165 ^ n3663);
assign n10853 = ~(n10819 ^ n2776);
assign n450 = ~(n1797 | n8525);
assign n10249 = ~(n5139 | n5385);
assign n5239 = ~n7428;
assign n12637 = ~(n7042 ^ n10717);
assign n647 = ~(n12315 ^ n1277);
assign n6617 = ~n10163;
assign n1128 = ~n4199;
assign n11481 = ~n6688;
assign n10867 = n11867 & n6075;
assign n11271 = n8114 | n12902;
assign n12020 = ~(n467 ^ n10549);
assign n5872 = ~(n7308 ^ n12751);
assign n6679 = ~(n3010 | n3702);
assign n1912 = ~(n4980 ^ n6139);
assign n3335 = n6577 | n5538;
assign n4470 = ~(n4880 ^ n7931);
assign n1261 = ~n9592;
assign n8358 = ~(n10740 ^ n4444);
assign n11548 = ~(n10615 | n4699);
assign n1022 = ~n10643;
assign n2083 = n3862 & n57;
assign n10173 = n7078 | n12905;
assign n7804 = n12878 | n10906;
assign n3519 = n5125 & n7598;
assign n2234 = ~(n4278 | n9769);
assign n12119 = ~n4805;
assign n3123 = n10339 | n8109;
assign n9644 = ~n9482;
assign n1070 = ~n2968;
assign n11217 = ~(n4613 ^ n10352);
assign n6088 = n11193 | n5636;
assign n2822 = n6036 | n707;
assign n9664 = n11849 | n7971;
assign n5957 = n784 | n4440;
assign n8385 = ~(n9810 ^ n7183);
assign n5152 = n1699 | n5468;
assign n12372 = n852 ^ n9711;
assign n10 = ~n10987;
assign n2537 = n4828 & n1512;
assign n4343 = ~n4938;
assign n4850 = n12241 & n9235;
assign n8786 = n12119 | n12441;
assign n10071 = ~(n10377 | n6673);
assign n7872 = n6486 | n1464;
assign n2681 = n5010 | n2080;
assign n3370 = ~n12106;
assign n12301 = n529 | n8272;
assign n3698 = n5181 | n3410;
assign n2886 = ~(n2997 | n6848);
assign n4737 = ~(n547 | n2487);
assign n1762 = n889 & n6430;
assign n953 = n2564 & n11662;
assign n8982 = ~n3517;
assign n3506 = n386 | n9354;
assign n7102 = ~(n7769 ^ n1970);
assign n4269 = ~(n10139 ^ n3615);
assign n4838 = n9010 & n10988;
assign n5236 = n6877 & n2024;
assign n1820 = n9372 & n3358;
assign n4814 = n8512 | n3286;
assign n4508 = n18 | n9599;
assign n737 = n10196 | n3606;
assign n3807 = n2217 | n4474;
assign n6133 = n10750 | n7136;
assign n1297 = ~n12280;
assign n927 = ~(n6673 ^ n12863);
assign n12821 = ~n8487;
assign n5458 = n252 | n3957;
assign n2020 = ~n10990;
assign n403 = ~n7748;
assign n3138 = ~(n8548 | n6380);
assign n10996 = ~n9263;
assign n8450 = n890 & n2327;
assign n2160 = ~(n9699 | n4684);
assign n9655 = ~(n5207 ^ n7367);
assign n1834 = ~n5614;
assign n12604 = n3743 | n3599;
assign n11450 = n8870 | n7928;
assign n7737 = ~(n9922 ^ n7669);
assign n4790 = n4778 | n1932;
assign n6652 = n11433 | n11775;
assign n4575 = ~(n12949 | n8289);
assign n12579 = ~n9711;
assign n10955 = n7116 | n6169;
assign n10060 = ~(n12663 | n593);
assign n7469 = n3127 | n2358;
assign n2903 = ~(n8542 ^ n8434);
assign n12562 = ~(n8862 ^ n6630);
assign n12722 = n1177 & n5354;
assign n4325 = ~(n1596 ^ n2450);
assign n10112 = n12303 & n1394;
assign n12517 = ~(n10552 ^ n11925);
assign n7419 = ~(n4511 ^ n2623);
assign n11022 = n684 & n11483;
assign n11181 = n9373 | n3606;
assign n2334 = ~n2851;
assign n3071 = n12746 ^ n742;
assign n944 = ~(n1708 ^ n8882);
assign n10937 = n1323 | n11688;
assign n3651 = n147 & n12571;
assign n3687 = n9917 | n9958;
assign n10931 = n1449 & n1174;
assign n9059 = n6672 & n1529;
assign n12033 = n989 | n4242;
assign n6789 = n8613 | n5943;
assign n6992 = ~(n10697 ^ n3995);
assign n7371 = ~n8734;
assign n11044 = n989 | n12843;
assign n5903 = ~(n8605 | n2161);
assign n11618 = n7485 & n6576;
assign n611 = ~(n11109 | n80);
assign n9919 = ~(n12448 ^ n4930);
assign n9108 = n994 | n1915;
assign n4863 = n3127 | n6402;
assign n9415 = ~(n8361 ^ n9641);
assign n4543 = ~(n8147 ^ n5270);
assign n5677 = n7526 | n790;
assign n6082 = ~(n4738 | n2794);
assign n2106 = n8600 & n2445;
assign n3830 = n4995 & n1652;
assign n7296 = ~(n5967 ^ n7486);
assign n9242 = ~(n301 ^ n10285);
assign n11121 = n10822 | n4711;
assign n8176 = n5434 & n11354;
assign n4382 = n1867 | n7371;
assign n4262 = ~n2387;
assign n2258 = n365 | n5457;
assign n11810 = n6313 & n4816;
assign n11767 = n7299 | n2239;
assign n6984 = ~(n4147 | n9011);
assign n6306 = ~n2116;
assign n10293 = n7978 & n9566;
assign n6771 = ~(n10526 ^ n3458);
assign n5769 = n10835 | n4864;
assign n5025 = ~n6070;
assign n11025 = ~(n7098 ^ n2391);
assign n2813 = ~n7244;
assign n9800 = n12417 | n11590;
assign n1673 = n986 | n11426;
assign n6300 = ~(n6408 ^ n528);
assign n2539 = n2099 | n12754;
assign n6486 = n7449 | n10916;
assign n9172 = ~n11672;
assign n7226 = n11384 & n668;
assign n12271 = n5355 | n2076;
assign n1588 = ~(n7600 ^ n8463);
assign n9467 = ~(n8593 ^ n6511);
assign n5569 = n8870 | n530;
assign n11736 = ~n2402;
assign n693 = n897 | n4850;
assign n9488 = ~(n2563 | n2196);
assign n4054 = n9500 | n9964;
assign n10580 = ~(n10221 ^ n5461);
assign n10398 = n6078 | n2672;
assign n4854 = n4979 | n8884;
assign n2153 = ~(n6731 ^ n2283);
assign n8726 = ~(n12248 ^ n1573);
assign n11426 = n4213 & n6233;
assign n12131 = n95 & n6792;
assign n3363 = ~(n981 | n3296);
assign n9630 = ~(n6560 ^ n3741);
assign n875 = n7874 & n12918;
assign n1463 = n5183 & n6299;
assign n2195 = n9648 | n5802;
assign n485 = ~(n12670 | n8341);
assign n3373 = ~(n7919 | n5872);
assign n10500 = n11580 & n3823;
assign n2329 = n2456 | n12124;
assign n9276 = ~n662;
assign n7686 = n9389 | n7881;
assign n303 = n1404 | n10558;
assign n5698 = n10771 | n11045;
assign n8170 = ~(n2161 ^ n8605);
assign n3416 = ~(n10288 ^ n7900);
assign n8719 = ~(n1152 ^ n10123);
assign n10618 = ~(n12319 ^ n2030);
assign n5808 = n686 | n2815;
assign n3812 = ~(n9026 ^ n4683);
assign n6835 = ~(n9229 ^ n6762);
assign n5408 = n3743 | n9521;
assign n5608 = n2167 & n8413;
assign n4137 = ~(n5254 ^ n8264);
assign n5887 = n8583 | n4527;
assign n11927 = n10915 & n6020;
assign n11194 = n2976 & n11495;
assign n12498 = ~(n11450 ^ n10908);
assign n1105 = n5134 & n5477;
assign n5566 = ~(n3964 ^ n2981);
assign n10819 = ~(n2119 ^ n2264);
assign n795 = ~n8028;
assign n5802 = n8959 | n11775;
assign n2859 = ~(n9204 ^ n8693);
assign n762 = n2456 | n1932;
assign n7188 = n3096 | n6455;
assign n6203 = n4059 | n4242;
assign n8285 = ~n6441;
assign n3727 = ~(n2029 ^ n8500);
assign n1544 = ~(n10128 ^ n2451);
assign n1909 = n9656 | n12411;
assign n12880 = n9812 | n10836;
assign n10740 = n4662 | n8987;
assign n304 = ~n4484;
assign n4317 = n4547 & n7335;
assign n8390 = ~(n7200 ^ n7499);
assign n8526 = n4772 & n9470;
assign n8908 = n12361 | n10919;
assign n6624 = ~(n7365 ^ n1753);
assign n1861 = ~n4439;
assign n10624 = n12344 & n815;
assign n9682 = n2367 | n795;
assign n7688 = n4628 | n12686;
assign n8859 = ~n1835;
assign n10216 = n8159 | n5299;
assign n82 = ~(n12348 ^ n9399);
assign n746 = ~(n3437 ^ n12075);
assign n2775 = ~(n12052 ^ n6440);
assign n7308 = ~(n1631 ^ n7296);
assign n9531 = n10157 | n4654;
assign n4147 = ~(n9369 | n2952);
assign n11588 = ~(n11262 ^ n9056);
assign n7244 = n11552 | n4654;
assign n8120 = n5504 | n9925;
assign n3186 = n3930 & n4483;
assign n12024 = n9827 & n11599;
assign n657 = ~(n7662 ^ n1800);
assign n9856 = ~n1050;
assign n5854 = ~(n6472 | n2174);
assign n2629 = n5945 | n6455;
assign n3384 = ~(n7520 ^ n9133);
assign n8391 = ~(n1151 ^ n6998);
assign n5662 = n9498 | n3880;
assign n2449 = ~(n9155 ^ n3395);
assign n6591 = ~(n7790 ^ n6416);
assign n2251 = n6667 | n604;
assign n3839 = ~(n12443 ^ n1734);
assign n4896 = ~n4850;
assign n4211 = ~(n7916 | n2642);
assign n12199 = ~n1456;
assign n4036 = ~(n4588 | n7660);
assign n9136 = ~(n1228 ^ n7560);
assign n10338 = n2217 | n8643;
assign n3997 = n5809 | n4818;
assign n9722 = ~(n8617 ^ n2375);
assign n2159 = n6924 | n12527;
assign n1052 = n7024 | n4661;
assign n2994 = ~n3734;
assign n1696 = n8583 | n4474;
assign n5509 = ~(n1624 ^ n6194);
assign n1954 = ~(n5825 ^ n12620);
assign n4085 = ~n8760;
assign n9061 = n11714 | n5551;
assign n9772 = ~n5344;
assign n11704 = n191 | n130;
assign n11193 = ~n7416;
assign n5285 = n8416 | n2933;
assign n8790 = n752 | n2232;
assign n1790 = ~n8204;
assign n9072 = ~(n12287 ^ n241);
assign n10779 = ~(n10038 ^ n9451);
assign n6627 = ~n8094;
assign n9150 = n6577 | n12816;
assign n7683 = ~n11243;
assign n8045 = n5575 | n12357;
assign n3761 = n3127 | n12843;
assign n2149 = n4679 & n1668;
assign n4486 = ~(n12611 ^ n10753);
assign n10479 = ~n10402;
assign n11931 = n9171 | n9221;
assign n2365 = ~(n4991 ^ n7427);
assign n9810 = ~(n8275 ^ n9052);
assign n12552 = ~(n5948 ^ n233);
assign n7979 = n11255 & n2591;
assign n5742 = ~(n4465 ^ n475);
assign n8350 = ~(n5486 ^ n3662);
assign n11878 = n10611 | n7249;
assign n4546 = n7116 | n5012;
assign n1301 = ~(n262 ^ n5634);
assign n4057 = n5233 & n11201;
assign n11687 = n989 | n8524;
assign n12041 = n6042 | n576;
assign n635 = n3018 ^ n11831;
assign n7158 = n3976 & n12059;
assign n3195 = ~(n4908 | n6596);
assign n7605 = ~(n6153 ^ n9374);
assign n7273 = ~n3020;
assign n12398 = n7420 | n12475;
assign n1492 = ~(n12324 ^ n2736);
assign n12911 = ~(n4148 ^ n8399);
assign n2871 = n9634 & n1250;
assign n1641 = ~n633;
assign n8332 = n7052 | n1864;
assign n8363 = ~n9757;
assign n7253 = n1951 ^ n3432;
assign n2270 = n6516 | n4321;
assign n360 = ~(n178 ^ n5387);
assign n4624 = ~n1826;
assign n1706 = n2217 | n28;
assign n2384 = ~n6661;
assign n11991 = ~(n4595 | n5624);
assign n6058 = n6977 | n3468;
assign n3029 = n8354 | n4913;
assign n36 = n4387 & n4162;
assign n5600 = n7391 | n11746;
assign n8036 = ~(n4906 | n9830);
assign n4527 = ~n11876;
assign n7877 = ~(n4283 ^ n10925);
assign n2274 = n6017 | n7056;
assign n9567 = ~(n9203 ^ n66);
assign n5693 = ~(n6640 ^ n9463);
assign n6783 = n10749 | n7229;
assign n4327 = ~n6129;
assign n6745 = n6369 & n3522;
assign n3365 = ~(n8194 | n4035);
assign n207 = ~(n1811 ^ n829);
assign n9123 = n294 & n7023;
assign n11209 = ~(n1809 ^ n8290);
assign n593 = ~(n3441 | n2121);
assign n12921 = ~(n7189 ^ n3107);
assign n8901 = n1472 | n5;
assign n1322 = n5425 & n2245;
assign n10956 = n525 | n8058;
assign n12500 = ~(n9014 | n10933);
assign n7972 = ~(n9708 | n3779);
assign n9933 = n8267 | n11939;
assign n5388 = ~n2166;
assign n7089 = n5919 | n9242;
assign n8189 = n994 | n7424;
assign n1027 = ~(n9307 ^ n1948);
assign n5041 = ~(n6704 ^ n6428);
assign n2032 = ~(n8647 ^ n8408);
assign n8376 = n5205 & n1662;
assign n8715 = ~(n9469 ^ n10314);
assign n8300 = ~(n5323 ^ n9025);
assign n8914 = ~(n10483 ^ n7852);
assign n1275 = n7495 | n11827;
assign n4705 = ~(n5279 ^ n2147);
assign n9710 = ~n12089;
assign n751 = ~(n4301 ^ n11741);
assign n11813 = n5614 & n12895;
assign n7462 = n2099 | n12735;
assign n7251 = n8026 | n995;
assign n7084 = n752 | n11896;
assign n6067 = n7233 & n10059;
assign n3615 = n1514 & n1149;
assign n7919 = n2002 & n12342;
assign n2836 = ~(n196 ^ n11477);
assign n1923 = ~n7342;
assign n7256 = n9110 | n10628;
assign n5381 = ~(n2142 ^ n6216);
assign n518 = ~n2630;
assign n6009 = ~(n885 | n5836);
assign n8692 = n5765 | n8830;
assign n7071 = n10142 | n6402;
assign n2986 = n2982 & n4319;
assign n1260 = n7495 | n7341;
assign n8865 = n8295 & n5242;
assign n8706 = ~(n9450 ^ n11002);
assign n11533 = n10750 | n9586;
assign n8978 = n11026 | n12771;
assign n6251 = n2171 | n10445;
assign n7661 = n1598 | n5564;
assign n2112 = n12116 | n6938;
assign n7255 = ~(n9595 ^ n162);
assign n6427 = ~(n9785 ^ n7764);
assign n1479 = ~(n2542 ^ n12206);
assign n4883 = n7388 & n11876;
assign n1748 = n639 & n1669;
assign n7868 = ~(n5508 ^ n3349);
assign n11971 = n3032 & n281;
assign n5323 = n1764 | n3495;
assign n3157 = n1705 & n12251;
assign n11446 = n11416 & n2535;
assign n2189 = ~n2181;
assign n8286 = n8583 | n4654;
assign n9988 = ~(n3706 | n10461);
assign n4193 = ~n2858;
assign n1710 = n505 & n12592;
assign n883 = ~(n12210 | n601);
assign n11160 = ~(n1988 ^ n4194);
assign n1040 = ~(n6782 ^ n1503);
assign n1003 = ~(n8347 ^ n8488);
assign n5203 = n10697 | n4968;
assign n3488 = ~n11467;
assign n7905 = n5663 & n11387;
assign n9883 = n2466 & n10806;
assign n3451 = ~n1357;
assign n10371 = ~(n10563 ^ n7222);
assign n12349 = ~n11040;
assign n5622 = n11478 & n12925;
assign n9076 = n12227 | n11940;
assign n8305 = ~n8044;
assign n11731 = ~n1750;
assign n8866 = n282 | n7494;
assign n10713 = ~(n10381 ^ n2837);
assign n1106 = n12552 & n6989;
assign n8778 = n8583 | n9568;
assign n6847 = ~n9450;
assign n4573 = ~n6998;
assign n2299 = ~(n1223 ^ n9500);
assign n12028 = ~n8420;
assign n2242 = ~n12915;
assign n10201 = ~(n9476 | n10602);
assign n9201 = ~(n1321 ^ n10886);
assign n7524 = ~(n1921 ^ n12402);
assign n10038 = n191 | n6524;
assign n2747 = ~(n10318 | n10110);
assign n5286 = ~(n7616 ^ n1723);
assign n10025 = n8310 & n2912;
assign n8456 = n5858 | n3911;
assign n184 = ~n11423;
assign n9438 = ~(n2305 ^ n10643);
assign n9557 = ~(n4174 ^ n4470);
assign n8063 = n1699 | n8259;
assign n8772 = n10928 & n7946;
assign n933 = ~(n11413 ^ n5653);
assign n3805 = ~(n11637 ^ n11738);
assign n12671 = ~(n7311 ^ n10151);
assign n1332 = ~(n2842 ^ n6260);
assign n12007 = ~(n4154 | n5746);
assign n11495 = n989 | n6389;
assign n7995 = n6943 & n7182;
assign n3608 = n8622 & n6200;
assign n4050 = ~n1021;
assign n554 = n10774 & n6765;
assign n9353 = n10750 | n3224;
assign n7246 = ~n4005;
assign n7496 = ~(n551 ^ n7975);
assign n9735 = n4628 | n6071;
assign n9487 = ~(n12619 ^ n10166);
assign n4603 = ~(n2878 ^ n10786);
assign n3864 = ~n4678;
assign n5711 = n6740 & n9524;
assign n9784 = ~(n7331 ^ n1865);
assign n7149 = ~n6954;
assign n5574 = ~n7520;
assign n3784 = ~(n3659 | n4993);
assign n11307 = n1882 | n2043;
assign n1887 = n4647 | n11236;
assign n11811 = ~n7289;
assign n10495 = ~(n255 ^ n6879);
assign n3494 = n7662 | n1800;
assign n9827 = n10780 & n12942;
assign n7914 = n11958 | n7558;
assign n2514 = ~(n11664 ^ n8314);
assign n966 = n994 | n12843;
assign n5282 = n11433 | n2815;
assign n11332 = ~(n8376 | n1378);
assign n5076 = n11451 & n6466;
assign n824 = ~n6322;
assign n8472 = ~(n6730 ^ n7510);
assign n4435 = ~(n9263 ^ n8292);
assign n865 = ~(n10191 ^ n9654);
assign n8983 = n12871 & n5649;
assign n7384 = n7462 & n2105;
assign n5360 = n10381 & n6177;
assign n11696 = ~n10857;
assign n1960 = n989 | n1851;
assign n5568 = ~(n7020 ^ n5668);
assign n9341 = n3127 | n1915;
assign n5942 = ~(n11488 ^ n192);
assign n891 = n3820 | n4474;
assign n2430 = n12361 | n5540;
assign n10798 = n11552 | n9521;
assign n2363 = n191 | n12328;
assign n11867 = n9389 | n7341;
assign n2328 = ~(n8592 | n5609);
assign n1915 = ~n7456;
assign n1249 = n191 | n4242;
assign n7602 = ~(n8333 ^ n5446);
assign n3011 = n4805 & n1067;
assign n6708 = ~(n5035 ^ n4003);
assign n5922 = n11958 | n12274;
assign n8258 = n11534 & n483;
assign n9013 = n10389 | n9041;
assign n840 = ~(n11086 ^ n5120);
assign n4320 = ~n12733;
assign n8713 = ~(n9849 | n8268);
assign n9372 = n2312 | n3899;
assign n9232 = n12715 | n7065;
assign n5907 = ~(n4491 ^ n235);
assign n5083 = ~(n7899 ^ n10565);
assign n2637 = ~n11758;
assign n8899 = ~(n5894 ^ n9436);
assign n2359 = n12503 | n9160;
assign n11170 = n3464 & n8805;
assign n3456 = ~(n8160 ^ n7692);
assign n9742 = n6758 | n3387;
assign n7983 = n2456 | n9586;
assign n10519 = ~(n5888 ^ n12923);
assign n4127 = n10960 | n10315;
assign n2969 = ~n2;
assign n2230 = n994 | n561;
assign n4277 = n5510 | n6609;
assign n10611 = ~n5606;
assign n2915 = n4674 | n12535;
assign n10357 = ~(n6012 ^ n5440);
assign n3095 = ~n11594;
assign n12876 = ~(n6009 | n1613);
assign n8195 = n11887 | n8109;
assign n912 = ~(n10768 ^ n328);
assign n1033 = ~(n8146 ^ n5613);
assign n1753 = ~(n4576 ^ n8052);
assign n6162 = n3724 | n53;
assign n7994 = n11850 & n5458;
assign n9835 = ~n250;
assign n8081 = ~(n622 ^ n7987);
assign n774 = ~(n6316 ^ n210);
assign n2176 = ~(n2635 ^ n1232);
assign n9946 = n1699 | n8644;
assign n8774 = ~n6867;
assign n7026 = ~(n10052 | n7353);
assign n9303 = n6373 | n4864;
assign n1234 = ~(n5067 | n12236);
assign n11304 = ~n12573;
assign n11203 = n994 | n4775;
assign n7151 = ~(n8634 ^ n11370);
assign n2891 = ~(n5873 ^ n8867);
assign n2034 = ~n7983;
assign n6862 = ~(n7845 | n5222);
assign n7184 = n12244 | n9425;
assign n4081 = ~(n6919 | n4935);
assign n3496 = ~(n3585 | n6383);
assign n5491 = n7116 | n995;
assign n9441 = n8920 | n8547;
assign n857 = n6331 | n9550;
assign n2135 = ~n531;
assign n3241 = ~(n4806 | n10449);
assign n4740 = n10798 | n10133;
assign n12924 = ~n12266;
assign n4230 = ~(n5447 ^ n4621);
assign n11421 = ~n1810;
assign n2927 = ~n10834;
assign n9578 = ~(n1669 ^ n5142);
assign n10345 = ~(n12204 ^ n1858);
assign n10301 = ~n2321;
assign n35 = ~(n5570 ^ n8963);
assign n3408 = n8601 | n2737;
assign n3514 = ~(n2190 ^ n2663);
assign n9491 = ~(n12377 ^ n8881);
assign n9511 = ~(n10830 | n1631);
assign n9785 = n11552 | n4875;
assign n6583 = n9751 | n10758;
assign n1124 = ~(n1826 ^ n8280);
assign n10648 = n2380 & n8177;
assign n10717 = n10163 | n10321;
assign n9694 = ~n5845;
assign n11316 = ~n5978;
assign n9109 = ~(n1715 ^ n2961);
assign n12655 = ~n7442;
assign n2029 = ~(n3180 ^ n10086);
assign n11082 = ~n167;
assign n6186 = n8480 & n5865;
assign n9901 = ~(n4948 ^ n11275);
assign n6230 = n10424 | n7245;
assign n834 = ~n990;
assign n8694 = n7449 | n5502;
assign n7185 = n12119 | n8259;
assign n3573 = ~(n2 | n11783);
assign n10818 = n12263 | n9203;
assign n12919 = ~(n2570 ^ n5038);
assign n7535 = ~(n12286 ^ n11836);
assign n10191 = n9730 & n3306;
assign n6580 = ~(n10324 ^ n7333);
assign n6790 = n12341 | n3075;
assign n2739 = n12199 & n4028;
assign n8750 = n10762 & n11365;
assign n630 = n8598 & n5581;
assign n10790 = n1183 | n3224;
assign n10280 = n3066 & n8669;
assign n8549 = n2791 | n278;
assign n12396 = n11245 & n2673;
assign n3560 = n3905 & n2270;
assign n7655 = n10157 | n4864;
assign n8143 = n4916 | n1263;
assign n5 = ~(n11790 ^ n2280);
assign n11324 = n8026 | n7558;
assign n6661 = n1941 | n5540;
assign n6704 = n6373 | n9521;
assign n6749 = n58 & n12426;
assign n12224 = ~(n11721 ^ n4146);
assign n3056 = n5990 & n11078;
assign n3340 = n11026 | n1476;
assign n5781 = ~n1353;
assign n5048 = n10360 & n12013;
assign n6170 = ~n1306;
assign n11655 = ~n12219;
assign n5773 = ~n12520;
assign n4948 = n8870 | n5326;
assign n12384 = ~n11884;
assign n5974 = ~n7778;
assign n11387 = n9426 | n5790;
assign n651 = ~n8048;
assign n8608 = ~n7151;
assign n10993 = n6671 | n4526;
assign n6188 = ~(n8013 ^ n1075);
assign n8037 = ~(n8162 | n9845);
assign n3679 = ~n7187;
assign n12023 = n752 | n3421;
assign n11997 = n1796 & n10623;
assign n12445 = ~(n3794 ^ n12285);
assign n8342 = n2052 & n1367;
assign n4288 = ~n6879;
assign n3957 = n6738 & n11179;
assign n5968 = ~(n11182 ^ n4200);
assign n12061 = n1699 | n8109;
assign n2471 = ~(n1991 ^ n6692);
assign n3281 = ~(n8602 ^ n5897);
assign n2569 = n11511 & n6885;
assign n1645 = n12647 ^ n10665;
assign n7229 = ~(n12742 ^ n11768);
assign n12353 = ~(n8515 ^ n6760);
assign n5564 = n3892 | n10358;
assign n1502 = n11528 & n2654;
assign n12309 = ~(n11908 ^ n7578);
assign n6927 = ~(n8155 | n4408);
assign n12751 = ~(n9059 ^ n6865);
assign n11267 = n4056 & n2169;
assign n11585 = ~(n3837 ^ n9096);
assign n11840 = n10670 & n5488;
assign n4596 = n1100 | n7763;
assign n11785 = n7688 & n11465;
assign n11567 = n7587 | n2343;
assign n12830 = n2697 & n11348;
assign n11411 = ~n2470;
assign n11073 = ~(n1782 ^ n12598);
assign n12172 = ~n6660;
assign n3225 = ~(n10909 | n3496);
assign n9577 = ~(n1956 ^ n8570);
assign n3907 = n1993 | n5090;
assign n11747 = n5840 | n6614;
assign n5134 = n11036 | n8030;
assign n11210 = ~(n4489 ^ n7013);
assign n12598 = ~n4834;
assign n11037 = n8870 | n4913;
assign n2811 = n1653 & n10896;
assign n12030 = ~n4999;
assign n12324 = n11958 | n8768;
assign n5973 = n7889 & n11993;
assign n5421 = ~(n9764 ^ n3997);
assign n555 = n3011 & n8660;
assign n10054 = ~(n3369 | n9471);
assign n7422 = ~n10009;
assign n3308 = n7251 & n4264;
assign n12417 = n2045 & n11274;
assign n1521 = n4696 | n2475;
assign n6048 = ~n3824;
assign n2729 = ~(n9522 ^ n2205);
assign n1021 = n11283 | n12773;
assign n4205 = n1941 | n7876;
assign n11167 = ~(n10560 ^ n2889);
assign n7018 = ~(n4942 ^ n7580);
assign n1746 = n10835 | n8285;
assign n4834 = n2530 & n2802;
assign n5523 = ~n5291;
assign n5786 = n7283 | n5497;
assign n8696 = ~(n11029 ^ n10800);
assign n8590 = n8687 | n28;
assign n1163 = ~n11922;
assign n10298 = ~(n9489 | n8935);
assign n4295 = n167 | n408;
assign n6592 = n2025 | n5322;
assign n6115 = n12262 | n8253;
assign n3025 = ~n5728;
assign n3759 = ~n2714;
assign n12819 = n8949 | n6724;
assign n12297 = ~n7331;
assign n2214 = n8332 | n10866;
assign n7014 = n11550 | n7051;
assign n5494 = ~(n10257 | n8868);
assign n4049 = ~(n4212 ^ n1485);
assign n4769 = n4176 | n3948;
assign n11442 = ~(n6464 ^ n9143);
assign n7473 = n8848 | n1008;
assign n9322 = n6718 | n4474;
assign n794 = n2950 & n1164;
assign n11555 = ~(n12445 ^ n1351);
assign n8842 = ~n4028;
assign n375 = ~n11834;
assign n2127 = n10157 | n12771;
assign n3556 = ~n625;
assign n336 = ~(n7978 ^ n4997);
assign n7954 = n5283 & n521;
assign n950 = ~(n6221 ^ n11379);
assign n11184 = n3096 | n1413;
assign n43 = n925 & n1958;
assign n10902 = n9655 | n12580;
assign n6526 = ~n10243;
assign n11923 = ~n5314;
assign n3548 = ~n1822;
assign n12541 = n9400 & n10439;
assign n10527 = n3324 | n4527;
assign n8949 = n5575 | n3468;
assign n1535 = ~(n6954 ^ n3812);
assign n8110 = ~(n3079 ^ n9237);
assign n1600 = ~n1294;
assign n11856 = n8428 | n9741;
assign n8101 = n1760 & n2859;
assign n11188 = ~(n5277 ^ n6240);
assign n3723 = ~(n12354 ^ n7165);
assign n3873 = n6977 | n5538;
assign n11225 = n12069 & n1512;
assign n102 = n4734 & n11489;
assign n6318 = n1941 | n1413;
assign n8993 = ~(n10945 ^ n5348);
assign n5631 = ~n2030;
assign n10443 = n4150 & n4627;
assign n11903 = ~(n11831 | n12798);
assign n1253 = ~n812;
assign n11146 = ~(n12935 ^ n9808);
assign n8455 = n6411 & n4132;
assign n2905 = n8026 | n6114;
assign n7072 = ~(n2726 ^ n3289);
assign n12862 = n10712 | n5583;
assign n9193 = n1226 & n2750;
assign n1962 = n10135 | n9854;
assign n11321 = n4120 & n2805;
assign n9674 = n191 | n1738;
assign n7132 = ~(n3387 ^ n12334);
assign n8174 = ~(n2567 ^ n2455);
assign n3371 = ~(n2928 ^ n12650);
assign n11619 = ~n11017;
assign n1391 = ~n2937;
assign n11230 = n10772 & n10793;
assign n10273 = ~(n10997 ^ n10940);
assign n6500 = ~(n3936 ^ n1946);
assign n10264 = ~(n8176 ^ n324);
assign n3802 = ~(n10722 ^ n5535);
assign n2633 = n7084 & n9091;
assign n10929 = n3820 | n28;
assign n4581 = n3316 & n7888;
assign n11255 = n2155 | n11112;
assign n4204 = ~n3247;
assign n9038 = n2718 & n4611;
assign n577 = n8354 | n826;
assign n103 = ~(n3130 ^ n7555);
assign n4365 = ~n5263;
assign n10778 = n4383 | n6297;
assign n4812 = n10590 | n7821;
assign n1829 = n6373 | n7921;
assign n1517 = ~(n3970 ^ n7091);
assign n12663 = ~(n11080 | n12597);
assign n11473 = ~n3825;
assign n12957 = ~n7807;
assign n1208 = ~(n4788 | n9620);
assign n5987 = ~(n5492 ^ n10072);
assign n6495 = ~(n5921 ^ n7360);
assign n7476 = ~n6527;
assign n9074 = ~n5582;
assign n7934 = ~(n2993 ^ n6468);
assign n12539 = n7116 | n11896;
assign n4163 = ~(n9926 ^ n1969);
assign n7372 = ~(n9305 | n6205);
assign n5233 = n5964 & n2577;
assign n3659 = n5575 | n6114;
assign n11228 = ~n2443;
assign n12070 = n6893 & n1068;
assign n6240 = ~(n5087 ^ n5357);
assign n8779 = n8026 | n12816;
assign n11445 = ~(n9613 ^ n4425);
assign n9465 = n4312 & n7456;
assign n9413 = n11958 | n995;
assign n1203 = ~(n10703 ^ n12311);
assign n7197 = ~(n9438 | n8982);
assign n4076 = ~(n12176 ^ n7150);
assign n11392 = n6718 | n5502;
assign n12852 = ~(n9043 ^ n10840);
assign n6729 = n3848 & n4974;
assign n7769 = ~(n9643 | n10076);
assign n8054 = n1937 | n6169;
assign n10868 = n5832 & n6531;
assign n6815 = ~(n6341 ^ n4419);
assign n6463 = n3007 | n8561;
assign n60 = n11958 | n6084;
assign n478 = n8337 & n5622;
assign n2884 = ~(n10918 ^ n6420);
assign n8361 = ~(n9392 ^ n7263);
assign n9964 = n1223 & n2892;
assign n11638 = ~n12564;
assign n4699 = n11572 | n3192;
assign n10518 = n6718 | n9160;
assign n7687 = ~n2643;
assign n692 = ~n8694;
assign n5402 = ~n1481;
assign n12079 = ~n649;
assign n6853 = n962 | n28;
assign n9589 = ~n9725;
assign n5797 = n9370 | n1162;
assign n5971 = n6914 & n4447;
assign n1056 = ~(n2763 ^ n12633);
assign n11456 = n3617 | n10854;
assign n2685 = ~(n12960 ^ n10487);
assign n3680 = ~(n9722 ^ n3739);
assign n8156 = n9360 & n7633;
assign n2247 = n4859 & n2263;
assign n7565 = ~(n10615 ^ n4523);
assign n9331 = n7872 & n9468;
assign n2846 = n2099 | n4249;
assign n2461 = n8737 & n5874;
assign n12715 = ~(n10866 ^ n8332);
assign n10760 = ~n12360;
assign n6330 = ~(n12533 ^ n9996);
assign n7556 = ~(n1642 ^ n6707);
assign n3334 = ~(n5301 | n8701);
assign n1553 = ~(n8390 ^ n757);
assign n6636 = ~n11844;
assign n4196 = n12146 & n10609;
assign n1615 = ~(n9130 ^ n9279);
assign n10467 = n4628 | n12124;
assign n10272 = ~(n10769 ^ n2241);
assign n7886 = n10108 | n11746;
assign n3055 = ~(n8111 ^ n9012);
assign n10000 = ~(n6466 ^ n6079);
assign n12078 = ~n8913;
assign n12442 = ~n10560;
assign n348 = n5589 | n11291;
assign n6766 = n12256 | n195;
assign n6406 = n2968 ^ n4306;
assign n3540 = ~n382;
assign n9913 = n636 | n6071;
assign n5398 = n3389 & n10001;
assign n11281 = n12119 | n12754;
assign n7998 = n5575 | n11820;
assign n12267 = n9705 & n971;
assign n11410 = ~n10451;
assign n5676 = ~(n4500 ^ n3469);
assign n10245 = ~(n1331 ^ n12919);
assign n4020 = ~(n8920 ^ n295);
assign n12459 = ~(n7176 ^ n506);
assign n10156 = n7986 | n968;
assign n234 = ~(n8778 ^ n955);
assign n8010 = ~n83;
assign n4000 = ~(n10808 ^ n2529);
assign n2055 = n5876 & n5307;
assign n10406 = ~(n4387 ^ n4894);
assign n7689 = ~(n84 | n9350);
assign n5900 = ~(n1364 ^ n1517);
assign n9747 = ~(n885 ^ n5836);
assign n2028 = ~(n7672 ^ n220);
assign n792 = n7090 | n7255;
assign n7104 = ~(n1863 | n11916);
assign n8657 = ~(n10143 ^ n909);
assign n3879 = ~(n5736 ^ n9955);
assign n9493 = ~(n7088 ^ n2926);
assign n8076 = ~(n7775 ^ n8490);
assign n12483 = ~(n774 | n5608);
assign n12599 = n9389 | n7246;
assign n6607 = ~n12611;
assign n2244 = n1144 & n5210;
assign n4773 = ~n4390;
assign n12766 = n7169 & n1238;
assign n1026 = n1215 | n5055;
assign n11599 = ~n12893;
assign n2040 = n6073 | n8947;
assign n894 = n7449 | n9160;
assign n4680 = ~(n7355 ^ n5444);
assign n12233 = ~(n324 | n5686);
assign n6606 = n12361 | n8414;
assign n3277 = n11241 | n7689;
assign n2824 = n4805 & n5645;
assign n6517 = ~(n11268 ^ n3525);
assign n6443 = ~(n4570 ^ n9874);
assign n9593 = n6231 & n3444;
assign n4835 = ~n7784;
assign n174 = ~(n6575 | n9458);
assign n12146 = n1803 | n6421;
assign n2424 = n12119 | n7382;
assign n5315 = ~(n1315 ^ n2211);
assign n12838 = ~(n7112 ^ n12654);
assign n6564 = n3743 | n8745;
assign n7936 = ~(n4409 ^ n11220);
assign n10458 = n994 | n11746;
assign n1563 = n9519 & n9023;
assign n2453 = n4737 | n5932;
assign n1698 = ~(n1653 ^ n10896);
assign n11363 = n2072 & n3908;
assign n10426 = ~n12452;
assign n9476 = n10879 | n6389;
assign n8380 = n4697 & n6968;
assign n5032 = n6418 | n729;
assign n1711 = ~(n11056 | n1535);
assign n10999 = ~(n5194 | n8710);
assign n11843 = ~n12052;
assign n804 = n1937 | n10903;
assign n4463 = n5964 & n9956;
assign n9780 = n3995 | n482;
assign n8523 = ~n5353;
assign n1455 = ~n9956;
assign n4456 = ~n758;
assign n5754 = n6307 & n4636;
assign n9324 = ~(n11836 | n12286);
assign n1390 = ~(n10307 ^ n999);
assign n1235 = n4892 & n583;
assign n11108 = ~(n2640 ^ n12181);
assign n7878 = ~(n7130 ^ n11464);
assign n8325 = n3820 | n8830;
assign n5648 = ~(n386 ^ n9354);
assign n386 = n8026 | n7952;
assign n3646 = n1701 & n3338;
assign n11431 = n9180 | n11564;
assign n236 = n5530 | n6071;
assign n5498 = ~(n5608 ^ n774);
assign n11915 = ~(n2363 ^ n10097);
assign n6408 = n9644 & n4925;
assign n10372 = ~(n12737 | n1742);
assign n946 = ~(n4808 ^ n2166);
assign n2851 = n5283 & n6254;
assign n621 = n9878 | n8655;
assign n4977 = n7203 & n3304;
assign n83 = n6706 & n10702;
assign n5506 = ~n11972;
assign n8425 = ~(n3203 ^ n9601);
assign n10543 = ~(n3733 | n8200);
assign n4947 = n12610 & n7794;
assign n9328 = n10879 | n1851;
assign n561 = ~n10327;
assign n9116 = ~(n1082 ^ n11336);
assign n10206 = n12616 | n10627;
assign n7981 = ~(n11730 ^ n6215);
assign n12362 = n636 | n8648;
assign n844 = ~(n2607 ^ n5472);
assign n10584 = n5211 & n9287;
assign n7434 = n2456 | n12446;
assign n327 = ~(n788 ^ n12009);
assign n10334 = n12496 & n10286;
assign n8454 = ~n10870;
assign n292 = ~(n433 ^ n11705);
assign n658 = ~(n10146 ^ n1522);
assign n1248 = ~(n5382 ^ n2905);
assign n8066 = n4498 | n4400;
assign n6470 = n5530 | n12735;
assign n5104 = ~(n2922 | n5244);
assign n1942 = ~(n9124 ^ n11629);
assign n6324 = ~(n3145 ^ n1267);
assign n114 = ~n12753;
assign n9445 = ~n12562;
assign n2907 = n12061 | n10900;
assign n5849 = ~(n7762 ^ n1213);
assign n10405 = ~(n643 | n11979);
assign n11579 = n2313 | n2669;
assign n5578 = ~(n5021 ^ n1414);
assign n10660 = n3947 | n172;
assign n9041 = ~(n891 ^ n4598);
assign n1839 = n11245 | n2673;
assign n1776 = n9370 | n7703;
assign n12470 = n1941 | n10903;
assign n8880 = n10139 | n3615;
assign n7714 = ~n8160;
assign n10731 = n7337 | n3400;
assign n12569 = n9365 & n3307;
assign n439 = n596 | n5716;
assign n9551 = n5503 & n730;
assign n7644 = ~(n5214 ^ n2616);
assign n3852 = n4203 & n7354;
assign n5468 = ~n2498;
assign n7562 = n6003 | n11614;
assign n4940 = n6385 | n8468;
assign n10030 = n9112 | n8186;
assign n11472 = ~n7531;
assign n12422 = n1082 & n919;
assign n11600 = ~(n1662 ^ n6713);
assign n433 = ~(n5217 ^ n9200);
assign n932 = ~(n5039 ^ n12358);
assign n2688 = ~(n11714 ^ n4251);
assign n11831 = n6101 ^ n2023;
assign n11569 = n7391 | n1455;
assign n7472 = ~(n6584 ^ n12702);
assign n11427 = ~(n5685 ^ n5658);
assign n7838 = ~(n5761 ^ n5831);
assign n5199 = ~n2436;
assign n8457 = ~(n161 ^ n550);
assign n6891 = ~(n12362 ^ n9811);
assign n7409 = n1699 | n3224;
assign n11550 = ~(n6060 ^ n299);
assign n12609 = ~(n11633 ^ n9647);
assign n5738 = ~n8906;
assign n3970 = n5462 & n4080;
assign n7923 = ~(n9698 ^ n12540);
assign n12742 = n5530 | n8644;
assign n9311 = n3992 & n159;
assign n9002 = ~(n5899 | n2928);
assign n2935 = ~n2943;
assign n6061 = ~(n1750 ^ n2500);
assign n4877 = n4872 & n12374;
assign n12773 = n947 & n6533;
assign n2416 = ~(n2933 ^ n9760);
assign n12428 = ~(n1309 ^ n9602);
assign n9357 = n11626 | n12763;
assign n10979 = n12495 & n4729;
assign n7761 = ~(n5525 ^ n5552);
assign n7458 = n5945 | n12816;
assign n1548 = n5355 | n3911;
assign n11710 = n807 | n1413;
assign n12099 = n3872 & n2814;
assign n11980 = ~n4314;
assign n3547 = ~(n3790 ^ n4106);
assign n1412 = n6091 & n6855;
assign n11094 = ~(n10493 ^ n9947);
assign n4616 = ~(n9943 ^ n4488);
assign n5701 = n9190 & n8079;
assign n7250 = n6525 | n2860;
assign n9182 = n1990 | n7635;
assign n11168 = ~n3401;
assign n8343 = n9373 | n1476;
assign n12732 = ~(n8594 | n10081);
assign n9846 = n5355 | n8735;
assign n12302 = n7709 | n4474;
assign n9499 = n6876 & n6818;
assign n6515 = n8187 | n510;
assign n12284 = n2099 | n10422;
assign n11933 = n3974 & n2041;
assign n7817 = ~(n3210 | n10527);
assign n11846 = n7449 | n9568;
assign n10194 = n910 & n9852;
assign n4225 = n9002 | n2114;
assign n2383 = ~(n8811 ^ n9774);
assign n3735 = ~n8235;
assign n12462 = n4911 | n1546;
assign n7065 = ~(n1878 | n11494);
assign n6196 = n12447 | n4665;
assign n6706 = n5331 & n12489;
assign n1265 = n10542 & n5178;
assign n11519 = ~n12505;
assign n12108 = ~(n2482 ^ n2163);
assign n6313 = n11808 | n1838;
assign n6154 = ~n12448;
assign n1215 = n9389 | n1851;
assign n9789 = ~(n12368 | n7583);
assign n6969 = ~n11173;
assign n12404 = n11375 & n6144;
assign n3813 = ~n233;
assign n8862 = ~(n4002 ^ n6061);
assign n2385 = ~(n613 ^ n836);
assign n11545 = ~(n5164 ^ n513);
assign n8166 = ~(n434 | n11871);
assign n10532 = n5724 | n8890;
assign n11842 = n5530 | n10854;
assign n3940 = n12289 | n9253;
assign n4493 = ~n3852;
assign n10474 = n9803 | n6160;
assign n2697 = n2761 | n6288;
assign n3690 = ~n12480;
assign n10102 = n6249 | n251;
assign n2350 = n9208 & n12696;
assign n7659 = ~n10450;
assign n11793 = ~n10845;
assign n9790 = ~(n11335 ^ n12278);
assign n732 = ~n49;
assign n1192 = n12661 & n2753;
assign n3590 = ~n6974;
assign n7751 = ~(n3176 ^ n10322);
assign n152 = ~(n7446 ^ n1023);
assign n12118 = n5915 | n12735;
assign n11784 = ~(n11482 ^ n10635);
assign n7045 = ~(n12607 | n10204);
assign n515 = n4628 | n4818;
assign n8963 = n6577 | n7425;
assign n10169 = n10835 | n12120;
assign n6275 = n8103 | n5741;
assign n6647 = ~(n8550 ^ n10934);
assign n4744 = n11189 & n7922;
assign n2538 = ~n12122;
assign n6731 = ~(n7059 ^ n3835);
assign n734 = ~n10972;
assign n7682 = n3188 & n689;
assign n8944 = ~n3904;
assign n12577 = ~n1275;
assign n7790 = n2217 | n2020;
assign n1692 = ~(n6231 ^ n12103);
assign n5120 = ~(n10773 ^ n490);
assign n12828 = ~(n3795 ^ n8868);
assign n2834 = ~(n6539 ^ n47);
assign n12420 = ~(n3301 ^ n691);
assign n7784 = ~(n12933 ^ n8989);
assign n6503 = ~(n3544 ^ n3414);
assign n10337 = ~n1124;
assign n11539 = n5231 | n5217;
assign n9865 = ~(n8869 ^ n12806);
assign n12614 = ~n2305;
assign n12627 = ~(n2005 ^ n3331);
assign n11171 = n3096 | n7425;
assign n3495 = n693 & n3069;
assign n3439 = n240 & n983;
assign n3780 = n9098 | n2812;
assign n3914 = ~(n9198 ^ n8640);
assign n4917 = ~(n9479 ^ n12515);
assign n3906 = n191 | n5851;
assign n4139 = ~(n9042 ^ n11399);
assign n4637 = n5225 | n1625;
assign n4201 = n12284 | n663;
assign n685 = ~n6002;
assign n5659 = n11060 & n11247;
assign n9075 = ~(n11842 ^ n7027);
assign n12461 = n148 & n3927;
assign n2467 = ~(n772 ^ n2645);
assign n6870 = ~(n6800 | n8436);
assign n393 = n719 & n6314;
assign n10129 = ~(n8015 | n12716);
assign n6435 = ~(n2136 ^ n10652);
assign n12800 = ~(n8444 | n6693);
assign n6545 = ~(n6805 ^ n869);
assign n5615 = ~(n7122 ^ n746);
assign n3980 = n1126 | n4143;
assign n5118 = ~(n11240 | n3993);
assign n6260 = n10829 & n3589;
assign n3523 = n10835 | n3599;
assign n4385 = ~(n6939 ^ n208);
assign n10676 = ~(n203 ^ n8447);
assign n531 = ~(n6453 ^ n7412);
assign n120 = ~n8093;
assign n7907 = ~(n7567 ^ n11794);
assign n604 = n19 & n4533;
assign n11145 = n2014 & n9821;
assign n11601 = n4223 | n1819;
assign n2760 = n8459 & n11573;
assign n4644 = n3743 | n4875;
assign n10098 = ~n12047;
assign n7467 = ~(n6318 ^ n7064);
assign n4982 = ~(n11514 | n3012);
assign n9198 = n12485 | n7670;
assign n6554 = ~(n8231 ^ n11135);
assign n945 = n11195 & n9292;
assign n8317 = n9584 | n2020;
assign n3256 = n4846 | n11562;
assign n4736 = ~n578;
assign n11408 = ~(n12524 ^ n2088);
assign n9542 = ~(n12309 ^ n10651);
assign n10511 = n2170 & n1897;
assign n5712 = n11433 | n9741;
assign n672 = ~(n1346 ^ n5163);
assign n9940 = n10879 | n1162;
assign n11559 = ~(n10693 ^ n8709);
assign n11929 = ~(n9897 ^ n979);
assign n11476 = ~(n9486 | n1264);
assign n8449 = n8026 | n8768;
assign n10959 = ~(n7075 ^ n4746);
assign n6713 = ~(n5205 ^ n3949);
assign n6599 = n9389 | n1546;
assign n1878 = n11560 | n9658;
assign n12528 = n5516 & n6719;
assign n7978 = ~(n3283 ^ n2849);
assign n6125 = ~(n709 | n1568);
assign n2374 = n2832 | n5497;
assign n12668 = n7449 | n5914;
assign n9102 = n7690 & n2558;
assign n6397 = ~(n1028 | n5924);
assign n7345 = n8256 & n2373;
assign n11798 = ~(n11669 ^ n652);
assign n8436 = ~(n5532 ^ n8501);
assign n8647 = ~(n11514 ^ n7727);
assign n10144 = n12853 | n12535;
assign n9990 = n1475 | n4986;
assign n5094 = ~(n11491 ^ n12222);
assign n8294 = n11958 | n184;
assign n4132 = n6134 | n12401;
assign n6685 = ~(n3354 | n7607);
assign n7841 = ~n7631;
assign n5824 = n12864 | n9456;
assign n3524 = n11968 & n6;
assign n7200 = n989 | n12328;
assign n12727 = n10398 & n1601;
assign n11636 = ~(n722 ^ n10325);
assign n10556 = ~(n5079 ^ n10084);
assign n11598 = n7449 | n28;
assign n4028 = n2464 & n5105;
assign n2839 = n6782 & n7054;
assign n9815 = ~n820;
assign n4507 = ~(n688 ^ n7853);
assign n6253 = ~(n4907 ^ n8766);
assign n581 = n10945 & n7318;
assign n9909 = n9382 & n3760;
assign n9307 = n752 | n6169;
assign n10847 = n5355 | n1079;
assign n1324 = n8476 & n1564;
assign n4889 = ~(n6861 | n10985);
assign n4804 = n9313 & n190;
assign n4397 = n165 ^ n6990;
assign n9266 = n4628 | n12080;
assign n12215 = ~(n12603 ^ n8696);
assign n1677 = n8996 | n9518;
assign n923 = ~(n11800 ^ n7358);
assign n3279 = n12365 | n11406;
assign n3599 = ~n1906;
assign n11402 = n11493 | n8122;
assign n1589 = ~(n9391 ^ n5302);
assign n7194 = ~(n9114 ^ n11581);
assign n8245 = ~(n1205 ^ n5617);
assign n10284 = n11740 & n4969;
assign n5730 = ~(n3202 ^ n8683);
assign n8598 = ~(n2440 ^ n9261);
assign n11310 = n3243 & n5880;
assign n10963 = n1282 & n12458;
assign n1586 = ~(n8840 ^ n11315);
assign n7884 = n6656 | n9548;
assign n3504 = n7398 & n12219;
assign n12246 = n8738 | n9160;
assign n2212 = ~(n10112 | n12547);
assign n11746 = ~n3932;
assign n2171 = ~n8521;
assign n9001 = ~(n418 ^ n207);
assign n11808 = ~(n6954 | n4912);
assign n9261 = n12194 & n2351;
assign n5650 = n10835 | n6138;
assign n7387 = ~(n8737 ^ n6644);
assign n6522 = n6271 | n11420;
assign n5387 = n5858 | n4400;
assign n10211 = n10387 & n3019;
assign n10756 = n2010 & n2261;
assign n9929 = ~(n3694 ^ n1849);
assign n7815 = ~(n12071 ^ n11230);
assign n9257 = ~(n12177 ^ n2430);
assign n8592 = ~n6584;
assign n6490 = ~n5093;
assign n1095 = n12701 | n6897;
assign n10208 = n11547 & n6832;
assign n8910 = n6686 & n5407;
assign n2118 = n11162 & n1302;
assign n9403 = n11936 & n3346;
assign n8281 = n11478 & n1564;
assign n1109 = n9266 & n8711;
assign n8233 = n2319 & n10252;
assign n12166 = n4950 & n2596;
assign n11872 = ~(n8892 ^ n8906);
assign n7673 = ~n9348;
assign n6587 = n4741 ^ n7253;
assign n1147 = n12438 & n8185;
assign n10989 = ~(n10880 ^ n7361);
assign n12519 = ~(n7248 ^ n12159);
assign n3134 = n8516 ^ n4682;
assign n2571 = n7166 & n11163;
assign n5422 = n8010 | n12089;
assign n7607 = ~n4427;
assign n413 = n3381 | n10811;
assign n12427 = ~n10802;
assign n3643 = n8816 & n1084;
assign n12142 = n2456 | n7382;
assign n3508 = n5575 | n2589;
assign n1174 = n8959 | n5012;
assign n7507 = ~(n8389 ^ n10747);
assign n5628 = ~(n6008 ^ n4581);
assign n677 = n7452 | n8615;
assign n12729 = n443 & n10200;
assign n10508 = n7911 & n5323;
assign n3860 = ~(n23 | n7844);
assign n8591 = ~(n1438 ^ n6778);
assign n3843 = n114 | n5012;
assign n5375 = ~(n7230 | n11019);
assign n4092 = n10354 & n1502;
assign n3520 = n12853 | n5468;
assign n9164 = n4778 | n5468;
assign n6844 = n11887 | n10854;
assign n673 = ~n1317;
assign n8937 = n12220 & n6388;
assign n4346 = n1941 | n6197;
assign n1444 = n11851 | n9255;
assign n11346 = ~n12355;
assign n5097 = ~(n2411 | n8486);
assign n11759 = ~n4930;
assign n7590 = n6971 | n7178;
assign n8872 = ~(n6581 ^ n12820);
assign n9663 = ~(n11988 ^ n2374);
assign n1797 = ~(n8938 | n578);
assign n7423 = n4457 & n622;
assign n8921 = ~n2760;
assign n5894 = ~(n3481 ^ n575);
assign n4611 = ~n6838;
assign n1012 = n191 | n6402;
assign n12923 = ~(n2019 ^ n462);
assign n193 = ~(n8452 ^ n8978);
assign n4219 = n1449 | n1174;
assign n5184 = ~(n11442 ^ n728);
assign n7325 = n9373 | n9078;
assign n11995 = ~(n6594 | n6670);
assign n1411 = ~(n1924 ^ n10014);
assign n5075 = ~(n9718 ^ n3738);
assign n7559 = ~(n7325 ^ n8325);
assign n11671 = n3594 & n7156;
assign n7016 = ~(n3483 ^ n12894);
assign n10659 = n9421 & n1885;
assign n437 = n10429 | n7158;
assign n1802 = n10064 & n10905;
assign n7445 = n7537 | n4803;
assign n2421 = n5800 & n738;
assign n10227 = ~(n12198 ^ n4024);
assign n5570 = n8428 | n11122;
assign n8740 = ~n1067;
assign n11714 = n8870 | n12535;
assign n6738 = n9389 | n7424;
assign n3065 = n5809 | n3924;
assign n11755 = ~(n5327 ^ n11912);
assign n6494 = ~(n12895 ^ n1834);
assign n1882 = n3717 | n1894;
assign n4764 = ~n9072;
assign n703 = ~(n5049 ^ n958);
assign n11315 = ~(n3346 ^ n3242);
assign n6072 = n6718 | n9568;
assign n1740 = n8428 | n6114;
assign n12141 = n10512 & n2742;
assign n10986 = ~n9805;
assign n9939 = n6136 | n5835;
assign n4326 = ~(n5978 ^ n10597);
assign n7809 = n3628 | n894;
assign n3782 = n2608 & n4615;
assign n12383 = ~(n9258 ^ n2584);
assign n12615 = ~(n11490 ^ n10318);
assign n6493 = ~n9467;
assign n12080 = ~n5579;
assign n10330 = ~n1984;
assign n9508 = ~(n11208 ^ n1911);
assign n8532 = n1371 & n6392;
assign n10061 = ~(n11955 ^ n1819);
assign n4242 = ~n4370;
assign n7398 = ~n7206;
assign n4195 = n12186 | n6455;
assign n11563 = n10835 | n4654;
assign n362 = ~n3715;
assign n754 = ~(n10582 | n6998);
assign n1837 = n7773 & n1633;
assign n6754 = ~(n3711 ^ n912);
assign n12875 = n3240 & n8801;
assign n11221 = n10142 | n7424;
assign n4156 = ~(n1021 ^ n3502);
assign n6555 = ~(n1258 ^ n7250);
assign n12266 = n9739 & n7224;
assign n10725 = n9266 | n8711;
assign n1806 = n7839 | n5012;
assign n1796 = ~n6370;
assign n11863 = ~n12292;
assign n2869 = ~(n11575 ^ n9057);
assign n1783 = n12891 | n11506;
assign n2763 = n5355 | n1851;
assign n5311 = ~n783;
assign n11857 = ~n11271;
assign n271 = n9389 | n12843;
assign n8055 = n191 | n10419;
assign n3180 = n10879 | n7341;
assign n11787 = n12525 & n3298;
assign n4851 = n8327 & n2701;
assign n9454 = n4600 & n410;
assign n5397 = n5809 | n6513;
assign n10047 = n8720 & n12064;
assign n10126 = ~(n7653 ^ n4688);
assign n12661 = n914 | n2429;
assign n12951 = ~(n2539 ^ n5910);
assign n4953 = n5305 & n5212;
assign n6007 = n12051 & n3091;
assign n10899 = n5501 | n4792;
assign n3422 = n12070 | n2621;
assign n1988 = n6158 | n3052;
assign n3896 = n9081 & n6258;
assign n998 = n11324 | n12756;
assign n11372 = ~(n7793 ^ n536);
assign n12840 = n7865 | n12338;
assign n319 = ~(n9455 | n513);
assign n7990 = ~(n2058 ^ n4218);
assign n7699 = n12063 & n12149;
assign n10328 = ~(n1810 ^ n7990);
assign n6996 = ~(n10404 ^ n1132);
assign n2588 = ~(n9270 ^ n6356);
assign n1524 = n1516 & n2189;
assign n4090 = ~(n1371 ^ n690);
assign n10629 = ~n6760;
assign n10316 = ~n3094;
assign n6695 = n3746 | n5012;
assign n9757 = n12936 & n6796;
assign n1603 = ~(n9492 ^ n4546);
assign n6999 = ~n9167;
assign n9709 = ~n2089;
assign n6056 = ~(n1947 ^ n3151);
assign n12716 = n10093 | n12105;
assign n4840 = ~(n12198 | n1562);
assign n2324 = n6767 | n6250;
assign n7744 = ~(n6853 | n5076);
assign n12482 = ~(n9443 ^ n7377);
assign n2626 = n8428 | n11820;
assign n1864 = ~(n5907 ^ n5343);
assign n10070 = ~n10844;
assign n4266 = n1549 | n10856;
assign n9163 = ~(n3135 ^ n11057);
assign n8728 = ~(n2071 ^ n10323);
assign n12278 = n10157 | n7921;
assign n12115 = n9707 & n6526;
assign n11658 = n1779 | n4685;
assign n4497 = ~(n5661 ^ n7164);
assign n390 = n10962 & n9333;
assign n2178 = n1341 & n9522;
assign n9809 = ~(n11069 ^ n11128);
assign n9505 = ~n1240;
assign n12743 = n7709 | n4654;
assign n1493 = n9370 | n2358;
assign n867 = ~(n12269 | n7003);
assign n3347 = ~n10648;
assign n12045 = n8369 | n4108;
assign n9518 = n1699 | n826;
assign n793 = ~(n935 ^ n606);
assign n820 = n994 | n4400;
assign n11778 = n4237 | n10229;
assign n3167 = ~(n11339 ^ n9224);
assign n2067 = ~n20;
assign n4255 = n9037 | n448;
assign n11451 = n3820 | n3606;
assign n7594 = ~(n7756 | n4681);
assign n5205 = n8755 & n6648;
assign n11921 = ~(n12226 ^ n6340);
assign n11365 = n11892 & n7294;
assign n2651 = ~(n3353 | n5545);
assign n1994 = n5964 & n1798;
assign n10703 = ~(n11704 ^ n2368);
assign n9917 = ~n10488;
assign n4743 = ~(n8828 ^ n4123);
assign n4261 = n4911 | n4242;
assign n7356 = ~n3250;
assign n7421 = n4360 | n8396;
assign n7925 = n2186 & n12453;
assign n10043 = ~(n63 ^ n11595);
assign n12681 = n3480 & n2611;
assign n12756 = n1107 & n5287;
assign n3288 = ~(n3136 ^ n8886);
assign n107 = n12119 | n12080;
assign n7146 = n10520 & n543;
assign n8775 = ~(n7929 ^ n5588);
assign n10523 = ~(n2934 | n2353);
assign n4870 = n420 | n10308;
assign n7763 = ~(n11593 ^ n4128);
assign n9484 = ~n12934;
assign n4419 = ~(n7034 | n10058);
assign n1079 = ~n10223;
assign n2910 = n1465 & n6272;
assign n12592 = ~(n10231 ^ n993);
assign n4257 = n1246 & n4355;
assign n10920 = n7383 & n4893;
assign n9068 = n5765 | n5759;
assign n11717 = n6365 | n6285;
assign n4655 = ~(n9684 ^ n6936);
assign n12437 = ~n3011;
assign n9880 = n12208 | n10017;
assign n12550 = n2456 | n12883;
assign n12116 = n3984 & n3902;
assign n8295 = n5915 | n1932;
assign n3468 = ~n8717;
assign n3890 = n6707 | n9870;
assign n8104 = ~(n7348 ^ n1806);
assign n8833 = ~(n2773 ^ n1718);
assign n12178 = n7391 | n1546;
assign n7871 = n3127 | n510;
assign n2483 = ~n3742;
assign n8716 = ~(n4804 | n9957);
assign n1725 = ~(n8903 ^ n5834);
assign n1403 = ~n4734;
assign n1800 = n8583 | n28;
assign n12378 = ~(n23 ^ n1830);
assign n5668 = ~(n3676 ^ n3173);
assign n12929 = ~n38;
assign n3664 = n11546 & n4638;
assign n32 = ~(n7559 ^ n4712);
assign n6010 = n1406 | n12168;
assign n2173 = ~(n445 ^ n9866);
assign n7836 = ~(n1111 ^ n7959);
assign n4987 = ~(n4976 | n5657);
assign n1704 = ~n8270;
assign n1149 = n11147 | n12290;
assign n10889 = ~(n9965 ^ n6803);
assign n4683 = ~(n21 ^ n3705);
assign n7963 = n9600 & n7860;
assign n6854 = n3837 & n9096;
assign n7807 = n6770 & n4634;
assign n10536 = ~(n8445 | n8754);
assign n1892 = ~(n12770 | n8877);
assign n3387 = ~(n3215 ^ n567);
assign n11707 = ~(n6942 ^ n10303);
assign n6569 = n7839 | n6455;
assign n11491 = n8153 & n10266;
assign n7574 = n3820 | n4642;
assign n8229 = n10750 | n8655;
assign n7583 = ~(n7764 | n6710);
assign n10947 = n4312 & n4634;
assign n3153 = n10750 | n4913;
assign n8626 = ~n12794;
assign n2541 = ~(n298 ^ n4919);
assign n10686 = ~(n12506 ^ n2489);
assign n1774 = ~(n9269 | n9169);
assign n2974 = ~n10993;
assign n5364 = n3617 | n3224;
assign n10053 = n3667 | n5580;
assign n6169 = ~n7354;
assign n4796 = n6470 & n7392;
assign n5898 = ~(n5869 ^ n7231);
assign n1363 = ~(n6895 ^ n414);
assign n9003 = n3818 | n10716;
assign n6920 = ~(n3268 ^ n1045);
assign n3023 = n91 | n3162;
assign n2847 = n630 | n12394;
assign n3859 = ~n8573;
assign n1505 = n10781 & n4941;
assign n8803 = ~n8477;
assign n10694 = ~(n8161 ^ n8218);
assign n1536 = ~(n10984 ^ n11643);
assign n5481 = ~(n3984 ^ n3902);
assign n3628 = n10835 | n9144;
assign n10712 = ~n8605;
assign n25 = ~n12201;
assign n1533 = n4479 | n859;
assign n3962 = ~n7309;
assign n231 = n10049 & n1521;
assign n12167 = n7283 | n4775;
assign n1715 = n11026 | n795;
assign n636 = ~n7891;
assign n6596 = ~n2296;
assign n10577 = ~(n5928 | n3511);
assign n9233 = ~n3255;
assign n12325 = ~(n4696 ^ n416);
assign n1815 = n9657 & n1807;
assign n7124 = ~n3202;
assign n124 = n10055 | n12613;
assign n10602 = n2979 & n4298;
assign n8475 = n752 | n7876;
assign n11726 = n9179 & n9479;
assign n10735 = n10142 | n1915;
assign n2559 = n4193 | n12637;
assign n9289 = n6797 & n5645;
assign n11434 = n2677 & n9579;
assign n12311 = ~(n8036 ^ n10094);
assign n10512 = n5305 & n2509;
assign n9167 = n11923 | n8830;
assign n3974 = n12775 | n12913;
assign n4182 = n5858 | n11827;
assign n2721 = n5575 | n12816;
assign n8676 = n4741 & n4384;
assign n4110 = n11597 & n9573;
assign n7727 = ~(n392 ^ n9940);
assign n5723 = ~(n9553 ^ n1771);
assign n232 = n5848 & n3913;
assign n3307 = ~(n10473 ^ n10167);
assign n2505 = n11013 | n1346;
assign n6232 = ~(n6053 ^ n2118);
assign n11837 = ~(n10562 ^ n8250);
assign n8239 = ~(n1363 ^ n6438);
assign n8512 = n1026 & n11169;
assign n2687 = n183 | n10638;
assign n11826 = n2832 | n11746;
assign n5669 = ~(n7029 ^ n9249);
assign n790 = ~n9038;
assign n5508 = ~(n6384 | n12233);
assign n6785 = ~n6148;
assign n12701 = n6373 | n4527;
assign n1108 = ~(n12668 ^ n10462);
assign n10027 = ~n1440;
assign n11233 = ~n7057;
assign n6099 = ~(n3659 ^ n11250);
assign n12376 = n8954 | n10870;
assign n1127 = ~(n4202 | n9496);
assign n10294 = ~n8868;
assign n12081 = n9106 & n1488;
assign n8086 = ~(n1024 ^ n7498);
assign n1 = n2346 | n6228;
assign n8465 = ~(n8181 ^ n8485);
assign n10503 = ~(n6534 ^ n10826);
assign n7179 = ~(n2089 ^ n2015);
assign n10416 = ~(n2199 ^ n10954);
assign n11572 = ~(n3921 | n3199);
assign n2924 = n8476 & n6016;
assign n9912 = ~(n5274 ^ n2418);
assign n10815 = ~(n4205 ^ n8931);
assign n4767 = n8117 & n745;
assign n9213 = ~(n2144 | n2392);
assign n4208 = ~(n2479 ^ n8144);
assign n12107 = n12186 | n12816;
assign n10516 = n6577 | n10919;
assign n427 = n4338 | n10237;
assign n11912 = ~(n10378 ^ n7279);
assign n8996 = n12119 | n3924;
assign n5809 = ~n10545;
assign n8738 = ~n3986;
assign n8810 = n5765 | n4875;
assign n5146 = n3328 & n10633;
assign n3358 = n10637 | n3057;
assign n9760 = ~(n8416 ^ n5562);
assign n12861 = ~(n7521 ^ n4244);
assign n7505 = n12312 & n7063;
assign n84 = ~(n6535 ^ n1482);
assign n10077 = ~n3772;
assign n1447 = n4301 & n2204;
assign n12708 = n5383 | n10553;
assign n3909 = n11401 | n2666;
assign n578 = n11539 & n7445;
assign n5976 = n10095 & n6546;
assign n11046 = ~(n6064 | n7069);
assign n8748 = n10365 | n10723;
assign n602 = n752 | n8414;
assign n2019 = n10162 & n1558;
assign n12189 = n12503 | n9568;
assign n8013 = ~(n4373 ^ n5628);
assign n11331 = n2473 | n7782;
assign n4652 = n3072 & n8111;
assign n29 = ~(n7490 ^ n10974);
assign n4443 = n8964 | n5839;
assign n6343 = ~(n3726 ^ n277);
assign n8902 = ~(n2962 | n6955);
assign n3625 = n3743 | n10916;
assign n11490 = n10835 | n11698;
assign n6104 = n2656 | n5536;
assign n5671 = ~n11178;
assign n648 = n11712 | n9574;
assign n2674 = ~(n6041 | n6923);
assign n1738 = ~n9637;
assign n4121 = n2456 | n5326;
assign n8793 = n3261 & n11673;
assign n7083 = ~(n5652 ^ n12768);
assign n720 = n5452 & n6117;
assign n3317 = ~(n11250 | n5379);
assign n705 = n2217 | n7506;
assign n5776 = ~(n8133 ^ n10317);
assign n3600 = n2001 & n8698;
assign n10343 = n5530 | n12754;
assign n2657 = n6186 | n4998;
assign n7709 = ~n9457;
assign n2418 = ~(n3314 ^ n915);
assign n4760 = n4366 | n10752;
assign n7355 = ~(n361 ^ n7728);
assign n2981 = n7283 | n561;
assign n12065 = n4498 | n1546;
assign n609 = ~n5153;
assign n6928 = ~n2141;
assign n9666 = ~(n2608 ^ n4615);
assign n1935 = n2893 & n1014;
assign n7835 = n4808 & n5388;
assign n9580 = ~(n7311 | n2344);
assign n2919 = n9058 & n4197;
assign n7203 = n6270 | n3877;
assign n11112 = n4059 | n4400;
assign n8051 = n1685 | n11030;
assign n6774 = n4674 | n3224;
assign n9416 = n4702 & n3750;
assign n296 = n12503 | n3606;
assign n8175 = n6373 | n9144;
assign n1170 = ~(n895 | n290);
assign n12194 = n7185 | n2895;
assign n10777 = n4628 | n10422;
assign n9225 = ~n7976;
assign n4495 = ~(n5650 ^ n11675);
assign n9707 = n8241 & n8962;
assign n1997 = ~n12163;
assign n11038 = n9920 & n3932;
assign n3886 = n8216 & n10480;
assign n12315 = n12163 & n8684;
assign n5265 = n9734 | n900;
assign n3141 = n8026 | n11820;
assign n1058 = ~n2918;
assign n459 = ~(n1495 ^ n1506);
assign n6540 = n3310 | n2706;
assign n2923 = n10434 | n9894;
assign n5210 = ~n7499;
assign n9904 = ~(n5690 ^ n1607);
assign n12565 = ~(n6356 | n9270);
assign n3044 = ~(n9398 ^ n446);
assign n1159 = ~(n2583 ^ n954);
assign n6643 = n8428 | n10919;
assign n4483 = n4628 | n8740;
assign n9262 = ~n4722;
assign n4861 = ~(n6283 ^ n5838);
assign n6242 = n8552 | n12735;
assign n550 = n8428 | n6084;
assign n920 = n2056 & n10008;
assign n4430 = ~(n9267 ^ n9044);
assign n12750 = n8070 | n473;
assign n8415 = n8920 & n8547;
assign n8323 = n936 | n5520;
assign n9300 = ~(n4852 ^ n7868);
assign n50 = n9389 | n4775;
assign n9137 = ~(n12081 ^ n153);
assign n6514 = n962 | n9144;
assign n10006 = ~(n4084 | n2120);
assign n2976 = n10142 | n1079;
assign n12063 = n2838 | n6164;
assign n11240 = ~(n9647 | n11633);
assign n10832 = n8458 | n3761;
assign n1635 = ~(n7275 | n3788);
assign n2718 = ~n1548;
assign n2047 = n5082 & n8365;
assign n11285 = n8959 | n6455;
assign n3425 = ~n8776;
assign n3889 = ~(n11507 | n3685);
assign n12121 = n6940 | n7615;
assign n6387 = ~(n12703 ^ n8033);
assign n3489 = ~n5078;
assign n5744 = n6377 & n12854;
assign n1572 = ~(n7824 | n12880);
assign n2338 = n8687 | n4654;
assign n4490 = n1839 & n4585;
assign n10015 = ~(n12556 ^ n997);
assign n4381 = ~n11189;
assign n8990 = ~(n820 ^ n12499);
assign n3866 = n3414 | n5170;
assign n218 = ~(n4112 ^ n2282);
assign n8209 = ~(n4766 | n9346);
assign n12412 = ~(n9081 ^ n3026);
assign n5050 = n10211 | n8355;
assign n3089 = ~(n2197 ^ n2281);
assign n694 = n2191 & n3550;
assign n1205 = n8959 | n2815;
assign n9274 = n10835 | n5914;
assign n8811 = ~(n11149 ^ n7385);
assign n12255 = ~(n12550 ^ n9946);
assign n10035 = n2639 | n6420;
assign n8817 = ~n5059;
assign n12544 = ~(n2271 | n2399);
assign n6867 = n6776 & n10439;
assign n2401 = n989 | n9589;
assign n2511 = n6740 | n9524;
assign n2852 = n12853 | n10422;
assign n4667 = n6570 | n11756;
assign n5867 = ~n11840;
assign n6451 = n8959 | n5540;
assign n3116 = n5530 | n7136;
assign n538 = ~(n5386 ^ n12572);
assign n1868 = n12423 & n7303;
assign n8756 = ~n8784;
assign n2116 = n8959 | n7425;
assign n3441 = n3746 | n6084;
assign n8331 = ~(n7 ^ n4663);
assign n4783 = n3242 & n6957;
assign n2889 = ~(n8551 ^ n12230);
assign n12439 = ~n10841;
assign n11360 = ~(n12040 ^ n11349);
assign n717 = n9077 & n5332;
assign n11692 = ~(n758 | n2826);
assign n882 = n3617 | n12535;
assign n3874 = n11653 | n4524;
assign n10031 = ~(n6037 ^ n5347);
assign n8758 = n5355 | n9589;
assign n9516 = ~(n7602 ^ n1841);
assign n3008 = ~(n7115 ^ n2330);
assign n11506 = ~(n11460 | n12888);
assign n11962 = n8220 | n7838;
assign n12222 = ~(n3579 ^ n8300);
assign n5163 = ~(n11013 ^ n2022);
assign n3500 = ~(n8149 ^ n109);
assign n6027 = n660 | n2927;
assign n7856 = ~n953;
assign n7918 = ~(n9606 | n679);
assign n9131 = ~(n666 ^ n10519);
assign n4492 = n7854 & n4952;
assign n596 = ~(n5881 | n10150);
assign n8556 = n2393 & n7294;
assign n12478 = ~n2476;
assign n5176 = ~(n5660 ^ n6107);
assign n1221 = ~(n5898 ^ n3139);
assign n702 = ~(n8458 ^ n3761);
assign n6796 = n5369 | n4259;
assign n7299 = ~(n1864 ^ n10145);
assign n5171 = ~(n3910 | n6548);
assign n11308 = ~(n8914 ^ n11802);
assign n1705 = n5355 | n7424;
assign n1426 = n1848 & n1374;
assign n3372 = ~(n5635 ^ n4056);
assign n10723 = ~(n10448 ^ n6747);
assign n10668 = n6681 & n10894;
assign n10933 = n7765 & n4208;
assign n1751 = ~(n2459 ^ n4594);
assign n7499 = n9389 | n2358;
assign n6988 = n5283 & n7610;
assign n12229 = ~n12241;
assign n8871 = n8429 | n10376;
assign n5404 = n8187 | n7881;
assign n9957 = ~(n11659 | n11408);
assign n11605 = n5765 | n6922;
assign n12211 = ~n7850;
assign n8330 = ~n10689;
assign n9120 = n9702 | n4844;
assign n5352 = ~(n12539 ^ n10409);
assign n9325 = n2133 | n11530;
assign n767 = ~n9882;
assign n2653 = ~n10686;
assign n10840 = n8870 | n5468;
assign n9279 = ~n7668;
assign n5518 = ~n721;
assign n1476 = ~n6611;
assign n7903 = n5366 | n5004;
assign n8640 = n5108 ^ n8939;
assign n7111 = n6373 | n4654;
assign n4324 = n6098 | n1845;
assign n11613 = n3820 | n1047;
assign n8207 = n9687 & n11344;
assign n5443 = ~(n7012 ^ n3834);
assign n6510 = ~n7929;
assign n9239 = n7268 | n1767;
assign n10942 = ~n10214;
assign n282 = n9389 | n6389;
assign n4207 = ~n11323;
assign n1977 = ~(n10834 ^ n6624);
assign n8562 = ~(n9404 ^ n9679);
assign n8655 = ~n4826;
assign n10484 = ~(n7284 ^ n365);
assign n10881 = n11998 | n11648;
assign n2888 = ~(n4023 ^ n7696);
assign n6073 = n10142 | n4242;
assign n5657 = ~(n8117 | n745);
assign n5906 = ~(n9627 ^ n833);
assign n5525 = n7391 | n3911;
assign n11199 = ~n7370;
assign n11776 = ~(n11754 ^ n3814);
assign n7890 = n10531 & n1467;
assign n4995 = n10065 | n198;
assign n9788 = ~(n7666 ^ n11010);
assign n10576 = n5495 | n10986;
assign n11640 = ~(n12500 ^ n2829);
assign n10623 = ~n5408;
assign n11693 = ~(n5059 ^ n4099);
assign n2390 = n1064 | n4813;
assign n1030 = ~(n3381 ^ n10811);
assign n5470 = ~(n120 | n65);
assign n487 = ~(n12939 | n6858);
assign n443 = n6368 | n1309;
assign n6721 = ~(n7680 | n8662);
assign n12003 = ~(n822 ^ n7162);
assign n8905 = n12237 | n12735;
assign n11500 = n2997 & n6848;
assign n8145 = n9373 | n7506;
assign n7735 = n5331 & n1512;
assign n6218 = n8011 | n4866;
assign n9843 = n8310 | n2912;
assign n3155 = n357 | n5306;
assign n395 = ~(n7635 ^ n10300);
assign n1799 = ~n4914;
assign n1182 = n62 | n377;
assign n12673 = n5361 | n6282;
assign n12137 = ~(n10514 | n11187);
assign n12434 = ~(n4779 | n4890);
assign n7122 = ~(n7622 ^ n10067);
assign n4253 = ~(n7675 ^ n6828);
assign n2941 = n3962 & n4463;
assign n780 = ~(n5707 ^ n9944);
assign n6161 = n989 | n2076;
assign n3827 = ~(n6882 ^ n6622);
assign n10055 = ~n6773;
assign n11870 = ~(n6660 ^ n7096);
assign n3402 = ~(n2443 | n3859);
assign n142 = n5621 & n4075;
assign n6413 = n12133 & n6866;
assign n4256 = n5893 & n6088;
assign n5565 = ~(n1046 ^ n3683);
assign n919 = ~n11336;
assign n5278 = n5527 & n1217;
assign n11518 = n8273 | n4909;
assign n526 = ~n4292;
assign n9570 = n989 | n1915;
assign n261 = ~n8035;
assign n7531 = ~(n7614 ^ n471);
assign n8674 = n10157 | n10916;
assign n2500 = n4870 & n500;
assign n5030 = ~(n4323 ^ n7426);
assign n11187 = n2520 & n1745;
assign n10235 = ~(n8596 | n3584);
assign n3086 = ~(n720 ^ n12516);
assign n2343 = ~(n11396 ^ n4847);
assign n6630 = ~n6059;
assign n11789 = ~(n1461 ^ n7491);
assign n2865 = ~(n5715 | n7720);
assign n2607 = n1469 | n10489;
assign n4777 = n3743 | n5258;
assign n8112 = n966 | n11943;
assign n5982 = n8870 | n826;
assign n54 = n12361 | n6084;
assign n12898 = ~(n4511 | n8863);
assign n11224 = ~(n8267 ^ n11939);
assign n6991 = ~n12215;
assign n11370 = n989 | n3911;
assign n12858 = n3743 | n609;
assign n9115 = ~(n4289 ^ n3035);
assign n9941 = ~(n601 ^ n3269);
assign n1884 = ~(n577 ^ n8482);
assign n12560 = n4263 & n8131;
assign n9539 = ~(n8293 ^ n12519);
assign n7996 = n962 | n4654;
assign n6029 = n12443 & n1734;
assign n7564 = n10142 | n12328;
assign n7186 = ~n3313;
assign n5082 = n173 & n3686;
assign n1034 = ~(n10031 ^ n5467);
assign n5532 = n8687 | n2020;
assign n12235 = ~n3991;
assign n2282 = n11923 | n12771;
assign n8848 = n10196 | n2020;
assign n12913 = n4911 | n10066;
assign n10517 = n11311 & n2522;
assign n530 = ~n4970;
assign n3432 = ~(n2033 ^ n8014);
assign n3593 = n7358 & n466;
assign n4542 = ~(n4298 ^ n1001);
assign n2722 = n12423 | n7303;
assign n6243 = n1415 & n4630;
assign n7138 = ~n6121;
assign n1346 = ~(n4449 ^ n4391);
assign n6860 = ~(n12693 ^ n10616);
assign n5172 = n3533 & n5660;
assign n8031 = ~n4417;
assign n1697 = n5855 & n3487;
assign n3474 = n114 | n7876;
assign n4267 = ~n3807;
assign n3487 = n11051 | n9731;
assign n2524 = n3611 | n11027;
assign n7242 = ~(n3305 ^ n6890);
assign n8399 = ~(n10873 ^ n1950);
assign n6509 = n8480 | n5865;
assign n11565 = ~(n4442 ^ n11248);
assign n1157 = n1941 | n6455;
assign n10878 = n5363 & n3006;
assign n8605 = ~(n10814 ^ n7368);
assign n8423 = n11958 | n6197;
assign n4045 = n8557 & n7653;
assign n3641 = ~(n2061 ^ n1158);
assign n2855 = ~(n4755 ^ n11338);
assign n8615 = ~n9737;
assign n10464 = ~n9326;
assign n6653 = ~(n7480 ^ n1080);
assign n8044 = ~(n12526 ^ n5750);
assign n2858 = n6298 | n6721;
assign n10872 = n6077 & n11715;
assign n6111 = n3106 & n11945;
assign n2803 = ~(n2284 ^ n11102);
assign n7220 = ~(n4431 | n6243);
assign n11026 = ~n2393;
assign n2961 = ~(n5204 ^ n283);
assign n9804 = ~(n11782 ^ n5114);
assign n12218 = ~n12747;
assign n7558 = ~n2522;
assign n11425 = n2217 | n5258;
assign n4614 = ~(n8503 | n3889);
assign n5733 = ~(n10452 ^ n10676);
assign n11192 = n962 | n9160;
assign n9133 = ~(n11945 ^ n6487);
assign n8714 = ~n4603;
assign n2931 = ~n7490;
assign n7693 = ~(n129 ^ n9330);
assign n9702 = n2195 & n1101;
assign n6525 = ~(n391 | n1821);
assign n10914 = ~(n1644 ^ n11612);
assign n9183 = ~(n5503 | n730);
assign n7970 = ~n9727;
assign n679 = ~n7647;
assign n8333 = ~(n4866 ^ n8252);
assign n7739 = ~n11575;
assign n4880 = ~(n12305 ^ n3223);
assign n3700 = n1872 | n3556;
assign n11352 = n5575 | n7876;
assign n6235 = n4053 | n10130;
assign n1578 = ~(n1879 | n142);
assign n358 = n8959 | n2232;
assign n7090 = ~n12790;
assign n2625 = n10157 | n609;
assign n1032 = ~(n4690 ^ n8965);
assign n3163 = n7432 & n5058;
assign n11300 = ~(n9557 ^ n4574);
assign n3692 = n11475 & n7800;
assign n3463 = ~(n737 | n6132);
assign n7734 = n1172 & n3669;
assign n3818 = ~n9508;
assign n8360 = ~(n11588 ^ n9112);
assign n5389 = ~n1062;
assign n9050 = n11542 & n6333;
assign n7755 = ~n8533;
assign n5010 = n10594 & n6540;
assign n1158 = ~(n7297 ^ n7935);
assign n6224 = n10108 | n12843;
assign n12659 = n3743 | n5502;
assign n8215 = n11753 | n3341;
assign n2204 = n11719 | n11827;
assign n7321 = n8430 & n1452;
assign n1148 = ~n8460;
assign n7967 = n12023 | n7734;
assign n3857 = ~(n2881 | n7744);
assign n4799 = n6437 & n12847;
assign n5587 = ~(n1355 ^ n7273);
assign n5944 = n6718 | n4864;
assign n345 = ~(n6931 ^ n1197);
assign n9058 = n2427 | n1157;
assign n9248 = n7586 | n1505;
assign n211 = ~n3536;
assign n11414 = ~(n1784 ^ n11686);
assign n3611 = ~(n7856 ^ n2798);
assign n1393 = n7381 | n865;
assign n12806 = ~(n320 ^ n12447);
assign n7917 = ~(n11360 ^ n2803);
assign n1338 = n2101 & n3422;
assign n11056 = ~(n5269 | n12488);
assign n1066 = n8450 | n10025;
assign n1843 = ~n7652;
assign n5445 = n664 & n9991;
assign n6312 = n1699 | n4913;
assign n9884 = n994 | n7703;
assign n3145 = n5575 | n995;
assign n126 = ~n5789;
assign n3139 = ~(n849 ^ n329);
assign n12908 = ~(n3265 ^ n1454);
assign n11592 = n5393 | n6733;
assign n8609 = ~(n10516 ^ n778);
assign n5485 = n11026 | n4527;
assign n11264 = ~(n2673 ^ n2648);
assign n8278 = ~(n9616 ^ n5262);
assign n6030 = n3544 | n4715;
assign n6852 = ~n7419;
assign n12318 = n5575 | n184;
assign n5619 = n6171 | n7351;
assign n9654 = ~(n3921 ^ n429);
assign n4344 = ~(n2503 ^ n5908);
assign n2264 = ~(n8023 ^ n9300);
assign n11761 = ~(n2162 | n7307);
assign n2079 = ~n11633;
assign n4882 = n4791 & n5762;
assign n2386 = ~n10923;
assign n3130 = n3820 | n4654;
assign n147 = n12648 & n2802;
assign n7700 = ~(n10958 ^ n540);
assign n6982 = n12144 & n5251;
assign n5290 = ~(n2309 | n3798);
assign n7621 = ~(n10992 ^ n14);
assign n9840 = ~(n248 ^ n11837);
assign n6200 = ~n10457;
assign n1160 = ~n822;
assign n5705 = ~(n9481 ^ n12507);
assign n63 = ~(n12095 | n1578);
assign n6428 = ~(n5989 ^ n3457);
assign n3674 = ~n10877;
assign n11762 = n7329 | n8461;
assign n9016 = n12119 | n8109;
assign n606 = ~(n6121 ^ n2158);
assign n1420 = ~(n7278 ^ n598);
assign n8611 = ~n12628;
assign n1374 = n8019 | n9631;
assign n12497 = n209 | n4050;
assign n3773 = n10309 & n11180;
assign n9504 = n5530 | n8655;
assign n7960 = n810 & n2058;
assign n4983 = ~n7612;
assign n2966 = n11892 & n806;
assign n1178 = n4097 & n11394;
assign n9830 = n6478 & n3855;
assign n4112 = n5765 | n9568;
assign n10091 = n7116 | n11820;
assign n1905 = ~(n2858 ^ n5772);
assign n1277 = ~n2784;
assign n10861 = ~(n12715 ^ n11494);
assign n9751 = ~n5688;
assign n5502 = ~n159;
assign n257 = n11594 | n272;
assign n10688 = n5700 | n2958;
assign n2412 = ~n628;
assign n614 = n573 | n11044;
assign n10802 = n5479 & n8519;
assign n1860 = ~(n8070 ^ n473);
assign n6767 = ~(n8774 ^ n3152);
assign n6705 = ~(n10407 ^ n2755);
assign n10864 = ~(n11734 | n6862);
assign n11251 = ~n9007;
assign n12279 = ~(n5361 ^ n12729);
assign n5507 = ~n904;
assign n5658 = n10157 | n9160;
assign n1039 = n1518 & n211;
assign n5718 = n7391 | n6389;
assign n11279 = ~(n12782 ^ n2379);
assign n1707 = ~(n6536 ^ n6532);
assign n2999 = n255 & n4288;
assign n1123 = n752 | n9971;
assign n9256 = n3348 | n67;
assign n8881 = n5620 | n9864;
assign n11032 = ~(n2574 | n1190);
assign n4545 = n4214 & n7650;
assign n7879 = n8452 & n8978;
assign n4448 = ~n3914;
assign n962 = ~n1471;
assign n4454 = ~(n5856 ^ n10890);
assign n2288 = n4112 | n2282;
assign n11134 = ~(n5554 ^ n12161);
assign n4873 = ~n12939;
assign n9299 = n3160 | n1116;
assign n5090 = ~(n8103 ^ n5741);
assign n2601 = ~(n3235 | n407);
assign n6214 = n11413 | n937;
assign n1037 = ~(n6987 ^ n3200);
assign n6521 = n5195 & n4478;
assign n4766 = ~n10117;
assign n4331 = n9185 & n3250;
assign n1036 = n8453 & n4625;
assign n343 = ~(n11119 ^ n7274);
assign n942 = n1947 & n11587;
assign n7245 = n11073 & n5965;
assign n11323 = ~(n10096 ^ n4208);
assign n2100 = n9878 | n4913;
assign n7604 = n6854 | n2439;
assign n10050 = n612 | n9775;
assign n10521 = n10242 & n12660;
assign n6937 = ~(n1483 ^ n5676);
assign n1131 = n2456 | n7928;
assign n800 = n3361 | n1243;
assign n6610 = ~(n12739 ^ n6652);
assign n11823 = ~n4435;
assign n12018 = ~(n9899 | n3737);
assign n9127 = ~(n10738 ^ n6451);
assign n3686 = ~n11498;
assign n10817 = n12622 & n3919;
assign n9744 = n191 | n8859;
assign n5567 = ~n2376;
assign n12147 = ~n10918;
assign n2190 = n6977 | n6084;
assign n2823 = ~n1210;
assign n4374 = ~(n6557 ^ n11804);
assign n7793 = ~(n8872 ^ n11270);
assign n2025 = ~(n3372 | n6124);
assign n2929 = ~(n3633 ^ n3825);
assign n5289 = n9448 | n4181;
assign n9848 = ~(n11727 ^ n1119);
assign n7055 = ~(n9342 | n11970);
assign n5477 = n5252 | n3309;
assign n10750 = ~n12391;
assign n68 = ~(n7016 ^ n11437);
assign n11845 = ~(n656 | n10580);
assign n5478 = ~(n5243 ^ n11640);
assign n7511 = n8549 & n2493;
assign n11743 = n9054 | n10082;
assign n9855 = ~(n2859 ^ n2949);
assign n11689 = n9370 | n5497;
assign n4375 = n2254 & n10227;
assign n7211 = ~(n4759 ^ n929);
assign n9871 = n11923 | n9280;
assign n1973 = n11958 | n2232;
assign n3377 = n591 | n11790;
assign n6315 = ~(n95 ^ n5882);
assign n6809 = ~(n6700 ^ n6120);
assign n3779 = ~(n6212 ^ n10328);
assign n1362 = n12721 & n6196;
assign n12931 = ~(n8294 | n6316);
assign n6897 = n3628 & n894;
assign n12430 = ~(n4613 | n4098);
assign n10468 = ~n9608;
assign n2942 = ~(n8816 ^ n1217);
assign n5189 = n8928 ^ n2974;
assign n3544 = n11958 | n3421;
assign n11486 = ~(n9161 | n2531);
assign n6665 = n3998 & n608;
assign n1211 = ~(n2598 ^ n265);
assign n3329 = ~(n6782 | n7054);
assign n567 = ~(n3141 ^ n4721);
assign n10232 = ~(n6738 ^ n252);
assign n4458 = n12853 | n6513;
assign n3385 = ~(n5621 ^ n1879);
assign n4700 = n2923 & n7999;
assign n8641 = n1642 | n12325;
assign n2958 = ~(n5863 ^ n3149);
assign n11477 = n12758 & n7584;
assign n7811 = ~(n6750 ^ n3701);
assign n5727 = ~n3815;
assign n7443 = ~n6364;
assign n7052 = n9007 | n7956;
assign n8140 = n9105 & n1981;
assign n12573 = n7128 & n6684;
assign n4359 = ~(n12117 | n143);
assign n274 = n9453 & n9646;
assign n5180 = n7694 & n12015;
assign n4460 = n1699 | n12535;
assign n3108 = n807 | n6455;
assign n7366 = ~(n10619 ^ n11819);
assign n9833 = n3105 & n358;
assign n5699 = ~n7997;
assign n239 = ~n8864;
assign n6488 = ~(n5080 ^ n7917);
assign n6912 = ~(n11677 ^ n1025);
assign n697 = n8552 | n9188;
assign n2107 = ~n1113;
assign n8221 = n12853 | n1932;
assign n8970 = ~n11536;
assign n344 = n204 & n6608;
assign n4428 = n3110 & n4940;
assign n3211 = n10791 & n8508;
assign n4602 = n8858 & n4452;
assign n347 = n5685 | n5658;
assign n3513 = n5950 & n5359;
assign n10248 = ~n4181;
assign n1486 = ~n3326;
assign n9066 = n7468 | n271;
assign n10093 = ~(n6085 | n12029);
assign n2933 = n9878 | n826;
assign n4175 = n1024 & n7498;
assign n1482 = ~(n7621 ^ n8614);
assign n5937 = ~n11136;
assign n12780 = n1089 & n10310;
assign n4016 = n6637 | n461;
assign n11673 = n6739 | n9109;
assign n10846 = n7283 | n1851;
assign n2622 = ~(n9290 ^ n6049);
assign n2437 = ~n6539;
assign n8410 = n8702 | n8911;
assign n2357 = n2176 & n8516;
assign n1416 = n5158 & n7751;
assign n6122 = n6577 | n6084;
assign n5563 = ~(n6447 ^ n11891);
assign n7927 = n5671 | n1134;
assign n10607 = ~n8445;
assign n9180 = n3611 & n11027;
assign n9285 = n10148 & n7996;
assign n4649 = ~(n7493 | n8551);
assign n10069 = ~(n6470 ^ n7392);
assign n5221 = ~(n4981 ^ n12209);
assign n1334 = n4059 | n510;
assign n4843 = ~n11388;
assign n10130 = n8996 & n9518;
assign n5825 = ~(n12545 ^ n1180);
assign n9008 = ~(n10225 | n3598);
assign n10422 = ~n2551;
assign n10213 = ~(n11205 ^ n11622);
assign n8094 = n6439 | n6447;
assign n3530 = ~n3170;
assign n9371 = ~(n7380 ^ n11427);
assign n1668 = n3740 | n10116;
assign n9951 = ~(n8879 | n7199);
assign n7647 = n5330 & n1401;
assign n3941 = n11709 & n831;
assign n3926 = n11181 | n4268;
assign n9503 = ~(n10598 | n2601);
assign n11239 = n1409 & n12780;
assign n5557 = ~(n1629 ^ n5509);
assign n98 = ~(n7910 ^ n8706);
assign n6674 = ~n4746;
assign n6952 = n10142 | n6524;
assign n8781 = ~(n1341 | n9522);
assign n2194 = ~(n7433 | n1884);
assign n4424 = n6718 | n9280;
assign n9247 = ~n10742;
assign n9558 = ~(n12723 ^ n1584);
assign n11674 = n7449 | n4875;
assign n803 = ~(n3925 | n4797);
assign n10158 = ~(n11844 | n6991);
assign n11577 = n8276 & n2024;
assign n5927 = ~(n12227 ^ n11940);
assign n1950 = ~(n1530 ^ n1115);
assign n337 = n4628 | n7382;
assign n8335 = n12579 & n6506;
assign n9993 = n7231 & n6505;
assign n11935 = n11923 | n7506;
assign n9069 = ~(n9848 ^ n2568);
assign n2520 = n2730 | n3094;
assign n2490 = n4343 | n9188;
assign n5155 = ~(n7318 ^ n8993);
assign n1525 = n9369 & n2952;
assign n12734 = n6577 | n7558;
assign n2660 = n6181 | n10334;
assign n744 = ~(n9353 ^ n9243);
assign n11098 = n961 & n9553;
assign n7019 = n6373 | n5502;
assign n1772 = ~(n9735 | n12481);
assign n325 = n10196 | n4527;
assign n8764 = n9277 | n9473;
assign n11075 = ~(n11783 ^ n2);
assign n9811 = ~(n7393 ^ n11507);
assign n1925 = ~(n10169 ^ n2473);
assign n9333 = ~n6507;
assign n12179 = n885 & n5836;
assign n618 = ~(n5773 | n12664);
assign n5992 = ~(n8417 ^ n9857);
assign n7771 = n12150 | n538;
assign n12664 = n10763 & n11582;
assign n4813 = n2516 & n11559;
assign n8746 = ~n4919;
assign n8314 = ~(n675 ^ n2290);
assign n1653 = n2217 | n1047;
assign n2496 = n2252 | n8340;
assign n11111 = ~n10702;
assign n2901 = n515 | n5941;
assign n8517 = ~(n2605 ^ n11921);
assign n317 = n5355 | n8970;
assign n5244 = ~(n7054 ^ n1040);
assign n210 = ~(n8294 ^ n7317);
assign n11749 = n7512 | n12181;
assign n12534 = ~(n302 ^ n12214);
assign n11560 = n7299 & n2239;
assign n8338 = n4029 & n8834;
assign n11643 = ~(n11212 ^ n12002);
assign n8069 = n12825 & n8744;
assign n3192 = n404 & n429;
assign n10056 = n807 | n6169;
assign n12356 = ~n8823;
assign n690 = n7947 & n493;
assign n1078 = ~n9347;
assign n7051 = n6602 | n2951;
assign n1991 = ~(n10254 ^ n8833);
assign n4236 = ~(n3330 ^ n7693);
assign n2983 = n5915 | n6071;
assign n10927 = ~(n9456 ^ n3101);
assign n2466 = n1409 | n12780;
assign n5238 = ~(n8380 | n1786);
assign n1506 = n686 | n995;
assign n8220 = n1249 & n7963;
assign n2777 = ~(n4007 ^ n7095);
assign n1678 = n4643 | n8913;
assign n5679 = n2217 | n9568;
assign n7959 = n10157 | n28;
assign n8146 = ~(n8741 ^ n2942);
assign n2838 = n5575 | n5538;
assign n4293 = ~(n11317 ^ n916);
assign n4321 = n10347 & n12182;
assign n10414 = n7449 | n12120;
assign n11348 = ~(n532 ^ n480);
assign n410 = ~n1218;
assign n9399 = ~n8529;
assign n5207 = n994 | n3911;
assign n9849 = n1941 | n3903;
assign n6035 = ~(n9141 ^ n901);
assign n3226 = n586 & n6172;
assign n1417 = ~(n372 | n1060);
assign n12678 = n12471 & n6433;
assign n8087 = ~(n3044 ^ n7066);
assign n7420 = ~n478;
assign n12490 = ~(n2277 ^ n4865);
assign n2358 = ~n4634;
assign n8858 = ~n5157;
assign n8702 = n5008 | n6841;
assign n5035 = ~(n8085 ^ n11814);
assign n9411 = n12870 & n10107;
assign n10106 = ~(n3105 ^ n358);
assign n8733 = ~n6483;
assign n2904 = n3457 | n3786;
assign n4184 = n4457 | n622;
assign n1659 = n4001 & n592;
assign n10613 = n2217 | n1739;
assign n3473 = ~(n7373 | n1340);
assign n7875 = ~n12653;
assign n1916 = ~(n8992 ^ n5106);
assign n5497 = ~n5212;
assign n6648 = ~n6599;
assign n1636 = ~n4406;
assign n10772 = n722 | n3987;
assign n3183 = ~(n5208 | n4917);
assign n3887 = n7462 | n2105;
assign n1519 = ~n8449;
assign n12208 = n2456 | n1163;
assign n3007 = n3127 | n7341;
assign n8760 = n11293 & n6013;
assign n8218 = ~(n5288 | n3040);
assign n115 = ~n9512;
assign n5271 = ~(n331 | n11840);
assign n12389 = ~(n11798 ^ n11143);
assign n10793 = n10325 | n10127;
assign n5248 = n3906 & n11203;
assign n2819 = ~(n9551 | n4044);
assign n582 = n10750 | n12080;
assign n7935 = ~(n9559 ^ n5050);
assign n3953 = n1097 & n7456;
assign n12754 = ~n447;
assign n10342 = n11812 & n6879;
assign n5267 = ~(n135 | n11786);
assign n4095 = ~(n3045 ^ n8558);
assign n10549 = ~(n10551 ^ n7988);
assign n145 = ~(n9519 ^ n1648);
assign n10645 = n2455 | n2567;
assign n2700 = n8959 | n7952;
assign n1881 = ~n6415;
assign n1041 = n10277 | n6343;
assign n4690 = ~(n11113 ^ n1005);
assign n7131 = n686 | n6455;
assign n7569 = ~(n5437 ^ n7104);
assign n7548 = ~(n8757 ^ n5031);
assign n9897 = ~(n10948 | n4359);
assign n10612 = ~(n11050 ^ n1336);
assign n8877 = ~(n7091 | n5427);
assign n8888 = ~(n6880 ^ n12440);
assign n11141 = n2515 & n12489;
assign n11326 = n3722 ^ n11793;
assign n3403 = ~(n10590 ^ n7821);
assign n2089 = n692 & n8763;
assign n3649 = ~(n4956 ^ n10521);
assign n3934 = ~(n12470 ^ n4336);
assign n6558 = ~(n7791 ^ n1227);
assign n7003 = ~(n3335 | n5740);
assign n3961 = n240 | n983;
assign n11827 = ~n7265;
assign n4670 = ~n438;
assign n513 = ~(n5130 ^ n9831);
assign n1936 = ~n7469;
assign n1886 = n9050 | n2873;
assign n6511 = ~(n9797 ^ n2900);
assign n5810 = n1012 & n11537;
assign n3440 = n1543 & n1600;
assign n2103 = n1752 | n2688;
assign n7898 = ~(n11683 ^ n7110);
assign n12002 = n5915 | n12754;
assign n10943 = n7625 | n2709;
assign n11338 = n8405 | n6513;
assign n2917 = n6977 | n6455;
assign n5000 = ~(n1135 ^ n9409);
assign n8984 = n12611 | n1437;
assign n4060 = ~(n9806 | n8579);
assign n1526 = ~n5475;
assign n5882 = n6979 & n6404;
assign n6089 = ~(n7301 ^ n3237);
assign n7534 = ~n9647;
assign n9857 = ~(n5179 ^ n529);
assign n10410 = n8596 & n3584;
assign n8205 = n10750 | n5781;
assign n11752 = ~n5167;
assign n5038 = ~(n7869 ^ n12455);
assign n4962 = ~(n11690 ^ n1914);
assign n2798 = ~n10528;
assign n12526 = n6577 | n3421;
assign n7870 = ~(n11174 | n2863);
assign n9093 = n4415 | n325;
assign n8288 = ~(n12879 | n7792);
assign n7058 = n9107 | n2986;
assign n11919 = ~(n7081 ^ n1713);
assign n11014 = n636 | n5468;
assign n10794 = n9531 | n1436;
assign n2279 = ~(n4235 | n7828);
assign n4073 = ~n1821;
assign n2377 = n4167 & n6892;
assign n4120 = ~(n9733 ^ n10564);
assign n6331 = ~n1361;
assign n7418 = ~(n2146 ^ n2636);
assign n9838 = n4187 & n2024;
assign n10630 = ~(n1626 ^ n1376);
assign n7380 = n6718 | n4527;
assign n135 = n10831 & n10959;
assign n5493 = n428 & n244;
assign n3978 = n10727 & n5662;
assign n12624 = n1335 | n1440;
assign n6698 = n7138 | n935;
assign n1115 = n8263 | n4545;
assign n2761 = n2034 & n2851;
assign n10369 = ~n2966;
assign n5252 = n8641 & n3890;
assign n6728 = ~(n12831 ^ n2915);
assign n1367 = ~n1804;
assign n5160 = n9884 & n3411;
assign n4567 = ~(n10963 ^ n465);
assign n11716 = ~n6159;
assign n9179 = n5809 | n1932;
assign n2548 = n5856 & n10890;
assign n7069 = ~(n8555 | n11568);
assign n9037 = n4272 & n11833;
assign n9079 = n752 | n995;
assign n12940 = n10607 | n341;
assign n8708 = ~(n7005 | n1291);
assign n1875 = ~(n6903 | n8419);
assign n2448 = n5530 | n10422;
assign n5391 = n6373 | n2020;
assign n10125 = ~(n11834 ^ n6459);
assign n3801 = n3078 & n6895;
assign n1402 = n11984 | n6460;
assign n10571 = ~(n4217 | n11726);
assign n298 = ~(n9827 ^ n12893);
assign n1110 = ~(n3354 ^ n8604);
assign n9025 = ~(n7911 ^ n6753);
assign n11019 = n808 & n9934;
assign n4039 = ~(n6291 | n5035);
assign n2826 = n7745 & n11854;
assign n1074 = n9881 & n9474;
assign n3655 = n9437 & n7908;
assign n9282 = ~(n504 | n3873);
assign n8334 = ~n8159;
assign n12329 = n5915 | n8109;
assign n2517 = ~(n6133 ^ n9913);
assign n12197 = n4358 | n10165;
assign n10877 = n752 | n2815;
assign n3835 = ~(n12476 | n485);
assign n2678 = ~n7790;
assign n3156 = n7009 | n4534;
assign n8529 = n7236 & n9763;
assign n11195 = n2124 | n3553;
assign n12643 = n4859 | n2263;
assign n7154 = n8187 | n7424;
assign n301 = n7232 | n1013;
assign n1966 = n10104 & n10498;
assign n11333 = ~(n3876 ^ n10111);
assign n4229 = ~n3017;
assign n196 = n4628 | n12735;
assign n6856 = ~(n5107 ^ n258);
assign n9221 = ~(n1816 | n5037);
assign n10463 = n3622 | n7803;
assign n6722 = ~(n5099 ^ n570);
assign n5342 = n5902 | n10066;
assign n6002 = n6776 & n10451;
assign n4464 = n7391 | n12843;
assign n10797 = ~n1131;
assign n527 = n5655 | n2296;
assign n11458 = ~(n5394 ^ n5152);
assign n2053 = n9914 | n1573;
assign n9755 = ~(n843 | n717);
assign n7966 = ~(n5615 ^ n5717);
assign n7302 = n6374 & n5757;
assign n11623 = n3691 | n4315;
assign n8879 = ~(n3464 | n8805);
assign n1459 = n3571 & n4869;
assign n2743 = n11846 | n7117;
assign n4888 = n636 | n8644;
assign n12191 = ~n9590;
assign n7447 = ~n5206;
assign n2287 = n7663 | n11886;
assign n8957 = ~n10685;
assign n4354 = ~(n1160 | n7162);
assign n12333 = n9170 | n7703;
assign n725 = n4327 | n8059;
assign n295 = n1303 & n4754;
assign n12188 = n6286 | n424;
assign n6902 = n5562 | n4550;
assign n3175 = ~n5039;
assign n4004 = n8977 & n5040;
assign n12201 = ~(n7519 ^ n9371);
assign n7955 = n3038 | n11124;
assign n11679 = n5530 | n8109;
assign n8947 = n9685 & n1926;
assign n12237 = ~n4828;
assign n12317 = n1883 | n105;
assign n1162 = ~n2509;
assign n8537 = ~(n9440 ^ n7068);
assign n4787 = n10750 | n1163;
assign n9867 = ~(n7100 ^ n9714);
assign n208 = ~(n10399 ^ n1426);
assign n11095 = n4549 & n8215;
assign n4904 = ~(n1131 ^ n11159);
assign n8927 = ~(n8171 ^ n11111);
assign n4521 = n9784 & n6920;
assign n5108 = ~(n12405 ^ n3415);
assign n11396 = n4911 | n3911;
assign n4275 = n1333 & n9195;
assign n11262 = ~n12541;
assign n861 = ~(n51 ^ n3764);
assign n3894 = ~(n6591 ^ n10653);
assign n99 = ~(n4658 | n2723);
assign n12808 = n7620 & n1724;
assign n9107 = n2099 | n5326;
assign n10430 = ~(n10135 ^ n4632);
assign n2990 = n2848 & n3695;
assign n6813 = ~(n5500 ^ n393);
assign n10209 = ~(n10556 ^ n7390);
assign n4673 = ~(n1807 ^ n6477);
assign n9624 = n2544 | n9477;
assign n9550 = n12026 & n6104;
assign n8024 = n10135 & n9854;
assign n1244 = ~(n2097 ^ n8794);
assign n8318 = n6819 | n3191;
assign n8709 = ~(n284 ^ n5010);
assign n8038 = n4403 | n8198;
assign n11779 = n9632 & n9210;
assign n3789 = ~(n5189 | n7960);
assign n9999 = ~(n9729 ^ n1690);
assign n1119 = n7839 | n5540;
assign n11214 = n2774 | n1617;
assign n10620 = n5328 | n7647;
assign n7330 = n9352 & n11275;
assign n6907 = ~(n10592 ^ n216);
assign n9893 = ~(n1672 | n8513);
assign n8117 = n3833 & n11418;
assign n9791 = ~(n6086 ^ n2356);
assign n6842 = ~(n10387 ^ n3019);
assign n5621 = n3096 | n995;
assign n8160 = n1344 & n11207;
assign n4212 = n9536 & n6755;
assign n10151 = ~(n621 ^ n6844);
assign n2229 = n1560 | n12132;
assign n258 = n1183 | n8740;
assign n9617 = n7914 | n4351;
assign n10440 = n12729 | n552;
assign n3484 = ~(n4644 ^ n9531);
assign n7956 = ~(n1167 ^ n8971);
assign n5131 = ~n461;
assign n3947 = n5014 & n11938;
assign n4019 = ~(n7808 ^ n2306);
assign n10409 = n10122 & n11428;
assign n150 = n11153 & n9763;
assign n7382 = ~n12777;
assign n8546 = n5809 | n1163;
assign n980 = ~(n4932 ^ n6550);
assign n2446 = ~n5363;
assign n9480 = ~(n1313 ^ n5117);
assign n5385 = n7927 & n5358;
assign n9683 = ~(n7718 ^ n1933);
assign n1210 = n3986 & n10990;
assign n7312 = n3746 | n6455;
assign n9451 = n5902 | n4400;
assign n7082 = n6257 & n8845;
assign n11150 = ~n9284;
assign n5427 = ~(n3970 | n1364);
assign n11672 = ~(n11109 ^ n11391);
assign n11069 = n3096 | n7952;
assign n11151 = ~(n2129 ^ n7529);
assign n339 = n10339 | n4913;
assign n8366 = n8354 | n8109;
assign n157 = n2160 | n8725;
assign n4778 = ~n7690;
assign n2260 = ~n7783;
assign n5084 = n7310 | n11202;
assign n12252 = ~(n5014 | n11938);
assign n12264 = ~(n12010 ^ n7886);
assign n10854 = ~n7733;
assign n7969 = n3174 & n12043;
assign n7490 = n2099 | n10854;
assign n11596 = n4778 | n3924;
assign n9740 = n5159 | n2304;
assign n8179 = ~(n9206 ^ n293);
assign n2084 = ~(n5516 ^ n8517);
assign n2845 = ~n5909;
assign n4471 = ~n7276;
assign n10434 = n1937 | n7952;
assign n6575 = n8040 & n4677;
assign n12778 = n8560 & n4532;
assign n4642 = ~n2749;
assign n9691 = ~(n2443 ^ n3391);
assign n4666 = n10838 & n3060;
assign n849 = n5422 & n7885;
assign n1908 = n991 | n354;
assign n1497 = ~(n6452 ^ n8226);
assign n11090 = n7474 | n1681;
assign n4665 = n320 & n8869;
assign n6482 = n10504 | n6682;
assign n5889 = n3096 | n12816;
assign n11729 = n5945 | n11820;
assign n3452 = n752 | n2589;
assign n8584 = n4911 | n4400;
assign n6725 = ~(n5639 ^ n11146);
assign n1580 = n1699 | n1163;
assign n1811 = n5915 | n12080;
assign n6930 = ~(n9744 | n3963);
assign n8673 = ~n9199;
assign n76 = n6669 | n3568;
assign n321 = n8692 | n2421;
assign n12077 = ~(n3559 ^ n11725);
assign n5941 = n12752 & n1425;
assign n5193 = n4660 & n4399;
assign n10287 = ~(n2526 ^ n9331);
assign n9699 = ~n11108;
assign n3669 = n2157 | n8245;
assign n9078 = ~n12704;
assign n1185 = n5964 & n2585;
assign n3013 = ~n2771;
assign n7401 = n12119 | n5468;
assign n10812 = ~(n6415 | n2871);
assign n10745 = n8959 | n11820;
assign n1107 = n7251 | n4264;
assign n12559 = ~n9353;
assign n9997 = n989 | n5497;
assign n10496 = ~(n12463 ^ n3197);
assign n6189 = n6718 | n12771;
assign n6549 = ~(n3334 ^ n2580);
assign n6138 = ~n11999;
assign n955 = n2727 & n2735;
assign n7704 = ~n384;
assign n941 = ~(n289 ^ n11681);
assign n6081 = ~(n8213 ^ n12073);
assign n7530 = n10835 | n795;
assign n9552 = ~(n11702 ^ n4296);
assign n5623 = ~(n11362 | n2314);
assign n7439 = n3620 | n5718;
assign n1904 = ~(n2326 ^ n10869);
assign n476 = ~n12466;
assign n5452 = n5438 | n11986;
assign n6516 = n3096 | n7876;
assign n7513 = n4498 | n2358;
assign n1088 = n8574 & n8739;
assign n1940 = ~(n5830 ^ n6232);
assign n11215 = ~(n3844 ^ n3360);
assign n12510 = ~n11395;
assign n1752 = n1315 & n2211;
assign n10167 = n10671 & n4295;
assign n5338 = n1686 & n2898;
assign n10583 = ~(n8117 ^ n4976);
assign n4635 = n3820 | n9568;
assign n2619 = ~(n8357 ^ n3670);
assign n3502 = ~(n7936 ^ n8298);
assign n7619 = n2326 & n10869;
assign n3306 = ~n12265;
assign n2640 = n5558 & n316;
assign n10507 = ~(n1815 | n6225);
assign n1098 = ~(n3780 ^ n11357);
assign n1880 = ~(n3170 ^ n11583);
assign n2117 = ~(n4756 ^ n2323);
assign n9524 = n12361 | n1413;
assign n632 = n3771 | n3302;
assign n9270 = n3318 & n2675;
assign n6422 = n2136 & n10652;
assign n1932 = ~n533;
assign n9639 = ~n5317;
assign n2485 = n12786 & n5687;
assign n8471 = ~(n4850 ^ n8016);
assign n1501 = ~(n9385 ^ n12529);
assign n11540 = n10157 | n8285;
assign n5279 = n1937 | n9741;
assign n11158 = n1434 | n4887;
assign n4066 = ~(n4753 | n4851);
assign n4259 = ~(n4126 ^ n12608);
assign n1822 = n10344 & n8541;
assign n3605 = n5605 | n3745;
assign n2143 = ~(n5880 ^ n3243);
assign n5255 = ~(n11846 ^ n7117);
assign n4641 = n12322 | n10872;
assign n12631 = ~n585;
assign n12493 = n4692 & n4977;
assign n1252 = n1646 & n11866;
assign n4496 = ~(n7408 ^ n3547);
assign n6691 = n10991 | n6056;
assign n11100 = ~(n4783 | n8840);
assign n12038 = n3822 & n1071;
assign n3928 = ~(n4320 ^ n1840);
assign n863 = ~(n2514 ^ n12097);
assign n2275 = ~(n768 ^ n10131);
assign n12521 = n8251 | n6109;
assign n1068 = n2649 | n9926;
assign n2140 = ~(n1317 ^ n4386);
assign n1341 = n1941 | n9741;
assign n4387 = n752 | n8768;
assign n1011 = n589 | n12321;
assign n827 = ~n7672;
assign n6956 = ~(n10802 ^ n1122);
assign n7740 = ~(n2958 ^ n11663);
assign n12675 = n9544 | n9882;
assign n5741 = ~(n6917 ^ n990);
assign n6536 = ~(n7806 ^ n519);
assign n10554 = ~(n10548 ^ n1579);
assign n7723 = ~n6665;
assign n6717 = ~(n9591 ^ n10044);
assign n6446 = ~(n2248 | n5854);
assign n5949 = n10338 | n6123;
assign n11564 = ~(n10723 ^ n10858);
assign n11909 = ~(n7291 ^ n9523);
assign n10733 = n4219 & n1817;
assign n7586 = ~n3372;
assign n4580 = n3534 & n11350;
assign n8547 = ~(n9547 ^ n3194);
assign n7357 = ~n4554;
assign n7453 = n6231 | n3444;
assign n5583 = ~n2161;
assign n9385 = n2827 & n6170;
assign n1475 = n9389 | n1162;
assign n7860 = n7883 | n1595;
assign n6732 = n11087 | n7183;
assign n9435 = ~(n6178 ^ n6494);
assign n2 = ~(n548 ^ n10859);
assign n8388 = n2022 | n514;
assign n4217 = n4778 | n4913;
assign n4586 = n11307 | n1550;
assign n5951 = ~(n8853 | n9941);
assign n12225 = n347 & n5560;
assign n5158 = ~n6872;
assign n9141 = n752 | n3356;
assign n8791 = ~n2469;
assign n10395 = n3345 & n2925;
assign n3243 = ~(n1493 ^ n4216);
assign n6098 = n11958 | n5538;
assign n2164 = n12237 | n1163;
assign n11806 = ~(n11198 ^ n12166);
assign n11404 = ~(n9652 ^ n1766);
assign n7581 = ~(n1036 | n11520);
assign n1222 = ~n1251;
assign n11504 = ~(n7434 ^ n8063);
assign n8187 = ~n6770;
assign n3730 = n1508 | n9862;
assign n511 = ~n2128;
assign n9703 = ~(n11512 ^ n5065);
assign n4679 = ~(n718 ^ n7454);
assign n4083 = ~(n7171 ^ n1999);
assign n12484 = n1955 & n7008;
assign n9408 = n10506 | n7060;
assign n10154 = ~(n3920 ^ n11164);
assign n12067 = ~n866;
assign n10346 = ~(n6995 | n2405);
assign n1945 = n11097 & n2935;
assign n9661 = n4838 | n12102;
assign n8008 = n582 & n11014;
assign n6686 = n10196 | n4875;
assign n8157 = n5235 & n433;
assign n2699 = n8583 | n10916;
assign n3147 = n4632 | n8024;
assign n9927 = ~(n6167 | n8883);
assign n9584 = ~n4817;
assign n9513 = n12318 & n6900;
assign n3289 = ~(n11674 ^ n7111);
assign n11439 = n1186 & n12849;
assign n7542 = ~(n3964 | n1334);
assign n10368 = ~(n4362 ^ n5115);
assign n9483 = n12395 | n11818;
assign n958 = n1539 | n3911;
assign n3168 = n8127 | n6389;
assign n9254 = ~(n12262 ^ n8253);
assign n1422 = ~n9891;
assign n9825 = n3096 | n9741;
assign n3607 = n10912 & n6143;
assign n10540 = ~(n9379 ^ n5110);
assign n11992 = ~(n7383 | n4893);
assign n5833 = n8026 | n3356;
assign n11937 = ~(n5318 | n1327);
assign n1096 = n2064 & n5122;
assign n9854 = ~(n2695 ^ n9302);
assign n9022 = n8026 | n5012;
assign n525 = n8966 | n3960;
assign n1789 = n9878 | n1163;
assign n9030 = ~n9485;
assign n11354 = n5283 & n2802;
assign n9463 = ~(n7342 ^ n9839);
assign n6031 = ~n1655;
assign n10669 = ~(n9849 ^ n2664);
assign n7726 = n1962 & n3147;
assign n7289 = ~(n6339 ^ n10539);
assign n9007 = n7933 | n10989;
assign n4042 = n12503 | n28;
assign n11949 = ~n5598;
assign n3091 = n8344 | n1756;
assign n11724 = ~(n7592 ^ n2775);
assign n1278 = ~n7685;
assign n2165 = n2862 | n8865;
assign n11106 = n9370 | n7246;
assign n12458 = n12642 | n12185;
assign n9250 = n9170 | n7341;
assign n10415 = ~(n2619 ^ n4978);
assign n3661 = ~(n7051 ^ n12323);
assign n3891 = n8880 & n12629;
assign n481 = n12797 | n12816;
assign n5724 = ~n8381;
assign n352 = ~(n3534 ^ n10914);
assign n12907 = ~(n8562 | n11642);
assign n12841 = n752 | n10903;
assign n7876 = ~n6703;
assign n4858 = n2031 | n650;
assign n11317 = ~(n1304 ^ n7767);
assign n5515 = ~n1139;
assign n7399 = ~(n526 ^ n3690);
assign n4123 = ~(n9317 ^ n12645);
assign n1759 = n5599 & n7256;
assign n1617 = ~(n10647 | n7422);
assign n11744 = n11026 | n9144;
assign n4746 = n76 & n9323;
assign n6150 = n200 & n6906;
assign n4949 = ~(n701 ^ n7036);
assign n8634 = n10142 | n11746;
assign n2349 = ~n10762;
assign n5979 = ~n12657;
assign n12263 = n2217 | n3606;
assign n2130 = n12186 | n6169;
assign n7079 = ~(n8606 ^ n170);
assign n4918 = ~(n882 ^ n11209);
assign n1810 = ~(n4701 ^ n6811);
assign n188 = n11015 & n12578;
assign n6941 = ~n12712;
assign n8426 = ~n3722;
assign n263 = ~(n3503 ^ n11139);
assign n4901 = n131 | n1228;
assign n11202 = n636 | n8740;
assign n11163 = ~n7878;
assign n2452 = ~(n5595 ^ n8170);
assign n10351 = n1695 | n8066;
assign n3067 = n12361 | n6455;
assign n821 = ~(n4257 ^ n20);
assign n12153 = ~(n2730 ^ n10316);
assign n2181 = ~(n11956 ^ n1168);
assign n4153 = n8428 | n1413;
assign n765 = ~n11489;
assign n3726 = n7410 | n3763;
assign n12570 = ~(n144 ^ n7137);
assign n10088 = n7899 | n5485;
assign n2694 = n4498 | n4242;
assign n10353 = n749 | n8676;
assign n4721 = n6977 | n1413;
assign n4166 = n7391 | n10419;
assign n5293 = ~(n1322 ^ n2565);
assign n5910 = ~(n7428 ^ n1113);
assign n10318 = n7449 | n7921;
assign n7405 = ~(n10783 ^ n12039);
assign n3614 = ~n557;
assign n1025 = ~n10336;
assign n5258 = ~n11791;
assign n4101 = n9413 | n9022;
assign n5575 = ~n6877;
assign n3539 = ~(n1945 | n3972);
assign n11115 = ~n5459;
assign n2800 = n182 | n6267;
assign n2246 = ~(n797 ^ n12169);
assign n5863 = ~(n9798 ^ n11404);
assign n10375 = ~(n5681 ^ n4819);
assign n5377 = n8527 | n11948;
assign n1867 = ~(n3384 ^ n2550);
assign n1480 = ~(n10172 ^ n8119);
assign n7516 = ~(n3752 ^ n2920);
assign n3870 = n2834 | n10526;
assign n7880 = ~(n357 ^ n5306);
assign n8660 = n11478 & n5645;
assign n9240 = ~(n12741 ^ n4229);
assign n10739 = n2763 | n789;
assign n2736 = n8514 & n7406;
assign n12375 = ~(n9825 | n8469);
assign n4209 = n10511 | n484;
assign n10393 = ~(n1274 ^ n6492);
assign n200 = ~n10265;
assign n8347 = n2456 | n8648;
assign n12523 = ~(n3706 ^ n2625);
assign n3344 = ~n6575;
assign n2218 = ~(n1751 ^ n4178);
assign n1238 = n11446 | n9084;
assign n2767 = ~(n12266 | n10337);
assign n12910 = ~(n3492 ^ n698);
assign n1817 = n9228 | n10931;
assign n1992 = n8026 | n6084;
assign n1513 = ~(n1675 ^ n344);
assign n12300 = ~(n10033 | n11823);
assign n4500 = n4911 | n1851;
assign n4583 = n1052 & n266;
assign n5653 = ~(n10847 ^ n12626);
assign n11335 = n3743 | n11698;
assign n5816 = n10202 | n9729;
assign n8479 = ~n6766;
assign n9963 = ~n8628;
assign n8198 = ~(n7777 ^ n11872);
assign n5843 = ~(n12516 | n720);
assign n4660 = n2552 | n6974;
assign n9766 = ~(n8567 ^ n341);
assign n9720 = n12755 | n9954;
assign n7931 = ~(n3046 ^ n7201);
assign n4468 = n4414 & n3781;
assign n9898 = ~(n5155 ^ n1860);
assign n424 = ~n720;
assign n2552 = ~n10973;
assign n9130 = n8629 & n1498;
assign n465 = ~(n3642 ^ n7601);
assign n5085 = ~(n7383 ^ n12914);
assign n4040 = ~n390;
assign n11256 = ~(n2110 ^ n11776);
assign n620 = ~(n3442 ^ n2694);
assign n11013 = n8552 | n8655;
assign n8580 = n3303 & n1744;
assign n8955 = n1183 | n4913;
assign n8802 = ~(n1123 ^ n3729);
assign n10506 = n9373 | n4654;
assign n9166 = n7310 & n11202;
assign n12128 = ~(n7554 ^ n9792);
assign n12488 = n9977 | n4375;
assign n9779 = n11825 & n10592;
assign n7053 = n11902 & n6883;
assign n818 = ~(n4401 | n9629);
assign n9259 = ~n8418;
assign n10419 = ~n5320;
assign n6070 = n11592 & n12419;
assign n3208 = n9625 & n5937;
assign n6247 = n5423 | n1528;
assign n979 = ~(n7940 | n818);
assign n7773 = n2499 & n5418;
assign n4561 = n12119 | n5326;
assign n3497 = n4694 | n2768;
assign n1859 = n7839 | n12816;
assign n7314 = ~(n10850 | n9605);
assign n722 = ~(n4390 ^ n7748);
assign n3601 = n2464 & n11023;
assign n7218 = n6636 | n12215;
assign n11297 = n107 & n10880;
assign n4845 = n4354 | n11639;
assign n11854 = n3082 | n2875;
assign n3509 = n527 & n9816;
assign n8931 = ~(n12622 ^ n3919);
assign n4886 = ~(n9222 ^ n5162);
assign n6546 = n1086 | n123;
assign n6848 = n2236 & n3277;
assign n5607 = n4778 | n8109;
assign n2848 = n7774 | n7127;
assign n383 = n1887 & n7903;
assign n7190 = ~n4612;
assign n9669 = n656 & n10580;
assign n4631 = ~(n8348 ^ n111);
assign n678 = n3243 | n5880;
assign n9194 = n6621 & n10910;
assign n4433 = n284 | n10693;
assign n3094 = ~(n8577 ^ n8249);
assign n12 = n8412 & n3521;
assign n723 = ~(n4821 ^ n48);
assign n12336 = ~(n3232 ^ n5997);
assign n12134 = ~(n7305 | n8872);
assign n125 = ~n1948;
assign n3663 = ~(n10116 ^ n4679);
assign n8768 = ~n10439;
assign n764 = ~(n634 ^ n11178);
assign n4707 = n3772 | n4171;
assign n10321 = ~(n3799 ^ n4590);
assign n9928 = ~(n8584 ^ n7644);
assign n9406 = ~(n11839 ^ n12876);
assign n5905 = ~(n8455 ^ n6891);
assign n7962 = ~n2015;
assign n2930 = n9428 | n9981;
assign n3042 = n11182 & n4200;
assign n3697 = ~(n2819 ^ n11830);
assign n2723 = ~(n2787 | n1208);
assign n1972 = n11281 | n4629;
assign n5345 = n8959 | n7876;
assign n12405 = ~(n4715 ^ n6503);
assign n6683 = n1471 & n11876;
assign n6934 = n10738 | n3150;
assign n4926 = n5915 | n12535;
assign n12314 = n9564 ^ n7680;
assign n2125 = n6697 | n12225;
assign n9157 = ~(n2976 ^ n11495);
assign n2473 = n2188 & n8006;
assign n5064 = n11958 | n11820;
assign n12768 = ~n8504;
assign n7383 = n10142 | n7389;
assign n5139 = ~(n11178 | n634);
assign n1153 = n9273 & n11048;
assign n12605 = n5214 & n2616;
assign n7695 = ~(n12144 ^ n3153);
assign n7561 = n11165 & n352;
assign n10786 = ~(n12325 ^ n7556);
assign n3345 = n8704 | n5761;
assign n10143 = ~(n5412 ^ n12255);
assign n10200 = n12416 | n9961;
assign n6106 = ~n3499;
assign n879 = n326 & n2904;
assign n9923 = ~(n10788 ^ n8523);
assign n4323 = n4667 & n6199;
assign n8379 = ~(n4984 ^ n1153);
assign n223 = ~(n5627 ^ n1770);
assign n11226 = ~n2418;
assign n6100 = ~(n11378 | n11991);
assign n441 = n12267 | n12890;
assign n1585 = ~(n3386 | n129);
assign n9853 = ~n6618;
assign n3691 = n8699 | n228;
assign n7328 = n6219 & n4959;
assign n10197 = n1539 | n10066;
assign n9027 = ~(n10777 ^ n10171);
assign n3769 = ~(n6250 ^ n93);
assign n10452 = ~(n3972 ^ n4477);
assign n10803 = n4911 | n1915;
assign n9419 = ~(n9567 ^ n5754);
assign n8548 = n10265 & n11132;
assign n6432 = ~(n12618 ^ n10353);
assign n8129 = ~(n5606 ^ n7249);
assign n0 = n3743 | n9568;
assign n6484 = n5815 | n6018;
assign n11083 = n1474 | n9633;
assign n1081 = n792 | n2880;
assign n12618 = ~(n10917 | n6238);
assign n4441 = n2385 | n5803;
assign n4356 = n3501 | n4924;
assign n6524 = ~n6604;
assign n2422 = ~n3384;
assign n4867 = n12494 | n12719;
assign n10625 = ~n2104;
assign n5369 = n773 | n12405;
assign n8025 = n12733 & n5820;
assign n3140 = n191 | n2076;
assign n11302 = n7918 | n544;
assign n434 = ~(n12739 | n3108);
assign n11375 = n12946 & n8265;
assign n4140 = ~n6591;
assign n1688 = n10835 | n28;
assign n6255 = n11914 & n6839;
assign n9134 = n636 | n9586;
assign n5014 = ~(n12564 ^ n8003);
assign n426 = n3118 | n2203;
assign n6388 = ~n11062;
assign n5632 = ~(n8442 ^ n4745);
assign n3912 = n11588 | n5476;
assign n3252 = n6095 & n781;
assign n8043 = ~(n6981 ^ n9149);
assign n1046 = ~(n9837 ^ n12126);
assign n4260 = ~(n2746 ^ n7887);
assign n356 = ~(n12882 ^ n11249);
assign n12335 = ~n1577;
assign n11739 = n11433 | n7952;
assign n10962 = ~n2978;
assign n9452 = ~n3833;
assign n6001 = n3821 | n4701;
assign n6078 = n5915 | n7382;
assign n4438 = ~(n9995 ^ n10754);
assign n9148 = ~n3726;
assign n11862 = n2071 & n10323;
assign n272 = ~(n377 ^ n1492);
assign n5496 = ~n9016;
assign n2878 = n3692 & n7649;
assign n12620 = ~(n61 ^ n8393);
assign n4306 = ~(n1543 ^ n1294);
assign n4617 = ~n2665;
assign n3968 = n11090 & n7010;
assign n6468 = n4396 | n10296;
assign n8432 = ~n5756;
assign n6347 = n11958 | n10903;
assign n4712 = ~(n5812 ^ n5984);
assign n12653 = n4433 & n2681;
assign n8053 = n9241 & n7946;
assign n5958 = ~(n158 | n9260);
assign n7386 = ~(n407 ^ n4006);
assign n5414 = n989 | n7424;
assign n5490 = ~(n855 ^ n5190);
assign n2322 = n3650 | n1285;
assign n8495 = ~(n9101 ^ n9516);
assign n1877 = n12237 | n12686;
assign n8686 = n5748 | n5639;
assign n3558 = n5563 & n5749;
assign n4554 = n4111 & n4215;
assign n5169 = ~(n11095 ^ n10087);
assign n5415 = ~n5504;
assign n9342 = n8851 & n6768;
assign n9146 = ~(n1039 | n5611);
assign n8545 = ~(n7338 ^ n10267);
assign n1077 = ~n9281;
assign n10557 = ~(n10230 ^ n10273);
assign n3747 = n5530 | n9586;
assign n11020 = ~(n4254 ^ n5926);
assign n5847 = ~(n8509 | n3099);
assign n5431 = ~n6917;
assign n1055 = n4270 ^ n7579;
assign n10789 = ~(n3343 ^ n7849);
assign n2771 = n7364 & n1843;
assign n1325 = n4707 | n495;
assign n9831 = ~(n4838 ^ n5901);
assign n9284 = n7768 & n2631;
assign n4725 = n11773 & n7473;
assign n2396 = ~(n3050 ^ n11524);
assign n4517 = ~(n4577 ^ n4887);
assign n436 = n1664 & n6851;
assign n6055 = ~n4806;
assign n1016 = ~(n3419 ^ n4610);
assign n10578 = n2081 | n4068;
assign n11471 = n9170 | n1915;
assign n7497 = n4124 & n11935;
assign n2318 = n11779 & n2256;
assign n10160 = ~(n555 ^ n6841);
assign n7752 = n9170 | n11827;
assign n4600 = n8607 & n371;
assign n789 = n4059 | n3911;
assign n12143 = ~(n1651 | n12695);
assign n10650 = ~(n8277 ^ n9724);
assign n8543 = ~n2954;
assign n5300 = ~(n12293 ^ n5833);
assign n6913 = n11470 & n7264;
assign n333 = n1099 & n11183;
assign n5688 = n1619 & n3477;
assign n8739 = n9366 | n3709;
assign n11580 = n4787 | n1889;
assign n5234 = n6151 & n11219;
assign n11362 = n2446 & n11631;
assign n7952 = ~n1209;
assign n6049 = n4059 | n1738;
assign n8707 = ~(n6628 | n11372);
assign n1474 = ~(n7459 | n4490);
assign n11033 = n7777 | n11872;
assign n6424 = ~(n7182 ^ n5905);
assign n3776 = n7041 | n2932;
assign n6987 = ~(n10865 ^ n8849);
assign n11058 = n8704 & n5761;
assign n9801 = n1937 | n11775;
assign n1801 = ~(n12027 | n10176);
assign n2044 = n11846 & n7117;
assign n1257 = n4552 | n12184;
assign n3332 = n2946 & n7488;
assign n11464 = ~(n5089 ^ n10823);
assign n7545 = n9492 & n4420;
assign n2075 = ~(n5650 | n11675);
assign n136 = ~(n8140 | n9877);
assign n1427 = ~(n8531 ^ n11985);
assign n3963 = n994 | n1738;
assign n4263 = ~(n3971 ^ n10897);
assign n1136 = ~(n4587 ^ n4975);
assign n6947 = ~(n11115 ^ n3320);
assign n1597 = ~(n11052 ^ n7719);
assign n12120 = ~n7270;
assign n3902 = n2040 & n1605;
assign n1792 = ~(n7609 ^ n7907);
assign n12638 = n1728 | n7627;
assign n7338 = ~n5081;
assign n4383 = ~(n8714 | n9608);
assign n4732 = ~(n8491 ^ n10287);
assign n7498 = n1677 & n6235;
assign n7337 = n10566 & n6730;
assign n5266 = ~n2650;
assign n1386 = n5448 | n932;
assign n11750 = ~n5233;
assign n9271 = n10835 | n1476;
assign n2720 = n8354 | n10854;
assign n4420 = n3096 | n2815;
assign n8224 = ~(n237 | n4556);
assign n4329 = ~(n2011 ^ n6268);
assign n11742 = ~n2571;
assign n2323 = ~(n4552 ^ n12011);
assign n12209 = ~(n9695 ^ n10708);
assign n302 = n967 & n6615;
assign n4484 = ~(n5391 ^ n11320);
assign n5691 = ~n1878;
assign n8554 = ~n3070;
assign n2821 = ~(n8124 | n5367);
assign n12522 = n7709 | n4527;
assign n6765 = n1715 | n11329;
assign n1574 = n2071 | n10323;
assign n6075 = n9170 | n1455;
assign n6290 = ~n2109;
assign n10679 = ~(n9967 | n7357);
assign n5056 = ~(n9598 | n4395);
assign n10992 = n3127 | n1455;
assign n2481 = ~(n12112 ^ n12364);
assign n6140 = n12216 & n10672;
assign n7747 = n4728 | n10505;
assign n12337 = n12271 & n12707;
assign n831 = n6685 | n8604;
assign n7508 = ~n8018;
assign n9443 = ~(n12783 ^ n12943);
assign n772 = ~(n4506 ^ n345);
assign n10476 = ~(n12573 ^ n1610);
assign n7013 = ~(n2641 ^ n11574);
assign n665 = ~n12540;
assign n7248 = ~(n12338 ^ n2528);
assign n8206 = ~(n10178 ^ n9727);
assign n10013 = n587 & n12665;
assign n3901 = n994 | n11430;
assign n11138 = ~n11393;
assign n8755 = ~n11687;
assign n12700 = n11433 | n6455;
assign n2553 = ~(n7590 ^ n10490);
assign n569 = ~n1037;
assign n5476 = ~(n11614 ^ n7152);
assign n8934 = ~(n3319 ^ n516);
assign n5141 = n4873 | n11880;
assign n12564 = ~(n10181 ^ n10126);
assign n7855 = n10471 | n9765;
assign n4069 = ~(n11001 ^ n6528);
assign n1927 = ~(n4367 | n119);
assign n6697 = n3743 | n4642;
assign n10960 = n6373 | n1047;
assign n2015 = n4466 & n9793;
assign n8155 = ~(n9274 | n10814);
assign n7486 = n2260 & n2454;
assign n10994 = ~(n11879 ^ n7655);
assign n662 = ~(n6725 ^ n9344);
assign n7939 = n2456 | n5781;
assign n5200 = n8552 | n1932;
assign n10998 = n12025 & n11407;
assign n9455 = ~n5164;
assign n3414 = n9617 & n139;
assign n11524 = n7449 | n1509;
assign n5333 = ~(n60 ^ n11213);
assign n8127 = ~n11821;
assign n2413 = n137 & n2802;
assign n926 = n5345 | n5711;
assign n7849 = ~(n1890 ^ n6436);
assign n10930 = ~(n4855 | n6753);
assign n8675 = n6551 & n2086;
assign n1383 = ~n6056;
assign n6609 = ~(n12716 ^ n10524);
assign n9629 = ~(n10453 ^ n7597);
assign n1509 = ~n10848;
assign n8843 = ~(n10579 ^ n1888);
assign n4750 = n8870 | n10854;
assign n10564 = n8051 | n3966;
assign n9885 = ~n3194;
assign n1952 = n3512 | n10293;
assign n12793 = ~(n991 ^ n5664);
assign n9961 = n6368 & n1309;
assign n9635 = ~(n9231 ^ n6395);
assign n3557 = n8810 & n318;
assign n9424 = ~(n4337 ^ n6558);
assign n2529 = n9878 | n5326;
assign n2628 = ~(n10756 | n3373);
assign n10120 = ~(n573 ^ n11044);
assign n9609 = ~(n12234 | n7292);
assign n12590 = ~(n3810 | n3181);
assign n10882 = n5765 | n4654;
assign n3949 = n11571 & n5511;
assign n4539 = n6227 & n11129;
assign n12011 = ~(n1637 ^ n11325);
assign n8600 = n12705 & n2509;
assign n12406 = ~n2108;
assign n5005 = ~(n680 | n2996);
assign n10046 = ~(n5903 | n7119);
assign n12757 = n8476 & n11967;
assign n1831 = ~n12588;
assign n400 = ~(n1919 ^ n12615);
assign n6157 = n4365 & n4323;
assign n6174 = ~(n4165 ^ n6878);
assign n10856 = ~n11642;
assign n5411 = ~(n604 ^ n1329);
assign n4308 = ~n11365;
assign n2166 = ~(n2452 ^ n11298);
assign n342 = n10960 & n10315;
assign n8002 = n752 | n11410;
assign n4221 = ~n2364;
assign n6751 = ~(n769 ^ n3129);
assign n4808 = n4841 & n6456;
assign n6537 = n12365 & n11406;
assign n9434 = ~(n5640 ^ n6840);
assign n6015 = n6718 | n8830;
assign n11725 = ~(n5410 ^ n460);
assign n8049 = n12666 & n3624;
assign n4647 = n6577 | n995;
assign n9258 = n11518 & n878;
assign n6634 = ~n12533;
assign n10455 = n3687 & n532;
assign n12354 = ~(n450 ^ n11516);
assign n5226 = n7630 & n5736;
assign n12646 = n8405 | n3224;
assign n1873 = ~(n10637 ^ n12714);
assign n12886 = n4167 | n6892;
assign n248 = ~(n8104 ^ n7934);
assign n1189 = ~n4707;
assign n8898 = n3810 & n3181;
assign n284 = n7116 | n3903;
assign n6872 = n11033 & n8038;
assign n975 = n11719 | n5497;
assign n5521 = ~(n4120 ^ n10032);
assign n11968 = n8428 | n7952;
assign n6737 = n3773 | n12287;
assign n10489 = n6436 & n7645;
assign n10531 = n1937 | n6197;
assign n10441 = ~(n12303 ^ n6904);
assign n285 = ~(n3015 ^ n2294);
assign n8377 = n4283 | n5524;
assign n11632 = ~(n11501 ^ n11188);
assign n9053 = ~(n1503 | n2839);
assign n3855 = ~n5973;
assign n11625 = n5794 | n4340;
assign n11705 = ~(n5235 ^ n11927);
assign n7568 = ~(n1952 ^ n2092);
assign n7009 = n9311 & n9534;
assign n11614 = ~(n7131 ^ n8807);
assign n12304 = ~n8952;
assign n4310 = ~n8486;
assign n2144 = n1571 & n1422;
assign n8928 = ~(n12249 ^ n3613);
assign n8644 = ~n5069;
assign n6584 = ~(n3125 ^ n11199);
assign n9730 = ~n11352;
assign n5684 = n8759 & n12709;
assign n10122 = ~n12692;
assign n10127 = n722 & n3987;
assign n4113 = ~n1639;
assign n3525 = ~(n8221 ^ n5445);
assign n1850 = ~(n667 ^ n10978);
assign n6321 = ~(n6222 | n3323);
assign n6880 = n6577 | n7395;
assign n7805 = ~(n3163 ^ n8381);
assign n8262 = ~(n1241 ^ n492);
assign n5709 = ~(n10381 | n6177);
assign n3009 = n5945 | n5540;
assign n2627 = ~(n5776 ^ n10454);
assign n9470 = ~n6799;
assign n8924 = n9262 | n4527;
assign n11429 = ~n10512;
assign n12695 = ~(n12167 | n4774);
assign n7713 = n10750 | n1932;
assign n10502 = n10157 | n9568;
assign n5947 = ~(n5992 ^ n12384);
assign n1464 = n2743 & n8597;
assign n1933 = ~(n5679 ^ n2963);
assign n1938 = ~n5302;
assign n10095 = n3425 | n7938;
assign n7323 = n3681 | n7492;
assign n10944 = ~n10059;
assign n10852 = ~(n7665 ^ n4557);
assign n488 = ~n8015;
assign n11700 = n1183 | n8655;
assign n2459 = n2217 | n7921;
assign n11096 = ~(n4923 ^ n2693);
assign n9649 = ~(n6649 | n542);
assign n7360 = ~(n11132 ^ n200);
assign n2664 = n686 | n11775;
assign n7454 = ~(n5292 ^ n369);
assign n9149 = n11923 | n7921;
assign n5629 = ~(n12590 | n11035);
assign n7503 = ~(n3808 | n8460);
assign n5823 = n12237 | n826;
assign n6772 = n2766 | n1770;
assign n3201 = n10290 ^ n3732;
assign n10973 = ~(n6899 ^ n8856);
assign n2033 = ~(n9712 ^ n7511);
assign n507 = n4322 | n512;
assign n5012 = ~n2024;
assign n2432 = ~(n12530 ^ n12779);
assign n2382 = ~(n6478 ^ n5973);
assign n2543 = ~(n8307 | n3539);
assign n431 = n8552 | n10422;
assign n12181 = ~(n10505 ^ n11441);
assign n10493 = n11944 & n5389;
assign n2706 = n4116 & n7188;
assign n12725 = n1937 | n5538;
assign n9004 = ~(n1987 | n3049);
assign n3490 = ~(n1616 | n1002);
assign n7600 = ~(n2978 ^ n6507);
assign n9520 = n11120 | n12373;
assign n4623 = ~n10409;
assign n8320 = n3617 | n9188;
assign n738 = n3653 | n5764;
assign n1755 = n2073 & n12028;
assign n3353 = ~n7925;
assign n6299 = ~(n7292 ^ n4786);
assign n6472 = n6577 | n8768;
assign n4717 = n11552 | n9568;
assign n8524 = ~n2577;
assign n1347 = n5809 | n12535;
assign n12060 = ~(n9663 ^ n6623);
assign n10283 = n12767 & n6780;
assign n6492 = ~(n3251 ^ n6134);
assign n5915 = ~n2530;
assign n9305 = n11887 | n5468;
assign n3455 = n1708 | n12114;
assign n5801 = n1183 | n7382;
assign n11836 = ~(n9223 ^ n9747);
assign n2604 = n737 & n6132;
assign n11174 = ~(n8308 | n6581);
assign n3223 = ~(n2182 ^ n11106);
assign n3039 = n9196 | n8349;
assign n1093 = n6398 & n9442;
assign n3144 = ~n7327;
assign n192 = ~n8053;
assign n11050 = n5496 & n9603;
assign n1242 = n7283 | n4400;
assign n4738 = ~(n3140 | n3447);
assign n8623 = n7293 | n1641;
assign n4943 = n6098 & n1845;
assign n2737 = n3767 & n7600;
assign n9626 = ~(n2759 ^ n16);
assign n8121 = ~(n6653 ^ n2956);
assign n11849 = n1737 & n11299;
assign n9569 = ~(n8483 ^ n2495);
assign n3549 = n7704 | n9671;
assign n8643 = ~n217;
assign n5093 = n5314 & n2749;
assign n6457 = ~n2788;
assign n2841 = ~(n9024 | n10201);
assign n10834 = n12173 & n1405;
assign n11628 = ~(n308 ^ n1500);
assign n331 = ~n6717;
assign n4097 = n4904 | n701;
assign n7276 = n5439 & n8083;
assign n9255 = n3672 & n8255;
assign n11880 = ~n6858;
assign n11071 = n7839 | n11775;
assign n9955 = n10005 ^ n791;
assign n1125 = ~(n6974 ^ n5719);
assign n3996 = n589 & n12321;
assign n2177 = ~(n7442 ^ n568);
assign n12568 = ~n4257;
assign n9538 = n7116 | n6455;
assign n12834 = ~(n5522 ^ n115);
assign n5743 = ~(n2418 | n5274);
assign n6978 = ~(n2516 ^ n1064);
assign n7292 = n627 | n11964;
assign n12223 = n10142 | n8859;
assign n1685 = ~n12956;
assign n1963 = n4373 | n5628;
assign n9653 = ~n12198;
assign n897 = ~n6612;
assign n7410 = n12234 & n7292;
assign n8853 = ~n2055;
assign n10520 = ~n816;
assign n4779 = n1453 ^ n1000;
assign n8181 = n8026 | n11896;
assign n5051 = ~(n4914 ^ n10227);
assign n9677 = n12853 | n12735;
assign n7180 = ~n10642;
assign n30 = ~(n12089 ^ n5879);
assign n3258 = n273 & n9126;
assign n7171 = n6677 & n12175;
assign n10738 = n12361 | n7952;
assign n4726 = n2872 | n12816;
assign n4609 = ~(n2699 ^ n10941);
assign n108 = n12062 | n73;
assign n12394 = n3780 & n6329;
assign n2207 = n2740 | n2844;
assign n2555 = ~(n12866 ^ n194);
assign n22 = ~n5947;
assign n10111 = ~(n3448 ^ n12744);
assign n10147 = n9108 & n3983;
assign n7783 = n10196 | n4654;
assign n4806 = ~(n7289 ^ n12141);
assign n7639 = ~n8359;
assign n10242 = n128 | n5460;
assign n10212 = n2332 | n6034;
assign n7976 = ~(n5867 ^ n11522);
assign n3668 = ~n4432;
assign n2676 = ~n6980;
assign n6626 = ~(n1147 ^ n729);
assign n7375 = ~(n11309 ^ n7738);
assign n3973 = ~(n2578 ^ n5842);
assign n7885 = n5879 | n2940;
assign n12293 = ~(n3946 | n7724);
assign n3099 = ~(n11117 ^ n7628);
assign n4338 = n12853 | n10854;
assign n5827 = ~(n814 ^ n2847);
assign n10505 = ~(n5524 ^ n7877);
assign n7802 = n9905 | n10792;
assign n10276 = ~(n5539 ^ n7430);
assign n10488 = ~(n1061 ^ n2685);
assign n10413 = ~(n7783 ^ n3710);
assign n8835 = n10835 | n9078;
assign n2463 = n1044 & n6668;
assign n346 = n11958 | n8414;
assign n5243 = ~(n12109 ^ n3355);
assign n948 = n4900 | n2219;
assign n3299 = ~(n12584 | n5733);
assign n2442 = ~(n8085 | n5180);
assign n5461 = ~(n4490 ^ n7459);
assign n8364 = ~n11024;
assign n10826 = n6977 | n11775;
assign n2097 = n2099 | n7928;
assign n5065 = ~(n7651 ^ n10119);
assign n2431 = ~(n7618 ^ n12836);
assign n1291 = ~n11094;
assign n1306 = ~(n7327 ^ n2971);
assign n10683 = n11415 & n12606;
assign n2102 = ~(n6462 ^ n2094);
assign n1060 = ~(n4633 ^ n2255);
assign n10604 = n9878 | n8109;
assign n10107 = ~(n1652 ^ n5498);
assign n6248 = ~(n1524 | n8540);
assign n4990 = n5964 & n7265;
assign n2920 = ~(n2116 ^ n12452);
assign n3210 = n3820 | n9144;
assign n9915 = n6373 | n1476;
assign n9088 = ~(n12208 ^ n10017);
assign n10326 = ~n9060;
assign n12313 = n7591 | n1787;
assign n5080 = ~(n10630 ^ n12861);
assign n7097 = n11884 | n5992;
assign n233 = n6977 | n10903;
assign n11357 = ~(n8598 ^ n5581);
assign n3316 = n6283 | n3543;
assign n9190 = n5355 | n10419;
assign n2641 = ~(n6734 | n9049);
assign n3933 = n6534 | n10826;
assign n1709 = n7552 | n12553;
assign n8480 = ~(n1790 ^ n2016);
assign n8891 = n6162 | n12432;
assign n3298 = n8552 | n3224;
assign n5066 = ~(n6015 ^ n8673);
assign n8386 = n1183 | n3924;
assign n6621 = n6877 & n7946;
assign n10616 = ~(n8990 ^ n11496);
assign n7172 = n7804 & n10341;
assign n10799 = ~n1672;
assign n2587 = n3324 | n28;
assign n3350 = ~(n8585 ^ n12187);
assign n9980 = n1459 & n10330;
assign n256 = ~(n10245 ^ n8760);
assign n4792 = n1011 & n864;
assign n7678 = ~n1395;
assign n2528 = ~n7865;
assign n5664 = n10750 | n8109;
assign n4528 = n2332 & n6034;
assign n1207 = n989 | n7389;
assign n9178 = n7509 | n3117;
assign n5182 = n6504 | n3863;
assign n7489 = n9076 & n4032;
assign n3467 = ~(n6824 ^ n6614);
assign n3326 = n5331 & n1067;
assign n10880 = n1699 | n9188;
assign n377 = ~(n4440 ^ n6083);
assign n6818 = n11337 | n11092;
assign n9280 = ~n6359;
assign n870 = n5638 | n10767;
assign n5962 = n343 & n7278;
assign n6102 = n2330 & n6450;
assign n1183 = ~n2515;
assign n11587 = n6626 | n6106;
assign n3027 = ~(n7883 ^ n4341);
assign n7216 = ~(n5850 ^ n3218);
assign n11435 = ~(n3491 ^ n2954);
assign n4188 = ~(n5341 ^ n11947);
assign n6171 = ~n6865;
assign n2728 = n289 & n11772;
assign n4909 = n3282 & n2907;
assign n5247 = ~(n7463 ^ n5146);
assign n7715 = n2689 | n10649;
assign n11526 = n12392 | n2231;
assign n1676 = n10450 | n117;
assign n8095 = n5329 | n9898;
assign n6376 = ~n3574;
assign n11085 = n11225 & n12559;
assign n1378 = ~(n3949 | n5935);
assign n1465 = n9373 | n9568;
assign n3325 = n10350 | n7081;
assign n2031 = ~(n12437 ^ n11238);
assign n6586 = n3386 & n129;
assign n8636 = ~(n3159 ^ n3459);
assign n7506 = ~n12947;
assign n1599 = n11923 | n9568;
assign n11961 = n7495 | n5497;
assign n766 = n3944 & n334;
assign n4797 = n2496 & n10452;
assign n9888 = n5337 | n3492;
assign n8339 = n11552 | n4474;
assign n3606 = ~n1478;
assign n4759 = n4498 | n7341;
assign n11715 = ~(n7008 ^ n155);
assign n12625 = n3909 & n6105;
assign n11175 = ~n12895;
assign n12277 = ~(n3217 ^ n5669);
assign n2402 = n2403 & n6763;
assign n3477 = ~n8975;
assign n4715 = ~(n9113 ^ n12032);
assign n3261 = n6426 | n11009;
assign n6045 = ~(n12016 ^ n6082);
assign n4234 = n994 | n5497;
assign n2881 = ~(n11451 | n6466);
assign n901 = n3746 | n8414;
assign n7413 = ~n9651;
assign n1644 = ~(n7374 ^ n7805);
assign n12835 = ~n5032;
assign n8832 = ~n3691;
assign n910 = n7283 | n4242;
assign n2434 = ~(n1507 ^ n12153);
assign n1651 = ~(n4972 | n2542);
assign n329 = ~(n12949 ^ n8289);
assign n10113 = n9648 & n5802;
assign n9181 = ~(n9094 ^ n5113);
assign n667 = ~(n11608 ^ n3839);
assign n4698 = ~n1445;
assign n6724 = ~(n12106 ^ n8284);
assign n2665 = n7436 & n11023;
assign n10670 = n8969 | n10961;
assign n12916 = n9413 & n9022;
assign n11509 = ~(n3059 | n10126);
assign n5003 = n994 | n510;
assign n7571 = ~n186;
assign n684 = ~n12306;
assign n7774 = ~(n5003 ^ n892);
assign n4915 = ~(n8486 ^ n2411);
assign n8469 = n807 | n12816;
assign n8875 = n9383 & n8195;
assign n9731 = n1072 & n2975;
assign n501 = n6218 & n2156;
assign n12331 = ~(n5350 | n3540);
assign n1791 = ~n7527;
assign n5181 = n12119 | n12686;
assign n3828 = n10387 | n3019;
assign n4989 = n718 & n1643;
assign n12629 = n7951 | n7215;
assign n1369 = ~(n4166 ^ n4261);
assign n3764 = n10108 | n6389;
assign n3396 = n3096 | n11775;
assign n11701 = ~n7321;
assign n12411 = n2187 & n9061;
assign n2940 = ~(n83 | n9710);
assign n12894 = ~(n3109 ^ n1103);
assign n8254 = ~n11796;
assign n1675 = n3743 | n7506;
assign n9291 = ~n719;
assign n1042 = n9411 | n12408;
assign n8831 = ~(n10154 ^ n5955);
assign n6507 = n4778 | n826;
assign n132 = ~(n4026 | n12410);
assign n5649 = n2175 & n1709;
assign n451 = ~(n1126 ^ n6970);
assign n1541 = ~(n10222 ^ n6842);
assign n7237 = ~(n9055 | n8077);
assign n9697 = ~(n3906 | n11203);
assign n1240 = n3746 | n2815;
assign n11461 = ~(n4131 ^ n3973);
assign n10916 = ~n806;
assign n7640 = n6373 | n795;
assign n1075 = n3013 | n10567;
assign n8234 = ~(n4692 | n4977);
assign n7609 = ~(n12604 ^ n11118);
assign n564 = n6986 & n8595;
assign n12175 = n5399 | n5400;
assign n2451 = ~(n4635 ^ n12369);
assign n3240 = ~n6558;
assign n11272 = n12530 | n12779;
assign n4340 = ~(n6859 ^ n10268);
assign n11955 = n3504 & n524;
assign n9214 = ~n1580;
assign n8128 = ~(n2124 ^ n3553);
assign n11063 = n4207 & n3371;
assign n9071 = ~n5684;
assign n11875 = ~(n3297 ^ n10757);
assign n9313 = ~n8304;
assign n4933 = ~n11677;
assign n556 = n5200 | n1010;
assign n7541 = ~n3724;
assign n5275 = ~(n10730 | n11104);
assign n3381 = n191 | n1079;
assign n520 = ~(n905 ^ n3168);
assign n4252 = n12041 & n10416;
assign n5423 = n9373 | n9144;
assign n7986 = ~(n3347 | n8179);
assign n4082 = ~(n1820 ^ n3206);
assign n4125 = ~(n2202 | n8402);
assign n1258 = ~(n11503 | n10388);
assign n11956 = ~(n11479 ^ n4083);
assign n3493 = n5519 | n1441;
assign n1914 = n5945 | n995;
assign n5667 = n11455 | n7614;
assign n3125 = ~(n12959 ^ n6355);
assign n12269 = ~(n3570 | n9972);
assign n12127 = n9079 | n6414;
assign n10903 = ~n11023;
assign n9608 = ~(n5929 ^ n8196);
assign n829 = n8552 | n5468;
assign n11116 = ~(n12056 | n12678);
assign n1998 = n7534 | n2079;
assign n2366 = ~n7957;
assign n11963 = ~n7463;
assign n12507 = n5915 | n8259;
assign n6478 = ~(n1220 ^ n1410);
assign n10228 = ~(n3873 ^ n9320);
assign n8074 = n8836 | n3941;
assign n4830 = ~n7364;
assign n12305 = ~(n1468 ^ n9097);
assign n2013 = n4151 & n3840;
assign n6689 = ~(n7720 ^ n1732);
assign n6629 = n2824 & n10042;
assign n5643 = ~(n6983 ^ n10037);
assign n12574 = ~n4989;
assign n9124 = n5684 & n563;
assign n2799 = ~(n98 ^ n5768);
assign n1152 = ~(n5393 ^ n6733);
assign n8553 = ~(n12932 ^ n2320);
assign n5503 = n12776 & n12587;
assign n2240 = ~(n2965 ^ n5968);
assign n12694 = n3025 | n6054;
assign n8648 = ~n6806;
assign n10762 = n7388 & n12704;
assign n4102 = ~(n12003 ^ n10876);
assign n10595 = n7959 | n2725;
assign n12467 = ~n6356;
assign n10596 = n7539 & n1328;
assign n3929 = n6137 & n9404;
assign n9756 = ~(n3479 ^ n4505);
assign n8413 = n3560 | n3505;
assign n3453 = ~(n7739 | n9057);
assign n6958 = ~(n4316 ^ n943);
assign n10841 = ~(n11147 ^ n12850);
assign n6769 = n1156 | n871;
assign n7999 = n1362 | n8878;
assign n6454 = ~n1236;
assign n6366 = ~(n11172 ^ n4832);
assign n9850 = ~(n4250 ^ n7101);
assign n11097 = ~n10522;
assign n8867 = ~(n12785 ^ n3806);
assign n1930 = ~(n7366 ^ n10062);
assign n549 = ~(n337 ^ n12329);
assign n896 = ~n4119;
assign n5337 = n8373 | n1940;
assign n11745 = ~n1419;
assign n10823 = n4628 | n5468;
assign n5079 = ~(n1528 ^ n2273);
assign n8046 = n9308 & n9562;
assign n2290 = ~(n3132 ^ n435);
assign n8850 = ~(n7632 ^ n4518);
assign n7254 = ~(n7697 ^ n8566);
assign n1604 = ~(n11 | n10159);
assign n10190 = ~n3973;
assign n6348 = ~(n8235 | n4597);
assign n571 = ~(n6654 ^ n3765);
assign n10023 = ~(n5251 ^ n7695);
assign n2645 = ~(n11425 ^ n6025);
assign n3435 = ~n6195;
assign n5492 = ~(n2944 | n4398);
assign n713 = n2272 | n10258;
assign n2518 = ~(n6180 ^ n3678);
assign n8216 = n752 | n7952;
assign n12334 = ~(n6347 ^ n9890);
assign n8656 = n12069 & n5645;
assign n971 = n4671 | n8300;
assign n3542 = ~(n8831 | n3918);
assign n11941 = ~n11836;
assign n67 = n4856 & n10610;
assign n1065 = n10517 & n8799;
assign n9973 = ~(n3802 ^ n8151);
assign n10100 = n1923 & n6640;
assign n9544 = ~(n456 ^ n779);
assign n3881 = ~(n3121 ^ n2436);
assign n2875 = n10745 & n12072;
assign n954 = ~(n7914 ^ n4351);
assign n5450 = n11716 | n9460;
assign n1452 = n848 | n2910;
assign n3824 = ~(n6553 ^ n11062);
assign n11586 = n12327 & n1660;
assign n7613 = ~n2890;
assign n1631 = ~(n5407 ^ n5390);
assign n6019 = ~(n1515 | n4832);
assign n6750 = n3084 & n2801;
assign n3609 = n11851 & n9255;
assign n3965 = ~n6413;
assign n3647 = n3959 & n2008;
assign n2818 = ~(n6745 ^ n2888);
assign n7148 = ~(n4098 ^ n11217);
assign n5714 = ~(n1140 ^ n10543);
assign n4832 = ~n2218;
assign n1135 = ~(n334 ^ n9156);
assign n12717 = ~(n8688 | n7086);
assign n1318 = ~(n1814 ^ n5708);
assign n1084 = ~n1217;
assign n10901 = ~(n1072 ^ n11051);
assign n6215 = ~(n2532 ^ n1880);
assign n5717 = ~(n9546 ^ n5184);
assign n10314 = ~(n5456 ^ n87);
assign n12684 = ~(n6296 ^ n10197);
assign n7239 = ~(n11136 ^ n8370);
assign n10482 = n3682 | n8958;
assign n7241 = ~(n2593 ^ n8497);
assign n7474 = n8959 | n9741;
assign n332 = n5949 & n661;
assign n11319 = ~n2411;
assign n6394 = n11805 & n8047;
assign n2857 = ~(n6036 ^ n4348);
assign n1558 = n12855 | n9717;
assign n6966 = ~(n8736 | n12526);
assign n12525 = n4628 | n1932;
assign n12073 = ~(n8225 ^ n9202);
assign n359 = ~(n11656 | n1416);
assign n10758 = ~(n8245 ^ n8464);
assign n4626 = ~(n5596 ^ n9906);
assign n1114 = ~n4897;
assign n3120 = ~n7908;
assign n2735 = n8339 | n4450;
assign n5230 = n9151 | n951;
assign n2096 = ~(n9038 ^ n7623);
assign n6845 = ~(n1585 | n11269);
assign n9869 = n5355 | n6389;
assign n8105 = ~(n8320 | n232);
assign n1415 = n3096 | n11820;
assign n2527 = ~(n4290 ^ n12634);
assign n3291 = n12935 | n9808;
assign n4286 = ~(n197 ^ n10689);
assign n553 = ~(n8077 ^ n3575);
assign n11612 = ~(n4960 ^ n4851);
assign n4088 = ~(n2485 ^ n9542);
assign n11712 = n2099 | n2964;
assign n4011 = ~(n2790 | n666);
assign n12355 = n8642 | n259;
assign n8599 = ~n7286;
assign n10222 = n11635 | n3037;
assign n12446 = ~n4094;
assign n8003 = n6542 & n8891;
assign n1307 = ~(n4087 ^ n5451);
assign n4371 = n6458 & n9204;
assign n6158 = n7157 & n6746;
assign n11981 = ~(n6643 | n9092);
assign n3478 = n5240 & n4921;
assign n2301 = ~(n1663 ^ n7833);
assign n1176 = ~(n12246 | n287);
assign n2035 = ~(n11060 ^ n11247);
assign n1985 = n3236 | n3067;
assign n9092 = n8736 & n12526;
assign n10628 = n35 & n887;
assign n12086 = n4728 & n10505;
assign n151 = ~n10790;
assign n8067 = ~n11002;
assign n5820 = n11153 & n8433;
assign n8735 = ~n615;
assign n6346 = ~(n6078 ^ n2672);
assign n2698 = ~(n9186 | n7172);
assign n11741 = n7495 | n6389;
assign n2129 = ~(n1191 ^ n9630);
assign n12339 = ~(n8945 ^ n11068);
assign n6194 = ~(n4619 ^ n9932);
assign n9397 = ~n753;
assign n3849 = ~(n1265 ^ n4293);
assign n12669 = ~n7693;
assign n12112 = n9370 | n10066;
assign n4899 = n5915 | n9586;
assign n11727 = n752 | n5311;
assign n957 = ~n10770;
assign n12960 = n12119 | n5781;
assign n6271 = n6718 | n4654;
assign n9559 = ~(n2972 | n10888);
assign n12782 = ~(n12131 | n11647);
assign n12811 = n1731 & n2068;
assign n5442 = n8778 & n12718;
assign n8026 = ~n10928;
assign n1090 = n158 & n9260;
assign n5103 = ~(n5963 ^ n4102);
assign n3177 = ~(n9355 | n2065);
assign n6530 = ~n9345;
assign n9528 = n2739 & n1033;
assign n4703 = ~(n4232 ^ n12549);
assign n9700 = n4540 | n4448;
assign n3068 = ~(n11318 ^ n8924);
assign n1902 = ~(n10507 ^ n1484);
assign n2786 = n7713 | n4012;
assign n6258 = ~(n4612 ^ n2417);
assign n11485 = n12586 | n1320;
assign n8777 = n3630 | n6831;
assign n2783 = ~(n2311 | n5206);
assign n2224 = n1494 | n7198;
assign n11626 = ~(n791 | n5226);
assign n11361 = n11327 & n599;
assign n5272 = ~(n9122 ^ n430);
assign n5593 = n2036 | n2853;
assign n4745 = ~(n5014 ^ n11938);
assign n9527 = n8515 & n10629;
assign n12922 = ~(n3519 ^ n6751);
assign n8642 = ~(n12582 | n10891);
assign n1470 = n10364 | n5156;
assign n986 = n12845 & n260;
assign n7510 = n10566 ^ n2183;
assign n2642 = n989 | n11430;
assign n1664 = n6131 | n2060;
assign n7495 = ~n12025;
assign n5263 = ~(n11388 ^ n11314);
assign n9931 = n636 | n530;
assign n28 = ~n5760;
assign n3282 = n12142 | n4458;
assign n9723 = n11538 & n8798;
assign n5543 = n6654 | n8578;
assign n4646 = n2207 & n5795;
assign n391 = ~(n6472 ^ n8457);
assign n6916 = ~(n6310 ^ n1606);
assign n9715 = ~(n12855 ^ n11989);
assign n10302 = n3007 & n8561;
assign n1974 = ~(n8986 | n10680);
assign n4368 = ~(n11986 ^ n11644);
assign n3051 = ~(n4756 | n6010);
assign n1775 = ~(n4202 ^ n9497);
assign n7313 = ~(n10098 | n4004);
assign n11457 = ~n9778;
assign n10196 = ~n5860;
assign n4932 = ~(n10475 ^ n748);
assign n5361 = n12853 | n7382;
assign n847 = ~(n9150 ^ n5308);
assign n3959 = n3746 | n9741;
assign n7987 = ~(n4457 ^ n11041);
assign n5878 = ~n6269;
assign n4361 = ~(n4601 ^ n7093);
assign n7106 = ~(n10531 ^ n670);
assign n2472 = ~n952;
assign n8633 = n10835 | n5759;
assign n2186 = ~n2992;
assign n4844 = n6365 & n6285;
assign n250 = n5353 & n1171;
assign n1139 = n3820 | n9160;
assign n7637 = n2523 & n5753;
assign n10168 = ~(n1999 | n7171);
assign n2269 = n3367 & n3056;
assign n3715 = n8564 | n12226;
assign n4181 = ~(n6148 ^ n2748);
assign n9906 = ~(n9508 ^ n146);
assign n4972 = n5355 | n5851;
assign n902 = ~(n3596 | n7345);
assign n7760 = n7271 & n11263;
assign n7155 = ~(n4286 ^ n8472);
assign n8057 = n12227 & n11940;
assign n10631 = ~(n4513 ^ n2331);
assign n7746 = ~(n2057 ^ n1431);
assign n9729 = n9373 | n9521;
assign n3666 = ~n9440;
assign n1657 = ~n8671;
assign n2174 = n161 & n550;
assign n5001 = ~(n2892 ^ n2299);
assign n8177 = ~n4949;
assign n8601 = n5593 & n2800;
assign n1008 = n6857 & n4544;
assign n9614 = n807 | n5012;
assign n12872 = n8556 & n12794;
assign n5726 = ~(n6374 ^ n2230);
assign n6508 = n2763 & n789;
assign n6532 = ~(n5420 ^ n7855);
assign n9599 = ~(n25 | n3952);
assign n1894 = ~(n7085 ^ n1725);
assign n6139 = ~(n9383 ^ n8195);
assign n4892 = n2217 | n5914;
assign n6849 = ~n2878;
assign n5347 = n12907 | n12636;
assign n5806 = ~(n1686 ^ n860);
assign n5063 = ~(n4255 ^ n9501);
assign n6603 = ~(n3133 ^ n6541);
assign n12536 = n7932 & n6065;
assign n12408 = ~(n440 | n5986);
assign n4377 = n4047 & n7770;
assign n27 = ~n6896;
assign n12254 = ~(n11801 ^ n4071);
assign n8834 = n7611 | n1296;
assign n1929 = ~n12309;
assign n4572 = ~n2177;
assign n12535 = ~n12925;
assign n3795 = n10394 & n9265;
assign n6238 = n11011 & n3869;
assign n6418 = ~n1147;
assign n11048 = n796 | n6116;
assign n20 = ~(n8474 ^ n12570);
assign n229 = ~(n10627 ^ n3656);
assign n1409 = n12119 | n10422;
assign n11514 = n2832 | n10066;
assign n10145 = ~n7052;
assign n9642 = ~n8892;
assign n6087 = ~(n3047 ^ n11403);
assign n5794 = ~(n1550 ^ n7129);
assign n4961 = n8026 | n7425;
assign n5019 = n4904 & n701;
assign n6645 = ~(n10525 ^ n1245);
assign n10339 = ~n3146;
assign n11925 = n8428 | n184;
assign n8704 = n994 | n7881;
assign n4710 = n10750 | n12754;
assign n5636 = ~(n4868 | n11379);
assign n5191 = n2342 ^ n6926;
assign n8248 = ~(n10529 | n12337);
assign n1392 = n11958 | n12899;
assign n10229 = n9043 & n10840;
assign n3632 = n12208 & n10017;
assign n11440 = ~(n3150 ^ n9127);
assign n11178 = ~(n872 ^ n230);
assign n11942 = n7705 & n11863;
assign n2892 = ~(n6668 ^ n3637);
assign n10792 = n7449 | n12771;
assign n6462 = n10987 & n5526;
assign n1924 = ~(n9530 ^ n193);
assign n6350 = ~(n7105 ^ n6716);
assign n12630 = n4059 | n10419;
assign n10918 = ~(n6342 ^ n3655);
assign n7666 = ~(n9041 ^ n6276);
assign n6442 = n4911 | n7424;
assign n8809 = n5563 ^ n4367;
assign n8846 = ~(n8555 ^ n6064);
assign n2744 = ~(n1958 ^ n5232);
assign n551 = ~(n3982 ^ n6005);
assign n6012 = ~(n10368 ^ n7269);
assign n172 = ~(n8442 | n12252);
assign n10698 = n12098 | n5499;
assign n8396 = n8458 & n3761;
assign n5618 = ~(n2153 ^ n704);
assign n5977 = ~n804;
assign n4946 = ~n12315;
assign n3127 = ~n11757;
assign n3073 = ~n3814;
assign n3528 = ~(n10235 | n3427);
assign n308 = n12119 | n6513;
assign n7580 = ~(n4374 ^ n3595);
assign n951 = ~(n695 ^ n2389);
assign n5386 = n3096 | n6169;
assign n12382 = ~(n2999 | n7484);
assign n3069 = ~(n8102 ^ n3854);
assign n2208 = n8428 | n11775;
assign n11173 = ~(n9275 ^ n8402);
assign n12322 = ~(n12211 | n3394);
assign n1303 = n12327 | n1660;
assign n12399 = n9701 & n2799;
assign n12868 = ~n9728;
assign n2314 = ~(n6305 ^ n4761);
assign n11571 = n1031 | n8378;
assign n11907 = ~n4583;
assign n7125 = ~n8091;
assign n778 = n1937 | n3421;
assign n594 = ~(n3881 ^ n10612);
assign n10153 = ~(n6911 ^ n52);
assign n8849 = ~(n9082 ^ n7944);
assign n982 = n12053 | n4464;
assign n7061 = n2268 | n3351;
assign n11814 = ~(n7694 ^ n12015);
assign n3753 = ~(n4849 ^ n963);
assign n6404 = n11681 | n2728;
assign n3390 = ~(n7737 ^ n2000);
assign n10425 = n7461 & n7892;
assign n4955 = n3221 & n3314;
assign n2394 = n1833 | n9684;
assign n7706 = n10585 | n11862;
assign n6762 = ~(n6058 ^ n10182);
assign n3526 = ~(n3036 ^ n6549);
assign n12948 = ~(n4380 ^ n5245);
assign n3499 = ~(n9072 ^ n12574);
assign n3198 = ~n868;
assign n2648 = ~(n11245 ^ n4725);
assign n4860 = ~(n2846 ^ n7904);
assign n1827 = n10478 | n4055;
assign n12257 = ~(n3003 ^ n2843);
assign n5634 = ~(n11156 ^ n11906);
assign n4537 = n8618 | n2247;
assign n4935 = ~(n7655 | n9410);
assign n1567 = ~n3753;
assign n5952 = ~(n12525 ^ n6571);
assign n1054 = ~(n5128 | n5018);
assign n5812 = n10157 | n11698;
assign n1934 = n10750 | n5468;
assign n12818 = n6261 & n6732;
assign n3582 = n8959 | n5538;
assign n3561 = n11026 | n4654;
assign n2063 = ~(n7087 | n611);
assign n1449 = n12361 | n995;
assign n4388 = ~(n3399 ^ n4328);
assign n1984 = ~(n9594 ^ n2370);
assign n2542 = n4059 | n12328;
assign n6276 = ~(n8674 ^ n5642);
assign n7283 = ~n5964;
assign n9354 = n6977 | n5540;
assign n2124 = n3746 | n11896;
assign n2647 = ~(n2661 | n9511);
assign n4775 = ~n2253;
assign n414 = ~(n3078 ^ n6032);
assign n10661 = ~n6096;
assign n6616 = n9027 | n1588;
assign n10256 = n7912 & n4136;
assign n11029 = ~n8129;
assign n1395 = n168 & n6761;
assign n11484 = ~n10747;
assign n5073 = ~(n10932 ^ n8425);
assign n8646 = n5977 & n1716;
assign n7315 = n8813 & n9401;
assign n3732 = ~(n11777 ^ n470);
assign n11139 = n9713 | n9873;
assign n7915 = ~(n9260 ^ n3981);
assign n9540 = ~(n1599 ^ n11816);
assign n11503 = n6547 & n670;
assign n187 = n12299 & n8595;
assign n5966 = n2790 & n666;
assign n5034 = ~(n6390 ^ n322);
assign n1744 = n29 | n4027;
assign n3650 = n5530 | n3924;
assign n2198 = ~(n4279 ^ n3446);
assign n8632 = n8132 & n7867;
assign n7011 = ~(n5482 | n6960);
assign n8544 = n201 & n8695;
assign n2713 = n2843 & n3578;
assign n5985 = ~n1355;
assign n10757 = ~(n3140 ^ n3447);
assign n6417 = ~n2827;
assign n95 = n8091 & n3759;
assign n11889 = ~n3054;
assign n6973 = n9921 | n10533;
assign n6910 = ~(n871 ^ n2769);
assign n9563 = ~n3420;
assign n6932 = ~(n5259 ^ n828);
assign n6327 = ~n8392;
assign n12214 = ~n8844;
assign n1944 = n6423 | n7786;
assign n1100 = n6204 & n11735;
assign n8019 = n5429 & n7702;
assign n4794 = ~(n1696 ^ n218);
assign n2701 = n4062 | n5962;
assign n5130 = ~(n8956 ^ n12922);
assign n1613 = ~(n9223 | n12179);
assign n6305 = n8687 | n4527;
assign n12345 = ~(n2296 ^ n8206);
assign n12792 = n11527 | n8072;
assign n4304 = n8204 & n3064;
assign n8383 = n4066 | n8800;
assign n10759 = n1475 & n4986;
assign n959 = n8070 & n473;
assign n7480 = n10835 | n609;
assign n4729 = n10709 | n4822;
assign n11630 = ~(n335 | n6702);
assign n4788 = n5088 & n3636;
assign n2419 = n4343 | n12535;
assign n5147 = n7495 | n1851;
assign n1658 = ~(n11966 ^ n9847);
assign n11120 = n4519 & n7109;
assign n10952 = ~n7064;
assign n6543 = n3820 | n795;
assign n7115 = ~n1016;
assign n12473 = ~(n5499 ^ n6638);
assign n12170 = ~n11971;
assign n6434 = ~(n3371 ^ n11323);
assign n11231 = ~(n3639 ^ n6499);
assign n10814 = n6373 | n12120;
assign n2203 = ~(n3875 ^ n657);
assign n5273 = ~(n8770 | n8248);
assign n4111 = ~n8475;
assign n13 = n2832 | n1162;
assign n666 = n4016 & n9314;
assign n7533 = n6864 | n451;
assign n4093 = ~(n4042 | n11666);
assign n11895 = ~(n8145 ^ n3449);
assign n9110 = n5844 & n5938;
assign n5002 = ~n4752;
assign n8932 = ~(n2319 ^ n1874);
assign n2615 = n874 | n109;
assign n7086 = ~(n1178 | n3563);
assign n9211 = n8262 & n3085;
assign n9533 = ~(n10347 ^ n12182);
assign n675 = ~(n5556 ^ n642);
assign n4007 = ~(n8068 ^ n11566);
assign n11390 = n11958 | n9741;
assign n7238 = n3324 | n4654;
assign n6272 = ~(n5266 ^ n12868);
assign n12426 = n6977 | n6169;
assign n3160 = ~n4577;
assign n7219 = ~(n3901 | n3929);
assign n10026 = ~n9603;
assign n5029 = n6600 | n2074;
assign n6644 = n4127 & n5890;
assign n7889 = n12203 | n10593;
assign n4220 = n1812 & n10855;
assign n9568 = ~n3342;
assign n10987 = n12069 & n2498;
assign n259 = n7352 & n3893;
assign n5224 = n835 & n7979;
assign n5689 = n5518 | n3990;
assign n943 = n1165 | n1640;
assign n11607 = ~(n4138 | n4587);
assign n9396 = ~(n2401 ^ n11973);
assign n750 = ~(n8936 ^ n10192);
assign n1298 = n10735 & n4091;
assign n6185 = ~n10929;
assign n4551 = ~(n895 ^ n6206);
assign n3424 = n6718 | n5258;
assign n12207 = ~(n12920 ^ n2113);
assign n1283 = ~n5895;
assign n5886 = n3735 | n2325;
assign n1587 = n3530 & n11583;
assign n6252 = n10417 | n10146;
assign n4378 = ~(n12787 ^ n2960);
assign n6682 = ~(n1420 ^ n557);
assign n1371 = n8477 & n8952;
assign n8316 = n5064 & n8974;
assign n8219 = ~(n181 | n5375);
assign n8144 = ~(n10107 ^ n6156);
assign n573 = n10142 | n7341;
assign n6121 = ~(n1973 ^ n8779);
assign n9380 = n3728 | n7740;
assign n10198 = n699 | n7085;
assign n5764 = n3757 & n10363;
assign n1481 = n827 & n3264;
assign n838 = ~(n7998 ^ n4153);
assign n1830 = n9158 & n2390;
assign n8027 = n10635 & n8078;
assign n8337 = ~n8585;
assign n11960 = n8127 | n7424;
assign n6311 = n12275 | n12086;
assign n8341 = ~(n6569 ^ n4031);
assign n6658 = ~(n961 | n9553);
assign n1592 = n2526 & n8491;
assign n2000 = ~(n11116 ^ n10050);
assign n9199 = n3992 & n12704;
assign n1396 = n6808 | n9124;
assign n11280 = n11402 & n6953;
assign n2643 = n4989 & n4764;
assign n12799 = n1051 | n11896;
assign n1669 = n3033 & n1049;
assign n12882 = n10142 | n8970;
assign n8409 = n97 & n2129;
assign n10574 = n8428 | n12899;
assign n12842 = n0 | n9322;
assign n3215 = n7116 | n7876;
assign n11401 = n12119 | n8644;
assign n4162 = ~(n2527 ^ n7257);
assign n3833 = n1333 & n2585;
assign n9998 = ~(n6407 ^ n2208);
assign n2263 = ~(n1035 ^ n2836);
assign n5280 = ~(n8758 | n12630);
assign n7285 = n11552 | n9160;
assign n8344 = n7181 & n11962;
assign n2069 = n191 | n1851;
assign n5140 = ~(n4656 ^ n1781);
assign n10682 = ~(n12923 | n5966);
assign n9692 = ~n7758;
assign n12125 = ~(n6448 ^ n7570);
assign n5448 = ~(n2365 | n9612);
assign n7341 = ~n11917;
assign n854 = n5449 & n427;
assign n1607 = n8583 | n9160;
assign n5609 = n4154 & n5746;
assign n1826 = n12119 | n4913;
assign n1351 = ~(n12316 ^ n8576);
assign n5713 = n6993 & n9915;
assign n1173 = ~(n8216 ^ n4183);
assign n5440 = ~(n9415 ^ n9968);
assign n87 = n12477 & n9178;
assign n12959 = ~(n5790 ^ n12174);
assign n4874 = n3706 & n10461;
assign n10215 = ~(n2240 ^ n6127);
assign n4800 = ~(n6151 ^ n694);
assign n6316 = n6977 | n11410;
assign n4694 = ~(n3965 | n12778);
assign n9890 = n7282 & n11604;
assign n10246 = ~(n1003 ^ n6265);
assign n10608 = ~(n2917 ^ n2426);
assign n3062 = ~n5783;
assign n3368 = n8583 | n5502;
assign n6613 = n2599 & n10681;
assign n9673 = ~(n4787 ^ n1889);
assign n11570 = ~(n132 ^ n5637);
assign n7235 = n9048 & n5993;
assign n8533 = n4059 | n7703;
assign n3187 = ~(n4339 ^ n5246);
assign n11939 = n8870 | n8109;
assign n3429 = ~n3805;
assign n5832 = n752 | n11820;
assign n6149 = n6182 & n11336;
assign n9704 = ~(n10718 | n6585);
assign n5779 = n6881 | n6489;
assign n3314 = n4059 | n8524;
assign n6632 = n5548 | n9768;
assign n9143 = ~(n6387 ^ n1487);
assign n9782 = ~n5229;
assign n4598 = ~(n6072 ^ n5473);
assign n8980 = ~(n6881 ^ n6489);
assign n9386 = ~(n10002 ^ n2587);
assign n7633 = ~n4260;
assign n9176 = ~(n10304 ^ n6928);
assign n4533 = n4951 | n11496;
assign n5412 = ~(n10137 ^ n2179);
assign n5227 = n4648 & n10473;
assign n5590 = n10479 & n6884;
assign n6301 = ~n10692;
assign n10360 = n7212 & n8772;
assign n4053 = n2456 | n8740;
assign n7953 = ~(n6562 ^ n8861);
assign n4332 = n5691 | n6338;
assign n11576 = n9335 | n11031;
assign n4515 = n9172 | n11949;
assign n7538 = n11864 | n8943;
assign n5072 = ~(n710 ^ n12851);
assign n922 = ~(n3643 | n8741);
assign n8497 = ~(n5752 ^ n5930);
assign n5626 = ~(n7688 ^ n11465);
assign n10032 = ~n3975;
assign n1735 = ~(n5146 | n11963);
assign n8460 = n3498 & n6048;
assign n9018 = ~(n7919 ^ n10756);
assign n3012 = n392 & n9940;
assign n11101 = n10842 & n5823;
assign n8725 = n10485 & n2084;
assign n739 = n5005 | n1968;
assign n12164 = n305 | n3321;
assign n10975 = ~(n1373 ^ n1074);
assign n10483 = ~(n12072 ^ n6263);
assign n12413 = n5981 | n5661;
assign n10657 = n420 & n10308;
assign n8231 = ~(n7185 ^ n2895);
assign n2561 = ~(n4124 | n11935);
assign n1440 = ~(n9161 ^ n11766);
assign n8612 = n994 | n5851;
assign n4681 = n8127 | n11746;
assign n852 = n12790 ^ n7255;
assign n12418 = ~(n2427 ^ n9801);
assign n12699 = ~n1009;
assign n5920 = ~(n10566 | n6730);
assign n11288 = n5856 | n10890;
assign n10407 = ~(n3285 ^ n5513);
assign n12494 = ~(n1575 | n6521);
assign n8372 = ~(n10820 ^ n10737);
assign n467 = n1290 | n7002;
assign n8918 = ~(n183 ^ n10638);
assign n11009 = n9588 & n3832;
assign n2043 = ~(n10681 ^ n5433);
assign n8018 = ~(n11498 ^ n5766);
assign n5471 = n1766 | n1532;
assign n2595 = n6103 & n11603;
assign n7290 = ~(n4286 | n8472);
assign n12881 = n9782 | n7875;
assign n3767 = n8552 | n3924;
assign n1893 = ~(n9342 ^ n6052);
assign n3552 = n1726 | n3718;
assign n283 = n6373 | n1509;
assign n10946 = ~(n83 ^ n30);
assign n2646 = n3875 | n9585;
assign n12812 = ~(n6095 ^ n781);
assign n4158 = ~(n11016 | n3968);
assign n7691 = ~n11702;
assign n2754 = ~n1198;
assign n8808 = ~(n1278 ^ n8796);
assign n6618 = n5767 & n9111;
assign n3059 = ~n10181;
assign n2228 = n10835 | n9280;
assign n7874 = n989 | n7881;
assign n12093 = ~n6050;
assign n4762 = ~(n6575 ^ n840);
assign n9841 = n5969 & n1313;
assign n10289 = ~(n6113 | n4646);
assign n7144 = n10157 | n5914;
assign n37 = ~(n9444 ^ n9291);
assign n9062 = ~(n3570 ^ n9972);
assign n8510 = n9370 | n1851;
assign n2313 = n8428 | n2232;
assign n5460 = n2722 & n10136;
assign n9012 = ~(n3072 ^ n4750);
assign n1343 = ~(n4591 | n1235);
assign n9204 = ~(n5624 ^ n1450);
assign n1844 = n10514 & n11187;
assign n1514 = n9368 | n809;
assign n7425 = ~n8819;
assign n8514 = n8423 | n7315;
assign n10908 = n12237 | n5326;
assign n6338 = ~(n4871 ^ n12090);
assign n8103 = n5575 | n10919;
assign n4037 = ~(n8596 ^ n1007);
assign n9321 = n10142 | n10066;
assign n9991 = n1719 | n766;
assign n7526 = ~(n11411 ^ n3856);
assign n583 = n11923 | n12120;
assign n9462 = n757 | n3707;
assign n1204 = ~(n8223 ^ n988);
assign n1628 = n3407 | n1087;
assign n422 = n5355 | n561;
assign n6990 = ~(n1306 ^ n6417);
assign n5924 = ~(n12278 | n3853);
assign n8841 = ~(n11547 ^ n6832);
assign n4130 = n3680 | n777;
assign n4574 = ~(n2471 ^ n2662);
assign n7166 = n4280 & n7970;
assign n7038 = n12047 | n3803;
assign n10764 = ~(n759 ^ n10907);
assign n241 = ~(n10309 ^ n11180);
assign n3399 = n5530 | n12441;
assign n862 = ~n6910;
assign n6277 = n8510 | n8274;
assign n9564 = ~(n10321 ^ n6617);
assign n7909 = n10142 | n5497;
assign n9006 = ~(n9627 | n833);
assign n5174 = ~(n1328 ^ n9359);
assign n5326 = ~n521;
assign n4981 = ~(n11703 ^ n7648);
assign n5881 = n9520 & n12624;
assign n2536 = n191 | n7424;
assign n10297 = n4628 | n7136;
assign n2741 = n1372 | n1873;
assign n1756 = n8055 & n3802;
assign n6208 = n11487 & n4548;
assign n10236 = n12188 & n11081;
assign n10640 = n8276 & n3602;
assign n4936 = ~n12342;
assign n9713 = ~(n3098 | n6711);
assign n3438 = n5561 | n7682;
assign n7304 = n4498 | n1162;
assign n771 = n7449 | n11698;
assign n5409 = n5858 | n10066;
assign n7475 = n374 & n10595;
assign n9175 = n10530 & n1038;
assign n5981 = n989 | n1079;
assign n2368 = n5902 | n11827;
assign n7930 = n2430 | n640;
assign n9384 = ~(n6256 ^ n7489);
assign n2602 = n7391 | n7703;
assign n846 = ~n1956;
assign n97 = n2217 | n5502;
assign n2954 = n7413 & n10998;
assign n9960 = n12562 | n8048;
assign n3129 = ~(n5995 ^ n8594);
assign n12593 = ~(n763 ^ n5979);
assign n12432 = ~(n5793 ^ n798);
assign n5599 = n35 | n887;
assign n3262 = n191 | n11430;
assign n7394 = n6373 | n9280;
assign n12089 = ~(n3255 ^ n2398);
assign n6833 = n1683 | n667;
assign n10569 = ~n4210;
assign n389 = ~n9925;
assign n3553 = n4509 & n7930;
assign n11118 = n9262 | n795;
assign n1150 = ~n4168;
assign n12853 = ~n137;
assign n7264 = n3975 | n11321;
assign n5752 = ~(n11779 ^ n2007);
assign n11900 = n1572 | n12710;
assign n11890 = n4059 | n11746;
assign n8253 = n7202 & n4103;
assign n9393 = n6750 | n8346;
assign n752 = ~n8759;
assign n12472 = ~n12343;
assign n1284 = ~n3111;
assign n3642 = ~(n8918 ^ n8764);
assign n4138 = ~n9136;
assign n2953 = n2870 & n6700;
assign n11652 = ~n1330;
assign n6095 = ~(n1940 ^ n8889);
assign n12744 = ~(n6655 ^ n5827);
assign n4923 = ~(n10989 ^ n7716);
assign n10063 = ~n2897;
assign n3366 = ~(n12066 ^ n10179);
assign n8974 = n8026 | n1413;
assign n3066 = n107 | n10880;
assign n8142 = n12539 & n4623;
assign n9842 = ~(n10841 ^ n9560);
assign n4239 = n8570 & n846;
assign n12822 = n7088 | n7214;
assign n11242 = ~(n11401 ^ n2666);
assign n40 = n12691 & n6543;
assign n12787 = ~(n152 ^ n9181);
assign n6123 = n12261 & n3190;
assign n2887 = n11538 | n8798;
assign n12280 = n12648 & n7610;
assign n3362 = n686 | n2232;
assign n808 = ~(n1886 ^ n12641);
assign n5425 = n3845 | n10733;
assign n11286 = ~(n5861 ^ n9994);
assign n12803 = n12520 | n12307;
assign n8534 = ~(n2343 ^ n8930);
assign n3981 = ~(n158 ^ n11961);
assign n4547 = n6678 | n3267;
assign n3323 = ~n8484;
assign n10003 = ~n5369;
assign n1104 = n11821 & n9956;
assign n2289 = n2677 | n9579;
assign n5630 = ~(n11997 | n9582);
assign n4148 = ~(n11895 ^ n11157);
assign n5896 = ~(n3817 | n9276);
assign n3858 = ~(n11772 ^ n941);
assign n6699 = ~(n9504 ^ n11910);
assign n11790 = ~(n325 ^ n2609);
assign n9343 = n636 | n4913;
assign n11295 = ~(n8578 ^ n571);
assign n11005 = n2456 | n5468;
assign n10591 = ~(n6606 ^ n3582);
assign n11291 = n7809 & n1095;
assign n11841 = n639 | n1669;
assign n9414 = n11829 & n4571;
assign n9721 = n9834 & n7467;
assign n990 = n7107 & n12400;
assign n9089 = n1236 & n9289;
assign n5132 = ~(n4833 ^ n10496);
assign n9404 = n9370 | n10419;
assign n6995 = n9878 | n12080;
assign n3529 = ~(n5988 | n10706);
assign n5845 = n3992 & n9763;
assign n16 = ~(n10292 ^ n11368);
assign n8167 = ~n10322;
assign n5303 = n1012 | n11537;
assign n1503 = n8127 | n1162;
assign n8531 = n962 | n9568;
assign n1618 = ~n10941;
assign n1376 = ~(n10342 | n12382);
assign n9566 = n7025 | n8234;
assign n2991 = ~(n6074 ^ n1400);
assign n12104 = ~(n10694 ^ n11012);
assign n3792 = ~(n9001 ^ n1650);
assign n10548 = n2456 | n7136;
assign n6181 = ~(n3864 | n3246);
assign n10445 = ~(n2004 ^ n11398);
assign n10538 = n7686 & n6074;
assign n11989 = ~n327;
assign n7487 = n9389 | n1079;
assign n6353 = n9400 & n10451;
assign n6743 = n9416 | n12276;
assign n12403 = ~(n6681 ^ n10894);
assign n11064 = ~(n3845 ^ n10733);
assign n5499 = n10196 | n9521;
assign n850 = n7080 & n10509;
assign n8689 = ~(n1358 ^ n12462);
assign n10466 = n12069 & n12489;
assign n664 = n3944 | n334;
assign n10972 = n2515 & n2558;
assign n4291 = n10846 & n5525;
assign n731 = ~(n9308 ^ n9562);
assign n3498 = ~n9321;
assign n361 = ~(n12684 ^ n3697);
assign n3036 = ~(n803 ^ n743);
assign n3876 = ~(n72 ^ n9675);
assign n6131 = ~(n3205 ^ n12472);
assign n12932 = ~(n3423 ^ n8948);
assign n328 = n9370 | n561;
assign n701 = ~(n12834 ^ n9992);
assign n10074 = n4480 & n7866;
assign n12431 = n9791 & n10393;
assign n12460 = ~(n7369 ^ n4867);
assign n10581 = ~n11601;
assign n11800 = n2680 & n12577;
assign n4480 = n5530 | n530;
assign n934 = n11785 | n11284;
assign n4357 = n9389 | n10419;
assign n3733 = n2665 & n5931;
assign n4386 = n5765 | n4527;
assign n2885 = n4820 | n3789;
assign n12424 = n3140 & n3447;
assign n6622 = n1788 | n11990;
assign n12677 = ~(n9027 ^ n2081);
assign n11818 = n5200 & n1010;
assign n8052 = n10750 | n2964;
assign n9383 = n9878 | n7382;
assign n4862 = n695 | n2389;
assign n8092 = ~n11380;
assign n237 = ~(n3206 | n1820);
assign n5918 = n128 & n5460;
assign n4339 = ~(n10168 | n1895);
assign n2549 = n7469 & n12465;
assign n8439 = ~(n2841 ^ n7582);
assign n10575 = n12583 | n10333;
assign n213 = n1 | n4669;
assign n11830 = n4125 | n2655;
assign n8572 = n2447 | n9150;
assign n1364 = ~(n6495 ^ n2588);
assign n10138 = ~(n8964 ^ n10120);
assign n2725 = n1111 & n11177;
assign n5245 = n11881 & n10053;
assign n7478 = ~(n9529 ^ n7950);
assign n3119 = n7157 ^ n11079;
assign n139 = n11034 | n2583;
assign n10072 = ~(n6752 | n12017);
assign n1812 = n762 | n6312;
assign n6882 = ~(n794 | n2083);
assign n10664 = ~n5603;
assign n7206 = n191 | n1162;
assign n686 = ~n4203;
assign n6379 = ~(n1655 ^ n3787);
assign n7161 = ~n8102;
assign n7615 = n2984 & n7350;
assign n6736 = ~(n9369 ^ n2952);
assign n11045 = n5690 & n1607;
assign n9019 = ~(n12139 ^ n8043);
assign n8588 = n5945 | n9741;
assign n3232 = ~(n7304 ^ n11017);
assign n9678 = ~(n182 ^ n11549);
assign n11462 = ~(n2349 ^ n4308);
assign n8805 = n3746 | n3468;
assign n2829 = n11661 | n6279;
assign n11574 = n6921 | n8812;
assign n9978 = ~n12506;
assign n12906 = n10879 | n1079;
assign n11444 = ~(n8156 | n6908);
assign n1197 = n11923 | n28;
assign n287 = n10361 & n6305;
assign n4117 = n5007 | n2377;
assign n5216 = ~(n11873 | n1758);
assign n1423 = n9652 | n9798;
assign n5972 = n5102 & n10400;
assign n9601 = ~(n6446 ^ n10660);
assign n5262 = n2491 & n3725;
assign n3799 = ~(n5796 ^ n9673);
assign n10457 = ~(n6920 ^ n1262);
assign n1630 = ~n3478;
assign n8173 = ~n7012;
assign n674 = ~n10777;
assign n9873 = ~(n4196 | n11519);
assign n3445 = n9271 | n1866;
assign n5142 = ~(n639 ^ n88);
assign n12707 = n7283 | n7246;
assign n728 = ~(n9069 ^ n5785);
assign n5996 = n1802 | n1869;
assign n12457 = ~(n3528 ^ n4944);
assign n10551 = ~(n733 ^ n682);
assign n7167 = ~n9942;
assign n12855 = ~(n4711 ^ n10822);
assign n11654 = n9140 | n3592;
assign n4934 = ~n11164;
assign n11367 = ~n10862;
assign n12596 = ~n11099;
assign n7464 = n636 | n1163;
assign n4292 = ~(n8672 ^ n4538);
assign n5149 = n12361 | n5538;
assign n4913 = ~n1512;
assign n452 = n5530 | n2259;
assign n8056 = n9380 | n1671;
assign n3517 = n5042 & n125;
assign n4786 = n12234 ^ n9814;
assign n8753 = ~n5930;
assign n4218 = n5189 ^ n8537;
assign n6 = n6577 | n5540;
assign n4431 = n11433 | n1413;
assign n5751 = ~n12370;
assign n1432 = ~n9499;
assign n2997 = ~n3559;
assign n7670 = n11931 & n10576;
assign n9039 = ~(n12284 ^ n7329);
assign n8485 = n3506 & n2724;
assign n12026 = n12585 | n1077;
assign n2049 = ~n1850;
assign n8627 = ~(n3708 ^ n11253);
assign n8922 = ~(n9611 | n6178);
assign n3915 = ~(n8321 ^ n13);
assign n4566 = ~(n9282 | n5464);
assign n5796 = ~(n5823 ^ n565);
assign n5187 = ~(n5200 ^ n12395);
assign n1647 = ~(n9806 ^ n9164);
assign n6906 = ~n11132;
assign n6280 = ~(n7018 ^ n6735);
assign n11848 = ~(n9497 | n10472);
assign n9768 = n8619 & n2746;
assign n8954 = ~n7882;
assign n379 = ~(n10973 | n3590);
assign n10155 = ~(n3087 ^ n511);
assign n4143 = n4206 & n4303;
assign n12040 = n3096 | n10903;
assign n7374 = ~(n9605 ^ n2566);
assign n3930 = n2099 | n3924;
assign n12692 = n3096 | n5540;
assign n3446 = ~(n12108 ^ n1818);
assign n3778 = ~(n11926 | n6362);
assign n10894 = n3290 & n2989;
assign n8428 = ~n9400;
assign n5914 = ~n2507;
assign n735 = n11699 | n6262;
assign n1458 = n9085 & n5071;
assign n4487 = n2618 & n1654;
assign n4541 = ~(n6891 | n8455);
assign n5428 = ~(n8762 | n12509);
assign n7450 = n7154 & n10837;
assign n471 = ~(n5589 ^ n11291);
assign n2337 = n6977 | n8768;
assign n12436 = ~(n9840 ^ n3238);
assign n8021 = n78 & n1934;
assign n2406 = ~n7285;
assign n11920 = ~(n11942 ^ n11765);
assign n6146 = n8026 | n5540;
assign n12516 = ~(n5757 ^ n5726);
assign n7310 = n10750 | n3924;
assign n4968 = ~(n7743 ^ n10967);
assign n11996 = n4515 & n6220;
assign n4155 = n2209 ^ n7039;
assign n8039 = ~(n2279 ^ n7754);
assign n11511 = ~n9883;
assign n3126 = n7449 | n8643;
assign n5790 = ~(n10573 ^ n6026);
assign n3336 = n2116 & n10426;
assign n9899 = ~(n10148 | n7996);
assign n8033 = n11719 | n1162;
assign n7539 = ~(n5264 ^ n11803);
assign n11604 = n6175 | n8316;
assign n11351 = ~(n5052 ^ n5478);
assign n4427 = n5817 & n2053;
assign n11047 = n5959 | n8534;
assign n1413 = ~n9640;
assign n9587 = ~(n4241 ^ n7699);
assign n294 = ~n6945;
assign n10728 = ~(n8343 ^ n5706);
assign n5211 = n11968 | n6;
assign n11374 = ~n12734;
assign n3447 = n994 | n7246;
assign n1083 = n2936 & n10198;
assign n9468 = n11898 | n1924;
assign n1018 = n4151 | n3840;
assign n3312 = ~(n390 ^ n2483);
assign n7073 = ~(n5714 ^ n7985);
assign n10610 = ~(n11590 ^ n2778);
assign n3171 = n2128 & n12801;
assign n509 = n6066 | n5292;
assign n9627 = ~(n3960 ^ n6775);
assign n4871 = ~(n12858 ^ n8742);
assign n8557 = n2134 & n6988;
assign n5686 = ~(n8176 | n2388);
assign n7165 = ~(n8012 ^ n9789);
assign n617 = ~(n2739 ^ n3369);
assign n7598 = n103 | n7134;
assign n9144 = ~n3754;
assign n10824 = ~(n641 | n11230);
assign n8829 = n2111 & n7841;
assign n5343 = ~(n10354 ^ n1502);
assign n3921 = ~(n4381 ^ n26);
assign n9746 = n10750 | n8259;
assign n277 = ~(n3680 ^ n8031);
assign n2614 = ~(n6740 ^ n9524);
assign n10428 = ~(n505 ^ n854);
assign n9378 = n3739 | n9722;
assign n3324 = ~n7646;
assign n12351 = ~(n2265 ^ n7026);
assign n11148 = ~(n5874 ^ n7387);
assign n9610 = ~(n10955 ^ n5648);
assign n6553 = n11958 | n6169;
assign n4916 = ~(n6128 | n8784);
assign n9391 = ~(n9473 ^ n3292);
assign n10011 = n8839 & n10927;
assign n5647 = n5203 & n9780;
assign n3411 = n4931 & n4459;
assign n965 = ~n6008;
assign n5394 = n2456 | n12080;
assign n10691 = ~n12716;
assign n9334 = ~(n8767 ^ n1974);
assign n178 = n5355 | n6524;
assign n6410 = n8108 & n101;
assign n4839 = ~n5159;
assign n4956 = n12119 | n8648;
assign n11556 = n994 | n2358;
assign n11070 = ~n5570;
assign n5312 = ~(n11500 | n11725);
assign n6265 = n12217 & n4608;
assign n7630 = ~n10005;
assign n4215 = ~n12600;
assign n6761 = n7729 | n2303;
assign n10525 = n5249 & n10356;
assign n3037 = ~(n12937 | n2339);
assign n7519 = n2336 & n3775;
assign n363 = ~(n8224 ^ n6397);
assign n10684 = n7097 | n9115;
assign n559 = ~(n1015 ^ n10240);
assign n8731 = n1665 & n10889;
assign n8070 = n10157 | n5258;
assign n9336 = ~(n2565 | n1322);
assign n1824 = n1929 | n2485;
assign n12897 = ~(n9448 ^ n10248);
assign n9365 = ~(n57 ^ n9099);
assign n10171 = n5915 | n1163;
assign n2239 = ~(n9788 ^ n362);
assign n3781 = ~n5166;
assign n10039 = ~(n10812 | n5744);
assign n3313 = n8611 & n9015;
assign n9903 = ~(n9177 ^ n9386);
assign n8488 = ~n11354;
assign n12259 = ~(n8492 ^ n5296);
assign n2245 = n5942 | n8925;
assign n1273 = ~(n9688 ^ n8446);
assign n12608 = ~(n7957 ^ n9592);
assign n10390 = ~n6629;
assign n9562 = n11722 & n10186;
assign n1304 = ~(n3851 ^ n11091);
assign n8192 = n7287 & n8860;
assign n6320 = n5720 & n6565;
assign n7435 = ~n6583;
assign n11313 = n8197 | n1098;
assign n6876 = n3768 | n1611;
assign n2937 = n1229 & n6905;
assign n8161 = ~(n10233 | n1965);
assign n421 = n9893 | n2553;
assign n3444 = ~(n11440 ^ n8128);
assign n9474 = n6059 | n8862;
assign n3567 = n2124 & n3553;
assign n11152 = n3612 | n12676;
assign n5464 = ~(n8915 | n3956);
assign n8992 = ~(n7126 ^ n5154);
assign n8291 = n3126 | n188;
assign n5294 = ~(n9435 ^ n7535);
assign n12805 = n6028 & n9435;
assign n8164 = n2866 | n4742;
assign n6675 = ~(n1992 | n12212);
assign n3245 = ~(n9301 ^ n12244);
assign n12083 = n1083 | n6613;
assign n2939 = ~(n5559 ^ n9735);
assign n10325 = n1444 & n3951;
assign n11733 = ~n5450;
assign n10239 = n2400 | n2705;
assign n12952 = n7298 & n1325;
assign n153 = ~(n2385 ^ n8884);
assign n11799 = n5679 | n2963;
assign n3660 = ~n9242;
assign n4210 = ~(n10138 ^ n7773);
assign n627 = n8535 & n2410;
assign n3010 = ~(n1461 | n3374);
assign n10885 = ~(n12766 | n4704);
assign n9191 = ~n5276;
assign n11516 = ~(n8994 | n3041);
assign n8126 = ~(n785 | n3177);
assign n5256 = ~(n11130 ^ n3871);
assign n7922 = n9400 & n6703;
assign n5054 = ~n4010;
assign n4335 = n7004 | n3319;
assign n10707 = ~(n11266 ^ n8286);
assign n10837 = ~(n6096 ^ n9191);
assign n65 = ~(n2388 ^ n10264);
assign n12647 = n10951 | n9916;
assign n2411 = ~(n7114 ^ n44);
assign n11954 = ~(n3931 ^ n8047);
assign n10380 = ~(n12302 ^ n2462);
assign n4222 = n11759 | n6154;
assign n817 = n7391 | n11827;
assign n930 = ~(n3350 ^ n10262);
assign n9362 = ~(n6198 ^ n12567);
assign n787 = ~(n9689 ^ n7040);
assign n9418 = ~(n9364 | n1458);
assign n8939 = n2660 ^ n12812;
assign n8230 = n7378 | n5188;
assign n12532 = n1941 | n7425;
assign n11424 = n7192 | n7696;
assign n598 = ~(n343 ^ n4062);
assign n12006 = n7495 | n1079;
assign n3919 = n1937 | n1413;
assign n7049 = ~(n2560 | n6965);
assign n10984 = ~(n7870 ^ n2341);
assign n502 = n8287 | n1196;
assign n4706 = n11743 & n12004;
assign n2284 = n6977 | n7395;
assign n1921 = ~(n12281 ^ n4939);
assign n6014 = n1177 ^ n1645;
assign n619 = ~n147;
assign n2501 = ~(n910 ^ n9852);
assign n1766 = n9373 | n9160;
assign n8885 = n12813 & n946;
assign n11415 = n3746 | n6197;
assign n7280 = ~(n7225 ^ n5070);
assign n4633 = n5168 | n8997;
assign n3638 = ~n3509;
assign n2456 = ~n11478;
assign n12204 = ~(n8126 ^ n2692);
assign n3431 = n8026 | n2232;
assign n8416 = n1699 | n3924;
assign n11713 = ~(n5843 | n10236);
assign n623 = ~(n4368 ^ n7543);
assign n11965 = n714 | n3537;
assign n8923 = n5219 & n4926;
assign n4114 = ~(n10165 ^ n2276);
assign n8895 = n10683 | n2527;
assign n12645 = ~(n5290 ^ n11551);
assign n8661 = ~(n10852 ^ n11134);
assign n4041 = n6577 | n1413;
assign n5540 = ~n7500;
assign n7438 = n10717 | n7042;
assign n11932 = ~(n6473 ^ n1194);
assign n2494 = ~(n140 | n9737);
assign n2596 = n12366 | n1366;
assign n8597 = n5024 | n2044;
assign n981 = ~n1629;
assign n9611 = n1834 & n11175;
assign n12752 = n12525 | n3298;
assign n2444 = ~(n10361 | n6305);
assign n10260 = ~(n163 | n1093);
assign n7460 = ~(n1821 ^ n391);
assign n12232 = ~(n3430 ^ n579);
assign n645 = n6847 & n11002;
assign n8171 = ~n6706;
assign n3469 = n7495 | n11746;
assign n7350 = ~(n1460 ^ n12415);
assign n8162 = n12712 & n9872;
assign n2608 = n10835 | n6922;
assign n11911 = n4283 & n5524;
assign n7792 = n7839 | n7876;
assign n4549 = n2877 | n572;
assign n11318 = n3743 | n5086;
assign n2136 = n10157 | n1047;
assign n7010 = n7654 | n4482;
assign n11339 = ~(n12386 ^ n9257);
assign n797 = ~(n12557 ^ n1270);
assign n1336 = ~(n12846 ^ n7514);
assign n5128 = ~(n5688 ^ n10758);
assign n3955 = n1805 | n7072;
assign n12566 = ~(n4281 | n10380);
assign n5417 = n4717 & n12302;
assign n10721 = n3141 | n4721;
assign n1309 = n9878 | n6513;
assign n12101 = ~(n3959 ^ n2008);
assign n5049 = n10142 | n9397;
assign n7685 = n12069 & n12925;
assign n8747 = ~(n1445 ^ n3815);
assign n2325 = ~n4597;
assign n31 = ~(n7469 ^ n6723);
assign n9767 = ~(n12420 ^ n4309);
assign n11881 = n11221 | n3260;
assign n9223 = n5915 | n7928;
assign n4051 = ~n5900;
assign n3430 = ~(n10936 ^ n3631);
assign n9231 = ~(n8803 ^ n12304);
assign n7582 = ~(n7945 | n12927);
assign n4455 = ~(n10338 ^ n6123);
assign n2495 = ~(n9951 ^ n1649);
assign n12726 = ~(n5278 | n922);
assign n659 = ~(n6157 | n3657);
assign n12463 = ~(n12505 ^ n4196);
assign n939 = ~(n2222 ^ n8638);
assign n12367 = ~n312;
assign n7470 = ~n7248;
assign n6744 = n386 & n9354;
assign n11582 = n5196 | n8731;
assign n716 = ~(n12548 ^ n980);
assign n8473 = ~(n7694 | n12015);
assign n8287 = ~(n951 ^ n9151);
assign n605 = n8389 & n11484;
assign n1918 = n4250 & n7101;
assign n3104 = n8261 | n12473;
assign n11754 = n12764 & n4834;
assign n4160 = n3617 | n8109;
assign n1051 = ~n8276;
assign n1550 = ~(n10504 ^ n6682);
assign n7593 = n11142 | n10187;
assign n11783 = n6463 & n12738;
assign n7133 = n2099 | n1932;
assign n2059 = n12103 | n9593;
assign n6620 = ~(n2835 ^ n4033);
assign n6456 = ~n4732;
assign n4412 = ~(n3222 ^ n12228);
assign n1017 = ~(n10976 ^ n4526);
assign n3028 = ~n7486;
assign n7017 = ~(n4161 ^ n4888);
assign n3057 = n2312 & n3899;
assign n12103 = n8818 & n6967;
assign n5939 = ~(n5947 | n9539);
assign n8134 = n10678 & n6703;
assign n10491 = ~(n4879 ^ n4157);
assign n7579 = n3918 ^ n4922;
assign n58 = n11958 | n7952;
assign n12217 = n4536 | n4220;
assign n12619 = n21 & n10600;
assign n3137 = n5269 & n12488;
assign n3654 = ~(n1570 ^ n4680);
assign n8078 = ~n11482;
assign n3634 = n8733 & n5632;
assign n2297 = ~n4490;
assign n1462 = n191 | n561;
assign n318 = n11923 | n4654;
assign n2610 = n994 | n8524;
assign n5154 = n114 | n5540;
assign n5892 = ~(n9107 ^ n2986);
assign n10178 = n2099 | n5468;
assign n6086 = n636 | n4818;
assign n5655 = ~n4908;
assign n10763 = n1665 | n10889;
assign n3790 = ~(n7094 ^ n3900);
assign n1689 = n12237 | n8740;
assign n12248 = ~(n9869 ^ n11852);
assign n11765 = ~(n5213 ^ n6533);
assign n12587 = ~n7827;
assign n914 = ~(n8580 | n12078);
assign n2906 = n636 | n12535;
assign n7492 = n7014 & n5176;
assign n6671 = ~n10976;
assign n12440 = n1937 | n11410;
assign n5089 = n2099 | n12080;
assign n6040 = n1988 & n10674;
assign n2837 = n12119 | n12124;
assign n4115 = n357 & n5306;
assign n2661 = n5954 & n7486;
assign n5891 = n5861 | n9506;
assign n1313 = n10339 | n3224;
assign n8583 = ~n996;
assign n10021 = n616 & n2258;
assign n6180 = n5765 | n5914;
assign n9522 = n114 | n12816;
assign n6513 = ~n12489;
assign n3667 = n9389 | n10066;
assign n3096 = ~n1094;
assign n1761 = ~n2235;
assign n5145 = n3959 | n2008;
assign n9425 = n9301 & n2028;
assign n5785 = ~(n3535 ^ n11795);
assign n3742 = n12648 & n11922;
assign n2926 = ~(n6924 ^ n12527);
assign n6573 = ~(n12264 ^ n11385);
assign n420 = n10142 | n510;
assign n2992 = n8782 & n4555;
assign n12206 = ~(n4972 ^ n12167);
assign n7485 = n10625 | n11701;
assign n10241 = n413 & n7955;
assign n10976 = n6255 & n11481;
assign n11180 = n509 & n10385;
assign n6267 = n2036 & n2853;
assign n3576 = ~(n12592 ^ n10428);
assign n3845 = n8959 | n995;
assign n2755 = ~(n5730 ^ n4428);
assign n8568 = ~(n9496 ^ n1775);
assign n2266 = ~(n2104 | n7321);
assign n3588 = n7388 & n10990;
assign n7749 = n8397 & n9700;
assign n2868 = ~(n6759 | n3694);
assign n7845 = n385 & n6108;
assign n714 = n5963 & n4102;
assign n4664 = n1822 & n8375;
assign n12711 = ~n9712;
assign n11898 = n6486 & n1464;
assign n9118 = ~(n11192 | n1901);
assign n10524 = ~(n8015 ^ n11946);
assign n3464 = n752 | n6114;
assign n10969 = n7053 | n7346;
assign n121 = ~(n11515 ^ n8271);
assign n8072 = n2018 & n10383;
assign n1951 = n12560 | n6040;
assign n1805 = n8313 & n879;
assign n5363 = n2393 & n2749;
assign n631 = ~(n7846 | n4955);
assign n624 = n8988 & n8804;
assign n11699 = n8836 & n3941;
assign n9429 = n5974 & n4471;
assign n568 = ~n5053;
assign n11186 = n2626 & n4041;
assign n1554 = ~n11747;
assign n4026 = n5023 & n4063;
assign n9461 = ~(n927 | n2180);
assign n1869 = n10601 & n3576;
assign n4214 = n11144 | n2139;
assign n3179 = n11222 & n8433;
assign n10322 = ~(n1365 ^ n7787);
assign n776 = ~(n1449 ^ n1174);
assign n1143 = n8687 | n12771;
assign n6152 = n8405 | n826;
assign n1219 = ~(n3133 | n10313);
assign n371 = ~n11370;
assign n10478 = ~n1999;
assign n7044 = n9240 | n11264;
assign n12393 = ~(n5185 | n5410);
assign n7529 = ~(n97 ^ n3891);
assign n222 = n6347 | n9890;
assign n3136 = ~(n3298 ^ n5952);
assign n6018 = ~(n697 ^ n1295);
assign n5674 = n8757 | n3021;
assign n9671 = ~n5972;
assign n1665 = ~(n8533 ^ n6193);
assign n12076 = ~(n8958 ^ n1551);
assign n3346 = n1129 & n4967;
assign n8941 = ~(n8694 ^ n2582);
assign n5680 = ~n12242;
assign n11513 = ~(n4213 ^ n986);
assign n7662 = n11923 | n3606;
assign n6380 = ~(n6150 | n5921);
assign n9561 = ~n7146;
assign n6816 = n11007 & n1253;
assign n7858 = n11623 | n7632;
assign n10230 = ~(n12906 ^ n9889);
assign n10244 = ~n2990;
assign n12039 = ~n10051;
assign n11453 = n4759 & n1569;
assign n8518 = ~n2244;
assign n4008 = ~(n3712 ^ n10986);
assign n7675 = ~(n12872 | n10586);
assign n3247 = n11085 & n486;
assign n7025 = ~(n12493 | n3785);
assign n11617 = ~(n10863 ^ n4245);
assign n1543 = n1399 & n965;
assign n293 = ~(n5101 ^ n1178);
assign n4985 = n3623 | n8591;
assign n3694 = ~n10805;
assign n6778 = ~(n6590 ^ n11930);
assign n6593 = ~(n1682 ^ n9303);
assign n4171 = ~(n3444 ^ n1692);
assign n6519 = n7391 | n6402;
assign n12496 = n238 | n1813;
assign n11155 = ~(n9556 ^ n3043);
assign n8767 = ~(n11436 | n8632);
assign n10807 = ~(n4116 ^ n3310);
assign n12163 = n4187 & n11728;
assign n1571 = n8201 & n3922;
assign n9813 = ~n1493;
assign n6091 = ~n10012;
assign n7258 = n10587 | n10140;
assign n10150 = n11138 & n10218;
assign n9971 = ~n10217;
assign n6090 = n11923 | n795;
assign n2312 = n9373 | n1047;
assign n4301 = n4911 | n1079;
assign n249 = n7747 & n6311;
assign n9099 = n3940 & n9740;
assign n6466 = n3324 | n2020;
assign n2131 = ~(n6848 ^ n12077);
assign n8616 = ~(n10141 ^ n2223);
assign n12037 = ~(n10366 ^ n11185);
assign n2439 = n3618 & n3793;
assign n758 = ~(n7234 ^ n9234);
assign n6374 = n191 | n7389;
assign n2346 = n5199 | n3121;
assign n4865 = ~(n9403 | n11100);
assign n12395 = n970 & n2165;
assign n9698 = n8870 | n4818;
assign n7471 = n3220 & n9239;
assign n407 = ~(n10646 ^ n10375);
assign n6057 = ~n12463;
assign n9290 = n7283 | n8859;
assign n4742 = n6491 & n4169;
assign n2304 = ~(n12289 ^ n9253);
assign n6957 = ~n3346;
assign n2850 = n5456 & n87;
assign n3196 = ~(n11807 ^ n6092);
assign n8913 = ~(n6799 ^ n4772);
assign n11952 = ~n9828;
assign n9896 = n7862 & n5212;
assign n5100 = ~(n2435 ^ n10995);
assign n1765 = n8671 & n9485;
assign n9098 = n6554 & n5201;
assign n12161 = ~(n5794 ^ n4340);
assign n6216 = n8428 | n9971;
assign n8699 = ~n8027;
assign n11670 = n5601 | n8237;
assign n11018 = ~n8134;
assign n4552 = n7750 & n8004;
assign n736 = n779 | n456;
assign n11578 = n7495 | n7881;
endmodule
