module top( 2_n45 , 2_n112 , 2_n137 , 2_n159 , 2_n217 , 2_n226 , 2_n381 , 2_n397 , 2_n405 , 2_n447 , 2_n503 , 2_n521 , 2_n533 , 2_n615 , 2_n658 , 2_n671 , 2_n753 , 2_n783 , 2_n806 , 2_n837 , 2_n844 , 2_n911 , 2_n992 , 2_n996 , 2_n1020 , 2_n1067 , 2_n1094 , 2_n1097 , 2_n1136 , 2_n1138 , 2_n1198 , 2_n1199 , 2_n1209 , 2_n1269 , 2_n1333 , 2_n1353 , 2_n1357 , 2_n1471 , 2_n1478 , 2_n1510 , 2_n1512 , 2_n1523 , 2_n1564 , 2_n1576 , 2_n1658 , 2_n1798 , 2_n1835 , 2_n1847 , 2_n1906 , 2_n1980 , 2_n2024 , 2_n2087 , 2_n2096 , 2_n2131 , 2_n2226 , 2_n2253 , 2_n2278 , 2_n2301 , 2_n2316 , 2_n2347 , 2_n2383 , 2_n2393 , 2_n2425 , 2_n2431 , 2_n2433 , 2_n2434 , 2_n2464 , 2_n2498 , 2_n2507 , 2_n2508 , 2_n2509 , 2_n2512 , 2_n2515 , 2_n2522 , 2_n2530 , 2_n2551 , 2_n2558 , 2_n2564 , 2_n2577 , 2_n2581 , 2_n2585 , 2_n2624 , 2_n2679 , 2_n2708 , 2_n2749 , 2_n2802 , 2_n2818 , 2_n2879 , 2_n2902 , 2_n3022 , 2_n3071 , 2_n3124 , 2_n3146 , 2_n3172 , 2_n3214 , 2_n3230 , 2_n3272 , 2_n3287 , 2_n3339 , 2_n3342 , 2_n3456 , 2_n3602 , 2_n3616 , 2_n3627 , 2_n3654 , 2_n3661 , 2_n3677 , 2_n3719 , 2_n3754 , 2_n3842 , 2_n3849 , 2_n3865 , 2_n3932 , 2_n3986 , 2_n3992 , 2_n4005 , 2_n4086 , 2_n4088 , 2_n4094 , 2_n4141 , 2_n4155 , 2_n4159 , 2_n4187 , 2_n4189 , 2_n4190 , 2_n4203 , 2_n4226 , 2_n4230 , 2_n4300 , 2_n4312 , 2_n4326 , 2_n4333 , 2_n4370 , 2_n4378 , 2_n4397 , 2_n4436 , 2_n4499 , 2_n4516 , 2_n4553 , 2_n4634 , 2_n4686 , 2_n4689 , 2_n4722 , 2_n4733 , 2_n4757 , 2_n4805 , 2_n4817 , 2_n4826 , 2_n4828 , 2_n4903 , 2_n4921 , 2_n4928 , 2_n4938 , 2_n4970 , 2_n4971 , 2_n5030 , 2_n5034 , 2_n5069 , 2_n5094 , 2_n5105 , 2_n5132 , 2_n5153 , 2_n5191 , 2_n5198 , 2_n5212 , 2_n5240 , 2_n5257 , 2_n5283 , 2_n5305 , 2_n5314 , 2_n5319 , 2_n5320 , 2_n5331 , 2_n5411 , 2_n5435 , 2_n5579 , 2_n5641 , 2_n5645 , 2_n5670 , 2_n5693 , 2_n5694 , 2_n5760 , 2_n5767 , 2_n5798 , 2_n5814 , 2_n5857 , 2_n5860 , 2_n5934 , 2_n5964 , 2_n6016 , 2_n6038 , 2_n6089 , 2_n6126 , 2_n6192 , 2_n6254 , 2_n6273 , 2_n6294 , 2_n6358 , 2_n6359 , 2_n6429 , 2_n6431 , 2_n6441 , 2_n6445 , 2_n6578 , 2_n6604 , 2_n6611 , 2_n6645 , 2_n6687 , 2_n6689 , 2_n6703 , 2_n6742 , 2_n6770 , 2_n6776 , 2_n6797 , 2_n6806 , 2_n6809 , 2_n6822 , 2_n6826 , 2_n6860 , 2_n6877 , 2_n6986 , 2_n7159 , 2_n7160 , 2_n7193 , 2_n7236 , 2_n7265 , 2_n7270 , 2_n7294 , 2_n7320 , 2_n7354 , 2_n7388 , 2_n7436 , 2_n7456 , 2_n7500 , 2_n7523 , 2_n7546 , 2_n7568 , 2_n7610 , 2_n7646 , 2_n7676 , 2_n7690 , 2_n7730 , 2_n7733 , 2_n7823 , 2_n7862 , 2_n7891 , 2_n7946 , 2_n7965 , 2_n7966 , 2_n7981 , 2_n8028 , 2_n8065 , 2_n8100 , 2_n8138 , 2_n8202 , 2_n8236 , 2_n8276 , 2_n8303 , 2_n8336 , 2_n8384 , 2_n8398 , 2_n8433 , 2_n8476 , 2_n8595 , 2_n8665 , 2_n8717 , 2_n8759 , 2_n8819 , 2_n9080 , 2_n9111 , 2_n9137 , 2_n9189 , 2_n9195 , 2_n9241 , 2_n9387 , 2_n9400 , 2_n9457 , 2_n9571 , 2_n9578 , 2_n9583 , 2_n9637 , 2_n9640 , 2_n9706 , 2_n9725 , 2_n9756 , 2_n9763 , 2_n9767 , 2_n9820 , 2_n9920 , 2_n9938 , 2_n9956 , 2_n10022 , 2_n10174 , 2_n10217 , 2_n10223 , 2_n10278 , 2_n10327 , 2_n10391 , 2_n10439 , 2_n10451 , 2_n10476 , 2_n10510 , 2_n10545 , 2_n10547 , 2_n10589 , 2_n10644 , 2_n10678 , 2_n10685 , 2_n10695 , 2_n10789 , 2_n10848 , 2_n10851 , 2_n10898 , 2_n10913 , 2_n10928 , 2_n10949 , 2_n10965 , 2_n10990 , 2_n11023 , 2_n11153 , 2_n11216 , 2_n11222 , 2_n11257 , 2_n11296 , 2_n11311 , 2_n11326 , 2_n11407 , 2_n11423 , 2_n11478 , 2_n11536 , 2_n11662 , 2_n11707 , 2_n11728 , 2_n11755 , 2_n11757 , 2_n11780 , 2_n11791 , 2_n11821 , 2_n11876 , 2_n11877 , 2_n11892 , 2_n11917 , 2_n11919 , 2_n11922 , 2_n11967 , 2_n11999 , 2_n12000 , 2_n12005 , 2_n12014 , 2_n12020 , 2_n12025 , 2_n12044 , 2_n12069 , 2_n12076 , 2_n12111 , 2_n12145 , 2_n12221 , 2_n12247 , 2_n12299 , 2_n12391 , 2_n12444 , 2_n12489 , 2_n12511 , 2_n12591 , 2_n12648 , 2_n12704 , 2_n12705 , 2_n12706 , 2_n12709 , 2_n12720 , 2_n12753 , 2_n12777 , 2_n12807 , 2_n12826 , 2_n12925 , 2_n12947 );
    input 2_n45 , 2_n137 , 2_n159 , 2_n217 , 2_n405 , 2_n447 , 2_n503 , 2_n521 , 2_n533 , 2_n615 , 2_n753 , 2_n783 , 2_n806 , 2_n996 , 2_n1067 , 2_n1094 , 2_n1097 , 2_n1198 , 2_n1199 , 2_n1209 , 2_n1333 , 2_n1353 , 2_n1357 , 2_n1471 , 2_n1478 , 2_n1510 , 2_n1512 , 2_n1564 , 2_n1576 , 2_n1798 , 2_n1835 , 2_n1906 , 2_n1980 , 2_n2024 , 2_n2087 , 2_n2226 , 2_n2253 , 2_n2278 , 2_n2347 , 2_n2393 , 2_n2433 , 2_n2464 , 2_n2498 , 2_n2507 , 2_n2508 , 2_n2509 , 2_n2512 , 2_n2515 , 2_n2522 , 2_n2530 , 2_n2551 , 2_n2558 , 2_n2564 , 2_n2577 , 2_n2585 , 2_n2749 , 2_n2802 , 2_n2879 , 2_n3022 , 2_n3146 , 2_n3172 , 2_n3342 , 2_n3602 , 2_n3616 , 2_n3627 , 2_n3719 , 2_n3754 , 2_n3842 , 2_n3865 , 2_n3932 , 2_n3986 , 2_n3992 , 2_n4005 , 2_n4086 , 2_n4094 , 2_n4141 , 2_n4187 , 2_n4189 , 2_n4190 , 2_n4203 , 2_n4312 , 2_n4370 , 2_n4436 , 2_n4499 , 2_n4516 , 2_n4634 , 2_n4722 , 2_n4805 , 2_n4817 , 2_n4826 , 2_n4828 , 2_n4903 , 2_n4921 , 2_n4928 , 2_n4938 , 2_n4970 , 2_n5069 , 2_n5105 , 2_n5153 , 2_n5198 , 2_n5212 , 2_n5240 , 2_n5283 , 2_n5305 , 2_n5314 , 2_n5319 , 2_n5320 , 2_n5331 , 2_n5579 , 2_n5645 , 2_n5694 , 2_n5760 , 2_n5767 , 2_n5798 , 2_n5814 , 2_n5857 , 2_n5860 , 2_n5964 , 2_n6016 , 2_n6038 , 2_n6126 , 2_n6254 , 2_n6294 , 2_n6358 , 2_n6359 , 2_n6429 , 2_n6431 , 2_n6441 , 2_n6578 , 2_n6604 , 2_n6611 , 2_n6687 , 2_n6703 , 2_n6770 , 2_n6776 , 2_n6797 , 2_n6806 , 2_n6826 , 2_n6877 , 2_n6986 , 2_n7159 , 2_n7160 , 2_n7236 , 2_n7265 , 2_n7270 , 2_n7294 , 2_n7320 , 2_n7354 , 2_n7388 , 2_n7436 , 2_n7456 , 2_n7500 , 2_n7523 , 2_n7546 , 2_n7610 , 2_n7646 , 2_n7690 , 2_n7730 , 2_n7733 , 2_n7823 , 2_n7862 , 2_n7891 , 2_n7946 , 2_n7965 , 2_n8028 , 2_n8065 , 2_n8236 , 2_n8276 , 2_n8336 , 2_n8384 , 2_n8433 , 2_n8476 , 2_n8595 , 2_n8665 , 2_n8717 , 2_n8759 , 2_n8819 , 2_n9080 , 2_n9111 , 2_n9189 , 2_n9195 , 2_n9241 , 2_n9400 , 2_n9457 , 2_n9583 , 2_n9637 , 2_n9640 , 2_n9725 , 2_n9763 , 2_n9920 , 2_n9956 , 2_n10022 , 2_n10174 , 2_n10217 , 2_n10223 , 2_n10278 , 2_n10327 , 2_n10391 , 2_n10439 , 2_n10451 , 2_n10510 , 2_n10545 , 2_n10547 , 2_n10644 , 2_n10678 , 2_n10685 , 2_n10848 , 2_n10898 , 2_n10928 , 2_n10965 , 2_n10990 , 2_n11023 , 2_n11153 , 2_n11222 , 2_n11257 , 2_n11296 , 2_n11311 , 2_n11407 , 2_n11423 , 2_n11478 , 2_n11536 , 2_n11662 , 2_n11728 , 2_n11757 , 2_n11791 , 2_n11821 , 2_n11876 , 2_n11877 , 2_n11892 , 2_n11917 , 2_n11922 , 2_n11967 , 2_n11999 , 2_n12000 , 2_n12025 , 2_n12044 , 2_n12069 , 2_n12145 , 2_n12221 , 2_n12247 , 2_n12299 , 2_n12391 , 2_n12489 , 2_n12511 , 2_n12591 , 2_n12648 , 2_n12704 , 2_n12705 , 2_n12706 , 2_n12709 , 2_n12720 , 2_n12753 , 2_n12777 , 2_n12826 , 2_n12925 , 2_n12947 ;
    output 2_n112 , 2_n226 , 2_n381 , 2_n397 , 2_n658 , 2_n671 , 2_n837 , 2_n844 , 2_n911 , 2_n992 , 2_n1020 , 2_n1136 , 2_n1138 , 2_n1269 , 2_n1523 , 2_n1658 , 2_n1847 , 2_n2096 , 2_n2131 , 2_n2301 , 2_n2316 , 2_n2383 , 2_n2425 , 2_n2431 , 2_n2434 , 2_n2581 , 2_n2624 , 2_n2679 , 2_n2708 , 2_n2818 , 2_n2902 , 2_n3071 , 2_n3124 , 2_n3214 , 2_n3230 , 2_n3272 , 2_n3287 , 2_n3339 , 2_n3456 , 2_n3654 , 2_n3661 , 2_n3677 , 2_n3849 , 2_n4088 , 2_n4155 , 2_n4159 , 2_n4226 , 2_n4230 , 2_n4300 , 2_n4326 , 2_n4333 , 2_n4378 , 2_n4397 , 2_n4553 , 2_n4686 , 2_n4689 , 2_n4733 , 2_n4757 , 2_n4971 , 2_n5030 , 2_n5034 , 2_n5094 , 2_n5132 , 2_n5191 , 2_n5257 , 2_n5411 , 2_n5435 , 2_n5641 , 2_n5670 , 2_n5693 , 2_n5934 , 2_n6089 , 2_n6192 , 2_n6273 , 2_n6445 , 2_n6645 , 2_n6689 , 2_n6742 , 2_n6809 , 2_n6822 , 2_n6860 , 2_n7193 , 2_n7568 , 2_n7676 , 2_n7966 , 2_n7981 , 2_n8100 , 2_n8138 , 2_n8202 , 2_n8303 , 2_n8398 , 2_n9137 , 2_n9387 , 2_n9571 , 2_n9578 , 2_n9706 , 2_n9756 , 2_n9767 , 2_n9820 , 2_n9938 , 2_n10476 , 2_n10589 , 2_n10695 , 2_n10789 , 2_n10851 , 2_n10913 , 2_n10949 , 2_n11216 , 2_n11326 , 2_n11707 , 2_n11755 , 2_n11780 , 2_n11919 , 2_n12005 , 2_n12014 , 2_n12020 , 2_n12076 , 2_n12111 , 2_n12444 , 2_n12807 ;
    wire 2_n0 , 2_n1 , 2_n2 , 2_n3 , 2_n4 , 2_n5 , 2_n6 , 2_n7 , 2_n8 , 2_n9 , 2_n10 , 2_n11 , 2_n12 , 2_n13 , 2_n14 , 2_n15 , 2_n16 , 2_n17 , 2_n18 , 2_n19 , 2_n20 , 2_n21 , 2_n22 , 2_n23 , 2_n24 , 2_n25 , 2_n26 , 2_n27 , 2_n28 , 2_n29 , 2_n30 , 2_n31 , 2_n32 , 2_n33 , 2_n34 , 2_n35 , 2_n36 , 2_n37 , 2_n38 , 2_n39 , 2_n40 , 2_n41 , 2_n42 , 2_n43 , 2_n44 , 2_n46 , 2_n47 , 2_n48 , 2_n49 , 2_n50 , 2_n51 , 2_n52 , 2_n53 , 2_n54 , 2_n55 , 2_n56 , 2_n57 , 2_n58 , 2_n59 , 2_n60 , 2_n61 , 2_n62 , 2_n63 , 2_n64 , 2_n65 , 2_n66 , 2_n67 , 2_n68 , 2_n69 , 2_n70 , 2_n71 , 2_n72 , 2_n73 , 2_n74 , 2_n75 , 2_n76 , 2_n77 , 2_n78 , 2_n79 , 2_n80 , 2_n81 , 2_n82 , 2_n83 , 2_n84 , 2_n85 , 2_n86 , 2_n87 , 2_n88 , 2_n89 , 2_n90 , 2_n91 , 2_n92 , 2_n93 , 2_n94 , 2_n95 , 2_n96 , 2_n97 , 2_n98 , 2_n99 , 2_n100 , 2_n101 , 2_n102 , 2_n103 , 2_n104 , 2_n105 , 2_n106 , 2_n107 , 2_n108 , 2_n109 , 2_n110 , 2_n111 , 2_n113 , 2_n114 , 2_n115 , 2_n116 , 2_n117 , 2_n118 , 2_n119 , 2_n120 , 2_n121 , 2_n122 , 2_n123 , 2_n124 , 2_n125 , 2_n126 , 2_n127 , 2_n128 , 2_n129 , 2_n130 , 2_n131 , 2_n132 , 2_n133 , 2_n134 , 2_n135 , 2_n136 , 2_n138 , 2_n139 , 2_n140 , 2_n141 , 2_n142 , 2_n143 , 2_n144 , 2_n145 , 2_n146 , 2_n147 , 2_n148 , 2_n149 , 2_n150 , 2_n151 , 2_n152 , 2_n153 , 2_n154 , 2_n155 , 2_n156 , 2_n157 , 2_n158 , 2_n160 , 2_n161 , 2_n162 , 2_n163 , 2_n164 , 2_n165 , 2_n166 , 2_n167 , 2_n168 , 2_n169 , 2_n170 , 2_n171 , 2_n172 , 2_n173 , 2_n174 , 2_n175 , 2_n176 , 2_n177 , 2_n178 , 2_n179 , 2_n180 , 2_n181 , 2_n182 , 2_n183 , 2_n184 , 2_n185 , 2_n186 , 2_n187 , 2_n188 , 2_n189 , 2_n190 , 2_n191 , 2_n192 , 2_n193 , 2_n194 , 2_n195 , 2_n196 , 2_n197 , 2_n198 , 2_n199 , 2_n200 , 2_n201 , 2_n202 , 2_n203 , 2_n204 , 2_n205 , 2_n206 , 2_n207 , 2_n208 , 2_n209 , 2_n210 , 2_n211 , 2_n212 , 2_n213 , 2_n214 , 2_n215 , 2_n216 , 2_n218 , 2_n219 , 2_n220 , 2_n221 , 2_n222 , 2_n223 , 2_n224 , 2_n225 , 2_n227 , 2_n228 , 2_n229 , 2_n230 , 2_n231 , 2_n232 , 2_n233 , 2_n234 , 2_n235 , 2_n236 , 2_n237 , 2_n238 , 2_n239 , 2_n240 , 2_n241 , 2_n242 , 2_n243 , 2_n244 , 2_n245 , 2_n246 , 2_n247 , 2_n248 , 2_n249 , 2_n250 , 2_n251 , 2_n252 , 2_n253 , 2_n254 , 2_n255 , 2_n256 , 2_n257 , 2_n258 , 2_n259 , 2_n260 , 2_n261 , 2_n262 , 2_n263 , 2_n264 , 2_n265 , 2_n266 , 2_n267 , 2_n268 , 2_n269 , 2_n270 , 2_n271 , 2_n272 , 2_n273 , 2_n274 , 2_n275 , 2_n276 , 2_n277 , 2_n278 , 2_n279 , 2_n280 , 2_n281 , 2_n282 , 2_n283 , 2_n284 , 2_n285 , 2_n286 , 2_n287 , 2_n288 , 2_n289 , 2_n290 , 2_n291 , 2_n292 , 2_n293 , 2_n294 , 2_n295 , 2_n296 , 2_n297 , 2_n298 , 2_n299 , 2_n300 , 2_n301 , 2_n302 , 2_n303 , 2_n304 , 2_n305 , 2_n306 , 2_n307 , 2_n308 , 2_n309 , 2_n310 , 2_n311 , 2_n312 , 2_n313 , 2_n314 , 2_n315 , 2_n316 , 2_n317 , 2_n318 , 2_n319 , 2_n320 , 2_n321 , 2_n322 , 2_n323 , 2_n324 , 2_n325 , 2_n326 , 2_n327 , 2_n328 , 2_n329 , 2_n330 , 2_n331 , 2_n332 , 2_n333 , 2_n334 , 2_n335 , 2_n336 , 2_n337 , 2_n338 , 2_n339 , 2_n340 , 2_n341 , 2_n342 , 2_n343 , 2_n344 , 2_n345 , 2_n346 , 2_n347 , 2_n348 , 2_n349 , 2_n350 , 2_n351 , 2_n352 , 2_n353 , 2_n354 , 2_n355 , 2_n356 , 2_n357 , 2_n358 , 2_n359 , 2_n360 , 2_n361 , 2_n362 , 2_n363 , 2_n364 , 2_n365 , 2_n366 , 2_n367 , 2_n368 , 2_n369 , 2_n370 , 2_n371 , 2_n372 , 2_n373 , 2_n374 , 2_n375 , 2_n376 , 2_n377 , 2_n378 , 2_n379 , 2_n380 , 2_n382 , 2_n383 , 2_n384 , 2_n385 , 2_n386 , 2_n387 , 2_n388 , 2_n389 , 2_n390 , 2_n391 , 2_n392 , 2_n393 , 2_n394 , 2_n395 , 2_n396 , 2_n398 , 2_n399 , 2_n400 , 2_n401 , 2_n402 , 2_n403 , 2_n404 , 2_n406 , 2_n407 , 2_n408 , 2_n409 , 2_n410 , 2_n411 , 2_n412 , 2_n413 , 2_n414 , 2_n415 , 2_n416 , 2_n417 , 2_n418 , 2_n419 , 2_n420 , 2_n421 , 2_n422 , 2_n423 , 2_n424 , 2_n425 , 2_n426 , 2_n427 , 2_n428 , 2_n429 , 2_n430 , 2_n431 , 2_n432 , 2_n433 , 2_n434 , 2_n435 , 2_n436 , 2_n437 , 2_n438 , 2_n439 , 2_n440 , 2_n441 , 2_n442 , 2_n443 , 2_n444 , 2_n445 , 2_n446 , 2_n448 , 2_n449 , 2_n450 , 2_n451 , 2_n452 , 2_n453 , 2_n454 , 2_n455 , 2_n456 , 2_n457 , 2_n458 , 2_n459 , 2_n460 , 2_n461 , 2_n462 , 2_n463 , 2_n464 , 2_n465 , 2_n466 , 2_n467 , 2_n468 , 2_n469 , 2_n470 , 2_n471 , 2_n472 , 2_n473 , 2_n474 , 2_n475 , 2_n476 , 2_n477 , 2_n478 , 2_n479 , 2_n480 , 2_n481 , 2_n482 , 2_n483 , 2_n484 , 2_n485 , 2_n486 , 2_n487 , 2_n488 , 2_n489 , 2_n490 , 2_n491 , 2_n492 , 2_n493 , 2_n494 , 2_n495 , 2_n496 , 2_n497 , 2_n498 , 2_n499 , 2_n500 , 2_n501 , 2_n502 , 2_n504 , 2_n505 , 2_n506 , 2_n507 , 2_n508 , 2_n509 , 2_n510 , 2_n511 , 2_n512 , 2_n513 , 2_n514 , 2_n515 , 2_n516 , 2_n517 , 2_n518 , 2_n519 , 2_n520 , 2_n522 , 2_n523 , 2_n524 , 2_n525 , 2_n526 , 2_n527 , 2_n528 , 2_n529 , 2_n530 , 2_n531 , 2_n532 , 2_n534 , 2_n535 , 2_n536 , 2_n537 , 2_n538 , 2_n539 , 2_n540 , 2_n541 , 2_n542 , 2_n543 , 2_n544 , 2_n545 , 2_n546 , 2_n547 , 2_n548 , 2_n549 , 2_n550 , 2_n551 , 2_n552 , 2_n553 , 2_n554 , 2_n555 , 2_n556 , 2_n557 , 2_n558 , 2_n559 , 2_n560 , 2_n561 , 2_n562 , 2_n563 , 2_n564 , 2_n565 , 2_n566 , 2_n567 , 2_n568 , 2_n569 , 2_n570 , 2_n571 , 2_n572 , 2_n573 , 2_n574 , 2_n575 , 2_n576 , 2_n577 , 2_n578 , 2_n579 , 2_n580 , 2_n581 , 2_n582 , 2_n583 , 2_n584 , 2_n585 , 2_n586 , 2_n587 , 2_n588 , 2_n589 , 2_n590 , 2_n591 , 2_n592 , 2_n593 , 2_n594 , 2_n595 , 2_n596 , 2_n597 , 2_n598 , 2_n599 , 2_n600 , 2_n601 , 2_n602 , 2_n603 , 2_n604 , 2_n605 , 2_n606 , 2_n607 , 2_n608 , 2_n609 , 2_n610 , 2_n611 , 2_n612 , 2_n613 , 2_n614 , 2_n616 , 2_n617 , 2_n618 , 2_n619 , 2_n620 , 2_n621 , 2_n622 , 2_n623 , 2_n624 , 2_n625 , 2_n626 , 2_n627 , 2_n628 , 2_n629 , 2_n630 , 2_n631 , 2_n632 , 2_n633 , 2_n634 , 2_n635 , 2_n636 , 2_n637 , 2_n638 , 2_n639 , 2_n640 , 2_n641 , 2_n642 , 2_n643 , 2_n644 , 2_n645 , 2_n646 , 2_n647 , 2_n648 , 2_n649 , 2_n650 , 2_n651 , 2_n652 , 2_n653 , 2_n654 , 2_n655 , 2_n656 , 2_n657 , 2_n659 , 2_n660 , 2_n661 , 2_n662 , 2_n663 , 2_n664 , 2_n665 , 2_n666 , 2_n667 , 2_n668 , 2_n669 , 2_n670 , 2_n672 , 2_n673 , 2_n674 , 2_n675 , 2_n676 , 2_n677 , 2_n678 , 2_n679 , 2_n680 , 2_n681 , 2_n682 , 2_n683 , 2_n684 , 2_n685 , 2_n686 , 2_n687 , 2_n688 , 2_n689 , 2_n690 , 2_n691 , 2_n692 , 2_n693 , 2_n694 , 2_n695 , 2_n696 , 2_n697 , 2_n698 , 2_n699 , 2_n700 , 2_n701 , 2_n702 , 2_n703 , 2_n704 , 2_n705 , 2_n706 , 2_n707 , 2_n708 , 2_n709 , 2_n710 , 2_n711 , 2_n712 , 2_n713 , 2_n714 , 2_n715 , 2_n716 , 2_n717 , 2_n718 , 2_n719 , 2_n720 , 2_n721 , 2_n722 , 2_n723 , 2_n724 , 2_n725 , 2_n726 , 2_n727 , 2_n728 , 2_n729 , 2_n730 , 2_n731 , 2_n732 , 2_n733 , 2_n734 , 2_n735 , 2_n736 , 2_n737 , 2_n738 , 2_n739 , 2_n740 , 2_n741 , 2_n742 , 2_n743 , 2_n744 , 2_n745 , 2_n746 , 2_n747 , 2_n748 , 2_n749 , 2_n750 , 2_n751 , 2_n752 , 2_n754 , 2_n755 , 2_n756 , 2_n757 , 2_n758 , 2_n759 , 2_n760 , 2_n761 , 2_n762 , 2_n763 , 2_n764 , 2_n765 , 2_n766 , 2_n767 , 2_n768 , 2_n769 , 2_n770 , 2_n771 , 2_n772 , 2_n773 , 2_n774 , 2_n775 , 2_n776 , 2_n777 , 2_n778 , 2_n779 , 2_n780 , 2_n781 , 2_n782 , 2_n784 , 2_n785 , 2_n786 , 2_n787 , 2_n788 , 2_n789 , 2_n790 , 2_n791 , 2_n792 , 2_n793 , 2_n794 , 2_n795 , 2_n796 , 2_n797 , 2_n798 , 2_n799 , 2_n800 , 2_n801 , 2_n802 , 2_n803 , 2_n804 , 2_n805 , 2_n807 , 2_n808 , 2_n809 , 2_n810 , 2_n811 , 2_n812 , 2_n813 , 2_n814 , 2_n815 , 2_n816 , 2_n817 , 2_n818 , 2_n819 , 2_n820 , 2_n821 , 2_n822 , 2_n823 , 2_n824 , 2_n825 , 2_n826 , 2_n827 , 2_n828 , 2_n829 , 2_n830 , 2_n831 , 2_n832 , 2_n833 , 2_n834 , 2_n835 , 2_n836 , 2_n838 , 2_n839 , 2_n840 , 2_n841 , 2_n842 , 2_n843 , 2_n845 , 2_n846 , 2_n847 , 2_n848 , 2_n849 , 2_n850 , 2_n851 , 2_n852 , 2_n853 , 2_n854 , 2_n855 , 2_n856 , 2_n857 , 2_n858 , 2_n859 , 2_n860 , 2_n861 , 2_n862 , 2_n863 , 2_n864 , 2_n865 , 2_n866 , 2_n867 , 2_n868 , 2_n869 , 2_n870 , 2_n871 , 2_n872 , 2_n873 , 2_n874 , 2_n875 , 2_n876 , 2_n877 , 2_n878 , 2_n879 , 2_n880 , 2_n881 , 2_n882 , 2_n883 , 2_n884 , 2_n885 , 2_n886 , 2_n887 , 2_n888 , 2_n889 , 2_n890 , 2_n891 , 2_n892 , 2_n893 , 2_n894 , 2_n895 , 2_n896 , 2_n897 , 2_n898 , 2_n899 , 2_n900 , 2_n901 , 2_n902 , 2_n903 , 2_n904 , 2_n905 , 2_n906 , 2_n907 , 2_n908 , 2_n909 , 2_n910 , 2_n912 , 2_n913 , 2_n914 , 2_n915 , 2_n916 , 2_n917 , 2_n918 , 2_n919 , 2_n920 , 2_n921 , 2_n922 , 2_n923 , 2_n924 , 2_n925 , 2_n926 , 2_n927 , 2_n928 , 2_n929 , 2_n930 , 2_n931 , 2_n932 , 2_n933 , 2_n934 , 2_n935 , 2_n936 , 2_n937 , 2_n938 , 2_n939 , 2_n940 , 2_n941 , 2_n942 , 2_n943 , 2_n944 , 2_n945 , 2_n946 , 2_n947 , 2_n948 , 2_n949 , 2_n950 , 2_n951 , 2_n952 , 2_n953 , 2_n954 , 2_n955 , 2_n956 , 2_n957 , 2_n958 , 2_n959 , 2_n960 , 2_n961 , 2_n962 , 2_n963 , 2_n964 , 2_n965 , 2_n966 , 2_n967 , 2_n968 , 2_n969 , 2_n970 , 2_n971 , 2_n972 , 2_n973 , 2_n974 , 2_n975 , 2_n976 , 2_n977 , 2_n978 , 2_n979 , 2_n980 , 2_n981 , 2_n982 , 2_n983 , 2_n984 , 2_n985 , 2_n986 , 2_n987 , 2_n988 , 2_n989 , 2_n990 , 2_n991 , 2_n993 , 2_n994 , 2_n995 , 2_n997 , 2_n998 , 2_n999 , 2_n1000 , 2_n1001 , 2_n1002 , 2_n1003 , 2_n1004 , 2_n1005 , 2_n1006 , 2_n1007 , 2_n1008 , 2_n1009 , 2_n1010 , 2_n1011 , 2_n1012 , 2_n1013 , 2_n1014 , 2_n1015 , 2_n1016 , 2_n1017 , 2_n1018 , 2_n1019 , 2_n1021 , 2_n1022 , 2_n1023 , 2_n1024 , 2_n1025 , 2_n1026 , 2_n1027 , 2_n1028 , 2_n1029 , 2_n1030 , 2_n1031 , 2_n1032 , 2_n1033 , 2_n1034 , 2_n1035 , 2_n1036 , 2_n1037 , 2_n1038 , 2_n1039 , 2_n1040 , 2_n1041 , 2_n1042 , 2_n1043 , 2_n1044 , 2_n1045 , 2_n1046 , 2_n1047 , 2_n1048 , 2_n1049 , 2_n1050 , 2_n1051 , 2_n1052 , 2_n1053 , 2_n1054 , 2_n1055 , 2_n1056 , 2_n1057 , 2_n1058 , 2_n1059 , 2_n1060 , 2_n1061 , 2_n1062 , 2_n1063 , 2_n1064 , 2_n1065 , 2_n1066 , 2_n1068 , 2_n1069 , 2_n1070 , 2_n1071 , 2_n1072 , 2_n1073 , 2_n1074 , 2_n1075 , 2_n1076 , 2_n1077 , 2_n1078 , 2_n1079 , 2_n1080 , 2_n1081 , 2_n1082 , 2_n1083 , 2_n1084 , 2_n1085 , 2_n1086 , 2_n1087 , 2_n1088 , 2_n1089 , 2_n1090 , 2_n1091 , 2_n1092 , 2_n1093 , 2_n1095 , 2_n1096 , 2_n1098 , 2_n1099 , 2_n1100 , 2_n1101 , 2_n1102 , 2_n1103 , 2_n1104 , 2_n1105 , 2_n1106 , 2_n1107 , 2_n1108 , 2_n1109 , 2_n1110 , 2_n1111 , 2_n1112 , 2_n1113 , 2_n1114 , 2_n1115 , 2_n1116 , 2_n1117 , 2_n1118 , 2_n1119 , 2_n1120 , 2_n1121 , 2_n1122 , 2_n1123 , 2_n1124 , 2_n1125 , 2_n1126 , 2_n1127 , 2_n1128 , 2_n1129 , 2_n1130 , 2_n1131 , 2_n1132 , 2_n1133 , 2_n1134 , 2_n1135 , 2_n1137 , 2_n1139 , 2_n1140 , 2_n1141 , 2_n1142 , 2_n1143 , 2_n1144 , 2_n1145 , 2_n1146 , 2_n1147 , 2_n1148 , 2_n1149 , 2_n1150 , 2_n1151 , 2_n1152 , 2_n1153 , 2_n1154 , 2_n1155 , 2_n1156 , 2_n1157 , 2_n1158 , 2_n1159 , 2_n1160 , 2_n1161 , 2_n1162 , 2_n1163 , 2_n1164 , 2_n1165 , 2_n1166 , 2_n1167 , 2_n1168 , 2_n1169 , 2_n1170 , 2_n1171 , 2_n1172 , 2_n1173 , 2_n1174 , 2_n1175 , 2_n1176 , 2_n1177 , 2_n1178 , 2_n1179 , 2_n1180 , 2_n1181 , 2_n1182 , 2_n1183 , 2_n1184 , 2_n1185 , 2_n1186 , 2_n1187 , 2_n1188 , 2_n1189 , 2_n1190 , 2_n1191 , 2_n1192 , 2_n1193 , 2_n1194 , 2_n1195 , 2_n1196 , 2_n1197 , 2_n1200 , 2_n1201 , 2_n1202 , 2_n1203 , 2_n1204 , 2_n1205 , 2_n1206 , 2_n1207 , 2_n1208 , 2_n1210 , 2_n1211 , 2_n1212 , 2_n1213 , 2_n1214 , 2_n1215 , 2_n1216 , 2_n1217 , 2_n1218 , 2_n1219 , 2_n1220 , 2_n1221 , 2_n1222 , 2_n1223 , 2_n1224 , 2_n1225 , 2_n1226 , 2_n1227 , 2_n1228 , 2_n1229 , 2_n1230 , 2_n1231 , 2_n1232 , 2_n1233 , 2_n1234 , 2_n1235 , 2_n1236 , 2_n1237 , 2_n1238 , 2_n1239 , 2_n1240 , 2_n1241 , 2_n1242 , 2_n1243 , 2_n1244 , 2_n1245 , 2_n1246 , 2_n1247 , 2_n1248 , 2_n1249 , 2_n1250 , 2_n1251 , 2_n1252 , 2_n1253 , 2_n1254 , 2_n1255 , 2_n1256 , 2_n1257 , 2_n1258 , 2_n1259 , 2_n1260 , 2_n1261 , 2_n1262 , 2_n1263 , 2_n1264 , 2_n1265 , 2_n1266 , 2_n1267 , 2_n1268 , 2_n1270 , 2_n1271 , 2_n1272 , 2_n1273 , 2_n1274 , 2_n1275 , 2_n1276 , 2_n1277 , 2_n1278 , 2_n1279 , 2_n1280 , 2_n1281 , 2_n1282 , 2_n1283 , 2_n1284 , 2_n1285 , 2_n1286 , 2_n1287 , 2_n1288 , 2_n1289 , 2_n1290 , 2_n1291 , 2_n1292 , 2_n1293 , 2_n1294 , 2_n1295 , 2_n1296 , 2_n1297 , 2_n1298 , 2_n1299 , 2_n1300 , 2_n1301 , 2_n1302 , 2_n1303 , 2_n1304 , 2_n1305 , 2_n1306 , 2_n1307 , 2_n1308 , 2_n1309 , 2_n1310 , 2_n1311 , 2_n1312 , 2_n1313 , 2_n1314 , 2_n1315 , 2_n1316 , 2_n1317 , 2_n1318 , 2_n1319 , 2_n1320 , 2_n1321 , 2_n1322 , 2_n1323 , 2_n1324 , 2_n1325 , 2_n1326 , 2_n1327 , 2_n1328 , 2_n1329 , 2_n1330 , 2_n1331 , 2_n1332 , 2_n1334 , 2_n1335 , 2_n1336 , 2_n1337 , 2_n1338 , 2_n1339 , 2_n1340 , 2_n1341 , 2_n1342 , 2_n1343 , 2_n1344 , 2_n1345 , 2_n1346 , 2_n1347 , 2_n1348 , 2_n1349 , 2_n1350 , 2_n1351 , 2_n1352 , 2_n1354 , 2_n1355 , 2_n1356 , 2_n1358 , 2_n1359 , 2_n1360 , 2_n1361 , 2_n1362 , 2_n1363 , 2_n1364 , 2_n1365 , 2_n1366 , 2_n1367 , 2_n1368 , 2_n1369 , 2_n1370 , 2_n1371 , 2_n1372 , 2_n1373 , 2_n1374 , 2_n1375 , 2_n1376 , 2_n1377 , 2_n1378 , 2_n1379 , 2_n1380 , 2_n1381 , 2_n1382 , 2_n1383 , 2_n1384 , 2_n1385 , 2_n1386 , 2_n1387 , 2_n1388 , 2_n1389 , 2_n1390 , 2_n1391 , 2_n1392 , 2_n1393 , 2_n1394 , 2_n1395 , 2_n1396 , 2_n1397 , 2_n1398 , 2_n1399 , 2_n1400 , 2_n1401 , 2_n1402 , 2_n1403 , 2_n1404 , 2_n1405 , 2_n1406 , 2_n1407 , 2_n1408 , 2_n1409 , 2_n1410 , 2_n1411 , 2_n1412 , 2_n1413 , 2_n1414 , 2_n1415 , 2_n1416 , 2_n1417 , 2_n1418 , 2_n1419 , 2_n1420 , 2_n1421 , 2_n1422 , 2_n1423 , 2_n1424 , 2_n1425 , 2_n1426 , 2_n1427 , 2_n1428 , 2_n1429 , 2_n1430 , 2_n1431 , 2_n1432 , 2_n1433 , 2_n1434 , 2_n1435 , 2_n1436 , 2_n1437 , 2_n1438 , 2_n1439 , 2_n1440 , 2_n1441 , 2_n1442 , 2_n1443 , 2_n1444 , 2_n1445 , 2_n1446 , 2_n1447 , 2_n1448 , 2_n1449 , 2_n1450 , 2_n1451 , 2_n1452 , 2_n1453 , 2_n1454 , 2_n1455 , 2_n1456 , 2_n1457 , 2_n1458 , 2_n1459 , 2_n1460 , 2_n1461 , 2_n1462 , 2_n1463 , 2_n1464 , 2_n1465 , 2_n1466 , 2_n1467 , 2_n1468 , 2_n1469 , 2_n1470 , 2_n1472 , 2_n1473 , 2_n1474 , 2_n1475 , 2_n1476 , 2_n1477 , 2_n1479 , 2_n1480 , 2_n1481 , 2_n1482 , 2_n1483 , 2_n1484 , 2_n1485 , 2_n1486 , 2_n1487 , 2_n1488 , 2_n1489 , 2_n1490 , 2_n1491 , 2_n1492 , 2_n1493 , 2_n1494 , 2_n1495 , 2_n1496 , 2_n1497 , 2_n1498 , 2_n1499 , 2_n1500 , 2_n1501 , 2_n1502 , 2_n1503 , 2_n1504 , 2_n1505 , 2_n1506 , 2_n1507 , 2_n1508 , 2_n1509 , 2_n1511 , 2_n1513 , 2_n1514 , 2_n1515 , 2_n1516 , 2_n1517 , 2_n1518 , 2_n1519 , 2_n1520 , 2_n1521 , 2_n1522 , 2_n1524 , 2_n1525 , 2_n1526 , 2_n1527 , 2_n1528 , 2_n1529 , 2_n1530 , 2_n1531 , 2_n1532 , 2_n1533 , 2_n1534 , 2_n1535 , 2_n1536 , 2_n1537 , 2_n1538 , 2_n1539 , 2_n1540 , 2_n1541 , 2_n1542 , 2_n1543 , 2_n1544 , 2_n1545 , 2_n1546 , 2_n1547 , 2_n1548 , 2_n1549 , 2_n1550 , 2_n1551 , 2_n1552 , 2_n1553 , 2_n1554 , 2_n1555 , 2_n1556 , 2_n1557 , 2_n1558 , 2_n1559 , 2_n1560 , 2_n1561 , 2_n1562 , 2_n1563 , 2_n1565 , 2_n1566 , 2_n1567 , 2_n1568 , 2_n1569 , 2_n1570 , 2_n1571 , 2_n1572 , 2_n1573 , 2_n1574 , 2_n1575 , 2_n1577 , 2_n1578 , 2_n1579 , 2_n1580 , 2_n1581 , 2_n1582 , 2_n1583 , 2_n1584 , 2_n1585 , 2_n1586 , 2_n1587 , 2_n1588 , 2_n1589 , 2_n1590 , 2_n1591 , 2_n1592 , 2_n1593 , 2_n1594 , 2_n1595 , 2_n1596 , 2_n1597 , 2_n1598 , 2_n1599 , 2_n1600 , 2_n1601 , 2_n1602 , 2_n1603 , 2_n1604 , 2_n1605 , 2_n1606 , 2_n1607 , 2_n1608 , 2_n1609 , 2_n1610 , 2_n1611 , 2_n1612 , 2_n1613 , 2_n1614 , 2_n1615 , 2_n1616 , 2_n1617 , 2_n1618 , 2_n1619 , 2_n1620 , 2_n1621 , 2_n1622 , 2_n1623 , 2_n1624 , 2_n1625 , 2_n1626 , 2_n1627 , 2_n1628 , 2_n1629 , 2_n1630 , 2_n1631 , 2_n1632 , 2_n1633 , 2_n1634 , 2_n1635 , 2_n1636 , 2_n1637 , 2_n1638 , 2_n1639 , 2_n1640 , 2_n1641 , 2_n1642 , 2_n1643 , 2_n1644 , 2_n1645 , 2_n1646 , 2_n1647 , 2_n1648 , 2_n1649 , 2_n1650 , 2_n1651 , 2_n1652 , 2_n1653 , 2_n1654 , 2_n1655 , 2_n1656 , 2_n1657 , 2_n1659 , 2_n1660 , 2_n1661 , 2_n1662 , 2_n1663 , 2_n1664 , 2_n1665 , 2_n1666 , 2_n1667 , 2_n1668 , 2_n1669 , 2_n1670 , 2_n1671 , 2_n1672 , 2_n1673 , 2_n1674 , 2_n1675 , 2_n1676 , 2_n1677 , 2_n1678 , 2_n1679 , 2_n1680 , 2_n1681 , 2_n1682 , 2_n1683 , 2_n1684 , 2_n1685 , 2_n1686 , 2_n1687 , 2_n1688 , 2_n1689 , 2_n1690 , 2_n1691 , 2_n1692 , 2_n1693 , 2_n1694 , 2_n1695 , 2_n1696 , 2_n1697 , 2_n1698 , 2_n1699 , 2_n1700 , 2_n1701 , 2_n1702 , 2_n1703 , 2_n1704 , 2_n1705 , 2_n1706 , 2_n1707 , 2_n1708 , 2_n1709 , 2_n1710 , 2_n1711 , 2_n1712 , 2_n1713 , 2_n1714 , 2_n1715 , 2_n1716 , 2_n1717 , 2_n1718 , 2_n1719 , 2_n1720 , 2_n1721 , 2_n1722 , 2_n1723 , 2_n1724 , 2_n1725 , 2_n1726 , 2_n1727 , 2_n1728 , 2_n1729 , 2_n1730 , 2_n1731 , 2_n1732 , 2_n1733 , 2_n1734 , 2_n1735 , 2_n1736 , 2_n1737 , 2_n1738 , 2_n1739 , 2_n1740 , 2_n1741 , 2_n1742 , 2_n1743 , 2_n1744 , 2_n1745 , 2_n1746 , 2_n1747 , 2_n1748 , 2_n1749 , 2_n1750 , 2_n1751 , 2_n1752 , 2_n1753 , 2_n1754 , 2_n1755 , 2_n1756 , 2_n1757 , 2_n1758 , 2_n1759 , 2_n1760 , 2_n1761 , 2_n1762 , 2_n1763 , 2_n1764 , 2_n1765 , 2_n1766 , 2_n1767 , 2_n1768 , 2_n1769 , 2_n1770 , 2_n1771 , 2_n1772 , 2_n1773 , 2_n1774 , 2_n1775 , 2_n1776 , 2_n1777 , 2_n1778 , 2_n1779 , 2_n1780 , 2_n1781 , 2_n1782 , 2_n1783 , 2_n1784 , 2_n1785 , 2_n1786 , 2_n1787 , 2_n1788 , 2_n1789 , 2_n1790 , 2_n1791 , 2_n1792 , 2_n1793 , 2_n1794 , 2_n1795 , 2_n1796 , 2_n1797 , 2_n1799 , 2_n1800 , 2_n1801 , 2_n1802 , 2_n1803 , 2_n1804 , 2_n1805 , 2_n1806 , 2_n1807 , 2_n1808 , 2_n1809 , 2_n1810 , 2_n1811 , 2_n1812 , 2_n1813 , 2_n1814 , 2_n1815 , 2_n1816 , 2_n1817 , 2_n1818 , 2_n1819 , 2_n1820 , 2_n1821 , 2_n1822 , 2_n1823 , 2_n1824 , 2_n1825 , 2_n1826 , 2_n1827 , 2_n1828 , 2_n1829 , 2_n1830 , 2_n1831 , 2_n1832 , 2_n1833 , 2_n1834 , 2_n1836 , 2_n1837 , 2_n1838 , 2_n1839 , 2_n1840 , 2_n1841 , 2_n1842 , 2_n1843 , 2_n1844 , 2_n1845 , 2_n1846 , 2_n1848 , 2_n1849 , 2_n1850 , 2_n1851 , 2_n1852 , 2_n1853 , 2_n1854 , 2_n1855 , 2_n1856 , 2_n1857 , 2_n1858 , 2_n1859 , 2_n1860 , 2_n1861 , 2_n1862 , 2_n1863 , 2_n1864 , 2_n1865 , 2_n1866 , 2_n1867 , 2_n1868 , 2_n1869 , 2_n1870 , 2_n1871 , 2_n1872 , 2_n1873 , 2_n1874 , 2_n1875 , 2_n1876 , 2_n1877 , 2_n1878 , 2_n1879 , 2_n1880 , 2_n1881 , 2_n1882 , 2_n1883 , 2_n1884 , 2_n1885 , 2_n1886 , 2_n1887 , 2_n1888 , 2_n1889 , 2_n1890 , 2_n1891 , 2_n1892 , 2_n1893 , 2_n1894 , 2_n1895 , 2_n1896 , 2_n1897 , 2_n1898 , 2_n1899 , 2_n1900 , 2_n1901 , 2_n1902 , 2_n1903 , 2_n1904 , 2_n1905 , 2_n1907 , 2_n1908 , 2_n1909 , 2_n1910 , 2_n1911 , 2_n1912 , 2_n1913 , 2_n1914 , 2_n1915 , 2_n1916 , 2_n1917 , 2_n1918 , 2_n1919 , 2_n1920 , 2_n1921 , 2_n1922 , 2_n1923 , 2_n1924 , 2_n1925 , 2_n1926 , 2_n1927 , 2_n1928 , 2_n1929 , 2_n1930 , 2_n1931 , 2_n1932 , 2_n1933 , 2_n1934 , 2_n1935 , 2_n1936 , 2_n1937 , 2_n1938 , 2_n1939 , 2_n1940 , 2_n1941 , 2_n1942 , 2_n1943 , 2_n1944 , 2_n1945 , 2_n1946 , 2_n1947 , 2_n1948 , 2_n1949 , 2_n1950 , 2_n1951 , 2_n1952 , 2_n1953 , 2_n1954 , 2_n1955 , 2_n1956 , 2_n1957 , 2_n1958 , 2_n1959 , 2_n1960 , 2_n1961 , 2_n1962 , 2_n1963 , 2_n1964 , 2_n1965 , 2_n1966 , 2_n1967 , 2_n1968 , 2_n1969 , 2_n1970 , 2_n1971 , 2_n1972 , 2_n1973 , 2_n1974 , 2_n1975 , 2_n1976 , 2_n1977 , 2_n1978 , 2_n1979 , 2_n1981 , 2_n1982 , 2_n1983 , 2_n1984 , 2_n1985 , 2_n1986 , 2_n1987 , 2_n1988 , 2_n1989 , 2_n1990 , 2_n1991 , 2_n1992 , 2_n1993 , 2_n1994 , 2_n1995 , 2_n1996 , 2_n1997 , 2_n1998 , 2_n1999 , 2_n2000 , 2_n2001 , 2_n2002 , 2_n2003 , 2_n2004 , 2_n2005 , 2_n2006 , 2_n2007 , 2_n2008 , 2_n2009 , 2_n2010 , 2_n2011 , 2_n2012 , 2_n2013 , 2_n2014 , 2_n2015 , 2_n2016 , 2_n2017 , 2_n2018 , 2_n2019 , 2_n2020 , 2_n2021 , 2_n2022 , 2_n2023 , 2_n2025 , 2_n2026 , 2_n2027 , 2_n2028 , 2_n2029 , 2_n2030 , 2_n2031 , 2_n2032 , 2_n2033 , 2_n2034 , 2_n2035 , 2_n2036 , 2_n2037 , 2_n2038 , 2_n2039 , 2_n2040 , 2_n2041 , 2_n2042 , 2_n2043 , 2_n2044 , 2_n2045 , 2_n2046 , 2_n2047 , 2_n2048 , 2_n2049 , 2_n2050 , 2_n2051 , 2_n2052 , 2_n2053 , 2_n2054 , 2_n2055 , 2_n2056 , 2_n2057 , 2_n2058 , 2_n2059 , 2_n2060 , 2_n2061 , 2_n2062 , 2_n2063 , 2_n2064 , 2_n2065 , 2_n2066 , 2_n2067 , 2_n2068 , 2_n2069 , 2_n2070 , 2_n2071 , 2_n2072 , 2_n2073 , 2_n2074 , 2_n2075 , 2_n2076 , 2_n2077 , 2_n2078 , 2_n2079 , 2_n2080 , 2_n2081 , 2_n2082 , 2_n2083 , 2_n2084 , 2_n2085 , 2_n2086 , 2_n2088 , 2_n2089 , 2_n2090 , 2_n2091 , 2_n2092 , 2_n2093 , 2_n2094 , 2_n2095 , 2_n2097 , 2_n2098 , 2_n2099 , 2_n2100 , 2_n2101 , 2_n2102 , 2_n2103 , 2_n2104 , 2_n2105 , 2_n2106 , 2_n2107 , 2_n2108 , 2_n2109 , 2_n2110 , 2_n2111 , 2_n2112 , 2_n2113 , 2_n2114 , 2_n2115 , 2_n2116 , 2_n2117 , 2_n2118 , 2_n2119 , 2_n2120 , 2_n2121 , 2_n2122 , 2_n2123 , 2_n2124 , 2_n2125 , 2_n2126 , 2_n2127 , 2_n2128 , 2_n2129 , 2_n2130 , 2_n2132 , 2_n2133 , 2_n2134 , 2_n2135 , 2_n2136 , 2_n2137 , 2_n2138 , 2_n2139 , 2_n2140 , 2_n2141 , 2_n2142 , 2_n2143 , 2_n2144 , 2_n2145 , 2_n2146 , 2_n2147 , 2_n2148 , 2_n2149 , 2_n2150 , 2_n2151 , 2_n2152 , 2_n2153 , 2_n2154 , 2_n2155 , 2_n2156 , 2_n2157 , 2_n2158 , 2_n2159 , 2_n2160 , 2_n2161 , 2_n2162 , 2_n2163 , 2_n2164 , 2_n2165 , 2_n2166 , 2_n2167 , 2_n2168 , 2_n2169 , 2_n2170 , 2_n2171 , 2_n2172 , 2_n2173 , 2_n2174 , 2_n2175 , 2_n2176 , 2_n2177 , 2_n2178 , 2_n2179 , 2_n2180 , 2_n2181 , 2_n2182 , 2_n2183 , 2_n2184 , 2_n2185 , 2_n2186 , 2_n2187 , 2_n2188 , 2_n2189 , 2_n2190 , 2_n2191 , 2_n2192 , 2_n2193 , 2_n2194 , 2_n2195 , 2_n2196 , 2_n2197 , 2_n2198 , 2_n2199 , 2_n2200 , 2_n2201 , 2_n2202 , 2_n2203 , 2_n2204 , 2_n2205 , 2_n2206 , 2_n2207 , 2_n2208 , 2_n2209 , 2_n2210 , 2_n2211 , 2_n2212 , 2_n2213 , 2_n2214 , 2_n2215 , 2_n2216 , 2_n2217 , 2_n2218 , 2_n2219 , 2_n2220 , 2_n2221 , 2_n2222 , 2_n2223 , 2_n2224 , 2_n2225 , 2_n2227 , 2_n2228 , 2_n2229 , 2_n2230 , 2_n2231 , 2_n2232 , 2_n2233 , 2_n2234 , 2_n2235 , 2_n2236 , 2_n2237 , 2_n2238 , 2_n2239 , 2_n2240 , 2_n2241 , 2_n2242 , 2_n2243 , 2_n2244 , 2_n2245 , 2_n2246 , 2_n2247 , 2_n2248 , 2_n2249 , 2_n2250 , 2_n2251 , 2_n2252 , 2_n2254 , 2_n2255 , 2_n2256 , 2_n2257 , 2_n2258 , 2_n2259 , 2_n2260 , 2_n2261 , 2_n2262 , 2_n2263 , 2_n2264 , 2_n2265 , 2_n2266 , 2_n2267 , 2_n2268 , 2_n2269 , 2_n2270 , 2_n2271 , 2_n2272 , 2_n2273 , 2_n2274 , 2_n2275 , 2_n2276 , 2_n2277 , 2_n2279 , 2_n2280 , 2_n2281 , 2_n2282 , 2_n2283 , 2_n2284 , 2_n2285 , 2_n2286 , 2_n2287 , 2_n2288 , 2_n2289 , 2_n2290 , 2_n2291 , 2_n2292 , 2_n2293 , 2_n2294 , 2_n2295 , 2_n2296 , 2_n2297 , 2_n2298 , 2_n2299 , 2_n2300 , 2_n2302 , 2_n2303 , 2_n2304 , 2_n2305 , 2_n2306 , 2_n2307 , 2_n2308 , 2_n2309 , 2_n2310 , 2_n2311 , 2_n2312 , 2_n2313 , 2_n2314 , 2_n2315 , 2_n2317 , 2_n2318 , 2_n2319 , 2_n2320 , 2_n2321 , 2_n2322 , 2_n2323 , 2_n2324 , 2_n2325 , 2_n2326 , 2_n2327 , 2_n2328 , 2_n2329 , 2_n2330 , 2_n2331 , 2_n2332 , 2_n2333 , 2_n2334 , 2_n2335 , 2_n2336 , 2_n2337 , 2_n2338 , 2_n2339 , 2_n2340 , 2_n2341 , 2_n2342 , 2_n2343 , 2_n2344 , 2_n2345 , 2_n2346 , 2_n2348 , 2_n2349 , 2_n2350 , 2_n2351 , 2_n2352 , 2_n2353 , 2_n2354 , 2_n2355 , 2_n2356 , 2_n2357 , 2_n2358 , 2_n2359 , 2_n2360 , 2_n2361 , 2_n2362 , 2_n2363 , 2_n2364 , 2_n2365 , 2_n2366 , 2_n2367 , 2_n2368 , 2_n2369 , 2_n2370 , 2_n2371 , 2_n2372 , 2_n2373 , 2_n2374 , 2_n2375 , 2_n2376 , 2_n2377 , 2_n2378 , 2_n2379 , 2_n2380 , 2_n2381 , 2_n2382 , 2_n2384 , 2_n2385 , 2_n2386 , 2_n2387 , 2_n2388 , 2_n2389 , 2_n2390 , 2_n2391 , 2_n2392 , 2_n2394 , 2_n2395 , 2_n2396 , 2_n2397 , 2_n2398 , 2_n2399 , 2_n2400 , 2_n2401 , 2_n2402 , 2_n2403 , 2_n2404 , 2_n2405 , 2_n2406 , 2_n2407 , 2_n2408 , 2_n2409 , 2_n2410 , 2_n2411 , 2_n2412 , 2_n2413 , 2_n2414 , 2_n2415 , 2_n2416 , 2_n2417 , 2_n2418 , 2_n2419 , 2_n2420 , 2_n2421 , 2_n2422 , 2_n2423 , 2_n2424 , 2_n2426 , 2_n2427 , 2_n2428 , 2_n2429 , 2_n2430 , 2_n2432 , 2_n2435 , 2_n2436 , 2_n2437 , 2_n2438 , 2_n2439 , 2_n2440 , 2_n2441 , 2_n2442 , 2_n2443 , 2_n2444 , 2_n2445 , 2_n2446 , 2_n2447 , 2_n2448 , 2_n2449 , 2_n2450 , 2_n2451 , 2_n2452 , 2_n2453 , 2_n2454 , 2_n2455 , 2_n2456 , 2_n2457 , 2_n2458 , 2_n2459 , 2_n2460 , 2_n2461 , 2_n2462 , 2_n2463 , 2_n2465 , 2_n2466 , 2_n2467 , 2_n2468 , 2_n2469 , 2_n2470 , 2_n2471 , 2_n2472 , 2_n2473 , 2_n2474 , 2_n2475 , 2_n2476 , 2_n2477 , 2_n2478 , 2_n2479 , 2_n2480 , 2_n2481 , 2_n2482 , 2_n2483 , 2_n2484 , 2_n2485 , 2_n2486 , 2_n2487 , 2_n2488 , 2_n2489 , 2_n2490 , 2_n2491 , 2_n2492 , 2_n2493 , 2_n2494 , 2_n2495 , 2_n2496 , 2_n2497 , 2_n2499 , 2_n2500 , 2_n2501 , 2_n2502 , 2_n2503 , 2_n2504 , 2_n2505 , 2_n2506 , 2_n2510 , 2_n2511 , 2_n2513 , 2_n2514 , 2_n2516 , 2_n2517 , 2_n2518 , 2_n2519 , 2_n2520 , 2_n2521 , 2_n2523 , 2_n2524 , 2_n2525 , 2_n2526 , 2_n2527 , 2_n2528 , 2_n2529 , 2_n2531 , 2_n2532 , 2_n2533 , 2_n2534 , 2_n2535 , 2_n2536 , 2_n2537 , 2_n2538 , 2_n2539 , 2_n2540 , 2_n2541 , 2_n2542 , 2_n2543 , 2_n2544 , 2_n2545 , 2_n2546 , 2_n2547 , 2_n2548 , 2_n2549 , 2_n2550 , 2_n2552 , 2_n2553 , 2_n2554 , 2_n2555 , 2_n2556 , 2_n2557 , 2_n2559 , 2_n2560 , 2_n2561 , 2_n2562 , 2_n2563 , 2_n2565 , 2_n2566 , 2_n2567 , 2_n2568 , 2_n2569 , 2_n2570 , 2_n2571 , 2_n2572 , 2_n2573 , 2_n2574 , 2_n2575 , 2_n2576 , 2_n2578 , 2_n2579 , 2_n2580 , 2_n2582 , 2_n2583 , 2_n2584 , 2_n2586 , 2_n2587 , 2_n2588 , 2_n2589 , 2_n2590 , 2_n2591 , 2_n2592 , 2_n2593 , 2_n2594 , 2_n2595 , 2_n2596 , 2_n2597 , 2_n2598 , 2_n2599 , 2_n2600 , 2_n2601 , 2_n2602 , 2_n2603 , 2_n2604 , 2_n2605 , 2_n2606 , 2_n2607 , 2_n2608 , 2_n2609 , 2_n2610 , 2_n2611 , 2_n2612 , 2_n2613 , 2_n2614 , 2_n2615 , 2_n2616 , 2_n2617 , 2_n2618 , 2_n2619 , 2_n2620 , 2_n2621 , 2_n2622 , 2_n2623 , 2_n2625 , 2_n2626 , 2_n2627 , 2_n2628 , 2_n2629 , 2_n2630 , 2_n2631 , 2_n2632 , 2_n2633 , 2_n2634 , 2_n2635 , 2_n2636 , 2_n2637 , 2_n2638 , 2_n2639 , 2_n2640 , 2_n2641 , 2_n2642 , 2_n2643 , 2_n2644 , 2_n2645 , 2_n2646 , 2_n2647 , 2_n2648 , 2_n2649 , 2_n2650 , 2_n2651 , 2_n2652 , 2_n2653 , 2_n2654 , 2_n2655 , 2_n2656 , 2_n2657 , 2_n2658 , 2_n2659 , 2_n2660 , 2_n2661 , 2_n2662 , 2_n2663 , 2_n2664 , 2_n2665 , 2_n2666 , 2_n2667 , 2_n2668 , 2_n2669 , 2_n2670 , 2_n2671 , 2_n2672 , 2_n2673 , 2_n2674 , 2_n2675 , 2_n2676 , 2_n2677 , 2_n2678 , 2_n2680 , 2_n2681 , 2_n2682 , 2_n2683 , 2_n2684 , 2_n2685 , 2_n2686 , 2_n2687 , 2_n2688 , 2_n2689 , 2_n2690 , 2_n2691 , 2_n2692 , 2_n2693 , 2_n2694 , 2_n2695 , 2_n2696 , 2_n2697 , 2_n2698 , 2_n2699 , 2_n2700 , 2_n2701 , 2_n2702 , 2_n2703 , 2_n2704 , 2_n2705 , 2_n2706 , 2_n2707 , 2_n2709 , 2_n2710 , 2_n2711 , 2_n2712 , 2_n2713 , 2_n2714 , 2_n2715 , 2_n2716 , 2_n2717 , 2_n2718 , 2_n2719 , 2_n2720 , 2_n2721 , 2_n2722 , 2_n2723 , 2_n2724 , 2_n2725 , 2_n2726 , 2_n2727 , 2_n2728 , 2_n2729 , 2_n2730 , 2_n2731 , 2_n2732 , 2_n2733 , 2_n2734 , 2_n2735 , 2_n2736 , 2_n2737 , 2_n2738 , 2_n2739 , 2_n2740 , 2_n2741 , 2_n2742 , 2_n2743 , 2_n2744 , 2_n2745 , 2_n2746 , 2_n2747 , 2_n2748 , 2_n2750 , 2_n2751 , 2_n2752 , 2_n2753 , 2_n2754 , 2_n2755 , 2_n2756 , 2_n2757 , 2_n2758 , 2_n2759 , 2_n2760 , 2_n2761 , 2_n2762 , 2_n2763 , 2_n2764 , 2_n2765 , 2_n2766 , 2_n2767 , 2_n2768 , 2_n2769 , 2_n2770 , 2_n2771 , 2_n2772 , 2_n2773 , 2_n2774 , 2_n2775 , 2_n2776 , 2_n2777 , 2_n2778 , 2_n2779 , 2_n2780 , 2_n2781 , 2_n2782 , 2_n2783 , 2_n2784 , 2_n2785 , 2_n2786 , 2_n2787 , 2_n2788 , 2_n2789 , 2_n2790 , 2_n2791 , 2_n2792 , 2_n2793 , 2_n2794 , 2_n2795 , 2_n2796 , 2_n2797 , 2_n2798 , 2_n2799 , 2_n2800 , 2_n2801 , 2_n2803 , 2_n2804 , 2_n2805 , 2_n2806 , 2_n2807 , 2_n2808 , 2_n2809 , 2_n2810 , 2_n2811 , 2_n2812 , 2_n2813 , 2_n2814 , 2_n2815 , 2_n2816 , 2_n2817 , 2_n2819 , 2_n2820 , 2_n2821 , 2_n2822 , 2_n2823 , 2_n2824 , 2_n2825 , 2_n2826 , 2_n2827 , 2_n2828 , 2_n2829 , 2_n2830 , 2_n2831 , 2_n2832 , 2_n2833 , 2_n2834 , 2_n2835 , 2_n2836 , 2_n2837 , 2_n2838 , 2_n2839 , 2_n2840 , 2_n2841 , 2_n2842 , 2_n2843 , 2_n2844 , 2_n2845 , 2_n2846 , 2_n2847 , 2_n2848 , 2_n2849 , 2_n2850 , 2_n2851 , 2_n2852 , 2_n2853 , 2_n2854 , 2_n2855 , 2_n2856 , 2_n2857 , 2_n2858 , 2_n2859 , 2_n2860 , 2_n2861 , 2_n2862 , 2_n2863 , 2_n2864 , 2_n2865 , 2_n2866 , 2_n2867 , 2_n2868 , 2_n2869 , 2_n2870 , 2_n2871 , 2_n2872 , 2_n2873 , 2_n2874 , 2_n2875 , 2_n2876 , 2_n2877 , 2_n2878 , 2_n2880 , 2_n2881 , 2_n2882 , 2_n2883 , 2_n2884 , 2_n2885 , 2_n2886 , 2_n2887 , 2_n2888 , 2_n2889 , 2_n2890 , 2_n2891 , 2_n2892 , 2_n2893 , 2_n2894 , 2_n2895 , 2_n2896 , 2_n2897 , 2_n2898 , 2_n2899 , 2_n2900 , 2_n2901 , 2_n2903 , 2_n2904 , 2_n2905 , 2_n2906 , 2_n2907 , 2_n2908 , 2_n2909 , 2_n2910 , 2_n2911 , 2_n2912 , 2_n2913 , 2_n2914 , 2_n2915 , 2_n2916 , 2_n2917 , 2_n2918 , 2_n2919 , 2_n2920 , 2_n2921 , 2_n2922 , 2_n2923 , 2_n2924 , 2_n2925 , 2_n2926 , 2_n2927 , 2_n2928 , 2_n2929 , 2_n2930 , 2_n2931 , 2_n2932 , 2_n2933 , 2_n2934 , 2_n2935 , 2_n2936 , 2_n2937 , 2_n2938 , 2_n2939 , 2_n2940 , 2_n2941 , 2_n2942 , 2_n2943 , 2_n2944 , 2_n2945 , 2_n2946 , 2_n2947 , 2_n2948 , 2_n2949 , 2_n2950 , 2_n2951 , 2_n2952 , 2_n2953 , 2_n2954 , 2_n2955 , 2_n2956 , 2_n2957 , 2_n2958 , 2_n2959 , 2_n2960 , 2_n2961 , 2_n2962 , 2_n2963 , 2_n2964 , 2_n2965 , 2_n2966 , 2_n2967 , 2_n2968 , 2_n2969 , 2_n2970 , 2_n2971 , 2_n2972 , 2_n2973 , 2_n2974 , 2_n2975 , 2_n2976 , 2_n2977 , 2_n2978 , 2_n2979 , 2_n2980 , 2_n2981 , 2_n2982 , 2_n2983 , 2_n2984 , 2_n2985 , 2_n2986 , 2_n2987 , 2_n2988 , 2_n2989 , 2_n2990 , 2_n2991 , 2_n2992 , 2_n2993 , 2_n2994 , 2_n2995 , 2_n2996 , 2_n2997 , 2_n2998 , 2_n2999 , 2_n3000 , 2_n3001 , 2_n3002 , 2_n3003 , 2_n3004 , 2_n3005 , 2_n3006 , 2_n3007 , 2_n3008 , 2_n3009 , 2_n3010 , 2_n3011 , 2_n3012 , 2_n3013 , 2_n3014 , 2_n3015 , 2_n3016 , 2_n3017 , 2_n3018 , 2_n3019 , 2_n3020 , 2_n3021 , 2_n3023 , 2_n3024 , 2_n3025 , 2_n3026 , 2_n3027 , 2_n3028 , 2_n3029 , 2_n3030 , 2_n3031 , 2_n3032 , 2_n3033 , 2_n3034 , 2_n3035 , 2_n3036 , 2_n3037 , 2_n3038 , 2_n3039 , 2_n3040 , 2_n3041 , 2_n3042 , 2_n3043 , 2_n3044 , 2_n3045 , 2_n3046 , 2_n3047 , 2_n3048 , 2_n3049 , 2_n3050 , 2_n3051 , 2_n3052 , 2_n3053 , 2_n3054 , 2_n3055 , 2_n3056 , 2_n3057 , 2_n3058 , 2_n3059 , 2_n3060 , 2_n3061 , 2_n3062 , 2_n3063 , 2_n3064 , 2_n3065 , 2_n3066 , 2_n3067 , 2_n3068 , 2_n3069 , 2_n3070 , 2_n3072 , 2_n3073 , 2_n3074 , 2_n3075 , 2_n3076 , 2_n3077 , 2_n3078 , 2_n3079 , 2_n3080 , 2_n3081 , 2_n3082 , 2_n3083 , 2_n3084 , 2_n3085 , 2_n3086 , 2_n3087 , 2_n3088 , 2_n3089 , 2_n3090 , 2_n3091 , 2_n3092 , 2_n3093 , 2_n3094 , 2_n3095 , 2_n3096 , 2_n3097 , 2_n3098 , 2_n3099 , 2_n3100 , 2_n3101 , 2_n3102 , 2_n3103 , 2_n3104 , 2_n3105 , 2_n3106 , 2_n3107 , 2_n3108 , 2_n3109 , 2_n3110 , 2_n3111 , 2_n3112 , 2_n3113 , 2_n3114 , 2_n3115 , 2_n3116 , 2_n3117 , 2_n3118 , 2_n3119 , 2_n3120 , 2_n3121 , 2_n3122 , 2_n3123 , 2_n3125 , 2_n3126 , 2_n3127 , 2_n3128 , 2_n3129 , 2_n3130 , 2_n3131 , 2_n3132 , 2_n3133 , 2_n3134 , 2_n3135 , 2_n3136 , 2_n3137 , 2_n3138 , 2_n3139 , 2_n3140 , 2_n3141 , 2_n3142 , 2_n3143 , 2_n3144 , 2_n3145 , 2_n3147 , 2_n3148 , 2_n3149 , 2_n3150 , 2_n3151 , 2_n3152 , 2_n3153 , 2_n3154 , 2_n3155 , 2_n3156 , 2_n3157 , 2_n3158 , 2_n3159 , 2_n3160 , 2_n3161 , 2_n3162 , 2_n3163 , 2_n3164 , 2_n3165 , 2_n3166 , 2_n3167 , 2_n3168 , 2_n3169 , 2_n3170 , 2_n3171 , 2_n3173 , 2_n3174 , 2_n3175 , 2_n3176 , 2_n3177 , 2_n3178 , 2_n3179 , 2_n3180 , 2_n3181 , 2_n3182 , 2_n3183 , 2_n3184 , 2_n3185 , 2_n3186 , 2_n3187 , 2_n3188 , 2_n3189 , 2_n3190 , 2_n3191 , 2_n3192 , 2_n3193 , 2_n3194 , 2_n3195 , 2_n3196 , 2_n3197 , 2_n3198 , 2_n3199 , 2_n3200 , 2_n3201 , 2_n3202 , 2_n3203 , 2_n3204 , 2_n3205 , 2_n3206 , 2_n3207 , 2_n3208 , 2_n3209 , 2_n3210 , 2_n3211 , 2_n3212 , 2_n3213 , 2_n3215 , 2_n3216 , 2_n3217 , 2_n3218 , 2_n3219 , 2_n3220 , 2_n3221 , 2_n3222 , 2_n3223 , 2_n3224 , 2_n3225 , 2_n3226 , 2_n3227 , 2_n3228 , 2_n3229 , 2_n3231 , 2_n3232 , 2_n3233 , 2_n3234 , 2_n3235 , 2_n3236 , 2_n3237 , 2_n3238 , 2_n3239 , 2_n3240 , 2_n3241 , 2_n3242 , 2_n3243 , 2_n3244 , 2_n3245 , 2_n3246 , 2_n3247 , 2_n3248 , 2_n3249 , 2_n3250 , 2_n3251 , 2_n3252 , 2_n3253 , 2_n3254 , 2_n3255 , 2_n3256 , 2_n3257 , 2_n3258 , 2_n3259 , 2_n3260 , 2_n3261 , 2_n3262 , 2_n3263 , 2_n3264 , 2_n3265 , 2_n3266 , 2_n3267 , 2_n3268 , 2_n3269 , 2_n3270 , 2_n3271 , 2_n3273 , 2_n3274 , 2_n3275 , 2_n3276 , 2_n3277 , 2_n3278 , 2_n3279 , 2_n3280 , 2_n3281 , 2_n3282 , 2_n3283 , 2_n3284 , 2_n3285 , 2_n3286 , 2_n3288 , 2_n3289 , 2_n3290 , 2_n3291 , 2_n3292 , 2_n3293 , 2_n3294 , 2_n3295 , 2_n3296 , 2_n3297 , 2_n3298 , 2_n3299 , 2_n3300 , 2_n3301 , 2_n3302 , 2_n3303 , 2_n3304 , 2_n3305 , 2_n3306 , 2_n3307 , 2_n3308 , 2_n3309 , 2_n3310 , 2_n3311 , 2_n3312 , 2_n3313 , 2_n3314 , 2_n3315 , 2_n3316 , 2_n3317 , 2_n3318 , 2_n3319 , 2_n3320 , 2_n3321 , 2_n3322 , 2_n3323 , 2_n3324 , 2_n3325 , 2_n3326 , 2_n3327 , 2_n3328 , 2_n3329 , 2_n3330 , 2_n3331 , 2_n3332 , 2_n3333 , 2_n3334 , 2_n3335 , 2_n3336 , 2_n3337 , 2_n3338 , 2_n3340 , 2_n3341 , 2_n3343 , 2_n3344 , 2_n3345 , 2_n3346 , 2_n3347 , 2_n3348 , 2_n3349 , 2_n3350 , 2_n3351 , 2_n3352 , 2_n3353 , 2_n3354 , 2_n3355 , 2_n3356 , 2_n3357 , 2_n3358 , 2_n3359 , 2_n3360 , 2_n3361 , 2_n3362 , 2_n3363 , 2_n3364 , 2_n3365 , 2_n3366 , 2_n3367 , 2_n3368 , 2_n3369 , 2_n3370 , 2_n3371 , 2_n3372 , 2_n3373 , 2_n3374 , 2_n3375 , 2_n3376 , 2_n3377 , 2_n3378 , 2_n3379 , 2_n3380 , 2_n3381 , 2_n3382 , 2_n3383 , 2_n3384 , 2_n3385 , 2_n3386 , 2_n3387 , 2_n3388 , 2_n3389 , 2_n3390 , 2_n3391 , 2_n3392 , 2_n3393 , 2_n3394 , 2_n3395 , 2_n3396 , 2_n3397 , 2_n3398 , 2_n3399 , 2_n3400 , 2_n3401 , 2_n3402 , 2_n3403 , 2_n3404 , 2_n3405 , 2_n3406 , 2_n3407 , 2_n3408 , 2_n3409 , 2_n3410 , 2_n3411 , 2_n3412 , 2_n3413 , 2_n3414 , 2_n3415 , 2_n3416 , 2_n3417 , 2_n3418 , 2_n3419 , 2_n3420 , 2_n3421 , 2_n3422 , 2_n3423 , 2_n3424 , 2_n3425 , 2_n3426 , 2_n3427 , 2_n3428 , 2_n3429 , 2_n3430 , 2_n3431 , 2_n3432 , 2_n3433 , 2_n3434 , 2_n3435 , 2_n3436 , 2_n3437 , 2_n3438 , 2_n3439 , 2_n3440 , 2_n3441 , 2_n3442 , 2_n3443 , 2_n3444 , 2_n3445 , 2_n3446 , 2_n3447 , 2_n3448 , 2_n3449 , 2_n3450 , 2_n3451 , 2_n3452 , 2_n3453 , 2_n3454 , 2_n3455 , 2_n3457 , 2_n3458 , 2_n3459 , 2_n3460 , 2_n3461 , 2_n3462 , 2_n3463 , 2_n3464 , 2_n3465 , 2_n3466 , 2_n3467 , 2_n3468 , 2_n3469 , 2_n3470 , 2_n3471 , 2_n3472 , 2_n3473 , 2_n3474 , 2_n3475 , 2_n3476 , 2_n3477 , 2_n3478 , 2_n3479 , 2_n3480 , 2_n3481 , 2_n3482 , 2_n3483 , 2_n3484 , 2_n3485 , 2_n3486 , 2_n3487 , 2_n3488 , 2_n3489 , 2_n3490 , 2_n3491 , 2_n3492 , 2_n3493 , 2_n3494 , 2_n3495 , 2_n3496 , 2_n3497 , 2_n3498 , 2_n3499 , 2_n3500 , 2_n3501 , 2_n3502 , 2_n3503 , 2_n3504 , 2_n3505 , 2_n3506 , 2_n3507 , 2_n3508 , 2_n3509 , 2_n3510 , 2_n3511 , 2_n3512 , 2_n3513 , 2_n3514 , 2_n3515 , 2_n3516 , 2_n3517 , 2_n3518 , 2_n3519 , 2_n3520 , 2_n3521 , 2_n3522 , 2_n3523 , 2_n3524 , 2_n3525 , 2_n3526 , 2_n3527 , 2_n3528 , 2_n3529 , 2_n3530 , 2_n3531 , 2_n3532 , 2_n3533 , 2_n3534 , 2_n3535 , 2_n3536 , 2_n3537 , 2_n3538 , 2_n3539 , 2_n3540 , 2_n3541 , 2_n3542 , 2_n3543 , 2_n3544 , 2_n3545 , 2_n3546 , 2_n3547 , 2_n3548 , 2_n3549 , 2_n3550 , 2_n3551 , 2_n3552 , 2_n3553 , 2_n3554 , 2_n3555 , 2_n3556 , 2_n3557 , 2_n3558 , 2_n3559 , 2_n3560 , 2_n3561 , 2_n3562 , 2_n3563 , 2_n3564 , 2_n3565 , 2_n3566 , 2_n3567 , 2_n3568 , 2_n3569 , 2_n3570 , 2_n3571 , 2_n3572 , 2_n3573 , 2_n3574 , 2_n3575 , 2_n3576 , 2_n3577 , 2_n3578 , 2_n3579 , 2_n3580 , 2_n3581 , 2_n3582 , 2_n3583 , 2_n3584 , 2_n3585 , 2_n3586 , 2_n3587 , 2_n3588 , 2_n3589 , 2_n3590 , 2_n3591 , 2_n3592 , 2_n3593 , 2_n3594 , 2_n3595 , 2_n3596 , 2_n3597 , 2_n3598 , 2_n3599 , 2_n3600 , 2_n3601 , 2_n3603 , 2_n3604 , 2_n3605 , 2_n3606 , 2_n3607 , 2_n3608 , 2_n3609 , 2_n3610 , 2_n3611 , 2_n3612 , 2_n3613 , 2_n3614 , 2_n3615 , 2_n3617 , 2_n3618 , 2_n3619 , 2_n3620 , 2_n3621 , 2_n3622 , 2_n3623 , 2_n3624 , 2_n3625 , 2_n3626 , 2_n3628 , 2_n3629 , 2_n3630 , 2_n3631 , 2_n3632 , 2_n3633 , 2_n3634 , 2_n3635 , 2_n3636 , 2_n3637 , 2_n3638 , 2_n3639 , 2_n3640 , 2_n3641 , 2_n3642 , 2_n3643 , 2_n3644 , 2_n3645 , 2_n3646 , 2_n3647 , 2_n3648 , 2_n3649 , 2_n3650 , 2_n3651 , 2_n3652 , 2_n3653 , 2_n3655 , 2_n3656 , 2_n3657 , 2_n3658 , 2_n3659 , 2_n3660 , 2_n3662 , 2_n3663 , 2_n3664 , 2_n3665 , 2_n3666 , 2_n3667 , 2_n3668 , 2_n3669 , 2_n3670 , 2_n3671 , 2_n3672 , 2_n3673 , 2_n3674 , 2_n3675 , 2_n3676 , 2_n3678 , 2_n3679 , 2_n3680 , 2_n3681 , 2_n3682 , 2_n3683 , 2_n3684 , 2_n3685 , 2_n3686 , 2_n3687 , 2_n3688 , 2_n3689 , 2_n3690 , 2_n3691 , 2_n3692 , 2_n3693 , 2_n3694 , 2_n3695 , 2_n3696 , 2_n3697 , 2_n3698 , 2_n3699 , 2_n3700 , 2_n3701 , 2_n3702 , 2_n3703 , 2_n3704 , 2_n3705 , 2_n3706 , 2_n3707 , 2_n3708 , 2_n3709 , 2_n3710 , 2_n3711 , 2_n3712 , 2_n3713 , 2_n3714 , 2_n3715 , 2_n3716 , 2_n3717 , 2_n3718 , 2_n3720 , 2_n3721 , 2_n3722 , 2_n3723 , 2_n3724 , 2_n3725 , 2_n3726 , 2_n3727 , 2_n3728 , 2_n3729 , 2_n3730 , 2_n3731 , 2_n3732 , 2_n3733 , 2_n3734 , 2_n3735 , 2_n3736 , 2_n3737 , 2_n3738 , 2_n3739 , 2_n3740 , 2_n3741 , 2_n3742 , 2_n3743 , 2_n3744 , 2_n3745 , 2_n3746 , 2_n3747 , 2_n3748 , 2_n3749 , 2_n3750 , 2_n3751 , 2_n3752 , 2_n3753 , 2_n3755 , 2_n3756 , 2_n3757 , 2_n3758 , 2_n3759 , 2_n3760 , 2_n3761 , 2_n3762 , 2_n3763 , 2_n3764 , 2_n3765 , 2_n3766 , 2_n3767 , 2_n3768 , 2_n3769 , 2_n3770 , 2_n3771 , 2_n3772 , 2_n3773 , 2_n3774 , 2_n3775 , 2_n3776 , 2_n3777 , 2_n3778 , 2_n3779 , 2_n3780 , 2_n3781 , 2_n3782 , 2_n3783 , 2_n3784 , 2_n3785 , 2_n3786 , 2_n3787 , 2_n3788 , 2_n3789 , 2_n3790 , 2_n3791 , 2_n3792 , 2_n3793 , 2_n3794 , 2_n3795 , 2_n3796 , 2_n3797 , 2_n3798 , 2_n3799 , 2_n3800 , 2_n3801 , 2_n3802 , 2_n3803 , 2_n3804 , 2_n3805 , 2_n3806 , 2_n3807 , 2_n3808 , 2_n3809 , 2_n3810 , 2_n3811 , 2_n3812 , 2_n3813 , 2_n3814 , 2_n3815 , 2_n3816 , 2_n3817 , 2_n3818 , 2_n3819 , 2_n3820 , 2_n3821 , 2_n3822 , 2_n3823 , 2_n3824 , 2_n3825 , 2_n3826 , 2_n3827 , 2_n3828 , 2_n3829 , 2_n3830 , 2_n3831 , 2_n3832 , 2_n3833 , 2_n3834 , 2_n3835 , 2_n3836 , 2_n3837 , 2_n3838 , 2_n3839 , 2_n3840 , 2_n3841 , 2_n3843 , 2_n3844 , 2_n3845 , 2_n3846 , 2_n3847 , 2_n3848 , 2_n3850 , 2_n3851 , 2_n3852 , 2_n3853 , 2_n3854 , 2_n3855 , 2_n3856 , 2_n3857 , 2_n3858 , 2_n3859 , 2_n3860 , 2_n3861 , 2_n3862 , 2_n3863 , 2_n3864 , 2_n3866 , 2_n3867 , 2_n3868 , 2_n3869 , 2_n3870 , 2_n3871 , 2_n3872 , 2_n3873 , 2_n3874 , 2_n3875 , 2_n3876 , 2_n3877 , 2_n3878 , 2_n3879 , 2_n3880 , 2_n3881 , 2_n3882 , 2_n3883 , 2_n3884 , 2_n3885 , 2_n3886 , 2_n3887 , 2_n3888 , 2_n3889 , 2_n3890 , 2_n3891 , 2_n3892 , 2_n3893 , 2_n3894 , 2_n3895 , 2_n3896 , 2_n3897 , 2_n3898 , 2_n3899 , 2_n3900 , 2_n3901 , 2_n3902 , 2_n3903 , 2_n3904 , 2_n3905 , 2_n3906 , 2_n3907 , 2_n3908 , 2_n3909 , 2_n3910 , 2_n3911 , 2_n3912 , 2_n3913 , 2_n3914 , 2_n3915 , 2_n3916 , 2_n3917 , 2_n3918 , 2_n3919 , 2_n3920 , 2_n3921 , 2_n3922 , 2_n3923 , 2_n3924 , 2_n3925 , 2_n3926 , 2_n3927 , 2_n3928 , 2_n3929 , 2_n3930 , 2_n3931 , 2_n3933 , 2_n3934 , 2_n3935 , 2_n3936 , 2_n3937 , 2_n3938 , 2_n3939 , 2_n3940 , 2_n3941 , 2_n3942 , 2_n3943 , 2_n3944 , 2_n3945 , 2_n3946 , 2_n3947 , 2_n3948 , 2_n3949 , 2_n3950 , 2_n3951 , 2_n3952 , 2_n3953 , 2_n3954 , 2_n3955 , 2_n3956 , 2_n3957 , 2_n3958 , 2_n3959 , 2_n3960 , 2_n3961 , 2_n3962 , 2_n3963 , 2_n3964 , 2_n3965 , 2_n3966 , 2_n3967 , 2_n3968 , 2_n3969 , 2_n3970 , 2_n3971 , 2_n3972 , 2_n3973 , 2_n3974 , 2_n3975 , 2_n3976 , 2_n3977 , 2_n3978 , 2_n3979 , 2_n3980 , 2_n3981 , 2_n3982 , 2_n3983 , 2_n3984 , 2_n3985 , 2_n3987 , 2_n3988 , 2_n3989 , 2_n3990 , 2_n3991 , 2_n3993 , 2_n3994 , 2_n3995 , 2_n3996 , 2_n3997 , 2_n3998 , 2_n3999 , 2_n4000 , 2_n4001 , 2_n4002 , 2_n4003 , 2_n4004 , 2_n4006 , 2_n4007 , 2_n4008 , 2_n4009 , 2_n4010 , 2_n4011 , 2_n4012 , 2_n4013 , 2_n4014 , 2_n4015 , 2_n4016 , 2_n4017 , 2_n4018 , 2_n4019 , 2_n4020 , 2_n4021 , 2_n4022 , 2_n4023 , 2_n4024 , 2_n4025 , 2_n4026 , 2_n4027 , 2_n4028 , 2_n4029 , 2_n4030 , 2_n4031 , 2_n4032 , 2_n4033 , 2_n4034 , 2_n4035 , 2_n4036 , 2_n4037 , 2_n4038 , 2_n4039 , 2_n4040 , 2_n4041 , 2_n4042 , 2_n4043 , 2_n4044 , 2_n4045 , 2_n4046 , 2_n4047 , 2_n4048 , 2_n4049 , 2_n4050 , 2_n4051 , 2_n4052 , 2_n4053 , 2_n4054 , 2_n4055 , 2_n4056 , 2_n4057 , 2_n4058 , 2_n4059 , 2_n4060 , 2_n4061 , 2_n4062 , 2_n4063 , 2_n4064 , 2_n4065 , 2_n4066 , 2_n4067 , 2_n4068 , 2_n4069 , 2_n4070 , 2_n4071 , 2_n4072 , 2_n4073 , 2_n4074 , 2_n4075 , 2_n4076 , 2_n4077 , 2_n4078 , 2_n4079 , 2_n4080 , 2_n4081 , 2_n4082 , 2_n4083 , 2_n4084 , 2_n4085 , 2_n4087 , 2_n4089 , 2_n4090 , 2_n4091 , 2_n4092 , 2_n4093 , 2_n4095 , 2_n4096 , 2_n4097 , 2_n4098 , 2_n4099 , 2_n4100 , 2_n4101 , 2_n4102 , 2_n4103 , 2_n4104 , 2_n4105 , 2_n4106 , 2_n4107 , 2_n4108 , 2_n4109 , 2_n4110 , 2_n4111 , 2_n4112 , 2_n4113 , 2_n4114 , 2_n4115 , 2_n4116 , 2_n4117 , 2_n4118 , 2_n4119 , 2_n4120 , 2_n4121 , 2_n4122 , 2_n4123 , 2_n4124 , 2_n4125 , 2_n4126 , 2_n4127 , 2_n4128 , 2_n4129 , 2_n4130 , 2_n4131 , 2_n4132 , 2_n4133 , 2_n4134 , 2_n4135 , 2_n4136 , 2_n4137 , 2_n4138 , 2_n4139 , 2_n4140 , 2_n4142 , 2_n4143 , 2_n4144 , 2_n4145 , 2_n4146 , 2_n4147 , 2_n4148 , 2_n4149 , 2_n4150 , 2_n4151 , 2_n4152 , 2_n4153 , 2_n4154 , 2_n4156 , 2_n4157 , 2_n4158 , 2_n4160 , 2_n4161 , 2_n4162 , 2_n4163 , 2_n4164 , 2_n4165 , 2_n4166 , 2_n4167 , 2_n4168 , 2_n4169 , 2_n4170 , 2_n4171 , 2_n4172 , 2_n4173 , 2_n4174 , 2_n4175 , 2_n4176 , 2_n4177 , 2_n4178 , 2_n4179 , 2_n4180 , 2_n4181 , 2_n4182 , 2_n4183 , 2_n4184 , 2_n4185 , 2_n4186 , 2_n4188 , 2_n4191 , 2_n4192 , 2_n4193 , 2_n4194 , 2_n4195 , 2_n4196 , 2_n4197 , 2_n4198 , 2_n4199 , 2_n4200 , 2_n4201 , 2_n4202 , 2_n4204 , 2_n4205 , 2_n4206 , 2_n4207 , 2_n4208 , 2_n4209 , 2_n4210 , 2_n4211 , 2_n4212 , 2_n4213 , 2_n4214 , 2_n4215 , 2_n4216 , 2_n4217 , 2_n4218 , 2_n4219 , 2_n4220 , 2_n4221 , 2_n4222 , 2_n4223 , 2_n4224 , 2_n4225 , 2_n4227 , 2_n4228 , 2_n4229 , 2_n4231 , 2_n4232 , 2_n4233 , 2_n4234 , 2_n4235 , 2_n4236 , 2_n4237 , 2_n4238 , 2_n4239 , 2_n4240 , 2_n4241 , 2_n4242 , 2_n4243 , 2_n4244 , 2_n4245 , 2_n4246 , 2_n4247 , 2_n4248 , 2_n4249 , 2_n4250 , 2_n4251 , 2_n4252 , 2_n4253 , 2_n4254 , 2_n4255 , 2_n4256 , 2_n4257 , 2_n4258 , 2_n4259 , 2_n4260 , 2_n4261 , 2_n4262 , 2_n4263 , 2_n4264 , 2_n4265 , 2_n4266 , 2_n4267 , 2_n4268 , 2_n4269 , 2_n4270 , 2_n4271 , 2_n4272 , 2_n4273 , 2_n4274 , 2_n4275 , 2_n4276 , 2_n4277 , 2_n4278 , 2_n4279 , 2_n4280 , 2_n4281 , 2_n4282 , 2_n4283 , 2_n4284 , 2_n4285 , 2_n4286 , 2_n4287 , 2_n4288 , 2_n4289 , 2_n4290 , 2_n4291 , 2_n4292 , 2_n4293 , 2_n4294 , 2_n4295 , 2_n4296 , 2_n4297 , 2_n4298 , 2_n4299 , 2_n4301 , 2_n4302 , 2_n4303 , 2_n4304 , 2_n4305 , 2_n4306 , 2_n4307 , 2_n4308 , 2_n4309 , 2_n4310 , 2_n4311 , 2_n4313 , 2_n4314 , 2_n4315 , 2_n4316 , 2_n4317 , 2_n4318 , 2_n4319 , 2_n4320 , 2_n4321 , 2_n4322 , 2_n4323 , 2_n4324 , 2_n4325 , 2_n4327 , 2_n4328 , 2_n4329 , 2_n4330 , 2_n4331 , 2_n4332 , 2_n4334 , 2_n4335 , 2_n4336 , 2_n4337 , 2_n4338 , 2_n4339 , 2_n4340 , 2_n4341 , 2_n4342 , 2_n4343 , 2_n4344 , 2_n4345 , 2_n4346 , 2_n4347 , 2_n4348 , 2_n4349 , 2_n4350 , 2_n4351 , 2_n4352 , 2_n4353 , 2_n4354 , 2_n4355 , 2_n4356 , 2_n4357 , 2_n4358 , 2_n4359 , 2_n4360 , 2_n4361 , 2_n4362 , 2_n4363 , 2_n4364 , 2_n4365 , 2_n4366 , 2_n4367 , 2_n4368 , 2_n4369 , 2_n4371 , 2_n4372 , 2_n4373 , 2_n4374 , 2_n4375 , 2_n4376 , 2_n4377 , 2_n4379 , 2_n4380 , 2_n4381 , 2_n4382 , 2_n4383 , 2_n4384 , 2_n4385 , 2_n4386 , 2_n4387 , 2_n4388 , 2_n4389 , 2_n4390 , 2_n4391 , 2_n4392 , 2_n4393 , 2_n4394 , 2_n4395 , 2_n4396 , 2_n4398 , 2_n4399 , 2_n4400 , 2_n4401 , 2_n4402 , 2_n4403 , 2_n4404 , 2_n4405 , 2_n4406 , 2_n4407 , 2_n4408 , 2_n4409 , 2_n4410 , 2_n4411 , 2_n4412 , 2_n4413 , 2_n4414 , 2_n4415 , 2_n4416 , 2_n4417 , 2_n4418 , 2_n4419 , 2_n4420 , 2_n4421 , 2_n4422 , 2_n4423 , 2_n4424 , 2_n4425 , 2_n4426 , 2_n4427 , 2_n4428 , 2_n4429 , 2_n4430 , 2_n4431 , 2_n4432 , 2_n4433 , 2_n4434 , 2_n4435 , 2_n4437 , 2_n4438 , 2_n4439 , 2_n4440 , 2_n4441 , 2_n4442 , 2_n4443 , 2_n4444 , 2_n4445 , 2_n4446 , 2_n4447 , 2_n4448 , 2_n4449 , 2_n4450 , 2_n4451 , 2_n4452 , 2_n4453 , 2_n4454 , 2_n4455 , 2_n4456 , 2_n4457 , 2_n4458 , 2_n4459 , 2_n4460 , 2_n4461 , 2_n4462 , 2_n4463 , 2_n4464 , 2_n4465 , 2_n4466 , 2_n4467 , 2_n4468 , 2_n4469 , 2_n4470 , 2_n4471 , 2_n4472 , 2_n4473 , 2_n4474 , 2_n4475 , 2_n4476 , 2_n4477 , 2_n4478 , 2_n4479 , 2_n4480 , 2_n4481 , 2_n4482 , 2_n4483 , 2_n4484 , 2_n4485 , 2_n4486 , 2_n4487 , 2_n4488 , 2_n4489 , 2_n4490 , 2_n4491 , 2_n4492 , 2_n4493 , 2_n4494 , 2_n4495 , 2_n4496 , 2_n4497 , 2_n4498 , 2_n4500 , 2_n4501 , 2_n4502 , 2_n4503 , 2_n4504 , 2_n4505 , 2_n4506 , 2_n4507 , 2_n4508 , 2_n4509 , 2_n4510 , 2_n4511 , 2_n4512 , 2_n4513 , 2_n4514 , 2_n4515 , 2_n4517 , 2_n4518 , 2_n4519 , 2_n4520 , 2_n4521 , 2_n4522 , 2_n4523 , 2_n4524 , 2_n4525 , 2_n4526 , 2_n4527 , 2_n4528 , 2_n4529 , 2_n4530 , 2_n4531 , 2_n4532 , 2_n4533 , 2_n4534 , 2_n4535 , 2_n4536 , 2_n4537 , 2_n4538 , 2_n4539 , 2_n4540 , 2_n4541 , 2_n4542 , 2_n4543 , 2_n4544 , 2_n4545 , 2_n4546 , 2_n4547 , 2_n4548 , 2_n4549 , 2_n4550 , 2_n4551 , 2_n4552 , 2_n4554 , 2_n4555 , 2_n4556 , 2_n4557 , 2_n4558 , 2_n4559 , 2_n4560 , 2_n4561 , 2_n4562 , 2_n4563 , 2_n4564 , 2_n4565 , 2_n4566 , 2_n4567 , 2_n4568 , 2_n4569 , 2_n4570 , 2_n4571 , 2_n4572 , 2_n4573 , 2_n4574 , 2_n4575 , 2_n4576 , 2_n4577 , 2_n4578 , 2_n4579 , 2_n4580 , 2_n4581 , 2_n4582 , 2_n4583 , 2_n4584 , 2_n4585 , 2_n4586 , 2_n4587 , 2_n4588 , 2_n4589 , 2_n4590 , 2_n4591 , 2_n4592 , 2_n4593 , 2_n4594 , 2_n4595 , 2_n4596 , 2_n4597 , 2_n4598 , 2_n4599 , 2_n4600 , 2_n4601 , 2_n4602 , 2_n4603 , 2_n4604 , 2_n4605 , 2_n4606 , 2_n4607 , 2_n4608 , 2_n4609 , 2_n4610 , 2_n4611 , 2_n4612 , 2_n4613 , 2_n4614 , 2_n4615 , 2_n4616 , 2_n4617 , 2_n4618 , 2_n4619 , 2_n4620 , 2_n4621 , 2_n4622 , 2_n4623 , 2_n4624 , 2_n4625 , 2_n4626 , 2_n4627 , 2_n4628 , 2_n4629 , 2_n4630 , 2_n4631 , 2_n4632 , 2_n4633 , 2_n4635 , 2_n4636 , 2_n4637 , 2_n4638 , 2_n4639 , 2_n4640 , 2_n4641 , 2_n4642 , 2_n4643 , 2_n4644 , 2_n4645 , 2_n4646 , 2_n4647 , 2_n4648 , 2_n4649 , 2_n4650 , 2_n4651 , 2_n4652 , 2_n4653 , 2_n4654 , 2_n4655 , 2_n4656 , 2_n4657 , 2_n4658 , 2_n4659 , 2_n4660 , 2_n4661 , 2_n4662 , 2_n4663 , 2_n4664 , 2_n4665 , 2_n4666 , 2_n4667 , 2_n4668 , 2_n4669 , 2_n4670 , 2_n4671 , 2_n4672 , 2_n4673 , 2_n4674 , 2_n4675 , 2_n4676 , 2_n4677 , 2_n4678 , 2_n4679 , 2_n4680 , 2_n4681 , 2_n4682 , 2_n4683 , 2_n4684 , 2_n4685 , 2_n4687 , 2_n4688 , 2_n4690 , 2_n4691 , 2_n4692 , 2_n4693 , 2_n4694 , 2_n4695 , 2_n4696 , 2_n4697 , 2_n4698 , 2_n4699 , 2_n4700 , 2_n4701 , 2_n4702 , 2_n4703 , 2_n4704 , 2_n4705 , 2_n4706 , 2_n4707 , 2_n4708 , 2_n4709 , 2_n4710 , 2_n4711 , 2_n4712 , 2_n4713 , 2_n4714 , 2_n4715 , 2_n4716 , 2_n4717 , 2_n4718 , 2_n4719 , 2_n4720 , 2_n4721 , 2_n4723 , 2_n4724 , 2_n4725 , 2_n4726 , 2_n4727 , 2_n4728 , 2_n4729 , 2_n4730 , 2_n4731 , 2_n4732 , 2_n4734 , 2_n4735 , 2_n4736 , 2_n4737 , 2_n4738 , 2_n4739 , 2_n4740 , 2_n4741 , 2_n4742 , 2_n4743 , 2_n4744 , 2_n4745 , 2_n4746 , 2_n4747 , 2_n4748 , 2_n4749 , 2_n4750 , 2_n4751 , 2_n4752 , 2_n4753 , 2_n4754 , 2_n4755 , 2_n4756 , 2_n4758 , 2_n4759 , 2_n4760 , 2_n4761 , 2_n4762 , 2_n4763 , 2_n4764 , 2_n4765 , 2_n4766 , 2_n4767 , 2_n4768 , 2_n4769 , 2_n4770 , 2_n4771 , 2_n4772 , 2_n4773 , 2_n4774 , 2_n4775 , 2_n4776 , 2_n4777 , 2_n4778 , 2_n4779 , 2_n4780 , 2_n4781 , 2_n4782 , 2_n4783 , 2_n4784 , 2_n4785 , 2_n4786 , 2_n4787 , 2_n4788 , 2_n4789 , 2_n4790 , 2_n4791 , 2_n4792 , 2_n4793 , 2_n4794 , 2_n4795 , 2_n4796 , 2_n4797 , 2_n4798 , 2_n4799 , 2_n4800 , 2_n4801 , 2_n4802 , 2_n4803 , 2_n4804 , 2_n4806 , 2_n4807 , 2_n4808 , 2_n4809 , 2_n4810 , 2_n4811 , 2_n4812 , 2_n4813 , 2_n4814 , 2_n4815 , 2_n4816 , 2_n4818 , 2_n4819 , 2_n4820 , 2_n4821 , 2_n4822 , 2_n4823 , 2_n4824 , 2_n4825 , 2_n4827 , 2_n4829 , 2_n4830 , 2_n4831 , 2_n4832 , 2_n4833 , 2_n4834 , 2_n4835 , 2_n4836 , 2_n4837 , 2_n4838 , 2_n4839 , 2_n4840 , 2_n4841 , 2_n4842 , 2_n4843 , 2_n4844 , 2_n4845 , 2_n4846 , 2_n4847 , 2_n4848 , 2_n4849 , 2_n4850 , 2_n4851 , 2_n4852 , 2_n4853 , 2_n4854 , 2_n4855 , 2_n4856 , 2_n4857 , 2_n4858 , 2_n4859 , 2_n4860 , 2_n4861 , 2_n4862 , 2_n4863 , 2_n4864 , 2_n4865 , 2_n4866 , 2_n4867 , 2_n4868 , 2_n4869 , 2_n4870 , 2_n4871 , 2_n4872 , 2_n4873 , 2_n4874 , 2_n4875 , 2_n4876 , 2_n4877 , 2_n4878 , 2_n4879 , 2_n4880 , 2_n4881 , 2_n4882 , 2_n4883 , 2_n4884 , 2_n4885 , 2_n4886 , 2_n4887 , 2_n4888 , 2_n4889 , 2_n4890 , 2_n4891 , 2_n4892 , 2_n4893 , 2_n4894 , 2_n4895 , 2_n4896 , 2_n4897 , 2_n4898 , 2_n4899 , 2_n4900 , 2_n4901 , 2_n4902 , 2_n4904 , 2_n4905 , 2_n4906 , 2_n4907 , 2_n4908 , 2_n4909 , 2_n4910 , 2_n4911 , 2_n4912 , 2_n4913 , 2_n4914 , 2_n4915 , 2_n4916 , 2_n4917 , 2_n4918 , 2_n4919 , 2_n4920 , 2_n4922 , 2_n4923 , 2_n4924 , 2_n4925 , 2_n4926 , 2_n4927 , 2_n4929 , 2_n4930 , 2_n4931 , 2_n4932 , 2_n4933 , 2_n4934 , 2_n4935 , 2_n4936 , 2_n4937 , 2_n4939 , 2_n4940 , 2_n4941 , 2_n4942 , 2_n4943 , 2_n4944 , 2_n4945 , 2_n4946 , 2_n4947 , 2_n4948 , 2_n4949 , 2_n4950 , 2_n4951 , 2_n4952 , 2_n4953 , 2_n4954 , 2_n4955 , 2_n4956 , 2_n4957 , 2_n4958 , 2_n4959 , 2_n4960 , 2_n4961 , 2_n4962 , 2_n4963 , 2_n4964 , 2_n4965 , 2_n4966 , 2_n4967 , 2_n4968 , 2_n4969 , 2_n4972 , 2_n4973 , 2_n4974 , 2_n4975 , 2_n4976 , 2_n4977 , 2_n4978 , 2_n4979 , 2_n4980 , 2_n4981 , 2_n4982 , 2_n4983 , 2_n4984 , 2_n4985 , 2_n4986 , 2_n4987 , 2_n4988 , 2_n4989 , 2_n4990 , 2_n4991 , 2_n4992 , 2_n4993 , 2_n4994 , 2_n4995 , 2_n4996 , 2_n4997 , 2_n4998 , 2_n4999 , 2_n5000 , 2_n5001 , 2_n5002 , 2_n5003 , 2_n5004 , 2_n5005 , 2_n5006 , 2_n5007 , 2_n5008 , 2_n5009 , 2_n5010 , 2_n5011 , 2_n5012 , 2_n5013 , 2_n5014 , 2_n5015 , 2_n5016 , 2_n5017 , 2_n5018 , 2_n5019 , 2_n5020 , 2_n5021 , 2_n5022 , 2_n5023 , 2_n5024 , 2_n5025 , 2_n5026 , 2_n5027 , 2_n5028 , 2_n5029 , 2_n5031 , 2_n5032 , 2_n5033 , 2_n5035 , 2_n5036 , 2_n5037 , 2_n5038 , 2_n5039 , 2_n5040 , 2_n5041 , 2_n5042 , 2_n5043 , 2_n5044 , 2_n5045 , 2_n5046 , 2_n5047 , 2_n5048 , 2_n5049 , 2_n5050 , 2_n5051 , 2_n5052 , 2_n5053 , 2_n5054 , 2_n5055 , 2_n5056 , 2_n5057 , 2_n5058 , 2_n5059 , 2_n5060 , 2_n5061 , 2_n5062 , 2_n5063 , 2_n5064 , 2_n5065 , 2_n5066 , 2_n5067 , 2_n5068 , 2_n5070 , 2_n5071 , 2_n5072 , 2_n5073 , 2_n5074 , 2_n5075 , 2_n5076 , 2_n5077 , 2_n5078 , 2_n5079 , 2_n5080 , 2_n5081 , 2_n5082 , 2_n5083 , 2_n5084 , 2_n5085 , 2_n5086 , 2_n5087 , 2_n5088 , 2_n5089 , 2_n5090 , 2_n5091 , 2_n5092 , 2_n5093 , 2_n5095 , 2_n5096 , 2_n5097 , 2_n5098 , 2_n5099 , 2_n5100 , 2_n5101 , 2_n5102 , 2_n5103 , 2_n5104 , 2_n5106 , 2_n5107 , 2_n5108 , 2_n5109 , 2_n5110 , 2_n5111 , 2_n5112 , 2_n5113 , 2_n5114 , 2_n5115 , 2_n5116 , 2_n5117 , 2_n5118 , 2_n5119 , 2_n5120 , 2_n5121 , 2_n5122 , 2_n5123 , 2_n5124 , 2_n5125 , 2_n5126 , 2_n5127 , 2_n5128 , 2_n5129 , 2_n5130 , 2_n5131 , 2_n5133 , 2_n5134 , 2_n5135 , 2_n5136 , 2_n5137 , 2_n5138 , 2_n5139 , 2_n5140 , 2_n5141 , 2_n5142 , 2_n5143 , 2_n5144 , 2_n5145 , 2_n5146 , 2_n5147 , 2_n5148 , 2_n5149 , 2_n5150 , 2_n5151 , 2_n5152 , 2_n5154 , 2_n5155 , 2_n5156 , 2_n5157 , 2_n5158 , 2_n5159 , 2_n5160 , 2_n5161 , 2_n5162 , 2_n5163 , 2_n5164 , 2_n5165 , 2_n5166 , 2_n5167 , 2_n5168 , 2_n5169 , 2_n5170 , 2_n5171 , 2_n5172 , 2_n5173 , 2_n5174 , 2_n5175 , 2_n5176 , 2_n5177 , 2_n5178 , 2_n5179 , 2_n5180 , 2_n5181 , 2_n5182 , 2_n5183 , 2_n5184 , 2_n5185 , 2_n5186 , 2_n5187 , 2_n5188 , 2_n5189 , 2_n5190 , 2_n5192 , 2_n5193 , 2_n5194 , 2_n5195 , 2_n5196 , 2_n5197 , 2_n5199 , 2_n5200 , 2_n5201 , 2_n5202 , 2_n5203 , 2_n5204 , 2_n5205 , 2_n5206 , 2_n5207 , 2_n5208 , 2_n5209 , 2_n5210 , 2_n5211 , 2_n5213 , 2_n5214 , 2_n5215 , 2_n5216 , 2_n5217 , 2_n5218 , 2_n5219 , 2_n5220 , 2_n5221 , 2_n5222 , 2_n5223 , 2_n5224 , 2_n5225 , 2_n5226 , 2_n5227 , 2_n5228 , 2_n5229 , 2_n5230 , 2_n5231 , 2_n5232 , 2_n5233 , 2_n5234 , 2_n5235 , 2_n5236 , 2_n5237 , 2_n5238 , 2_n5239 , 2_n5241 , 2_n5242 , 2_n5243 , 2_n5244 , 2_n5245 , 2_n5246 , 2_n5247 , 2_n5248 , 2_n5249 , 2_n5250 , 2_n5251 , 2_n5252 , 2_n5253 , 2_n5254 , 2_n5255 , 2_n5256 , 2_n5258 , 2_n5259 , 2_n5260 , 2_n5261 , 2_n5262 , 2_n5263 , 2_n5264 , 2_n5265 , 2_n5266 , 2_n5267 , 2_n5268 , 2_n5269 , 2_n5270 , 2_n5271 , 2_n5272 , 2_n5273 , 2_n5274 , 2_n5275 , 2_n5276 , 2_n5277 , 2_n5278 , 2_n5279 , 2_n5280 , 2_n5281 , 2_n5282 , 2_n5284 , 2_n5285 , 2_n5286 , 2_n5287 , 2_n5288 , 2_n5289 , 2_n5290 , 2_n5291 , 2_n5292 , 2_n5293 , 2_n5294 , 2_n5295 , 2_n5296 , 2_n5297 , 2_n5298 , 2_n5299 , 2_n5300 , 2_n5301 , 2_n5302 , 2_n5303 , 2_n5304 , 2_n5306 , 2_n5307 , 2_n5308 , 2_n5309 , 2_n5310 , 2_n5311 , 2_n5312 , 2_n5313 , 2_n5315 , 2_n5316 , 2_n5317 , 2_n5318 , 2_n5321 , 2_n5322 , 2_n5323 , 2_n5324 , 2_n5325 , 2_n5326 , 2_n5327 , 2_n5328 , 2_n5329 , 2_n5330 , 2_n5332 , 2_n5333 , 2_n5334 , 2_n5335 , 2_n5336 , 2_n5337 , 2_n5338 , 2_n5339 , 2_n5340 , 2_n5341 , 2_n5342 , 2_n5343 , 2_n5344 , 2_n5345 , 2_n5346 , 2_n5347 , 2_n5348 , 2_n5349 , 2_n5350 , 2_n5351 , 2_n5352 , 2_n5353 , 2_n5354 , 2_n5355 , 2_n5356 , 2_n5357 , 2_n5358 , 2_n5359 , 2_n5360 , 2_n5361 , 2_n5362 , 2_n5363 , 2_n5364 , 2_n5365 , 2_n5366 , 2_n5367 , 2_n5368 , 2_n5369 , 2_n5370 , 2_n5371 , 2_n5372 , 2_n5373 , 2_n5374 , 2_n5375 , 2_n5376 , 2_n5377 , 2_n5378 , 2_n5379 , 2_n5380 , 2_n5381 , 2_n5382 , 2_n5383 , 2_n5384 , 2_n5385 , 2_n5386 , 2_n5387 , 2_n5388 , 2_n5389 , 2_n5390 , 2_n5391 , 2_n5392 , 2_n5393 , 2_n5394 , 2_n5395 , 2_n5396 , 2_n5397 , 2_n5398 , 2_n5399 , 2_n5400 , 2_n5401 , 2_n5402 , 2_n5403 , 2_n5404 , 2_n5405 , 2_n5406 , 2_n5407 , 2_n5408 , 2_n5409 , 2_n5410 , 2_n5412 , 2_n5413 , 2_n5414 , 2_n5415 , 2_n5416 , 2_n5417 , 2_n5418 , 2_n5419 , 2_n5420 , 2_n5421 , 2_n5422 , 2_n5423 , 2_n5424 , 2_n5425 , 2_n5426 , 2_n5427 , 2_n5428 , 2_n5429 , 2_n5430 , 2_n5431 , 2_n5432 , 2_n5433 , 2_n5434 , 2_n5436 , 2_n5437 , 2_n5438 , 2_n5439 , 2_n5440 , 2_n5441 , 2_n5442 , 2_n5443 , 2_n5444 , 2_n5445 , 2_n5446 , 2_n5447 , 2_n5448 , 2_n5449 , 2_n5450 , 2_n5451 , 2_n5452 , 2_n5453 , 2_n5454 , 2_n5455 , 2_n5456 , 2_n5457 , 2_n5458 , 2_n5459 , 2_n5460 , 2_n5461 , 2_n5462 , 2_n5463 , 2_n5464 , 2_n5465 , 2_n5466 , 2_n5467 , 2_n5468 , 2_n5469 , 2_n5470 , 2_n5471 , 2_n5472 , 2_n5473 , 2_n5474 , 2_n5475 , 2_n5476 , 2_n5477 , 2_n5478 , 2_n5479 , 2_n5480 , 2_n5481 , 2_n5482 , 2_n5483 , 2_n5484 , 2_n5485 , 2_n5486 , 2_n5487 , 2_n5488 , 2_n5489 , 2_n5490 , 2_n5491 , 2_n5492 , 2_n5493 , 2_n5494 , 2_n5495 , 2_n5496 , 2_n5497 , 2_n5498 , 2_n5499 , 2_n5500 , 2_n5501 , 2_n5502 , 2_n5503 , 2_n5504 , 2_n5505 , 2_n5506 , 2_n5507 , 2_n5508 , 2_n5509 , 2_n5510 , 2_n5511 , 2_n5512 , 2_n5513 , 2_n5514 , 2_n5515 , 2_n5516 , 2_n5517 , 2_n5518 , 2_n5519 , 2_n5520 , 2_n5521 , 2_n5522 , 2_n5523 , 2_n5524 , 2_n5525 , 2_n5526 , 2_n5527 , 2_n5528 , 2_n5529 , 2_n5530 , 2_n5531 , 2_n5532 , 2_n5533 , 2_n5534 , 2_n5535 , 2_n5536 , 2_n5537 , 2_n5538 , 2_n5539 , 2_n5540 , 2_n5541 , 2_n5542 , 2_n5543 , 2_n5544 , 2_n5545 , 2_n5546 , 2_n5547 , 2_n5548 , 2_n5549 , 2_n5550 , 2_n5551 , 2_n5552 , 2_n5553 , 2_n5554 , 2_n5555 , 2_n5556 , 2_n5557 , 2_n5558 , 2_n5559 , 2_n5560 , 2_n5561 , 2_n5562 , 2_n5563 , 2_n5564 , 2_n5565 , 2_n5566 , 2_n5567 , 2_n5568 , 2_n5569 , 2_n5570 , 2_n5571 , 2_n5572 , 2_n5573 , 2_n5574 , 2_n5575 , 2_n5576 , 2_n5577 , 2_n5578 , 2_n5580 , 2_n5581 , 2_n5582 , 2_n5583 , 2_n5584 , 2_n5585 , 2_n5586 , 2_n5587 , 2_n5588 , 2_n5589 , 2_n5590 , 2_n5591 , 2_n5592 , 2_n5593 , 2_n5594 , 2_n5595 , 2_n5596 , 2_n5597 , 2_n5598 , 2_n5599 , 2_n5600 , 2_n5601 , 2_n5602 , 2_n5603 , 2_n5604 , 2_n5605 , 2_n5606 , 2_n5607 , 2_n5608 , 2_n5609 , 2_n5610 , 2_n5611 , 2_n5612 , 2_n5613 , 2_n5614 , 2_n5615 , 2_n5616 , 2_n5617 , 2_n5618 , 2_n5619 , 2_n5620 , 2_n5621 , 2_n5622 , 2_n5623 , 2_n5624 , 2_n5625 , 2_n5626 , 2_n5627 , 2_n5628 , 2_n5629 , 2_n5630 , 2_n5631 , 2_n5632 , 2_n5633 , 2_n5634 , 2_n5635 , 2_n5636 , 2_n5637 , 2_n5638 , 2_n5639 , 2_n5640 , 2_n5642 , 2_n5643 , 2_n5644 , 2_n5646 , 2_n5647 , 2_n5648 , 2_n5649 , 2_n5650 , 2_n5651 , 2_n5652 , 2_n5653 , 2_n5654 , 2_n5655 , 2_n5656 , 2_n5657 , 2_n5658 , 2_n5659 , 2_n5660 , 2_n5661 , 2_n5662 , 2_n5663 , 2_n5664 , 2_n5665 , 2_n5666 , 2_n5667 , 2_n5668 , 2_n5669 , 2_n5671 , 2_n5672 , 2_n5673 , 2_n5674 , 2_n5675 , 2_n5676 , 2_n5677 , 2_n5678 , 2_n5679 , 2_n5680 , 2_n5681 , 2_n5682 , 2_n5683 , 2_n5684 , 2_n5685 , 2_n5686 , 2_n5687 , 2_n5688 , 2_n5689 , 2_n5690 , 2_n5691 , 2_n5692 , 2_n5695 , 2_n5696 , 2_n5697 , 2_n5698 , 2_n5699 , 2_n5700 , 2_n5701 , 2_n5702 , 2_n5703 , 2_n5704 , 2_n5705 , 2_n5706 , 2_n5707 , 2_n5708 , 2_n5709 , 2_n5710 , 2_n5711 , 2_n5712 , 2_n5713 , 2_n5714 , 2_n5715 , 2_n5716 , 2_n5717 , 2_n5718 , 2_n5719 , 2_n5720 , 2_n5721 , 2_n5722 , 2_n5723 , 2_n5724 , 2_n5725 , 2_n5726 , 2_n5727 , 2_n5728 , 2_n5729 , 2_n5730 , 2_n5731 , 2_n5732 , 2_n5733 , 2_n5734 , 2_n5735 , 2_n5736 , 2_n5737 , 2_n5738 , 2_n5739 , 2_n5740 , 2_n5741 , 2_n5742 , 2_n5743 , 2_n5744 , 2_n5745 , 2_n5746 , 2_n5747 , 2_n5748 , 2_n5749 , 2_n5750 , 2_n5751 , 2_n5752 , 2_n5753 , 2_n5754 , 2_n5755 , 2_n5756 , 2_n5757 , 2_n5758 , 2_n5759 , 2_n5761 , 2_n5762 , 2_n5763 , 2_n5764 , 2_n5765 , 2_n5766 , 2_n5768 , 2_n5769 , 2_n5770 , 2_n5771 , 2_n5772 , 2_n5773 , 2_n5774 , 2_n5775 , 2_n5776 , 2_n5777 , 2_n5778 , 2_n5779 , 2_n5780 , 2_n5781 , 2_n5782 , 2_n5783 , 2_n5784 , 2_n5785 , 2_n5786 , 2_n5787 , 2_n5788 , 2_n5789 , 2_n5790 , 2_n5791 , 2_n5792 , 2_n5793 , 2_n5794 , 2_n5795 , 2_n5796 , 2_n5797 , 2_n5799 , 2_n5800 , 2_n5801 , 2_n5802 , 2_n5803 , 2_n5804 , 2_n5805 , 2_n5806 , 2_n5807 , 2_n5808 , 2_n5809 , 2_n5810 , 2_n5811 , 2_n5812 , 2_n5813 , 2_n5815 , 2_n5816 , 2_n5817 , 2_n5818 , 2_n5819 , 2_n5820 , 2_n5821 , 2_n5822 , 2_n5823 , 2_n5824 , 2_n5825 , 2_n5826 , 2_n5827 , 2_n5828 , 2_n5829 , 2_n5830 , 2_n5831 , 2_n5832 , 2_n5833 , 2_n5834 , 2_n5835 , 2_n5836 , 2_n5837 , 2_n5838 , 2_n5839 , 2_n5840 , 2_n5841 , 2_n5842 , 2_n5843 , 2_n5844 , 2_n5845 , 2_n5846 , 2_n5847 , 2_n5848 , 2_n5849 , 2_n5850 , 2_n5851 , 2_n5852 , 2_n5853 , 2_n5854 , 2_n5855 , 2_n5856 , 2_n5858 , 2_n5859 , 2_n5861 , 2_n5862 , 2_n5863 , 2_n5864 , 2_n5865 , 2_n5866 , 2_n5867 , 2_n5868 , 2_n5869 , 2_n5870 , 2_n5871 , 2_n5872 , 2_n5873 , 2_n5874 , 2_n5875 , 2_n5876 , 2_n5877 , 2_n5878 , 2_n5879 , 2_n5880 , 2_n5881 , 2_n5882 , 2_n5883 , 2_n5884 , 2_n5885 , 2_n5886 , 2_n5887 , 2_n5888 , 2_n5889 , 2_n5890 , 2_n5891 , 2_n5892 , 2_n5893 , 2_n5894 , 2_n5895 , 2_n5896 , 2_n5897 , 2_n5898 , 2_n5899 , 2_n5900 , 2_n5901 , 2_n5902 , 2_n5903 , 2_n5904 , 2_n5905 , 2_n5906 , 2_n5907 , 2_n5908 , 2_n5909 , 2_n5910 , 2_n5911 , 2_n5912 , 2_n5913 , 2_n5914 , 2_n5915 , 2_n5916 , 2_n5917 , 2_n5918 , 2_n5919 , 2_n5920 , 2_n5921 , 2_n5922 , 2_n5923 , 2_n5924 , 2_n5925 , 2_n5926 , 2_n5927 , 2_n5928 , 2_n5929 , 2_n5930 , 2_n5931 , 2_n5932 , 2_n5933 , 2_n5935 , 2_n5936 , 2_n5937 , 2_n5938 , 2_n5939 , 2_n5940 , 2_n5941 , 2_n5942 , 2_n5943 , 2_n5944 , 2_n5945 , 2_n5946 , 2_n5947 , 2_n5948 , 2_n5949 , 2_n5950 , 2_n5951 , 2_n5952 , 2_n5953 , 2_n5954 , 2_n5955 , 2_n5956 , 2_n5957 , 2_n5958 , 2_n5959 , 2_n5960 , 2_n5961 , 2_n5962 , 2_n5963 , 2_n5965 , 2_n5966 , 2_n5967 , 2_n5968 , 2_n5969 , 2_n5970 , 2_n5971 , 2_n5972 , 2_n5973 , 2_n5974 , 2_n5975 , 2_n5976 , 2_n5977 , 2_n5978 , 2_n5979 , 2_n5980 , 2_n5981 , 2_n5982 , 2_n5983 , 2_n5984 , 2_n5985 , 2_n5986 , 2_n5987 , 2_n5988 , 2_n5989 , 2_n5990 , 2_n5991 , 2_n5992 , 2_n5993 , 2_n5994 , 2_n5995 , 2_n5996 , 2_n5997 , 2_n5998 , 2_n5999 , 2_n6000 , 2_n6001 , 2_n6002 , 2_n6003 , 2_n6004 , 2_n6005 , 2_n6006 , 2_n6007 , 2_n6008 , 2_n6009 , 2_n6010 , 2_n6011 , 2_n6012 , 2_n6013 , 2_n6014 , 2_n6015 , 2_n6017 , 2_n6018 , 2_n6019 , 2_n6020 , 2_n6021 , 2_n6022 , 2_n6023 , 2_n6024 , 2_n6025 , 2_n6026 , 2_n6027 , 2_n6028 , 2_n6029 , 2_n6030 , 2_n6031 , 2_n6032 , 2_n6033 , 2_n6034 , 2_n6035 , 2_n6036 , 2_n6037 , 2_n6039 , 2_n6040 , 2_n6041 , 2_n6042 , 2_n6043 , 2_n6044 , 2_n6045 , 2_n6046 , 2_n6047 , 2_n6048 , 2_n6049 , 2_n6050 , 2_n6051 , 2_n6052 , 2_n6053 , 2_n6054 , 2_n6055 , 2_n6056 , 2_n6057 , 2_n6058 , 2_n6059 , 2_n6060 , 2_n6061 , 2_n6062 , 2_n6063 , 2_n6064 , 2_n6065 , 2_n6066 , 2_n6067 , 2_n6068 , 2_n6069 , 2_n6070 , 2_n6071 , 2_n6072 , 2_n6073 , 2_n6074 , 2_n6075 , 2_n6076 , 2_n6077 , 2_n6078 , 2_n6079 , 2_n6080 , 2_n6081 , 2_n6082 , 2_n6083 , 2_n6084 , 2_n6085 , 2_n6086 , 2_n6087 , 2_n6088 , 2_n6090 , 2_n6091 , 2_n6092 , 2_n6093 , 2_n6094 , 2_n6095 , 2_n6096 , 2_n6097 , 2_n6098 , 2_n6099 , 2_n6100 , 2_n6101 , 2_n6102 , 2_n6103 , 2_n6104 , 2_n6105 , 2_n6106 , 2_n6107 , 2_n6108 , 2_n6109 , 2_n6110 , 2_n6111 , 2_n6112 , 2_n6113 , 2_n6114 , 2_n6115 , 2_n6116 , 2_n6117 , 2_n6118 , 2_n6119 , 2_n6120 , 2_n6121 , 2_n6122 , 2_n6123 , 2_n6124 , 2_n6125 , 2_n6127 , 2_n6128 , 2_n6129 , 2_n6130 , 2_n6131 , 2_n6132 , 2_n6133 , 2_n6134 , 2_n6135 , 2_n6136 , 2_n6137 , 2_n6138 , 2_n6139 , 2_n6140 , 2_n6141 , 2_n6142 , 2_n6143 , 2_n6144 , 2_n6145 , 2_n6146 , 2_n6147 , 2_n6148 , 2_n6149 , 2_n6150 , 2_n6151 , 2_n6152 , 2_n6153 , 2_n6154 , 2_n6155 , 2_n6156 , 2_n6157 , 2_n6158 , 2_n6159 , 2_n6160 , 2_n6161 , 2_n6162 , 2_n6163 , 2_n6164 , 2_n6165 , 2_n6166 , 2_n6167 , 2_n6168 , 2_n6169 , 2_n6170 , 2_n6171 , 2_n6172 , 2_n6173 , 2_n6174 , 2_n6175 , 2_n6176 , 2_n6177 , 2_n6178 , 2_n6179 , 2_n6180 , 2_n6181 , 2_n6182 , 2_n6183 , 2_n6184 , 2_n6185 , 2_n6186 , 2_n6187 , 2_n6188 , 2_n6189 , 2_n6190 , 2_n6191 , 2_n6193 , 2_n6194 , 2_n6195 , 2_n6196 , 2_n6197 , 2_n6198 , 2_n6199 , 2_n6200 , 2_n6201 , 2_n6202 , 2_n6203 , 2_n6204 , 2_n6205 , 2_n6206 , 2_n6207 , 2_n6208 , 2_n6209 , 2_n6210 , 2_n6211 , 2_n6212 , 2_n6213 , 2_n6214 , 2_n6215 , 2_n6216 , 2_n6217 , 2_n6218 , 2_n6219 , 2_n6220 , 2_n6221 , 2_n6222 , 2_n6223 , 2_n6224 , 2_n6225 , 2_n6226 , 2_n6227 , 2_n6228 , 2_n6229 , 2_n6230 , 2_n6231 , 2_n6232 , 2_n6233 , 2_n6234 , 2_n6235 , 2_n6236 , 2_n6237 , 2_n6238 , 2_n6239 , 2_n6240 , 2_n6241 , 2_n6242 , 2_n6243 , 2_n6244 , 2_n6245 , 2_n6246 , 2_n6247 , 2_n6248 , 2_n6249 , 2_n6250 , 2_n6251 , 2_n6252 , 2_n6253 , 2_n6255 , 2_n6256 , 2_n6257 , 2_n6258 , 2_n6259 , 2_n6260 , 2_n6261 , 2_n6262 , 2_n6263 , 2_n6264 , 2_n6265 , 2_n6266 , 2_n6267 , 2_n6268 , 2_n6269 , 2_n6270 , 2_n6271 , 2_n6272 , 2_n6274 , 2_n6275 , 2_n6276 , 2_n6277 , 2_n6278 , 2_n6279 , 2_n6280 , 2_n6281 , 2_n6282 , 2_n6283 , 2_n6284 , 2_n6285 , 2_n6286 , 2_n6287 , 2_n6288 , 2_n6289 , 2_n6290 , 2_n6291 , 2_n6292 , 2_n6293 , 2_n6295 , 2_n6296 , 2_n6297 , 2_n6298 , 2_n6299 , 2_n6300 , 2_n6301 , 2_n6302 , 2_n6303 , 2_n6304 , 2_n6305 , 2_n6306 , 2_n6307 , 2_n6308 , 2_n6309 , 2_n6310 , 2_n6311 , 2_n6312 , 2_n6313 , 2_n6314 , 2_n6315 , 2_n6316 , 2_n6317 , 2_n6318 , 2_n6319 , 2_n6320 , 2_n6321 , 2_n6322 , 2_n6323 , 2_n6324 , 2_n6325 , 2_n6326 , 2_n6327 , 2_n6328 , 2_n6329 , 2_n6330 , 2_n6331 , 2_n6332 , 2_n6333 , 2_n6334 , 2_n6335 , 2_n6336 , 2_n6337 , 2_n6338 , 2_n6339 , 2_n6340 , 2_n6341 , 2_n6342 , 2_n6343 , 2_n6344 , 2_n6345 , 2_n6346 , 2_n6347 , 2_n6348 , 2_n6349 , 2_n6350 , 2_n6351 , 2_n6352 , 2_n6353 , 2_n6354 , 2_n6355 , 2_n6356 , 2_n6357 , 2_n6360 , 2_n6361 , 2_n6362 , 2_n6363 , 2_n6364 , 2_n6365 , 2_n6366 , 2_n6367 , 2_n6368 , 2_n6369 , 2_n6370 , 2_n6371 , 2_n6372 , 2_n6373 , 2_n6374 , 2_n6375 , 2_n6376 , 2_n6377 , 2_n6378 , 2_n6379 , 2_n6380 , 2_n6381 , 2_n6382 , 2_n6383 , 2_n6384 , 2_n6385 , 2_n6386 , 2_n6387 , 2_n6388 , 2_n6389 , 2_n6390 , 2_n6391 , 2_n6392 , 2_n6393 , 2_n6394 , 2_n6395 , 2_n6396 , 2_n6397 , 2_n6398 , 2_n6399 , 2_n6400 , 2_n6401 , 2_n6402 , 2_n6403 , 2_n6404 , 2_n6405 , 2_n6406 , 2_n6407 , 2_n6408 , 2_n6409 , 2_n6410 , 2_n6411 , 2_n6412 , 2_n6413 , 2_n6414 , 2_n6415 , 2_n6416 , 2_n6417 , 2_n6418 , 2_n6419 , 2_n6420 , 2_n6421 , 2_n6422 , 2_n6423 , 2_n6424 , 2_n6425 , 2_n6426 , 2_n6427 , 2_n6428 , 2_n6430 , 2_n6432 , 2_n6433 , 2_n6434 , 2_n6435 , 2_n6436 , 2_n6437 , 2_n6438 , 2_n6439 , 2_n6440 , 2_n6442 , 2_n6443 , 2_n6444 , 2_n6446 , 2_n6447 , 2_n6448 , 2_n6449 , 2_n6450 , 2_n6451 , 2_n6452 , 2_n6453 , 2_n6454 , 2_n6455 , 2_n6456 , 2_n6457 , 2_n6458 , 2_n6459 , 2_n6460 , 2_n6461 , 2_n6462 , 2_n6463 , 2_n6464 , 2_n6465 , 2_n6466 , 2_n6467 , 2_n6468 , 2_n6469 , 2_n6470 , 2_n6471 , 2_n6472 , 2_n6473 , 2_n6474 , 2_n6475 , 2_n6476 , 2_n6477 , 2_n6478 , 2_n6479 , 2_n6480 , 2_n6481 , 2_n6482 , 2_n6483 , 2_n6484 , 2_n6485 , 2_n6486 , 2_n6487 , 2_n6488 , 2_n6489 , 2_n6490 , 2_n6491 , 2_n6492 , 2_n6493 , 2_n6494 , 2_n6495 , 2_n6496 , 2_n6497 , 2_n6498 , 2_n6499 , 2_n6500 , 2_n6501 , 2_n6502 , 2_n6503 , 2_n6504 , 2_n6505 , 2_n6506 , 2_n6507 , 2_n6508 , 2_n6509 , 2_n6510 , 2_n6511 , 2_n6512 , 2_n6513 , 2_n6514 , 2_n6515 , 2_n6516 , 2_n6517 , 2_n6518 , 2_n6519 , 2_n6520 , 2_n6521 , 2_n6522 , 2_n6523 , 2_n6524 , 2_n6525 , 2_n6526 , 2_n6527 , 2_n6528 , 2_n6529 , 2_n6530 , 2_n6531 , 2_n6532 , 2_n6533 , 2_n6534 , 2_n6535 , 2_n6536 , 2_n6537 , 2_n6538 , 2_n6539 , 2_n6540 , 2_n6541 , 2_n6542 , 2_n6543 , 2_n6544 , 2_n6545 , 2_n6546 , 2_n6547 , 2_n6548 , 2_n6549 , 2_n6550 , 2_n6551 , 2_n6552 , 2_n6553 , 2_n6554 , 2_n6555 , 2_n6556 , 2_n6557 , 2_n6558 , 2_n6559 , 2_n6560 , 2_n6561 , 2_n6562 , 2_n6563 , 2_n6564 , 2_n6565 , 2_n6566 , 2_n6567 , 2_n6568 , 2_n6569 , 2_n6570 , 2_n6571 , 2_n6572 , 2_n6573 , 2_n6574 , 2_n6575 , 2_n6576 , 2_n6577 , 2_n6579 , 2_n6580 , 2_n6581 , 2_n6582 , 2_n6583 , 2_n6584 , 2_n6585 , 2_n6586 , 2_n6587 , 2_n6588 , 2_n6589 , 2_n6590 , 2_n6591 , 2_n6592 , 2_n6593 , 2_n6594 , 2_n6595 , 2_n6596 , 2_n6597 , 2_n6598 , 2_n6599 , 2_n6600 , 2_n6601 , 2_n6602 , 2_n6603 , 2_n6605 , 2_n6606 , 2_n6607 , 2_n6608 , 2_n6609 , 2_n6610 , 2_n6612 , 2_n6613 , 2_n6614 , 2_n6615 , 2_n6616 , 2_n6617 , 2_n6618 , 2_n6619 , 2_n6620 , 2_n6621 , 2_n6622 , 2_n6623 , 2_n6624 , 2_n6625 , 2_n6626 , 2_n6627 , 2_n6628 , 2_n6629 , 2_n6630 , 2_n6631 , 2_n6632 , 2_n6633 , 2_n6634 , 2_n6635 , 2_n6636 , 2_n6637 , 2_n6638 , 2_n6639 , 2_n6640 , 2_n6641 , 2_n6642 , 2_n6643 , 2_n6644 , 2_n6646 , 2_n6647 , 2_n6648 , 2_n6649 , 2_n6650 , 2_n6651 , 2_n6652 , 2_n6653 , 2_n6654 , 2_n6655 , 2_n6656 , 2_n6657 , 2_n6658 , 2_n6659 , 2_n6660 , 2_n6661 , 2_n6662 , 2_n6663 , 2_n6664 , 2_n6665 , 2_n6666 , 2_n6667 , 2_n6668 , 2_n6669 , 2_n6670 , 2_n6671 , 2_n6672 , 2_n6673 , 2_n6674 , 2_n6675 , 2_n6676 , 2_n6677 , 2_n6678 , 2_n6679 , 2_n6680 , 2_n6681 , 2_n6682 , 2_n6683 , 2_n6684 , 2_n6685 , 2_n6686 , 2_n6688 , 2_n6690 , 2_n6691 , 2_n6692 , 2_n6693 , 2_n6694 , 2_n6695 , 2_n6696 , 2_n6697 , 2_n6698 , 2_n6699 , 2_n6700 , 2_n6701 , 2_n6702 , 2_n6704 , 2_n6705 , 2_n6706 , 2_n6707 , 2_n6708 , 2_n6709 , 2_n6710 , 2_n6711 , 2_n6712 , 2_n6713 , 2_n6714 , 2_n6715 , 2_n6716 , 2_n6717 , 2_n6718 , 2_n6719 , 2_n6720 , 2_n6721 , 2_n6722 , 2_n6723 , 2_n6724 , 2_n6725 , 2_n6726 , 2_n6727 , 2_n6728 , 2_n6729 , 2_n6730 , 2_n6731 , 2_n6732 , 2_n6733 , 2_n6734 , 2_n6735 , 2_n6736 , 2_n6737 , 2_n6738 , 2_n6739 , 2_n6740 , 2_n6741 , 2_n6743 , 2_n6744 , 2_n6745 , 2_n6746 , 2_n6747 , 2_n6748 , 2_n6749 , 2_n6750 , 2_n6751 , 2_n6752 , 2_n6753 , 2_n6754 , 2_n6755 , 2_n6756 , 2_n6757 , 2_n6758 , 2_n6759 , 2_n6760 , 2_n6761 , 2_n6762 , 2_n6763 , 2_n6764 , 2_n6765 , 2_n6766 , 2_n6767 , 2_n6768 , 2_n6769 , 2_n6771 , 2_n6772 , 2_n6773 , 2_n6774 , 2_n6775 , 2_n6777 , 2_n6778 , 2_n6779 , 2_n6780 , 2_n6781 , 2_n6782 , 2_n6783 , 2_n6784 , 2_n6785 , 2_n6786 , 2_n6787 , 2_n6788 , 2_n6789 , 2_n6790 , 2_n6791 , 2_n6792 , 2_n6793 , 2_n6794 , 2_n6795 , 2_n6796 , 2_n6798 , 2_n6799 , 2_n6800 , 2_n6801 , 2_n6802 , 2_n6803 , 2_n6804 , 2_n6805 , 2_n6807 , 2_n6808 , 2_n6810 , 2_n6811 , 2_n6812 , 2_n6813 , 2_n6814 , 2_n6815 , 2_n6816 , 2_n6817 , 2_n6818 , 2_n6819 , 2_n6820 , 2_n6821 , 2_n6823 , 2_n6824 , 2_n6825 , 2_n6827 , 2_n6828 , 2_n6829 , 2_n6830 , 2_n6831 , 2_n6832 , 2_n6833 , 2_n6834 , 2_n6835 , 2_n6836 , 2_n6837 , 2_n6838 , 2_n6839 , 2_n6840 , 2_n6841 , 2_n6842 , 2_n6843 , 2_n6844 , 2_n6845 , 2_n6846 , 2_n6847 , 2_n6848 , 2_n6849 , 2_n6850 , 2_n6851 , 2_n6852 , 2_n6853 , 2_n6854 , 2_n6855 , 2_n6856 , 2_n6857 , 2_n6858 , 2_n6859 , 2_n6861 , 2_n6862 , 2_n6863 , 2_n6864 , 2_n6865 , 2_n6866 , 2_n6867 , 2_n6868 , 2_n6869 , 2_n6870 , 2_n6871 , 2_n6872 , 2_n6873 , 2_n6874 , 2_n6875 , 2_n6876 , 2_n6878 , 2_n6879 , 2_n6880 , 2_n6881 , 2_n6882 , 2_n6883 , 2_n6884 , 2_n6885 , 2_n6886 , 2_n6887 , 2_n6888 , 2_n6889 , 2_n6890 , 2_n6891 , 2_n6892 , 2_n6893 , 2_n6894 , 2_n6895 , 2_n6896 , 2_n6897 , 2_n6898 , 2_n6899 , 2_n6900 , 2_n6901 , 2_n6902 , 2_n6903 , 2_n6904 , 2_n6905 , 2_n6906 , 2_n6907 , 2_n6908 , 2_n6909 , 2_n6910 , 2_n6911 , 2_n6912 , 2_n6913 , 2_n6914 , 2_n6915 , 2_n6916 , 2_n6917 , 2_n6918 , 2_n6919 , 2_n6920 , 2_n6921 , 2_n6922 , 2_n6923 , 2_n6924 , 2_n6925 , 2_n6926 , 2_n6927 , 2_n6928 , 2_n6929 , 2_n6930 , 2_n6931 , 2_n6932 , 2_n6933 , 2_n6934 , 2_n6935 , 2_n6936 , 2_n6937 , 2_n6938 , 2_n6939 , 2_n6940 , 2_n6941 , 2_n6942 , 2_n6943 , 2_n6944 , 2_n6945 , 2_n6946 , 2_n6947 , 2_n6948 , 2_n6949 , 2_n6950 , 2_n6951 , 2_n6952 , 2_n6953 , 2_n6954 , 2_n6955 , 2_n6956 , 2_n6957 , 2_n6958 , 2_n6959 , 2_n6960 , 2_n6961 , 2_n6962 , 2_n6963 , 2_n6964 , 2_n6965 , 2_n6966 , 2_n6967 , 2_n6968 , 2_n6969 , 2_n6970 , 2_n6971 , 2_n6972 , 2_n6973 , 2_n6974 , 2_n6975 , 2_n6976 , 2_n6977 , 2_n6978 , 2_n6979 , 2_n6980 , 2_n6981 , 2_n6982 , 2_n6983 , 2_n6984 , 2_n6985 , 2_n6987 , 2_n6988 , 2_n6989 , 2_n6990 , 2_n6991 , 2_n6992 , 2_n6993 , 2_n6994 , 2_n6995 , 2_n6996 , 2_n6997 , 2_n6998 , 2_n6999 , 2_n7000 , 2_n7001 , 2_n7002 , 2_n7003 , 2_n7004 , 2_n7005 , 2_n7006 , 2_n7007 , 2_n7008 , 2_n7009 , 2_n7010 , 2_n7011 , 2_n7012 , 2_n7013 , 2_n7014 , 2_n7015 , 2_n7016 , 2_n7017 , 2_n7018 , 2_n7019 , 2_n7020 , 2_n7021 , 2_n7022 , 2_n7023 , 2_n7024 , 2_n7025 , 2_n7026 , 2_n7027 , 2_n7028 , 2_n7029 , 2_n7030 , 2_n7031 , 2_n7032 , 2_n7033 , 2_n7034 , 2_n7035 , 2_n7036 , 2_n7037 , 2_n7038 , 2_n7039 , 2_n7040 , 2_n7041 , 2_n7042 , 2_n7043 , 2_n7044 , 2_n7045 , 2_n7046 , 2_n7047 , 2_n7048 , 2_n7049 , 2_n7050 , 2_n7051 , 2_n7052 , 2_n7053 , 2_n7054 , 2_n7055 , 2_n7056 , 2_n7057 , 2_n7058 , 2_n7059 , 2_n7060 , 2_n7061 , 2_n7062 , 2_n7063 , 2_n7064 , 2_n7065 , 2_n7066 , 2_n7067 , 2_n7068 , 2_n7069 , 2_n7070 , 2_n7071 , 2_n7072 , 2_n7073 , 2_n7074 , 2_n7075 , 2_n7076 , 2_n7077 , 2_n7078 , 2_n7079 , 2_n7080 , 2_n7081 , 2_n7082 , 2_n7083 , 2_n7084 , 2_n7085 , 2_n7086 , 2_n7087 , 2_n7088 , 2_n7089 , 2_n7090 , 2_n7091 , 2_n7092 , 2_n7093 , 2_n7094 , 2_n7095 , 2_n7096 , 2_n7097 , 2_n7098 , 2_n7099 , 2_n7100 , 2_n7101 , 2_n7102 , 2_n7103 , 2_n7104 , 2_n7105 , 2_n7106 , 2_n7107 , 2_n7108 , 2_n7109 , 2_n7110 , 2_n7111 , 2_n7112 , 2_n7113 , 2_n7114 , 2_n7115 , 2_n7116 , 2_n7117 , 2_n7118 , 2_n7119 , 2_n7120 , 2_n7121 , 2_n7122 , 2_n7123 , 2_n7124 , 2_n7125 , 2_n7126 , 2_n7127 , 2_n7128 , 2_n7129 , 2_n7130 , 2_n7131 , 2_n7132 , 2_n7133 , 2_n7134 , 2_n7135 , 2_n7136 , 2_n7137 , 2_n7138 , 2_n7139 , 2_n7140 , 2_n7141 , 2_n7142 , 2_n7143 , 2_n7144 , 2_n7145 , 2_n7146 , 2_n7147 , 2_n7148 , 2_n7149 , 2_n7150 , 2_n7151 , 2_n7152 , 2_n7153 , 2_n7154 , 2_n7155 , 2_n7156 , 2_n7157 , 2_n7158 , 2_n7161 , 2_n7162 , 2_n7163 , 2_n7164 , 2_n7165 , 2_n7166 , 2_n7167 , 2_n7168 , 2_n7169 , 2_n7170 , 2_n7171 , 2_n7172 , 2_n7173 , 2_n7174 , 2_n7175 , 2_n7176 , 2_n7177 , 2_n7178 , 2_n7179 , 2_n7180 , 2_n7181 , 2_n7182 , 2_n7183 , 2_n7184 , 2_n7185 , 2_n7186 , 2_n7187 , 2_n7188 , 2_n7189 , 2_n7190 , 2_n7191 , 2_n7192 , 2_n7194 , 2_n7195 , 2_n7196 , 2_n7197 , 2_n7198 , 2_n7199 , 2_n7200 , 2_n7201 , 2_n7202 , 2_n7203 , 2_n7204 , 2_n7205 , 2_n7206 , 2_n7207 , 2_n7208 , 2_n7209 , 2_n7210 , 2_n7211 , 2_n7212 , 2_n7213 , 2_n7214 , 2_n7215 , 2_n7216 , 2_n7217 , 2_n7218 , 2_n7219 , 2_n7220 , 2_n7221 , 2_n7222 , 2_n7223 , 2_n7224 , 2_n7225 , 2_n7226 , 2_n7227 , 2_n7228 , 2_n7229 , 2_n7230 , 2_n7231 , 2_n7232 , 2_n7233 , 2_n7234 , 2_n7235 , 2_n7237 , 2_n7238 , 2_n7239 , 2_n7240 , 2_n7241 , 2_n7242 , 2_n7243 , 2_n7244 , 2_n7245 , 2_n7246 , 2_n7247 , 2_n7248 , 2_n7249 , 2_n7250 , 2_n7251 , 2_n7252 , 2_n7253 , 2_n7254 , 2_n7255 , 2_n7256 , 2_n7257 , 2_n7258 , 2_n7259 , 2_n7260 , 2_n7261 , 2_n7262 , 2_n7263 , 2_n7264 , 2_n7266 , 2_n7267 , 2_n7268 , 2_n7269 , 2_n7271 , 2_n7272 , 2_n7273 , 2_n7274 , 2_n7275 , 2_n7276 , 2_n7277 , 2_n7278 , 2_n7279 , 2_n7280 , 2_n7281 , 2_n7282 , 2_n7283 , 2_n7284 , 2_n7285 , 2_n7286 , 2_n7287 , 2_n7288 , 2_n7289 , 2_n7290 , 2_n7291 , 2_n7292 , 2_n7293 , 2_n7295 , 2_n7296 , 2_n7297 , 2_n7298 , 2_n7299 , 2_n7300 , 2_n7301 , 2_n7302 , 2_n7303 , 2_n7304 , 2_n7305 , 2_n7306 , 2_n7307 , 2_n7308 , 2_n7309 , 2_n7310 , 2_n7311 , 2_n7312 , 2_n7313 , 2_n7314 , 2_n7315 , 2_n7316 , 2_n7317 , 2_n7318 , 2_n7319 , 2_n7321 , 2_n7322 , 2_n7323 , 2_n7324 , 2_n7325 , 2_n7326 , 2_n7327 , 2_n7328 , 2_n7329 , 2_n7330 , 2_n7331 , 2_n7332 , 2_n7333 , 2_n7334 , 2_n7335 , 2_n7336 , 2_n7337 , 2_n7338 , 2_n7339 , 2_n7340 , 2_n7341 , 2_n7342 , 2_n7343 , 2_n7344 , 2_n7345 , 2_n7346 , 2_n7347 , 2_n7348 , 2_n7349 , 2_n7350 , 2_n7351 , 2_n7352 , 2_n7353 , 2_n7355 , 2_n7356 , 2_n7357 , 2_n7358 , 2_n7359 , 2_n7360 , 2_n7361 , 2_n7362 , 2_n7363 , 2_n7364 , 2_n7365 , 2_n7366 , 2_n7367 , 2_n7368 , 2_n7369 , 2_n7370 , 2_n7371 , 2_n7372 , 2_n7373 , 2_n7374 , 2_n7375 , 2_n7376 , 2_n7377 , 2_n7378 , 2_n7379 , 2_n7380 , 2_n7381 , 2_n7382 , 2_n7383 , 2_n7384 , 2_n7385 , 2_n7386 , 2_n7387 , 2_n7389 , 2_n7390 , 2_n7391 , 2_n7392 , 2_n7393 , 2_n7394 , 2_n7395 , 2_n7396 , 2_n7397 , 2_n7398 , 2_n7399 , 2_n7400 , 2_n7401 , 2_n7402 , 2_n7403 , 2_n7404 , 2_n7405 , 2_n7406 , 2_n7407 , 2_n7408 , 2_n7409 , 2_n7410 , 2_n7411 , 2_n7412 , 2_n7413 , 2_n7414 , 2_n7415 , 2_n7416 , 2_n7417 , 2_n7418 , 2_n7419 , 2_n7420 , 2_n7421 , 2_n7422 , 2_n7423 , 2_n7424 , 2_n7425 , 2_n7426 , 2_n7427 , 2_n7428 , 2_n7429 , 2_n7430 , 2_n7431 , 2_n7432 , 2_n7433 , 2_n7434 , 2_n7435 , 2_n7437 , 2_n7438 , 2_n7439 , 2_n7440 , 2_n7441 , 2_n7442 , 2_n7443 , 2_n7444 , 2_n7445 , 2_n7446 , 2_n7447 , 2_n7448 , 2_n7449 , 2_n7450 , 2_n7451 , 2_n7452 , 2_n7453 , 2_n7454 , 2_n7455 , 2_n7457 , 2_n7458 , 2_n7459 , 2_n7460 , 2_n7461 , 2_n7462 , 2_n7463 , 2_n7464 , 2_n7465 , 2_n7466 , 2_n7467 , 2_n7468 , 2_n7469 , 2_n7470 , 2_n7471 , 2_n7472 , 2_n7473 , 2_n7474 , 2_n7475 , 2_n7476 , 2_n7477 , 2_n7478 , 2_n7479 , 2_n7480 , 2_n7481 , 2_n7482 , 2_n7483 , 2_n7484 , 2_n7485 , 2_n7486 , 2_n7487 , 2_n7488 , 2_n7489 , 2_n7490 , 2_n7491 , 2_n7492 , 2_n7493 , 2_n7494 , 2_n7495 , 2_n7496 , 2_n7497 , 2_n7498 , 2_n7499 , 2_n7501 , 2_n7502 , 2_n7503 , 2_n7504 , 2_n7505 , 2_n7506 , 2_n7507 , 2_n7508 , 2_n7509 , 2_n7510 , 2_n7511 , 2_n7512 , 2_n7513 , 2_n7514 , 2_n7515 , 2_n7516 , 2_n7517 , 2_n7518 , 2_n7519 , 2_n7520 , 2_n7521 , 2_n7522 , 2_n7524 , 2_n7525 , 2_n7526 , 2_n7527 , 2_n7528 , 2_n7529 , 2_n7530 , 2_n7531 , 2_n7532 , 2_n7533 , 2_n7534 , 2_n7535 , 2_n7536 , 2_n7537 , 2_n7538 , 2_n7539 , 2_n7540 , 2_n7541 , 2_n7542 , 2_n7543 , 2_n7544 , 2_n7545 , 2_n7547 , 2_n7548 , 2_n7549 , 2_n7550 , 2_n7551 , 2_n7552 , 2_n7553 , 2_n7554 , 2_n7555 , 2_n7556 , 2_n7557 , 2_n7558 , 2_n7559 , 2_n7560 , 2_n7561 , 2_n7562 , 2_n7563 , 2_n7564 , 2_n7565 , 2_n7566 , 2_n7567 , 2_n7569 , 2_n7570 , 2_n7571 , 2_n7572 , 2_n7573 , 2_n7574 , 2_n7575 , 2_n7576 , 2_n7577 , 2_n7578 , 2_n7579 , 2_n7580 , 2_n7581 , 2_n7582 , 2_n7583 , 2_n7584 , 2_n7585 , 2_n7586 , 2_n7587 , 2_n7588 , 2_n7589 , 2_n7590 , 2_n7591 , 2_n7592 , 2_n7593 , 2_n7594 , 2_n7595 , 2_n7596 , 2_n7597 , 2_n7598 , 2_n7599 , 2_n7600 , 2_n7601 , 2_n7602 , 2_n7603 , 2_n7604 , 2_n7605 , 2_n7606 , 2_n7607 , 2_n7608 , 2_n7609 , 2_n7611 , 2_n7612 , 2_n7613 , 2_n7614 , 2_n7615 , 2_n7616 , 2_n7617 , 2_n7618 , 2_n7619 , 2_n7620 , 2_n7621 , 2_n7622 , 2_n7623 , 2_n7624 , 2_n7625 , 2_n7626 , 2_n7627 , 2_n7628 , 2_n7629 , 2_n7630 , 2_n7631 , 2_n7632 , 2_n7633 , 2_n7634 , 2_n7635 , 2_n7636 , 2_n7637 , 2_n7638 , 2_n7639 , 2_n7640 , 2_n7641 , 2_n7642 , 2_n7643 , 2_n7644 , 2_n7645 , 2_n7647 , 2_n7648 , 2_n7649 , 2_n7650 , 2_n7651 , 2_n7652 , 2_n7653 , 2_n7654 , 2_n7655 , 2_n7656 , 2_n7657 , 2_n7658 , 2_n7659 , 2_n7660 , 2_n7661 , 2_n7662 , 2_n7663 , 2_n7664 , 2_n7665 , 2_n7666 , 2_n7667 , 2_n7668 , 2_n7669 , 2_n7670 , 2_n7671 , 2_n7672 , 2_n7673 , 2_n7674 , 2_n7675 , 2_n7677 , 2_n7678 , 2_n7679 , 2_n7680 , 2_n7681 , 2_n7682 , 2_n7683 , 2_n7684 , 2_n7685 , 2_n7686 , 2_n7687 , 2_n7688 , 2_n7689 , 2_n7691 , 2_n7692 , 2_n7693 , 2_n7694 , 2_n7695 , 2_n7696 , 2_n7697 , 2_n7698 , 2_n7699 , 2_n7700 , 2_n7701 , 2_n7702 , 2_n7703 , 2_n7704 , 2_n7705 , 2_n7706 , 2_n7707 , 2_n7708 , 2_n7709 , 2_n7710 , 2_n7711 , 2_n7712 , 2_n7713 , 2_n7714 , 2_n7715 , 2_n7716 , 2_n7717 , 2_n7718 , 2_n7719 , 2_n7720 , 2_n7721 , 2_n7722 , 2_n7723 , 2_n7724 , 2_n7725 , 2_n7726 , 2_n7727 , 2_n7728 , 2_n7729 , 2_n7731 , 2_n7732 , 2_n7734 , 2_n7735 , 2_n7736 , 2_n7737 , 2_n7738 , 2_n7739 , 2_n7740 , 2_n7741 , 2_n7742 , 2_n7743 , 2_n7744 , 2_n7745 , 2_n7746 , 2_n7747 , 2_n7748 , 2_n7749 , 2_n7750 , 2_n7751 , 2_n7752 , 2_n7753 , 2_n7754 , 2_n7755 , 2_n7756 , 2_n7757 , 2_n7758 , 2_n7759 , 2_n7760 , 2_n7761 , 2_n7762 , 2_n7763 , 2_n7764 , 2_n7765 , 2_n7766 , 2_n7767 , 2_n7768 , 2_n7769 , 2_n7770 , 2_n7771 , 2_n7772 , 2_n7773 , 2_n7774 , 2_n7775 , 2_n7776 , 2_n7777 , 2_n7778 , 2_n7779 , 2_n7780 , 2_n7781 , 2_n7782 , 2_n7783 , 2_n7784 , 2_n7785 , 2_n7786 , 2_n7787 , 2_n7788 , 2_n7789 , 2_n7790 , 2_n7791 , 2_n7792 , 2_n7793 , 2_n7794 , 2_n7795 , 2_n7796 , 2_n7797 , 2_n7798 , 2_n7799 , 2_n7800 , 2_n7801 , 2_n7802 , 2_n7803 , 2_n7804 , 2_n7805 , 2_n7806 , 2_n7807 , 2_n7808 , 2_n7809 , 2_n7810 , 2_n7811 , 2_n7812 , 2_n7813 , 2_n7814 , 2_n7815 , 2_n7816 , 2_n7817 , 2_n7818 , 2_n7819 , 2_n7820 , 2_n7821 , 2_n7822 , 2_n7824 , 2_n7825 , 2_n7826 , 2_n7827 , 2_n7828 , 2_n7829 , 2_n7830 , 2_n7831 , 2_n7832 , 2_n7833 , 2_n7834 , 2_n7835 , 2_n7836 , 2_n7837 , 2_n7838 , 2_n7839 , 2_n7840 , 2_n7841 , 2_n7842 , 2_n7843 , 2_n7844 , 2_n7845 , 2_n7846 , 2_n7847 , 2_n7848 , 2_n7849 , 2_n7850 , 2_n7851 , 2_n7852 , 2_n7853 , 2_n7854 , 2_n7855 , 2_n7856 , 2_n7857 , 2_n7858 , 2_n7859 , 2_n7860 , 2_n7861 , 2_n7863 , 2_n7864 , 2_n7865 , 2_n7866 , 2_n7867 , 2_n7868 , 2_n7869 , 2_n7870 , 2_n7871 , 2_n7872 , 2_n7873 , 2_n7874 , 2_n7875 , 2_n7876 , 2_n7877 , 2_n7878 , 2_n7879 , 2_n7880 , 2_n7881 , 2_n7882 , 2_n7883 , 2_n7884 , 2_n7885 , 2_n7886 , 2_n7887 , 2_n7888 , 2_n7889 , 2_n7890 , 2_n7892 , 2_n7893 , 2_n7894 , 2_n7895 , 2_n7896 , 2_n7897 , 2_n7898 , 2_n7899 , 2_n7900 , 2_n7901 , 2_n7902 , 2_n7903 , 2_n7904 , 2_n7905 , 2_n7906 , 2_n7907 , 2_n7908 , 2_n7909 , 2_n7910 , 2_n7911 , 2_n7912 , 2_n7913 , 2_n7914 , 2_n7915 , 2_n7916 , 2_n7917 , 2_n7918 , 2_n7919 , 2_n7920 , 2_n7921 , 2_n7922 , 2_n7923 , 2_n7924 , 2_n7925 , 2_n7926 , 2_n7927 , 2_n7928 , 2_n7929 , 2_n7930 , 2_n7931 , 2_n7932 , 2_n7933 , 2_n7934 , 2_n7935 , 2_n7936 , 2_n7937 , 2_n7938 , 2_n7939 , 2_n7940 , 2_n7941 , 2_n7942 , 2_n7943 , 2_n7944 , 2_n7945 , 2_n7947 , 2_n7948 , 2_n7949 , 2_n7950 , 2_n7951 , 2_n7952 , 2_n7953 , 2_n7954 , 2_n7955 , 2_n7956 , 2_n7957 , 2_n7958 , 2_n7959 , 2_n7960 , 2_n7961 , 2_n7962 , 2_n7963 , 2_n7964 , 2_n7967 , 2_n7968 , 2_n7969 , 2_n7970 , 2_n7971 , 2_n7972 , 2_n7973 , 2_n7974 , 2_n7975 , 2_n7976 , 2_n7977 , 2_n7978 , 2_n7979 , 2_n7980 , 2_n7982 , 2_n7983 , 2_n7984 , 2_n7985 , 2_n7986 , 2_n7987 , 2_n7988 , 2_n7989 , 2_n7990 , 2_n7991 , 2_n7992 , 2_n7993 , 2_n7994 , 2_n7995 , 2_n7996 , 2_n7997 , 2_n7998 , 2_n7999 , 2_n8000 , 2_n8001 , 2_n8002 , 2_n8003 , 2_n8004 , 2_n8005 , 2_n8006 , 2_n8007 , 2_n8008 , 2_n8009 , 2_n8010 , 2_n8011 , 2_n8012 , 2_n8013 , 2_n8014 , 2_n8015 , 2_n8016 , 2_n8017 , 2_n8018 , 2_n8019 , 2_n8020 , 2_n8021 , 2_n8022 , 2_n8023 , 2_n8024 , 2_n8025 , 2_n8026 , 2_n8027 , 2_n8029 , 2_n8030 , 2_n8031 , 2_n8032 , 2_n8033 , 2_n8034 , 2_n8035 , 2_n8036 , 2_n8037 , 2_n8038 , 2_n8039 , 2_n8040 , 2_n8041 , 2_n8042 , 2_n8043 , 2_n8044 , 2_n8045 , 2_n8046 , 2_n8047 , 2_n8048 , 2_n8049 , 2_n8050 , 2_n8051 , 2_n8052 , 2_n8053 , 2_n8054 , 2_n8055 , 2_n8056 , 2_n8057 , 2_n8058 , 2_n8059 , 2_n8060 , 2_n8061 , 2_n8062 , 2_n8063 , 2_n8064 , 2_n8066 , 2_n8067 , 2_n8068 , 2_n8069 , 2_n8070 , 2_n8071 , 2_n8072 , 2_n8073 , 2_n8074 , 2_n8075 , 2_n8076 , 2_n8077 , 2_n8078 , 2_n8079 , 2_n8080 , 2_n8081 , 2_n8082 , 2_n8083 , 2_n8084 , 2_n8085 , 2_n8086 , 2_n8087 , 2_n8088 , 2_n8089 , 2_n8090 , 2_n8091 , 2_n8092 , 2_n8093 , 2_n8094 , 2_n8095 , 2_n8096 , 2_n8097 , 2_n8098 , 2_n8099 , 2_n8101 , 2_n8102 , 2_n8103 , 2_n8104 , 2_n8105 , 2_n8106 , 2_n8107 , 2_n8108 , 2_n8109 , 2_n8110 , 2_n8111 , 2_n8112 , 2_n8113 , 2_n8114 , 2_n8115 , 2_n8116 , 2_n8117 , 2_n8118 , 2_n8119 , 2_n8120 , 2_n8121 , 2_n8122 , 2_n8123 , 2_n8124 , 2_n8125 , 2_n8126 , 2_n8127 , 2_n8128 , 2_n8129 , 2_n8130 , 2_n8131 , 2_n8132 , 2_n8133 , 2_n8134 , 2_n8135 , 2_n8136 , 2_n8137 , 2_n8139 , 2_n8140 , 2_n8141 , 2_n8142 , 2_n8143 , 2_n8144 , 2_n8145 , 2_n8146 , 2_n8147 , 2_n8148 , 2_n8149 , 2_n8150 , 2_n8151 , 2_n8152 , 2_n8153 , 2_n8154 , 2_n8155 , 2_n8156 , 2_n8157 , 2_n8158 , 2_n8159 , 2_n8160 , 2_n8161 , 2_n8162 , 2_n8163 , 2_n8164 , 2_n8165 , 2_n8166 , 2_n8167 , 2_n8168 , 2_n8169 , 2_n8170 , 2_n8171 , 2_n8172 , 2_n8173 , 2_n8174 , 2_n8175 , 2_n8176 , 2_n8177 , 2_n8178 , 2_n8179 , 2_n8180 , 2_n8181 , 2_n8182 , 2_n8183 , 2_n8184 , 2_n8185 , 2_n8186 , 2_n8187 , 2_n8188 , 2_n8189 , 2_n8190 , 2_n8191 , 2_n8192 , 2_n8193 , 2_n8194 , 2_n8195 , 2_n8196 , 2_n8197 , 2_n8198 , 2_n8199 , 2_n8200 , 2_n8201 , 2_n8203 , 2_n8204 , 2_n8205 , 2_n8206 , 2_n8207 , 2_n8208 , 2_n8209 , 2_n8210 , 2_n8211 , 2_n8212 , 2_n8213 , 2_n8214 , 2_n8215 , 2_n8216 , 2_n8217 , 2_n8218 , 2_n8219 , 2_n8220 , 2_n8221 , 2_n8222 , 2_n8223 , 2_n8224 , 2_n8225 , 2_n8226 , 2_n8227 , 2_n8228 , 2_n8229 , 2_n8230 , 2_n8231 , 2_n8232 , 2_n8233 , 2_n8234 , 2_n8235 , 2_n8237 , 2_n8238 , 2_n8239 , 2_n8240 , 2_n8241 , 2_n8242 , 2_n8243 , 2_n8244 , 2_n8245 , 2_n8246 , 2_n8247 , 2_n8248 , 2_n8249 , 2_n8250 , 2_n8251 , 2_n8252 , 2_n8253 , 2_n8254 , 2_n8255 , 2_n8256 , 2_n8257 , 2_n8258 , 2_n8259 , 2_n8260 , 2_n8261 , 2_n8262 , 2_n8263 , 2_n8264 , 2_n8265 , 2_n8266 , 2_n8267 , 2_n8268 , 2_n8269 , 2_n8270 , 2_n8271 , 2_n8272 , 2_n8273 , 2_n8274 , 2_n8275 , 2_n8277 , 2_n8278 , 2_n8279 , 2_n8280 , 2_n8281 , 2_n8282 , 2_n8283 , 2_n8284 , 2_n8285 , 2_n8286 , 2_n8287 , 2_n8288 , 2_n8289 , 2_n8290 , 2_n8291 , 2_n8292 , 2_n8293 , 2_n8294 , 2_n8295 , 2_n8296 , 2_n8297 , 2_n8298 , 2_n8299 , 2_n8300 , 2_n8301 , 2_n8302 , 2_n8304 , 2_n8305 , 2_n8306 , 2_n8307 , 2_n8308 , 2_n8309 , 2_n8310 , 2_n8311 , 2_n8312 , 2_n8313 , 2_n8314 , 2_n8315 , 2_n8316 , 2_n8317 , 2_n8318 , 2_n8319 , 2_n8320 , 2_n8321 , 2_n8322 , 2_n8323 , 2_n8324 , 2_n8325 , 2_n8326 , 2_n8327 , 2_n8328 , 2_n8329 , 2_n8330 , 2_n8331 , 2_n8332 , 2_n8333 , 2_n8334 , 2_n8335 , 2_n8337 , 2_n8338 , 2_n8339 , 2_n8340 , 2_n8341 , 2_n8342 , 2_n8343 , 2_n8344 , 2_n8345 , 2_n8346 , 2_n8347 , 2_n8348 , 2_n8349 , 2_n8350 , 2_n8351 , 2_n8352 , 2_n8353 , 2_n8354 , 2_n8355 , 2_n8356 , 2_n8357 , 2_n8358 , 2_n8359 , 2_n8360 , 2_n8361 , 2_n8362 , 2_n8363 , 2_n8364 , 2_n8365 , 2_n8366 , 2_n8367 , 2_n8368 , 2_n8369 , 2_n8370 , 2_n8371 , 2_n8372 , 2_n8373 , 2_n8374 , 2_n8375 , 2_n8376 , 2_n8377 , 2_n8378 , 2_n8379 , 2_n8380 , 2_n8381 , 2_n8382 , 2_n8383 , 2_n8385 , 2_n8386 , 2_n8387 , 2_n8388 , 2_n8389 , 2_n8390 , 2_n8391 , 2_n8392 , 2_n8393 , 2_n8394 , 2_n8395 , 2_n8396 , 2_n8397 , 2_n8399 , 2_n8400 , 2_n8401 , 2_n8402 , 2_n8403 , 2_n8404 , 2_n8405 , 2_n8406 , 2_n8407 , 2_n8408 , 2_n8409 , 2_n8410 , 2_n8411 , 2_n8412 , 2_n8413 , 2_n8414 , 2_n8415 , 2_n8416 , 2_n8417 , 2_n8418 , 2_n8419 , 2_n8420 , 2_n8421 , 2_n8422 , 2_n8423 , 2_n8424 , 2_n8425 , 2_n8426 , 2_n8427 , 2_n8428 , 2_n8429 , 2_n8430 , 2_n8431 , 2_n8432 , 2_n8434 , 2_n8435 , 2_n8436 , 2_n8437 , 2_n8438 , 2_n8439 , 2_n8440 , 2_n8441 , 2_n8442 , 2_n8443 , 2_n8444 , 2_n8445 , 2_n8446 , 2_n8447 , 2_n8448 , 2_n8449 , 2_n8450 , 2_n8451 , 2_n8452 , 2_n8453 , 2_n8454 , 2_n8455 , 2_n8456 , 2_n8457 , 2_n8458 , 2_n8459 , 2_n8460 , 2_n8461 , 2_n8462 , 2_n8463 , 2_n8464 , 2_n8465 , 2_n8466 , 2_n8467 , 2_n8468 , 2_n8469 , 2_n8470 , 2_n8471 , 2_n8472 , 2_n8473 , 2_n8474 , 2_n8475 , 2_n8477 , 2_n8478 , 2_n8479 , 2_n8480 , 2_n8481 , 2_n8482 , 2_n8483 , 2_n8484 , 2_n8485 , 2_n8486 , 2_n8487 , 2_n8488 , 2_n8489 , 2_n8490 , 2_n8491 , 2_n8492 , 2_n8493 , 2_n8494 , 2_n8495 , 2_n8496 , 2_n8497 , 2_n8498 , 2_n8499 , 2_n8500 , 2_n8501 , 2_n8502 , 2_n8503 , 2_n8504 , 2_n8505 , 2_n8506 , 2_n8507 , 2_n8508 , 2_n8509 , 2_n8510 , 2_n8511 , 2_n8512 , 2_n8513 , 2_n8514 , 2_n8515 , 2_n8516 , 2_n8517 , 2_n8518 , 2_n8519 , 2_n8520 , 2_n8521 , 2_n8522 , 2_n8523 , 2_n8524 , 2_n8525 , 2_n8526 , 2_n8527 , 2_n8528 , 2_n8529 , 2_n8530 , 2_n8531 , 2_n8532 , 2_n8533 , 2_n8534 , 2_n8535 , 2_n8536 , 2_n8537 , 2_n8538 , 2_n8539 , 2_n8540 , 2_n8541 , 2_n8542 , 2_n8543 , 2_n8544 , 2_n8545 , 2_n8546 , 2_n8547 , 2_n8548 , 2_n8549 , 2_n8550 , 2_n8551 , 2_n8552 , 2_n8553 , 2_n8554 , 2_n8555 , 2_n8556 , 2_n8557 , 2_n8558 , 2_n8559 , 2_n8560 , 2_n8561 , 2_n8562 , 2_n8563 , 2_n8564 , 2_n8565 , 2_n8566 , 2_n8567 , 2_n8568 , 2_n8569 , 2_n8570 , 2_n8571 , 2_n8572 , 2_n8573 , 2_n8574 , 2_n8575 , 2_n8576 , 2_n8577 , 2_n8578 , 2_n8579 , 2_n8580 , 2_n8581 , 2_n8582 , 2_n8583 , 2_n8584 , 2_n8585 , 2_n8586 , 2_n8587 , 2_n8588 , 2_n8589 , 2_n8590 , 2_n8591 , 2_n8592 , 2_n8593 , 2_n8594 , 2_n8596 , 2_n8597 , 2_n8598 , 2_n8599 , 2_n8600 , 2_n8601 , 2_n8602 , 2_n8603 , 2_n8604 , 2_n8605 , 2_n8606 , 2_n8607 , 2_n8608 , 2_n8609 , 2_n8610 , 2_n8611 , 2_n8612 , 2_n8613 , 2_n8614 , 2_n8615 , 2_n8616 , 2_n8617 , 2_n8618 , 2_n8619 , 2_n8620 , 2_n8621 , 2_n8622 , 2_n8623 , 2_n8624 , 2_n8625 , 2_n8626 , 2_n8627 , 2_n8628 , 2_n8629 , 2_n8630 , 2_n8631 , 2_n8632 , 2_n8633 , 2_n8634 , 2_n8635 , 2_n8636 , 2_n8637 , 2_n8638 , 2_n8639 , 2_n8640 , 2_n8641 , 2_n8642 , 2_n8643 , 2_n8644 , 2_n8645 , 2_n8646 , 2_n8647 , 2_n8648 , 2_n8649 , 2_n8650 , 2_n8651 , 2_n8652 , 2_n8653 , 2_n8654 , 2_n8655 , 2_n8656 , 2_n8657 , 2_n8658 , 2_n8659 , 2_n8660 , 2_n8661 , 2_n8662 , 2_n8663 , 2_n8664 , 2_n8666 , 2_n8667 , 2_n8668 , 2_n8669 , 2_n8670 , 2_n8671 , 2_n8672 , 2_n8673 , 2_n8674 , 2_n8675 , 2_n8676 , 2_n8677 , 2_n8678 , 2_n8679 , 2_n8680 , 2_n8681 , 2_n8682 , 2_n8683 , 2_n8684 , 2_n8685 , 2_n8686 , 2_n8687 , 2_n8688 , 2_n8689 , 2_n8690 , 2_n8691 , 2_n8692 , 2_n8693 , 2_n8694 , 2_n8695 , 2_n8696 , 2_n8697 , 2_n8698 , 2_n8699 , 2_n8700 , 2_n8701 , 2_n8702 , 2_n8703 , 2_n8704 , 2_n8705 , 2_n8706 , 2_n8707 , 2_n8708 , 2_n8709 , 2_n8710 , 2_n8711 , 2_n8712 , 2_n8713 , 2_n8714 , 2_n8715 , 2_n8716 , 2_n8718 , 2_n8719 , 2_n8720 , 2_n8721 , 2_n8722 , 2_n8723 , 2_n8724 , 2_n8725 , 2_n8726 , 2_n8727 , 2_n8728 , 2_n8729 , 2_n8730 , 2_n8731 , 2_n8732 , 2_n8733 , 2_n8734 , 2_n8735 , 2_n8736 , 2_n8737 , 2_n8738 , 2_n8739 , 2_n8740 , 2_n8741 , 2_n8742 , 2_n8743 , 2_n8744 , 2_n8745 , 2_n8746 , 2_n8747 , 2_n8748 , 2_n8749 , 2_n8750 , 2_n8751 , 2_n8752 , 2_n8753 , 2_n8754 , 2_n8755 , 2_n8756 , 2_n8757 , 2_n8758 , 2_n8760 , 2_n8761 , 2_n8762 , 2_n8763 , 2_n8764 , 2_n8765 , 2_n8766 , 2_n8767 , 2_n8768 , 2_n8769 , 2_n8770 , 2_n8771 , 2_n8772 , 2_n8773 , 2_n8774 , 2_n8775 , 2_n8776 , 2_n8777 , 2_n8778 , 2_n8779 , 2_n8780 , 2_n8781 , 2_n8782 , 2_n8783 , 2_n8784 , 2_n8785 , 2_n8786 , 2_n8787 , 2_n8788 , 2_n8789 , 2_n8790 , 2_n8791 , 2_n8792 , 2_n8793 , 2_n8794 , 2_n8795 , 2_n8796 , 2_n8797 , 2_n8798 , 2_n8799 , 2_n8800 , 2_n8801 , 2_n8802 , 2_n8803 , 2_n8804 , 2_n8805 , 2_n8806 , 2_n8807 , 2_n8808 , 2_n8809 , 2_n8810 , 2_n8811 , 2_n8812 , 2_n8813 , 2_n8814 , 2_n8815 , 2_n8816 , 2_n8817 , 2_n8818 , 2_n8820 , 2_n8821 , 2_n8822 , 2_n8823 , 2_n8824 , 2_n8825 , 2_n8826 , 2_n8827 , 2_n8828 , 2_n8829 , 2_n8830 , 2_n8831 , 2_n8832 , 2_n8833 , 2_n8834 , 2_n8835 , 2_n8836 , 2_n8837 , 2_n8838 , 2_n8839 , 2_n8840 , 2_n8841 , 2_n8842 , 2_n8843 , 2_n8844 , 2_n8845 , 2_n8846 , 2_n8847 , 2_n8848 , 2_n8849 , 2_n8850 , 2_n8851 , 2_n8852 , 2_n8853 , 2_n8854 , 2_n8855 , 2_n8856 , 2_n8857 , 2_n8858 , 2_n8859 , 2_n8860 , 2_n8861 , 2_n8862 , 2_n8863 , 2_n8864 , 2_n8865 , 2_n8866 , 2_n8867 , 2_n8868 , 2_n8869 , 2_n8870 , 2_n8871 , 2_n8872 , 2_n8873 , 2_n8874 , 2_n8875 , 2_n8876 , 2_n8877 , 2_n8878 , 2_n8879 , 2_n8880 , 2_n8881 , 2_n8882 , 2_n8883 , 2_n8884 , 2_n8885 , 2_n8886 , 2_n8887 , 2_n8888 , 2_n8889 , 2_n8890 , 2_n8891 , 2_n8892 , 2_n8893 , 2_n8894 , 2_n8895 , 2_n8896 , 2_n8897 , 2_n8898 , 2_n8899 , 2_n8900 , 2_n8901 , 2_n8902 , 2_n8903 , 2_n8904 , 2_n8905 , 2_n8906 , 2_n8907 , 2_n8908 , 2_n8909 , 2_n8910 , 2_n8911 , 2_n8912 , 2_n8913 , 2_n8914 , 2_n8915 , 2_n8916 , 2_n8917 , 2_n8918 , 2_n8919 , 2_n8920 , 2_n8921 , 2_n8922 , 2_n8923 , 2_n8924 , 2_n8925 , 2_n8926 , 2_n8927 , 2_n8928 , 2_n8929 , 2_n8930 , 2_n8931 , 2_n8932 , 2_n8933 , 2_n8934 , 2_n8935 , 2_n8936 , 2_n8937 , 2_n8938 , 2_n8939 , 2_n8940 , 2_n8941 , 2_n8942 , 2_n8943 , 2_n8944 , 2_n8945 , 2_n8946 , 2_n8947 , 2_n8948 , 2_n8949 , 2_n8950 , 2_n8951 , 2_n8952 , 2_n8953 , 2_n8954 , 2_n8955 , 2_n8956 , 2_n8957 , 2_n8958 , 2_n8959 , 2_n8960 , 2_n8961 , 2_n8962 , 2_n8963 , 2_n8964 , 2_n8965 , 2_n8966 , 2_n8967 , 2_n8968 , 2_n8969 , 2_n8970 , 2_n8971 , 2_n8972 , 2_n8973 , 2_n8974 , 2_n8975 , 2_n8976 , 2_n8977 , 2_n8978 , 2_n8979 , 2_n8980 , 2_n8981 , 2_n8982 , 2_n8983 , 2_n8984 , 2_n8985 , 2_n8986 , 2_n8987 , 2_n8988 , 2_n8989 , 2_n8990 , 2_n8991 , 2_n8992 , 2_n8993 , 2_n8994 , 2_n8995 , 2_n8996 , 2_n8997 , 2_n8998 , 2_n8999 , 2_n9000 , 2_n9001 , 2_n9002 , 2_n9003 , 2_n9004 , 2_n9005 , 2_n9006 , 2_n9007 , 2_n9008 , 2_n9009 , 2_n9010 , 2_n9011 , 2_n9012 , 2_n9013 , 2_n9014 , 2_n9015 , 2_n9016 , 2_n9017 , 2_n9018 , 2_n9019 , 2_n9020 , 2_n9021 , 2_n9022 , 2_n9023 , 2_n9024 , 2_n9025 , 2_n9026 , 2_n9027 , 2_n9028 , 2_n9029 , 2_n9030 , 2_n9031 , 2_n9032 , 2_n9033 , 2_n9034 , 2_n9035 , 2_n9036 , 2_n9037 , 2_n9038 , 2_n9039 , 2_n9040 , 2_n9041 , 2_n9042 , 2_n9043 , 2_n9044 , 2_n9045 , 2_n9046 , 2_n9047 , 2_n9048 , 2_n9049 , 2_n9050 , 2_n9051 , 2_n9052 , 2_n9053 , 2_n9054 , 2_n9055 , 2_n9056 , 2_n9057 , 2_n9058 , 2_n9059 , 2_n9060 , 2_n9061 , 2_n9062 , 2_n9063 , 2_n9064 , 2_n9065 , 2_n9066 , 2_n9067 , 2_n9068 , 2_n9069 , 2_n9070 , 2_n9071 , 2_n9072 , 2_n9073 , 2_n9074 , 2_n9075 , 2_n9076 , 2_n9077 , 2_n9078 , 2_n9079 , 2_n9081 , 2_n9082 , 2_n9083 , 2_n9084 , 2_n9085 , 2_n9086 , 2_n9087 , 2_n9088 , 2_n9089 , 2_n9090 , 2_n9091 , 2_n9092 , 2_n9093 , 2_n9094 , 2_n9095 , 2_n9096 , 2_n9097 , 2_n9098 , 2_n9099 , 2_n9100 , 2_n9101 , 2_n9102 , 2_n9103 , 2_n9104 , 2_n9105 , 2_n9106 , 2_n9107 , 2_n9108 , 2_n9109 , 2_n9110 , 2_n9112 , 2_n9113 , 2_n9114 , 2_n9115 , 2_n9116 , 2_n9117 , 2_n9118 , 2_n9119 , 2_n9120 , 2_n9121 , 2_n9122 , 2_n9123 , 2_n9124 , 2_n9125 , 2_n9126 , 2_n9127 , 2_n9128 , 2_n9129 , 2_n9130 , 2_n9131 , 2_n9132 , 2_n9133 , 2_n9134 , 2_n9135 , 2_n9136 , 2_n9138 , 2_n9139 , 2_n9140 , 2_n9141 , 2_n9142 , 2_n9143 , 2_n9144 , 2_n9145 , 2_n9146 , 2_n9147 , 2_n9148 , 2_n9149 , 2_n9150 , 2_n9151 , 2_n9152 , 2_n9153 , 2_n9154 , 2_n9155 , 2_n9156 , 2_n9157 , 2_n9158 , 2_n9159 , 2_n9160 , 2_n9161 , 2_n9162 , 2_n9163 , 2_n9164 , 2_n9165 , 2_n9166 , 2_n9167 , 2_n9168 , 2_n9169 , 2_n9170 , 2_n9171 , 2_n9172 , 2_n9173 , 2_n9174 , 2_n9175 , 2_n9176 , 2_n9177 , 2_n9178 , 2_n9179 , 2_n9180 , 2_n9181 , 2_n9182 , 2_n9183 , 2_n9184 , 2_n9185 , 2_n9186 , 2_n9187 , 2_n9188 , 2_n9190 , 2_n9191 , 2_n9192 , 2_n9193 , 2_n9194 , 2_n9196 , 2_n9197 , 2_n9198 , 2_n9199 , 2_n9200 , 2_n9201 , 2_n9202 , 2_n9203 , 2_n9204 , 2_n9205 , 2_n9206 , 2_n9207 , 2_n9208 , 2_n9209 , 2_n9210 , 2_n9211 , 2_n9212 , 2_n9213 , 2_n9214 , 2_n9215 , 2_n9216 , 2_n9217 , 2_n9218 , 2_n9219 , 2_n9220 , 2_n9221 , 2_n9222 , 2_n9223 , 2_n9224 , 2_n9225 , 2_n9226 , 2_n9227 , 2_n9228 , 2_n9229 , 2_n9230 , 2_n9231 , 2_n9232 , 2_n9233 , 2_n9234 , 2_n9235 , 2_n9236 , 2_n9237 , 2_n9238 , 2_n9239 , 2_n9240 , 2_n9242 , 2_n9243 , 2_n9244 , 2_n9245 , 2_n9246 , 2_n9247 , 2_n9248 , 2_n9249 , 2_n9250 , 2_n9251 , 2_n9252 , 2_n9253 , 2_n9254 , 2_n9255 , 2_n9256 , 2_n9257 , 2_n9258 , 2_n9259 , 2_n9260 , 2_n9261 , 2_n9262 , 2_n9263 , 2_n9264 , 2_n9265 , 2_n9266 , 2_n9267 , 2_n9268 , 2_n9269 , 2_n9270 , 2_n9271 , 2_n9272 , 2_n9273 , 2_n9274 , 2_n9275 , 2_n9276 , 2_n9277 , 2_n9278 , 2_n9279 , 2_n9280 , 2_n9281 , 2_n9282 , 2_n9283 , 2_n9284 , 2_n9285 , 2_n9286 , 2_n9287 , 2_n9288 , 2_n9289 , 2_n9290 , 2_n9291 , 2_n9292 , 2_n9293 , 2_n9294 , 2_n9295 , 2_n9296 , 2_n9297 , 2_n9298 , 2_n9299 , 2_n9300 , 2_n9301 , 2_n9302 , 2_n9303 , 2_n9304 , 2_n9305 , 2_n9306 , 2_n9307 , 2_n9308 , 2_n9309 , 2_n9310 , 2_n9311 , 2_n9312 , 2_n9313 , 2_n9314 , 2_n9315 , 2_n9316 , 2_n9317 , 2_n9318 , 2_n9319 , 2_n9320 , 2_n9321 , 2_n9322 , 2_n9323 , 2_n9324 , 2_n9325 , 2_n9326 , 2_n9327 , 2_n9328 , 2_n9329 , 2_n9330 , 2_n9331 , 2_n9332 , 2_n9333 , 2_n9334 , 2_n9335 , 2_n9336 , 2_n9337 , 2_n9338 , 2_n9339 , 2_n9340 , 2_n9341 , 2_n9342 , 2_n9343 , 2_n9344 , 2_n9345 , 2_n9346 , 2_n9347 , 2_n9348 , 2_n9349 , 2_n9350 , 2_n9351 , 2_n9352 , 2_n9353 , 2_n9354 , 2_n9355 , 2_n9356 , 2_n9357 , 2_n9358 , 2_n9359 , 2_n9360 , 2_n9361 , 2_n9362 , 2_n9363 , 2_n9364 , 2_n9365 , 2_n9366 , 2_n9367 , 2_n9368 , 2_n9369 , 2_n9370 , 2_n9371 , 2_n9372 , 2_n9373 , 2_n9374 , 2_n9375 , 2_n9376 , 2_n9377 , 2_n9378 , 2_n9379 , 2_n9380 , 2_n9381 , 2_n9382 , 2_n9383 , 2_n9384 , 2_n9385 , 2_n9386 , 2_n9388 , 2_n9389 , 2_n9390 , 2_n9391 , 2_n9392 , 2_n9393 , 2_n9394 , 2_n9395 , 2_n9396 , 2_n9397 , 2_n9398 , 2_n9399 , 2_n9401 , 2_n9402 , 2_n9403 , 2_n9404 , 2_n9405 , 2_n9406 , 2_n9407 , 2_n9408 , 2_n9409 , 2_n9410 , 2_n9411 , 2_n9412 , 2_n9413 , 2_n9414 , 2_n9415 , 2_n9416 , 2_n9417 , 2_n9418 , 2_n9419 , 2_n9420 , 2_n9421 , 2_n9422 , 2_n9423 , 2_n9424 , 2_n9425 , 2_n9426 , 2_n9427 , 2_n9428 , 2_n9429 , 2_n9430 , 2_n9431 , 2_n9432 , 2_n9433 , 2_n9434 , 2_n9435 , 2_n9436 , 2_n9437 , 2_n9438 , 2_n9439 , 2_n9440 , 2_n9441 , 2_n9442 , 2_n9443 , 2_n9444 , 2_n9445 , 2_n9446 , 2_n9447 , 2_n9448 , 2_n9449 , 2_n9450 , 2_n9451 , 2_n9452 , 2_n9453 , 2_n9454 , 2_n9455 , 2_n9456 , 2_n9458 , 2_n9459 , 2_n9460 , 2_n9461 , 2_n9462 , 2_n9463 , 2_n9464 , 2_n9465 , 2_n9466 , 2_n9467 , 2_n9468 , 2_n9469 , 2_n9470 , 2_n9471 , 2_n9472 , 2_n9473 , 2_n9474 , 2_n9475 , 2_n9476 , 2_n9477 , 2_n9478 , 2_n9479 , 2_n9480 , 2_n9481 , 2_n9482 , 2_n9483 , 2_n9484 , 2_n9485 , 2_n9486 , 2_n9487 , 2_n9488 , 2_n9489 , 2_n9490 , 2_n9491 , 2_n9492 , 2_n9493 , 2_n9494 , 2_n9495 , 2_n9496 , 2_n9497 , 2_n9498 , 2_n9499 , 2_n9500 , 2_n9501 , 2_n9502 , 2_n9503 , 2_n9504 , 2_n9505 , 2_n9506 , 2_n9507 , 2_n9508 , 2_n9509 , 2_n9510 , 2_n9511 , 2_n9512 , 2_n9513 , 2_n9514 , 2_n9515 , 2_n9516 , 2_n9517 , 2_n9518 , 2_n9519 , 2_n9520 , 2_n9521 , 2_n9522 , 2_n9523 , 2_n9524 , 2_n9525 , 2_n9526 , 2_n9527 , 2_n9528 , 2_n9529 , 2_n9530 , 2_n9531 , 2_n9532 , 2_n9533 , 2_n9534 , 2_n9535 , 2_n9536 , 2_n9537 , 2_n9538 , 2_n9539 , 2_n9540 , 2_n9541 , 2_n9542 , 2_n9543 , 2_n9544 , 2_n9545 , 2_n9546 , 2_n9547 , 2_n9548 , 2_n9549 , 2_n9550 , 2_n9551 , 2_n9552 , 2_n9553 , 2_n9554 , 2_n9555 , 2_n9556 , 2_n9557 , 2_n9558 , 2_n9559 , 2_n9560 , 2_n9561 , 2_n9562 , 2_n9563 , 2_n9564 , 2_n9565 , 2_n9566 , 2_n9567 , 2_n9568 , 2_n9569 , 2_n9570 , 2_n9572 , 2_n9573 , 2_n9574 , 2_n9575 , 2_n9576 , 2_n9577 , 2_n9579 , 2_n9580 , 2_n9581 , 2_n9582 , 2_n9584 , 2_n9585 , 2_n9586 , 2_n9587 , 2_n9588 , 2_n9589 , 2_n9590 , 2_n9591 , 2_n9592 , 2_n9593 , 2_n9594 , 2_n9595 , 2_n9596 , 2_n9597 , 2_n9598 , 2_n9599 , 2_n9600 , 2_n9601 , 2_n9602 , 2_n9603 , 2_n9604 , 2_n9605 , 2_n9606 , 2_n9607 , 2_n9608 , 2_n9609 , 2_n9610 , 2_n9611 , 2_n9612 , 2_n9613 , 2_n9614 , 2_n9615 , 2_n9616 , 2_n9617 , 2_n9618 , 2_n9619 , 2_n9620 , 2_n9621 , 2_n9622 , 2_n9623 , 2_n9624 , 2_n9625 , 2_n9626 , 2_n9627 , 2_n9628 , 2_n9629 , 2_n9630 , 2_n9631 , 2_n9632 , 2_n9633 , 2_n9634 , 2_n9635 , 2_n9636 , 2_n9638 , 2_n9639 , 2_n9641 , 2_n9642 , 2_n9643 , 2_n9644 , 2_n9645 , 2_n9646 , 2_n9647 , 2_n9648 , 2_n9649 , 2_n9650 , 2_n9651 , 2_n9652 , 2_n9653 , 2_n9654 , 2_n9655 , 2_n9656 , 2_n9657 , 2_n9658 , 2_n9659 , 2_n9660 , 2_n9661 , 2_n9662 , 2_n9663 , 2_n9664 , 2_n9665 , 2_n9666 , 2_n9667 , 2_n9668 , 2_n9669 , 2_n9670 , 2_n9671 , 2_n9672 , 2_n9673 , 2_n9674 , 2_n9675 , 2_n9676 , 2_n9677 , 2_n9678 , 2_n9679 , 2_n9680 , 2_n9681 , 2_n9682 , 2_n9683 , 2_n9684 , 2_n9685 , 2_n9686 , 2_n9687 , 2_n9688 , 2_n9689 , 2_n9690 , 2_n9691 , 2_n9692 , 2_n9693 , 2_n9694 , 2_n9695 , 2_n9696 , 2_n9697 , 2_n9698 , 2_n9699 , 2_n9700 , 2_n9701 , 2_n9702 , 2_n9703 , 2_n9704 , 2_n9705 , 2_n9707 , 2_n9708 , 2_n9709 , 2_n9710 , 2_n9711 , 2_n9712 , 2_n9713 , 2_n9714 , 2_n9715 , 2_n9716 , 2_n9717 , 2_n9718 , 2_n9719 , 2_n9720 , 2_n9721 , 2_n9722 , 2_n9723 , 2_n9724 , 2_n9726 , 2_n9727 , 2_n9728 , 2_n9729 , 2_n9730 , 2_n9731 , 2_n9732 , 2_n9733 , 2_n9734 , 2_n9735 , 2_n9736 , 2_n9737 , 2_n9738 , 2_n9739 , 2_n9740 , 2_n9741 , 2_n9742 , 2_n9743 , 2_n9744 , 2_n9745 , 2_n9746 , 2_n9747 , 2_n9748 , 2_n9749 , 2_n9750 , 2_n9751 , 2_n9752 , 2_n9753 , 2_n9754 , 2_n9755 , 2_n9757 , 2_n9758 , 2_n9759 , 2_n9760 , 2_n9761 , 2_n9762 , 2_n9764 , 2_n9765 , 2_n9766 , 2_n9768 , 2_n9769 , 2_n9770 , 2_n9771 , 2_n9772 , 2_n9773 , 2_n9774 , 2_n9775 , 2_n9776 , 2_n9777 , 2_n9778 , 2_n9779 , 2_n9780 , 2_n9781 , 2_n9782 , 2_n9783 , 2_n9784 , 2_n9785 , 2_n9786 , 2_n9787 , 2_n9788 , 2_n9789 , 2_n9790 , 2_n9791 , 2_n9792 , 2_n9793 , 2_n9794 , 2_n9795 , 2_n9796 , 2_n9797 , 2_n9798 , 2_n9799 , 2_n9800 , 2_n9801 , 2_n9802 , 2_n9803 , 2_n9804 , 2_n9805 , 2_n9806 , 2_n9807 , 2_n9808 , 2_n9809 , 2_n9810 , 2_n9811 , 2_n9812 , 2_n9813 , 2_n9814 , 2_n9815 , 2_n9816 , 2_n9817 , 2_n9818 , 2_n9819 , 2_n9821 , 2_n9822 , 2_n9823 , 2_n9824 , 2_n9825 , 2_n9826 , 2_n9827 , 2_n9828 , 2_n9829 , 2_n9830 , 2_n9831 , 2_n9832 , 2_n9833 , 2_n9834 , 2_n9835 , 2_n9836 , 2_n9837 , 2_n9838 , 2_n9839 , 2_n9840 , 2_n9841 , 2_n9842 , 2_n9843 , 2_n9844 , 2_n9845 , 2_n9846 , 2_n9847 , 2_n9848 , 2_n9849 , 2_n9850 , 2_n9851 , 2_n9852 , 2_n9853 , 2_n9854 , 2_n9855 , 2_n9856 , 2_n9857 , 2_n9858 , 2_n9859 , 2_n9860 , 2_n9861 , 2_n9862 , 2_n9863 , 2_n9864 , 2_n9865 , 2_n9866 , 2_n9867 , 2_n9868 , 2_n9869 , 2_n9870 , 2_n9871 , 2_n9872 , 2_n9873 , 2_n9874 , 2_n9875 , 2_n9876 , 2_n9877 , 2_n9878 , 2_n9879 , 2_n9880 , 2_n9881 , 2_n9882 , 2_n9883 , 2_n9884 , 2_n9885 , 2_n9886 , 2_n9887 , 2_n9888 , 2_n9889 , 2_n9890 , 2_n9891 , 2_n9892 , 2_n9893 , 2_n9894 , 2_n9895 , 2_n9896 , 2_n9897 , 2_n9898 , 2_n9899 , 2_n9900 , 2_n9901 , 2_n9902 , 2_n9903 , 2_n9904 , 2_n9905 , 2_n9906 , 2_n9907 , 2_n9908 , 2_n9909 , 2_n9910 , 2_n9911 , 2_n9912 , 2_n9913 , 2_n9914 , 2_n9915 , 2_n9916 , 2_n9917 , 2_n9918 , 2_n9919 , 2_n9921 , 2_n9922 , 2_n9923 , 2_n9924 , 2_n9925 , 2_n9926 , 2_n9927 , 2_n9928 , 2_n9929 , 2_n9930 , 2_n9931 , 2_n9932 , 2_n9933 , 2_n9934 , 2_n9935 , 2_n9936 , 2_n9937 , 2_n9939 , 2_n9940 , 2_n9941 , 2_n9942 , 2_n9943 , 2_n9944 , 2_n9945 , 2_n9946 , 2_n9947 , 2_n9948 , 2_n9949 , 2_n9950 , 2_n9951 , 2_n9952 , 2_n9953 , 2_n9954 , 2_n9955 , 2_n9957 , 2_n9958 , 2_n9959 , 2_n9960 , 2_n9961 , 2_n9962 , 2_n9963 , 2_n9964 , 2_n9965 , 2_n9966 , 2_n9967 , 2_n9968 , 2_n9969 , 2_n9970 , 2_n9971 , 2_n9972 , 2_n9973 , 2_n9974 , 2_n9975 , 2_n9976 , 2_n9977 , 2_n9978 , 2_n9979 , 2_n9980 , 2_n9981 , 2_n9982 , 2_n9983 , 2_n9984 , 2_n9985 , 2_n9986 , 2_n9987 , 2_n9988 , 2_n9989 , 2_n9990 , 2_n9991 , 2_n9992 , 2_n9993 , 2_n9994 , 2_n9995 , 2_n9996 , 2_n9997 , 2_n9998 , 2_n9999 , 2_n10000 , 2_n10001 , 2_n10002 , 2_n10003 , 2_n10004 , 2_n10005 , 2_n10006 , 2_n10007 , 2_n10008 , 2_n10009 , 2_n10010 , 2_n10011 , 2_n10012 , 2_n10013 , 2_n10014 , 2_n10015 , 2_n10016 , 2_n10017 , 2_n10018 , 2_n10019 , 2_n10020 , 2_n10021 , 2_n10023 , 2_n10024 , 2_n10025 , 2_n10026 , 2_n10027 , 2_n10028 , 2_n10029 , 2_n10030 , 2_n10031 , 2_n10032 , 2_n10033 , 2_n10034 , 2_n10035 , 2_n10036 , 2_n10037 , 2_n10038 , 2_n10039 , 2_n10040 , 2_n10041 , 2_n10042 , 2_n10043 , 2_n10044 , 2_n10045 , 2_n10046 , 2_n10047 , 2_n10048 , 2_n10049 , 2_n10050 , 2_n10051 , 2_n10052 , 2_n10053 , 2_n10054 , 2_n10055 , 2_n10056 , 2_n10057 , 2_n10058 , 2_n10059 , 2_n10060 , 2_n10061 , 2_n10062 , 2_n10063 , 2_n10064 , 2_n10065 , 2_n10066 , 2_n10067 , 2_n10068 , 2_n10069 , 2_n10070 , 2_n10071 , 2_n10072 , 2_n10073 , 2_n10074 , 2_n10075 , 2_n10076 , 2_n10077 , 2_n10078 , 2_n10079 , 2_n10080 , 2_n10081 , 2_n10082 , 2_n10083 , 2_n10084 , 2_n10085 , 2_n10086 , 2_n10087 , 2_n10088 , 2_n10089 , 2_n10090 , 2_n10091 , 2_n10092 , 2_n10093 , 2_n10094 , 2_n10095 , 2_n10096 , 2_n10097 , 2_n10098 , 2_n10099 , 2_n10100 , 2_n10101 , 2_n10102 , 2_n10103 , 2_n10104 , 2_n10105 , 2_n10106 , 2_n10107 , 2_n10108 , 2_n10109 , 2_n10110 , 2_n10111 , 2_n10112 , 2_n10113 , 2_n10114 , 2_n10115 , 2_n10116 , 2_n10117 , 2_n10118 , 2_n10119 , 2_n10120 , 2_n10121 , 2_n10122 , 2_n10123 , 2_n10124 , 2_n10125 , 2_n10126 , 2_n10127 , 2_n10128 , 2_n10129 , 2_n10130 , 2_n10131 , 2_n10132 , 2_n10133 , 2_n10134 , 2_n10135 , 2_n10136 , 2_n10137 , 2_n10138 , 2_n10139 , 2_n10140 , 2_n10141 , 2_n10142 , 2_n10143 , 2_n10144 , 2_n10145 , 2_n10146 , 2_n10147 , 2_n10148 , 2_n10149 , 2_n10150 , 2_n10151 , 2_n10152 , 2_n10153 , 2_n10154 , 2_n10155 , 2_n10156 , 2_n10157 , 2_n10158 , 2_n10159 , 2_n10160 , 2_n10161 , 2_n10162 , 2_n10163 , 2_n10164 , 2_n10165 , 2_n10166 , 2_n10167 , 2_n10168 , 2_n10169 , 2_n10170 , 2_n10171 , 2_n10172 , 2_n10173 , 2_n10175 , 2_n10176 , 2_n10177 , 2_n10178 , 2_n10179 , 2_n10180 , 2_n10181 , 2_n10182 , 2_n10183 , 2_n10184 , 2_n10185 , 2_n10186 , 2_n10187 , 2_n10188 , 2_n10189 , 2_n10190 , 2_n10191 , 2_n10192 , 2_n10193 , 2_n10194 , 2_n10195 , 2_n10196 , 2_n10197 , 2_n10198 , 2_n10199 , 2_n10200 , 2_n10201 , 2_n10202 , 2_n10203 , 2_n10204 , 2_n10205 , 2_n10206 , 2_n10207 , 2_n10208 , 2_n10209 , 2_n10210 , 2_n10211 , 2_n10212 , 2_n10213 , 2_n10214 , 2_n10215 , 2_n10216 , 2_n10218 , 2_n10219 , 2_n10220 , 2_n10221 , 2_n10222 , 2_n10224 , 2_n10225 , 2_n10226 , 2_n10227 , 2_n10228 , 2_n10229 , 2_n10230 , 2_n10231 , 2_n10232 , 2_n10233 , 2_n10234 , 2_n10235 , 2_n10236 , 2_n10237 , 2_n10238 , 2_n10239 , 2_n10240 , 2_n10241 , 2_n10242 , 2_n10243 , 2_n10244 , 2_n10245 , 2_n10246 , 2_n10247 , 2_n10248 , 2_n10249 , 2_n10250 , 2_n10251 , 2_n10252 , 2_n10253 , 2_n10254 , 2_n10255 , 2_n10256 , 2_n10257 , 2_n10258 , 2_n10259 , 2_n10260 , 2_n10261 , 2_n10262 , 2_n10263 , 2_n10264 , 2_n10265 , 2_n10266 , 2_n10267 , 2_n10268 , 2_n10269 , 2_n10270 , 2_n10271 , 2_n10272 , 2_n10273 , 2_n10274 , 2_n10275 , 2_n10276 , 2_n10277 , 2_n10279 , 2_n10280 , 2_n10281 , 2_n10282 , 2_n10283 , 2_n10284 , 2_n10285 , 2_n10286 , 2_n10287 , 2_n10288 , 2_n10289 , 2_n10290 , 2_n10291 , 2_n10292 , 2_n10293 , 2_n10294 , 2_n10295 , 2_n10296 , 2_n10297 , 2_n10298 , 2_n10299 , 2_n10300 , 2_n10301 , 2_n10302 , 2_n10303 , 2_n10304 , 2_n10305 , 2_n10306 , 2_n10307 , 2_n10308 , 2_n10309 , 2_n10310 , 2_n10311 , 2_n10312 , 2_n10313 , 2_n10314 , 2_n10315 , 2_n10316 , 2_n10317 , 2_n10318 , 2_n10319 , 2_n10320 , 2_n10321 , 2_n10322 , 2_n10323 , 2_n10324 , 2_n10325 , 2_n10326 , 2_n10328 , 2_n10329 , 2_n10330 , 2_n10331 , 2_n10332 , 2_n10333 , 2_n10334 , 2_n10335 , 2_n10336 , 2_n10337 , 2_n10338 , 2_n10339 , 2_n10340 , 2_n10341 , 2_n10342 , 2_n10343 , 2_n10344 , 2_n10345 , 2_n10346 , 2_n10347 , 2_n10348 , 2_n10349 , 2_n10350 , 2_n10351 , 2_n10352 , 2_n10353 , 2_n10354 , 2_n10355 , 2_n10356 , 2_n10357 , 2_n10358 , 2_n10359 , 2_n10360 , 2_n10361 , 2_n10362 , 2_n10363 , 2_n10364 , 2_n10365 , 2_n10366 , 2_n10367 , 2_n10368 , 2_n10369 , 2_n10370 , 2_n10371 , 2_n10372 , 2_n10373 , 2_n10374 , 2_n10375 , 2_n10376 , 2_n10377 , 2_n10378 , 2_n10379 , 2_n10380 , 2_n10381 , 2_n10382 , 2_n10383 , 2_n10384 , 2_n10385 , 2_n10386 , 2_n10387 , 2_n10388 , 2_n10389 , 2_n10390 , 2_n10392 , 2_n10393 , 2_n10394 , 2_n10395 , 2_n10396 , 2_n10397 , 2_n10398 , 2_n10399 , 2_n10400 , 2_n10401 , 2_n10402 , 2_n10403 , 2_n10404 , 2_n10405 , 2_n10406 , 2_n10407 , 2_n10408 , 2_n10409 , 2_n10410 , 2_n10411 , 2_n10412 , 2_n10413 , 2_n10414 , 2_n10415 , 2_n10416 , 2_n10417 , 2_n10418 , 2_n10419 , 2_n10420 , 2_n10421 , 2_n10422 , 2_n10423 , 2_n10424 , 2_n10425 , 2_n10426 , 2_n10427 , 2_n10428 , 2_n10429 , 2_n10430 , 2_n10431 , 2_n10432 , 2_n10433 , 2_n10434 , 2_n10435 , 2_n10436 , 2_n10437 , 2_n10438 , 2_n10440 , 2_n10441 , 2_n10442 , 2_n10443 , 2_n10444 , 2_n10445 , 2_n10446 , 2_n10447 , 2_n10448 , 2_n10449 , 2_n10450 , 2_n10452 , 2_n10453 , 2_n10454 , 2_n10455 , 2_n10456 , 2_n10457 , 2_n10458 , 2_n10459 , 2_n10460 , 2_n10461 , 2_n10462 , 2_n10463 , 2_n10464 , 2_n10465 , 2_n10466 , 2_n10467 , 2_n10468 , 2_n10469 , 2_n10470 , 2_n10471 , 2_n10472 , 2_n10473 , 2_n10474 , 2_n10475 , 2_n10477 , 2_n10478 , 2_n10479 , 2_n10480 , 2_n10481 , 2_n10482 , 2_n10483 , 2_n10484 , 2_n10485 , 2_n10486 , 2_n10487 , 2_n10488 , 2_n10489 , 2_n10490 , 2_n10491 , 2_n10492 , 2_n10493 , 2_n10494 , 2_n10495 , 2_n10496 , 2_n10497 , 2_n10498 , 2_n10499 , 2_n10500 , 2_n10501 , 2_n10502 , 2_n10503 , 2_n10504 , 2_n10505 , 2_n10506 , 2_n10507 , 2_n10508 , 2_n10509 , 2_n10511 , 2_n10512 , 2_n10513 , 2_n10514 , 2_n10515 , 2_n10516 , 2_n10517 , 2_n10518 , 2_n10519 , 2_n10520 , 2_n10521 , 2_n10522 , 2_n10523 , 2_n10524 , 2_n10525 , 2_n10526 , 2_n10527 , 2_n10528 , 2_n10529 , 2_n10530 , 2_n10531 , 2_n10532 , 2_n10533 , 2_n10534 , 2_n10535 , 2_n10536 , 2_n10537 , 2_n10538 , 2_n10539 , 2_n10540 , 2_n10541 , 2_n10542 , 2_n10543 , 2_n10544 , 2_n10546 , 2_n10548 , 2_n10549 , 2_n10550 , 2_n10551 , 2_n10552 , 2_n10553 , 2_n10554 , 2_n10555 , 2_n10556 , 2_n10557 , 2_n10558 , 2_n10559 , 2_n10560 , 2_n10561 , 2_n10562 , 2_n10563 , 2_n10564 , 2_n10565 , 2_n10566 , 2_n10567 , 2_n10568 , 2_n10569 , 2_n10570 , 2_n10571 , 2_n10572 , 2_n10573 , 2_n10574 , 2_n10575 , 2_n10576 , 2_n10577 , 2_n10578 , 2_n10579 , 2_n10580 , 2_n10581 , 2_n10582 , 2_n10583 , 2_n10584 , 2_n10585 , 2_n10586 , 2_n10587 , 2_n10588 , 2_n10590 , 2_n10591 , 2_n10592 , 2_n10593 , 2_n10594 , 2_n10595 , 2_n10596 , 2_n10597 , 2_n10598 , 2_n10599 , 2_n10600 , 2_n10601 , 2_n10602 , 2_n10603 , 2_n10604 , 2_n10605 , 2_n10606 , 2_n10607 , 2_n10608 , 2_n10609 , 2_n10610 , 2_n10611 , 2_n10612 , 2_n10613 , 2_n10614 , 2_n10615 , 2_n10616 , 2_n10617 , 2_n10618 , 2_n10619 , 2_n10620 , 2_n10621 , 2_n10622 , 2_n10623 , 2_n10624 , 2_n10625 , 2_n10626 , 2_n10627 , 2_n10628 , 2_n10629 , 2_n10630 , 2_n10631 , 2_n10632 , 2_n10633 , 2_n10634 , 2_n10635 , 2_n10636 , 2_n10637 , 2_n10638 , 2_n10639 , 2_n10640 , 2_n10641 , 2_n10642 , 2_n10643 , 2_n10645 , 2_n10646 , 2_n10647 , 2_n10648 , 2_n10649 , 2_n10650 , 2_n10651 , 2_n10652 , 2_n10653 , 2_n10654 , 2_n10655 , 2_n10656 , 2_n10657 , 2_n10658 , 2_n10659 , 2_n10660 , 2_n10661 , 2_n10662 , 2_n10663 , 2_n10664 , 2_n10665 , 2_n10666 , 2_n10667 , 2_n10668 , 2_n10669 , 2_n10670 , 2_n10671 , 2_n10672 , 2_n10673 , 2_n10674 , 2_n10675 , 2_n10676 , 2_n10677 , 2_n10679 , 2_n10680 , 2_n10681 , 2_n10682 , 2_n10683 , 2_n10684 , 2_n10686 , 2_n10687 , 2_n10688 , 2_n10689 , 2_n10690 , 2_n10691 , 2_n10692 , 2_n10693 , 2_n10694 , 2_n10696 , 2_n10697 , 2_n10698 , 2_n10699 , 2_n10700 , 2_n10701 , 2_n10702 , 2_n10703 , 2_n10704 , 2_n10705 , 2_n10706 , 2_n10707 , 2_n10708 , 2_n10709 , 2_n10710 , 2_n10711 , 2_n10712 , 2_n10713 , 2_n10714 , 2_n10715 , 2_n10716 , 2_n10717 , 2_n10718 , 2_n10719 , 2_n10720 , 2_n10721 , 2_n10722 , 2_n10723 , 2_n10724 , 2_n10725 , 2_n10726 , 2_n10727 , 2_n10728 , 2_n10729 , 2_n10730 , 2_n10731 , 2_n10732 , 2_n10733 , 2_n10734 , 2_n10735 , 2_n10736 , 2_n10737 , 2_n10738 , 2_n10739 , 2_n10740 , 2_n10741 , 2_n10742 , 2_n10743 , 2_n10744 , 2_n10745 , 2_n10746 , 2_n10747 , 2_n10748 , 2_n10749 , 2_n10750 , 2_n10751 , 2_n10752 , 2_n10753 , 2_n10754 , 2_n10755 , 2_n10756 , 2_n10757 , 2_n10758 , 2_n10759 , 2_n10760 , 2_n10761 , 2_n10762 , 2_n10763 , 2_n10764 , 2_n10765 , 2_n10766 , 2_n10767 , 2_n10768 , 2_n10769 , 2_n10770 , 2_n10771 , 2_n10772 , 2_n10773 , 2_n10774 , 2_n10775 , 2_n10776 , 2_n10777 , 2_n10778 , 2_n10779 , 2_n10780 , 2_n10781 , 2_n10782 , 2_n10783 , 2_n10784 , 2_n10785 , 2_n10786 , 2_n10787 , 2_n10788 , 2_n10790 , 2_n10791 , 2_n10792 , 2_n10793 , 2_n10794 , 2_n10795 , 2_n10796 , 2_n10797 , 2_n10798 , 2_n10799 , 2_n10800 , 2_n10801 , 2_n10802 , 2_n10803 , 2_n10804 , 2_n10805 , 2_n10806 , 2_n10807 , 2_n10808 , 2_n10809 , 2_n10810 , 2_n10811 , 2_n10812 , 2_n10813 , 2_n10814 , 2_n10815 , 2_n10816 , 2_n10817 , 2_n10818 , 2_n10819 , 2_n10820 , 2_n10821 , 2_n10822 , 2_n10823 , 2_n10824 , 2_n10825 , 2_n10826 , 2_n10827 , 2_n10828 , 2_n10829 , 2_n10830 , 2_n10831 , 2_n10832 , 2_n10833 , 2_n10834 , 2_n10835 , 2_n10836 , 2_n10837 , 2_n10838 , 2_n10839 , 2_n10840 , 2_n10841 , 2_n10842 , 2_n10843 , 2_n10844 , 2_n10845 , 2_n10846 , 2_n10847 , 2_n10849 , 2_n10850 , 2_n10852 , 2_n10853 , 2_n10854 , 2_n10855 , 2_n10856 , 2_n10857 , 2_n10858 , 2_n10859 , 2_n10860 , 2_n10861 , 2_n10862 , 2_n10863 , 2_n10864 , 2_n10865 , 2_n10866 , 2_n10867 , 2_n10868 , 2_n10869 , 2_n10870 , 2_n10871 , 2_n10872 , 2_n10873 , 2_n10874 , 2_n10875 , 2_n10876 , 2_n10877 , 2_n10878 , 2_n10879 , 2_n10880 , 2_n10881 , 2_n10882 , 2_n10883 , 2_n10884 , 2_n10885 , 2_n10886 , 2_n10887 , 2_n10888 , 2_n10889 , 2_n10890 , 2_n10891 , 2_n10892 , 2_n10893 , 2_n10894 , 2_n10895 , 2_n10896 , 2_n10897 , 2_n10899 , 2_n10900 , 2_n10901 , 2_n10902 , 2_n10903 , 2_n10904 , 2_n10905 , 2_n10906 , 2_n10907 , 2_n10908 , 2_n10909 , 2_n10910 , 2_n10911 , 2_n10912 , 2_n10914 , 2_n10915 , 2_n10916 , 2_n10917 , 2_n10918 , 2_n10919 , 2_n10920 , 2_n10921 , 2_n10922 , 2_n10923 , 2_n10924 , 2_n10925 , 2_n10926 , 2_n10927 , 2_n10929 , 2_n10930 , 2_n10931 , 2_n10932 , 2_n10933 , 2_n10934 , 2_n10935 , 2_n10936 , 2_n10937 , 2_n10938 , 2_n10939 , 2_n10940 , 2_n10941 , 2_n10942 , 2_n10943 , 2_n10944 , 2_n10945 , 2_n10946 , 2_n10947 , 2_n10948 , 2_n10950 , 2_n10951 , 2_n10952 , 2_n10953 , 2_n10954 , 2_n10955 , 2_n10956 , 2_n10957 , 2_n10958 , 2_n10959 , 2_n10960 , 2_n10961 , 2_n10962 , 2_n10963 , 2_n10964 , 2_n10966 , 2_n10967 , 2_n10968 , 2_n10969 , 2_n10970 , 2_n10971 , 2_n10972 , 2_n10973 , 2_n10974 , 2_n10975 , 2_n10976 , 2_n10977 , 2_n10978 , 2_n10979 , 2_n10980 , 2_n10981 , 2_n10982 , 2_n10983 , 2_n10984 , 2_n10985 , 2_n10986 , 2_n10987 , 2_n10988 , 2_n10989 , 2_n10991 , 2_n10992 , 2_n10993 , 2_n10994 , 2_n10995 , 2_n10996 , 2_n10997 , 2_n10998 , 2_n10999 , 2_n11000 , 2_n11001 , 2_n11002 , 2_n11003 , 2_n11004 , 2_n11005 , 2_n11006 , 2_n11007 , 2_n11008 , 2_n11009 , 2_n11010 , 2_n11011 , 2_n11012 , 2_n11013 , 2_n11014 , 2_n11015 , 2_n11016 , 2_n11017 , 2_n11018 , 2_n11019 , 2_n11020 , 2_n11021 , 2_n11022 , 2_n11024 , 2_n11025 , 2_n11026 , 2_n11027 , 2_n11028 , 2_n11029 , 2_n11030 , 2_n11031 , 2_n11032 , 2_n11033 , 2_n11034 , 2_n11035 , 2_n11036 , 2_n11037 , 2_n11038 , 2_n11039 , 2_n11040 , 2_n11041 , 2_n11042 , 2_n11043 , 2_n11044 , 2_n11045 , 2_n11046 , 2_n11047 , 2_n11048 , 2_n11049 , 2_n11050 , 2_n11051 , 2_n11052 , 2_n11053 , 2_n11054 , 2_n11055 , 2_n11056 , 2_n11057 , 2_n11058 , 2_n11059 , 2_n11060 , 2_n11061 , 2_n11062 , 2_n11063 , 2_n11064 , 2_n11065 , 2_n11066 , 2_n11067 , 2_n11068 , 2_n11069 , 2_n11070 , 2_n11071 , 2_n11072 , 2_n11073 , 2_n11074 , 2_n11075 , 2_n11076 , 2_n11077 , 2_n11078 , 2_n11079 , 2_n11080 , 2_n11081 , 2_n11082 , 2_n11083 , 2_n11084 , 2_n11085 , 2_n11086 , 2_n11087 , 2_n11088 , 2_n11089 , 2_n11090 , 2_n11091 , 2_n11092 , 2_n11093 , 2_n11094 , 2_n11095 , 2_n11096 , 2_n11097 , 2_n11098 , 2_n11099 , 2_n11100 , 2_n11101 , 2_n11102 , 2_n11103 , 2_n11104 , 2_n11105 , 2_n11106 , 2_n11107 , 2_n11108 , 2_n11109 , 2_n11110 , 2_n11111 , 2_n11112 , 2_n11113 , 2_n11114 , 2_n11115 , 2_n11116 , 2_n11117 , 2_n11118 , 2_n11119 , 2_n11120 , 2_n11121 , 2_n11122 , 2_n11123 , 2_n11124 , 2_n11125 , 2_n11126 , 2_n11127 , 2_n11128 , 2_n11129 , 2_n11130 , 2_n11131 , 2_n11132 , 2_n11133 , 2_n11134 , 2_n11135 , 2_n11136 , 2_n11137 , 2_n11138 , 2_n11139 , 2_n11140 , 2_n11141 , 2_n11142 , 2_n11143 , 2_n11144 , 2_n11145 , 2_n11146 , 2_n11147 , 2_n11148 , 2_n11149 , 2_n11150 , 2_n11151 , 2_n11152 , 2_n11154 , 2_n11155 , 2_n11156 , 2_n11157 , 2_n11158 , 2_n11159 , 2_n11160 , 2_n11161 , 2_n11162 , 2_n11163 , 2_n11164 , 2_n11165 , 2_n11166 , 2_n11167 , 2_n11168 , 2_n11169 , 2_n11170 , 2_n11171 , 2_n11172 , 2_n11173 , 2_n11174 , 2_n11175 , 2_n11176 , 2_n11177 , 2_n11178 , 2_n11179 , 2_n11180 , 2_n11181 , 2_n11182 , 2_n11183 , 2_n11184 , 2_n11185 , 2_n11186 , 2_n11187 , 2_n11188 , 2_n11189 , 2_n11190 , 2_n11191 , 2_n11192 , 2_n11193 , 2_n11194 , 2_n11195 , 2_n11196 , 2_n11197 , 2_n11198 , 2_n11199 , 2_n11200 , 2_n11201 , 2_n11202 , 2_n11203 , 2_n11204 , 2_n11205 , 2_n11206 , 2_n11207 , 2_n11208 , 2_n11209 , 2_n11210 , 2_n11211 , 2_n11212 , 2_n11213 , 2_n11214 , 2_n11215 , 2_n11217 , 2_n11218 , 2_n11219 , 2_n11220 , 2_n11221 , 2_n11223 , 2_n11224 , 2_n11225 , 2_n11226 , 2_n11227 , 2_n11228 , 2_n11229 , 2_n11230 , 2_n11231 , 2_n11232 , 2_n11233 , 2_n11234 , 2_n11235 , 2_n11236 , 2_n11237 , 2_n11238 , 2_n11239 , 2_n11240 , 2_n11241 , 2_n11242 , 2_n11243 , 2_n11244 , 2_n11245 , 2_n11246 , 2_n11247 , 2_n11248 , 2_n11249 , 2_n11250 , 2_n11251 , 2_n11252 , 2_n11253 , 2_n11254 , 2_n11255 , 2_n11256 , 2_n11258 , 2_n11259 , 2_n11260 , 2_n11261 , 2_n11262 , 2_n11263 , 2_n11264 , 2_n11265 , 2_n11266 , 2_n11267 , 2_n11268 , 2_n11269 , 2_n11270 , 2_n11271 , 2_n11272 , 2_n11273 , 2_n11274 , 2_n11275 , 2_n11276 , 2_n11277 , 2_n11278 , 2_n11279 , 2_n11280 , 2_n11281 , 2_n11282 , 2_n11283 , 2_n11284 , 2_n11285 , 2_n11286 , 2_n11287 , 2_n11288 , 2_n11289 , 2_n11290 , 2_n11291 , 2_n11292 , 2_n11293 , 2_n11294 , 2_n11295 , 2_n11297 , 2_n11298 , 2_n11299 , 2_n11300 , 2_n11301 , 2_n11302 , 2_n11303 , 2_n11304 , 2_n11305 , 2_n11306 , 2_n11307 , 2_n11308 , 2_n11309 , 2_n11310 , 2_n11312 , 2_n11313 , 2_n11314 , 2_n11315 , 2_n11316 , 2_n11317 , 2_n11318 , 2_n11319 , 2_n11320 , 2_n11321 , 2_n11322 , 2_n11323 , 2_n11324 , 2_n11325 , 2_n11327 , 2_n11328 , 2_n11329 , 2_n11330 , 2_n11331 , 2_n11332 , 2_n11333 , 2_n11334 , 2_n11335 , 2_n11336 , 2_n11337 , 2_n11338 , 2_n11339 , 2_n11340 , 2_n11341 , 2_n11342 , 2_n11343 , 2_n11344 , 2_n11345 , 2_n11346 , 2_n11347 , 2_n11348 , 2_n11349 , 2_n11350 , 2_n11351 , 2_n11352 , 2_n11353 , 2_n11354 , 2_n11355 , 2_n11356 , 2_n11357 , 2_n11358 , 2_n11359 , 2_n11360 , 2_n11361 , 2_n11362 , 2_n11363 , 2_n11364 , 2_n11365 , 2_n11366 , 2_n11367 , 2_n11368 , 2_n11369 , 2_n11370 , 2_n11371 , 2_n11372 , 2_n11373 , 2_n11374 , 2_n11375 , 2_n11376 , 2_n11377 , 2_n11378 , 2_n11379 , 2_n11380 , 2_n11381 , 2_n11382 , 2_n11383 , 2_n11384 , 2_n11385 , 2_n11386 , 2_n11387 , 2_n11388 , 2_n11389 , 2_n11390 , 2_n11391 , 2_n11392 , 2_n11393 , 2_n11394 , 2_n11395 , 2_n11396 , 2_n11397 , 2_n11398 , 2_n11399 , 2_n11400 , 2_n11401 , 2_n11402 , 2_n11403 , 2_n11404 , 2_n11405 , 2_n11406 , 2_n11408 , 2_n11409 , 2_n11410 , 2_n11411 , 2_n11412 , 2_n11413 , 2_n11414 , 2_n11415 , 2_n11416 , 2_n11417 , 2_n11418 , 2_n11419 , 2_n11420 , 2_n11421 , 2_n11422 , 2_n11424 , 2_n11425 , 2_n11426 , 2_n11427 , 2_n11428 , 2_n11429 , 2_n11430 , 2_n11431 , 2_n11432 , 2_n11433 , 2_n11434 , 2_n11435 , 2_n11436 , 2_n11437 , 2_n11438 , 2_n11439 , 2_n11440 , 2_n11441 , 2_n11442 , 2_n11443 , 2_n11444 , 2_n11445 , 2_n11446 , 2_n11447 , 2_n11448 , 2_n11449 , 2_n11450 , 2_n11451 , 2_n11452 , 2_n11453 , 2_n11454 , 2_n11455 , 2_n11456 , 2_n11457 , 2_n11458 , 2_n11459 , 2_n11460 , 2_n11461 , 2_n11462 , 2_n11463 , 2_n11464 , 2_n11465 , 2_n11466 , 2_n11467 , 2_n11468 , 2_n11469 , 2_n11470 , 2_n11471 , 2_n11472 , 2_n11473 , 2_n11474 , 2_n11475 , 2_n11476 , 2_n11477 , 2_n11479 , 2_n11480 , 2_n11481 , 2_n11482 , 2_n11483 , 2_n11484 , 2_n11485 , 2_n11486 , 2_n11487 , 2_n11488 , 2_n11489 , 2_n11490 , 2_n11491 , 2_n11492 , 2_n11493 , 2_n11494 , 2_n11495 , 2_n11496 , 2_n11497 , 2_n11498 , 2_n11499 , 2_n11500 , 2_n11501 , 2_n11502 , 2_n11503 , 2_n11504 , 2_n11505 , 2_n11506 , 2_n11507 , 2_n11508 , 2_n11509 , 2_n11510 , 2_n11511 , 2_n11512 , 2_n11513 , 2_n11514 , 2_n11515 , 2_n11516 , 2_n11517 , 2_n11518 , 2_n11519 , 2_n11520 , 2_n11521 , 2_n11522 , 2_n11523 , 2_n11524 , 2_n11525 , 2_n11526 , 2_n11527 , 2_n11528 , 2_n11529 , 2_n11530 , 2_n11531 , 2_n11532 , 2_n11533 , 2_n11534 , 2_n11535 , 2_n11537 , 2_n11538 , 2_n11539 , 2_n11540 , 2_n11541 , 2_n11542 , 2_n11543 , 2_n11544 , 2_n11545 , 2_n11546 , 2_n11547 , 2_n11548 , 2_n11549 , 2_n11550 , 2_n11551 , 2_n11552 , 2_n11553 , 2_n11554 , 2_n11555 , 2_n11556 , 2_n11557 , 2_n11558 , 2_n11559 , 2_n11560 , 2_n11561 , 2_n11562 , 2_n11563 , 2_n11564 , 2_n11565 , 2_n11566 , 2_n11567 , 2_n11568 , 2_n11569 , 2_n11570 , 2_n11571 , 2_n11572 , 2_n11573 , 2_n11574 , 2_n11575 , 2_n11576 , 2_n11577 , 2_n11578 , 2_n11579 , 2_n11580 , 2_n11581 , 2_n11582 , 2_n11583 , 2_n11584 , 2_n11585 , 2_n11586 , 2_n11587 , 2_n11588 , 2_n11589 , 2_n11590 , 2_n11591 , 2_n11592 , 2_n11593 , 2_n11594 , 2_n11595 , 2_n11596 , 2_n11597 , 2_n11598 , 2_n11599 , 2_n11600 , 2_n11601 , 2_n11602 , 2_n11603 , 2_n11604 , 2_n11605 , 2_n11606 , 2_n11607 , 2_n11608 , 2_n11609 , 2_n11610 , 2_n11611 , 2_n11612 , 2_n11613 , 2_n11614 , 2_n11615 , 2_n11616 , 2_n11617 , 2_n11618 , 2_n11619 , 2_n11620 , 2_n11621 , 2_n11622 , 2_n11623 , 2_n11624 , 2_n11625 , 2_n11626 , 2_n11627 , 2_n11628 , 2_n11629 , 2_n11630 , 2_n11631 , 2_n11632 , 2_n11633 , 2_n11634 , 2_n11635 , 2_n11636 , 2_n11637 , 2_n11638 , 2_n11639 , 2_n11640 , 2_n11641 , 2_n11642 , 2_n11643 , 2_n11644 , 2_n11645 , 2_n11646 , 2_n11647 , 2_n11648 , 2_n11649 , 2_n11650 , 2_n11651 , 2_n11652 , 2_n11653 , 2_n11654 , 2_n11655 , 2_n11656 , 2_n11657 , 2_n11658 , 2_n11659 , 2_n11660 , 2_n11661 , 2_n11663 , 2_n11664 , 2_n11665 , 2_n11666 , 2_n11667 , 2_n11668 , 2_n11669 , 2_n11670 , 2_n11671 , 2_n11672 , 2_n11673 , 2_n11674 , 2_n11675 , 2_n11676 , 2_n11677 , 2_n11678 , 2_n11679 , 2_n11680 , 2_n11681 , 2_n11682 , 2_n11683 , 2_n11684 , 2_n11685 , 2_n11686 , 2_n11687 , 2_n11688 , 2_n11689 , 2_n11690 , 2_n11691 , 2_n11692 , 2_n11693 , 2_n11694 , 2_n11695 , 2_n11696 , 2_n11697 , 2_n11698 , 2_n11699 , 2_n11700 , 2_n11701 , 2_n11702 , 2_n11703 , 2_n11704 , 2_n11705 , 2_n11706 , 2_n11708 , 2_n11709 , 2_n11710 , 2_n11711 , 2_n11712 , 2_n11713 , 2_n11714 , 2_n11715 , 2_n11716 , 2_n11717 , 2_n11718 , 2_n11719 , 2_n11720 , 2_n11721 , 2_n11722 , 2_n11723 , 2_n11724 , 2_n11725 , 2_n11726 , 2_n11727 , 2_n11729 , 2_n11730 , 2_n11731 , 2_n11732 , 2_n11733 , 2_n11734 , 2_n11735 , 2_n11736 , 2_n11737 , 2_n11738 , 2_n11739 , 2_n11740 , 2_n11741 , 2_n11742 , 2_n11743 , 2_n11744 , 2_n11745 , 2_n11746 , 2_n11747 , 2_n11748 , 2_n11749 , 2_n11750 , 2_n11751 , 2_n11752 , 2_n11753 , 2_n11754 , 2_n11756 , 2_n11758 , 2_n11759 , 2_n11760 , 2_n11761 , 2_n11762 , 2_n11763 , 2_n11764 , 2_n11765 , 2_n11766 , 2_n11767 , 2_n11768 , 2_n11769 , 2_n11770 , 2_n11771 , 2_n11772 , 2_n11773 , 2_n11774 , 2_n11775 , 2_n11776 , 2_n11777 , 2_n11778 , 2_n11779 , 2_n11781 , 2_n11782 , 2_n11783 , 2_n11784 , 2_n11785 , 2_n11786 , 2_n11787 , 2_n11788 , 2_n11789 , 2_n11790 , 2_n11792 , 2_n11793 , 2_n11794 , 2_n11795 , 2_n11796 , 2_n11797 , 2_n11798 , 2_n11799 , 2_n11800 , 2_n11801 , 2_n11802 , 2_n11803 , 2_n11804 , 2_n11805 , 2_n11806 , 2_n11807 , 2_n11808 , 2_n11809 , 2_n11810 , 2_n11811 , 2_n11812 , 2_n11813 , 2_n11814 , 2_n11815 , 2_n11816 , 2_n11817 , 2_n11818 , 2_n11819 , 2_n11820 , 2_n11822 , 2_n11823 , 2_n11824 , 2_n11825 , 2_n11826 , 2_n11827 , 2_n11828 , 2_n11829 , 2_n11830 , 2_n11831 , 2_n11832 , 2_n11833 , 2_n11834 , 2_n11835 , 2_n11836 , 2_n11837 , 2_n11838 , 2_n11839 , 2_n11840 , 2_n11841 , 2_n11842 , 2_n11843 , 2_n11844 , 2_n11845 , 2_n11846 , 2_n11847 , 2_n11848 , 2_n11849 , 2_n11850 , 2_n11851 , 2_n11852 , 2_n11853 , 2_n11854 , 2_n11855 , 2_n11856 , 2_n11857 , 2_n11858 , 2_n11859 , 2_n11860 , 2_n11861 , 2_n11862 , 2_n11863 , 2_n11864 , 2_n11865 , 2_n11866 , 2_n11867 , 2_n11868 , 2_n11869 , 2_n11870 , 2_n11871 , 2_n11872 , 2_n11873 , 2_n11874 , 2_n11875 , 2_n11878 , 2_n11879 , 2_n11880 , 2_n11881 , 2_n11882 , 2_n11883 , 2_n11884 , 2_n11885 , 2_n11886 , 2_n11887 , 2_n11888 , 2_n11889 , 2_n11890 , 2_n11891 , 2_n11893 , 2_n11894 , 2_n11895 , 2_n11896 , 2_n11897 , 2_n11898 , 2_n11899 , 2_n11900 , 2_n11901 , 2_n11902 , 2_n11903 , 2_n11904 , 2_n11905 , 2_n11906 , 2_n11907 , 2_n11908 , 2_n11909 , 2_n11910 , 2_n11911 , 2_n11912 , 2_n11913 , 2_n11914 , 2_n11915 , 2_n11916 , 2_n11918 , 2_n11920 , 2_n11921 , 2_n11923 , 2_n11924 , 2_n11925 , 2_n11926 , 2_n11927 , 2_n11928 , 2_n11929 , 2_n11930 , 2_n11931 , 2_n11932 , 2_n11933 , 2_n11934 , 2_n11935 , 2_n11936 , 2_n11937 , 2_n11938 , 2_n11939 , 2_n11940 , 2_n11941 , 2_n11942 , 2_n11943 , 2_n11944 , 2_n11945 , 2_n11946 , 2_n11947 , 2_n11948 , 2_n11949 , 2_n11950 , 2_n11951 , 2_n11952 , 2_n11953 , 2_n11954 , 2_n11955 , 2_n11956 , 2_n11957 , 2_n11958 , 2_n11959 , 2_n11960 , 2_n11961 , 2_n11962 , 2_n11963 , 2_n11964 , 2_n11965 , 2_n11966 , 2_n11968 , 2_n11969 , 2_n11970 , 2_n11971 , 2_n11972 , 2_n11973 , 2_n11974 , 2_n11975 , 2_n11976 , 2_n11977 , 2_n11978 , 2_n11979 , 2_n11980 , 2_n11981 , 2_n11982 , 2_n11983 , 2_n11984 , 2_n11985 , 2_n11986 , 2_n11987 , 2_n11988 , 2_n11989 , 2_n11990 , 2_n11991 , 2_n11992 , 2_n11993 , 2_n11994 , 2_n11995 , 2_n11996 , 2_n11997 , 2_n11998 , 2_n12001 , 2_n12002 , 2_n12003 , 2_n12004 , 2_n12006 , 2_n12007 , 2_n12008 , 2_n12009 , 2_n12010 , 2_n12011 , 2_n12012 , 2_n12013 , 2_n12015 , 2_n12016 , 2_n12017 , 2_n12018 , 2_n12019 , 2_n12021 , 2_n12022 , 2_n12023 , 2_n12024 , 2_n12026 , 2_n12027 , 2_n12028 , 2_n12029 , 2_n12030 , 2_n12031 , 2_n12032 , 2_n12033 , 2_n12034 , 2_n12035 , 2_n12036 , 2_n12037 , 2_n12038 , 2_n12039 , 2_n12040 , 2_n12041 , 2_n12042 , 2_n12043 , 2_n12045 , 2_n12046 , 2_n12047 , 2_n12048 , 2_n12049 , 2_n12050 , 2_n12051 , 2_n12052 , 2_n12053 , 2_n12054 , 2_n12055 , 2_n12056 , 2_n12057 , 2_n12058 , 2_n12059 , 2_n12060 , 2_n12061 , 2_n12062 , 2_n12063 , 2_n12064 , 2_n12065 , 2_n12066 , 2_n12067 , 2_n12068 , 2_n12070 , 2_n12071 , 2_n12072 , 2_n12073 , 2_n12074 , 2_n12075 , 2_n12077 , 2_n12078 , 2_n12079 , 2_n12080 , 2_n12081 , 2_n12082 , 2_n12083 , 2_n12084 , 2_n12085 , 2_n12086 , 2_n12087 , 2_n12088 , 2_n12089 , 2_n12090 , 2_n12091 , 2_n12092 , 2_n12093 , 2_n12094 , 2_n12095 , 2_n12096 , 2_n12097 , 2_n12098 , 2_n12099 , 2_n12100 , 2_n12101 , 2_n12102 , 2_n12103 , 2_n12104 , 2_n12105 , 2_n12106 , 2_n12107 , 2_n12108 , 2_n12109 , 2_n12110 , 2_n12112 , 2_n12113 , 2_n12114 , 2_n12115 , 2_n12116 , 2_n12117 , 2_n12118 , 2_n12119 , 2_n12120 , 2_n12121 , 2_n12122 , 2_n12123 , 2_n12124 , 2_n12125 , 2_n12126 , 2_n12127 , 2_n12128 , 2_n12129 , 2_n12130 , 2_n12131 , 2_n12132 , 2_n12133 , 2_n12134 , 2_n12135 , 2_n12136 , 2_n12137 , 2_n12138 , 2_n12139 , 2_n12140 , 2_n12141 , 2_n12142 , 2_n12143 , 2_n12144 , 2_n12146 , 2_n12147 , 2_n12148 , 2_n12149 , 2_n12150 , 2_n12151 , 2_n12152 , 2_n12153 , 2_n12154 , 2_n12155 , 2_n12156 , 2_n12157 , 2_n12158 , 2_n12159 , 2_n12160 , 2_n12161 , 2_n12162 , 2_n12163 , 2_n12164 , 2_n12165 , 2_n12166 , 2_n12167 , 2_n12168 , 2_n12169 , 2_n12170 , 2_n12171 , 2_n12172 , 2_n12173 , 2_n12174 , 2_n12175 , 2_n12176 , 2_n12177 , 2_n12178 , 2_n12179 , 2_n12180 , 2_n12181 , 2_n12182 , 2_n12183 , 2_n12184 , 2_n12185 , 2_n12186 , 2_n12187 , 2_n12188 , 2_n12189 , 2_n12190 , 2_n12191 , 2_n12192 , 2_n12193 , 2_n12194 , 2_n12195 , 2_n12196 , 2_n12197 , 2_n12198 , 2_n12199 , 2_n12200 , 2_n12201 , 2_n12202 , 2_n12203 , 2_n12204 , 2_n12205 , 2_n12206 , 2_n12207 , 2_n12208 , 2_n12209 , 2_n12210 , 2_n12211 , 2_n12212 , 2_n12213 , 2_n12214 , 2_n12215 , 2_n12216 , 2_n12217 , 2_n12218 , 2_n12219 , 2_n12220 , 2_n12222 , 2_n12223 , 2_n12224 , 2_n12225 , 2_n12226 , 2_n12227 , 2_n12228 , 2_n12229 , 2_n12230 , 2_n12231 , 2_n12232 , 2_n12233 , 2_n12234 , 2_n12235 , 2_n12236 , 2_n12237 , 2_n12238 , 2_n12239 , 2_n12240 , 2_n12241 , 2_n12242 , 2_n12243 , 2_n12244 , 2_n12245 , 2_n12246 , 2_n12248 , 2_n12249 , 2_n12250 , 2_n12251 , 2_n12252 , 2_n12253 , 2_n12254 , 2_n12255 , 2_n12256 , 2_n12257 , 2_n12258 , 2_n12259 , 2_n12260 , 2_n12261 , 2_n12262 , 2_n12263 , 2_n12264 , 2_n12265 , 2_n12266 , 2_n12267 , 2_n12268 , 2_n12269 , 2_n12270 , 2_n12271 , 2_n12272 , 2_n12273 , 2_n12274 , 2_n12275 , 2_n12276 , 2_n12277 , 2_n12278 , 2_n12279 , 2_n12280 , 2_n12281 , 2_n12282 , 2_n12283 , 2_n12284 , 2_n12285 , 2_n12286 , 2_n12287 , 2_n12288 , 2_n12289 , 2_n12290 , 2_n12291 , 2_n12292 , 2_n12293 , 2_n12294 , 2_n12295 , 2_n12296 , 2_n12297 , 2_n12298 , 2_n12300 , 2_n12301 , 2_n12302 , 2_n12303 , 2_n12304 , 2_n12305 , 2_n12306 , 2_n12307 , 2_n12308 , 2_n12309 , 2_n12310 , 2_n12311 , 2_n12312 , 2_n12313 , 2_n12314 , 2_n12315 , 2_n12316 , 2_n12317 , 2_n12318 , 2_n12319 , 2_n12320 , 2_n12321 , 2_n12322 , 2_n12323 , 2_n12324 , 2_n12325 , 2_n12326 , 2_n12327 , 2_n12328 , 2_n12329 , 2_n12330 , 2_n12331 , 2_n12332 , 2_n12333 , 2_n12334 , 2_n12335 , 2_n12336 , 2_n12337 , 2_n12338 , 2_n12339 , 2_n12340 , 2_n12341 , 2_n12342 , 2_n12343 , 2_n12344 , 2_n12345 , 2_n12346 , 2_n12347 , 2_n12348 , 2_n12349 , 2_n12350 , 2_n12351 , 2_n12352 , 2_n12353 , 2_n12354 , 2_n12355 , 2_n12356 , 2_n12357 , 2_n12358 , 2_n12359 , 2_n12360 , 2_n12361 , 2_n12362 , 2_n12363 , 2_n12364 , 2_n12365 , 2_n12366 , 2_n12367 , 2_n12368 , 2_n12369 , 2_n12370 , 2_n12371 , 2_n12372 , 2_n12373 , 2_n12374 , 2_n12375 , 2_n12376 , 2_n12377 , 2_n12378 , 2_n12379 , 2_n12380 , 2_n12381 , 2_n12382 , 2_n12383 , 2_n12384 , 2_n12385 , 2_n12386 , 2_n12387 , 2_n12388 , 2_n12389 , 2_n12390 , 2_n12392 , 2_n12393 , 2_n12394 , 2_n12395 , 2_n12396 , 2_n12397 , 2_n12398 , 2_n12399 , 2_n12400 , 2_n12401 , 2_n12402 , 2_n12403 , 2_n12404 , 2_n12405 , 2_n12406 , 2_n12407 , 2_n12408 , 2_n12409 , 2_n12410 , 2_n12411 , 2_n12412 , 2_n12413 , 2_n12414 , 2_n12415 , 2_n12416 , 2_n12417 , 2_n12418 , 2_n12419 , 2_n12420 , 2_n12421 , 2_n12422 , 2_n12423 , 2_n12424 , 2_n12425 , 2_n12426 , 2_n12427 , 2_n12428 , 2_n12429 , 2_n12430 , 2_n12431 , 2_n12432 , 2_n12433 , 2_n12434 , 2_n12435 , 2_n12436 , 2_n12437 , 2_n12438 , 2_n12439 , 2_n12440 , 2_n12441 , 2_n12442 , 2_n12443 , 2_n12445 , 2_n12446 , 2_n12447 , 2_n12448 , 2_n12449 , 2_n12450 , 2_n12451 , 2_n12452 , 2_n12453 , 2_n12454 , 2_n12455 , 2_n12456 , 2_n12457 , 2_n12458 , 2_n12459 , 2_n12460 , 2_n12461 , 2_n12462 , 2_n12463 , 2_n12464 , 2_n12465 , 2_n12466 , 2_n12467 , 2_n12468 , 2_n12469 , 2_n12470 , 2_n12471 , 2_n12472 , 2_n12473 , 2_n12474 , 2_n12475 , 2_n12476 , 2_n12477 , 2_n12478 , 2_n12479 , 2_n12480 , 2_n12481 , 2_n12482 , 2_n12483 , 2_n12484 , 2_n12485 , 2_n12486 , 2_n12487 , 2_n12488 , 2_n12490 , 2_n12491 , 2_n12492 , 2_n12493 , 2_n12494 , 2_n12495 , 2_n12496 , 2_n12497 , 2_n12498 , 2_n12499 , 2_n12500 , 2_n12501 , 2_n12502 , 2_n12503 , 2_n12504 , 2_n12505 , 2_n12506 , 2_n12507 , 2_n12508 , 2_n12509 , 2_n12510 , 2_n12512 , 2_n12513 , 2_n12514 , 2_n12515 , 2_n12516 , 2_n12517 , 2_n12518 , 2_n12519 , 2_n12520 , 2_n12521 , 2_n12522 , 2_n12523 , 2_n12524 , 2_n12525 , 2_n12526 , 2_n12527 , 2_n12528 , 2_n12529 , 2_n12530 , 2_n12531 , 2_n12532 , 2_n12533 , 2_n12534 , 2_n12535 , 2_n12536 , 2_n12537 , 2_n12538 , 2_n12539 , 2_n12540 , 2_n12541 , 2_n12542 , 2_n12543 , 2_n12544 , 2_n12545 , 2_n12546 , 2_n12547 , 2_n12548 , 2_n12549 , 2_n12550 , 2_n12551 , 2_n12552 , 2_n12553 , 2_n12554 , 2_n12555 , 2_n12556 , 2_n12557 , 2_n12558 , 2_n12559 , 2_n12560 , 2_n12561 , 2_n12562 , 2_n12563 , 2_n12564 , 2_n12565 , 2_n12566 , 2_n12567 , 2_n12568 , 2_n12569 , 2_n12570 , 2_n12571 , 2_n12572 , 2_n12573 , 2_n12574 , 2_n12575 , 2_n12576 , 2_n12577 , 2_n12578 , 2_n12579 , 2_n12580 , 2_n12581 , 2_n12582 , 2_n12583 , 2_n12584 , 2_n12585 , 2_n12586 , 2_n12587 , 2_n12588 , 2_n12589 , 2_n12590 , 2_n12592 , 2_n12593 , 2_n12594 , 2_n12595 , 2_n12596 , 2_n12597 , 2_n12598 , 2_n12599 , 2_n12600 , 2_n12601 , 2_n12602 , 2_n12603 , 2_n12604 , 2_n12605 , 2_n12606 , 2_n12607 , 2_n12608 , 2_n12609 , 2_n12610 , 2_n12611 , 2_n12612 , 2_n12613 , 2_n12614 , 2_n12615 , 2_n12616 , 2_n12617 , 2_n12618 , 2_n12619 , 2_n12620 , 2_n12621 , 2_n12622 , 2_n12623 , 2_n12624 , 2_n12625 , 2_n12626 , 2_n12627 , 2_n12628 , 2_n12629 , 2_n12630 , 2_n12631 , 2_n12632 , 2_n12633 , 2_n12634 , 2_n12635 , 2_n12636 , 2_n12637 , 2_n12638 , 2_n12639 , 2_n12640 , 2_n12641 , 2_n12642 , 2_n12643 , 2_n12644 , 2_n12645 , 2_n12646 , 2_n12647 , 2_n12649 , 2_n12650 , 2_n12651 , 2_n12652 , 2_n12653 , 2_n12654 , 2_n12655 , 2_n12656 , 2_n12657 , 2_n12658 , 2_n12659 , 2_n12660 , 2_n12661 , 2_n12662 , 2_n12663 , 2_n12664 , 2_n12665 , 2_n12666 , 2_n12667 , 2_n12668 , 2_n12669 , 2_n12670 , 2_n12671 , 2_n12672 , 2_n12673 , 2_n12674 , 2_n12675 , 2_n12676 , 2_n12677 , 2_n12678 , 2_n12679 , 2_n12680 , 2_n12681 , 2_n12682 , 2_n12683 , 2_n12684 , 2_n12685 , 2_n12686 , 2_n12687 , 2_n12688 , 2_n12689 , 2_n12690 , 2_n12691 , 2_n12692 , 2_n12693 , 2_n12694 , 2_n12695 , 2_n12696 , 2_n12697 , 2_n12698 , 2_n12699 , 2_n12700 , 2_n12701 , 2_n12702 , 2_n12703 , 2_n12707 , 2_n12708 , 2_n12710 , 2_n12711 , 2_n12712 , 2_n12713 , 2_n12714 , 2_n12715 , 2_n12716 , 2_n12717 , 2_n12718 , 2_n12719 , 2_n12721 , 2_n12722 , 2_n12723 , 2_n12724 , 2_n12725 , 2_n12726 , 2_n12727 , 2_n12728 , 2_n12729 , 2_n12730 , 2_n12731 , 2_n12732 , 2_n12733 , 2_n12734 , 2_n12735 , 2_n12736 , 2_n12737 , 2_n12738 , 2_n12739 , 2_n12740 , 2_n12741 , 2_n12742 , 2_n12743 , 2_n12744 , 2_n12745 , 2_n12746 , 2_n12747 , 2_n12748 , 2_n12749 , 2_n12750 , 2_n12751 , 2_n12752 , 2_n12754 , 2_n12755 , 2_n12756 , 2_n12757 , 2_n12758 , 2_n12759 , 2_n12760 , 2_n12761 , 2_n12762 , 2_n12763 , 2_n12764 , 2_n12765 , 2_n12766 , 2_n12767 , 2_n12768 , 2_n12769 , 2_n12770 , 2_n12771 , 2_n12772 , 2_n12773 , 2_n12774 , 2_n12775 , 2_n12776 , 2_n12778 , 2_n12779 , 2_n12780 , 2_n12781 , 2_n12782 , 2_n12783 , 2_n12784 , 2_n12785 , 2_n12786 , 2_n12787 , 2_n12788 , 2_n12789 , 2_n12790 , 2_n12791 , 2_n12792 , 2_n12793 , 2_n12794 , 2_n12795 , 2_n12796 , 2_n12797 , 2_n12798 , 2_n12799 , 2_n12800 , 2_n12801 , 2_n12802 , 2_n12803 , 2_n12804 , 2_n12805 , 2_n12806 , 2_n12808 , 2_n12809 , 2_n12810 , 2_n12811 , 2_n12812 , 2_n12813 , 2_n12814 , 2_n12815 , 2_n12816 , 2_n12817 , 2_n12818 , 2_n12819 , 2_n12820 , 2_n12821 , 2_n12822 , 2_n12823 , 2_n12824 , 2_n12825 , 2_n12827 , 2_n12828 , 2_n12829 , 2_n12830 , 2_n12831 , 2_n12832 , 2_n12833 , 2_n12834 , 2_n12835 , 2_n12836 , 2_n12837 , 2_n12838 , 2_n12839 , 2_n12840 , 2_n12841 , 2_n12842 , 2_n12843 , 2_n12844 , 2_n12845 , 2_n12846 , 2_n12847 , 2_n12848 , 2_n12849 , 2_n12850 , 2_n12851 , 2_n12852 , 2_n12853 , 2_n12854 , 2_n12855 , 2_n12856 , 2_n12857 , 2_n12858 , 2_n12859 , 2_n12860 , 2_n12861 , 2_n12862 , 2_n12863 , 2_n12864 , 2_n12865 , 2_n12866 , 2_n12867 , 2_n12868 , 2_n12869 , 2_n12870 , 2_n12871 , 2_n12872 , 2_n12873 , 2_n12874 , 2_n12875 , 2_n12876 , 2_n12877 , 2_n12878 , 2_n12879 , 2_n12880 , 2_n12881 , 2_n12882 , 2_n12883 , 2_n12884 , 2_n12885 , 2_n12886 , 2_n12887 , 2_n12888 , 2_n12889 , 2_n12890 , 2_n12891 , 2_n12892 , 2_n12893 , 2_n12894 , 2_n12895 , 2_n12896 , 2_n12897 , 2_n12898 , 2_n12899 , 2_n12900 , 2_n12901 , 2_n12902 , 2_n12903 , 2_n12904 , 2_n12905 , 2_n12906 , 2_n12907 , 2_n12908 , 2_n12909 , 2_n12910 , 2_n12911 , 2_n12912 , 2_n12913 , 2_n12914 , 2_n12915 , 2_n12916 , 2_n12917 , 2_n12918 , 2_n12919 , 2_n12920 , 2_n12921 , 2_n12922 , 2_n12923 , 2_n12924 , 2_n12926 , 2_n12927 , 2_n12928 , 2_n12929 , 2_n12930 , 2_n12931 , 2_n12932 , 2_n12933 , 2_n12934 , 2_n12935 , 2_n12936 , 2_n12937 , 2_n12938 , 2_n12939 , 2_n12940 , 2_n12941 , 2_n12942 , 2_n12943 , 2_n12944 , 2_n12945 , 2_n12946 , 2_n12948 , 2_n12949 , 2_n12950 , 2_n12951 , 2_n12952 , 2_n12953 , 2_n12954 , 2_n12955 , 2_n12956 , 2_n12957 , 2_n12958 , 2_n12959 , 2_n12960 ;
assign 2_n2141 = 2_n2530 & 2_n521;
assign 2_n206 = ~(2_n491 ^ 2_n5906);
assign 2_n3102 = 2_n4112 & 2_n2282;
assign 2_n2523 = 2_n12144 | 2_n5251;
assign 2_n2468 = 2_n491 | 2_n9006;
assign 2_n5935 = ~(2_n5205 | 2_n1662);
assign 2_n12452 = 2_n3831 & 2_n6309;
assign 2_n3584 = 2_n9389 | 2_n6402;
assign 2_n12769 = ~(2_n12488 ^ 2_n2077);
assign 2_n9132 = ~(2_n8037 ^ 2_n4937);
assign 2_n8628 = ~(2_n8093 ^ 2_n65);
assign 2_n7698 = ~(2_n8387 ^ 2_n966);
assign 2_n490 = ~2_n5531;
assign 2_n999 = 2_n9750 | 2_n4371;
assign 2_n5811 = ~(2_n7893 | 2_n291);
assign 2_n4271 = ~(2_n3168 | 2_n10348);
assign 2_n12068 = 2_n636 | 2_n12735;
assign 2_n2076 = ~2_n12706;
assign 2_n10627 = ~(2_n9510 ^ 2_n851);
assign 2_n8741 = ~(2_n5885 ^ 2_n10164);
assign 2_n6963 = 2_n9723 | 2_n12736;
assign 2_n5770 = 2_n10925 | 2_n11911;
assign 2_n2237 = ~(2_n6664 ^ 2_n8627);
assign 2_n7708 = ~2_n10979;
assign 2_n8228 = 2_n6073 & 2_n8947;
assign 2_n8420 = ~(2_n6208 ^ 2_n6269);
assign 2_n1335 = ~2_n12713;
assign 2_n6572 = ~(2_n1342 | 2_n7497);
assign 2_n12308 = ~(2_n5629 ^ 2_n8716);
assign 2_n3369 = 2_n12792 & 2_n2220;
assign 2_n3113 = ~(2_n9048 ^ 2_n5993);
assign 2_n5819 = ~(2_n10889 ^ 2_n7455);
assign 2_n5150 = ~(2_n7321 ^ 2_n2104);
assign 2_n6886 = 2_n9202 & 2_n7379;
assign 2_n6118 = ~(2_n10013 ^ 2_n9298);
assign 2_n171 = ~2_n8009;
assign 2_n10492 = 2_n638 & 2_n7227;
assign 2_n9668 = ~(2_n2213 ^ 2_n1443);
assign 2_n10042 = 2_n7236 & 2_n11876;
assign 2_n12212 = 2_n1392 & 2_n2337;
assign 2_n3581 = 2_n11073 | 2_n5965;
assign 2_n6875 = 2_n246 & 2_n5633;
assign 2_n12285 = ~(2_n1762 | 2_n5238);
assign 2_n2936 = 2_n8903 | 2_n5834;
assign 2_n8724 = ~(2_n11543 ^ 2_n924);
assign 2_n11838 = 2_n989 | 2_n1546;
assign 2_n4629 = ~(2_n11708 ^ 2_n11243);
assign 2_n4319 = 2_n7130 | 2_n2371;
assign 2_n8111 = 2_n12237 | 2_n12535;
assign 2_n6562 = ~(2_n11596 ^ 2_n5864);
assign 2_n2487 = 2_n1989 & 2_n3600;
assign 2_n6692 = ~(2_n10970 ^ 2_n11448);
assign 2_n3458 = ~(2_n2834 ^ 2_n2017);
assign 2_n10494 = ~(2_n638 ^ 2_n1446);
assign 2_n2545 = ~(2_n9828 ^ 2_n952);
assign 2_n9965 = ~(2_n5371 ^ 2_n1780);
assign 2_n8178 = ~(2_n5532 | 2_n2604);
assign 2_n11147 = 2_n11923 | 2_n4527;
assign 2_n1622 = ~(2_n4430 ^ 2_n2054);
assign 2_n1082 = 2_n11026 | 2_n10916;
assign 2_n8348 = 2_n2099 | 2_n1163;
assign 2_n8486 = 2_n3207 & 2_n10957;
assign 2_n1757 = 2_n7749 | 2_n8602;
assign 2_n10124 = 2_n4250 | 2_n7101;
assign 2_n2478 = ~(2_n3943 | 2_n7708);
assign 2_n1228 = ~(2_n9428 ^ 2_n9981);
assign 2_n4157 = ~(2_n8423 ^ 2_n7315);
assign 2_n8463 = ~(2_n3767 ^ 2_n8601);
assign 2_n9317 = ~(2_n2340 ^ 2_n6152);
assign 2_n8303 = 2_n5732 ^ 2_n5336;
assign 2_n10085 = 2_n9122 & 2_n4460;
assign 2_n8631 = 2_n242 | 2_n12250;
assign 2_n10958 = ~(2_n3380 | 2_n4252);
assign 2_n1579 = 2_n1699 | 2_n6071;
assign 2_n5316 = 2_n4358 & 2_n10165;
assign 2_n10473 = ~(2_n9382 ^ 2_n3001);
assign 2_n2321 = 2_n8428 | 2_n2815;
assign 2_n4965 = 2_n9271 & 2_n1866;
assign 2_n3103 = 2_n7916 & 2_n2642;
assign 2_n8152 = ~2_n5213;
assign 2_n3034 = ~(2_n8018 ^ 2_n744);
assign 2_n10839 = 2_n9370 | 2_n12328;
assign 2_n10454 = ~(2_n1661 ^ 2_n6545);
assign 2_n10310 = 2_n4175 | 2_n457;
assign 2_n6142 = 2_n1653 | 2_n10896;
assign 2_n4910 = ~(2_n6400 ^ 2_n2360);
assign 2_n8690 = ~2_n7121;
assign 2_n10461 = 2_n6718 | 2_n12120;
assign 2_n11803 = ~2_n6866;
assign 2_n372 = 2_n5350 & 2_n3540;
assign 2_n9377 = ~2_n6787;
assign 2_n4958 = 2_n9561 | 2_n11702;
assign 2_n6911 = 2_n1937 | 2_n12816;
assign 2_n8730 = 2_n6510 | 2_n49;
assign 2_n2061 = ~(2_n5956 ^ 2_n2369);
assign 2_n11117 = ~(2_n1930 ^ 2_n9047);
assign 2_n2307 = 2_n3655 & 2_n4653;
assign 2_n12594 = ~(2_n7659 | 2_n9923);
assign 2_n8651 = ~(2_n6335 ^ 2_n5728);
assign 2_n7187 = 2_n8623 & 2_n7113;
assign 2_n2050 = ~2_n8938;
assign 2_n3442 = 2_n3127 | 2_n10419;
assign 2_n5257 = ~(2_n10357 ^ 2_n5568);
assign 2_n5834 = 2_n5489 & 2_n10173;
assign 2_n2462 = ~(2_n4717 ^ 2_n12433);
assign 2_n7483 = ~(2_n3418 ^ 2_n2490);
assign 2_n7076 = 2_n3218 | 2_n3846;
assign 2_n4520 = ~(2_n1033 ^ 2_n617);
assign 2_n5455 = ~2_n11016;
assign 2_n9277 = 2_n12138 | 2_n7132;
assign 2_n12377 = ~(2_n11098 | 2_n2315);
assign 2_n11028 = ~(2_n1179 | 2_n7664);
assign 2_n1103 = ~(2_n12125 ^ 2_n1204);
assign 2_n12342 = 2_n11892 & 2_n217;
assign 2_n6480 = ~(2_n2246 ^ 2_n9569);
assign 2_n9422 = ~2_n8937;
assign 2_n4639 = ~(2_n3509 | 2_n727);
assign 2_n221 = ~(2_n5107 | 2_n258);
assign 2_n9126 = 2_n2956 | 2_n6653;
assign 2_n11397 = ~(2_n842 ^ 2_n10764);
assign 2_n1049 = 2_n12442 | 2_n10382;
assign 2_n3740 = ~2_n6165;
assign 2_n1169 = 2_n4760 & 2_n10105;
assign 2_n12150 = 2_n8181 & 2_n8485;
assign 2_n4048 = ~2_n11265;
assign 2_n2984 = 2_n10904 | 2_n126;
assign 2_n8290 = 2_n1183 | 2_n10854;
assign 2_n8158 = ~2_n5745;
assign 2_n6389 = ~2_n2879;
assign 2_n7837 = 2_n295 | 2_n8415;
assign 2_n9153 = ~(2_n9388 ^ 2_n6619);
assign 2_n5683 = ~2_n4809;
assign 2_n3724 = 2_n12398 | 2_n4655;
assign 2_n1355 = 2_n9512 & 2_n5173;
assign 2_n8260 = 2_n3127 | 2_n8524;
assign 2_n12831 = 2_n2099 | 2_n12441;
assign 2_n8029 = ~(2_n6075 ^ 2_n12581);
assign 2_n7347 = 2_n2671 | 2_n9678;
assign 2_n8443 = ~(2_n4210 | 2_n5871);
assign 2_n8006 = 2_n1146 | 2_n8593;
assign 2_n12126 = ~(2_n7468 ^ 2_n271);
assign 2_n7882 = ~(2_n8058 ^ 2_n6323);
assign 2_n4258 = ~(2_n8581 ^ 2_n4231);
assign 2_n8100 = ~(2_n750 ^ 2_n863);
assign 2_n2201 = 2_n6577 | 2_n8414;
assign 2_n1179 = ~2_n7009;
assign 2_n9690 = 2_n8042 | 2_n1905;
assign 2_n9775 = 2_n7843 & 2_n3005;
assign 2_n8929 = ~2_n2945;
assign 2_n8182 = ~(2_n2474 | 2_n6830);
assign 2_n1955 = 2_n4456 | 2_n10442;
assign 2_n11129 = 2_n5659 | 2_n366;
assign 2_n7119 = 2_n12862 & 2_n5595;
assign 2_n661 = 2_n6349 | 2_n8350;
assign 2_n3565 = 2_n4744 & 2_n171;
assign 2_n3098 = ~2_n9572;
assign 2_n7791 = 2_n11923 | 2_n9078;
assign 2_n8763 = 2_n11892 & 2_n2749;
assign 2_n9184 = ~(2_n9621 ^ 2_n1490);
assign 2_n1142 = ~(2_n2600 | 2_n12332);
assign 2_n10231 = 2_n9878 | 2_n10854;
assign 2_n6119 = 2_n7046 & 2_n11778;
assign 2_n3993 = 2_n1998 & 2_n6081;
assign 2_n9684 = ~(2_n10144 ^ 2_n10484);
assign 2_n7261 = 2_n10546 | 2_n1307;
assign 2_n5800 = 2_n3757 | 2_n10363;
assign 2_n12481 = 2_n5559 & 2_n496;
assign 2_n2007 = ~(2_n2086 ^ 2_n7547);
assign 2_n6659 = ~(2_n7359 ^ 2_n8616);
assign 2_n11289 = 2_n4498 | 2_n5497;
assign 2_n10195 = ~(2_n2608 | 2_n4615);
assign 2_n1467 = ~2_n670;
assign 2_n12265 = ~(2_n11377 ^ 2_n4052);
assign 2_n9114 = 2_n3096 | 2_n6197;
assign 2_n12106 = ~(2_n887 ^ 2_n8942);
assign 2_n12785 = ~(2_n9065 ^ 2_n141);
assign 2_n11886 = ~(2_n4999 ^ 2_n4897);
assign 2_n2345 = ~(2_n3978 ^ 2_n3515);
assign 2_n11694 = 2_n7391 | 2_n1851;
assign 2_n1064 = 2_n118 & 2_n5957;
assign 2_n11474 = ~2_n7519;
assign 2_n6846 = 2_n2125 & 2_n9796;
assign 2_n12160 = ~(2_n5177 ^ 2_n4626);
assign 2_n9081 = 2_n11026 | 2_n9568;
assign 2_n9402 = ~2_n5697;
assign 2_n5261 = ~2_n9539;
assign 2_n4451 = 2_n1941 | 2_n11820;
assign 2_n12075 = ~(2_n747 ^ 2_n4069);
assign 2_n1443 = 2_n5436 & 2_n6471;
assign 2_n676 = ~2_n9677;
assign 2_n7897 = 2_n12406 & 2_n5121;
assign 2_n9592 = 2_n6030 & 2_n3866;
assign 2_n6858 = ~(2_n5377 ^ 2_n10765);
assign 2_n1968 = ~(2_n1557 | 2_n7030);
assign 2_n10924 = ~(2_n176 ^ 2_n6873);
assign 2_n10008 = ~(2_n1689 ^ 2_n9950);
assign 2_n1682 = 2_n7449 | 2_n6922;
assign 2_n4784 = 2_n9978 | 2_n2489;
assign 2_n2632 = 2_n3992 & 2_n8433;
assign 2_n5703 = 2_n8535 | 2_n2410;
assign 2_n9494 = ~(2_n4980 | 2_n8875);
assign 2_n9082 = 2_n7391 | 2_n7881;
assign 2_n4696 = 2_n7116 | 2_n12816;
assign 2_n7725 = ~2_n716;
assign 2_n11913 = 2_n1161 & 2_n134;
assign 2_n12192 = 2_n11434 | 2_n10153;
assign 2_n3185 = ~(2_n12347 | 2_n9480);
assign 2_n1397 = 2_n10545 & 2_n7159;
assign 2_n3564 = ~(2_n10959 ^ 2_n3879);
assign 2_n8596 = 2_n10142 | 2_n2076;
assign 2_n500 = 2_n10657 | 2_n11861;
assign 2_n9942 = 2_n7363 & 2_n10684;
assign 2_n3555 = 2_n9004 | 2_n3164;
assign 2_n8213 = ~(2_n10527 ^ 2_n4227);
assign 2_n2670 = 2_n994 | 2_n1162;
assign 2_n1528 = ~(2_n1139 ^ 2_n5098);
assign 2_n5190 = 2_n11969 & 2_n5585;
assign 2_n5526 = 2_n12391 & 2_n2558;
assign 2_n6193 = ~2_n1185;
assign 2_n12583 = 2_n5395 & 2_n1952;
assign 2_n10722 = ~(2_n8066 ^ 2_n9294);
assign 2_n8639 = ~(2_n4777 ^ 2_n7475);
assign 2_n10497 = ~(2_n6177 ^ 2_n10713);
assign 2_n141 = ~(2_n9073 ^ 2_n4641);
assign 2_n7553 = ~2_n270;
assign 2_n3900 = 2_n3562 | 2_n10796;
assign 2_n7127 = 2_n6601 & 2_n7223;
assign 2_n5167 = 2_n11736 & 2_n569;
assign 2_n7230 = 2_n12675 & 2_n11381;
assign 2_n10258 = 2_n11204 & 2_n243;
assign 2_n6464 = ~(2_n12351 ^ 2_n5804);
assign 2_n4032 = 2_n3967 | 2_n8057;
assign 2_n6740 = 2_n3746 | 2_n11820;
assign 2_n9773 = 2_n4966 & 2_n5161;
assign 2_n442 = ~(2_n690 | 2_n11084);
assign 2_n1693 = ~(2_n12004 ^ 2_n5033);
assign 2_n9719 = ~(2_n4012 ^ 2_n1971);
assign 2_n5673 = 2_n9199 & 2_n2302;
assign 2_n2623 = ~(2_n8863 ^ 2_n7766);
assign 2_n839 = 2_n6590 | 2_n11930;
assign 2_n11893 = ~2_n9547;
assign 2_n7577 = 2_n4787 & 2_n1889;
assign 2_n3734 = 2_n7810 | 2_n4538;
assign 2_n9652 = 2_n6718 | 2_n9144;
assign 2_n9954 = 2_n2995 & 2_n10800;
assign 2_n1130 = ~2_n1584;
assign 2_n6681 = 2_n5530 | 2_n5326;
assign 2_n7139 = 2_n12803 & 2_n11117;
assign 2_n12032 = ~(2_n11324 ^ 2_n12756);
assign 2_n639 = ~(2_n2381 ^ 2_n8506);
assign 2_n1461 = 2_n2456 | 2_n6071;
assign 2_n3623 = 2_n10435 & 2_n4895;
assign 2_n11001 = ~(2_n8123 ^ 2_n6774);
assign 2_n10036 = ~(2_n9152 ^ 2_n9509);
assign 2_n5449 = 2_n7906 | 2_n9794;
assign 2_n2236 = 2_n12930 | 2_n6947;
assign 2_n886 = ~(2_n2837 | 2_n5360);
assign 2_n8020 = 2_n4960 | 2_n4945;
assign 2_n5473 = 2_n9373 | 2_n12771;
assign 2_n1311 = ~2_n1594;
assign 2_n186 = 2_n12705 & 2_n3932;
assign 2_n10142 = ~2_n6687;
assign 2_n9203 = 2_n11923 | 2_n2020;
assign 2_n9070 = 2_n2056 | 2_n10008;
assign 2_n10747 = ~(2_n5294 ^ 2_n4748);
assign 2_n2654 = 2_n4579 | 2_n1167;
assign 2_n11602 = 2_n8216 | 2_n10480;
assign 2_n9159 = 2_n5160 | 2_n9283;
assign 2_n1496 = ~(2_n6993 ^ 2_n8633);
assign 2_n5652 = 2_n4628 | 2_n530;
assign 2_n1005 = ~(2_n11813 | 2_n8922);
assign 2_n64 = 2_n2842 & 2_n6424;
assign 2_n10675 = 2_n6032 | 2_n3801;
assign 2_n8405 = ~2_n6578;
assign 2_n11788 = ~(2_n11610 ^ 2_n2547);
assign 2_n4774 = 2_n4972 & 2_n2542;
assign 2_n11068 = 2_n5945 | 2_n2232;
assign 2_n8169 = 2_n2382 | 2_n948;
assign 2_n4396 = ~(2_n5092 | 2_n3074);
assign 2_n1714 = 2_n12610 | 2_n7794;
assign 2_n11266 = 2_n11923 | 2_n4875;
assign 2_n11608 = 2_n3127 | 2_n11827;
assign 2_n8210 = ~2_n8772;
assign 2_n9482 = 2_n12273 & 2_n9256;
assign 2_n6458 = 2_n5788 | 2_n7673;
assign 2_n7728 = ~(2_n2009 ^ 2_n12921);
assign 2_n5978 = 2_n4481 & 2_n10634;
assign 2_n4176 = ~2_n6751;
assign 2_n6028 = 2_n11941 | 2_n4793;
assign 2_n12190 = ~(2_n9490 | 2_n767);
assign 2_n1730 = ~(2_n5559 | 2_n496);
assign 2_n11371 = ~(2_n6067 | 2_n8182);
assign 2_n1151 = 2_n4275 & 2_n9813;
assign 2_n7449 = ~2_n7388;
assign 2_n3704 = ~(2_n6984 ^ 2_n2543);
assign 2_n1366 = ~(2_n4714 ^ 2_n1118);
assign 2_n5735 = ~2_n10425;
assign 2_n8668 = ~(2_n10743 ^ 2_n8721);
assign 2_n8135 = 2_n288 | 2_n11386;
assign 2_n10134 = 2_n3829 | 2_n10384;
assign 2_n12158 = ~(2_n1091 ^ 2_n10497);
assign 2_n7652 = ~(2_n4794 ^ 2_n7799);
assign 2_n3389 = 2_n4247 | 2_n554;
assign 2_n4228 = 2_n10196 | 2_n8643;
assign 2_n1547 = 2_n10824 | 2_n6501;
assign 2_n2262 = ~2_n10831;
assign 2_n2825 = ~(2_n5454 ^ 2_n9125);
assign 2_n1686 = 2_n1261 & 2_n2366;
assign 2_n12867 = 2_n7683 & 2_n12954;
assign 2_n10831 = 2_n2093 | 2_n6102;
assign 2_n3359 = 2_n9829 & 2_n5541;
assign 2_n4421 = ~2_n5207;
assign 2_n11610 = ~(2_n5784 ^ 2_n10591);
assign 2_n9902 = ~(2_n8484 ^ 2_n4363);
assign 2_n5983 = ~(2_n11624 ^ 2_n3484);
assign 2_n2045 = 2_n8428 | 2_n6197;
assign 2_n5276 = 2_n3627 & 2_n6038;
assign 2_n8357 = ~(2_n6135 ^ 2_n12459);
assign 2_n4122 = ~(2_n12931 | 2_n9495);
assign 2_n8649 = 2_n27 | 2_n1050;
assign 2_n8783 = ~(2_n6467 ^ 2_n11860);
assign 2_n3278 = 2_n11923 | 2_n4864;
assign 2_n7199 = ~(2_n4512 | 2_n11170);
assign 2_n10118 = 2_n5765 | 2_n9144;
assign 2_n2353 = ~(2_n2549 | 2_n1680);
assign 2_n2093 = ~(2_n7115 | 2_n310);
assign 2_n5045 = ~2_n7464;
assign 2_n8328 = ~(2_n5647 | 2_n10263);
assign 2_n2589 = ~2_n2278;
assign 2_n4046 = 2_n6072 | 2_n891;
assign 2_n12401 = 2_n3251 & 2_n1274;
assign 2_n3705 = ~(2_n2906 ^ 2_n6699);
assign 2_n1292 = 2_n12722 | 2_n1763;
assign 2_n12759 = 2_n3491 & 2_n8543;
assign 2_n12122 = 2_n2099 | 2_n9188;
assign 2_n10981 = ~(2_n5109 ^ 2_n12295);
assign 2_n2187 = 2_n8229 | 2_n1276;
assign 2_n416 = ~(2_n7504 ^ 2_n224);
assign 2_n12307 = ~2_n12664;
assign 2_n2949 = ~(2_n1760 ^ 2_n12766);
assign 2_n7022 = ~2_n4386;
assign 2_n8096 = 2_n11552 | 2_n8830;
assign 2_n2795 = 2_n9379 & 2_n1356;
assign 2_n2663 = 2_n7116 | 2_n8768;
assign 2_n9745 = ~(2_n2314 ^ 2_n268);
assign 2_n2765 = ~(2_n2644 ^ 2_n12810);
assign 2_n6843 = 2_n7283 | 2_n9589;
assign 2_n1239 = 2_n7243 | 2_n2460;
assign 2_n6803 = ~(2_n8118 ^ 2_n11933);
assign 2_n10530 = 2_n8583 | 2_n9144;
assign 2_n1494 = 2_n4347 & 2_n6375;
assign 2_n1602 = 2_n4369 & 2_n467;
assign 2_n8141 = ~(2_n4717 | 2_n12302);
assign 2_n2705 = 2_n11328 & 2_n6043;
assign 2_n11482 = ~(2_n7551 ^ 2_n9867);
assign 2_n5091 = ~(2_n8163 | 2_n3914);
assign 2_n12323 = ~(2_n11550 ^ 2_n5176);
assign 2_n6479 = ~(2_n1654 ^ 2_n8571);
assign 2_n2455 = 2_n6574 | 2_n8331;
assign 2_n7550 = 2_n10843 | 2_n11295;
assign 2_n2352 = ~(2_n11617 ^ 2_n8400);
assign 2_n8505 = ~2_n2500;
assign 2_n2119 = ~(2_n10456 ^ 2_n32);
assign 2_n3216 = ~2_n9437;
assign 2_n2113 = 2_n4059 | 2_n561;
assign 2_n307 = 2_n4492 | 2_n11901;
assign 2_n11355 = 2_n9905 & 2_n10792;
assign 2_n10096 = 2_n2687 & 2_n7153;
assign 2_n10752 = 2_n2159 & 2_n12822;
assign 2_n12184 = ~(2_n1637 | 2_n11325);
assign 2_n163 = ~(2_n10497 | 2_n1091);
assign 2_n1819 = ~(2_n7763 ^ 2_n185);
assign 2_n2988 = 2_n12727 | 2_n8005;
assign 2_n6836 = 2_n2217 | 2_n1476;
assign 2_n12416 = 2_n12853 | 2_n8109;
assign 2_n7622 = ~(2_n4137 ^ 2_n4640);
assign 2_n11950 = 2_n12699 & 2_n4113;
assign 2_n10182 = 2_n7116 | 2_n11122;
assign 2_n4842 = 2_n9136 | 2_n7642;
assign 2_n3749 = ~(2_n2674 ^ 2_n11847);
assign 2_n4558 = ~(2_n3769 ^ 2_n3070);
assign 2_n7215 = ~(2_n5887 ^ 2_n11904);
assign 2_n11812 = ~2_n255;
assign 2_n3757 = 2_n5765 | 2_n1047;
assign 2_n11320 = ~(2_n9000 ^ 2_n11598);
assign 2_n12746 = 2_n5355 | 2_n4400;
assign 2_n9672 = ~(2_n11646 ^ 2_n1203);
assign 2_n826 = ~2_n5645;
assign 2_n2185 = ~(2_n10639 | 2_n6479);
assign 2_n9950 = ~2_n4967;
assign 2_n42 = ~(2_n12508 ^ 2_n2994);
assign 2_n409 = ~(2_n715 ^ 2_n4000);
assign 2_n6489 = 2_n1985 & 2_n4186;
assign 2_n7796 = ~(2_n2307 ^ 2_n12902);
assign 2_n12480 = ~(2_n3541 ^ 2_n11067);
assign 2_n11720 = ~(2_n817 ^ 2_n9361);
assign 2_n6409 = 2_n6642 & 2_n1893;
assign 2_n7063 = ~2_n10556;
assign 2_n10319 = ~(2_n6580 ^ 2_n5304);
assign 2_n11105 = ~(2_n11280 ^ 2_n8825);
assign 2_n2679 = ~(2_n68 ^ 2_n1876);
assign 2_n8406 = ~(2_n11983 ^ 2_n1036);
assign 2_n4978 = ~(2_n4669 ^ 2_n9650);
assign 2_n2004 = ~(2_n3148 ^ 2_n6821);
assign 2_n7775 = ~(2_n5983 ^ 2_n9347);
assign 2_n260 = 2_n10208 | 2_n11932;
assign 2_n1400 = ~(2_n7686 ^ 2_n10079);
assign 2_n10621 = 2_n41 & 2_n1255;
assign 2_n10953 = 2_n9529 & 2_n7950;
assign 2_n8567 = ~(2_n2432 ^ 2_n213);
assign 2_n9812 = 2_n5108 & 2_n9198;
assign 2_n878 = 2_n756 | 2_n12428;
assign 2_n3433 = ~2_n4270;
assign 2_n12098 = 2_n6373 | 2_n4875;
assign 2_n12419 = 2_n6001 | 2_n1152;
assign 2_n584 = 2_n4994 | 2_n2980;
assign 2_n534 = ~(2_n6889 ^ 2_n6179);
assign 2_n8356 = 2_n3627 & 2_n11407;
assign 2_n4467 = ~(2_n7684 | 2_n12162);
assign 2_n7743 = ~(2_n2717 ^ 2_n5282);
assign 2_n8151 = ~(2_n8055 ^ 2_n8344);
assign 2_n727 = ~2_n7528;
assign 2_n724 = 2_n3275 | 2_n9293;
assign 2_n9475 = 2_n8753 & 2_n5752;
assign 2_n3448 = ~(2_n3068 ^ 2_n12058);
assign 2_n7346 = 2_n4716 & 2_n7;
assign 2_n1120 = ~(2_n633 ^ 2_n1221);
assign 2_n1220 = 2_n5960 & 2_n10664;
assign 2_n12316 = 2_n994 | 2_n9589;
assign 2_n5113 = ~(2_n9903 ^ 2_n7362);
assign 2_n5603 = ~(2_n6964 ^ 2_n2143);
assign 2_n11455 = 2_n5589 & 2_n11291;
assign 2_n906 = 2_n4453 | 2_n4706;
assign 2_n9658 = 2_n11535 & 2_n11767;
assign 2_n4061 = 2_n10750 | 2_n6071;
assign 2_n8378 = ~(2_n9863 ^ 2_n12860);
assign 2_n7033 = 2_n921 | 2_n8298;
assign 2_n6069 = 2_n2838 & 2_n6164;
assign 2_n1019 = 2_n9389 | 2_n11746;
assign 2_n3815 = 2_n10640 & 2_n5223;
assign 2_n7778 = 2_n6358 & 2_n217;
assign 2_n545 = 2_n333 | 2_n487;
assign 2_n8987 = 2_n8490 & 2_n5321;
assign 2_n7813 = 2_n8945 & 2_n1859;
assign 2_n3337 = 2_n8158 & 2_n5616;
assign 2_n11399 = ~(2_n6515 ^ 2_n11471);
assign 2_n4013 = 2_n2045 | 2_n11274;
assign 2_n3333 = 2_n0 & 2_n9322;
assign 2_n7378 = 2_n4911 | 2_n1455;
assign 2_n425 = ~(2_n75 ^ 2_n1823);
assign 2_n8933 = 2_n8363 & 2_n5806;
assign 2_n8407 = ~2_n2695;
assign 2_n8451 = 2_n12924 | 2_n1124;
assign 2_n4891 = 2_n10843 & 2_n11295;
assign 2_n11833 = ~(2_n408 ^ 2_n11082);
assign 2_n813 = 2_n7306 & 2_n10584;
assign 2_n10366 = ~(2_n2457 ^ 2_n2517);
assign 2_n2667 = 2_n2266 | 2_n11618;
assign 2_n5722 = ~(2_n11021 ^ 2_n9660);
assign 2_n6945 = 2_n8583 | 2_n8830;
assign 2_n2085 = 2_n12299 & 2_n8819;
assign 2_n3413 = ~(2_n9709 | 2_n2015);
assign 2_n10485 = 2_n11108 | 2_n11637;
assign 2_n779 = 2_n10642 | 2_n9973;
assign 2_n12774 = ~(2_n11137 | 2_n470);
assign 2_n10176 = 2_n8758 & 2_n12630;
assign 2_n523 = 2_n2367 | 2_n4474;
assign 2_n2252 = ~2_n8447;
assign 2_n3269 = ~(2_n12210 ^ 2_n12536);
assign 2_n9535 = ~(2_n1062 ^ 2_n12811);
assign 2_n11902 = 2_n5466 | 2_n4578;
assign 2_n5663 = 2_n1808 | 2_n2210;
assign 2_n11496 = ~(2_n4742 ^ 2_n8621);
assign 2_n6113 = ~(2_n9298 | 2_n10013);
assign 2_n9436 = ~(2_n6161 ^ 2_n12599);
assign 2_n938 = 2_n10354 | 2_n1502;
assign 2_n6696 = ~2_n9391;
assign 2_n4526 = ~(2_n9493 ^ 2_n10069);
assign 2_n428 = 2_n4121 | 2_n11975;
assign 2_n6093 = 2_n2013 | 2_n8542;
assign 2_n4749 = ~(2_n9079 ^ 2_n6695);
assign 2_n7024 = ~(2_n1242 ^ 2_n6378);
assign 2_n12728 = ~(2_n3225 ^ 2_n7099);
assign 2_n2814 = 2_n11358 | 2_n6201;
assign 2_n7169 = 2_n11416 | 2_n2535;
assign 2_n9803 = 2_n11832 & 2_n9681;
assign 2_n12148 = ~(2_n4703 ^ 2_n11570);
assign 2_n9925 = 2_n9802 | 2_n9220;
assign 2_n12850 = ~(2_n9368 ^ 2_n809);
assign 2_n2695 = 2_n12503 | 2_n2020;
assign 2_n10909 = ~(2_n7441 | 2_n3009);
assign 2_n8765 = ~(2_n11563 ^ 2_n5192);
assign 2_n8034 = ~(2_n7579 | 2_n10073);
assign 2_n3538 = ~2_n733;
assign 2_n3101 = ~(2_n5016 ^ 2_n12202);
assign 2_n3434 = ~2_n3443;
assign 2_n4231 = ~(2_n771 ^ 2_n1829);
assign 2_n12242 = 2_n10835 | 2_n9160;
assign 2_n3793 = 2_n3837 | 2_n9096;
assign 2_n9797 = 2_n10835 | 2_n10916;
assign 2_n4610 = ~2_n4784;
assign 2_n8264 = 2_n5847 | 2_n136;
assign 2_n6933 = ~(2_n645 | 2_n4043);
assign 2_n1184 = ~2_n6474;
assign 2_n6893 = 2_n10874 | 2_n1300;
assign 2_n2764 = ~(2_n11538 ^ 2_n8798);
assign 2_n12610 = ~(2_n12118 ^ 2_n3721);
assign 2_n2369 = ~(2_n522 ^ 2_n8401);
assign 2_n3050 = 2_n10835 | 2_n1047;
assign 2_n9670 = 2_n5384 & 2_n12652;
assign 2_n5592 = 2_n8115 | 2_n1106;
assign 2_n2351 = 2_n8467 | 2_n8231;
assign 2_n7266 = 2_n11271 | 2_n8239;
assign 2_n9060 = 2_n9119 & 2_n1182;
assign 2_n1542 = 2_n10326 & 2_n9618;
assign 2_n10619 = 2_n11719 | 2_n10066;
assign 2_n5902 = ~2_n6826;
assign 2_n9345 = 2_n9236 & 2_n1559;
assign 2_n1538 = ~(2_n11605 ^ 2_n3278);
assign 2_n9235 = ~2_n3460;
assign 2_n1976 = ~(2_n10746 | 2_n10577);
assign 2_n11124 = 2_n3381 & 2_n10811;
assign 2_n5218 = ~(2_n11548 | 2_n4523);
assign 2_n11467 = ~(2_n6907 ^ 2_n3610);
assign 2_n8434 = ~(2_n3840 ^ 2_n4151);
assign 2_n4333 = ~(2_n8792 ^ 2_n6372);
assign 2_n9794 = 2_n9878 | 2_n12535;
assign 2_n8962 = ~2_n8732;
assign 2_n2012 = ~2_n8790;
assign 2_n3522 = ~2_n1027;
assign 2_n1661 = ~(2_n2063 ^ 2_n7466);
assign 2_n1445 = 2_n8959 | 2_n6197;
assign 2_n10573 = 2_n12237 | 2_n3224;
assign 2_n5617 = ~(2_n12195 ^ 2_n4622);
assign 2_n10225 = 2_n10336 & 2_n11677;
assign 2_n11469 = ~(2_n1248 ^ 2_n8440);
assign 2_n11350 = ~2_n10914;
assign 2_n10641 = ~2_n9738;
assign 2_n6556 = ~(2_n3085 ^ 2_n2554);
assign 2_n947 = 2_n8152 | 2_n11942;
assign 2_n9432 = 2_n5355 | 2_n7703;
assign 2_n1168 = ~(2_n6413 ^ 2_n12778);
assign 2_n8107 = ~(2_n9358 ^ 2_n547);
assign 2_n8956 = ~(2_n7092 ^ 2_n4030);
assign 2_n1871 = ~2_n3978;
assign 2_n10673 = 2_n5384 | 2_n12652;
assign 2_n2221 = ~2_n1611;
assign 2_n837 = ~(2_n5483 ^ 2_n5072);
assign 2_n1043 = 2_n6577 | 2_n9741;
assign 2_n7768 = 2_n2097 | 2_n3792;
assign 2_n1406 = ~(2_n6889 | 2_n9422);
assign 2_n12290 = 2_n9368 & 2_n809;
assign 2_n12928 = ~(2_n11234 ^ 2_n2359);
assign 2_n4284 = ~(2_n2069 ^ 2_n10458);
assign 2_n5851 = ~2_n3865;
assign 2_n5772 = ~(2_n8287 ^ 2_n10188);
assign 2_n2600 = 2_n12119 | 2_n12446;
assign 2_n9689 = ~(2_n7070 | 2_n10571);
assign 2_n3765 = 2_n9933 & 2_n8729;
assign 2_n8705 = 2_n3771 & 2_n3302;
assign 2_n11299 = 2_n2497 | 2_n9001;
assign 2_n566 = 2_n6934 & 2_n1377;
assign 2_n6799 = ~(2_n4926 ^ 2_n2745);
assign 2_n1038 = ~(2_n7285 ^ 2_n6498);
assign 2_n11093 = 2_n3766 & 2_n11974;
assign 2_n1917 = 2_n849 | 2_n4575;
assign 2_n3814 = 2_n3581 & 2_n6230;
assign 2_n2441 = 2_n3236 & 2_n3067;
assign 2_n7696 = ~(2_n3517 ^ 2_n823);
assign 2_n3751 = ~(2_n1252 | 2_n9565);
assign 2_n8854 = 2_n196 & 2_n11477;
assign 2_n5829 = ~(2_n6794 | 2_n3545);
assign 2_n3652 = 2_n6550 | 2_n5792;
assign 2_n10418 = 2_n8071 | 2_n7595;
assign 2_n8137 = 2_n5850 | 2_n1347;
assign 2_n4264 = 2_n6977 | 2_n5012;
assign 2_n11031 = ~2_n11501;
assign 2_n3405 = 2_n1051 | 2_n12816;
assign 2_n11775 = ~2_n3602;
assign 2_n5594 = ~2_n6087;
assign 2_n1520 = ~(2_n11112 ^ 2_n5123);
assign 2_n12843 = ~2_n4921;
assign 2_n7279 = ~(2_n9194 ^ 2_n2480);
assign 2_n1911 = 2_n7735 & 2_n1324;
assign 2_n4801 = ~(2_n7817 | 2_n9118);
assign 2_n7096 = 2_n10742 & 2_n12001;
assign 2_n10101 = ~2_n1515;
assign 2_n3739 = 2_n6766 | 2_n395;
assign 2_n3214 = ~(2_n4583 ^ 2_n4276);
assign 2_n7326 = ~2_n12710;
assign 2_n3301 = ~(2_n7746 ^ 2_n4743);
assign 2_n1317 = 2_n2217 | 2_n9160;
assign 2_n270 = 2_n12531 | 2_n5565;
assign 2_n2395 = 2_n5915 | 2_n3224;
assign 2_n3166 = 2_n10142 | 2_n4400;
assign 2_n5192 = 2_n7449 | 2_n9521;
assign 2_n6287 = 2_n9570 & 2_n12050;
assign 2_n4849 = 2_n4059 | 2_n1455;
assign 2_n11369 = ~2_n12632;
assign 2_n6942 = ~(2_n3985 ^ 2_n5112);
assign 2_n4369 = 2_n10551 | 2_n7988;
assign 2_n8282 = 2_n6977 | 2_n8414;
assign 2_n8459 = 2_n9896 & 2_n9815;
assign 2_n3151 = ~(2_n11343 ^ 2_n6106);
assign 2_n10632 = 2_n9262 | 2_n4474;
assign 2_n6602 = ~(2_n10525 | 2_n9466);
assign 2_n8684 = ~2_n7143;
assign 2_n9783 = ~(2_n12142 ^ 2_n12061);
assign 2_n11232 = 2_n3746 | 2_n7395;
assign 2_n6985 = ~2_n4079;
assign 2_n10472 = 2_n4202 & 2_n9496;
assign 2_n11794 = 2_n3324 | 2_n1509;
assign 2_n1348 = ~(2_n9063 | 2_n9580);
assign 2_n1201 = ~(2_n3584 ^ 2_n4037);
assign 2_n5606 = 2_n11950 & 2_n5127;
assign 2_n3465 = 2_n4187 & 2_n3602;
assign 2_n2277 = ~(2_n221 | 2_n3529);
assign 2_n1448 = ~2_n10904;
assign 2_n12409 = ~(2_n2912 ^ 2_n4192);
assign 2_n9882 = 2_n11152 & 2_n10482;
assign 2_n469 = ~(2_n6220 ^ 2_n59);
assign 2_n12589 = ~(2_n10983 ^ 2_n91);
assign 2_n11505 = 2_n10108 | 2_n11827;
assign 2_n12407 = ~(2_n5424 | 2_n9337);
assign 2_n9433 = 2_n7221 | 2_n6453;
assign 2_n10312 = 2_n2593 | 2_n8497;
assign 2_n12268 = ~(2_n7386 ^ 2_n8651);
assign 2_n8606 = ~(2_n3077 ^ 2_n2627);
assign 2_n3272 = ~(2_n5354 ^ 2_n6014);
assign 2_n10562 = ~(2_n1785 ^ 2_n12143);
assign 2_n2387 = ~(2_n2637 ^ 2_n8950);
assign 2_n4771 = ~(2_n6090 ^ 2_n1698);
assign 2_n2982 = 2_n5089 | 2_n10823;
assign 2_n3589 = 2_n7905 | 2_n12431;
assign 2_n10384 = ~(2_n721 | 2_n9327);
assign 2_n12094 = ~(2_n7483 ^ 2_n5297);
assign 2_n10980 = ~(2_n4541 | 2_n7995);
assign 2_n10128 = 2_n3324 | 2_n4474;
assign 2_n3541 = 2_n10508 | 2_n10930;
assign 2_n10636 = 2_n10199 | 2_n7637;
assign 2_n6597 = ~(2_n9446 | 2_n9051);
assign 2_n11384 = 2_n1705 | 2_n12251;
assign 2_n11501 = 2_n12815 & 2_n10109;
assign 2_n6127 = ~(2_n10744 ^ 2_n5913);
assign 2_n9874 = ~(2_n9145 ^ 2_n12649);
assign 2_n4887 = ~(2_n9499 ^ 2_n11096);
assign 2_n4414 = 2_n12069 & 2_n1564;
assign 2_n4668 = 2_n3265 & 2_n1454;
assign 2_n323 = 2_n12879 & 2_n7792;
assign 2_n7512 = ~2_n2640;
assign 2_n9278 = ~(2_n2011 | 2_n4899);
assign 2_n10087 = 2_n6087 ^ 2_n3134;
assign 2_n5106 = ~(2_n6168 ^ 2_n4418);
assign 2_n10741 = 2_n5289 & 2_n6166;
assign 2_n12363 = ~2_n11842;
assign 2_n9112 = 2_n4013 & 2_n9800;
assign 2_n382 = ~(2_n8140 ^ 2_n10253);
assign 2_n11508 = 2_n6776 & 2_n6703;
assign 2_n3426 = 2_n3693 | 2_n12795;
assign 2_n9989 = ~(2_n4930 | 2_n12448);
assign 2_n5098 = ~2_n6683;
assign 2_n10704 = ~(2_n9278 | 2_n12352);
assign 2_n10681 = ~(2_n10815 ^ 2_n9254);
assign 2_n5217 = ~(2_n7244 ^ 2_n2890);
assign 2_n5541 = ~2_n11256;
assign 2_n7287 = 2_n11425 | 2_n6025;
assign 2_n11768 = ~(2_n5846 ^ 2_n12628);
assign 2_n9796 = 2_n12283 | 2_n8333;
assign 2_n691 = ~(2_n7496 ^ 2_n3436);
assign 2_n10843 = ~(2_n11533 ^ 2_n12068);
assign 2_n3367 = ~(2_n2488 ^ 2_n6203);
assign 2_n9806 = 2_n5809 | 2_n12080;
assign 2_n8191 = 2_n7283 | 2_n2076;
assign 2_n4803 = 2_n5231 & 2_n5217;
assign 2_n12449 = ~(2_n8313 ^ 2_n879);
assign 2_n4238 = 2_n10735 | 2_n4091;
assign 2_n3285 = ~(2_n3884 ^ 2_n734);
assign 2_n8084 = ~(2_n12203 ^ 2_n10593);
assign 2_n4034 = 2_n3274 & 2_n3755;
assign 2_n350 = ~(2_n1065 | 2_n4039);
assign 2_n8900 = 2_n7236 & 2_n5760;
assign 2_n8782 = 2_n7271 | 2_n11263;
assign 2_n2639 = ~(2_n10918 | 2_n12900);
assign 2_n1561 = 2_n5020 & 2_n3916;
assign 2_n5721 = ~(2_n12873 ^ 2_n10513);
assign 2_n6384 = 2_n8176 & 2_n2388;
assign 2_n8789 = 2_n5575 | 2_n11896;
assign 2_n7437 = 2_n4428 | 2_n8797;
assign 2_n1745 = 2_n1507 | 2_n9168;
assign 2_n134 = 2_n10521 | 2_n1828;
assign 2_n699 = 2_n8903 & 2_n5834;
assign 2_n10822 = 2_n3666 | 2_n7068;
assign 2_n12100 = ~(2_n10091 ^ 2_n3560);
assign 2_n12091 = ~(2_n6195 ^ 2_n7571);
assign 2_n1551 = ~(2_n5284 ^ 2_n12676);
assign 2_n12443 = 2_n994 | 2_n1079;
assign 2_n4052 = ~2_n10042;
assign 2_n2188 = 2_n9797 | 2_n2900;
assign 2_n8293 = ~2_n10741;
assign 2_n1361 = ~(2_n8027 ^ 2_n228);
assign 2_n5325 = ~(2_n1408 ^ 2_n11875);
assign 2_n7395 = ~2_n10278;
assign 2_n10075 = 2_n11462 | 2_n11148;
assign 2_n976 = 2_n2651 | 2_n4394;
assign 2_n9636 = ~2_n10080;
assign 2_n3536 = ~(2_n11568 ^ 2_n8846);
assign 2_n3729 = 2_n3746 | 2_n10919;
assign 2_n4453 = ~(2_n6485 | 2_n1187);
assign 2_n368 = ~(2_n1571 ^ 2_n9891);
assign 2_n10633 = 2_n4522 | 2_n4656;
assign 2_n10774 = 2_n5204 | 2_n283;
assign 2_n7705 = ~2_n5432;
assign 2_n7653 = ~(2_n5795 ^ 2_n6118);
assign 2_n7846 = 2_n7283 | 2_n1738;
assign 2_n5846 = ~(2_n10393 ^ 2_n2540);
assign 2_n5932 = ~(2_n1989 | 2_n3600);
assign 2_n10024 = ~(2_n10457 ^ 2_n7820);
assign 2_n893 = 2_n5026 & 2_n9139;
assign 2_n4466 = 2_n8941 | 2_n1418;
assign 2_n7776 = 2_n12658 & 2_n6327;
assign 2_n1931 = ~2_n7312;
assign 2_n4811 = ~2_n10517;
assign 2_n3546 = ~(2_n11267 ^ 2_n4751);
assign 2_n4952 = ~2_n6203;
assign 2_n11358 = 2_n7168 | 2_n3047;
assign 2_n10742 = 2_n9920 & 2_n4921;
assign 2_n2145 = 2_n991 & 2_n354;
assign 2_n5376 = 2_n1215 & 2_n5055;
assign 2_n8744 = ~(2_n7146 ^ 2_n9552);
assign 2_n11377 = ~2_n2824;
assign 2_n4841 = ~2_n8773;
assign 2_n9471 = ~(2_n2739 | 2_n1033);
assign 2_n5651 = ~(2_n6857 ^ 2_n4544);
assign 2_n3017 = 2_n11892 & 2_n11791;
assign 2_n9534 = ~2_n11468;
assign 2_n11200 = 2_n10332 | 2_n12934;
assign 2_n6539 = 2_n3746 | 2_n11122;
assign 2_n11394 = 2_n5493 | 2_n5019;
assign 2_n2849 = ~2_n4;
assign 2_n7674 = 2_n9075 | 2_n4840;
assign 2_n512 = ~(2_n4233 ^ 2_n11553);
assign 2_n7820 = 2_n7453 & 2_n2059;
assign 2_n7040 = ~(2_n3651 | 2_n3183);
assign 2_n8535 = ~(2_n4655 ^ 2_n4825);
assign 2_n8528 = 2_n2427 & 2_n1157;
assign 2_n7636 = ~(2_n1050 ^ 2_n2544);
assign 2_n10907 = ~(2_n10297 ^ 2_n2983);
assign 2_n3618 = 2_n12474 | 2_n881;
assign 2_n5317 = ~(2_n7844 ^ 2_n12378);
assign 2_n6499 = ~(2_n5501 ^ 2_n4792);
assign 2_n6588 = ~(2_n5848 ^ 2_n3913);
assign 2_n4864 = ~2_n1510;
assign 2_n454 = ~(2_n10904 ^ 2_n5789);
assign 2_n8255 = 2_n817 | 2_n9817;
assign 2_n6110 = ~(2_n12867 ^ 2_n3443);
assign 2_n4128 = ~(2_n8189 ^ 2_n5797);
assign 2_n1750 = ~(2_n11564 ^ 2_n5015);
assign 2_n2388 = ~(2_n5009 ^ 2_n821);
assign 2_n4105 = 2_n3992 & 2_n8028;
assign 2_n8172 = ~(2_n2272 ^ 2_n10258);
assign 2_n6332 = ~(2_n2625 | 2_n4874);
assign 2_n5522 = 2_n11887 | 2_n9188;
assign 2_n5625 = 2_n4780 | 2_n10436;
assign 2_n2227 = 2_n12680 & 2_n3783;
assign 2_n3758 = ~(2_n775 ^ 2_n11071);
assign 2_n516 = ~(2_n11417 ^ 2_n1314);
assign 2_n195 = ~(2_n9999 ^ 2_n7478);
assign 2_n4998 = ~(2_n5942 ^ 2_n11064);
assign 2_n6444 = 2_n3964 & 2_n1334;
assign 2_n80 = 2_n6801 & 2_n6011;
assign 2_n11212 = 2_n4628 | 2_n5781;
assign 2_n3944 = 2_n1699 | 2_n1932;
assign 2_n9192 = 2_n213 | 2_n2432;
assign 2_n8540 = 2_n11422 & 2_n10028;
assign 2_n3019 = ~(2_n10441 ^ 2_n12904);
assign 2_n10424 = 2_n2901 & 2_n2938;
assign 2_n4689 = ~(2_n595 ^ 2_n10785);
assign 2_n2590 = 2_n12723 & 2_n1130;
assign 2_n4678 = ~(2_n669 ^ 2_n10559);
assign 2_n5457 = 2_n7284 & 2_n10144;
assign 2_n7803 = ~2_n12162;
assign 2_n11708 = ~(2_n3592 ^ 2_n12383);
assign 2_n1001 = ~(2_n2979 ^ 2_n9476);
assign 2_n8296 = ~(2_n7608 ^ 2_n10632);
assign 2_n6633 = ~(2_n3600 ^ 2_n8107);
assign 2_n10263 = ~(2_n610 | 2_n469);
assign 2_n6176 = ~(2_n6098 ^ 2_n1845);
assign 2_n5840 = ~2_n6824;
assign 2_n7358 = ~2_n10947;
assign 2_n9595 = ~(2_n4886 ^ 2_n5135);
assign 2_n7150 = ~(2_n12875 | 2_n6875);
assign 2_n8060 = ~(2_n11036 ^ 2_n5252);
assign 2_n12612 = ~(2_n9244 | 2_n4025);
assign 2_n11850 = 2_n6738 | 2_n11179;
assign 2_n2738 = 2_n11259 & 2_n6119;
assign 2_n5561 = 2_n4184 & 2_n3169;
assign 2_n5704 = ~2_n5236;
assign 2_n11412 = ~(2_n6945 ^ 2_n7023);
assign 2_n5016 = 2_n8026 | 2_n10903;
assign 2_n10730 = 2_n7839 | 2_n2815;
assign 2_n4524 = ~(2_n1366 ^ 2_n8351);
assign 2_n3303 = 2_n7161 | 2_n8765;
assign 2_n10888 = ~(2_n901 | 2_n11252);
assign 2_n4459 = 2_n11593 | 2_n4584;
assign 2_n2659 = 2_n5915 | 2_n826;
assign 2_n9889 = 2_n2832 | 2_n6389;
assign 2_n12810 = ~(2_n4413 ^ 2_n10803);
assign 2_n10254 = ~(2_n9649 ^ 2_n12726);
assign 2_n8804 = ~(2_n2611 ^ 2_n286);
assign 2_n5956 = ~(2_n3523 ^ 2_n9682);
assign 2_n9228 = 2_n1051 | 2_n2815;
assign 2_n9858 = 2_n4828 & 2_n2498;
assign 2_n3064 = 2_n12299 & 2_n2522;
assign 2_n12737 = 2_n7668 & 2_n9130;
assign 2_n1342 = 2_n5765 | 2_n8285;
assign 2_n367 = 2_n9795 | 2_n9719;
assign 2_n3320 = ~(2_n8092 ^ 2_n8358);
assign 2_n2409 = 2_n6590 & 2_n11930;
assign 2_n9914 = ~(2_n12294 | 2_n6665);
assign 2_n586 = 2_n10838 | 2_n3060;
assign 2_n8757 = 2_n10157 | 2_n3606;
assign 2_n5970 = ~2_n5192;
assign 2_n10658 = ~(2_n8790 ^ 2_n4089);
assign 2_n1857 = ~2_n1949;
assign 2_n8108 = 2_n6931 | 2_n4506;
assign 2_n9638 = 2_n11028 | 2_n8;
assign 2_n7632 = ~(2_n2874 ^ 2_n9587);
assign 2_n5774 = 2_n222 & 2_n9742;
assign 2_n1286 = ~2_n12159;
assign 2_n10462 = 2_n6373 | 2_n609;
assign 2_n7428 = ~(2_n7794 ^ 2_n11888);
assign 2_n2916 = 2_n8011 & 2_n4866;
assign 2_n6285 = ~(2_n2629 ^ 2_n8062);
assign 2_n2417 = ~2_n7043;
assign 2_n4848 = ~2_n11878;
assign 2_n1672 = ~(2_n8712 ^ 2_n10344);
assign 2_n809 = 2_n5765 | 2_n9160;
assign 2_n92 = 2_n7407 | 2_n10662;
assign 2_n12034 = ~2_n6520;
assign 2_n6760 = ~(2_n10580 ^ 2_n9095);
assign 2_n11182 = 2_n8428 | 2_n7425;
assign 2_n9972 = 2_n8428 | 2_n8414;
assign 2_n12682 = ~(2_n11694 ^ 2_n4377);
assign 2_n5165 = ~(2_n12772 ^ 2_n9264);
assign 2_n6974 = 2_n7826 & 2_n12034;
assign 2_n10306 = 2_n12797 | 2_n7876;
assign 2_n268 = ~(2_n3006 ^ 2_n2446);
assign 2_n2620 = ~2_n5327;
assign 2_n5346 = 2_n8844 & 2_n302;
assign 2_n3457 = 2_n7449 | 2_n4654;
assign 2_n1360 = 2_n9331 | 2_n1592;
assign 2_n5715 = ~2_n7024;
assign 2_n4416 = ~(2_n11995 ^ 2_n8168);
assign 2_n9497 = 2_n8738 | 2_n12771;
assign 2_n12849 = 2_n12260 | 2_n1501;
assign 2_n5214 = 2_n4059 | 2_n7881;
assign 2_n9545 = ~(2_n9749 ^ 2_n7513);
assign 2_n6817 = 2_n4498 | 2_n1915;
assign 2_n2945 = 2_n12237 | 2_n8109;
assign 2_n9619 = 2_n12731 & 2_n2110;
assign 2_n8610 = 2_n4815 | 2_n5729;
assign 2_n1281 = ~(2_n12736 ^ 2_n2764);
assign 2_n3885 = 2_n1051 | 2_n10903;
assign 2_n4730 = ~(2_n3704 ^ 2_n9396);
assign 2_n5513 = ~(2_n11259 ^ 2_n6119);
assign 2_n2092 = ~(2_n4469 ^ 2_n1428);
assign 2_n8119 = 2_n5809 | 2_n5326;
assign 2_n5026 = ~(2_n11750 ^ 2_n10935);
assign 2_n2909 = ~(2_n12911 ^ 2_n2198);
assign 2_n11734 = 2_n7082 & 2_n10579;
assign 2_n5215 = 2_n1675 | 2_n344;
assign 2_n6684 = 2_n3241 | 2_n6236;
assign 2_n9234 = ~(2_n5542 ^ 2_n11232);
assign 2_n3 = ~(2_n1451 ^ 2_n9676);
assign 2_n6668 = ~(2_n7035 ^ 2_n11168);
assign 2_n7975 = ~(2_n12490 ^ 2_n6916);
assign 2_n9573 = 2_n11172 | 2_n6019;
assign 2_n10643 = 2_n3746 | 2_n6169;
assign 2_n7623 = ~(2_n7526 ^ 2_n4988);
assign 2_n6166 = 2_n7001 | 2_n6401;
assign 2_n3295 = 2_n10565 | 2_n10570;
assign 2_n10926 = 2_n4059 | 2_n1851;
assign 2_n138 = 2_n6589 & 2_n4049;
assign 2_n6601 = 2_n9108 | 2_n3983;
assign 2_n2882 = ~(2_n5931 ^ 2_n4617);
assign 2_n8319 = 2_n7832 & 2_n11869;
assign 2_n4897 = 2_n4201 & 2_n11762;
assign 2_n4731 = 2_n113 | 2_n10259;
assign 2_n9602 = ~(2_n6368 ^ 2_n12416);
assign 2_n1270 = 2_n2367 | 2_n2020;
assign 2_n7282 = 2_n5064 | 2_n8974;
assign 2_n9448 = ~2_n7779;
assign 2_n216 = ~(2_n8035 ^ 2_n6322);
assign 2_n5068 = ~2_n12319;
assign 2_n4170 = ~(2_n9794 ^ 2_n4954);
assign 2_n10017 = 2_n4531 & 2_n4885;
assign 2_n1394 = ~2_n6904;
assign 2_n3738 = ~(2_n459 ^ 2_n8609);
assign 2_n3327 = 2_n8555 & 2_n11568;
assign 2_n11771 = ~(2_n4366 ^ 2_n10752);
assign 2_n7677 = ~(2_n10160 ^ 2_n12201);
assign 2_n5913 = 2_n2289 & 2_n12192;
assign 2_n5697 = 2_n9472 & 2_n9462;
assign 2_n6307 = ~2_n1706;
assign 2_n761 = ~(2_n6244 ^ 2_n4042);
assign 2_n1245 = ~(2_n11246 ^ 2_n7814);
assign 2_n9154 = ~(2_n808 ^ 2_n5849);
assign 2_n6011 = 2_n8026 | 2_n10919;
assign 2_n12241 = 2_n8759 & 2_n3719;
assign 2_n11428 = ~2_n11882;
assign 2_n11465 = 2_n3455 & 2_n5392;
assign 2_n6781 = 2_n7626 & 2_n7913;
assign 2_n12893 = ~(2_n745 ^ 2_n10583);
assign 2_n2215 = 2_n2099 | 2_n12686;
assign 2_n9944 = ~(2_n4860 ^ 2_n1497);
assign 2_n4489 = ~(2_n5022 ^ 2_n2864);
assign 2_n7772 = ~(2_n4790 ^ 2_n3029);
assign 2_n5548 = ~(2_n7710 | 2_n3531);
assign 2_n4606 = ~(2_n7874 ^ 2_n4992);
assign 2_n4478 = 2_n2269 | 2_n6987;
assign 2_n5318 = 2_n3337 & 2_n10736;
assign 2_n181 = ~(2_n808 | 2_n9934);
assign 2_n1623 = 2_n2003 | 2_n12762;
assign 2_n6866 = 2_n7891 & 2_n7610;
assign 2_n3984 = 2_n10142 | 2_n10419;
assign 2_n2348 = 2_n11694 & 2_n4377;
assign 2_n5740 = 2_n3570 & 2_n9972;
assign 2_n5194 = 2_n3219 & 2_n1956;
assign 2_n3743 = ~2_n7236;
assign 2_n10365 = 2_n8187 | 2_n1851;
assign 2_n5383 = ~2_n6367;
assign 2_n11512 = ~(2_n12006 ^ 2_n5953);
assign 2_n3971 = ~(2_n2791 ^ 2_n278);
assign 2_n10968 = ~(2_n7154 ^ 2_n7994);
assign 2_n3622 = ~2_n7684;
assign 2_n4194 = ~(2_n4263 ^ 2_n8131);
assign 2_n9667 = 2_n499 | 2_n819;
assign 2_n12205 = 2_n1417 | 2_n12331;
assign 2_n7136 = ~2_n10965;
assign 2_n7032 = 2_n4778 | 2_n8740;
assign 2_n7853 = 2_n5945 | 2_n5012;
assign 2_n10811 = 2_n994 | 2_n6389;
assign 2_n1358 = 2_n7391 | 2_n8524;
assign 2_n12827 = ~(2_n7958 ^ 2_n9537);
assign 2_n10528 = 2_n4189 & 2_n7456;
assign 2_n4394 = ~(2_n7511 | 2_n12711);
assign 2_n6794 = 2_n6425 & 2_n10409;
assign 2_n6233 = ~(2_n103 ^ 2_n1273);
assign 2_n5302 = ~(2_n706 ^ 2_n12314);
assign 2_n12441 = ~2_n7546;
assign 2_n2973 = 2_n11742 | 2_n11342;
assign 2_n2147 = 2_n11680 & 2_n5625;
assign 2_n4098 = 2_n8687 | 2_n795;
assign 2_n5654 = 2_n2127 | 2_n3333;
assign 2_n7411 = ~(2_n10999 ^ 2_n1976);
assign 2_n9712 = ~(2_n7925 ^ 2_n5545);
assign 2_n4403 = 2_n6583 | 2_n10700;
assign 2_n2914 = ~(2_n12053 ^ 2_n4464);
assign 2_n12809 = ~2_n290;
assign 2_n10317 = ~(2_n12189 ^ 2_n4476);
assign 2_n12837 = 2_n1044 | 2_n6668;
assign 2_n3832 = 2_n7640 | 2_n1489;
assign 2_n1652 = ~(2_n7484 ^ 2_n10495);
assign 2_n6361 = 2_n3171 & 2_n8421;
assign 2_n6223 = ~(2_n8913 ^ 2_n4605);
assign 2_n10964 = 2_n10692 & 2_n1210;
assign 2_n10714 = 2_n6044 & 2_n12521;
assign 2_n1958 = ~(2_n10012 ^ 2_n5837);
assign 2_n12213 = 2_n9878 | 2_n12735;
assign 2_n5696 = 2_n6287 | 2_n10666;
assign 2_n9040 = ~(2_n7217 | 2_n11996);
assign 2_n5329 = 2_n1675 & 2_n344;
assign 2_n8617 = 2_n3743 | 2_n9280;
assign 2_n3014 = 2_n3115 | 2_n8324;
assign 2_n12216 = ~(2_n7166 ^ 2_n7878);
assign 2_n9525 = ~2_n2346;
assign 2_n1732 = ~(2_n7024 ^ 2_n1942);
assign 2_n3436 = ~(2_n703 ^ 2_n9491);
assign 2_n11554 = 2_n11272 & 2_n9192;
assign 2_n10961 = ~2_n6010;
assign 2_n4043 = ~(2_n4475 | 2_n7910);
assign 2_n6052 = ~(2_n8122 ^ 2_n1466);
assign 2_n3304 = 2_n12461 | 2_n8212;
assign 2_n11748 = ~2_n3831;
assign 2_n12844 = 2_n6901 & 2_n12638;
assign 2_n9446 = ~(2_n7693 | 2_n3330);
assign 2_n2575 = 2_n4001 | 2_n592;
assign 2_n6225 = ~(2_n7969 | 2_n3357);
assign 2_n6143 = 2_n11799 & 2_n8502;
assign 2_n2336 = 2_n7236 & 2_n10898;
assign 2_n12274 = ~2_n7823;
assign 2_n7627 = ~(2_n10837 ^ 2_n10968);
assign 2_n6589 = ~2_n11554;
assign 2_n6954 = 2_n9875 & 2_n7674;
assign 2_n12611 = 2_n4104 & 2_n8504;
assign 2_n411 = 2_n5925 | 2_n4882;
assign 2_n11543 = 2_n2357 | 2_n12434;
assign 2_n7466 = 2_n10622 | 2_n4876;
assign 2_n4986 = 2_n8187 | 2_n10066;
assign 2_n7794 = ~(2_n10140 ^ 2_n11763);
assign 2_n2276 = ~(2_n4358 ^ 2_n10715);
assign 2_n224 = 2_n6977 | 2_n2232;
assign 2_n12392 = ~(2_n7929 | 2_n732);
assign 2_n11631 = ~2_n3006;
assign 2_n3911 = ~2_n1798;
assign 2_n1852 = 2_n686 | 2_n1413;
assign 2_n11364 = 2_n9319 | 2_n5751;
assign 2_n4186 = 2_n1057 | 2_n2441;
assign 2_n5550 = 2_n9584 | 2_n795;
assign 2_n7753 = ~(2_n9976 ^ 2_n11224);
assign 2_n10985 = ~(2_n9701 | 2_n2799);
assign 2_n4055 = ~2_n7171;
assign 2_n3111 = ~(2_n1515 ^ 2_n6366);
assign 2_n8653 = 2_n6461 & 2_n3148;
assign 2_n3774 = 2_n144 & 2_n7137;
assign 2_n9368 = 2_n2217 | 2_n9144;
assign 2_n9532 = ~2_n492;
assign 2_n12660 = 2_n5918 | 2_n11409;
assign 2_n3688 = 2_n2069 | 2_n10458;
assign 2_n10653 = ~2_n4727;
assign 2_n8373 = 2_n9218 | 2_n10559;
assign 2_n12545 = 2_n8583 | 2_n7506;
assign 2_n2631 = 2_n8794 | 2_n2257;
assign 2_n5748 = 2_n12935 & 2_n9808;
assign 2_n4714 = ~(2_n11179 ^ 2_n10232);
assign 2_n2071 = 2_n12361 | 2_n11820;
assign 2_n10568 = 2_n8127 | 2_n7881;
assign 2_n10049 = 2_n7504 | 2_n224;
assign 2_n6904 = ~(2_n10537 ^ 2_n9412);
assign 2_n8906 = 2_n7967 & 2_n7261;
assign 2_n12755 = ~(2_n11029 | 2_n11685);
assign 2_n12064 = ~(2_n9829 ^ 2_n11256);
assign 2_n8857 = ~(2_n7980 ^ 2_n6183);
assign 2_n10465 = ~2_n7209;
assign 2_n9054 = 2_n10270 & 2_n6999;
assign 2_n6283 = 2_n2217 | 2_n12120;
assign 2_n1227 = ~(2_n10555 ^ 2_n2162);
assign 2_n11190 = ~(2_n3375 ^ 2_n1986);
assign 2_n4243 = 2_n12071 | 2_n9046;
assign 2_n7377 = 2_n11047 & 2_n7479;
assign 2_n4363 = ~(2_n6985 ^ 2_n11077);
assign 2_n10860 = 2_n9878 | 2_n12686;
assign 2_n9862 = 2_n6767 & 2_n6250;
assign 2_n10646 = 2_n8354 | 2_n12535;
assign 2_n11589 = 2_n8583 | 2_n12120;
assign 2_n11847 = ~(2_n590 | 2_n9762);
assign 2_n6144 = ~2_n11414;
assign 2_n9450 = 2_n8583 | 2_n4642;
assign 2_n4299 = 2_n5690 | 2_n1607;
assign 2_n281 = 2_n8374 | 2_n7235;
assign 2_n3379 = 2_n11154 | 2_n9405;
assign 2_n484 = 2_n7587 & 2_n2343;
assign 2_n1926 = 2_n9997 | 2_n12576;
assign 2_n7971 = 2_n9176 & 2_n12409;
assign 2_n4534 = ~2_n7664;
assign 2_n7243 = 2_n3743 | 2_n12120;
assign 2_n6538 = 2_n12147 | 2_n85;
assign 2_n12169 = ~(2_n4676 ^ 2_n8590);
assign 2_n9312 = ~2_n12404;
assign 2_n9177 = ~(2_n6564 ^ 2_n2896);
assign 2_n11131 = 2_n11674 & 2_n2726;
assign 2_n4939 = 2_n4674 | 2_n6513;
assign 2_n1059 = ~(2_n8899 ^ 2_n8565);
assign 2_n1165 = ~(2_n4461 | 2_n10766);
assign 2_n9921 = 2_n1423 & 2_n5471;
assign 2_n10533 = 2_n5423 & 2_n1528;
assign 2_n4902 = ~(2_n9205 | 2_n8089);
assign 2_n1670 = 2_n7661 & 2_n8724;
assign 2_n12017 = ~(2_n1874 | 2_n8233);
assign 2_n6642 = 2_n4782 | 2_n4554;
assign 2_n2621 = 2_n2448 & 2_n3799;
assign 2_n3797 = 2_n8025 & 2_n3280;
assign 2_n3267 = ~2_n6548;
assign 2_n5883 = 2_n807 | 2_n11775;
assign 2_n4770 = 2_n896 | 2_n10155;
assign 2_n4659 = 2_n12404 & 2_n6493;
assign 2_n5177 = ~(2_n2752 ^ 2_n9236);
assign 2_n9949 = 2_n3569 | 2_n2707;
assign 2_n5850 = 2_n5915 | 2_n8655;
assign 2_n11002 = 2_n2406 & 2_n8073;
assign 2_n2644 = ~(2_n5147 ^ 2_n8691);
assign 2_n4991 = ~(2_n789 ^ 2_n1056);
assign 2_n9937 = 2_n8127 | 2_n7341;
assign 2_n9688 = 2_n9373 | 2_n4875;
assign 2_n5359 = ~2_n10608;
assign 2_n8266 = ~(2_n9683 ^ 2_n6559);
assign 2_n12176 = ~(2_n2192 | 2_n11761);
assign 2_n180 = 2_n7209 | 2_n6807;
assign 2_n6951 = ~2_n2385;
assign 2_n10579 = ~(2_n10416 ^ 2_n4569);
assign 2_n11303 = ~(2_n9196 ^ 2_n4996);
assign 2_n1866 = ~(2_n12473 ^ 2_n10784);
assign 2_n12644 = ~(2_n8526 ^ 2_n12250);
assign 2_n12327 = 2_n9370 | 2_n1079;
assign 2_n7808 = ~(2_n1121 | 2_n11510);
assign 2_n3708 = ~(2_n4045 | 2_n1635);
assign 2_n12791 = ~(2_n5959 ^ 2_n10748);
assign 2_n3595 = ~(2_n7939 ^ 2_n11065);
assign 2_n12369 = 2_n962 | 2_n12771;
assign 2_n3706 = 2_n3743 | 2_n5914;
assign 2_n2300 = 2_n9148 | 2_n4417;
assign 2_n9138 = ~2_n1338;
assign 2_n2154 = ~(2_n11834 | 2_n12355);
assign 2_n370 = 2_n12119 | 2_n2259;
assign 2_n5116 = ~(2_n11233 | 2_n5078);
assign 2_n8058 = ~(2_n11928 ^ 2_n11308);
assign 2_n19 = 2_n8990 | 2_n1720;
assign 2_n4274 = ~(2_n6944 | 2_n8783);
assign 2_n4124 = 2_n2217 | 2_n6138;
assign 2_n6623 = ~(2_n8139 ^ 2_n1473);
assign 2_n5060 = 2_n11927 | 2_n8157;
assign 2_n5429 = 2_n9308 | 2_n9562;
assign 2_n129 = 2_n636 | 2_n10422;
assign 2_n2870 = 2_n2541 | 2_n10427;
assign 2_n11356 = 2_n191 | 2_n8735;
assign 2_n1331 = ~(2_n9854 ^ 2_n10430);
assign 2_n11959 = 2_n7283 | 2_n5851;
assign 2_n7787 = ~(2_n4304 ^ 2_n3074);
assign 2_n8292 = ~(2_n11372 ^ 2_n6918);
assign 2_n5379 = 2_n3659 & 2_n4993;
assign 2_n6690 = ~(2_n6579 ^ 2_n9997);
assign 2_n8011 = 2_n10157 | 2_n9144;
assign 2_n6334 = ~(2_n2600 ^ 2_n12332);
assign 2_n9421 = 2_n6174 | 2_n157;
assign 2_n4693 = 2_n3625 | 2_n9031;
assign 2_n3237 = ~(2_n6636 ^ 2_n6991);
assign 2_n6735 = ~(2_n10779 ^ 2_n1902);
assign 2_n7110 = ~(2_n9924 | 2_n2185);
assign 2_n3899 = 2_n11874 & 2_n6793;
assign 2_n7902 = 2_n3078 | 2_n6895;
assign 2_n7080 = ~(2_n3171 ^ 2_n2831);
assign 2_n10638 = ~(2_n10362 ^ 2_n1251);
assign 2_n6092 = 2_n8946 & 2_n1593;
assign 2_n9844 = ~2_n3546;
assign 2_n10977 = ~(2_n2064 ^ 2_n2267);
assign 2_n3082 = 2_n1574 & 2_n7706;
assign 2_n1487 = ~(2_n6519 ^ 2_n5549);
assign 2_n3357 = ~(2_n9657 | 2_n1807);
assign 2_n6881 = 2_n752 | 2_n6197;
assign 2_n212 = ~(2_n1759 | 2_n11817);
assign 2_n892 = ~2_n11166;
assign 2_n6483 = ~(2_n4010 ^ 2_n6300);
assign 2_n8920 = 2_n3127 | 2_n1079;
assign 2_n4630 = 2_n807 | 2_n7876;
assign 2_n4615 = 2_n7449 | 2_n4864;
assign 2_n7893 = 2_n2832 | 2_n3911;
assign 2_n7030 = 2_n5027 & 2_n10477;
assign 2_n10083 = ~(2_n11613 ^ 2_n5928);
assign 2_n4044 = ~(2_n12844 | 2_n9183);
assign 2_n355 = ~(2_n4492 ^ 2_n6521);
assign 2_n5159 = 2_n8631 | 2_n1453;
assign 2_n7452 = ~(2_n12956 ^ 2_n11030);
assign 2_n11660 = ~(2_n11959 ^ 2_n8659);
assign 2_n11114 = ~(2_n5216 ^ 2_n8306);
assign 2_n2972 = ~(2_n9141 | 2_n5149);
assign 2_n11633 = 2_n6247 & 2_n6973;
assign 2_n7719 = ~(2_n8897 ^ 2_n9213);
assign 2_n5943 = 2_n7037 & 2_n3232;
assign 2_n599 = 2_n7057 | 2_n3489;
assign 2_n2703 = ~(2_n7267 | 2_n8470);
assign 2_n8864 = 2_n2047 & 2_n12130;
assign 2_n244 = 2_n9754 | 2_n4491;
assign 2_n8352 = ~(2_n330 | 2_n2628);
assign 2_n10435 = 2_n191 | 2_n1915;
assign 2_n8893 = ~(2_n7133 ^ 2_n9918);
assign 2_n41 = 2_n1937 | 2_n995;
assign 2_n7681 = 2_n9240 & 2_n11264;
assign 2_n9752 = 2_n962 | 2_n4875;
assign 2_n11136 = ~(2_n939 ^ 2_n12824);
assign 2_n5334 = ~2_n9739;
assign 2_n6168 = 2_n2872 | 2_n6169;
assign 2_n8419 = ~(2_n3619 | 2_n7592);
assign 2_n1302 = 2_n10668 | 2_n2397;
assign 2_n6281 = ~(2_n10352 | 2_n8815);
assign 2_n5168 = 2_n8120 & 2_n4248;
assign 2_n9297 = 2_n9807 & 2_n6295;
assign 2_n466 = ~2_n11800;
assign 2_n7391 = ~2_n4312;
assign 2_n2784 = 2_n11311 & 2_n8819;
assign 2_n6715 = ~(2_n2626 ^ 2_n4041);
assign 2_n6297 = 2_n301 & 2_n3154;
assign 2_n2785 = ~(2_n12759 | 2_n7915);
assign 2_n2656 = ~(2_n11784 | 2_n9281);
assign 2_n3415 = ~2_n773;
assign 2_n6823 = 2_n1978 & 2_n5237;
assign 2_n6568 = ~(2_n4859 ^ 2_n8618);
assign 2_n687 = 2_n8793 | 2_n7736;
assign 2_n6396 = ~2_n5174;
assign 2_n5229 = ~(2_n2337 ^ 2_n9930);
assign 2_n8464 = ~(2_n7992 ^ 2_n8569);
assign 2_n4074 = 2_n8173 & 2_n3834;
assign 2_n3118 = 2_n4510 & 2_n6410;
assign 2_n11663 = ~(2_n12659 ^ 2_n6846);
assign 2_n1441 = 2_n12647 & 2_n11313;
assign 2_n2128 = 2_n12069 & 2_n1067;
assign 2_n7757 = 2_n11347 | 2_n6405;
assign 2_n11521 = 2_n11443 | 2_n11237;
assign 2_n597 = 2_n870 & 2_n1257;
assign 2_n12595 = ~(2_n3954 ^ 2_n8955);
assign 2_n6720 = 2_n5455 | 2_n7785;
assign 2_n7130 = 2_n5915 | 2_n9188;
assign 2_n445 = ~(2_n12491 ^ 2_n6657);
assign 2_n11282 = ~2_n9438;
assign 2_n4914 = ~(2_n5582 ^ 2_n1691);
assign 2_n8952 = 2_n5314 & 2_n806;
assign 2_n10020 = 2_n1031 & 2_n8378;
assign 2_n1629 = ~(2_n3216 ^ 2_n3120);
assign 2_n6976 = ~(2_n4057 | 2_n176);
assign 2_n1708 = 2_n4628 | 2_n8655;
assign 2_n6304 = 2_n1298 | 2_n11303;
assign 2_n8412 = ~(2_n1850 ^ 2_n12356);
assign 2_n1469 = 2_n1890 & 2_n3343;
assign 2_n6595 = ~2_n3000;
assign 2_n11340 = ~(2_n9836 ^ 2_n249);
assign 2_n9620 = ~(2_n7867 ^ 2_n2545);
assign 2_n8801 = ~2_n4337;
assign 2_n7844 = ~(2_n10884 ^ 2_n3143);
assign 2_n7116 = ~2_n2226;
assign 2_n11385 = ~(2_n7871 ^ 2_n6817);
assign 2_n10253 = ~(2_n2533 ^ 2_n3099);
assign 2_n5362 = ~2_n8670;
assign 2_n5558 = 2_n5236 & 2_n10301;
assign 2_n9938 = ~(2_n7323 ^ 2_n7518);
assign 2_n11525 = 2_n1432 | 2_n4923;
assign 2_n4798 = 2_n7774 & 2_n7127;
assign 2_n4461 = ~(2_n3196 | 2_n2274);
assign 2_n7309 = 2_n5355 | 2_n12843;
assign 2_n435 = ~(2_n2234 ^ 2_n12414);
assign 2_n7189 = ~(2_n10980 ^ 2_n4614);
assign 2_n12895 = 2_n2476 & 2_n9102;
assign 2_n7481 = ~(2_n9383 | 2_n8195);
assign 2_n1995 = 2_n686 | 2_n5540;
assign 2_n2787 = 2_n7550 & 2_n12390;
assign 2_n2655 = ~(2_n8603 | 2_n6969);
assign 2_n4103 = 2_n11905 | 2_n11186;
assign 2_n1293 = ~(2_n12914 | 2_n10920);
assign 2_n5374 = 2_n11292 | 2_n9517;
assign 2_n10291 = 2_n2784 & 2_n12315;
assign 2_n10746 = ~(2_n11613 | 2_n10710);
assign 2_n8397 = 2_n11966 | 2_n5091;
assign 2_n6354 = ~2_n6318;
assign 2_n2082 = ~2_n7699;
assign 2_n2533 = 2_n1825 & 2_n3229;
assign 2_n10331 = ~2_n9130;
assign 2_n11873 = 2_n4057 & 2_n176;
assign 2_n5994 = ~2_n2610;
assign 2_n4816 = 2_n9487 | 2_n3897;
assign 2_n12009 = 2_n10993 | 2_n8928;
assign 2_n12177 = 2_n3746 | 2_n7952;
assign 2_n1939 = ~(2_n3646 ^ 2_n1201);
assign 2_n4993 = 2_n6577 | 2_n11122;
assign 2_n7951 = 2_n10139 & 2_n3615;
assign 2_n5588 = ~(2_n4908 ^ 2_n12345);
assign 2_n7591 = 2_n10535 | 2_n1457;
assign 2_n3302 = 2_n4018 & 2_n9159;
assign 2_n4513 = ~(2_n5241 ^ 2_n245);
assign 2_n2712 = 2_n8034 | 2_n5868;
assign 2_n9442 = ~(2_n9337 ^ 2_n5587);
assign 2_n1876 = ~(2_n11760 ^ 2_n1301);
assign 2_n3537 = ~(2_n2684 | 2_n9962);
assign 2_n61 = 2_n5765 | 2_n6138;
assign 2_n6903 = 2_n11843 & 2_n6440;
assign 2_n9420 = ~2_n6899;
assign 2_n144 = 2_n12119 | 2_n12883;
assign 2_n1329 = ~(2_n7563 ^ 2_n6609);
assign 2_n9948 = 2_n9918 | 2_n7575;
assign 2_n9717 = ~(2_n2885 | 2_n11989);
assign 2_n6929 = 2_n10835 | 2_n5086;
assign 2_n7672 = 2_n4911 | 2_n12843;
assign 2_n5370 = 2_n11887 | 2_n1932;
assign 2_n10753 = 2_n2606 & 2_n11485;
assign 2_n5454 = ~(2_n452 ^ 2_n12646);
assign 2_n2199 = ~(2_n8180 ^ 2_n761);
assign 2_n8500 = ~(2_n9974 ^ 2_n3392);
assign 2_n479 = ~(2_n679 ^ 2_n9045);
assign 2_n8511 = 2_n7944 | 2_n2594;
assign 2_n7750 = 2_n10729 | 2_n8018;
assign 2_n5803 = ~2_n12081;
assign 2_n4879 = ~(2_n9538 ^ 2_n10503);
assign 2_n9479 = 2_n8354 | 2_n3224;
assign 2_n2808 = 2_n3018 & 2_n6810;
assign 2_n8159 = ~(2_n2043 ^ 2_n7717);
assign 2_n3822 = 2_n6560 | 2_n3741;
assign 2_n4491 = ~(2_n4815 ^ 2_n10041);
assign 2_n11926 = ~2_n7984;
assign 2_n10550 = ~(2_n3131 ^ 2_n10813);
assign 2_n4250 = 2_n8428 | 2_n3903;
assign 2_n5129 = ~(2_n1123 | 2_n396);
assign 2_n1144 = ~2_n7200;
assign 2_n3511 = 2_n11613 & 2_n10710;
assign 2_n6582 = 2_n319 | 2_n1234;
assign 2_n10590 = 2_n2217 | 2_n9280;
assign 2_n5560 = 2_n7380 | 2_n1634;
assign 2_n10251 = ~(2_n11280 | 2_n6141);
assign 2_n8302 = ~2_n1213;
assign 2_n4898 = ~(2_n6248 ^ 2_n3497);
assign 2_n4472 = 2_n2424 & 2_n12846;
assign 2_n9770 = 2_n2217 | 2_n3451;
assign 2_n4818 = ~2_n2802;
assign 2_n4682 = 2_n2176 ^ 2_n4779;
assign 2_n7451 = ~(2_n1598 ^ 2_n8724);
assign 2_n5865 = 2_n1272 & 2_n8761;
assign 2_n2854 = 2_n12853 | 2_n3924;
assign 2_n175 = 2_n1659 | 2_n4714;
assign 2_n6199 = 2_n5365 | 2_n479;
assign 2_n2691 = ~(2_n11499 ^ 2_n1216);
assign 2_n5782 = ~2_n4233;
assign 2_n11984 = 2_n191 | 2_n1546;
assign 2_n12465 = ~2_n6723;
assign 2_n8194 = 2_n9170 | 2_n1851;
assign 2_n2616 = 2_n7391 | 2_n5497;
assign 2_n5185 = ~2_n1339;
assign 2_n3816 = 2_n5828 | 2_n5186;
assign 2_n1340 = ~(2_n8052 | 2_n7989);
assign 2_n9881 = 2_n4002 | 2_n6061;
assign 2_n9330 = ~(2_n3386 ^ 2_n9746);
assign 2_n6375 = 2_n9459 | 2_n2193;
assign 2_n4772 = 2_n2931 & 2_n4376;
assign 2_n5059 = 2_n12541 & 2_n12031;
assign 2_n11479 = ~(2_n4918 ^ 2_n1268);
assign 2_n10935 = ~2_n11201;
assign 2_n3085 = ~(2_n6892 ^ 2_n12469);
assign 2_n7910 = ~(2_n12522 ^ 2_n12928);
assign 2_n7107 = 2_n9836 | 2_n8081;
assign 2_n2734 = ~2_n8702;
assign 2_n5281 = 2_n2872 | 2_n6455;
assign 2_n1057 = 2_n3746 | 2_n11775;
assign 2_n8555 = 2_n5895 & 2_n11374;
assign 2_n91 = 2_n3127 | 2_n1162;
assign 2_n3888 = ~(2_n1590 ^ 2_n1954);
assign 2_n1549 = ~2_n8562;
assign 2_n6557 = ~(2_n7481 | 2_n9494);
assign 2_n8570 = ~2_n3219;
assign 2_n11982 = ~(2_n8159 ^ 2_n2238);
assign 2_n12512 = 2_n2534 | 2_n4747;
assign 2_n1295 = ~(2_n9266 ^ 2_n8711);
assign 2_n560 = 2_n2140 | 2_n12656;
assign 2_n4475 = 2_n9450 & 2_n8067;
assign 2_n2758 = ~(2_n3943 ^ 2_n4262);
assign 2_n10202 = 2_n10157 | 2_n4875;
assign 2_n8754 = ~(2_n5604 ^ 2_n8837);
assign 2_n5446 = ~(2_n6697 ^ 2_n12225);
assign 2_n7349 = ~(2_n610 ^ 2_n5647);
assign 2_n8926 = 2_n9670 | 2_n10048;
assign 2_n10389 = 2_n8674 & 2_n5642;
assign 2_n11499 = ~(2_n9153 ^ 2_n8379);
assign 2_n3209 = ~(2_n4730 ^ 2_n12060);
assign 2_n859 = ~(2_n12355 ^ 2_n10125);
assign 2_n2372 = ~(2_n5267 ^ 2_n9406);
assign 2_n1666 = ~(2_n2359 | 2_n3212);
assign 2_n12182 = 2_n7116 | 2_n1413;
assign 2_n6527 = 2_n191 | 2_n11827;
assign 2_n12558 = 2_n11134 & 2_n401;
assign 2_n1000 = ~2_n8631;
assign 2_n11609 = ~(2_n4905 ^ 2_n620);
assign 2_n5527 = ~2_n8816;
assign 2_n1768 = ~(2_n3689 | 2_n9332);
assign 2_n11447 = ~(2_n4961 ^ 2_n231);
assign 2_n10845 = 2_n7862 & 2_n1798;
assign 2_n7974 = ~2_n1241;
assign 2_n11343 = ~2_n6626;
assign 2_n10288 = 2_n9373 | 2_n12120;
assign 2_n3193 = 2_n10040 | 2_n7990;
assign 2_n1138 = ~(2_n12461 ^ 2_n12672);
assign 2_n9023 = ~2_n1648;
assign 2_n3319 = ~(2_n10585 ^ 2_n8728);
assign 2_n11936 = 2_n7160 & 2_n11922;
assign 2_n12272 = ~(2_n6929 ^ 2_n275);
assign 2_n11398 = ~(2_n6836 ^ 2_n332);
assign 2_n8571 = ~(2_n2618 ^ 2_n4564);
assign 2_n2342 = ~(2_n2721 ^ 2_n11628);
assign 2_n3268 = ~(2_n12306 ^ 2_n9351);
assign 2_n8183 = ~2_n3689;
assign 2_n5406 = ~2_n7096;
assign 2_n5682 = 2_n8175 | 2_n11003;
assign 2_n12021 = ~2_n11275;
assign 2_n3154 = 2_n4603 | 2_n10468;
assign 2_n8437 = ~(2_n2677 ^ 2_n9579);
assign 2_n7982 = 2_n9301 | 2_n2028;
assign 2_n1660 = 2_n3127 | 2_n6389;
assign 2_n2056 = 2_n8870 | 2_n3924;
assign 2_n989 = ~2_n2564;
assign 2_n2709 = 2_n6625 & 2_n12959;
assign 2_n6390 = 2_n11278 & 2_n441;
assign 2_n1690 = ~(2_n10202 ^ 2_n6271);
assign 2_n8427 = ~(2_n3538 | 2_n682);
assign 2_n2952 = 2_n10879 | 2_n5497;
assign 2_n11918 = ~(2_n3689 ^ 2_n206);
assign 2_n11378 = 2_n4314 & 2_n9089;
assign 2_n5463 = ~2_n8990;
assign 2_n1187 = 2_n1337 & 2_n4054;
assign 2_n2014 = 2_n3252 | 2_n12542;
assign 2_n8148 = 2_n337 & 2_n12329;
assign 2_n463 = ~2_n1872;
assign 2_n3274 = 2_n8737 | 2_n5874;
assign 2_n625 = 2_n3648 & 2_n9664;
assign 2_n8365 = ~2_n4771;
assign 2_n9512 = 2_n6294 & 2_n2498;
assign 2_n5433 = ~(2_n2599 ^ 2_n1083);
assign 2_n3577 = 2_n10463 & 2_n5119;
assign 2_n12582 = ~(2_n3062 ^ 2_n2242);
assign 2_n6619 = ~(2_n3007 ^ 2_n8561);
assign 2_n322 = ~(2_n5169 ^ 2_n42);
assign 2_n313 = 2_n5765 | 2_n2020;
assign 2_n4697 = 2_n3127 | 2_n4242;
assign 2_n6465 = 2_n4085 & 2_n6000;
assign 2_n7933 = ~2_n7716;
assign 2_n2489 = ~(2_n11530 ^ 2_n8625);
assign 2_n7906 = 2_n1699 | 2_n8655;
assign 2_n4296 = ~(2_n8732 ^ 2_n1280);
assign 2_n12029 = ~2_n4742;
assign 2_n10749 = 2_n7370 | 2_n3125;
assign 2_n1674 = ~(2_n1953 ^ 2_n10276);
assign 2_n7307 = 2_n10555 & 2_n7791;
assign 2_n10706 = 2_n5107 & 2_n258;
assign 2_n10810 = 2_n994 | 2_n8859;
assign 2_n104 = ~(2_n1687 ^ 2_n3785);
assign 2_n10470 = 2_n1461 & 2_n3374;
assign 2_n937 = 2_n10847 & 2_n12626;
assign 2_n11345 = 2_n1102 & 2_n468;
assign 2_n7390 = 2_n12518 & 2_n10688;
assign 2_n7432 = 2_n9834 | 2_n7467;
assign 2_n10873 = ~(2_n3857 ^ 2_n9008);
assign 2_n2172 = ~(2_n5144 ^ 2_n5705);
assign 2_n9910 = ~(2_n2250 ^ 2_n1977);
assign 2_n3937 = 2_n7978 | 2_n9566;
assign 2_n3063 = ~(2_n969 ^ 2_n5046);
assign 2_n3170 = 2_n11290 & 2_n497;
assign 2_n4550 = 2_n8416 & 2_n2933;
assign 2_n8308 = 2_n5809 | 2_n7382;
assign 2_n12786 = 2_n10378 | 2_n2620;
assign 2_n908 = 2_n279 & 2_n2876;
assign 2_n7100 = 2_n5575 | 2_n7952;
assign 2_n1743 = 2_n12881 & 2_n10884;
assign 2_n10737 = 2_n8354 | 2_n5468;
assign 2_n2880 = ~(2_n4846 ^ 2_n11562);
assign 2_n6228 = ~(2_n1029 ^ 2_n8639);
assign 2_n9208 = 2_n1746 | 2_n2404;
assign 2_n9174 = 2_n6078 & 2_n2672;
assign 2_n1557 = ~2_n6834;
assign 2_n1101 = 2_n4290 | 2_n10113;
assign 2_n4553 = 2_n253 ^ 2_n11227;
assign 2_n6628 = 2_n12757 & 2_n5057;
assign 2_n7863 = ~(2_n7407 ^ 2_n10662);
assign 2_n2950 = 2_n5735 & 2_n1058;
assign 2_n5166 = 2_n2217 | 2_n795;
assign 2_n5291 = 2_n8276 & 2_n9640;
assign 2_n1758 = ~(2_n908 | 2_n6976);
assign 2_n8769 = ~(2_n12033 ^ 2_n6781);
assign 2_n10776 = ~(2_n5333 ^ 2_n257);
assign 2_n9826 = ~2_n9662;
assign 2_n2332 = 2_n5765 | 2_n10916;
assign 2_n7782 = 2_n10169 & 2_n1411;
assign 2_n10014 = ~(2_n6486 ^ 2_n1464);
assign 2_n198 = ~2_n5608;
assign 2_n79 = ~(2_n8295 ^ 2_n2862);
assign 2_n8197 = ~(2_n352 ^ 2_n8973);
assign 2_n6714 = 2_n4635 & 2_n12369;
assign 2_n4149 = ~2_n3775;
assign 2_n2454 = ~2_n3710;
assign 2_n12935 = 2_n2217 | 2_n8830;
assign 2_n11966 = 2_n2822 & 2_n5265;
assign 2_n1737 = 2_n7864 | 2_n8099;
assign 2_n2048 = ~(2_n5108 | 2_n9198);
assign 2_n12642 = 2_n10620 & 2_n11302;
assign 2_n12571 = 2_n4145 & 2_n11459;
assign 2_n7318 = 2_n3820 | 2_n2020;
assign 2_n670 = 2_n3465 & 2_n9147;
assign 2_n10666 = ~(2_n1899 ^ 2_n9575);
assign 2_n7514 = ~(2_n2424 ^ 2_n8822);
assign 2_n7643 = 2_n11958 | 2_n6114;
assign 2_n2568 = ~(2_n2130 ^ 2_n2037);
assign 2_n1116 = ~2_n10423;
assign 2_n12479 = ~2_n10255;
assign 2_n9265 = 2_n8384 & 2_n806;
assign 2_n3131 = 2_n2099 | 2_n530;
assign 2_n5260 = ~(2_n3030 ^ 2_n8394);
assign 2_n8453 = 2_n9674 | 2_n2691;
assign 2_n9604 = ~(2_n5229 | 2_n12653);
assign 2_n2233 = ~(2_n8591 ^ 2_n3731);
assign 2_n1477 = ~(2_n8960 | 2_n12466);
assign 2_n8232 = 2_n8026 | 2_n3468;
assign 2_n1085 = 2_n4943 | 2_n3189;
assign 2_n49 = 2_n3674 & 2_n1636;
assign 2_n6655 = ~(2_n9638 ^ 2_n3555);
assign 2_n4988 = ~(2_n4554 ^ 2_n3935);
assign 2_n1429 = ~(2_n11641 ^ 2_n6333);
assign 2_n3598 = ~(2_n11353 | 2_n10000);
assign 2_n6871 = 2_n11285 | 2_n6537;
assign 2_n3290 = 2_n78 | 2_n1934;
assign 2_n12703 = 2_n7495 | 2_n7424;
assign 2_n6909 = 2_n3591 | 2_n8082;
assign 2_n6360 = ~2_n3330;
assign 2_n7940 = 2_n12172 & 2_n7096;
assign 2_n967 = ~2_n2717;
assign 2_n3364 = 2_n5171 | 2_n4317;
assign 2_n5196 = 2_n10103 & 2_n411;
assign 2_n1967 = ~2_n12087;
assign 2_n6914 = 2_n3746 | 2_n7425;
assign 2_n3853 = 2_n11335 & 2_n6518;
assign 2_n6983 = ~(2_n1206 ^ 2_n5300);
assign 2_n9776 = 2_n11433 | 2_n2232;
assign 2_n1779 = ~(2_n2557 | 2_n10923);
assign 2_n9032 = ~(2_n128 ^ 2_n5460);
assign 2_n2120 = ~2_n157;
assign 2_n9246 = 2_n7388 & 2_n12947;
assign 2_n5842 = ~(2_n11745 ^ 2_n4969);
assign 2_n6786 = 2_n12391 & 2_n6806;
assign 2_n7527 = 2_n8583 | 2_n8643;
assign 2_n5595 = ~(2_n8568 ^ 2_n9116);
assign 2_n7980 = ~(2_n12901 | 2_n8105);
assign 2_n8691 = 2_n11719 | 2_n11746;
assign 2_n2801 = 2_n4445 | 2_n11105;
assign 2_n1769 = ~(2_n6500 ^ 2_n6593);
assign 2_n9886 = ~2_n8284;
assign 2_n5793 = 2_n12119 | 2_n6071;
assign 2_n1785 = ~(2_n5310 | 2_n5912);
assign 2_n3419 = ~(2_n6669 ^ 2_n3568);
assign 2_n4079 = 2_n11222 & 2_n9111;
assign 2_n983 = ~(2_n12795 ^ 2_n9407);
assign 2_n11103 = ~2_n3296;
assign 2_n2809 = ~(2_n6292 | 2_n9824);
assign 2_n3535 = ~(2_n5273 ^ 2_n108);
assign 2_n3351 = 2_n1726 & 2_n3718;
assign 2_n2791 = 2_n3743 | 2_n7921;
assign 2_n11389 = ~2_n5048;
assign 2_n290 = 2_n10006 | 2_n10659;
assign 2_n123 = ~(2_n3509 ^ 2_n1188);
assign 2_n2669 = 2_n2447 & 2_n9150;
assign 2_n8827 = ~(2_n787 ^ 2_n12944);
assign 2_n4002 = 2_n10142 | 2_n561;
assign 2_n9105 = 2_n6777 | 2_n2908;
assign 2_n52 = ~(2_n11856 ^ 2_n11998);
assign 2_n7217 = 2_n9172 & 2_n11949;
assign 2_n7174 = ~(2_n2285 ^ 2_n7801);
assign 2_n3194 = 2_n8127 | 2_n11827;
assign 2_n8382 = 2_n7123 | 2_n10074;
assign 2_n1161 = 2_n4956 | 2_n5000;
assign 2_n3662 = ~(2_n8810 ^ 2_n318);
assign 2_n2727 = 2_n1599 | 2_n11816;
assign 2_n8035 = 2_n3939 & 2_n1368;
assign 2_n2132 = ~(2_n12457 ^ 2_n3366);
assign 2_n5096 = 2_n9000 & 2_n5391;
assign 2_n4555 = 2_n7760 | 2_n11617;
assign 2_n10402 = 2_n12237 | 2_n10854;
assign 2_n6859 = 2_n2808 | 2_n11903;
assign 2_n905 = 2_n4498 | 2_n1079;
assign 2_n8874 = ~(2_n99 ^ 2_n11008);
assign 2_n8812 = 2_n9900 & 2_n5063;
assign 2_n306 = 2_n9373 | 2_n1509;
assign 2_n7143 = 2_n686 | 2_n12816;
assign 2_n6065 = 2_n4824 | 2_n11273;
assign 2_n6531 = 2_n3746 | 2_n1413;
assign 2_n9370 = ~2_n3172;
assign 2_n10324 = ~(2_n12165 ^ 2_n2720);
assign 2_n10421 = ~(2_n3189 ^ 2_n6176);
assign 2_n8784 = 2_n10572 & 2_n2741;
assign 2_n4929 = 2_n5739 | 2_n10241;
assign 2_n3428 = 2_n3096 | 2_n2232;
assign 2_n5520 = ~(2_n6449 | 2_n4626);
assign 2_n3031 = ~(2_n856 ^ 2_n7324);
assign 2_n2379 = 2_n12797 | 2_n6169;
assign 2_n1795 = ~(2_n9925 ^ 2_n8658);
assign 2_n12798 = ~(2_n3018 | 2_n6810);
assign 2_n7234 = 2_n12361 | 2_n11410;
assign 2_n12958 = ~2_n8912;
assign 2_n4782 = ~2_n9967;
assign 2_n4713 = 2_n6718 | 2_n609;
assign 2_n12848 = ~(2_n4741 | 2_n4384);
assign 2_n811 = 2_n5224 | 2_n3851;
assign 2_n4197 = 2_n9801 | 2_n8528;
assign 2_n5480 = ~(2_n12691 ^ 2_n306);
assign 2_n9576 = 2_n11552 | 2_n8643;
assign 2_n6649 = ~(2_n6129 | 2_n4700);
assign 2_n5687 = 2_n8498 | 2_n7279;
assign 2_n6000 = ~2_n10245;
assign 2_n4823 = ~(2_n1730 | 2_n1772);
assign 2_n7816 = ~2_n3204;
assign 2_n8329 = 2_n9690 & 2_n5546;
assign 2_n9263 = 2_n2107 & 2_n5239;
assign 2_n2484 = ~(2_n9296 ^ 2_n2712);
assign 2_n8538 = 2_n12231 & 2_n3958;
assign 2_n2696 = 2_n7912 | 2_n4136;
assign 2_n12504 = 2_n4668 | 2_n5572;
assign 2_n5928 = 2_n962 | 2_n1509;
assign 2_n4868 = ~(2_n3513 ^ 2_n10491);
assign 2_n106 = ~(2_n5947 ^ 2_n5261);
assign 2_n8346 = ~(2_n6379 | 2_n9484);
assign 2_n8133 = ~(2_n10613 ^ 2_n12740);
assign 2_n8208 = 2_n11958 | 2_n2754;
assign 2_n7873 = ~(2_n219 ^ 2_n10523);
assign 2_n12794 = 2_n10770 & 2_n4048;
assign 2_n8506 = 2_n11747 | 2_n4058;
assign 2_n8279 = 2_n37 | 2_n11316;
assign 2_n11016 = ~(2_n4512 ^ 2_n9986);
assign 2_n8015 = ~(2_n847 ^ 2_n11950);
assign 2_n8446 = 2_n9758 & 2_n9408;
assign 2_n8306 = 2_n931 | 2_n1735;
assign 2_n10635 = 2_n9420 & 2_n5665;
assign 2_n11882 = 2_n11433 | 2_n6169;
assign 2_n6212 = ~2_n10778;
assign 2_n11418 = ~2_n1776;
assign 2_n10189 = ~(2_n8677 ^ 2_n1369);
assign 2_n2389 = ~(2_n4462 ^ 2_n11363);
assign 2_n10286 = 2_n4678 | 2_n10234;
assign 2_n1583 = 2_n1670 | 2_n8700;
assign 2_n2586 = ~(2_n9865 ^ 2_n8654);
assign 2_n7342 = ~(2_n7566 ^ 2_n2932);
assign 2_n3182 = ~(2_n5998 ^ 2_n9577);
assign 2_n11276 = ~(2_n9205 ^ 2_n1069);
assign 2_n4192 = ~(2_n8310 ^ 2_n8450);
assign 2_n4847 = ~(2_n10926 ^ 2_n5600);
assign 2_n12740 = 2_n9584 | 2_n4474;
assign 2_n6371 = 2_n855 & 2_n10699;
assign 2_n8289 = ~(2_n4484 ^ 2_n1777);
assign 2_n6445 = ~(2_n9566 ^ 2_n336);
assign 2_n3844 = ~(2_n9937 ^ 2_n6224);
assign 2_n2810 = 2_n3746 | 2_n184;
assign 2_n9220 = ~(2_n4649 | 2_n8075);
assign 2_n4963 = ~(2_n8536 ^ 2_n1656);
assign 2_n4584 = 2_n8189 & 2_n5797;
assign 2_n590 = 2_n4434 & 2_n1584;
assign 2_n6798 = 2_n8757 & 2_n3021;
assign 2_n4807 = ~(2_n2948 ^ 2_n11083);
assign 2_n683 = 2_n12853 | 2_n12080;
assign 2_n9171 = 2_n7501 & 2_n1628;
assign 2_n496 = 2_n5915 | 2_n530;
assign 2_n802 = 2_n9887 & 2_n9226;
assign 2_n5206 = 2_n7258 & 2_n2988;
assign 2_n5021 = ~(2_n1552 ^ 2_n2091);
assign 2_n11874 = 2_n12691 | 2_n6543;
assign 2_n3040 = ~(2_n1563 | 2_n7062);
assign 2_n286 = ~(2_n4070 ^ 2_n4017);
assign 2_n4937 = ~(2_n7118 | 2_n4093);
assign 2_n146 = ~(2_n10243 ^ 2_n9707);
assign 2_n1399 = ~2_n4581;
assign 2_n10218 = ~(2_n1439 ^ 2_n4412);
assign 2_n12902 = ~(2_n4497 ^ 2_n731);
assign 2_n3872 = 2_n12180 | 2_n4558;
assign 2_n5017 = ~2_n6328;
assign 2_n11871 = ~(2_n6652 | 2_n6046);
assign 2_n6939 = 2_n10142 | 2_n4775;
assign 2_n8964 = 2_n9389 | 2_n1455;
assign 2_n6059 = 2_n4843 | 2_n11314;
assign 2_n10243 = ~(2_n7640 ^ 2_n2396);
assign 2_n6625 = 2_n5530 | 2_n8648;
assign 2_n3250 = 2_n6797 & 2_n12489;
assign 2_n4119 = 2_n8656 & 2_n3144;
assign 2_n2249 = 2_n2703 | 2_n850;
assign 2_n1816 = ~(2_n7501 | 2_n1628);
assign 2_n7232 = 2_n11400 & 2_n7590;
assign 2_n341 = ~2_n8754;
assign 2_n408 = ~(2_n2228 ^ 2_n5286);
assign 2_n968 = ~(2_n10795 | 2_n12909);
assign 2_n12557 = 2_n10835 | 2_n8745;
assign 2_n12765 = ~(2_n11140 ^ 2_n7163);
assign 2_n7173 = 2_n11445 & 2_n247;
assign 2_n755 = ~(2_n9674 ^ 2_n2691);
assign 2_n12502 = 2_n9341 & 2_n8154;
assign 2_n12688 = 2_n2693 & 2_n11525;
assign 2_n1784 = 2_n6373 | 2_n4474;
assign 2_n5707 = ~(2_n8372 ^ 2_n1480);
assign 2_n5841 = 2_n6977 | 2_n7425;
assign 2_n5807 = ~(2_n1088 ^ 2_n1479);
assign 2_n2360 = ~(2_n1398 ^ 2_n2338);
assign 2_n5598 = 2_n4022 & 2_n9318;
assign 2_n3093 = 2_n9389 | 2_n4400;
assign 2_n10183 = ~2_n8743;
assign 2_n8272 = 2_n5179 & 2_n8417;
assign 2_n6994 = ~(2_n3368 ^ 2_n1326);
assign 2_n12555 = ~2_n10493;
assign 2_n9821 = 2_n12910 | 2_n5296;
assign 2_n1285 = 2_n928 & 2_n6381;
assign 2_n85 = 2_n7895 & 2_n89;
assign 2_n6764 = ~2_n9872;
assign 2_n5092 = ~2_n4304;
assign 2_n3683 = ~(2_n589 ^ 2_n12321);
assign 2_n8711 = 2_n5915 | 2_n5468;
assign 2_n5138 = ~(2_n10070 | 2_n7997);
assign 2_n10412 = 2_n8894 | 2_n10256;
assign 2_n4023 = ~(2_n11429 ^ 2_n9761);
assign 2_n12770 = 2_n3970 & 2_n1364;
assign 2_n650 = ~(2_n12601 ^ 2_n4149);
assign 2_n7091 = 2_n1305 & 2_n1928;
assign 2_n885 = 2_n2099 | 2_n12124;
assign 2_n12451 = ~2_n10448;
assign 2_n6173 = 2_n2711 & 2_n2807;
assign 2_n6192 = ~(2_n7079 ^ 2_n9911);
assign 2_n8001 = ~(2_n11741 | 2_n1447);
assign 2_n12613 = ~2_n9419;
assign 2_n12942 = ~2_n2828;
assign 2_n10941 = 2_n6618 & 2_n12588;
assign 2_n2710 = ~(2_n392 | 2_n9940);
assign 2_n1216 = 2_n12197 & 2_n8637;
assign 2_n10397 = 2_n8896 & 2_n4710;
assign 2_n6349 = 2_n10338 & 2_n6123;
assign 2_n8542 = ~(2_n4268 ^ 2_n5586);
assign 2_n5950 = 2_n9074 & 2_n972;
assign 2_n11606 = ~(2_n3336 | 2_n3752);
assign 2_n11706 = 2_n12694 & 2_n7386;
assign 2_n11865 = ~(2_n7146 | 2_n7691);
assign 2_n5539 = ~(2_n9034 ^ 2_n11359);
assign 2_n12016 = ~(2_n7819 | 2_n7339);
assign 2_n12814 = 2_n8118 | 2_n9965;
assign 2_n11438 = 2_n111 | 2_n4618;
assign 2_n12546 = ~2_n6556;
assign 2_n12295 = ~(2_n6746 ^ 2_n3119);
assign 2_n5960 = ~2_n11345;
assign 2_n4763 = 2_n10339 | 2_n8740;
assign 2_n11376 = ~2_n6262;
assign 2_n11086 = ~(2_n9016 ^ 2_n10026);
assign 2_n9162 = ~(2_n8268 ^ 2_n10669);
assign 2_n7257 = ~(2_n11415 ^ 2_n12606);
assign 2_n5862 = ~2_n9380;
assign 2_n5877 = ~(2_n7620 | 2_n1724);
assign 2_n8625 = ~(2_n2400 ^ 2_n2705);
assign 2_n8007 = ~(2_n10403 | 2_n6870);
assign 2_n10374 = 2_n5355 | 2_n11430;
assign 2_n4876 = ~(2_n6406 | 2_n3542);
assign 2_n312 = 2_n2762 & 2_n5782;
assign 2_n3543 = ~(2_n6187 ^ 2_n7403);
assign 2_n12833 = ~(2_n6390 | 2_n8238);
assign 2_n8507 = 2_n1396 & 2_n10946;
assign 2_n7223 = 2_n10147 | 2_n12838;
assign 2_n6006 = 2_n9079 & 2_n6414;
assign 2_n8917 = ~(2_n2957 ^ 2_n3671);
assign 2_n5058 = 2_n11043 | 2_n9721;
assign 2_n6878 = ~2_n11749;
assign 2_n6998 = 2_n678 & 2_n1703;
assign 2_n3423 = ~(2_n4346 ^ 2_n1308);
assign 2_n8681 = ~(2_n10036 ^ 2_n3526);
assign 2_n11172 = ~(2_n7229 ^ 2_n10749);
assign 2_n5426 = ~2_n1373;
assign 2_n12400 = 2_n249 | 2_n11480;
assign 2_n12008 = ~(2_n6081 ^ 2_n12609);
assign 2_n7463 = ~(2_n9581 ^ 2_n10924);
assign 2_n887 = ~(2_n12258 ^ 2_n4705);
assign 2_n5348 = 2_n9373 | 2_n28;
assign 2_n12623 = 2_n5303 & 2_n3393;
assign 2_n4075 = 2_n807 | 2_n2815;
assign 2_n12397 = ~2_n3895;
assign 2_n5220 = ~(2_n229 ^ 2_n11915);
assign 2_n1433 = 2_n1941 | 2_n11896;
assign 2_n10045 = 2_n2459 | 2_n4594;
assign 2_n7081 = 2_n5677 & 2_n11125;
assign 2_n3863 = ~(2_n6237 ^ 2_n12917);
assign 2_n3315 = ~(2_n12308 ^ 2_n227);
assign 2_n11515 = ~(2_n8999 ^ 2_n11371);
assign 2_n9553 = ~(2_n11724 ^ 2_n9919);
assign 2_n3510 = 2_n2602 & 2_n4014;
assign 2_n11979 = ~(2_n5277 | 2_n7517);
assign 2_n5613 = ~(2_n4700 ^ 2_n6129);
assign 2_n10404 = 2_n3326 & 2_n2364;
assign 2_n11337 = ~(2_n7401 ^ 2_n6412);
assign 2_n5135 = ~(2_n4247 ^ 2_n554);
assign 2_n2599 = 2_n5575 | 2_n11410;
assign 2_n3752 = ~(2_n1859 ^ 2_n12339);
assign 2_n6748 = ~(2_n1878 ^ 2_n10861);
assign 2_n12873 = 2_n7449 | 2_n6138;
assign 2_n2708 = ~(2_n7749 ^ 2_n3281);
assign 2_n12056 = 2_n4602 & 2_n2676;
assign 2_n11801 = 2_n11026 | 2_n4875;
assign 2_n2532 = ~(2_n1722 ^ 2_n1055);
assign 2_n773 = 2_n11389 | 2_n1159;
assign 2_n9302 = ~2_n7177;
assign 2_n460 = ~(2_n1339 ^ 2_n6299);
assign 2_n4025 = ~(2_n6569 | 2_n12796);
assign 2_n4 = 2_n270 | 2_n11231;
assign 2_n8966 = 2_n6031 | 2_n3787;
assign 2_n6438 = ~(2_n7564 ^ 2_n8019);
assign 2_n7544 = 2_n1966 | 2_n7784;
assign 2_n7262 = ~(2_n1672 ^ 2_n2553);
assign 2_n3942 = ~(2_n2345 ^ 2_n8444);
assign 2_n3173 = ~(2_n2555 ^ 2_n12042);
assign 2_n204 = 2_n4777 | 2_n7475;
assign 2_n7367 = ~2_n3604;
assign 2_n2597 = 2_n7688 | 2_n11465;
assign 2_n10582 = ~2_n1151;
assign 2_n1099 = 2_n763 | 2_n5976;
assign 2_n5057 = ~2_n12118;
assign 2_n4692 = ~2_n1687;
assign 2_n1891 = ~(2_n3048 | 2_n5978);
assign 2_n6791 = ~(2_n2854 ^ 2_n7701);
assign 2_n7821 = ~(2_n292 ^ 2_n2428);
assign 2_n11381 = 2_n8438 | 2_n12190;
assign 2_n11011 = ~2_n6209;
assign 2_n6497 = ~(2_n1348 ^ 2_n10372);
assign 2_n4599 = ~2_n8963;
assign 2_n784 = 2_n8481 & 2_n1048;
assign 2_n9579 = 2_n8572 & 2_n11579;
assign 2_n11534 = 2_n3558 | 2_n1927;
assign 2_n3260 = 2_n989 | 2_n1162;
assign 2_n12888 = ~2_n39;
assign 2_n378 = ~2_n10155;
assign 2_n9168 = ~(2_n10061 | 2_n10316);
assign 2_n9417 = ~2_n10362;
assign 2_n9994 = ~(2_n3620 ^ 2_n5718);
assign 2_n4733 = ~(2_n12019 ^ 2_n8661);
assign 2_n10605 = ~(2_n12464 ^ 2_n2122);
assign 2_n1582 = 2_n1871 & 2_n3515;
assign 2_n5504 = ~(2_n495 ^ 2_n1189);
assign 2_n2840 = 2_n5414 | 2_n10759;
assign 2_n109 = ~2_n5517;
assign 2_n4523 = ~(2_n4514 ^ 2_n7677);
assign 2_n2770 = ~(2_n2842 | 2_n6424);
assign 2_n9045 = ~(2_n5328 ^ 2_n2683);
assign 2_n695 = 2_n2217 | 2_n4864;
assign 2_n9389 = ~2_n4189;
assign 2_n12022 = 2_n12960 & 2_n10487;
assign 2_n542 = 2_n725 & 2_n8146;
assign 2_n3569 = 2_n5765 | 2_n28;
assign 2_n4341 = ~(2_n10180 ^ 2_n4234);
assign 2_n5046 = 2_n7439 & 2_n5891;
assign 2_n12600 = ~(2_n10226 ^ 2_n9680);
assign 2_n6861 = 2_n607 & 2_n419;
assign 2_n5435 = ~(2_n1385 ^ 2_n4009);
assign 2_n4213 = ~(2_n588 ^ 2_n156);
assign 2_n3048 = ~2_n37;
assign 2_n314 = ~(2_n8789 ^ 2_n1733);
assign 2_n11468 = 2_n6718 | 2_n4642;
assign 2_n9147 = ~2_n7131;
assign 2_n11611 = ~2_n1865;
assign 2_n7786 = ~2_n1264;
assign 2_n179 = ~(2_n5023 ^ 2_n10401);
assign 2_n7920 = 2_n11220 & 2_n7829;
assign 2_n11786 = ~(2_n3879 | 2_n10499);
assign 2_n9014 = 2_n2479 & 2_n2317;
assign 2_n4587 = ~2_n7642;
assign 2_n11884 = 2_n4565 | 2_n1281;
assign 2_n11191 = ~2_n2861;
assign 2_n5757 = 2_n9370 | 2_n510;
assign 2_n9817 = 2_n24 & 2_n7334;
assign 2_n9769 = ~(2_n8232 | 2_n7679);
assign 2_n6326 = ~(2_n6233 ^ 2_n11513);
assign 2_n2273 = ~(2_n5423 ^ 2_n9921);
assign 2_n11930 = 2_n9370 | 2_n11746;
assign 2_n10966 = ~2_n2311;
assign 2_n5339 = ~2_n7775;
assign 2_n1650 = ~(2_n7864 ^ 2_n8099);
assign 2_n3310 = 2_n7116 | 2_n11775;
assign 2_n7393 = 2_n5530 | 2_n12883;
assign 2_n8863 = ~(2_n6694 ^ 2_n11733);
assign 2_n11639 = ~(2_n10876 | 2_n10982);
assign 2_n5884 = 2_n5679 & 2_n2963;
assign 2_n4164 = ~2_n4920;
assign 2_n12779 = ~(2_n2903 ^ 2_n10734);
assign 2_n6534 = 2_n8026 | 2_n3903;
assign 2_n6392 = ~(2_n10341 ^ 2_n6357);
assign 2_n4422 = ~(2_n5090 ^ 2_n1993);
assign 2_n9453 = ~(2_n12658 ^ 2_n8392);
assign 2_n10453 = 2_n2832 | 2_n1455;
assign 2_n3645 = ~(2_n4580 | 2_n7561);
assign 2_n9348 = 2_n7028 & 2_n898;
assign 2_n9911 = ~(2_n3811 ^ 2_n7135);
assign 2_n6114 = ~2_n7730;
assign 2_n6474 = 2_n9052 & 2_n2716;
assign 2_n2163 = 2_n4343 | 2_n6513;
assign 2_n2429 = 2_n4605 & 2_n1678;
assign 2_n6900 = 2_n8428 | 2_n7395;
assign 2_n2205 = ~(2_n1341 ^ 2_n3362);
assign 2_n2778 = ~(2_n2045 ^ 2_n11274);
assign 2_n7284 = 2_n2456 | 2_n8655;
assign 2_n7767 = ~2_n4529;
assign 2_n12783 = ~(2_n12091 ^ 2_n12682);
assign 2_n6322 = ~(2_n5149 ^ 2_n6035);
assign 2_n4875 = ~2_n4086;
assign 2_n6430 = 2_n7834 & 2_n8364;
assign 2_n5235 = ~(2_n7121 ^ 2_n8944);
assign 2_n2036 = 2_n5915 | 2_n3924;
assign 2_n688 = 2_n1051 | 2_n995;
assign 2_n6485 = ~2_n9054;
assign 2_n4068 = 2_n9027 & 2_n1588;
assign 2_n1726 = 2_n10142 | 2_n1851;
assign 2_n3238 = ~(2_n12563 ^ 2_n9703);
assign 2_n4429 = ~(2_n1411 ^ 2_n1925);
assign 2_n12042 = ~(2_n12035 ^ 2_n6063);
assign 2_n6551 = 2_n8690 & 2_n3904;
assign 2_n4942 = ~(2_n8219 ^ 2_n6815);
assign 2_n12513 = 2_n7449 | 2_n609;
assign 2_n909 = ~(2_n4525 ^ 2_n11382);
assign 2_n11353 = 2_n1025 & 2_n4933;
assign 2_n9216 = 2_n15 | 2_n5218;
assign 2_n11298 = ~(2_n3665 ^ 2_n9355);
assign 2_n5870 = ~(2_n12571 ^ 2_n619);
assign 2_n9020 = ~(2_n1583 ^ 2_n4473);
assign 2_n2305 = 2_n752 | 2_n5540;
assign 2_n5624 = ~(2_n940 ^ 2_n9984);
assign 2_n11680 = 2_n1043 | 2_n11532;
assign 2_n1530 = ~(2_n1754 | 2_n2291);
assign 2_n7656 = 2_n11576 & 2_n1712;
assign 2_n9711 = ~(2_n8331 ^ 2_n5351);
assign 2_n5459 = 2_n12497 & 2_n7033;
assign 2_n4984 = ~(2_n2610 ^ 2_n9541);
assign 2_n7303 = 2_n2456 | 2_n4913;
assign 2_n7964 = 2_n2136 | 2_n10652;
assign 2_n11718 = ~(2_n7448 | 2_n3231);
assign 2_n8257 = ~2_n12571;
assign 2_n5308 = ~(2_n2447 ^ 2_n2313);
assign 2_n9996 = 2_n5680 & 2_n4883;
assign 2_n9868 = ~(2_n7487 ^ 2_n8251);
assign 2_n6298 = 2_n9564 & 2_n706;
assign 2_n4980 = 2_n10339 | 2_n6513;
assign 2_n10708 = ~(2_n9245 ^ 2_n8383);
assign 2_n12231 = 2_n3989 & 2_n5970;
assign 2_n10934 = 2_n5765 | 2_n9280;
assign 2_n7599 = 2_n8738 | 2_n4654;
assign 2_n7271 = 2_n3743 | 2_n9078;
assign 2_n10900 = 2_n12142 & 2_n4458;
assign 2_n6814 = 2_n5355 | 2_n1738;
assign 2_n1539 = ~2_n2087;
assign 2_n11709 = 2_n6863 | 2_n4427;
assign 2_n6219 = 2_n2376 | 2_n3679;
assign 2_n2630 = 2_n12748 | 2_n1336;
assign 2_n4992 = 2_n9389 | 2_n5497;
assign 2_n267 = ~(2_n956 ^ 2_n8680);
assign 2_n3176 = 2_n5738 & 2_n9642;
assign 2_n1821 = 2_n7562 & 2_n12889;
assign 2_n8776 = ~(2_n8975 ^ 2_n1619);
assign 2_n12425 = 2_n7713 & 2_n4012;
assign 2_n6506 = 2_n5689 & 2_n10134;
assign 2_n11380 = ~(2_n7920 ^ 2_n8715);
assign 2_n4411 = ~2_n1723;
assign 2_n266 = 2_n2865 | 2_n1942;
assign 2_n3041 = ~(2_n4446 | 2_n1491);
assign 2_n5011 = 2_n4559 | 2_n10651;
assign 2_n493 = 2_n6395 | 2_n2806;
assign 2_n643 = ~(2_n5087 | 2_n5357);
assign 2_n558 = 2_n11069 & 2_n10056;
assign 2_n7113 = 2_n7624 | 2_n3139;
assign 2_n8424 = ~(2_n5673 ^ 2_n8784);
assign 2_n4519 = 2_n22 | 2_n5261;
assign 2_n12303 = 2_n8211 & 2_n12745;
assign 2_n11278 = 2_n526 | 2_n12480;
assign 2_n2241 = ~(2_n122 ^ 2_n11504);
assign 2_n3276 = 2_n1886 & 2_n4382;
assign 2_n8586 = ~(2_n3749 ^ 2_n8995);
assign 2_n3263 = ~(2_n140 ^ 2_n7811);
assign 2_n7442 = ~(2_n3807 ^ 2_n1967);
assign 2_n7947 = 2_n9231 | 2_n6051;
assign 2_n1134 = ~2_n634;
assign 2_n6857 = 2_n6373 | 2_n3606;
assign 2_n9597 = ~(2_n694 | 2_n1527);
assign 2_n11052 = ~(2_n4122 ^ 2_n4225);
assign 2_n634 = 2_n556 & 2_n9483;
assign 2_n3846 = 2_n5850 & 2_n1347;
assign 2_n9603 = 2_n11478 & 2_n12489;
assign 2_n8301 = ~2_n1242;
assign 2_n613 = 2_n10142 | 2_n12843;
assign 2_n406 = ~2_n8914;
assign 2_n11544 = 2_n10157 | 2_n6922;
assign 2_n8064 = 2_n5542 & 2_n7234;
assign 2_n11081 = ~(2_n11276 ^ 2_n5298);
assign 2_n9795 = 2_n10199 & 2_n7637;
assign 2_n12617 = ~2_n9519;
assign 2_n10875 = ~(2_n2781 ^ 2_n2132);
assign 2_n2544 = ~(2_n11679 ^ 2_n1702);
assign 2_n12538 = ~(2_n3065 | 2_n577);
assign 2_n10105 = 2_n5999 | 2_n7753;
assign 2_n4276 = ~(2_n12788 ^ 2_n1120);
assign 2_n969 = 2_n7391 | 2_n1079;
assign 2_n7103 = ~(2_n9887 ^ 2_n9226);
assign 2_n6377 = 2_n1881 | 2_n3482;
assign 2_n5488 = 2_n3051 | 2_n2323;
assign 2_n12227 = 2_n4628 | 2_n3924;
assign 2_n12186 = ~2_n10644;
assign 2_n5946 = ~2_n935;
assign 2_n353 = ~(2_n8242 ^ 2_n6266);
assign 2_n8440 = ~(2_n3138 ^ 2_n5747);
assign 2_n4087 = ~(2_n9228 ^ 2_n776);
assign 2_n3966 = ~(2_n8534 ^ 2_n12791);
assign 2_n1425 = 2_n6571 | 2_n11787;
assign 2_n417 = ~(2_n7501 ^ 2_n5037);
assign 2_n4540 = ~2_n8163;
assign 2_n10917 = 2_n8097 & 2_n3621;
assign 2_n11522 = ~(2_n331 ^ 2_n9121);
assign 2_n10146 = 2_n9431 & 2_n421;
assign 2_n6351 = 2_n6635 & 2_n9863;
assign 2_n10995 = 2_n12797 | 2_n2815;
assign 2_n881 = 2_n12933 & 2_n4152;
assign 2_n1847 = ~(2_n3521 ^ 2_n6605);
assign 2_n11327 = 2_n10251 | 2_n7741;
assign 2_n9507 = 2_n10551 & 2_n7988;
assign 2_n1262 = ~(2_n9784 ^ 2_n945);
assign 2_n4727 = 2_n8336 & 2_n12709;
assign 2_n6824 = 2_n12141 & 2_n11811;
assign 2_n2223 = 2_n5809 | 2_n12735;
assign 2_n8519 = ~2_n4650;
assign 2_n9485 = 2_n11821 & 2_n1798;
assign 2_n12174 = ~(2_n1808 ^ 2_n2210);
assign 2_n1846 = ~(2_n3474 | 2_n5126);
assign 2_n6512 = ~(2_n4017 | 2_n4070);
assign 2_n338 = 2_n11782 & 2_n5114;
assign 2_n12270 = ~(2_n5791 ^ 2_n3300);
assign 2_n9104 = ~2_n6988;
assign 2_n158 = 2_n4911 | 2_n7881;
assign 2_n11858 = 2_n3196 ^ 2_n10766;
assign 2_n8903 = 2_n5575 | 2_n10903;
assign 2_n1717 = ~2_n5948;
assign 2_n11678 = 2_n4961 & 2_n231;
assign 2_n11627 = ~2_n9395;
assign 2_n10642 = 2_n8921 | 2_n1555;
assign 2_n1072 = 2_n5355 | 2_n6402;
assign 2_n6501 = 2_n4243 & 2_n8520;
assign 2_n921 = ~(2_n7936 | 2_n1021);
assign 2_n5642 = 2_n3756 & 2_n2970;
assign 2_n9530 = 2_n10196 | 2_n4474;
assign 2_n5771 = 2_n1462 | 2_n10617;
assign 2_n9572 = 2_n6376 & 2_n7343;
assign 2_n12499 = ~2_n9896;
assign 2_n6448 = ~(2_n8675 | 2_n9295);
assign 2_n8392 = 2_n6888 & 2_n11121;
assign 2_n8794 = 2_n7058 & 2_n6484;
assign 2_n9647 = ~(2_n11392 ^ 2_n10994);
assign 2_n6405 = ~(2_n2303 ^ 2_n6676);
assign 2_n7277 = 2_n11126 & 2_n687;
assign 2_n8969 = ~2_n4756;
assign 2_n9786 = 2_n2595 | 2_n920;
assign 2_n11109 = 2_n6977 | 2_n3421;
assign 2_n3218 = 2_n8552 | 2_n10854;
assign 2_n9646 = ~(2_n11094 ^ 2_n7005);
assign 2_n11258 = ~(2_n9176 ^ 2_n11849);
assign 2_n3575 = ~(2_n7527 ^ 2_n5344);
assign 2_n899 = 2_n10157 | 2_n5759;
assign 2_n2378 = 2_n1663 & 2_n4964;
assign 2_n1490 = ~(2_n3403 ^ 2_n3675);
assign 2_n4347 = 2_n12841 | 2_n6563;
assign 2_n7912 = 2_n7283 | 2_n7881;
assign 2_n8048 = 2_n659 | 2_n2151;
assign 2_n2110 = ~(2_n5358 ^ 2_n764);
assign 2_n9872 = 2_n7177 & 2_n8407;
assign 2_n11561 = ~(2_n9894 ^ 2_n5047);
assign 2_n12863 = ~(2_n10377 ^ 2_n11);
assign 2_n4827 = 2_n6931 & 2_n4506;
assign 2_n2209 = 2_n5355 | 2_n11827;
assign 2_n4908 = 2_n2538 & 2_n2861;
assign 2_n8585 = 2_n12119 | 2_n10854;
assign 2_n12576 = 2_n6579 & 2_n3093;
assign 2_n5340 = 2_n8371 | 2_n4073;
assign 2_n6178 = ~(2_n8579 ^ 2_n1647);
assign 2_n1439 = 2_n6743 & 2_n4503;
assign 2_n9875 = 2_n9653 | 2_n3928;
assign 2_n9356 = ~(2_n4949 ^ 2_n3083);
assign 2_n4096 = ~2_n5380;
assign 2_n8483 = ~(2_n9799 ^ 2_n12802);
assign 2_n3087 = 2_n10750 | 2_n826;
assign 2_n3954 = 2_n12237 | 2_n1932;
assign 2_n9139 = ~(2_n2028 ^ 2_n3245);
assign 2_n8930 = ~(2_n7587 ^ 2_n10511);
assign 2_n12072 = ~(2_n5523 ^ 2_n12349);
assign 2_n11238 = ~2_n8660;
assign 2_n9151 = 2_n9835 | 2_n11151;
assign 2_n254 = ~2_n4135;
assign 2_n10570 = 2_n7899 & 2_n5485;
assign 2_n12580 = ~2_n3945;
assign 2_n11887 = ~2_n6797;
assign 2_n1194 = ~(2_n12155 ^ 2_n10506);
assign 2_n7916 = 2_n10142 | 2_n9589;
assign 2_n7797 = 2_n9849 & 2_n8268;
assign 2_n8444 = ~(2_n4110 ^ 2_n11565);
assign 2_n1856 = 2_n6277 & 2_n8368;
assign 2_n6505 = ~2_n5869;
assign 2_n6116 = ~(2_n4360 ^ 2_n702);
assign 2_n7247 = ~(2_n11899 ^ 2_n477);
assign 2_n11074 = 2_n4932 | 2_n12548;
assign 2_n11388 = 2_n9454 & 2_n6302;
assign 2_n3794 = ~(2_n5877 | 2_n653);
assign 2_n2807 = 2_n11608 | 2_n6029;
assign 2_n2816 = 2_n8617 | 2_n2375;
assign 2_n10290 = 2_n11521 & 2_n7438;
assign 2_n5351 = ~2_n6574;
assign 2_n11711 = 2_n3197 & 2_n6057;
assign 2_n10639 = 2_n12178 & 2_n5402;
assign 2_n11653 = 2_n2579 | 2_n4751;
assign 2_n3275 = ~2_n4664;
assign 2_n3636 = ~2_n12068;
assign 2_n7718 = 2_n11923 | 2_n4474;
assign 2_n12665 = 2_n854 | 2_n1710;
assign 2_n9590 = 2_n12299 & 2_n11023;
assign 2_n6132 = 2_n8738 | 2_n28;
assign 2_n798 = ~(2_n1853 ^ 2_n1577);
assign 2_n710 = ~(2_n2777 ^ 2_n10319);
assign 2_n8892 = ~(2_n4998 ^ 2_n6646);
assign 2_n10214 = ~(2_n82 ^ 2_n3917);
assign 2_n7895 = 2_n1629 | 2_n11103;
assign 2_n4974 = 2_n3461 | 2_n8923;
assign 2_n11781 = ~(2_n3471 ^ 2_n355);
assign 2_n9320 = ~(2_n504 ^ 2_n8915);
assign 2_n9824 = ~2_n2869;
assign 2_n4687 = ~(2_n7144 ^ 2_n4713);
assign 2_n3053 = ~2_n3396;
assign 2_n7424 = ~2_n12720;
assign 2_n5778 = 2_n264 | 2_n3350;
assign 2_n11647 = ~(2_n5882 | 2_n786);
assign 2_n11864 = 2_n12853 | 2_n9188;
assign 2_n7731 = ~2_n7401;
assign 2_n3716 = 2_n12501 & 2_n7631;
assign 2_n4648 = ~2_n10167;
assign 2_n6741 = 2_n5466 & 2_n4578;
assign 2_n2220 = 2_n876 | 2_n11561;
assign 2_n5330 = 2_n375 | 2_n11346;
assign 2_n9251 = ~(2_n12632 ^ 2_n2990);
assign 2_n8870 = ~2_n7160;
assign 2_n2261 = 2_n4488 | 2_n11502;
assign 2_n1164 = ~2_n7252;
assign 2_n11227 = ~(2_n6239 ^ 2_n8808);
assign 2_n5554 = 2_n3587 | 2_n2295;
assign 2_n12219 = 2_n1333 & 2_n6038;
assign 2_n10299 = ~(2_n7916 ^ 2_n2642);
assign 2_n12860 = ~(2_n6635 ^ 2_n9193);
assign 2_n12055 = ~(2_n11303 ^ 2_n1614);
assign 2_n3821 = 2_n6849 | 2_n10786;
assign 2_n7198 = 2_n8002 & 2_n8934;
assign 2_n9472 = 2_n8390 | 2_n2744;
assign 2_n1069 = ~(2_n7756 ^ 2_n4681);
assign 2_n9230 = ~(2_n1260 ^ 2_n1053);
assign 2_n11383 = ~(2_n2073 ^ 2_n8420);
assign 2_n1154 = 2_n2217 | 2_n5086;
assign 2_n11140 = ~(2_n5801 ^ 2_n4160);
assign 2_n10535 = 2_n10938 | 2_n5356;
assign 2_n7252 = ~(2_n12268 ^ 2_n4486);
assign 2_n113 = 2_n2033 & 2_n8014;
assign 2_n11839 = ~(2_n9324 | 2_n12805);
assign 2_n11454 = ~(2_n7083 ^ 2_n12586);
assign 2_n4089 = 2_n3746 | 2_n12816;
assign 2_n3159 = ~(2_n8143 ^ 2_n976);
assign 2_n903 = 2_n5940 & 2_n6495;
assign 2_n3437 = ~(2_n12387 ^ 2_n4258);
assign 2_n11642 = 2_n12886 & 2_n4117;
assign 2_n8904 = ~(2_n5428 ^ 2_n2647);
assign 2_n2492 = ~(2_n8193 ^ 2_n4752);
assign 2_n7351 = ~2_n9059;
assign 2_n7415 = ~(2_n2704 ^ 2_n6163);
assign 2_n5313 = ~(2_n11080 ^ 2_n3441);
assign 2_n11041 = 2_n8377 & 2_n5770;
assign 2_n5750 = ~(2_n8736 ^ 2_n6643);
assign 2_n6678 = ~2_n3910;
assign 2_n1214 = 2_n5650 & 2_n11675;
assign 2_n9459 = 2_n12841 & 2_n6563;
assign 2_n1259 = 2_n4633 & 2_n6062;
assign 2_n2835 = ~(2_n2779 | 2_n8001);
assign 2_n10566 = ~(2_n2869 ^ 2_n6292);
assign 2_n8168 = ~(2_n10320 | 2_n2747);
assign 2_n5479 = ~2_n2100;
assign 2_n2980 = 2_n9370 | 2_n12843;
assign 2_n8771 = ~(2_n5023 | 2_n4063);
assign 2_n6756 = 2_n2906 | 2_n6213;
assign 2_n2693 = ~(2_n9778 ^ 2_n4240);
assign 2_n10333 = 2_n4469 & 2_n1428;
assign 2_n12938 = 2_n9563 | 2_n3881;
assign 2_n340 = ~(2_n8795 ^ 2_n12151);
assign 2_n5277 = 2_n9389 | 2_n12328;
assign 2_n1804 = ~(2_n5122 ^ 2_n10977);
assign 2_n4734 = 2_n6770 & 2_n2508;
assign 2_n936 = 2_n5177 & 2_n10438;
assign 2_n5534 = ~(2_n7684 ^ 2_n12162);
assign 2_n9560 = 2_n673 & 2_n7022;
assign 2_n2310 = ~(2_n2502 ^ 2_n11123);
assign 2_n9680 = ~2_n6768;
assign 2_n1625 = 2_n10612 & 2_n12938;
assign 2_n4781 = 2_n4212 & 2_n4350;
assign 2_n11868 = ~2_n4991;
assign 2_n8578 = ~(2_n2945 ^ 2_n5725);
assign 2_n7046 = 2_n9043 | 2_n10840;
assign 2_n5581 = ~(2_n2897 ^ 2_n12421);
assign 2_n11816 = 2_n8583 | 2_n12771;
assign 2_n1241 = 2_n994 | 2_n10419;
assign 2_n6385 = 2_n9616 & 2_n5262;
assign 2_n8670 = 2_n1239 & 2_n5737;
assign 2_n5510 = ~(2_n7563 | 2_n9272);
assign 2_n472 = ~(2_n2761 ^ 2_n1190);
assign 2_n220 = ~2_n3264;
assign 2_n9641 = ~(2_n10728 ^ 2_n8985);
assign 2_n5297 = ~(2_n12717 ^ 2_n10156);
assign 2_n3923 = ~(2_n7310 ^ 2_n11202);
assign 2_n2405 = 2_n10339 | 2_n9188;
assign 2_n12173 = 2_n11259 | 2_n6119;
assign 2_n2531 = ~2_n12276;
assign 2_n7777 = 2_n752 | 2_n10919;
assign 2_n4379 = ~(2_n11957 ^ 2_n7460);
assign 2_n6071 = ~2_n503;
assign 2_n992 = ~(2_n4977 ^ 2_n104);
assign 2_n7446 = ~(2_n11555 ^ 2_n11609);
assign 2_n3585 = 2_n7839 | 2_n6169;
assign 2_n7041 = ~2_n7566;
assign 2_n10040 = ~(2_n1810 | 2_n10778);
assign 2_n7913 = 2_n4992 | 2_n875;
assign 2_n10788 = ~(2_n7215 ^ 2_n4269);
assign 2_n2027 = ~(2_n6567 ^ 2_n11161);
assign 2_n3394 = 2_n4675 & 2_n5818;
assign 2_n5940 = 2_n12467 | 2_n918;
assign 2_n3987 = ~(2_n9366 ^ 2_n3063);
assign 2_n4654 = ~2_n405;
assign 2_n3090 = ~(2_n11221 ^ 2_n3260);
assign 2_n12666 = 2_n4180 & 2_n4990;
assign 2_n8530 = ~2_n2342;
assign 2_n12691 = 2_n6718 | 2_n1047;
assign 2_n2339 = 2_n12479 & 2_n8174;
assign 2_n11904 = ~(2_n10118 ^ 2_n5601);
assign 2_n10188 = ~2_n12637;
assign 2_n11780 = ~(2_n11241 ^ 2_n2062);
assign 2_n8274 = 2_n3127 | 2_n11746;
assign 2_n626 = ~(2_n12271 ^ 2_n12707);
assign 2_n4748 = ~(2_n1872 ^ 2_n625);
assign 2_n8710 = ~(2_n4239 | 2_n5998);
assign 2_n12366 = 2_n7071 & 2_n8338;
assign 2_n10367 = 2_n8870 | 2_n10422;
assign 2_n6944 = ~2_n9487;
assign 2_n1747 = 2_n349 | 2_n3520;
assign 2_n4180 = ~2_n9869;
assign 2_n5178 = 2_n4294 | 2_n1120;
assign 2_n10674 = 2_n4263 | 2_n8131;
assign 2_n4447 = 2_n5145 & 2_n1247;
assign 2_n10219 = ~(2_n9445 | 2_n651);
assign 2_n10925 = 2_n6577 | 2_n5012;
assign 2_n1621 = 2_n5038 & 2_n2570;
assign 2_n1117 = ~2_n3074;
assign 2_n10341 = ~(2_n10380 ^ 2_n4609);
assign 2_n6033 = 2_n11887 | 2_n8740;
assign 2_n9958 = ~2_n6039;
assign 2_n10509 = 2_n3322 | 2_n9842;
assign 2_n8695 = ~2_n8808;
assign 2_n3004 = ~(2_n223 ^ 2_n4172);
assign 2_n4450 = 2_n1599 & 2_n11816;
assign 2_n9340 = ~(2_n6952 ^ 2_n4592);
assign 2_n1731 = 2_n3747 | 2_n12249;
assign 2_n7278 = ~(2_n7467 ^ 2_n1063);
assign 2_n11834 = ~(2_n812 ^ 2_n11007);
assign 2_n1388 = ~(2_n9261 | 2_n9726);
assign 2_n10092 = ~(2_n11234 | 2_n12522);
assign 2_n8016 = ~(2_n6612 ^ 2_n3069);
assign 2_n2957 = 2_n11887 | 2_n8655;
assign 2_n4595 = 2_n11980 & 2_n3142;
assign 2_n1851 = ~2_n12591;
assign 2_n11498 = 2_n5765 | 2_n795;
assign 2_n9701 = 2_n11796 & 2_n5093;
assign 2_n1004 = ~2_n11208;
assign 2_n7612 = 2_n8026 | 2_n3421;
assign 2_n7566 = 2_n6474 & 2_n10755;
assign 2_n10477 = 2_n12 | 2_n3805;
assign 2_n7501 = ~(2_n5742 ^ 2_n10360);
assign 2_n10411 = 2_n9365 | 2_n3307;
assign 2_n12114 = 2_n8552 | 2_n12535;
assign 2_n3640 = 2_n7038 & 2_n6907;
assign 2_n7373 = ~(2_n4576 | 2_n7365);
assign 2_n6730 = 2_n4504 | 2_n12036;
assign 2_n4997 = ~(2_n3577 ^ 2_n4372);
assign 2_n12132 = 2_n288 & 2_n11386;
assign 2_n11008 = 2_n9693 | 2_n8708;
assign 2_n1807 = ~(2_n3626 ^ 2_n5062);
assign 2_n1256 = 2_n1542 & 2_n9639;
assign 2_n2546 = ~(2_n9677 ^ 2_n4331);
assign 2_n8576 = 2_n9370 | 2_n11430;
assign 2_n3117 = 2_n6407 & 2_n2208;
assign 2_n506 = 2_n6325 & 2_n12504;
assign 2_n11417 = 2_n3746 | 2_n10903;
assign 2_n9500 = 2_n321 & 2_n3426;
assign 2_n7468 = 2_n989 | 2_n7341;
assign 2_n3610 = ~(2_n12047 ^ 2_n4004);
assign 2_n9392 = ~(2_n1959 ^ 2_n5349);
assign 2_n8561 = 2_n10832 & 2_n7421;
assign 2_n8541 = ~2_n8712;
assign 2_n1421 = 2_n236 | 2_n3770;
assign 2_n6289 = ~(2_n3208 ^ 2_n6757);
assign 2_n3803 = ~2_n4004;
assign 2_n5173 = ~2_n5522;
assign 2_n7570 = ~(2_n2318 | 2_n9475);
assign 2_n1141 = ~(2_n2598 | 2_n7576);
assign 2_n8896 = 2_n5530 | 2_n5781;
assign 2_n3684 = 2_n8187 | 2_n6402;
assign 2_n6993 = 2_n7449 | 2_n9280;
assign 2_n11091 = ~(2_n835 ^ 2_n7979);
assign 2_n7163 = ~(2_n4723 ^ 2_n8905);
assign 2_n7822 = 2_n3467 | 2_n11304;
assign 2_n1243 = ~2_n833;
assign 2_n1975 = 2_n6306 & 2_n12452;
assign 2_n11475 = ~2_n1973;
assign 2_n7416 = 2_n3137 | 2_n1711;
assign 2_n4793 = ~2_n12286;
assign 2_n832 = 2_n3920 & 2_n4934;
assign 2_n4612 = 2_n8738 | 2_n4474;
assign 2_n3696 = ~(2_n11971 ^ 2_n10228);
assign 2_n4822 = ~2_n3779;
assign 2_n12202 = 2_n10721 & 2_n8976;
assign 2_n5353 = 2_n9560 & 2_n12439;
assign 2_n8742 = ~(2_n716 ^ 2_n8670);
assign 2_n7694 = 2_n1941 | 2_n995;
assign 2_n11379 = ~2_n9851;
assign 2_n21 = 2_n12363 & 2_n9142;
assign 2_n3527 = 2_n7801 | 2_n6651;
assign 2_n12117 = 2_n10879 | 2_n12843;
assign 2_n3006 = 2_n6364 & 2_n8599;
assign 2_n6710 = 2_n9785 & 2_n574;
assign 2_n1456 = 2_n8428 | 2_n5538;
assign 2_n12758 = 2_n337 | 2_n12329;
assign 2_n10135 = 2_n8583 | 2_n3606;
assign 2_n11646 = ~(2_n12054 ^ 2_n2173);
assign 2_n11166 = 2_n3172 & 2_n7456;
assign 2_n4021 = ~(2_n11700 ^ 2_n11456);
assign 2_n8886 = ~(2_n5466 ^ 2_n4578);
assign 2_n956 = ~(2_n12918 ^ 2_n4606);
assign 2_n191 = ~2_n7862;
assign 2_n2355 = ~(2_n12200 | 2_n6975);
assign 2_n12180 = 2_n752 | 2_n6084;
assign 2_n1981 = 2_n8506 | 2_n2381;
assign 2_n143 = 2_n9250 & 2_n10453;
assign 2_n10876 = 2_n12955 & 2_n873;
assign 2_n6369 = 2_n5305 & 2_n6038;
assign 2_n7567 = 2_n962 | 2_n1047;
assign 2_n10082 = ~2_n1187;
assign 2_n12051 = 2_n8055 | 2_n3802;
assign 2_n6439 = 2_n2612 | 2_n10166;
assign 2_n2376 = ~(2_n9993 ^ 2_n1281);
assign 2_n12338 = ~(2_n2263 ^ 2_n6568);
assign 2_n10828 = ~(2_n2333 ^ 2_n9209);
assign 2_n7536 = 2_n6560 & 2_n3741;
assign 2_n1970 = ~(2_n8663 | 2_n5056);
assign 2_n10544 = ~(2_n12544 ^ 2_n9334);
assign 2_n11568 = ~(2_n6708 ^ 2_n7781);
assign 2_n6758 = 2_n6347 & 2_n9890;
assign 2_n5274 = 2_n7982 & 2_n7184;
assign 2_n2780 = 2_n4343 | 2_n3224;
assign 2_n8894 = 2_n7391 | 2_n4400;
assign 2_n2652 = ~(2_n11120 ^ 2_n280);
assign 2_n3868 = ~2_n1520;
assign 2_n9523 = 2_n3746 | 2_n9971;
assign 2_n8887 = 2_n10992 | 2_n12749;
assign 2_n1841 = ~2_n1511;
assign 2_n10185 = 2_n11671 | 2_n7681;
assign 2_n9205 = 2_n10108 | 2_n3911;
assign 2_n4556 = 2_n5374 & 2_n3182;
assign 2_n7012 = 2_n3127 | 2_n7703;
assign 2_n2769 = ~2_n1156;
assign 2_n760 = ~(2_n5000 ^ 2_n3649);
assign 2_n3205 = 2_n989 | 2_n10419;
assign 2_n9879 = ~(2_n9909 | 2_n5227);
assign 2_n3239 = ~(2_n12023 ^ 2_n7734);
assign 2_n5208 = 2_n619 & 2_n8257;
assign 2_n1224 = 2_n6836 | 2_n2004;
assign 2_n8985 = ~(2_n899 ^ 2_n4424);
assign 2_n8478 = ~2_n479;
assign 2_n10456 = ~(2_n363 ^ 2_n7411);
assign 2_n438 = 2_n8428 | 2_n6455;
assign 2_n9294 = ~(2_n1695 ^ 2_n276);
assign 2_n7504 = 2_n8026 | 2_n9741;
assign 2_n11211 = 2_n3188 | 2_n689;
assign 2_n10361 = 2_n10196 | 2_n9144;
assign 2_n3026 = 2_n726 & 2_n3800;
assign 2_n1922 = 2_n7449 | 2_n4474;
assign 2_n1598 = ~(2_n6201 ^ 2_n1957);
assign 2_n12149 = 2_n6069 | 2_n2586;
assign 2_n1044 = 2_n8583 | 2_n1047;
assign 2_n10450 = ~(2_n6361 ^ 2_n4163);
assign 2_n9985 = ~(2_n6598 ^ 2_n10704);
assign 2_n6917 = ~(2_n689 ^ 2_n12152);
assign 2_n8023 = ~(2_n841 ^ 2_n7242);
assign 2_n51 = 2_n8127 | 2_n1079;
assign 2_n10358 = ~(2_n5646 | 2_n3134);
assign 2_n2280 = ~(2_n11142 ^ 2_n10187);
assign 2_n117 = ~2_n9923;
assign 2_n6694 = ~(2_n5769 ^ 2_n7239);
assign 2_n8093 = 2_n629 & 2_n8432;
assign 2_n4237 = 2_n12237 | 2_n9188;
assign 2_n2294 = ~(2_n9390 ^ 2_n9482);
assign 2_n1518 = 2_n834 & 2_n5431;
assign 2_n2447 = 2_n5575 | 2_n9741;
assign 2_n5821 = ~(2_n9103 ^ 2_n11114);
assign 2_n12492 = ~(2_n8666 ^ 2_n10557);
assign 2_n2719 = ~2_n1624;
assign 2_n5999 = 2_n4366 & 2_n10752;
assign 2_n12283 = 2_n6697 & 2_n12225;
assign 2_n1380 = 2_n8183 | 2_n4720;
assign 2_n10065 = ~2_n774;
assign 2_n9351 = 2_n5945 | 2_n6169;
assign 2_n3181 = 2_n1183 | 2_n8109;
assign 2_n5365 = 2_n6570 & 2_n11756;
assign 2_n9295 = ~(2_n8243 | 2_n2510);
assign 2_n440 = 2_n3796 & 2_n5592;
assign 2_n8683 = ~2_n4307;
assign 2_n6308 = ~(2_n10056 ^ 2_n9809);
assign 2_n255 = 2_n7116 | 2_n10903;
assign 2_n1507 = 2_n9622 & 2_n2782;
assign 2_n9227 = ~(2_n3116 | 2_n9931);
assign 2_n11102 = 2_n7116 | 2_n11410;
assign 2_n12918 = 2_n8187 | 2_n4400;
assign 2_n11815 = ~(2_n2019 | 2_n11218);
assign 2_n4756 = ~(2_n38 ^ 2_n6317);
assign 2_n275 = 2_n2367 | 2_n4527;
assign 2_n11413 = 2_n4059 | 2_n11827;
assign 2_n5552 = ~(2_n10846 ^ 2_n11890);
assign 2_n5357 = 2_n989 | 2_n4775;
assign 2_n1724 = 2_n10108 | 2_n4400;
assign 2_n9206 = ~(2_n9442 ^ 2_n12158);
assign 2_n11254 = 2_n4961 | 2_n231;
assign 2_n11637 = ~2_n4684;
assign 2_n4136 = 2_n4059 | 2_n5497;
assign 2_n10801 = 2_n3632 | 2_n2416;
assign 2_n4457 = 2_n8428 | 2_n7558;
assign 2_n6975 = ~(2_n1586 ^ 2_n4236);
assign 2_n745 = ~(2_n845 ^ 2_n5325);
assign 2_n11825 = 2_n824 | 2_n261;
assign 2_n7977 = 2_n10751 | 2_n4114;
assign 2_n10821 = ~(2_n4124 ^ 2_n1342);
assign 2_n11021 = ~(2_n6004 ^ 2_n7204);
assign 2_n1389 = ~(2_n7194 ^ 2_n3514);
assign 2_n10383 = 2_n813 | 2_n9865;
assign 2_n1029 = ~(2_n3021 ^ 2_n7548);
assign 2_n698 = ~2_n5337;
assign 2_n884 = 2_n5501 & 2_n4792;
assign 2_n1385 = 2_n8279 & 2_n3861;
assign 2_n2827 = 2_n8336 & 2_n6703;
assign 2_n10436 = 2_n1043 & 2_n11532;
assign 2_n2947 = 2_n9878 | 2_n3924;
assign 2_n3002 = 2_n1795 | 2_n1748;
assign 2_n1091 = 2_n8269 & 2_n5528;
assign 2_n12251 = 2_n7283 | 2_n1162;
assign 2_n4070 = 2_n9441 & 2_n7837;
assign 2_n7596 = ~(2_n3829 ^ 2_n8150);
assign 2_n6167 = 2_n10075 & 2_n4837;
assign 2_n8975 = ~(2_n6414 ^ 2_n4749);
assign 2_n1200 = ~2_n6535;
assign 2_n9309 = 2_n12429 | 2_n6135;
assign 2_n2873 = 2_n11641 & 2_n12379;
assign 2_n12258 = ~(2_n7143 ^ 2_n1997);
assign 2_n6340 = ~2_n8564;
assign 2_n8976 = 2_n3215 | 2_n2682;
assign 2_n2812 = 2_n6859 & 2_n8559;
assign 2_n1786 = ~(2_n1724 ^ 2_n3122);
assign 2_n1289 = ~(2_n2292 ^ 2_n9276);
assign 2_n4651 = 2_n1421 & 2_n1254;
assign 2_n12469 = ~(2_n4167 ^ 2_n5007);
assign 2_n9430 = 2_n3405 | 2_n9833;
assign 2_n2820 = ~(2_n10238 ^ 2_n3850);
assign 2_n1191 = ~(2_n10771 ^ 2_n9904);
assign 2_n6263 = ~(2_n10745 ^ 2_n3082);
assign 2_n161 = 2_n5575 | 2_n12899;
assign 2_n12321 = 2_n614 & 2_n4443;
assign 2_n4512 = 2_n12361 | 2_n11122;
assign 2_n8484 = ~(2_n10 ^ 2_n11277);
assign 2_n10842 = 2_n636 | 2_n3924;
assign 2_n9738 = 2_n4324 & 2_n1085;
assign 2_n8226 = 2_n7606 | 2_n9822;
assign 2_n1626 = ~(2_n12483 | 2_n3830);
assign 2_n8200 = ~(2_n8806 | 2_n110);
assign 2_n9975 = ~(2_n5709 | 2_n886);
assign 2_n8752 = 2_n1937 | 2_n6455;
assign 2_n7676 = ~(2_n4439 ^ 2_n9375);
assign 2_n11213 = ~(2_n3762 ^ 2_n9060);
assign 2_n12634 = ~(2_n9648 ^ 2_n5802);
assign 2_n2863 = ~(2_n5607 | 2_n7712);
assign 2_n10401 = 2_n6616 & 2_n10578;
assign 2_n8697 = 2_n6265 | 2_n8041;
assign 2_n8186 = 2_n11588 & 2_n5476;
assign 2_n4131 = ~(2_n2233 ^ 2_n1184);
assign 2_n8299 = 2_n12853 | 2_n530;
assign 2_n3670 = ~2_n6948;
assign 2_n1287 = 2_n12237 | 2_n4818;
assign 2_n7926 = ~(2_n3116 ^ 2_n4061);
assign 2_n4249 = ~2_n1576;
assign 2_n3772 = 2_n6530 | 2_n3167;
assign 2_n3338 = 2_n7994 | 2_n7450;
assign 2_n10079 = 2_n8187 | 2_n5497;
assign 2_n4754 = 2_n9510 | 2_n11586;
assign 2_n12352 = ~(2_n6268 | 2_n2420);
assign 2_n9716 = 2_n8406 & 2_n2607;
assign 2_n11924 = ~2_n7097;
assign 2_n6278 = 2_n6066 & 2_n5292;
assign 2_n11206 = ~(2_n1012 ^ 2_n5547);
assign 2_n4400 = ~2_n11407;
assign 2_n1703 = 2_n11310 | 2_n6964;
assign 2_n12095 = ~(2_n5621 | 2_n4075);
assign 2_n10016 = ~(2_n8908 ^ 2_n3736);
assign 2_n9748 = 2_n994 | 2_n4242;
assign 2_n3766 = 2_n9748 | 2_n10395;
assign 2_n8277 = ~2_n9319;
assign 2_n10335 = 2_n10975 & 2_n2152;
assign 2_n9634 = 2_n5279 | 2_n12258;
assign 2_n464 = 2_n7396 & 2_n5885;
assign 2_n8071 = 2_n2215 & 2_n6729;
assign 2_n12236 = ~2_n11545;
assign 2_n3121 = ~(2_n11177 ^ 2_n7836);
assign 2_n505 = 2_n12853 | 2_n8655;
assign 2_n5465 = 2_n12742 | 2_n11768;
assign 2_n6663 = 2_n5355 | 2_n9397;
assign 2_n6915 = ~(2_n4510 ^ 2_n6410);
assign 2_n6579 = 2_n10142 | 2_n7881;
assign 2_n6302 = ~2_n12055;
assign 2_n6064 = 2_n11211 & 2_n3438;
assign 2_n1320 = 2_n7083 & 2_n672;
assign 2_n10329 = 2_n5279 & 2_n12258;
assign 2_n11807 = ~(2_n1542 ^ 2_n5317);
assign 2_n7944 = 2_n5923 & 2_n412;
assign 2_n8785 = 2_n10374 | 2_n3898;
assign 2_n12005 = ~(2_n9737 ^ 2_n3263);
assign 2_n6420 = ~(2_n1628 ^ 2_n417);
assign 2_n3061 = ~(2_n1312 ^ 2_n2518);
assign 2_n9103 = ~(2_n317 ^ 2_n4065);
assign 2_n4330 = ~(2_n3362 | 2_n2178);
assign 2_n10373 = ~2_n6086;
assign 2_n6241 = 2_n7133 | 2_n2395;
assign 2_n12650 = ~(2_n5899 ^ 2_n3201);
assign 2_n9621 = ~(2_n12865 ^ 2_n6627);
assign 2_n11084 = ~(2_n1371 | 2_n6392);
assign 2_n7392 = 2_n1908 & 2_n315;
assign 2_n9519 = 2_n3127 | 2_n1546;
assign 2_n8297 = ~2_n10535;
assign 2_n2946 = 2_n3603 | 2_n2715;
assign 2_n880 = ~2_n8719;
assign 2_n11667 = ~(2_n8474 | 2_n3774);
assign 2_n3030 = 2_n11026 | 2_n12120;
assign 2_n5483 = ~(2_n8668 ^ 2_n2206);
assign 2_n11641 = ~(2_n9405 ^ 2_n1794);
assign 2_n3079 = ~2_n7074;
assign 2_n5916 = 2_n1777 & 2_n304;
assign 2_n9478 = ~(2_n2535 ^ 2_n11416);
assign 2_n10697 = ~(2_n7612 ^ 2_n10080);
assign 2_n3681 = 2_n11550 & 2_n7051;
assign 2_n1818 = ~(2_n1774 ^ 2_n3777);
assign 2_n4885 = 2_n10656 | 2_n7948;
assign 2_n10164 = ~(2_n7396 ^ 2_n1995);
assign 2_n12310 = 2_n3105 | 2_n358;
assign 2_n310 = ~2_n1979;
assign 2_n7798 = 2_n3742 & 2_n390;
assign 2_n12506 = 2_n8049 & 2_n12510;
assign 2_n6919 = ~(2_n11879 | 2_n11392);
assign 2_n6148 = ~(2_n1608 ^ 2_n9668);
assign 2_n9086 = 2_n8169 & 2_n6633;
assign 2_n1767 = ~(2_n1457 ^ 2_n8297);
assign 2_n4505 = ~(2_n4210 ^ 2_n12769);
assign 2_n7968 = ~2_n6289;
assign 2_n3975 = ~(2_n8454 ^ 2_n5734);
assign 2_n2283 = ~(2_n12612 ^ 2_n5537);
assign 2_n12763 = ~(2_n7630 | 2_n5736);
assign 2_n9839 = ~(2_n6234 ^ 2_n11982);
assign 2_n1643 = ~2_n7454;
assign 2_n10857 = 2_n10902 & 2_n1393;
assign 2_n4144 = 2_n9370 | 2_n1738;
assign 2_n9155 = 2_n11026 | 2_n7506;
assign 2_n10855 = 2_n11076 | 2_n7067;
assign 2_n5018 = ~2_n5976;
assign 2_n3867 = ~2_n3858;
assign 2_n7834 = ~2_n11289;
assign 2_n6426 = 2_n10835 | 2_n8830;
assign 2_n5033 = ~(2_n9054 ^ 2_n1187);
assign 2_n489 = ~(2_n5542 | 2_n7234);
assign 2_n7353 = ~(2_n3510 | 2_n7366);
assign 2_n5909 = 2_n4134 & 2_n1943;
assign 2_n3882 = ~(2_n9429 | 2_n7092);
assign 2_n11143 = ~(2_n6246 ^ 2_n10345);
assign 2_n1719 = 2_n12853 | 2_n4913;
assign 2_n8797 = 2_n5730 & 2_n10407;
assign 2_n1511 = 2_n11474 | 2_n9371;
assign 2_n1028 = ~(2_n11335 | 2_n6518);
assign 2_n9269 = 2_n12867 & 2_n3434;
assign 2_n9011 = ~(2_n8682 | 2_n1525);
assign 2_n4107 = 2_n1183 | 2_n1932;
assign 2_n4557 = ~2_n3776;
assign 2_n10121 = 2_n11682 | 2_n12092;
assign 2_n4663 = ~(2_n4716 ^ 2_n7053);
assign 2_n10572 = 2_n5066 | 2_n3226;
assign 2_n9864 = ~(2_n1074 | 2_n5426);
assign 2_n11978 = ~2_n3877;
assign 2_n10967 = ~(2_n5491 ^ 2_n3664);
assign 2_n7054 = 2_n10108 | 2_n10066;
assign 2_n11443 = 2_n5530 | 2_n8259;
assign 2_n3717 = ~2_n3565;
assign 2_n8948 = ~(2_n6122 ^ 2_n189);
assign 2_n504 = 2_n11958 | 2_n3356;
assign 2_n11055 = 2_n7862 & 2_n2879;
assign 2_n4159 = ~(2_n4766 ^ 2_n3635);
assign 2_n5295 = ~(2_n7251 ^ 2_n4264);
assign 2_n1552 = ~(2_n10046 ^ 2_n6927);
assign 2_n7228 = 2_n10104 | 2_n10498;
assign 2_n5287 = 2_n10269 | 2_n3308;
assign 2_n12832 = ~(2_n905 | 2_n11505);
assign 2_n6372 = ~(2_n9708 ^ 2_n4822);
assign 2_n9352 = ~2_n4948;
assign 2_n11651 = ~(2_n1611 ^ 2_n11337);
assign 2_n6885 = ~2_n11373;
assign 2_n2370 = ~(2_n2244 ^ 2_n5697);
assign 2_n1897 = 2_n11890 | 2_n4291;
assign 2_n7400 = 2_n12361 | 2_n3468;
assign 2_n5585 = 2_n5889 | 2_n802;
assign 2_n3895 = 2_n752 | 2_n1413;
assign 2_n8734 = ~(2_n8124 ^ 2_n3270);
assign 2_n5747 = 2_n12565 | 2_n903;
assign 2_n12358 = ~(2_n3988 ^ 2_n11105);
assign 2_n11265 = 2_n8738 | 2_n795;
assign 2_n5835 = ~(2_n1017 | 2_n4853);
assign 2_n3257 = 2_n8336 & 2_n7500;
assign 2_n2267 = 2_n11254 & 2_n7847;
assign 2_n12140 = ~(2_n11462 ^ 2_n5398);
assign 2_n5577 = 2_n10641 & 2_n3867;
assign 2_n6079 = ~(2_n11451 ^ 2_n6853);
assign 2_n4564 = 2_n7495 | 2_n12843;
assign 2_n455 = 2_n8752 | 2_n1918;
assign 2_n10350 = ~2_n2365;
assign 2_n5419 = ~2_n7304;
assign 2_n4029 = 2_n4380 | 2_n5245;
assign 2_n5795 = ~(2_n12671 ^ 2_n1615);
assign 2_n12151 = 2_n12136 | 2_n9779;
assign 2_n12374 = ~(2_n9745 ^ 2_n3112);
assign 2_n12456 = 2_n12503 | 2_n4875;
assign 2_n11551 = 2_n12774 | 2_n2423;
assign 2_n9936 = ~(2_n6367 | 2_n987);
assign 2_n2779 = ~(2_n4301 | 2_n2204);
assign 2_n12652 = 2_n12839 & 2_n1279;
assign 2_n12731 = 2_n11754 | 2_n3073;
assign 2_n10513 = 2_n6373 | 2_n8285;
assign 2_n8089 = 2_n7756 & 2_n4681;
assign 2_n11552 = ~2_n5767;
assign 2_n7616 = ~(2_n9035 ^ 2_n4616);
assign 2_n11395 = ~(2_n11720 ^ 2_n11089);
assign 2_n9863 = ~(2_n9247 ^ 2_n9033);
assign 2_n2967 = ~(2_n1612 | 2_n4673);
assign 2_n2772 = 2_n12245 | 2_n300;
assign 2_n2293 = 2_n11928 | 2_n11308;
assign 2_n11294 = ~2_n7658;
assign 2_n6780 = 2_n8854 | 2_n1035;
assign 2_n6046 = 2_n12739 & 2_n3108;
assign 2_n4951 = ~(2_n5463 | 2_n12693);
assign 2_n718 = 2_n7074 & 2_n4105;
assign 2_n1842 = 2_n6625 | 2_n12959;
assign 2_n12429 = 2_n7176 & 2_n506;
assign 2_n5438 = 2_n3127 | 2_n1851;
assign 2_n8371 = ~2_n391;
assign 2_n11312 = ~(2_n3416 ^ 2_n4687);
assign 2_n6036 = ~2_n7796;
assign 2_n1720 = ~2_n12693;
assign 2_n12933 = 2_n7173 | 2_n8125;
assign 2_n8824 = ~(2_n3405 ^ 2_n10106);
assign 2_n11494 = ~2_n6338;
assign 2_n2438 = ~(2_n1124 ^ 2_n8110);
assign 2_n5959 = 2_n5355 | 2_n510;
assign 2_n2579 = ~2_n11267;
assign 2_n1614 = ~(2_n10735 ^ 2_n4091);
assign 2_n5309 = ~(2_n3628 ^ 2_n894);
assign 2_n8989 = ~(2_n862 ^ 2_n2668);
assign 2_n5366 = 2_n1941 | 2_n2815;
assign 2_n10718 = 2_n12214 & 2_n4423;
assign 2_n11624 = 2_n6718 | 2_n9521;
assign 2_n8620 = 2_n12009 | 2_n788;
assign 2_n12162 = ~(2_n5749 ^ 2_n8809);
assign 2_n11492 = 2_n8294 & 2_n6316;
assign 2_n5403 = ~(2_n1412 ^ 2_n12957);
assign 2_n4462 = ~(2_n11824 ^ 2_n1545);
assign 2_n10094 = 2_n754 | 2_n624;
assign 2_n3931 = ~(2_n10215 ^ 2_n4848);
assign 2_n6137 = 2_n191 | 2_n9589;
assign 2_n6319 = 2_n6003 & 2_n11614;
assign 2_n4619 = ~(2_n5758 ^ 2_n8210);
assign 2_n8995 = ~(2_n8972 ^ 2_n2667);
assign 2_n9410 = 2_n11879 & 2_n11392;
assign 2_n2965 = ~(2_n11532 ^ 2_n1195);
assign 2_n8327 = 2_n343 | 2_n7278;
assign 2_n3568 = ~(2_n11053 ^ 2_n5745);
assign 2_n8022 = ~(2_n1803 ^ 2_n6421);
assign 2_n9358 = ~(2_n11723 ^ 2_n8487);
assign 2_n1229 = 2_n10545 & 2_n7733;
assign 2_n9218 = ~2_n669;
assign 2_n3811 = ~(2_n1707 ^ 2_n700);
assign 2_n8624 = ~2_n1132;
assign 2_n4071 = 2_n10698 & 2_n7208;
assign 2_n11934 = 2_n12814 & 2_n8431;
assign 2_n12621 = ~2_n1410;
assign 2_n10109 = 2_n10714 | 2_n43;
assign 2_n2898 = ~2_n860;
assign 2_n3015 = 2_n5575 | 2_n6084;
assign 2_n7062 = ~(2_n1569 ^ 2_n7211);
assign 2_n3969 = ~(2_n11042 | 2_n6350);
assign 2_n3033 = 2_n9286 | 2_n2889;
assign 2_n12370 = 2_n12393 | 2_n1463;
assign 2_n11835 = ~(2_n6097 ^ 2_n4496);
assign 2_n4446 = 2_n11923 | 2_n1476;
assign 2_n649 = 2_n191 | 2_n10066;
assign 2_n11065 = 2_n1699 | 2_n12754;
assign 2_n3829 = 2_n9003 & 2_n7006;
assign 2_n8123 = 2_n2099 | 2_n2259;
assign 2_n11259 = 2_n8870 | 2_n12080;
assign 2_n4723 = 2_n8870 | 2_n9586;
assign 2_n4407 = 2_n6720 & 2_n7516;
assign 2_n9095 = ~(2_n656 ^ 2_n3516);
assign 2_n3400 = ~(2_n2183 | 2_n5920);
assign 2_n7901 = 2_n1230 & 2_n811;
assign 2_n388 = ~2_n3646;
assign 2_n173 = 2_n11222 & 2_n10848;
assign 2_n1438 = 2_n3127 | 2_n3911;
assign 2_n7866 = ~(2_n3055 ^ 2_n10950);
assign 2_n11260 = ~(2_n5632 ^ 2_n6483);
assign 2_n3884 = ~2_n9858;
assign 2_n10863 = ~(2_n6543 ^ 2_n5480);
assign 2_n2853 = 2_n8552 | 2_n8740;
assign 2_n9315 = ~2_n11499;
assign 2_n5535 = ~(2_n9748 ^ 2_n10395);
assign 2_n1010 = ~(2_n11088 ^ 2_n9952);
assign 2_n11629 = ~(2_n10658 ^ 2_n10946);
assign 2_n4776 = ~(2_n6423 ^ 2_n1125);
assign 2_n8938 = ~(2_n4446 ^ 2_n6647);
assign 2_n1848 = 2_n7564 | 2_n1363;
assign 2_n5020 = 2_n6470 | 2_n7392;
assign 2_n6548 = 2_n11691 & 2_n8511;
assign 2_n2570 = 2_n4831 & 2_n426;
assign 2_n10447 = ~(2_n7762 | 2_n8302);
assign 2_n1451 = 2_n3926 & 2_n10474;
assign 2_n11883 = 2_n3088 | 2_n8080;
assign 2_n4334 = ~(2_n2111 ^ 2_n7631);
assign 2_n5087 = 2_n10142 | 2_n5851;
assign 2_n1532 = 2_n9652 & 2_n9798;
assign 2_n1349 = 2_n9621 & 2_n1490;
assign 2_n3199 = ~2_n10191;
assign 2_n10379 = 2_n8738 | 2_n9144;
assign 2_n916 = ~2_n12553;
assign 2_n2139 = ~2_n1451;
assign 2_n6883 = 2_n6741 | 2_n3136;
assign 2_n6739 = 2_n6426 & 2_n11009;
assign 2_n8909 = ~2_n4883;
assign 2_n3080 = ~2_n7977;
assign 2_n66 = ~(2_n12263 ^ 2_n3569);
assign 2_n6888 = 2_n7322 | 2_n256;
assign 2_n12035 = ~(2_n9117 ^ 2_n3266);
assign 2_n7710 = ~2_n3804;
assign 2_n10177 = ~(2_n1923 | 2_n6640);
assign 2_n2122 = ~2_n8356;
assign 2_n2788 = 2_n5413 & 2_n10170;
assign 2_n1186 = 2_n7151 | 2_n7714;
assign 2_n601 = ~(2_n7488 ^ 2_n8876);
assign 2_n5390 = ~(2_n6686 ^ 2_n7599);
assign 2_n3755 = 2_n6644 | 2_n2461;
assign 2_n4244 = 2_n8026 | 2_n184;
assign 2_n6382 = ~2_n1324;
assign 2_n9236 = 2_n12614 & 2_n1022;
assign 2_n8736 = 2_n5575 | 2_n9971;
assign 2_n4920 = 2_n10835 | 2_n9521;
assign 2_n6961 = ~(2_n4076 ^ 2_n10213);
assign 2_n9543 = 2_n6868 | 2_n793;
assign 2_n12385 = ~2_n2350;
assign 2_n7225 = ~(2_n9336 | 2_n11463);
assign 2_n6680 = 2_n12223 & 2_n7114;
assign 2_n12019 = 2_n12183 | 2_n10177;
assign 2_n6850 = ~(2_n2664 | 2_n7797);
assign 2_n6147 = 2_n4387 | 2_n4162;
assign 2_n5720 = ~(2_n6110 ^ 2_n4199);
assign 2_n11480 = 2_n9836 & 2_n8081;
assign 2_n5371 = 2_n7495 | 2_n10066;
assign 2_n3283 = ~(2_n4322 ^ 2_n512);
assign 2_n6386 = 2_n10744 | 2_n2240;
assign 2_n5378 = 2_n1003 | 2_n6517;
assign 2_n1499 = ~(2_n9752 ^ 2_n7238);
assign 2_n9 = ~(2_n12538 | 2_n10690);
assign 2_n544 = ~(2_n2249 ^ 2_n9983);
assign 2_n4353 = ~(2_n11356 ^ 2_n5342);
assign 2_n12686 = ~2_n7610;
assign 2_n3736 = 2_n8959 | 2_n3421;
assign 2_n9021 = 2_n10018 & 2_n10021;
assign 2_n11430 = ~2_n12000;
assign 2_n1263 = 2_n1679 & 2_n10359;
assign 2_n6979 = 2_n289 | 2_n11772;
assign 2_n805 = 2_n9335 & 2_n11031;
assign 2_n9823 = ~(2_n10195 | 2_n3161);
assign 2_n235 = ~(2_n4121 ^ 2_n11975);
assign 2_n11386 = 2_n8583 | 2_n1509;
assign 2_n4701 = ~(2_n8030 ^ 2_n8060);
assign 2_n8727 = 2_n9504 | 2_n11910;
assign 2_n7293 = ~2_n5898;
assign 2_n9347 = 2_n12218 & 2_n2632;
assign 2_n3228 = ~(2_n6624 | 2_n10834);
assign 2_n3515 = ~(2_n5577 ^ 2_n3204);
assign 2_n4576 = 2_n5530 | 2_n12124;
assign 2_n2183 = 2_n10004 ^ 2_n6289;
assign 2_n6821 = ~(2_n6461 ^ 2_n3211);
assign 2_n12584 = 2_n81 & 2_n12343;
assign 2_n1898 = 2_n2003 & 2_n12762;
assign 2_n7748 = 2_n4059 | 2_n2358;
assign 2_n12761 = 2_n989 | 2_n5851;
assign 2_n3105 = 2_n12361 | 2_n9741;
assign 2_n7595 = ~(2_n12114 ^ 2_n944);
assign 2_n11470 = 2_n4120 | 2_n2805;
assign 2_n4270 = ~(2_n9757 ^ 2_n5806);
assign 2_n4129 = 2_n7941 | 2_n9113;
assign 2_n7164 = ~(2_n5981 ^ 2_n282);
assign 2_n6164 = 2_n1073 & 2_n6790;
assign 2_n10770 = 2_n5860 & 2_n10848;
assign 2_n3808 = ~2_n7405;
assign 2_n12567 = 2_n2286 | 2_n7581;
assign 2_n5736 = 2_n7544 & 2_n7228;
assign 2_n11944 = ~2_n12811;
assign 2_n8959 = ~2_n7436;
assign 2_n1466 = ~(2_n1486 ^ 2_n4221);
assign 2_n7178 = 2_n6698 & 2_n2158;
assign 2_n4172 = ~(2_n1330 ^ 2_n106);
assign 2_n486 = ~2_n10023;
assign 2_n4161 = 2_n10750 | 2_n12883;
assign 2_n1959 = ~(2_n12887 | 2_n539);
assign 2_n9555 = ~(2_n11284 ^ 2_n5626);
assign 2_n8482 = ~(2_n3065 ^ 2_n7032);
assign 2_n7175 = ~(2_n8776 ^ 2_n123);
assign 2_n8404 = 2_n3096 | 2_n11896;
assign 2_n10354 = 2_n12119 | 2_n7928;
assign 2_n12054 = ~(2_n10809 ^ 2_n11107);
assign 2_n11162 = 2_n6681 | 2_n10894;
assign 2_n11219 = ~(2_n815 ^ 2_n11075);
assign 2_n1372 = 2_n5066 & 2_n3226;
assign 2_n9318 = 2_n3664 | 2_n6712;
assign 2_n4709 = ~(2_n2215 ^ 2_n6729);
assign 2_n3058 = ~2_n4838;
assign 2_n12014 = ~(2_n2805 ^ 2_n5521);
assign 2_n10991 = ~(2_n1361 | 2_n8577);
assign 2_n6654 = 2_n8870 | 2_n7382;
assign 2_n2689 = ~2_n1479;
assign 2_n8165 = 2_n23 & 2_n7844;
assign 2_n825 = ~(2_n11745 | 2_n2578);
assign 2_n3229 = ~2_n5819;
assign 2_n3391 = ~(2_n9281 ^ 2_n8563);
assign 2_n1971 = ~(2_n7713 ^ 2_n9343);
assign 2_n4964 = 2_n10975 | 2_n2152;
assign 2_n4674 = ~2_n4499;
assign 2_n7818 = ~(2_n705 ^ 2_n8192);
assign 2_n10480 = 2_n12361 | 2_n6169;
assign 2_n3354 = ~(2_n933 ^ 2_n12666);
assign 2_n9932 = ~(2_n6222 ^ 2_n9902);
assign 2_n4802 = ~2_n1880;
assign 2_n2565 = ~(2_n396 ^ 2_n8802);
assign 2_n8408 = ~(2_n11489 ^ 2_n1403);
assign 2_n7943 = ~2_n12700;
assign 2_n9169 = 2_n1128 & 2_n6110;
assign 2_n7482 = ~(2_n2382 ^ 2_n6633);
assign 2_n8090 = ~2_n8799;
assign 2_n7887 = ~(2_n3804 ^ 2_n3531);
assign 2_n4676 = 2_n8738 | 2_n3606;
assign 2_n11721 = ~(2_n3327 | 2_n11046);
assign 2_n10982 = ~2_n12003;
assign 2_n243 = 2_n6146 | 2_n6749;
assign 2_n12856 = 2_n9370 | 2_n1455;
assign 2_n11547 = 2_n10157 | 2_n8643;
assign 2_n2790 = ~2_n5888;
assign 2_n2922 = 2_n7012 & 2_n2026;
assign 2_n10957 = 2_n9193 | 2_n6351;
assign 2_n12097 = ~(2_n3209 ^ 2_n8681);
assign 2_n78 = 2_n5530 | 2_n12080;
assign 2_n12733 = 2_n11222 & 2_n405;
assign 2_n770 = 2_n6348 | 2_n10175;
assign 2_n1053 = 2_n11719 | 2_n12843;
assign 2_n9536 = ~2_n10734;
assign 2_n3689 = ~(2_n3966 ^ 2_n11977);
assign 2_n1266 = 2_n6577 | 2_n2815;
assign 2_n12693 = 2_n508 & 2_n8530;
assign 2_n1712 = ~(2_n4542 ^ 2_n5403);
assign 2_n8569 = 2_n12127 & 2_n3081;
assign 2_n10773 = ~2_n8900;
assign 2_n7766 = ~(2_n1787 ^ 2_n7591);
assign 2_n11249 = 2_n1539 | 2_n1455;
assign 2_n4206 = 2_n7283 | 2_n7424;
assign 2_n2296 = ~(2_n8353 ^ 2_n1922);
assign 2_n7108 = 2_n6650 | 2_n5386;
assign 2_n10359 = ~(2_n3182 ^ 2_n4082);
assign 2_n8098 = 2_n6111 | 2_n212;
assign 2_n1485 = ~(2_n10313 ^ 2_n6603);
assign 2_n10910 = ~2_n82;
assign 2_n7465 = 2_n8026 | 2_n11775;
assign 2_n1736 = 2_n646 & 2_n494;
assign 2_n7370 = 2_n4204 | 2_n5028;
assign 2_n6023 = ~(2_n12884 ^ 2_n4139);
assign 2_n8847 = 2_n12119 | 2_n2964;
assign 2_n5462 = ~2_n3284;
assign 2_n6291 = 2_n4811 & 2_n8090;
assign 2_n8138 = ~(2_n8460 ^ 2_n5610);
assign 2_n5533 = ~(2_n11935 ^ 2_n10821);
assign 2_n8659 = 2_n4059 | 2_n4775;
assign 2_n9510 = 2_n4498 | 2_n11827;
assign 2_n11292 = ~2_n3206;
assign 2_n9335 = ~2_n11188;
assign 2_n5831 = ~(2_n8704 ^ 2_n11689);
assign 2_n10808 = 2_n12853 | 2_n7928;
assign 2_n3682 = ~2_n5284;
assign 2_n5880 = 2_n8587 & 2_n10206;
assign 2_n6702 = ~(2_n8320 ^ 2_n6588);
assign 2_n2804 = ~2_n742;
assign 2_n9947 = ~(2_n9620 ^ 2_n9238);
assign 2_n2932 = ~(2_n1356 ^ 2_n10540);
assign 2_n6533 = ~(2_n11997 ^ 2_n930);
assign 2_n8680 = ~(2_n6073 ^ 2_n8947);
assign 2_n5350 = 2_n11841 & 2_n3002;
assign 2_n10974 = 2_n4628 | 2_n12535;
assign 2_n8945 = 2_n1051 | 2_n9741;
assign 2_n4686 = 2_n1027 ^ 2_n3950;
assign 2_n10157 = ~2_n3992;
assign 2_n7029 = ~(2_n10878 | 2_n5623);
assign 2_n10559 = ~(2_n2397 ^ 2_n12403);
assign 2_n10587 = 2_n8552 | 2_n7382;
assign 2_n6701 = 2_n11445 | 2_n247;
assign 2_n985 = ~(2_n1266 ^ 2_n6324);
assign 2_n2672 = 2_n8552 | 2_n8109;
assign 2_n7426 = ~(2_n5263 ^ 2_n3657);
assign 2_n365 = 2_n1699 | 2_n10854;
assign 2_n10403 = 2_n1594 & 2_n10964;
assign 2_n5486 = 2_n8583 | 2_n9521;
assign 2_n4445 = ~(2_n3988 | 2_n5039);
assign 2_n8237 = 2_n10118 & 2_n5887;
assign 2_n1854 = 2_n11226 | 2_n2658;
assign 2_n3356 = ~2_n8236;
assign 2_n1319 = ~(2_n4718 | 2_n3634);
assign 2_n4278 = ~(2_n7643 | 2_n913);
assign 2_n7275 = 2_n637 & 2_n5996;
assign 2_n8878 = 2_n10434 & 2_n9894;
assign 2_n6024 = 2_n197 & 2_n8330;
assign 2_n6398 = 2_n3713 | 2_n3227;
assign 2_n1323 = ~(2_n6865 | 2_n9059);
assign 2_n11119 = ~2_n6353;
assign 2_n6117 = 2_n1856 | 2_n3748;
assign 2_n6581 = 2_n8354 | 2_n6513;
assign 2_n1177 = ~(2_n12471 ^ 2_n535);
assign 2_n11035 = ~(2_n12524 | 2_n8898);
assign 2_n7067 = 2_n762 & 2_n6312;
assign 2_n7301 = 2_n2251 & 2_n4277;
assign 2_n2196 = ~(2_n7897 | 2_n4918);
assign 2_n3124 = ~(2_n12267 ^ 2_n7399);
assign 2_n9753 = 2_n9279 & 2_n10331;
assign 2_n5844 = 2_n11182 | 2_n4200;
assign 2_n600 = ~(2_n3906 ^ 2_n11203);
assign 2_n7222 = ~(2_n1536 ^ 2_n12651);
assign 2_n11284 = ~(2_n1347 ^ 2_n7216);
assign 2_n5517 = ~(2_n9467 ^ 2_n9312);
assign 2_n4856 = 2_n5575 | 2_n8768;
assign 2_n1639 = 2_n8428 | 2_n12816;
assign 2_n4348 = ~2_n707;
assign 2_n8844 = 2_n2226 & 2_n2522;
assign 2_n9586 = ~2_n11967;
assign 2_n10711 = ~(2_n10724 ^ 2_n10581);
assign 2_n9887 = 2_n6977 | 2_n9741;
assign 2_n4919 = 2_n2930 & 2_n4901;
assign 2_n5251 = 2_n636 | 2_n3224;
assign 2_n2707 = 2_n12263 & 2_n9203;
assign 2_n10705 = ~(2_n582 ^ 2_n11014);
assign 2_n2796 = ~(2_n3976 ^ 2_n10429);
assign 2_n8211 = ~2_n7277;
assign 2_n6182 = ~2_n1082;
assign 2_n2320 = ~(2_n4191 ^ 2_n6555);
assign 2_n10693 = ~(2_n3396 ^ 2_n12700);
assign 2_n10606 = ~2_n10171;
assign 2_n12088 = ~(2_n6894 | 2_n7105);
assign 2_n12628 = 2_n1842 & 2_n10943;
assign 2_n12058 = ~(2_n6514 ^ 2_n5373);
assign 2_n11246 = ~(2_n4597 ^ 2_n394);
assign 2_n458 = ~(2_n1873 ^ 2_n11223);
assign 2_n8751 = 2_n10835 | 2_n1739;
assign 2_n1428 = ~(2_n2274 ^ 2_n11858);
assign 2_n6226 = 2_n7243 & 2_n2460;
assign 2_n3869 = ~(2_n8097 ^ 2_n4520);
assign 2_n10192 = ~(2_n3888 ^ 2_n10029);
assign 2_n12689 = 2_n116 & 2_n5826;
assign 2_n7540 = 2_n9656 & 2_n12411;
assign 2_n10259 = 2_n1951 & 2_n11244;
assign 2_n5099 = ~(2_n9461 | 2_n6363);
assign 2_n9962 = ~(2_n5963 | 2_n4102);
assign 2_n112 = 2_n9321 ^ 2_n3824;
assign 2_n12943 = ~(2_n8545 ^ 2_n4824);
assign 2_n11973 = 2_n9389 | 2_n11430;
assign 2_n4469 = ~(2_n1949 ^ 2_n12487);
assign 2_n9405 = ~(2_n8949 ^ 2_n6724);
assign 2_n11263 = 2_n8322 & 2_n6737;
assign 2_n12887 = ~(2_n6751 | 2_n3519);
assign 2_n1112 = 2_n1051 | 2_n7425;
assign 2_n4675 = 2_n2613 | 2_n3826;
assign 2_n1118 = ~(2_n4001 ^ 2_n592);
assign 2_n2398 = 2_n4628 | 2_n6513;
assign 2_n5304 = ~(2_n6728 ^ 2_n3827);
assign 2_n6938 = ~(2_n2991 ^ 2_n8769);
assign 2_n540 = ~(2_n2561 | 2_n6572);
assign 2_n3100 = ~(2_n9230 ^ 2_n8689);
assign 2_n6834 = ~(2_n4437 ^ 2_n5220);
assign 2_n1379 = ~(2_n1127 | 2_n11848);
assign 2_n482 = 2_n10697 & 2_n4968;
assign 2_n9613 = ~(2_n3792 ^ 2_n1244);
assign 2_n5555 = ~(2_n7009 ^ 2_n7664);
assign 2_n12912 = 2_n11887 | 2_n12080;
assign 2_n6520 = ~(2_n5334 ^ 2_n4884);
assign 2_n11804 = ~(2_n5335 | 2_n9207);
assign 2_n3046 = ~(2_n11960 ^ 2_n3273);
assign 2_n2414 = 2_n3145 | 2_n1267;
assign 2_n2584 = ~(2_n7983 ^ 2_n2334);
assign 2_n5109 = ~(2_n4315 ^ 2_n8832);
assign 2_n6037 = ~(2_n10203 | 2_n7219);
assign 2_n8840 = ~(2_n5988 ^ 2_n6856);
assign 2_n6341 = ~(2_n6874 | 2_n10455);
assign 2_n2146 = ~(2_n8635 ^ 2_n2698);
assign 2_n8942 = ~(2_n35 ^ 2_n9110);
assign 2_n9502 = ~(2_n9432 ^ 2_n7226);
assign 2_n7781 = ~(2_n8319 ^ 2_n8044);
assign 2_n2445 = ~2_n5371;
assign 2_n11216 = ~(2_n7230 ^ 2_n9154);
assign 2_n10247 = ~(2_n8092 | 2_n5459);
assign 2_n12111 = ~(2_n7708 ^ 2_n2758);
assign 2_n4384 = 2_n1288 | 2_n2868;
assign 2_n10486 = 2_n2854 & 2_n1961;
assign 2_n9210 = ~2_n292;
assign 2_n9622 = 2_n11228 | 2_n8573;
assign 2_n6560 = 2_n5765 | 2_n4642;
assign 2_n4024 = ~(2_n3928 ^ 2_n9075);
assign 2_n5859 = ~(2_n8254 ^ 2_n6490);
assign 2_n4058 = ~(2_n2975 ^ 2_n10901);
assign 2_n1468 = ~(2_n3329 | 2_n9053);
assign 2_n2861 = 2_n7965 & 2_n9763;
assign 2_n4538 = ~(2_n10048 ^ 2_n9129);
assign 2_n9643 = ~(2_n3954 | 2_n8955);
assign 2_n10727 = 2_n346 | 2_n7721;
assign 2_n11905 = 2_n1937 | 2_n7876;
assign 2_n8946 = 2_n60 | 2_n11213;
assign 2_n1267 = 2_n8428 | 2_n5012;
assign 2_n2893 = 2_n5355 | 2_n7341;
assign 2_n5986 = ~(2_n12870 | 2_n10107);
assign 2_n3617 = ~2_n1199;
assign 2_n4994 = 2_n994 | 2_n7341;
assign 2_n2874 = 2_n5575 | 2_n8414;
assign 2_n2134 = ~2_n6946;
assign 2_n1566 = 2_n10010 | 2_n10815;
assign 2_n2436 = 2_n8900 & 2_n5531;
assign 2_n5639 = ~(2_n3653 ^ 2_n2021);
assign 2_n7552 = 2_n11317 & 2_n1265;
assign 2_n8102 = 2_n10464 & 2_n4164;
assign 2_n1305 = 2_n2064 | 2_n5122;
assign 2_n11133 = 2_n2619 | 2_n4978;
assign 2_n3785 = ~(2_n4256 ^ 2_n5534);
assign 2_n5006 = ~2_n8765;
assign 2_n1024 = 2_n12119 | 2_n1163;
assign 2_n6455 = ~2_n3719;
assign 2_n2716 = ~2_n8275;
assign 2_n5589 = 2_n10835 | 2_n4642;
assign 2_n12090 = 2_n3715 | 2_n9788;
assign 2_n1695 = 2_n9370 | 2_n7881;
assign 2_n8981 = 2_n5059 | 2_n11994;
assign 2_n7008 = ~(2_n110 ^ 2_n2882);
assign 2_n269 = ~2_n9581;
assign 2_n8991 = 2_n2850 | 2_n9469;
assign 2_n11732 = 2_n2408 & 2_n1931;
assign 2_n10210 = 2_n4778 | 2_n7382;
assign 2_n12857 = ~(2_n9907 | 2_n9927);
assign 2_n8621 = ~(2_n6085 ^ 2_n4762);
assign 2_n5997 = ~(2_n7037 ^ 2_n8613);
assign 2_n9196 = 2_n8187 | 2_n3911;
assign 2_n7417 = ~(2_n6165 | 2_n8787);
assign 2_n7039 = ~(2_n10877 ^ 2_n4406);
assign 2_n1531 = 2_n7195 & 2_n7793;
assign 2_n230 = ~(2_n7457 ^ 2_n9017);
assign 2_n10724 = ~(2_n11537 ^ 2_n11206);
assign 2_n8883 = ~(2_n8750 | 2_n10537);
assign 2_n4941 = 2_n7503 | 2_n11066;
assign 2_n5121 = ~2_n5590;
assign 2_n5117 = ~(2_n5969 ^ 2_n11591);
assign 2_n7509 = 2_n6577 | 2_n6455;
assign 2_n7121 = 2_n5765 | 2_n1476;
assign 2_n5732 = 2_n191 | 2_n1455;
assign 2_n12508 = ~(2_n12059 ^ 2_n2796);
assign 2_n1900 = 2_n6131 & 2_n2060;
assign 2_n12680 = 2_n8406 | 2_n2607;
assign 2_n2060 = 2_n3486 & 2_n7825;
assign 2_n8953 = ~(2_n12761 ^ 2_n50);
assign 2_n3731 = ~(2_n10435 ^ 2_n4895);
assign 2_n9412 = ~(2_n8750 ^ 2_n6167);
assign 2_n5156 = ~2_n8289;
assign 2_n11777 = 2_n9138 & 2_n2135;
assign 2_n265 = ~2_n7576;
assign 2_n2162 = 2_n5765 | 2_n7921;
assign 2_n2732 = 2_n7149 | 2_n9026;
assign 2_n8050 = 2_n12385 & 2_n12353;
assign 2_n12326 = 2_n4500 & 2_n1483;
assign 2_n3763 = ~(2_n9814 | 2_n9609);
assign 2_n3321 = 2_n6650 & 2_n5386;
assign 2_n11169 = 2_n1899 | 2_n5376;
assign 2_n101 = 2_n1197 | 2_n4827;
assign 2_n12238 = ~(2_n2227 | 2_n9716);
assign 2_n10542 = 2_n8496 | 2_n4583;
assign 2_n1047 = ~2_n1980;
assign 2_n1102 = 2_n2363 | 2_n229;
assign 2_n12491 = ~(2_n10346 | 2_n7372);
assign 2_n8603 = 2_n5077 & 2_n12350;
assign 2_n10382 = ~2_n5029;
assign 2_n3597 = ~2_n11953;
assign 2_n7634 = ~2_n3881;
assign 2_n4254 = 2_n11958 | 2_n5311;
assign 2_n10654 = ~(2_n5569 ^ 2_n1877);
assign 2_n3450 = ~(2_n9108 ^ 2_n3983);
assign 2_n1175 = ~2_n11198;
assign 2_n830 = 2_n6090 | 2_n2811;
assign 2_n2806 = 2_n9231 & 2_n6051;
assign 2_n12603 = ~2_n11685;
assign 2_n1575 = ~2_n4492;
assign 2_n5453 = 2_n2217 | 2_n3599;
assign 2_n9739 = 2_n4805 & 2_n1564;
assign 2_n5948 = 2_n8026 | 2_n11410;
assign 2_n8470 = ~2_n9842;
assign 2_n1146 = 2_n9797 & 2_n2900;
assign 2_n3898 = ~(2_n1037 ^ 2_n2402);
assign 2_n10806 = 2_n11239 | 2_n5980;
assign 2_n6128 = ~2_n5673;
assign 2_n9792 = ~(2_n7827 ^ 2_n711);
assign 2_n4289 = 2_n752 | 2_n3468;
assign 2_n3678 = 2_n11923 | 2_n609;
assign 2_n10081 = 2_n5995 & 2_n769;
assign 2_n3630 = ~(2_n8817 | 2_n4099);
assign 2_n7259 = ~(2_n9655 ^ 2_n865);
assign 2_n2326 = 2_n7449 | 2_n3606;
assign 2_n170 = ~(2_n12492 ^ 2_n425);
assign 2_n4305 = ~2_n3257;
assign 2_n4973 = ~2_n3428;
assign 2_n3676 = ~(2_n12104 ^ 2_n11215);
assign 2_n7334 = 2_n4059 | 2_n6389;
assign 2_n9726 = ~2_n2440;
assign 2_n7114 = 2_n9389 | 2_n8524;
assign 2_n1941 = ~2_n4187;
assign 2_n3619 = 2_n12052 & 2_n9818;
assign 2_n1218 = ~(2_n2268 ^ 2_n7047);
assign 2_n11234 = 2_n11552 | 2_n9144;
assign 2_n7560 = ~2_n131;
assign 2_n11998 = 2_n6577 | 2_n2232;
assign 2_n8979 = ~(2_n10730 ^ 2_n4507);
assign 2_n8375 = ~2_n267;
assign 2_n628 = 2_n3097 | 2_n7281;
assign 2_n2375 = ~(2_n6326 ^ 2_n6631);
assign 2_n4900 = 2_n1814 & 2_n739;
assign 2_n3280 = ~2_n5405;
assign 2_n8729 = 2_n9976 | 2_n1638;
assign 2_n9000 = 2_n10835 | 2_n3606;
assign 2_n4010 = 2_n2562 & 2_n5484;
assign 2_n48 = ~(2_n11025 ^ 2_n6958);
assign 2_n9908 = 2_n2213 | 2_n1443;
assign 2_n8256 = 2_n973 | 2_n12170;
assign 2_n12048 = ~(2_n12879 ^ 2_n10887);
assign 2_n5911 = ~(2_n54 ^ 2_n11751);
assign 2_n7680 = 2_n250 ^ 2_n11151;
assign 2_n10599 = ~(2_n10018 ^ 2_n10021);
assign 2_n7205 = 2_n1471 & 2_n8028;
assign 2_n9367 = 2_n7268 & 2_n1767;
assign 2_n11252 = 2_n9141 & 2_n5149;
assign 2_n10827 = ~2_n7233;
assign 2_n449 = 2_n10532 & 2_n7374;
assign 2_n1232 = 2_n8538 & 2_n1504;
assign 2_n6244 = 2_n11552 | 2_n3606;
assign 2_n8919 = 2_n5577 & 2_n7816;
assign 2_n8971 = ~(2_n4561 ^ 2_n10280);
assign 2_n12239 = ~(2_n12775 ^ 2_n12157);
assign 2_n5133 = ~(2_n7605 ^ 2_n3031);
assign 2_n6631 = 2_n9182 & 2_n6245;
assign 2_n10309 = 2_n3743 | 2_n8830;
assign 2_n12435 = 2_n1708 & 2_n12114;
assign 2_n11621 = 2_n6413 | 2_n166;
assign 2_n6742 = 2_n3166 ^ 2_n3894;
assign 2_n6600 = ~(2_n12129 | 2_n12573);
assign 2_n3038 = 2_n9370 | 2_n11827;
assign 2_n10567 = ~(2_n3543 ^ 2_n4861);
assign 2_n1166 = 2_n11433 | 2_n12816;
assign 2_n9283 = ~(2_n2817 ^ 2_n12589);
assign 2_n6436 = ~(2_n12370 ^ 2_n10650);
assign 2_n1943 = 2_n2118 | 2_n1155;
assign 2_n169 = ~(2_n11073 ^ 2_n10424);
assign 2_n3075 = ~(2_n8054 ^ 2_n9338);
assign 2_n385 = 2_n5038 | 2_n2570;
assign 2_n1996 = ~2_n7035;
assign 2_n1137 = 2_n1233 | 2_n6330;
assign 2_n10220 = 2_n2536 & 2_n12112;
assign 2_n5505 = 2_n2067 | 2_n12568;
assign 2_n10481 = ~(2_n7332 ^ 2_n6932);
assign 2_n9308 = 2_n10142 | 2_n2358;
assign 2_n12350 = 2_n3874 | 2_n6060;
assign 2_n7128 = 2_n6055 | 2_n6997;
assign 2_n11293 = 2_n705 | 2_n1310;
assign 2_n6868 = ~(2_n9692 | 2_n4439);
assign 2_n2046 = ~2_n1104;
assign 2_n2243 = 2_n10390 | 2_n10883;
assign 2_n10364 = ~2_n12949;
assign 2_n10417 = ~(2_n267 ^ 2_n3548);
assign 2_n9388 = ~(2_n1630 ^ 2_n2046);
assign 2_n305 = 2_n6977 | 2_n7952;
assign 2_n12607 = ~(2_n6993 | 2_n9915);
assign 2_n4235 = ~(2_n8945 | 2_n1859);
assign 2_n11382 = 2_n6080 | 2_n2953;
assign 2_n10005 = ~(2_n6872 ^ 2_n7751);
assign 2_n11441 = ~(2_n4728 ^ 2_n12275);
assign 2_n11879 = 2_n3743 | 2_n6922;
assign 2_n11531 = 2_n2593 & 2_n8497;
assign 2_n3998 = ~2_n2209;
assign 2_n8828 = ~(2_n978 ^ 2_n977);
assign 2_n4118 = ~(2_n3372 ^ 2_n5322);
assign 2_n4367 = 2_n8521 ^ 2_n10445;
assign 2_n3572 = ~(2_n3302 ^ 2_n3771);
assign 2_n7376 = 2_n11958 | 2_n3903;
assign 2_n11897 = ~(2_n6722 ^ 2_n8318);
assign 2_n5988 = 2_n3617 | 2_n826;
assign 2_n5328 = ~2_n9606;
assign 2_n9793 = 2_n215 | 2_n939;
assign 2_n7779 = ~(2_n2788 ^ 2_n12627);
assign 2_n2556 = 2_n9584 | 2_n9521;
assign 2_n4627 = 2_n12091 | 2_n2348;
assign 2_n3871 = ~(2_n11444 ^ 2_n439);
assign 2_n6469 = ~(2_n1646 ^ 2_n11022);
assign 2_n3164 = ~(2_n12421 | 2_n10063);
assign 2_n11888 = ~(2_n12610 ^ 2_n10283);
assign 2_n9326 = 2_n2099 | 2_n12535;
assign 2_n12183 = ~(2_n10100 | 2_n9839);
assign 2_n351 = ~2_n400;
assign 2_n11860 = ~2_n3797;
assign 2_n5537 = 2_n3746 | 2_n12899;
assign 2_n2603 = 2_n6027 & 2_n2250;
assign 2_n9077 = ~2_n12952;
assign 2_n3702 = ~(2_n7491 | 2_n10470);
assign 2_n3271 = 2_n10663 | 2_n8937;
assign 2_n11290 = 2_n6939 | 2_n208;
assign 2_n11974 = 2_n8203 | 2_n10722;
assign 2_n9750 = ~(2_n7667 | 2_n9348);
assign 2_n7162 = ~(2_n3404 ^ 2_n12828);
assign 2_n3374 = 2_n1699 | 2_n530;
assign 2_n8353 = 2_n10835 | 2_n12771;
assign 2_n3032 = 2_n9048 | 2_n5993;
assign 2_n12854 = ~(2_n2729 ^ 2_n647);
assign 2_n6053 = 2_n5530 | 2_n7928;
assign 2_n11373 = ~(2_n9084 ^ 2_n9478);
assign 2_n4303 = 2_n4059 | 2_n1162;
assign 2_n2341 = ~(2_n3376 | 2_n12134);
assign 2_n3135 = ~(2_n7542 | 2_n12896);
assign 2_n4498 = ~2_n5240;
assign 2_n4894 = 2_n5779 & 2_n10102;
assign 2_n473 = 2_n5674 & 2_n11330;
assign 2_n12230 = ~(2_n7493 ^ 2_n8075);
assign 2_n10939 = ~2_n3424;
assign 2_n10269 = 2_n7116 | 2_n2815;
assign 2_n9306 = 2_n2292 | 2_n662;
assign 2_n4395 = ~(2_n5364 ^ 2_n12595);
assign 2_n588 = 2_n6718 | 2_n8643;
assign 2_n12859 = ~2_n4325;
assign 2_n10830 = 2_n5967 & 2_n3028;
assign 2_n9444 = 2_n994 | 2_n1455;
assign 2_n4474 = ~2_n9763;
assign 2_n7948 = 2_n5441 & 2_n1862;
assign 2_n6017 = ~(2_n3577 | 2_n46);
assign 2_n7654 = 2_n12310 & 2_n9430;
assign 2_n1121 = 2_n3133 & 2_n10313;
assign 2_n10561 = ~2_n3769;
assign 2_n6964 = ~(2_n8547 ^ 2_n4020);
assign 2_n6401 = ~(2_n7779 | 2_n10248);
assign 2_n3903 = ~2_n6126;
assign 2_n10303 = ~(2_n12436 ^ 2_n12389);
assign 2_n12635 = ~(2_n7170 | 2_n9038);
assign 2_n9935 = ~(2_n1537 | 2_n8188);
assign 2_n2037 = 2_n7313 | 2_n3640;
assign 2_n10651 = ~(2_n10423 ^ 2_n4517);
assign 2_n8441 = 2_n2686 | 2_n10618;
assign 2_n11273 = 2_n8545 & 2_n12783;
assign 2_n3924 = ~2_n8665;
assign 2_n819 = 2_n11744 & 2_n2222;
assign 2_n1472 = 2_n10761 & 2_n3234;
assign 2_n7629 = 2_n3984 | 2_n3902;
assign 2_n4014 = ~2_n2106;
assign 2_n3220 = 2_n5116 | 2_n11361;
assign 2_n3470 = 2_n4299 & 2_n5698;
assign 2_n3122 = ~(2_n7620 ^ 2_n1181);
assign 2_n3658 = ~2_n6631;
assign 2_n8826 = ~(2_n3221 | 2_n3314);
assign 2_n11957 = ~(2_n9162 ^ 2_n7106);
assign 2_n2733 = 2_n12818 | 2_n541;
assign 2_n10266 = 2_n5138 | 2_n8471;
assign 2_n6084 = ~2_n8065;
assign 2_n9607 = ~2_n4659;
assign 2_n2316 = ~(2_n11439 ^ 2_n1609);
assign 2_n3471 = ~(2_n7335 ^ 2_n8466);
assign 2_n12944 = ~(2_n4246 ^ 2_n4265);
assign 2_n6165 = 2_n8451 & 2_n5430;
assign 2_n1264 = 2_n12079 & 2_n1704;
assign 2_n8225 = 2_n5515 & 2_n6683;
assign 2_n9286 = ~(2_n10560 | 2_n5029);
assign 2_n11 = 2_n4628 | 2_n8259;
assign 2_n10785 = ~(2_n9844 ^ 2_n9225);
assign 2_n357 = 2_n7283 | 2_n7341;
assign 2_n592 = 2_n9990 & 2_n2840;
assign 2_n495 = ~(2_n602 ^ 2_n10024);
assign 2_n2458 = ~(2_n10289 ^ 2_n6679);
assign 2_n633 = 2_n9554 | 2_n8507;
assign 2_n3049 = ~(2_n12008 ^ 2_n5555);
assign 2_n209 = ~2_n7936;
assign 2_n833 = ~(2_n3220 ^ 2_n5675);
assign 2_n10442 = ~2_n2826;
assign 2_n1986 = ~(2_n5571 ^ 2_n537);
assign 2_n57 = ~(2_n2950 ^ 2_n7252);
assign 2_n3673 = 2_n1623 & 2_n7323;
assign 2_n9541 = 2_n9370 | 2_n1546;
assign 2_n5416 = 2_n6256 | 2_n7489;
assign 2_n5815 = 2_n9107 & 2_n2986;
assign 2_n10729 = ~2_n4468;
assign 2_n18 = ~(2_n4514 | 2_n9659);
assign 2_n11832 = 2_n10945 | 2_n7318;
assign 2_n3563 = ~(2_n5101 | 2_n9206);
assign 2_n7210 = ~(2_n8273 ^ 2_n4909);
assign 2_n2319 = 2_n2217 | 2_n6922;
assign 2_n7088 = 2_n8870 | 2_n6513;
assign 2_n10012 = 2_n9170 | 2_n6389;
assign 2_n11769 = 2_n1075 | 2_n8013;
assign 2_n4151 = ~(2_n6050 ^ 2_n3424);
assign 2_n5368 = 2_n309 & 2_n8529;
assign 2_n7042 = ~(2_n11443 ^ 2_n11237);
assign 2_n5031 = 2_n6718 | 2_n28;
assign 2_n3760 = ~2_n3001;
assign 2_n12527 = 2_n636 | 2_n8109;
assign 2_n10699 = ~(2_n3428 ^ 2_n1166);
assign 2_n1794 = ~2_n11154;
assign 2_n6190 = ~(2_n832 | 2_n3178);
assign 2_n2684 = 2_n4332 & 2_n9232;
assign 2_n10199 = 2_n5530 | 2_n4818;
assign 2_n12866 = ~(2_n8045 ^ 2_n7557);
assign 2_n929 = 2_n8127 | 2_n12843;
assign 2_n8658 = ~(2_n5415 ^ 2_n4248);
assign 2_n2179 = ~(2_n9064 | 2_n3185);
assign 2_n1581 = 2_n3976 | 2_n12059;
assign 2_n6711 = ~(2_n5733 ^ 2_n1237);
assign 2_n4636 = ~2_n313;
assign 2_n8280 = ~2_n8281;
assign 2_n2921 = 2_n6948 | 2_n8357;
assign 2_n10805 = 2_n11061 | 2_n9759;
assign 2_n1527 = ~(2_n6151 | 2_n11219);
assign 2_n6141 = ~2_n6330;
assign 2_n5424 = 2_n7273 & 2_n5985;
assign 2_n11792 = 2_n6072 & 2_n891;
assign 2_n5938 = 2_n3042 | 2_n2965;
assign 2_n6646 = ~(2_n5865 ^ 2_n8480);
assign 2_n276 = 2_n3127 | 2_n5497;
assign 2_n9575 = ~(2_n1215 ^ 2_n5055);
assign 2_n9456 = ~(2_n6516 ^ 2_n9533);
assign 2_n2491 = 2_n582 | 2_n11014;
assign 2_n715 = ~(2_n12912 ^ 2_n8916);
assign 2_n4372 = ~(2_n10776 ^ 2_n4809);
assign 2_n3078 = 2_n989 | 2_n2358;
assign 2_n6660 = 2_n8187 | 2_n1546;
assign 2_n5358 = ~(2_n4917 ^ 2_n5870);
assign 2_n12851 = ~(2_n11397 ^ 2_n5821);
assign 2_n11208 = ~(2_n2395 ^ 2_n8893);
assign 2_n3786 = 2_n5989 & 2_n6704;
assign 2_n10315 = 2_n11026 | 2_n1509;
assign 2_n11985 = 2_n3324 | 2_n12771;
assign 2_n845 = ~(2_n5244 ^ 2_n5443);
assign 2_n7865 = 2_n6457 | 2_n12627;
assign 2_n12448 = 2_n8748 & 2_n4814;
assign 2_n9287 = 2_n8054 | 2_n3524;
assign 2_n876 = 2_n11527 & 2_n8072;
assign 2_n2913 = 2_n4862 & 2_n5230;
assign 2_n1087 = 2_n9212 & 2_n9932;
assign 2_n12171 = 2_n5473 | 2_n11792;
assign 2_n11164 = ~(2_n9910 ^ 2_n4795);
assign 2_n3507 = 2_n1695 & 2_n8066;
assign 2_n1825 = ~2_n1697;
assign 2_n309 = ~2_n12348;
assign 2_n4912 = ~2_n9026;
assign 2_n11764 = 2_n9432 | 2_n7226;
assign 2_n3088 = 2_n8649 & 2_n9624;
assign 2_n7614 = ~(2_n5485 ^ 2_n5083);
assign 2_n898 = 2_n7701 | 2_n10486;
assign 2_n1662 = ~(2_n5161 ^ 2_n4915);
assign 2_n6293 = 2_n9389 | 2_n11827;
assign 2_n9598 = 2_n9698 & 2_n665;
assign 2_n11994 = ~2_n4099;
assign 2_n8193 = 2_n8554 & 2_n10561;
assign 2_n10862 = 2_n8326 | 2_n10044;
assign 2_n5213 = ~(2_n438 ^ 2_n12631);
assign 2_n5963 = ~(2_n9819 ^ 2_n10795);
assign 2_n381 = ~(2_n3941 ^ 2_n11054);
assign 2_n12836 = ~(2_n5247 ^ 2_n9020);
assign 2_n11301 = ~(2_n4034 ^ 2_n400);
assign 2_n4657 = 2_n7687 | 2_n2352;
assign 2_n8884 = ~(2_n8544 ^ 2_n5051);
assign 2_n10433 = ~(2_n4500 | 2_n1483);
assign 2_n3880 = ~(2_n346 ^ 2_n7721);
assign 2_n2078 = 2_n1909 & 2_n1773;
assign 2_n9249 = ~(2_n2444 | 2_n1176);
assign 2_n1442 = ~2_n7909;
assign 2_n9253 = ~(2_n2918 ^ 2_n10425);
assign 2_n8097 = 2_n2082 & 2_n7007;
assign 2_n205 = ~(2_n6966 | 2_n11981);
assign 2_n7336 = ~2_n10751;
assign 2_n637 = 2_n10601 | 2_n3576;
assign 2_n12877 = 2_n10196 | 2_n8830;
assign 2_n5430 = 2_n8110 | 2_n2767;
assign 2_n5912 = 2_n7715 & 2_n3883;
assign 2_n8564 = 2_n11457 | 2_n4240;
assign 2_n11122 = ~2_n2433;
assign 2_n12543 = ~2_n10998;
assign 2_n4819 = 2_n4778 | 2_n10854;
assign 2_n6130 = 2_n8305 | 2_n1667;
assign 2_n6096 = 2_n9170 | 2_n1162;
assign 2_n9437 = 2_n6687 & 2_n2879;
assign 2_n3951 = 2_n3609 | 2_n11286;
assign 2_n7037 = 2_n3127 | 2_n7424;
assign 2_n9605 = ~(2_n3474 ^ 2_n8780);
assign 2_n7000 = ~(2_n11233 ^ 2_n3489);
assign 2_n7070 = ~(2_n9179 | 2_n9479);
assign 2_n9847 = ~(2_n8163 ^ 2_n4448);
assign 2_n4640 = ~(2_n9846 ^ 2_n5409);
assign 2_n9301 = 2_n7391 | 2_n7341;
assign 2_n12845 = 2_n11547 | 2_n6832;
assign 2_n2281 = ~(2_n11390 ^ 2_n3431);
assign 2_n167 = 2_n8345 | 2_n2635;
assign 2_n1987 = ~2_n7505;
assign 2_n5124 = ~(2_n3864 ^ 2_n10234);
assign 2_n5765 = ~2_n11153;
assign 2_n4662 = ~(2_n4135 | 2_n5339);
assign 2_n1872 = 2_n2924 & 2_n2141;
assign 2_n3701 = ~(2_n10332 ^ 2_n9484);
assign 2_n3580 = ~2_n9194;
assign 2_n2115 = ~(2_n4480 ^ 2_n7123);
assign 2_n4199 = 2_n1972 & 2_n3977;
assign 2_n860 = ~(2_n469 ^ 2_n7349);
assign 2_n12540 = 2_n2537 & 2_n151;
assign 2_n5616 = ~2_n11053;
assign 2_n12495 = 2_n8792 | 2_n7972;
assign 2_n6421 = ~(2_n11155 ^ 2_n3574);
assign 2_n5545 = ~(2_n10359 ^ 2_n8424);
assign 2_n1111 = 2_n3743 | 2_n3606;
assign 2_n5562 = 2_n12853 | 2_n8740;
assign 2_n10170 = ~2_n10034;
assign 2_n3043 = ~(2_n2060 ^ 2_n6131);
assign 2_n2612 = ~2_n12619;
assign 2_n4625 = 2_n7977 | 2_n755;
assign 2_n6373 = ~2_n11892;
assign 2_n1246 = 2_n8221 | 2_n11268;
assign 2_n4833 = 2_n12683 & 2_n6552;
assign 2_n8354 = ~2_n3616;
assign 2_n2219 = 2_n5708 & 2_n12892;
assign 2_n2908 = ~(2_n5819 ^ 2_n1697);
assign 2_n7227 = ~(2_n4170 ^ 2_n10599);
assign 2_n709 = 2_n6628 & 2_n11372;
assign 2_n6222 = 2_n12087 & 2_n4267;
assign 2_n4857 = ~(2_n3885 ^ 2_n11729);
assign 2_n2202 = ~2_n9275;
assign 2_n7193 = ~(2_n1505 ^ 2_n4118);
assign 2_n11156 = ~(2_n4021 ^ 2_n10654);
assign 2_n9044 = ~(2_n7295 | 2_n2785);
assign 2_n9244 = ~(2_n7316 | 2_n9090);
assign 2_n8429 = ~2_n7824;
assign 2_n2993 = 2_n12186 | 2_n2815;
assign 2_n2593 = ~(2_n10028 ^ 2_n4651);
assign 2_n2557 = ~2_n9982;
assign 2_n4568 = 2_n10852 & 2_n12019;
assign 2_n3672 = 2_n24 | 2_n7334;
assign 2_n5292 = 2_n6718 | 2_n795;
assign 2_n7352 = 2_n4100 | 2_n9385;
assign 2_n5042 = ~2_n9307;
assign 2_n1326 = 2_n11552 | 2_n4642;
assign 2_n5706 = 2_n3820 | 2_n8643;
assign 2_n1190 = 2_n7788 & 2_n11654;
assign 2_n4065 = 2_n5858 | 2_n1455;
assign 2_n6552 = 2_n2478 | 2_n2387;
assign 2_n93 = ~(2_n6767 ^ 2_n1508);
assign 2_n4360 = 2_n4498 | 2_n1455;
assign 2_n6273 = ~(2_n10382 ^ 2_n11167);
assign 2_n5081 = 2_n5964 & 2_n11662;
assign 2_n9982 = 2_n7124 & 2_n4307;
assign 2_n7408 = ~(2_n12272 ^ 2_n6950);
assign 2_n11730 = 2_n1757 & 2_n303;
assign 2_n6805 = ~(2_n8532 | 2_n442);
assign 2_n10090 = ~(2_n6995 ^ 2_n9305);
assign 2_n12273 = 2_n4856 | 2_n10610;
assign 2_n6356 = ~(2_n913 ^ 2_n8493);
assign 2_n4442 = 2_n10647 ^ 2_n10009;
assign 2_n2428 = 2_n1224 & 2_n8422;
assign 2_n11463 = 2_n10078 & 2_n8652;
assign 2_n3711 = ~(2_n6962 ^ 2_n7049);
assign 2_n8204 = 2_n6776 & 2_n12145;
assign 2_n4859 = 2_n2099 | 2_n9586;
assign 2_n11753 = ~2_n3541;
assign 2_n10667 = 2_n2217 | 2_n8745;
assign 2_n10665 = ~(2_n8197 ^ 2_n1098);
assign 2_n380 = ~2_n9698;
assign 2_n8321 = 2_n10879 | 2_n7424;
assign 2_n4405 = ~2_n4070;
assign 2_n6802 = 2_n9806 & 2_n8579;
assign 2_n10420 = ~(2_n3365 | 2_n5811);
assign 2_n9799 = ~(2_n9669 | 2_n12196);
assign 2_n9145 = ~(2_n1622 ^ 2_n10189);
assign 2_n1813 = 2_n2102 & 2_n517;
assign 2_n1787 = ~(2_n7663 ^ 2_n11886);
assign 2_n11666 = 2_n6244 & 2_n8180;
assign 2_n7028 = 2_n2854 | 2_n1961;
assign 2_n397 = 2_n649 ^ 2_n8270;
assign 2_n12220 = ~2_n6553;
assign 2_n3378 = 2_n4272 | 2_n11833;
assign 2_n88 = ~2_n1795;
assign 2_n9094 = ~(2_n7254 ^ 2_n11190);
assign 2_n4418 = 2_n9528 | 2_n10054;
assign 2_n3665 = 2_n3819 & 2_n2966;
assign 2_n11113 = ~(2_n4060 | 2_n2225);
assign 2_n9083 = ~2_n4463;
assign 2_n10553 = ~2_n987;
assign 2_n12795 = ~(2_n1560 ^ 2_n12697);
assign 2_n12275 = 2_n2414 & 2_n1920;
assign 2_n10089 = 2_n8959 | 2_n11122;
assign 2_n11076 = 2_n12853 | 2_n3224;
assign 2_n12062 = ~(2_n4273 | 2_n11934);
assign 2_n3361 = ~2_n9627;
assign 2_n2021 = ~(2_n3757 ^ 2_n10363);
assign 2_n4976 = 2_n632 & 2_n4881;
assign 2_n12685 = ~(2_n2230 | 2_n7302);
assign 2_n7984 = ~(2_n5332 ^ 2_n12952);
assign 2_n6889 = ~(2_n5380 ^ 2_n4305);
assign 2_n3074 = 2_n6509 & 2_n2657;
assign 2_n4146 = 2_n2872 | 2_n2815;
assign 2_n5179 = 2_n752 | 2_n11122;
assign 2_n5137 = ~(2_n7418 ^ 2_n3061);
assign 2_n9736 = ~2_n5931;
assign 2_n4202 = 2_n10196 | 2_n9568;
assign 2_n11928 = 2_n752 | 2_n7395;
assign 2_n5144 = ~(2_n9 ^ 2_n12486);
assign 2_n7129 = ~2_n11307;
assign 2_n5702 = ~(2_n9340 ^ 2_n263);
assign 2_n4503 = 2_n9945 | 2_n11486;
assign 2_n9097 = ~(2_n4074 | 2_n5104);
assign 2_n3750 = 2_n10741 | 2_n10149;
assign 2_n6364 = 2_n5860 & 2_n10898;
assign 2_n9695 = ~(2_n3508 ^ 2_n12096);
assign 2_n9260 = 2_n11719 | 2_n4400;
assign 2_n815 = ~(2_n7062 ^ 2_n145);
assign 2_n2636 = ~(2_n2098 ^ 2_n6959);
assign 2_n12762 = ~(2_n1458 ^ 2_n3942);
assign 2_n6229 = ~(2_n3228 | 2_n2603);
assign 2_n12563 = ~(2_n6620 ^ 2_n11660);
assign 2_n418 = 2_n5809 | 2_n9188;
assign 2_n11686 = ~(2_n9905 ^ 2_n10792);
assign 2_n9537 = ~(2_n861 ^ 2_n9545);
assign 2_n2928 = 2_n2559 & 2_n502;
assign 2_n15 = 2_n10615 & 2_n4699;
assign 2_n2480 = ~(2_n4349 ^ 2_n4927);
assign 2_n6043 = 2_n5061 | 2_n11720;
assign 2_n6325 = 2_n3265 | 2_n1454;
assign 2_n2022 = 2_n8137 & 2_n7076;
assign 2_n8525 = 2_n2833 & 2_n553;
assign 2_n44 = ~(2_n12223 ^ 2_n4389);
assign 2_n9986 = ~(2_n3464 ^ 2_n8805);
assign 2_n2255 = ~(2_n7984 ^ 2_n6362);
assign 2_n10137 = ~(2_n3233 | 2_n4402);
assign 2_n10141 = 2_n8552 | 2_n9586;
assign 2_n1889 = 2_n5084 & 2_n562;
assign 2_n10954 = ~(2_n9872 ^ 2_n6941);
assign 2_n376 = 2_n959 | 2_n5155;
assign 2_n12344 = 2_n2969 | 2_n11072;
assign 2_n1009 = 2_n5575 | 2_n2232;
assign 2_n3491 = 2_n7391 | 2_n4242;
assign 2_n5641 = 2_n1548 ^ 2_n6838;
assign 2_n6345 = 2_n4178 | 2_n1751;
assign 2_n10377 = 2_n2099 | 2_n12446;
assign 2_n5542 = 2_n752 | 2_n184;
assign 2_n2866 = ~2_n6085;
assign 2_n9390 = ~(2_n5476 ^ 2_n8360);
assign 2_n1993 = 2_n11749 | 2_n4165;
assign 2_n6160 = 2_n11181 & 2_n4268;
assign 2_n8212 = ~(2_n12537 | 2_n11978);
assign 2_n4178 = 2_n239 | 2_n8788;
assign 2_n10720 = ~(2_n1059 ^ 2_n10875);
assign 2_n11953 = 2_n5032 | 2_n760;
assign 2_n11684 = ~(2_n489 | 2_n10184);
assign 2_n12059 = ~(2_n366 ^ 2_n2035);
assign 2_n8560 = 2_n7539 | 2_n1328;
assign 2_n2003 = ~(2_n11173 ^ 2_n8603);
assign 2_n9743 = ~2_n1853;
assign 2_n3486 = 2_n12033 | 2_n6781;
assign 2_n11947 = 2_n584 & 2_n8887;
assign 2_n12687 = ~2_n1166;
assign 2_n4565 = ~2_n9993;
assign 2_n12402 = ~(2_n6125 ^ 2_n2867);
assign 2_n4337 = 2_n12837 & 2_n12554;
assign 2_n396 = 2_n12361 | 2_n3421;
assign 2_n164 = 2_n11856 | 2_n6911;
assign 2_n1290 = ~(2_n12859 | 2_n2412);
assign 2_n3070 = 2_n6147 & 2_n9876;
assign 2_n2510 = ~(2_n6551 | 2_n2086);
assign 2_n7020 = ~(2_n8553 ^ 2_n5073);
assign 2_n5228 = 2_n10833 | 2_n7761;
assign 2_n1568 = ~(2_n1424 | 2_n8707);
assign 2_n4971 = ~(2_n12818 ^ 2_n11461);
assign 2_n7528 = ~(2_n11414 ^ 2_n11375);
assign 2_n12312 = ~2_n7390;
assign 2_n5013 = ~2_n1688;
assign 2_n6177 = 2_n1699 | 2_n7928;
assign 2_n6997 = 2_n6795 & 2_n11424;
assign 2_n8961 = 2_n11421 | 2_n6212;
assign 2_n10108 = ~2_n9080;
assign 2_n5559 = 2_n2099 | 2_n7136;
assign 2_n2650 = 2_n5198 & 2_n9111;
assign 2_n3983 = 2_n839 & 2_n69;
assign 2_n9188 = ~2_n2558;
assign 2_n8481 = 2_n8026 | 2_n6197;
assign 2_n7831 = ~(2_n8022 ^ 2_n724);
assign 2_n2516 = ~(2_n8449 ^ 2_n4758);
assign 2_n11824 = ~(2_n1038 ^ 2_n3466);
assign 2_n3762 = ~(2_n11559 ^ 2_n6978);
assign 2_n7669 = 2_n5902 | 2_n3911;
assign 2_n7333 = ~(2_n7021 ^ 2_n10726);
assign 2_n4688 = ~(2_n8557 ^ 2_n7275);
assign 2_n6175 = 2_n6977 | 2_n7876;
assign 2_n7269 = ~(2_n4963 ^ 2_n9362);
assign 2_n491 = 2_n11200 & 2_n9393;
assign 2_n1642 = 2_n11958 | 2_n7425;
assign 2_n5864 = 2_n8354 | 2_n8740;
assign 2_n514 = 2_n11013 & 2_n1346;
assign 2_n1780 = ~2_n8600;
assign 2_n6777 = 2_n5355 | 2_n7246;
assign 2_n10710 = 2_n3324 | 2_n795;
assign 2_n10637 = ~(2_n9395 ^ 2_n10386);
assign 2_n11644 = ~(2_n5438 ^ 2_n1856);
assign 2_n3190 = 2_n10882 | 2_n9665;
assign 2_n12789 = 2_n9433 & 2_n11196;
assign 2_n8269 = 2_n683 | 2_n12834;
assign 2_n5335 = 2_n676 & 2_n4331;
assign 2_n1534 = 2_n8387 | 2_n12856;
assign 2_n653 = ~(2_n1181 | 2_n12808);
assign 2_n12869 = ~2_n4331;
assign 2_n3112 = ~(2_n987 ^ 2_n6367);
assign 2_n6335 = 2_n2505 & 2_n8388;
assign 2_n9777 = 2_n7176 | 2_n506;
assign 2_n1126 = 2_n7391 | 2_n10066;
assign 2_n8589 = 2_n11584 | 2_n4156;
assign 2_n11634 = 2_n4311 | 2_n2572;
assign 2_n8307 = 2_n10522 & 2_n2943;
assign 2_n7295 = 2_n1387 & 2_n2954;
assign 2_n6775 = ~2_n8966;
assign 2_n6808 = ~2_n10658;
assign 2_n1213 = ~(2_n2519 ^ 2_n4673);
assign 2_n12234 = ~(2_n53 ^ 2_n7541);
assign 2_n2675 = 2_n5190 | 2_n6371;
assign 2_n11562 = ~(2_n9381 ^ 2_n7277);
assign 2_n8821 = 2_n298 & 2_n8746;
assign 2_n7603 = ~(2_n12730 ^ 2_n3123);
assign 2_n9759 = ~(2_n9615 | 2_n5253);
assign 2_n4739 = ~(2_n4451 | 2_n1852);
assign 2_n6491 = ~2_n2721;
assign 2_n8579 = 2_n8354 | 2_n9188;
assign 2_n4015 = 2_n11266 | 2_n8286;
assign 2_n9554 = ~(2_n10658 | 2_n2513);
assign 2_n6565 = ~(2_n4049 ^ 2_n11554);
assign 2_n73 = 2_n7884 & 2_n1930;
assign 2_n4702 = 2_n7470 | 2_n1286;
assign 2_n6800 = 2_n1311 & 2_n799;
assign 2_n6250 = ~(2_n6285 ^ 2_n7515);
assign 2_n7457 = 2_n2099 | 2_n12883;
assign 2_n1701 = 2_n7154 | 2_n10837;
assign 2_n2211 = 2_n8727 & 2_n6756;
assign 2_n9106 = ~2_n253;
assign 2_n6004 = 2_n5575 | 2_n2754;
assign 2_n7260 = ~2_n5500;
assign 2_n928 = 2_n10750 | 2_n8740;
assign 2_n7135 = ~(2_n5137 ^ 2_n7340);
assign 2_n4476 = 2_n7709 | 2_n12771;
assign 2_n2064 = ~(2_n3284 ^ 2_n5841);
assign 2_n8395 = 2_n5915 | 2_n6513;
assign 2_n935 = 2_n4727 & 2_n4140;
assign 2_n6155 = ~(2_n10843 ^ 2_n1169);
assign 2_n5310 = ~(2_n1479 | 2_n1088);
assign 2_n8227 = 2_n3743 | 2_n4864;
assign 2_n7663 = 2_n2099 | 2_n8259;
assign 2_n415 = 2_n3776 | 2_n7665;
assign 2_n7989 = 2_n4576 & 2_n7365;
assign 2_n2180 = 2_n1684 & 2_n3408;
assign 2_n3656 = ~(2_n11556 ^ 2_n6173);
assign 2_n3158 = 2_n6654 & 2_n8578;
assign 2_n11760 = ~(2_n12037 ^ 2_n8968);
assign 2_n2364 = 2_n8476 & 2_n5645;
assign 2_n9645 = 2_n5179 | 2_n8417;
assign 2_n8873 = ~(2_n548 | 2_n2184);
assign 2_n574 = 2_n7709 | 2_n9521;
assign 2_n3206 = ~(2_n6518 ^ 2_n9790);
assign 2_n663 = ~(2_n9678 ^ 2_n9384);
assign 2_n3927 = 2_n8443 | 2_n12769;
assign 2_n4142 = ~(2_n11400 | 2_n7590);
assign 2_n402 = ~(2_n1299 ^ 2_n11634);
assign 2_n8466 = ~(2_n6548 ^ 2_n3910);
assign 2_n11987 = 2_n8441 & 2_n10645;
assign 2_n1611 = ~(2_n3213 ^ 2_n9694);
assign 2_n11051 = 2_n11764 & 2_n7533;
assign 2_n757 = 2_n7902 & 2_n10675;
assign 2_n2090 = 2_n3145 & 2_n1267;
assign 2_n10067 = ~(2_n8827 ^ 2_n364);
assign 2_n1365 = ~(2_n8652 ^ 2_n5293);
assign 2_n11795 = ~(2_n9755 ^ 2_n10274);
assign 2_n5246 = ~(2_n9227 | 2_n11615);
assign 2_n10307 = ~(2_n1142 | 2_n5933);
assign 2_n5700 = 2_n12659 & 2_n6846;
assign 2_n5571 = 2_n6577 | 2_n3468;
assign 2_n2427 = 2_n6577 | 2_n3903;
assign 2_n5620 = ~(2_n4719 | 2_n5723);
assign 2_n10066 = ~2_n6038;
assign 2_n12914 = 2_n989 | 2_n561;
assign 2_n1863 = 2_n9465 & 2_n3003;
assign 2_n8242 = ~(2_n5118 ^ 2_n4081);
assign 2_n1593 = 2_n257 | 2_n5333;
assign 2_n10490 = ~(2_n11400 ^ 2_n4691);
assign 2_n4509 = 2_n12177 | 2_n12386;
assign 2_n5418 = 2_n2564 & 2_n9956;
assign 2_n1573 = ~(2_n49 ^ 2_n8775);
assign 2_n7183 = ~(2_n4699 ^ 2_n7565);
assign 2_n3349 = 2_n5470 | 2_n4672;
assign 2_n5037 = ~(2_n4799 ^ 2_n4607);
assign 2_n11773 = 2_n6857 | 2_n4544;
assign 2_n6094 = ~(2_n9615 ^ 2_n10981);
assign 2_n1288 = 2_n9376 & 2_n11160;
assign 2_n3466 = ~(2_n10530 ^ 2_n3470);
assign 2_n10086 = 2_n2832 | 2_n12843;
assign 2_n9369 = 2_n9170 | 2_n7881;
assign 2_n10617 = ~(2_n623 ^ 2_n5157);
assign 2_n11546 = 2_n9492 | 2_n4420;
assign 2_n2519 = 2_n10534 & 2_n12546;
assign 2_n1687 = ~(2_n11231 ^ 2_n7553);
assign 2_n6895 = ~(2_n7752 ^ 2_n9868);
assign 2_n3476 = ~(2_n5242 ^ 2_n79);
assign 2_n6712 = 2_n5491 & 2_n7743;
assign 2_n7142 = ~(2_n762 ^ 2_n6312);
assign 2_n8340 = ~2_n203;
assign 2_n10378 = ~(2_n8912 ^ 2_n7830);
assign 2_n3420 = 2_n9895 & 2_n1832;
assign 2_n3533 = ~(2_n3880 ^ 2_n9498);
assign 2_n1840 = ~2_n5820;
assign 2_n1076 = 2_n3291 & 2_n8686;
assign 2_n8240 = ~2_n2680;
assign 2_n11908 = ~(2_n3038 ^ 2_n1030);
assign 2_n6145 = 2_n8959 | 2_n12816;
assign 2_n2955 = ~(2_n12939 ^ 2_n6858);
assign 2_n6759 = ~2_n8850;
assign 2_n2074 = 2_n7822 & 2_n5165;
assign 2_n4530 = ~(2_n11248 | 2_n7525);
assign 2_n5791 = 2_n5530 | 2_n4249;
assign 2_n3224 = ~2_n1564;
assign 2_n11943 = 2_n8387 & 2_n12856;
assign 2_n12245 = ~(2_n12367 | 2_n11600);
assign 2_n12926 = ~(2_n5564 ^ 2_n7451);
assign 2_n10560 = ~(2_n4058 ^ 2_n1554);
assign 2_n7057 = ~(2_n3016 ^ 2_n5356);
assign 2_n1949 = ~(2_n312 ^ 2_n11600);
assign 2_n2989 = 2_n10922 | 2_n8021;
assign 2_n8091 = 2_n10928 & 2_n4141;
assign 2_n3626 = ~(2_n1786 ^ 2_n10971);
assign 2_n4279 = ~(2_n7603 ^ 2_n11951);
assign 2_n1435 = ~(2_n5346 | 2_n9704);
assign 2_n3485 = 2_n3765 | 2_n3158;
assign 2_n2774 = ~(2_n7186 | 2_n11809);
assign 2_n9355 = 2_n8679 & 2_n1360;
assign 2_n997 = ~(2_n8646 | 2_n7314);
assign 2_n7213 = 2_n11569 | 2_n4115;
assign 2_n5254 = 2_n618 | 2_n7139;
assign 2_n6355 = ~(2_n6625 ^ 2_n7625);
assign 2_n7525 = 2_n4442 & 2_n4110;
assign 2_n8222 = 2_n3024 & 2_n7596;
assign 2_n12909 = ~2_n9819;
assign 2_n572 = ~(2_n12661 ^ 2_n1211);
assign 2_n1113 = 2_n12643 & 2_n4537;
assign 2_n8720 = ~2_n11987;
assign 2_n6477 = ~(2_n9657 ^ 2_n7969);
assign 2_n12010 = 2_n8127 | 2_n1851;
assign 2_n1373 = ~(2_n2150 ^ 2_n5723);
assign 2_n2617 = ~(2_n9825 ^ 2_n9776);
assign 2_n8988 = 2_n1151 | 2_n4573;
assign 2_n7335 = ~(2_n7915 ^ 2_n11435);
assign 2_n8214 = ~2_n9810;
assign 2_n4959 = ~(2_n7001 ^ 2_n12897);
assign 2_n494 = 2_n6718 | 2_n7506;
assign 2_n12683 = 2_n7831 | 2_n10979;
assign 2_n10064 = 2_n10018 | 2_n10021;
assign 2_n10563 = ~(2_n12460 ^ 2_n360);
assign 2_n2062 = ~(2_n12930 ^ 2_n9350);
assign 2_n11127 = 2_n3131 & 2_n10813;
assign 2_n10161 = ~(2_n1975 | 2_n11606);
assign 2_n4604 = ~2_n4437;
assign 2_n6204 = 2_n191 | 2_n7703;
assign 2_n10796 = ~(2_n10004 | 2_n7968);
assign 2_n3024 = 2_n868 | 2_n8323;
assign 2_n6060 = ~(2_n3791 ^ 2_n11806);
assign 2_n10526 = ~(2_n1681 ^ 2_n7048);
assign 2_n9057 = ~(2_n4063 ^ 2_n179);
assign 2_n297 = ~(2_n1830 | 2_n3860);
assign 2_n1983 = ~2_n9567;
assign 2_n8079 = ~(2_n9928 ^ 2_n2501);
assign 2_n5661 = 2_n8187 | 2_n11827;
assign 2_n6784 = 2_n1315 | 2_n2211;
assign 2_n10446 = ~(2_n1439 | 2_n9427);
assign 2_n5195 = 2_n3367 | 2_n3056;
assign 2_n6054 = ~2_n6335;
assign 2_n10104 = ~(2_n8198 ^ 2_n4403);
assign 2_n11697 = ~(2_n5574 | 2_n9133);
assign 2_n11695 = 2_n3617 | 2_n4913;
assign 2_n10363 = 2_n11923 | 2_n1509;
assign 2_n11669 = ~(2_n7280 ^ 2_n11909);
assign 2_n6032 = 2_n12413 & 2_n8866;
assign 2_n4154 = ~2_n12702;
assign 2_n5597 = 2_n2638 & 2_n8358;
assign 2_n9952 = ~2_n11459;
assign 2_n6707 = 2_n4560 & 2_n11334;
assign 2_n5998 = ~(2_n10710 ^ 2_n10083);
assign 2_n696 = ~(2_n8174 ^ 2_n12937);
assign 2_n1223 = ~(2_n1354 ^ 2_n9167);
assign 2_n5495 = ~(2_n5048 ^ 2_n1159);
assign 2_n707 = ~(2_n11931 ^ 2_n4008);
assign 2_n557 = 2_n12346 & 2_n12083;
assign 2_n11309 = ~(2_n1352 ^ 2_n7851);
assign 2_n5501 = 2_n10142 | 2_n8524;
assign 2_n10988 = ~2_n588;
assign 2_n2781 = ~(2_n11279 ^ 2_n11020);
assign 2_n8856 = ~2_n5665;
assign 2_n2938 = 2_n10132 | 2_n3476;
assign 2_n843 = 2_n3608 & 2_n3488;
assign 2_n4465 = 2_n6977 | 2_n2815;
assign 2_n8298 = ~(2_n4135 ^ 2_n8076);
assign 2_n10400 = 2_n3470 | 2_n9175;
assign 2_n2371 = 2_n5089 & 2_n10823;
assign 2_n3534 = 2_n3614 & 2_n8539;
assign 2_n7684 = ~(2_n272 ^ 2_n3095);
assign 2_n4198 = ~(2_n74 | 2_n7776);
assign 2_n940 = 2_n10339 | 2_n826;
assign 2_n6487 = ~(2_n3106 ^ 2_n1759);
assign 2_n8838 = 2_n11838 & 2_n7344;
assign 2_n9395 = 2_n3820 | 2_n1509;
assign 2_n8761 = 2_n7196 | 2_n4087;
assign 2_n10622 = 2_n8831 & 2_n3918;
assign 2_n3328 = 2_n6814 | 2_n2929;
assign 2_n904 = 2_n10750 | 2_n10422;
assign 2_n7904 = 2_n4674 | 2_n9188;
assign 2_n1778 = ~(2_n10839 | 2_n5248);
assign 2_n9632 = ~2_n2428;
assign 2_n4589 = ~(2_n1632 | 2_n11730);
assign 2_n1907 = 2_n8217 & 2_n10941;
assign 2_n12934 = ~(2_n11327 ^ 2_n7000);
assign 2_n10936 = 2_n12119 | 2_n8957;
assign 2_n816 = 2_n2099 | 2_n3224;
assign 2_n12228 = ~(2_n4435 ^ 2_n10033);
assign 2_n9046 = ~2_n11230;
assign 2_n3592 = ~(2_n6282 ^ 2_n12279);
assign 2_n6667 = ~2_n7563;
assign 2_n7958 = ~(2_n7873 ^ 2_n9771);
assign 2_n5489 = 2_n7998 | 2_n4153;
assign 2_n5660 = 2_n5886 & 2_n770;
assign 2_n8487 = 2_n6275 & 2_n3907;
assign 2_n2690 = ~(2_n8429 ^ 2_n7326);
assign 2_n242 = ~2_n8526;
assign 2_n10234 = ~2_n3246;
assign 2_n10110 = 2_n11490 & 2_n1919;
assign 2_n6344 = ~(2_n8194 ^ 2_n4035);
assign 2_n8477 = 2_n11153 & 2_n7270;
assign 2_n7551 = 2_n6577 | 2_n6169;
assign 2_n4134 = 2_n6053 | 2_n5830;
assign 2_n9805 = ~(2_n12496 ^ 2_n5124);
assign 2_n8669 = 2_n11005 | 2_n11297;
assign 2_n5219 = 2_n2099 | 2_n8655;
assign 2_n12386 = 2_n8959 | 2_n6169;
assign 2_n5633 = ~(2_n6350 ^ 2_n11412);
assign 2_n7717 = ~2_n1882;
assign 2_n10034 = ~(2_n8395 ^ 2_n7863);
assign 2_n4535 = 2_n10157 | 2_n4642;
assign 2_n6955 = 2_n5054 & 2_n6300;
assign 2_n3294 = ~(2_n8520 ^ 2_n7815);
assign 2_n3212 = 2_n11234 & 2_n12522;
assign 2_n10166 = ~(2_n2688 ^ 2_n5315);
assign 2_n291 = 2_n8194 & 2_n4035;
assign 2_n6779 = ~(2_n5975 | 2_n2362);
assign 2_n2254 = 2_n1799 | 2_n8544;
assign 2_n2005 = ~(2_n9304 ^ 2_n549);
assign 2_n9329 = 2_n6544 | 2_n6422;
assign 2_n7176 = 2_n12119 | 2_n9586;
assign 2_n9047 = ~(2_n11934 ^ 2_n4273);
assign 2_n12760 = 2_n6941 & 2_n6764;
assign 2_n7249 = ~(2_n10153 ^ 2_n8437);
assign 2_n918 = ~2_n9270;
assign 2_n5516 = 2_n603 | 2_n12688;
assign 2_n1145 = 2_n1696 | 2_n3102;
assign 2_n8414 = ~2_n4928;
assign 2_n10340 = 2_n10732 | 2_n476;
assign 2_n8499 = 2_n9373 | 2_n5502;
assign 2_n2962 = 2_n6408 & 2_n5787;
assign 2_n6959 = ~(2_n8141 | 2_n12804);
assign 2_n5993 = 2_n7108 & 2_n12164;
assign 2_n5547 = 2_n8411 & 2_n4596;
assign 2_n4837 = 2_n5398 | 2_n3248;
assign 2_n2618 = 2_n4911 | 2_n7341;
assign 2_n11437 = ~(2_n2138 ^ 2_n723);
assign 2_n11220 = 2_n585 & 2_n4670;
assign 2_n8795 = ~(2_n9514 | 2_n3751);
assign 2_n154 = ~(2_n9017 | 2_n8199);
assign 2_n2943 = 2_n6709 & 2_n8356;
assign 2_n8587 = 2_n11556 | 2_n6173;
assign 2_n11247 = 2_n3155 & 2_n7213;
assign 2_n10594 = 2_n4116 | 2_n7188;
assign 2_n8431 = 2_n11933 | 2_n11322;
assign 2_n8270 = ~(2_n6520 ^ 2_n5991);
assign 2_n5756 = ~(2_n6517 ^ 2_n10246);
assign 2_n9215 = 2_n8221 & 2_n11268;
assign 2_n10754 = 2_n3617 | 2_n5468;
assign 2_n6227 = 2_n11060 | 2_n11247;
assign 2_n8814 = 2_n10157 | 2_n1509;
assign 2_n11243 = 2_n9777 & 2_n9309;
assign 2_n10471 = ~(2_n8518 | 2_n5697);
assign 2_n9375 = ~(2_n7758 ^ 2_n793);
assign 2_n7182 = ~(2_n4395 ^ 2_n7923);
assign 2_n9808 = 2_n6142 & 2_n830;
assign 2_n3988 = ~(2_n9197 ^ 2_n12110);
assign 2_n12776 = 2_n2564 & 2_n2585;
assign 2_n2292 = ~2_n3817;
assign 2_n877 = ~(2_n12178 ^ 2_n1481);
assign 2_n5384 = 2_n5355 | 2_n1546;
assign 2_n461 = ~(2_n2885 ^ 2_n9715);
assign 2_n8250 = ~(2_n359 ^ 2_n9357);
assign 2_n130 = ~2_n2512;
assign 2_n1713 = ~(2_n2365 ^ 2_n932);
assign 2_n39 = ~(2_n10152 ^ 2_n1693);
assign 2_n3775 = 2_n3992 & 2_n11876;
assign 2_n536 = ~(2_n5206 ^ 2_n2311);
assign 2_n2443 = ~(2_n2481 ^ 2_n3504);
assign 2_n480 = ~(2_n6039 ^ 2_n10488);
assign 2_n11409 = ~(2_n11076 ^ 2_n7142);
assign 2_n11852 = ~2_n4990;
assign 2_n3092 = ~(2_n10844 ^ 2_n8471);
assign 2_n10891 = ~2_n9385;
assign 2_n5675 = ~(2_n7268 ^ 2_n1767);
assign 2_n5783 = 2_n8336 & 2_n9640;
assign 2_n3722 = ~(2_n11352 ^ 2_n12265);
assign 2_n3152 = ~2_n187;
assign 2_n2065 = ~(2_n3665 | 2_n2452);
assign 2_n654 = ~(2_n8282 ^ 2_n12298);
assign 2_n3737 = ~(2_n11405 | 2_n9285);
assign 2_n8061 = ~(2_n1031 ^ 2_n9297);
assign 2_n2526 = ~(2_n10414 ^ 2_n10369);
assign 2_n7311 = 2_n10339 | 2_n12535;
assign 2_n10537 = ~(2_n4829 ^ 2_n11301);
assign 2_n7327 = 2_n2217 | 2_n4527;
assign 2_n2692 = ~(2_n7835 | 2_n8885);
assign 2_n6830 = ~(2_n3108 ^ 2_n6610);
assign 2_n354 = 2_n636 | 2_n6513;
assign 2_n836 = ~2_n5418;
assign 2_n4080 = ~2_n5841;
assign 2_n10386 = ~2_n7205;
assign 2_n8243 = 2_n2792 & 2_n5060;
assign 2_n2830 = ~2_n4017;
assign 2_n2750 = 2_n6475 | 2_n10867;
assign 2_n7852 = ~(2_n3826 ^ 2_n2613);
assign 2_n4072 = ~(2_n6556 ^ 2_n6007);
assign 2_n7724 = ~(2_n11128 | 2_n558);
assign 2_n10614 = 2_n6914 | 2_n4447;
assign 2_n26 = ~2_n7922;
assign 2_n4577 = ~(2_n985 ^ 2_n5558);
assign 2_n11405 = 2_n3324 | 2_n9521;
assign 2_n6901 = 2_n9792 | 2_n7554;
assign 2_n2407 = ~(2_n1844 | 2_n6094);
assign 2_n4824 = 2_n11567 & 2_n4209;
assign 2_n4594 = ~(2_n5001 ^ 2_n6787);
assign 2_n9866 = ~(2_n2329 ^ 2_n8000);
assign 2_n9758 = 2_n12155 | 2_n6473;
assign 2_n5989 = 2_n10835 | 2_n4875;
assign 2_n9687 = 2_n9529 | 2_n7950;
assign 2_n7601 = ~2_n1905;
assign 2_n1274 = ~(2_n10790 ^ 2_n11235);
assign 2_n12244 = 2_n982 & 2_n8230;
assign 2_n1749 = 2_n10129 | 2_n11946;
assign 2_n10308 = 2_n4238 & 2_n6304;
assign 2_n11583 = ~(2_n1459 ^ 2_n1984);
assign 2_n1771 = ~(2_n961 ^ 2_n1359);
assign 2_n2023 = ~2_n8410;
assign 2_n12547 = 2_n8309 & 2_n10441;
assign 2_n6605 = ~(2_n8412 ^ 2_n3429);
assign 2_n2649 = 2_n10874 & 2_n1300;
assign 2_n5551 = 2_n8229 & 2_n1276;
assign 2_n2911 = ~(2_n4442 | 2_n4110);
assign 2_n7668 = 2_n137 & 2_n7610;
assign 2_n3621 = ~2_n4520;
assign 2_n8447 = ~(2_n4357 ^ 2_n10299);
assign 2_n4109 = ~(2_n240 ^ 2_n1076);
assign 2_n10140 = ~(2_n5044 ^ 2_n7639);
assign 2_n6310 = 2_n10750 | 2_n12446;
assign 2_n12509 = ~(2_n7599 | 2_n8910);
assign 2_n4272 = ~(2_n2304 ^ 2_n4839);
assign 2_n8201 = ~2_n11363;
assign 2_n6570 = ~(2_n12055 ^ 2_n8246);
assign 2_n2486 = ~(2_n2838 ^ 2_n6164);
assign 2_n72 = ~(2_n10015 ^ 2_n12517);
assign 2_n316 = ~2_n985;
assign 2_n2715 = ~2_n10443;
assign 2_n11218 = ~(2_n9453 | 2_n9646);
assign 2_n888 = 2_n610 & 2_n469;
assign 2_n12585 = ~2_n11784;
assign 2_n9440 = 2_n399 & 2_n7949;
assign 2_n8349 = 2_n1960 & 2_n1019;
assign 2_n4376 = ~2_n10974;
assign 2_n4417 = ~(2_n12432 ^ 2_n6162);
assign 2_n712 = ~(2_n644 ^ 2_n9966);
assign 2_n8185 = ~2_n6935;
assign 2_n6083 = ~(2_n8481 ^ 2_n1048);
assign 2_n2006 = 2_n10893 & 2_n9121;
assign 2_n6237 = 2_n9373 | 2_n4474;
assign 2_n10487 = 2_n2456 | 2_n12754;
assign 2_n6559 = 2_n4079 & 2_n150;
assign 2_n1788 = ~(2_n6607 | 2_n10753);
assign 2_n7027 = 2_n10750 | 2_n12535;
assign 2_n2613 = ~(2_n685 ^ 2_n12191);
assign 2_n5638 = ~2_n1637;
assign 2_n9229 = ~(2_n11171 ^ 2_n5712);
assign 2_n9916 = 2_n5794 & 2_n4340;
assign 2_n5400 = 2_n10057 & 2_n5822;
assign 2_n11036 = 2_n11958 | 2_n11122;
assign 2_n12129 = ~2_n3467;
assign 2_n4313 = 2_n7301 | 2_n10158;
assign 2_n3110 = 2_n9616 | 2_n5262;
assign 2_n1156 = 2_n2973 | 2_n9613;
assign 2_n6201 = ~(2_n12180 ^ 2_n4558);
assign 2_n3819 = ~2_n10414;
assign 2_n1910 = 2_n5404 | 2_n6823;
assign 2_n6672 = 2_n11801 | 2_n10413;
assign 2_n5836 = 2_n4628 | 2_n2964;
assign 2_n11553 = 2_n10899 & 2_n7532;
assign 2_n11591 = 2_n11887 | 2_n4913;
assign 2_n10923 = 2_n6481 & 2_n7437;
assign 2_n7231 = 2_n2012 & 2_n11497;
assign 2_n11972 = ~(2_n3067 ^ 2_n1793);
assign 2_n11042 = 2_n6945 & 2_n423;
assign 2_n6220 = ~(2_n6585 ^ 2_n12534);
assign 2_n11573 = ~2_n3027;
assign 2_n2330 = ~(2_n10498 ^ 2_n7857);
assign 2_n11328 = 2_n5780 | 2_n960;
assign 2_n6108 = 2_n1621 | 2_n1331;
assign 2_n8977 = 2_n9784 | 2_n6920;
assign 2_n7477 = 2_n4567 & 2_n9960;
assign 2_n12622 = 2_n6577 | 2_n11820;
assign 2_n5070 = ~(2_n3716 | 2_n3586);
assign 2_n6908 = 2_n7167 & 2_n2477;
assign 2_n4605 = ~(2_n12231 ^ 2_n5041);
assign 2_n7431 = ~2_n12166;
assign 2_n6097 = ~(2_n7073 ^ 2_n9628);
assign 2_n4945 = ~2_n4851;
assign 2_n5115 = ~(2_n6497 ^ 2_n10554);
assign 2_n4927 = ~(2_n5368 ^ 2_n11651);
assign 2_n11906 = ~(2_n4388 ^ 2_n4898);
assign 2_n7679 = 2_n7643 & 2_n913;
assign 2_n7840 = 2_n1854 & 2_n4620;
assign 2_n11400 = ~(2_n3089 ^ 2_n3692);
assign 2_n6314 = ~2_n9444;
assign 2_n6063 = ~(2_n8902 ^ 2_n12784);
assign 2_n1408 = 2_n9394 & 2_n6789;
assign 2_n10117 = 2_n12833 | 2_n984;
assign 2_n6810 = 2_n4724 | 2_n7896;
assign 2_n8393 = 2_n11923 | 2_n8285;
assign 2_n11964 = 2_n10740 & 2_n5703;
assign 2_n10849 = 2_n3930 | 2_n4483;
assign 2_n11099 = 2_n1911 & 2_n1004;
assign 2_n3197 = ~2_n9131;
assign 2_n7543 = ~(2_n7127 ^ 2_n7774);
assign 2_n786 = ~(2_n95 | 2_n6792);
assign 2_n392 = 2_n9170 | 2_n7424;
assign 2_n12874 = 2_n9005 | 2_n1608;
assign 2_n3709 = 2_n969 & 2_n5046;
assign 2_n4866 = 2_n9373 | 2_n4527;
assign 2_n10692 = 2_n5860 & 2_n5760;
assign 2_n11951 = ~(2_n7502 ^ 2_n12213);
assign 2_n1368 = 2_n566 | 2_n5656;
assign 2_n6669 = 2_n5355 | 2_n4775;
assign 2_n4362 = ~(2_n2458 ^ 2_n12238);
assign 2_n9009 = 2_n9343 | 2_n12425;
assign 2_n2101 = 2_n2448 | 2_n3799;
assign 2_n10068 = ~2_n11653;
assign 2_n6504 = 2_n3625 & 2_n9031;
assign 2_n11128 = 2_n11433 | 2_n5540;
assign 2_n7 = ~(2_n3476 ^ 2_n1193);
assign 2_n12087 = 2_n12069 & 2_n2558;
assign 2_n12240 = ~(2_n12318 ^ 2_n6900);
assign 2_n1596 = ~(2_n10374 ^ 2_n3898);
assign 2_n5899 = 2_n2913 ^ 2_n368;
assign 2_n11336 = 2_n7043 & 2_n7190;
assign 2_n3162 = 2_n10983 & 2_n2817;
assign 2_n3309 = 2_n11036 & 2_n8030;
assign 2_n1140 = ~(2_n11692 | 2_n12484);
assign 2_n8693 = ~(2_n9348 ^ 2_n7667);
assign 2_n1946 = 2_n10196 | 2_n4642;
assign 2_n8766 = 2_n9389 | 2_n1738;
assign 2_n4718 = 2_n1041 & 2_n11364;
assign 2_n4569 = ~(2_n7726 ^ 2_n5533);
assign 2_n7626 = 2_n7874 | 2_n12918;
assign 2_n8890 = ~2_n3163;
assign 2_n5162 = ~(2_n10960 ^ 2_n10315);
assign 2_n1619 = 2_n8743 & 2_n9505;
assign 2_n4018 = 2_n9884 | 2_n3411;
assign 2_n682 = 2_n8785 & 2_n6021;
assign 2_n10123 = ~2_n6001;
assign 2_n3106 = 2_n11070 & 2_n4599;
assign 2_n5027 = 2_n8412 | 2_n3521;
assign 2_n10874 = 2_n5530 | 2_n1163;
assign 2_n11702 = ~(2_n3397 ^ 2_n6382);
assign 2_n5341 = 2_n994 | 2_n1546;
assign 2_n2740 = ~2_n9298;
assign 2_n1722 = 2_n11900 & 2_n8871;
assign 2_n2426 = ~(2_n7376 ^ 2_n7465);
assign 2_n7306 = 2_n8428 | 2_n11896;
assign 2_n9515 = ~(2_n7585 ^ 2_n8283);
assign 2_n9401 = 2_n2917 | 2_n2465;
assign 2_n6008 = ~(2_n6051 ^ 2_n9635);
assign 2_n12485 = ~(2_n3712 | 2_n9805);
assign 2_n6210 = ~(2_n1884 ^ 2_n3312);
assign 2_n12735 = ~2_n6254;
assign 2_n8075 = ~(2_n6506 ^ 2_n12372);
assign 2_n8737 = 2_n11026 | 2_n1047;
assign 2_n10949 = ~(2_n948 ^ 2_n7482);
assign 2_n6159 = 2_n8418 & 2_n11472;
assign 2_n10734 = 2_n5215 & 2_n8095;
assign 2_n11802 = 2_n9970 & 2_n2224;
assign 2_n6303 = 2_n4604 | 2_n5220;
assign 2_n6205 = 2_n6995 & 2_n2405;
assign 2_n3721 = ~2_n12757;
assign 2_n6013 = 2_n8192 | 2_n10193;
assign 2_n6807 = ~(2_n10610 ^ 2_n1855);
assign 2_n4479 = ~(2_n2109 | 2_n6274);
assign 2_n4342 = ~2_n11491;
assign 2_n3265 = 2_n12119 | 2_n12735;
assign 2_n12549 = 2_n4674 | 2_n826;
assign 2_n12816 = ~2_n12709;
assign 2_n2298 = 2_n5573 & 2_n7618;
assign 2_n2951 = ~(2_n7732 | 2_n11246);
assign 2_n2302 = ~2_n6015;
assign 2_n9705 = 2_n10396 | 2_n11491;
assign 2_n2789 = ~(2_n9515 ^ 2_n2825);
assign 2_n12920 = 2_n7283 | 2_n7389;
assign 2_n1990 = 2_n3743 | 2_n1476;
assign 2_n9814 = 2_n395 ^ 2_n8479;
assign 2_n7322 = 2_n2217 | 2_n8285;
assign 2_n5917 = 2_n1446 | 2_n10492;
assign 2_n8077 = ~(2_n574 ^ 2_n6427);
assign 2_n6656 = ~2_n4273;
assign 2_n580 = ~2_n6242;
assign 2_n11054 = ~(2_n8836 ^ 2_n11376);
assign 2_n4502 = 2_n2272 & 2_n10258;
assign 2_n3284 = 2_n8026 | 2_n11122;
assign 2_n987 = 2_n7617 & 2_n9667;
assign 2_n2753 = 2_n12644 | 2_n265;
assign 2_n1247 = 2_n6145 | 2_n3647;
assign 2_n6195 = 2_n7495 | 2_n3911;
assign 2_n4613 = 2_n10196 | 2_n1047;
assign 2_n8614 = ~(2_n11984 ^ 2_n6460);
assign 2_n6949 = ~(2_n10155 ^ 2_n2140);
assign 2_n6855 = 2_n3627 & 2_n7265;
assign 2_n8241 = 2_n7965 & 2_n10848;
assign 2_n8490 = ~(2_n478 ^ 2_n12475);
assign 2_n1308 = 2_n686 | 2_n3903;
assign 2_n7191 = ~(2_n11343 | 2_n3499);
assign 2_n10851 = 2_n11557 ^ 2_n12360;
assign 2_n12195 = 2_n3746 | 2_n995;
assign 2_n11683 = ~(2_n9987 | 2_n2361);
assign 2_n6664 = ~(2_n8786 ^ 2_n2419);
assign 2_n3741 = 2_n5151 & 2_n11670;
assign 2_n6172 = 2_n4666 | 2_n10863;
assign 2_n10522 = 2_n6770 & 2_n4370;
assign 2_n8438 = ~2_n12123;
assign 2_n9314 = 2_n880 | 2_n11758;
assign 2_n6940 = ~(2_n1448 | 2_n5789);
assign 2_n9381 = ~(2_n11148 ^ 2_n12140);
assign 2_n7120 = 2_n2017 | 2_n2883;
assign 2_n8273 = 2_n2456 | 2_n12735;
assign 2_n3505 = 2_n10091 & 2_n100;
assign 2_n12870 = 2_n1717 & 2_n3813;
assign 2_n9878 = ~2_n6294;
assign 2_n1129 = ~2_n1689;
assign 2_n9859 = 2_n636 | 2_n2964;
assign 2_n7788 = 2_n2584 | 2_n9258;
assign 2_n6047 = ~(2_n6033 | 2_n214);
assign 2_n2843 = ~2_n9465;
assign 2_n7224 = 2_n7236 & 2_n8028;
assign 2_n8 = 2_n3156 & 2_n12008;
assign 2_n2902 = ~(2_n11187 ^ 2_n7671);
assign 2_n1515 = 2_n12007 | 2_n2328;
assign 2_n9764 = 2_n8552 | 2_n8648;
assign 2_n2268 = 2_n9389 | 2_n3911;
assign 2_n10585 = 2_n1051 | 2_n7876;
assign 2_n4869 = ~2_n10399;
assign 2_n11620 = ~(2_n7898 ^ 2_n2622);
assign 2_n4855 = ~(2_n7911 | 2_n5323);
assign 2_n12900 = ~2_n85;
assign 2_n5456 = 2_n5575 | 2_n6197;
assign 2_n3532 = ~(2_n1409 ^ 2_n12780);
assign 2_n2327 = 2_n418 | 2_n7924;
assign 2_n2306 = ~(2_n4781 | 2_n138);
assign 2_n2970 = 2_n6237 | 2_n9526;
assign 2_n7092 = ~(2_n11405 ^ 2_n11665);
assign 2_n1865 = 2_n12361 | 2_n11896;
assign 2_n7888 = 2_n5838 | 2_n10892;
assign 2_n7645 = 2_n1890 | 2_n3343;
assign 2_n4591 = 2_n5765 | 2_n609;
assign 2_n5804 = ~(2_n8191 ^ 2_n11176);
assign 2_n166 = ~2_n12778;
assign 2_n8965 = ~(2_n10467 ^ 2_n12288);
assign 2_n11975 = 2_n11668 & 2_n7538;
assign 2_n12203 = 2_n191 | 2_n4775;
assign 2_n228 = ~(2_n3075 ^ 2_n314);
assign 2_n11648 = 2_n11856 & 2_n6911;
assign 2_n2521 = 2_n3026 | 2_n3896;
assign 2_n3976 = 2_n5355 | 2_n8524;
assign 2_n1002 = 2_n6894 & 2_n7105;
assign 2_n3516 = 2_n7044 & 2_n10185;
assign 2_n2008 = 2_n12361 | 2_n2232;
assign 2_n6416 = ~2_n10466;
assign 2_n12749 = 2_n4994 & 2_n2980;
assign 2_n6261 = 2_n8214 | 2_n10857;
assign 2_n5984 = 2_n6718 | 2_n7921;
assign 2_n546 = ~(2_n10019 | 2_n11667);
assign 2_n5753 = 2_n3153 | 2_n6982;
assign 2_n4233 = ~(2_n8378 ^ 2_n8061);
assign 2_n5482 = 2_n2067 & 2_n12568;
assign 2_n1855 = ~(2_n4856 ^ 2_n3348);
assign 2_n6755 = ~2_n2903;
assign 2_n3960 = ~(2_n8934 ^ 2_n10460);
assign 2_n3410 = 2_n444 & 2_n12829;
assign 2_n9506 = 2_n3620 & 2_n5718;
assign 2_n3449 = 2_n3820 | 2_n5258;
assign 2_n2121 = 2_n11080 & 2_n12597;
assign 2_n9316 = ~(2_n10059 ^ 2_n10827);
assign 2_n10265 = 2_n2226 & 2_n8819;
assign 2_n7385 = ~(2_n12827 ^ 2_n1674);
assign 2_n14 = ~(2_n4994 ^ 2_n2980);
assign 2_n1436 = 2_n4644 & 2_n11624;
assign 2_n12371 = ~2_n1322;
assign 2_n6863 = ~2_n3354;
assign 2_n3905 = 2_n10347 | 2_n12182;
assign 2_n6391 = 2_n5016 | 2_n12202;
assign 2_n5441 = 2_n2456 | 2_n3924;
assign 2_n9625 = ~2_n8370;
assign 2_n11530 = ~(2_n11286 ^ 2_n12320);
assign 2_n3388 = 2_n5404 & 2_n6823;
assign 2_n9588 = 2_n3050 | 2_n11524;
assign 2_n4821 = ~(2_n7247 ^ 2_n199);
assign 2_n9207 = ~(2_n1350 | 2_n1912);
assign 2_n1071 = 2_n7536 | 2_n1191;
assign 2_n1754 = ~(2_n646 | 2_n494);
assign 2_n858 = ~(2_n1746 ^ 2_n2404);
assign 2_n10320 = ~(2_n11490 | 2_n1919);
assign 2_n3233 = ~(2_n5969 | 2_n1313);
assign 2_n10139 = 2_n2217 | 2_n4642;
assign 2_n11391 = ~(2_n6801 ^ 2_n6011);
assign 2_n177 = ~2_n9289;
assign 2_n133 = 2_n10108 | 2_n5497;
assign 2_n11763 = ~(2_n10587 ^ 2_n12727);
assign 2_n7298 = 2_n602 | 2_n10024;
assign 2_n6333 = ~(2_n8445 ^ 2_n9766);
assign 2_n871 = ~(2_n11712 ^ 2_n9574);
assign 2_n6129 = ~(2_n3335 ^ 2_n9062);
assign 2_n8645 = 2_n2244 | 2_n9402;
assign 2_n62 = 2_n12324 & 2_n2736;
assign 2_n3143 = ~(2_n12653 ^ 2_n5229);
assign 2_n11244 = 2_n2033 | 2_n8014;
assign 2_n4432 = 2_n989 | 2_n4400;
assign 2_n10838 = 2_n10157 | 2_n8830;
assign 2_n644 = ~(2_n8116 ^ 2_n9576);
assign 2_n7002 = 2_n2652 & 2_n3518;
assign 2_n12084 = ~(2_n2899 ^ 2_n4182);
assign 2_n2098 = ~(2_n1907 | 2_n12566);
assign 2_n5576 = ~(2_n5584 ^ 2_n5672);
assign 2_n4173 = 2_n2874 | 2_n9587;
assign 2_n8575 = 2_n12698 | 2_n2298;
assign 2_n446 = ~(2_n9363 ^ 2_n4807);
assign 2_n11012 = ~(2_n10810 ^ 2_n4144);
assign 2_n7532 = 2_n884 | 2_n3639;
assign 2_n11891 = ~2_n6439;
assign 2_n9895 = 2_n3344 | 2_n11086;
assign 2_n3382 = 2_n10343 | 2_n9535;
assign 2_n10940 = 2_n9170 | 2_n2358;
assign 2_n5367 = ~(2_n5720 | 2_n6565);
assign 2_n10501 = 2_n9908 & 2_n12874;
assign 2_n1947 = 2_n7417 | 2_n2149;
assign 2_n4452 = ~2_n623;
assign 2_n9373 = ~2_n6358;
assign 2_n2759 = ~(2_n1154 ^ 2_n10804);
assign 2_n10997 = 2_n8187 | 2_n12328;
assign 2_n9665 = 2_n432 & 2_n9549;
assign 2_n12739 = 2_n3096 | 2_n3903;
assign 2_n6753 = ~(2_n8580 ^ 2_n6223);
assign 2_n9293 = ~(2_n6938 ^ 2_n5481);
assign 2_n8950 = ~(2_n880 ^ 2_n5131);
assign 2_n5528 = 2_n12953 | 2_n4878;
assign 2_n1483 = 2_n11719 | 2_n3911;
assign 2_n12102 = ~2_n5901;
assign 2_n11161 = 2_n6320 | 2_n2821;
assign 2_n1727 = 2_n2539 | 2_n5910;
assign 2_n6184 = 2_n9101 | 2_n9516;
assign 2_n11853 = ~(2_n12200 ^ 2_n12789);
assign 2_n10132 = 2_n515 & 2_n5941;
assign 2_n6217 = ~(2_n4791 ^ 2_n5925);
assign 2_n1269 = ~(2_n10631 ^ 2_n2095);
assign 2_n55 = 2_n4984 & 2_n9153;
assign 2_n2070 = ~(2_n646 ^ 2_n11540);
assign 2_n6782 = 2_n4498 | 2_n7424;
assign 2_n9819 = ~(2_n10648 ^ 2_n8179);
assign 2_n2611 = ~(2_n1680 ^ 2_n31);
assign 2_n335 = 2_n4948 & 2_n12021;
assign 2_n8462 = 2_n3262 | 2_n4072;
assign 2_n11916 = ~(2_n2713 | 2_n6937);
assign 2_n5136 = 2_n3617 | 2_n8740;
assign 2_n7268 = ~(2_n9460 ^ 2_n6159);
assign 2_n12690 = 2_n9274 & 2_n10814;
assign 2_n4352 = ~(2_n10279 | 2_n9855);
assign 2_n11977 = ~2_n8051;
assign 2_n10313 = ~(2_n7650 ^ 2_n3);
assign 2_n524 = ~2_n2481;
assign 2_n3107 = 2_n1898 | 2_n3673;
assign 2_n9807 = 2_n11838 | 2_n7344;
assign 2_n11722 = 2_n2976 | 2_n11495;
assign 2_n4248 = ~(2_n10255 ^ 2_n696);
assign 2_n8700 = 2_n1598 & 2_n5564;
assign 2_n1885 = ~(2_n11535 ^ 2_n8403);
assign 2_n1048 = 2_n3933 & 2_n3406;
assign 2_n3648 = 2_n9176 | 2_n12409;
assign 2_n4285 = ~2_n4414;
assign 2_n11368 = 2_n7709 | 2_n9160;
assign 2_n4349 = ~(2_n2321 ^ 2_n5704);
assign 2_n6473 = 2_n3820 | 2_n9521;
assign 2_n6752 = ~(2_n2319 | 2_n10252);
assign 2_n2574 = ~2_n2761;
assign 2_n199 = ~(2_n11517 ^ 2_n5883);
assign 2_n5749 = 2_n4274 | 2_n11810;
assign 2_n6107 = ~(2_n3533 ^ 2_n1284);
assign 2_n11681 = 2_n4957 & 2_n7771;
assign 2_n10084 = ~(2_n4747 ^ 2_n2534);
assign 2_n4544 = 2_n11026 | 2_n28;
assign 2_n591 = 2_n11142 & 2_n10187;
assign 2_n2894 = 2_n10738 & 2_n3150;
assign 2_n12718 = ~(2_n9853 ^ 2_n1831);
assign 2_n2493 = 2_n4657 | 2_n3971;
assign 2_n4884 = ~2_n7224;
assign 2_n3427 = ~(2_n1007 | 2_n10410);
assign 2_n4350 = ~2_n1485;
assign 2_n6841 = ~(2_n9518 ^ 2_n5197);
assign 2_n8326 = ~2_n9591;
assign 2_n8565 = ~(2_n3915 ^ 2_n11558);
assign 2_n10237 = 2_n7906 & 2_n9794;
assign 2_n8911 = ~(2_n457 ^ 2_n8086);
assign 2_n6074 = 2_n9170 | 2_n4400;
assign 2_n5739 = 2_n191 | 2_n2358;
assign 2_n585 = 2_n6877 & 2_n3602;
assign 2_n7157 = ~(2_n2352 ^ 2_n2643);
assign 2_n10970 = ~(2_n1433 ^ 2_n5853);
assign 2_n4716 = 2_n2099 | 2_n8648;
assign 2_n6498 = 2_n12503 | 2_n4527;
assign 2_n12260 = ~(2_n8608 | 2_n8160);
assign 2_n11542 = 2_n11641 | 2_n12379;
assign 2_n6793 = 2_n306 | 2_n40;
assign 2_n10252 = 2_n11923 | 2_n5502;
assign 2_n3165 = 2_n4352 | 2_n1388;
assign 2_n4001 = 2_n989 | 2_n7703;
assign 2_n1691 = ~2_n972;
assign 2_n2792 = 2_n5235 | 2_n433;
assign 2_n12155 = 2_n6718 | 2_n4875;
assign 2_n12289 = 2_n2099 | 2_n6071;
assign 2_n4311 = ~(2_n4224 | 2_n7290);
assign 2_n7941 = 2_n11324 & 2_n12756;
assign 2_n9379 = 2_n191 | 2_n510;
assign 2_n2333 = ~(2_n8499 ^ 2_n7574);
assign 2_n2095 = ~(2_n3184 ^ 2_n11333);
assign 2_n7707 = 2_n4183 | 2_n3886;
assign 2_n12885 = ~(2_n6174 ^ 2_n1885);
assign 2_n6066 = 2_n3743 | 2_n1047;
assign 2_n11703 = ~(2_n11713 ^ 2_n4695);
assign 2_n3945 = 2_n10845 & 2_n8426;
assign 2_n4825 = ~2_n12398;
assign 2_n9659 = ~2_n10160;
assign 2_n5447 = ~(2_n11835 ^ 2_n2891);
assign 2_n8666 = ~(2_n8439 ^ 2_n8953);
assign 2_n8845 = ~2_n12455;
assign 2_n10978 = ~(2_n5739 ^ 2_n10241);
assign 2_n4409 = ~(2_n7509 ^ 2_n9998);
assign 2_n8180 = 2_n7709 | 2_n2020;
assign 2_n2217 = ~2_n11222;
assign 2_n10279 = ~2_n2569;
assign 2_n5047 = ~(2_n10434 ^ 2_n1362);
assign 2_n8188 = ~(2_n8290 | 2_n5095);
assign 2_n12332 = 2_n2456 | 2_n8259;
assign 2_n10295 = 2_n5209 & 2_n10312;
assign 2_n8635 = ~(2_n6393 | 2_n1343);
assign 2_n3950 = ~2_n6369;
assign 2_n9970 = 2_n8002 | 2_n8934;
assign 2_n9660 = ~(2_n4726 ^ 2_n8098);
assign 2_n2257 = 2_n2097 & 2_n3792;
assign 2_n5665 = 2_n9400 & 2_n7354;
assign 2_n12721 = 2_n320 | 2_n8869;
assign 2_n11433 = ~2_n10678;
assign 2_n5420 = ~(2_n9980 | 2_n1587);
assign 2_n5355 = ~2_n5305;
assign 2_n7711 = ~(2_n9701 ^ 2_n6861);
assign 2_n2828 = ~(2_n12336 ^ 2_n3572);
assign 2_n12662 = ~2_n3513;
assign 2_n9762 = ~(2_n2590 | 2_n1544);
assign 2_n5204 = 2_n7449 | 2_n1047;
assign 2_n7869 = 2_n5765 | 2_n7506;
assign 2_n4413 = 2_n7391 | 2_n510;
assign 2_n4078 = 2_n597 | 2_n5896;
assign 2_n6827 = 2_n3383 | 2_n2297;
assign 2_n3746 = ~2_n6776;
assign 2_n6723 = 2_n11893 & 2_n9885;
assign 2_n11772 = ~(2_n8374 ^ 2_n3113);
assign 2_n11268 = ~(2_n2100 ^ 2_n4650);
assign 2_n10866 = ~(2_n8847 ^ 2_n9356);
assign 2_n5500 = ~(2_n12856 ^ 2_n7698);
assign 2_n1437 = ~2_n10753;
assign 2_n10355 = 2_n4535 & 2_n501;
assign 2_n9310 = ~(2_n1435 ^ 2_n9040);
assign 2_n5734 = ~(2_n8954 ^ 2_n6852);
assign 2_n9026 = ~(2_n5405 ^ 2_n8025);
assign 2_n9934 = ~2_n5849;
assign 2_n2017 = 2_n10614 & 2_n7859;
assign 2_n3809 = ~(2_n3968 ^ 2_n11016);
assign 2_n4695 = ~(2_n11419 | 2_n12685);
assign 2_n246 = 2_n3240 | 2_n8801;
assign 2_n11593 = 2_n3127 | 2_n10066;
assign 2_n8047 = ~(2_n2308 ^ 2_n10415);
assign 2_n3418 = 2_n12119 | 2_n4249;
assign 2_n4027 = ~(2_n8102 | 2_n5006);
assign 2_n11366 = 2_n1791 & 2_n5344;
assign 2_n11422 = ~2_n4651;
assign 2_n2291 = ~(2_n11540 | 2_n1736);
assign 2_n7331 = 2_n3746 | 2_n5538;
assign 2_n2213 = 2_n10835 | 2_n5258;
assign 2_n10349 = ~(2_n5567 | 2_n7187);
assign 2_n4510 = 2_n5765 | 2_n5258;
assign 2_n4795 = ~(2_n9982 ^ 2_n10923);
assign 2_n11144 = ~2_n9676;
assign 2_n8851 = 2_n5331 & 2_n5645;
assign 2_n7810 = ~2_n8672;
assign 2_n10423 = 2_n3838 | 2_n5529;
assign 2_n8249 = ~(2_n6331 ^ 2_n1383);
assign 2_n10850 = 2_n804 & 2_n3714;
assign 2_n11179 = 2_n9170 | 2_n10066;
assign 2_n4390 = 2_n7283 | 2_n12328;
assign 2_n11575 = 2_n1114 & 2_n12030;
assign 2_n2404 = ~(2_n5475 ^ 2_n1395);
assign 2_n6811 = ~2_n3821;
assign 2_n12294 = ~2_n12248;
assign 2_n4820 = ~(2_n810 | 2_n2058);
assign 2_n4719 = ~2_n2150;
assign 2_n4152 = 2_n6910 | 2_n2668;
assign 2_n7274 = ~2_n3601;
assign 2_n4038 = 2_n12340 | 2_n1385;
assign 2_n1061 = 2_n1699 | 2_n9586;
assign 2_n3893 = ~(2_n4119 ^ 2_n6949);
assign 2_n2367 = ~2_n45;
assign 2_n6481 = 2_n5730 | 2_n10407;
assign 2_n10715 = 2_n1402 & 2_n5866;
assign 2_n7123 = 2_n6784 & 2_n2103;
assign 2_n127 = 2_n5832 | 2_n6531;
assign 2_n2077 = ~(2_n5269 ^ 2_n1535);
assign 2_n2138 = ~(2_n1694 ^ 2_n3727);
assign 2_n11159 = ~2_n7954;
assign 2_n4003 = ~(2_n8799 ^ 2_n4811);
assign 2_n8703 = ~2_n3588;
assign 2_n9466 = 2_n7732 & 2_n11246;
assign 2_n4653 = ~2_n6342;
assign 2_n3395 = 2_n10196 | 2_n5258;
assign 2_n759 = ~(2_n4036 ^ 2_n9503);
assign 2_n10044 = ~(2_n9610 ^ 2_n8172);
assign 2_n1560 = 2_n11552 | 2_n795;
assign 2_n12817 = 2_n3747 & 2_n12249;
assign 2_n2680 = 2_n12705 & 2_n2879;
assign 2_n608 = ~2_n7039;
assign 2_n5601 = 2_n11923 | 2_n9160;
assign 2_n1565 = 2_n4750 | 2_n4652;
assign 2_n6726 = ~2_n8130;
assign 2_n1577 = 2_n949 & 2_n5917;
assign 2_n2899 = 2_n5355 | 2_n130;
assign 2_n5990 = 2_n910 | 2_n9852;
assign 2_n12475 = ~(2_n4460 ^ 2_n5272);
assign 2_n4232 = 2_n2099 | 2_n8957;
assign 2_n70 = ~(2_n3758 ^ 2_n7031);
assign 2_n168 = 2_n11305 | 2_n10501;
assign 2_n1377 = 2_n6451 | 2_n2894;
assign 2_n8265 = ~2_n1922;
assign 2_n1254 = 2_n8094 | 2_n12865;
assign 2_n5395 = 2_n4469 | 2_n1428;
assign 2_n2506 = ~2_n6092;
assign 2_n6268 = 2_n2099 | 2_n5781;
assign 2_n7021 = 2_n8552 | 2_n530;
assign 2_n3184 = ~(2_n5221 ^ 2_n8032);
assign 2_n4735 = ~2_n8049;
assign 2_n1823 = ~(2_n7942 ^ 2_n2484);
assign 2_n12340 = ~2_n6813;
assign 2_n12043 = 2_n11093 | 2_n9211;
assign 2_n10600 = ~2_n3705;
assign 2_n6266 = ~(2_n6779 ^ 2_n4801);
assign 2_n1601 = 2_n5397 | 2_n9174;
assign 2_n9582 = ~2_n3350;
assign 2_n4671 = ~(2_n3579 | 2_n4342);
assign 2_n12542 = 2_n2660 & 2_n10205;
assign 2_n8367 = ~2_n1201;
assign 2_n86 = ~(2_n10964 ^ 2_n1311);
assign 2_n7785 = ~2_n3968;
assign 2_n6965 = ~(2_n12502 | 2_n11276);
assign 2_n519 = 2_n1539 | 2_n11827;
assign 2_n2133 = 2_n2400 & 2_n2705;
assign 2_n3512 = 2_n4997 & 2_n3937;
assign 2_n7348 = 2_n752 | 2_n12274;
assign 2_n1196 = ~(2_n2858 | 2_n10188);
assign 2_n6792 = ~(2_n2373 ^ 2_n3696);
assign 2_n9360 = 2_n9826 & 2_n3979;
assign 2_n6076 = ~2_n42;
assign 2_n9394 = 2_n7037 | 2_n3232;
assign 2_n12157 = 2_n7391 | 2_n1162;
assign 2_n9458 = ~2_n11086;
assign 2_n3979 = ~2_n6771;
assign 2_n5519 = 2_n8197 & 2_n1098;
assign 2_n2979 = 2_n9170 | 2_n1079;
assign 2_n8685 = ~2_n2632;
assign 2_n9165 = 2_n1277 & 2_n4946;
assign 2_n10152 = 2_n9377 & 2_n6523;
assign 2_n5897 = ~2_n10558;
assign 2_n3925 = ~(2_n8447 | 2_n203);
assign 2_n9200 = ~(2_n5231 ^ 2_n7537);
assign 2_n10387 = ~(2_n12064 ^ 2_n11987);
assign 2_n1545 = ~(2_n5859 ^ 2_n12038);
assign 2_n6317 = 2_n3257 & 2_n4096;
assign 2_n6887 = ~2_n3894;
assign 2_n8313 = 2_n10835 | 2_n8643;
assign 2_n2256 = ~2_n2007;
assign 2_n995 = ~2_n9189;
assign 2_n3360 = ~(2_n8260 ^ 2_n12065);
assign 2_n245 = ~(2_n8362 ^ 2_n12232);
assign 2_n1359 = 2_n2524 & 2_n11431;
assign 2_n3189 = ~(2_n538 ^ 2_n8465);
assign 2_n11253 = 2_n11509 | 2_n6804;
assign 2_n4890 = ~(2_n2176 | 2_n8516);
assign 2_n12601 = ~2_n2336;
assign 2_n11774 = ~(2_n7912 ^ 2_n4136);
assign 2_n4620 = ~(2_n6479 ^ 2_n877);
assign 2_n12292 = ~(2_n6370 ^ 2_n5408);
assign 2_n10175 = ~(2_n5746 ^ 2_n7472);
assign 2_n6183 = ~(2_n7330 | 2_n11630);
assign 2_n8998 = ~(2_n4823 ^ 2_n7140);
assign 2_n1633 = ~2_n10138;
assign 2_n823 = ~(2_n9438 ^ 2_n8744);
assign 2_n9135 = ~(2_n1249 ^ 2_n7963);
assign 2_n12667 = ~(2_n4392 ^ 2_n11710);
assign 2_n5242 = 2_n5809 | 2_n3224;
assign 2_n1080 = ~(2_n4732 ^ 2_n8773);
assign 2_n4297 = 2_n8567 | 2_n10536;
assign 2_n5127 = ~2_n847;
assign 2_n9974 = 2_n8187 | 2_n8524;
assign 2_n5614 = 2_n12648 & 2_n521;
assign 2_n320 = 2_n6577 | 2_n7952;
assign 2_n12168 = 2_n3271 & 2_n6179;
assign 2_n7324 = 2_n7116 | 2_n3421;
assign 2_n7233 = 2_n2226 & 2_n8595;
assign 2_n9600 = 2_n10180 | 2_n4234;
assign 2_n6719 = 2_n2605 | 2_n11921;
assign 2_n730 = ~(2_n2032 ^ 2_n1939);
assign 2_n1387 = ~2_n3491;
assign 2_n2435 = ~(2_n888 | 2_n8328);
assign 2_n4168 = 2_n6687 & 2_n7265;
assign 2_n7801 = 2_n3746 | 2_n2232;
assign 2_n12930 = ~2_n84;
assign 2_n9662 = 2_n9645 & 2_n12301;
assign 2_n75 = ~(2_n5100 ^ 2_n6264);
assign 2_n3531 = 2_n3870 & 2_n7120;
assign 2_n7288 = 2_n5494 | 2_n5401;
assign 2_n11341 = ~2_n6222;
assign 2_n9648 = 2_n12361 | 2_n3903;
assign 2_n7957 = ~(2_n4968 ^ 2_n6992);
assign 2_n5746 = 2_n9306 & 2_n4078;
assign 2_n8551 = 2_n11466 | 2_n8222;
assign 2_n1540 = ~(2_n12823 ^ 2_n1143);
assign 2_n1849 = ~(2_n6759 ^ 2_n11160);
assign 2_n10767 = ~2_n11325;
assign 2_n5611 = 2_n11723 & 2_n12821;
assign 2_n3412 = 2_n3020 & 2_n1355;
assign 2_n10114 = 2_n4589 | 2_n9128;
assign 2_n140 = ~2_n7452;
assign 2_n6839 = ~2_n1702;
assign 2_n11080 = 2_n752 | 2_n12899;
assign 2_n6865 = ~(2_n9915 ^ 2_n1496);
assign 2_n8496 = ~2_n12788;
assign 2_n8762 = ~(2_n6686 | 2_n5407);
assign 2_n5817 = 2_n12248 | 2_n7723;
assign 2_n2373 = ~(2_n6308 ^ 2_n5352);
assign 2_n264 = ~2_n11997;
assign 2_n12423 = 2_n12119 | 2_n1932;
assign 2_n10205 = 2_n6095 | 2_n781;
assign 2_n5164 = 2_n3658 & 2_n10207;
assign 2_n12110 = 2_n12397 & 2_n11508;
assign 2_n2862 = 2_n8552 | 2_n4913;
assign 2_n5472 = ~(2_n8406 ^ 2_n3783);
assign 2_n10238 = ~(2_n11312 ^ 2_n8586);
assign 2_n9158 = 2_n2516 | 2_n11559;
assign 2_n4226 = 2_n6527 ^ 2_n10214;
assign 2_n12606 = 2_n3279 & 2_n6871;
assign 2_n4836 = ~(2_n12552 ^ 2_n8115);
assign 2_n7894 = ~2_n10152;
assign 2_n782 = 2_n11476 | 2_n1125;
assign 2_n8498 = ~(2_n7861 | 2_n5327);
assign 2_n1953 = ~(2_n12224 ^ 2_n5268);
assign 2_n4165 = ~(2_n8081 ^ 2_n11340);
assign 2_n4628 = ~2_n8476;
assign 2_n11236 = 2_n1937 | 2_n5012;
assign 2_n9323 = 2_n4784 | 2_n3419;
assign 2_n3273 = 2_n10108 | 2_n1162;
assign 2_n11198 = ~(2_n7627 ^ 2_n12128);
assign 2_n10696 = 2_n9389 | 2_n561;
assign 2_n1181 = 2_n8127 | 2_n5497;
assign 2_n781 = ~(2_n10567 ^ 2_n2771);
assign 2_n911 = ~(2_n11756 ^ 2_n10459);
assign 2_n3021 = 2_n9373 | 2_n2020;
assign 2_n890 = 2_n1811 | 2_n829;
assign 2_n11347 = ~2_n7440;
assign 2_n6763 = 2_n7901 | 2_n5701;
assign 2_n7430 = ~(2_n9146 ^ 2_n2453);
assign 2_n10592 = ~(2_n9565 ^ 2_n6469);
assign 2_n6639 = ~(2_n251 ^ 2_n8980);
assign 2_n11828 = ~(2_n9310 ^ 2_n10043);
assign 2_n11819 = ~(2_n6442 ^ 2_n3462);
assign 2_n3999 = ~(2_n10887 | 2_n323);
assign 2_n5061 = 2_n5780 & 2_n960;
assign 2_n8743 = 2_n8759 & 2_n2024;
assign 2_n5344 = 2_n2813 & 2_n7613;
assign 2_n2259 = ~2_n5694;
assign 2_n4511 = 2_n9367 | 2_n7471;
assign 2_n1729 = ~2_n11508;
assign 2_n457 = ~(2_n10656 ^ 2_n12903);
assign 2_n6245 = 2_n8207 | 2_n8650;
assign 2_n8925 = 2_n3845 & 2_n10733;
assign 2_n5830 = ~(2_n8468 ^ 2_n8278);
assign 2_n9616 = 2_n10750 | 2_n5326;
assign 2_n3848 = 2_n5219 | 2_n4926;
assign 2_n11595 = 2_n8026 | 2_n9971;
assign 2_n2686 = 2_n2099 | 2_n8644;
assign 2_n1964 = ~(2_n5404 ^ 2_n6823);
assign 2_n5646 = 2_n5594 & 2_n11095;
assign 2_n8199 = 2_n7457 & 2_n872;
assign 2_n7606 = ~(2_n463 | 2_n625);
assign 2_n12468 = 2_n488 | 2_n10691;
assign 2_n8852 = 2_n6718 | 2_n8285;
assign 2_n2971 = ~2_n8656;
assign 2_n7147 = ~2_n8266;
assign 2_n8324 = ~(2_n2467 ^ 2_n311);
assign 2_n10656 = 2_n12853 | 2_n826;
assign 2_n247 = ~(2_n4429 ^ 2_n4659);
assign 2_n6412 = ~2_n3472;
assign 2_n11894 = 2_n9837 | 2_n6529;
assign 2_n10515 = 2_n5681 & 2_n10646;
assign 2_n7134 = 2_n9688 & 2_n8446;
assign 2_n7101 = 2_n6577 | 2_n11775;
assign 2_n2704 = 2_n3743 | 2_n3451;
assign 2_n11017 = 2_n8127 | 2_n10066;
assign 2_n7839 = ~2_n10510;
assign 2_n10615 = ~(2_n8009 ^ 2_n4744);
assign 2_n10179 = 2_n12800 | 2_n9418;
assign 2_n12185 = ~(2_n9391 | 2_n5302);
assign 2_n680 = 2_n1557 & 2_n7030;
assign 2_n11089 = ~(2_n5780 ^ 2_n960);
assign 2_n1321 = 2_n1051 | 2_n6197;
assign 2_n6068 = 2_n11822 & 2_n8382;
assign 2_n7745 = 2_n10745 | 2_n12072;
assign 2_n11751 = 2_n8959 | 2_n8768;
assign 2_n2111 = 2_n8959 | 2_n7558;
assign 2_n8118 = 2_n7391 | 2_n7424;
assign 2_n2477 = ~(2_n9360 ^ 2_n4260);
assign 2_n1491 = 2_n8550 & 2_n10934;
assign 2_n6475 = 2_n8187 | 2_n12843;
assign 2_n4373 = 2_n2217 | 2_n609;
assign 2_n4789 = 2_n8395 | 2_n10588;
assign 2_n7950 = 2_n11110 & 2_n10794;
assign 2_n7812 = ~(2_n7429 ^ 2_n4344);
assign 2_n6923 = ~(2_n10128 | 2_n6714);
assign 2_n7625 = 2_n10636 & 2_n367;
assign 2_n2157 = 2_n7992 & 2_n8569;
assign 2_n8310 = 2_n8552 | 2_n12080;
assign 2_n11053 = ~(2_n3987 ^ 2_n11636);
assign 2_n6896 = 2_n10466 & 2_n2678;
assign 2_n8283 = ~(2_n12046 ^ 2_n1287);
assign 2_n11829 = 2_n8778 | 2_n12718;
assign 2_n8550 = 2_n2217 | 2_n5759;
assign 2_n11287 = ~2_n9720;
assign 2_n11657 = 2_n4205 | 2_n10817;
assign 2_n8513 = ~2_n917;
assign 2_n12092 = 2_n9661 & 2_n5130;
assign 2_n4658 = 2_n4788 & 2_n9620;
assign 2_n12187 = ~2_n5622;
assign 2_n4035 = 2_n10879 | 2_n11746;
assign 2_n517 = 2_n4179 | 2_n8266;
assign 2_n548 = 2_n9370 | 2_n8524;
assign 2_n4030 = ~(2_n7276 ^ 2_n5974);
assign 2_n9319 = ~(2_n285 ^ 2_n180);
assign 2_n5755 = 2_n1070 & 2_n4306;
assign 2_n5868 = ~(2_n3433 | 2_n1722);
assign 2_n10078 = 2_n3836 | 2_n12371;
assign 2_n9129 = ~(2_n5384 ^ 2_n12652);
assign 2_n11043 = 2_n1382 & 2_n11657;
assign 2_n4145 = 2_n10545 & 2_n1512;
assign 2_n6414 = 2_n12361 | 2_n2815;
assign 2_n6395 = 2_n10212 & 2_n907;
assign 2_n4704 = ~(2_n1760 | 2_n2859);
assign 2_n6336 = ~(2_n12579 | 2_n6506);
assign 2_n4747 = 2_n10224 & 2_n11452;
assign 2_n11004 = ~(2_n805 | 2_n7656);
assign 2_n3579 = ~(2_n3753 ^ 2_n2941);
assign 2_n6156 = ~(2_n12870 ^ 2_n440);
assign 2_n9861 = ~(2_n2947 | 2_n940);
assign 2_n5269 = ~(2_n10608 ^ 2_n5950);
assign 2_n9481 = 2_n4628 | 2_n12446;
assign 2_n5088 = ~2_n11533;
assign 2_n12052 = 2_n8187 | 2_n1915;
assign 2_n11665 = ~(2_n10148 ^ 2_n7996);
assign 2_n5731 = ~(2_n9626 ^ 2_n1597);
assign 2_n3459 = ~(2_n867 ^ 2_n4731);
assign 2_n334 = 2_n9878 | 2_n3224;
assign 2_n7692 = ~(2_n7151 ^ 2_n1501);
assign 2_n6039 = 2_n12673 & 2_n10440;
assign 2_n5125 = 2_n9688 | 2_n8446;
assign 2_n5439 = ~2_n3130;
assign 2_n9686 = ~(2_n12123 ^ 2_n9490);
assign 2_n1741 = ~2_n7920;
assign 2_n11274 = 2_n10124 & 2_n455;
assign 2_n9113 = ~(2_n4420 ^ 2_n1603);
assign 2_n492 = 2_n9370 | 2_n4242;
assign 2_n3920 = 2_n2845 & 2_n4177;
assign 2_n5556 = ~(2_n10667 ^ 2_n8317);
assign 2_n8251 = 2_n8187 | 2_n6389;
assign 2_n89 = 2_n3363 | 2_n5509;
assign 2_n7814 = ~(2_n4524 ^ 2_n10068);
assign 2_n6734 = 2_n8193 & 2_n5002;
assign 2_n9876 = 2_n4894 | 2_n36;
assign 2_n1608 = ~(2_n9787 ^ 2_n1904);
assign 2_n10539 = ~(2_n1705 ^ 2_n12251);
assign 2_n8577 = ~2_n9550;
assign 2_n5259 = ~(2_n1112 ^ 2_n8588);
assign 2_n10057 = 2_n8870 | 2_n8655;
assign 2_n2897 = ~(2_n7505 ^ 2_n3049);
assign 2_n3128 = ~(2_n9339 ^ 2_n4763);
assign 2_n10184 = ~(2_n11232 | 2_n8064);
assign 2_n10041 = ~(2_n349 ^ 2_n3520);
assign 2_n6812 = ~(2_n8522 | 2_n3882);
assign 2_n6370 = 2_n12119 | 2_n12535;
assign 2_n9820 = ~(2_n1264 ^ 2_n4776);
assign 2_n4785 = 2_n9379 | 2_n1356;
assign 2_n851 = ~(2_n12327 ^ 2_n1660);
assign 2_n5231 = 2_n8583 | 2_n4875;
assign 2_n812 = ~(2_n6175 ^ 2_n11006);
assign 2_n1562 = ~2_n3928;
assign 2_n2285 = 2_n752 | 2_n9741;
assign 2_n11245 = 2_n11026 | 2_n3606;
assign 2_n11010 = ~(2_n7243 ^ 2_n2460);
assign 2_n7095 = ~(2_n8904 ^ 2_n12193);
assign 2_n9651 = 2_n4911 | 2_n5497;
assign 2_n11948 = 2_n9029 & 2_n2615;
assign 2_n6450 = 2_n1016 | 2_n1979;
assign 2_n3375 = ~(2_n12532 ^ 2_n1620);
assign 2_n11896 = ~2_n5105;
assign 2_n7657 = ~2_n1216;
assign 2_n9028 = ~2_n9655;
assign 2_n2073 = ~(2_n4224 ^ 2_n7155);
assign 2_n8830 = ~2_n7294;
assign 2_n689 = ~(2_n1255 ^ 2_n10444);
assign 2_n3948 = ~2_n3519;
assign 2_n12748 = ~2_n11050;
assign 2_n9732 = 2_n3795 | 2_n10294;
assign 2_n4810 = ~(2_n1475 ^ 2_n5414);
assign 2_n6124 = ~2_n1505;
assign 2_n1450 = ~(2_n9089 ^ 2_n11980);
assign 2_n7402 = ~(2_n5832 ^ 2_n6531);
assign 2_n10813 = 2_n681 & 2_n10418;
assign 2_n373 = ~2_n3921;
assign 2_n10115 = ~(2_n1721 ^ 2_n10114);
assign 2_n12649 = ~(2_n7375 ^ 2_n5256);
assign 2_n917 = 2_n7588 & 2_n9543;
assign 2_n6234 = ~2_n5299;
assign 2_n7075 = ~(2_n3337 ^ 2_n3294);
assign 2_n8042 = 2_n3642 & 2_n10963;
assign 2_n5336 = ~(2_n5432 ^ 2_n12292);
assign 2_n11126 = 2_n8835 | 2_n9595;
assign 2_n8958 = 2_n7218 & 2_n4313;
assign 2_n8839 = 2_n11958 | 2_n11410;
assign 2_n3207 = 2_n6635 | 2_n9863;
assign 2_n5393 = 2_n11958 | 2_n3468;
assign 2_n6747 = ~2_n11038;
assign 2_n8972 = ~(2_n9988 | 2_n6332);
assign 2_n6105 = 2_n11953 | 2_n11242;
assign 2_n4741 = ~(2_n3869 ^ 2_n6209);
assign 2_n11419 = ~(2_n6374 | 2_n5757);
assign 2_n6153 = 2_n3096 | 2_n7558;
assign 2_n11822 = 2_n4480 | 2_n7866;
assign 2_n603 = ~(2_n9499 | 2_n17);
assign 2_n1013 = ~(2_n4142 | 2_n4691);
assign 2_n10945 = 2_n6718 | 2_n3606;
assign 2_n2842 = 2_n6786 & 2_n10373;
assign 2_n12261 = 2_n432 | 2_n9549;
assign 2_n3787 = ~(2_n2193 ^ 2_n4708);
assign 2_n3393 = 2_n5547 | 2_n5810;
assign 2_n8520 = ~(2_n3883 ^ 2_n5807);
assign 2_n10769 = ~(2_n1390 ^ 2_n1292);
assign 2_n6021 = 2_n6772 | 2_n1596;
assign 2_n7701 = 2_n5285 & 2_n6902;
assign 2_n3991 = 2_n7657 & 2_n9315;
assign 2_n2225 = ~(2_n9164 | 2_n6802);
assign 2_n5784 = ~(2_n12799 ^ 2_n12253);
assign 2_n1956 = 2_n11627 & 2_n7205;
assign 2_n575 = ~(2_n102 | 2_n5875);
assign 2_n873 = 2_n12090 | 2_n4871;
assign 2_n12588 = 2_n5319 & 2_n9763;
assign 2_n12790 = 2_n12115 & 2_n1761;
assign 2_n11740 = 2_n1419 | 2_n9216;
assign 2_n214 = 2_n2947 & 2_n940;
assign 2_n841 = ~(2_n5370 ^ 2_n339);
assign 2_n5967 = 2_n11026 | 2_n8643;
assign 2_n6657 = ~(2_n3412 | 2_n12407);
assign 2_n9212 = 2_n12941 | 2_n1624;
assign 2_n1663 = 2_n10219 | 2_n7477;
assign 2_n5475 = ~(2_n11264 ^ 2_n3744);
assign 2_n11466 = ~(2_n3198 | 2_n12772);
assign 2_n6851 = 2_n1900 | 2_n9556;
assign 2_n12698 = 2_n5247 & 2_n9020;
assign 2_n7993 = 2_n7236 & 2_n9111;
assign 2_n9851 = ~(2_n6313 ^ 2_n498);
assign 2_n3045 = ~(2_n12950 | 2_n1381);
assign 2_n2072 = 2_n97 | 2_n2129;
assign 2_n4975 = ~(2_n4138 ^ 2_n9929);
assign 2_n4724 = 2_n9101 & 2_n9516;
assign 2_n1654 = 2_n11719 | 2_n1455;
assign 2_n2948 = ~(2_n2075 | 2_n6972);
assign 2_n100 = ~(2_n11184 ^ 2_n11018);
assign 2_n10449 = ~2_n6997;
assign 2_n5856 = ~(2_n5324 ^ 2_n518);
assign 2_n4108 = 2_n2069 & 2_n10458;
assign 2_n2766 = ~2_n5627;
assign 2_n10751 = 2_n1200 | 2_n1482;
assign 2_n9822 = 2_n3700 & 2_n5294;
assign 2_n10904 = 2_n6867 & 2_n187;
assign 2_n1694 = ~(2_n11929 ^ 2_n6253);
assign 2_n4966 = 2_n11319 | 2_n4310;
assign 2_n3492 = ~(2_n5605 ^ 2_n3745);
assign 2_n9765 = 2_n8645 & 2_n9594;
assign 2_n3404 = ~(2_n6576 ^ 2_n5150);
assign 2_n4177 = ~2_n6705;
assign 2_n1646 = 2_n8959 | 2_n11896;
assign 2_n12954 = ~2_n11708;
assign 2_n9090 = 2_n5945 | 2_n11775;
assign 2_n11060 = 2_n7283 | 2_n1546;
assign 2_n8916 = 2_n10339 | 2_n5468;
assign 2_n10136 = 2_n7409 | 2_n1868;
assign 2_n419 = 2_n12038 | 2_n1913;
assign 2_n5888 = ~(2_n6070 ^ 2_n56);
assign 2_n12771 = ~2_n9111;
assign 2_n11676 = ~(2_n6190 ^ 2_n11658);
assign 2_n6476 = ~(2_n4647 ^ 2_n11236);
assign 2_n3840 = 2_n12750 & 2_n376;
assign 2_n7440 = 2_n5916 & 2_n6785;
assign 2_n5885 = 2_n114 | 2_n6169;
assign 2_n12343 = 2_n4189 & 2_n4370;
assign 2_n8501 = ~(2_n737 ^ 2_n6132);
assign 2_n8445 = 2_n1316 | 2_n6898;
assign 2_n2805 = 2_n12135 & 2_n1380;
assign 2_n9366 = ~(2_n1275 ^ 2_n8240);
assign 2_n4437 = 2_n8823 & 2_n2049;
assign 2_n10913 = ~(2_n10857 ^ 2_n8385);
assign 2_n8073 = ~2_n6498;
assign 2_n278 = ~(2_n458 ^ 2_n2992);
assign 2_n8068 = ~(2_n3340 ^ 2_n4228);
assign 2_n10392 = 2_n8839 | 2_n10927;
assign 2_n11283 = ~(2_n5213 | 2_n12602);
assign 2_n5512 = 2_n807 | 2_n2232;
assign 2_n2315 = ~(2_n1359 | 2_n6658);
assign 2_n9197 = ~(2_n3076 ^ 2_n7402);
assign 2_n6080 = 2_n2541 & 2_n10427;
assign 2_n1457 = ~(2_n663 ^ 2_n9039);
assign 2_n11899 = ~(2_n8165 | 2_n297);
assign 2_n3571 = ~2_n1426;
assign 2_n1484 = 2_n2967 | 2_n10447;
assign 2_n2408 = 2_n8759 & 2_n3602;
assign 2_n3406 = 2_n9538 | 2_n4064;
assign 2_n7209 = 2_n1741 | 2_n8715;
assign 2_n9049 = 2_n12388 & 2_n2492;
assign 2_n10634 = ~2_n5336;
assign 2_n11851 = 2_n7283 | 2_n2358;
assign 2_n11723 = ~(2_n1518 ^ 2_n3536);
assign 2_n8940 = 2_n10247 | 2_n5597;
assign 2_n9067 = 2_n4255 & 2_n10411;
assign 2_n5853 = 2_n686 | 2_n7952;
assign 2_n1195 = ~(2_n1043 ^ 2_n4780);
assign 2_n9469 = ~(2_n8752 ^ 2_n9850);
assign 2_n9029 = 2_n4639 | 2_n6140;
assign 2_n7697 = ~(2_n10039 ^ 2_n5591);
assign 2_n7991 = ~(2_n12859 ^ 2_n2652);
assign 2_n4607 = ~(2_n8266 ^ 2_n2102);
assign 2_n6042 = ~2_n5533;
assign 2_n3266 = 2_n3573 | 2_n10624;
assign 2_n2867 = 2_n11059 | 2_n12300;
assign 2_n6134 = 2_n10626 & 2_n12317;
assign 2_n2344 = 2_n621 & 2_n6844;
assign 2_n6362 = ~2_n1541;
assign 2_n10593 = ~(2_n5603 ^ 2_n11345);
assign 2_n10677 = 2_n2534 & 2_n4747;
assign 2_n8430 = 2_n1465 | 2_n6272;
assign 2_n7406 = 2_n8136 | 2_n4879;
assign 2_n9449 = ~(2_n3546 | 2_n9225);
assign 2_n1634 = 2_n5685 & 2_n5658;
assign 2_n12466 = 2_n11717 & 2_n9120;
assign 2_n9657 = 2_n7974 & 2_n9532;
assign 2_n11248 = 2_n11460 ^ 2_n39;
assign 2_n5923 = 2_n5214 | 2_n2616;
assign 2_n3587 = ~(2_n8334 | 2_n6234);
assign 2_n9431 = 2_n10799 | 2_n917;
assign 2_n6296 = 2_n10142 | 2_n8735;
assign 2_n2668 = ~2_n8121;
assign 2_n11487 = 2_n422 | 2_n12482;
assign 2_n10716 = ~2_n146;
assign 2_n1454 = 2_n1627 & 2_n5813;
assign 2_n5656 = 2_n2700 & 2_n3268;
assign 2_n10709 = ~2_n9708;
assign 2_n5126 = 2_n4451 & 2_n1852;
assign 2_n7059 = ~(2_n1477 | 2_n11049);
assign 2_n5605 = 2_n5530 | 2_n2964;
assign 2_n7729 = 2_n11305 & 2_n10501;
assign 2_n1031 = ~(2_n11687 ^ 2_n6599);
assign 2_n7738 = ~(2_n12107 ^ 2_n6632);
assign 2_n12651 = ~(2_n9985 ^ 2_n5777);
assign 2_n7908 = 2_n2564 & 2_n7265;
assign 2_n4425 = ~2_n2973;
assign 2_n8618 = 2_n3887 & 2_n3583;
assign 2_n5737 = 2_n6226 | 2_n7666;
assign 2_n47 = ~2_n2085;
assign 2_n6943 = 2_n7015 | 2_n9959;
assign 2_n12654 = ~(2_n8510 ^ 2_n8274);
assign 2_n9273 = 2_n5341 | 2_n11947;
assign 2_n1233 = ~2_n11280;
assign 2_n8403 = ~(2_n7299 ^ 2_n2239);
assign 2_n12253 = 2_n5945 | 2_n7952;
assign 2_n10332 = ~2_n6379;
assign 2_n5413 = 2_n9233 & 2_n8244;
assign 2_n12710 = ~(2_n2014 ^ 2_n12259);
assign 2_n2465 = 2_n7376 & 2_n7465;
assign 2_n12823 = 2_n8738 | 2_n9568;
assign 2_n5777 = 2_n9507 | 2_n1602;
assign 2_n8861 = ~(2_n431 ^ 2_n8546);
assign 2_n11237 = ~(2_n531 ^ 2_n1338);
assign 2_n5895 = 2_n9400 & 2_n12145;
assign 2_n711 = ~2_n12776;
assign 2_n5572 = ~(2_n4458 ^ 2_n9783);
assign 2_n74 = 2_n6465 & 2_n4645;
assign 2_n4281 = 2_n2699 & 2_n1618;
assign 2_n7635 = ~(2_n11932 ^ 2_n8841);
assign 2_n7851 = 2_n7839 | 2_n2232;
assign 2_n5399 = 2_n3878 & 2_n1565;
assign 2_n5591 = ~(2_n10291 | 2_n11261);
assign 2_n5122 = ~(2_n10699 ^ 2_n5490);
assign 2_n2726 = 2_n11026 | 2_n9521;
assign 2_n5848 = 2_n12237 | 2_n12080;
assign 2_n8527 = ~(2_n8149 | 2_n5517);
assign 2_n3483 = ~(2_n121 ^ 2_n1389);
assign 2_n668 = 2_n6339 | 2_n3157;
assign 2_n1679 = 2_n5673 | 2_n8756;
assign 2_n4240 = ~(2_n9322 ^ 2_n3475);
assign 2_n11796 = 2_n11153 & 2_n159;
assign 2_n5761 = 2_n3127 | 2_n4400;
assign 2_n3653 = 2_n8583 | 2_n795;
assign 2_n2860 = 2_n5340 & 2_n11957;
assign 2_n756 = 2_n8273 & 2_n4909;
assign 2_n9237 = ~2_n4105;
assign 2_n1957 = ~2_n11358;
assign 2_n4444 = ~(2_n8535 ^ 2_n2410);
assign 2_n12165 = 2_n4778 | 2_n8655;
assign 2_n2535 = 2_n9880 & 2_n10801;
assign 2_n116 = 2_n12195 | 2_n4622;
assign 2_n9073 = 2_n12186 | 2_n7876;
assign 2_n7479 = 2_n10748 | 2_n2039;
assign 2_n7702 = 2_n8046 | 2_n4497;
assign 2_n6970 = ~(2_n4206 ^ 2_n4303);
assign 2_n3322 = ~2_n7267;
assign 2_n8973 = 2_n6482 & 2_n4586;
assign 2_n399 = 2_n5754 & 2_n1983;
assign 2_n11306 = ~(2_n11718 ^ 2_n350);
assign 2_n5301 = 2_n8342 & 2_n4051;
assign 2_n5930 = 2_n4812 & 2_n2573;
assign 2_n4906 = 2_n1220 & 2_n12621;
assign 2_n7363 = 2_n4289 | 2_n3035;
assign 2_n7397 = ~2_n5003;
assign 2_n2959 = ~2_n12178;
assign 2_n2038 = ~(2_n583 ^ 2_n6202);
assign 2_n3877 = ~(2_n7416 ^ 2_n950);
assign 2_n4174 = ~(2_n1916 ^ 2_n655);
assign 2_n8448 = ~(2_n4158 | 2_n4407);
assign 2_n9268 = ~(2_n5728 | 2_n6335);
assign 2_n4761 = ~(2_n10361 ^ 2_n12246);
assign 2_n12474 = ~(2_n862 | 2_n8121);
assign 2_n12031 = 2_n2464 & 2_n8595;
assign 2_n1434 = ~(2_n4577 | 2_n10423);
assign 2_n2776 = ~(2_n9832 ^ 2_n8657);
assign 2_n8238 = 2_n6076 & 2_n5169;
assign 2_n7281 = ~(2_n12871 | 2_n5649);
assign 2_n5253 = ~(2_n5109 | 2_n12295);
assign 2_n3217 = ~(2_n12639 ^ 2_n9823);
assign 2_n11805 = 2_n3931 | 2_n9720;
assign 2_n12438 = 2_n4624 & 2_n8281;
assign 2_n12641 = ~(2_n1867 ^ 2_n8734);
assign 2_n2105 = 2_n92 & 2_n4789;
assign 2_n6103 = 2_n10842 | 2_n5823;
assign 2_n7005 = 2_n3382 & 2_n8620;
assign 2_n203 = 2_n1910 & 2_n3114;
assign 2_n8080 = ~(2_n6773 | 2_n9419);
assign 2_n535 = 2_n5771 & 2_n415;
assign 2_n7196 = 2_n4562 & 2_n12689;
assign 2_n12807 = ~(2_n310 ^ 2_n3008);
assign 2_n5929 = ~2_n6136;
assign 2_n4439 = 2_n1345 & 2_n6887;
assign 2_n10598 = 2_n12280 & 2_n2937;
assign 2_n10938 = ~2_n3016;
assign 2_n6795 = 2_n4023 | 2_n1870;
assign 2_n3851 = ~(2_n8894 ^ 2_n11774);
assign 2_n12639 = ~(2_n9936 | 2_n2634);
assign 2_n12486 = ~(2_n7798 | 2_n2194);
assign 2_n9498 = 2_n10862 | 2_n10421;
assign 2_n1268 = ~(2_n5590 ^ 2_n12406);
assign 2_n4251 = ~(2_n8229 ^ 2_n1276);
assign 2_n6529 = 2_n7468 & 2_n271;
assign 2_n11510 = ~(2_n6541 | 2_n1219);
assign 2_n5232 = ~(2_n925 ^ 2_n10714);
assign 2_n7650 = ~(2_n10000 ^ 2_n6912);
assign 2_n11197 = 2_n12775 & 2_n12913;
assign 2_n10062 = ~(2_n2602 ^ 2_n2106);
assign 2_n7433 = 2_n2483 & 2_n4040;
assign 2_n11675 = 2_n7449 | 2_n8285;
assign 2_n7549 = 2_n8583 | 2_n9078;
assign 2_n6236 = ~(2_n10438 ^ 2_n12160);
assign 2_n12518 = 2_n12659 | 2_n6846;
assign 2_n1684 = 2_n3767 | 2_n7600;
assign 2_n2460 = 2_n4693 & 2_n5182;
assign 2_n2009 = ~(2_n7102 ^ 2_n7017);
assign 2_n10262 = ~(2_n12747 ^ 2_n8685);
assign 2_n9187 = ~(2_n9770 ^ 2_n2556);
assign 2_n5531 = 2_n3992 & 2_n10990;
assign 2_n977 = ~(2_n10367 ^ 2_n2164);
assign 2_n190 = 2_n8929 & 2_n11141;
assign 2_n7671 = ~(2_n10711 ^ 2_n6094);
assign 2_n2362 = ~(2_n6886 | 2_n8213);
assign 2_n5161 = ~(2_n9629 ^ 2_n11870);
assign 2_n5995 = 2_n10157 | 2_n9280;
assign 2_n10835 = ~2_n7965;
assign 2_n7240 = 2_n6442 & 2_n10619;
assign 2_n9924 = 2_n2959 & 2_n1481;
assign 2_n2200 = ~(2_n5026 ^ 2_n4539);
assign 2_n641 = ~2_n12071;
assign 2_n6518 = 2_n6718 | 2_n9078;
assign 2_n10695 = ~(2_n6665 ^ 2_n8726);
assign 2_n2782 = 2_n3402 | 2_n3391;
assign 2_n12804 = ~(2_n12433 | 2_n5417);
assign 2_n8122 = ~(2_n12242 ^ 2_n8909);
assign 2_n7369 = 2_n6022 | 2_n8427;
assign 2_n10983 = 2_n9370 | 2_n7424;
assign 2_n12939 = ~(2_n10700 ^ 2_n7435);
assign 2_n7145 = 2_n4498 | 2_n7703;
assign 2_n6041 = ~(2_n4635 | 2_n12369);
assign 2_n777 = ~(2_n3726 | 2_n8031);
assign 2_n12719 = 2_n307 & 2_n3471;
assign 2_n5407 = 2_n8687 | 2_n9521;
assign 2_n788 = ~(2_n10343 ^ 2_n9535);
assign 2_n925 = 2_n8187 | 2_n1079;
assign 2_n5826 = 2_n1205 | 2_n4282;
assign 2_n7842 = ~(2_n12945 ^ 2_n9859);
assign 2_n8370 = 2_n7780 & 2_n8901;
assign 2_n2317 = ~2_n8144;
assign 2_n10858 = ~(2_n10365 ^ 2_n8512);
assign 2_n9574 = ~(2_n8130 ^ 2_n9284);
assign 2_n7921 = ~2_n5814;
assign 2_n4440 = ~(2_n7188 ^ 2_n10807);
assign 2_n2168 = 2_n2326 | 2_n10869;
assign 2_n7911 = ~(2_n11972 ^ 2_n11732);
assign 2_n197 = ~(2_n12012 ^ 2_n3054);
assign 2_n7077 = 2_n9900 | 2_n5063;
assign 2_n5249 = 2_n9844 | 2_n7976;
assign 2_n10163 = 2_n5372 | 2_n4163;
assign 2_n12152 = ~(2_n3188 ^ 2_n5561);
assign 2_n10270 = ~2_n1354;
assign 2_n12936 = 2_n4126 | 2_n12608;
assign 2_n8637 = 2_n10715 | 2_n5316;
assign 2_n4133 = ~(2_n578 ^ 2_n8938);
assign 2_n10911 = 2_n5774 | 2_n10011;
assign 2_n12531 = ~2_n1837;
assign 2_n1495 = 2_n1941 | 2_n7558;
assign 2_n10498 = 2_n5141 & 2_n545;
assign 2_n587 = 2_n505 | 2_n12592;
assign 2_n8411 = 2_n6204 | 2_n11735;
assign 2_n7494 = 2_n5981 & 2_n5661;
assign 2_n5327 = 2_n7476 & 2_n10942;
assign 2_n4059 = ~2_n1097;
assign 2_n12047 = 2_n12297 & 2_n11611;
assign 2_n3417 = ~(2_n8733 | 2_n5632);
assign 2_n12764 = 2_n8476 & 2_n6806;
assign 2_n9492 = 2_n6977 | 2_n995;
assign 2_n81 = ~2_n3205;
assign 2_n4562 = 2_n3746 | 2_n7558;
assign 2_n8275 = ~(2_n8369 ^ 2_n4284);
assign 2_n8629 = ~2_n10231;
assign 2_n2560 = 2_n3352 & 2_n1765;
assign 2_n8418 = 2_n9996 & 2_n6634;
assign 2_n5908 = 2_n7709 | 2_n1509;
assign 2_n6005 = ~(2_n10335 | 2_n2378);
assign 2_n7152 = ~(2_n6003 ^ 2_n2919);
assign 2_n11460 = 2_n10045 & 2_n6345;
assign 2_n1760 = 2_n12067 & 2_n9214;
assign 2_n4944 = ~(2_n7300 | 2_n9252);
assign 2_n10647 = 2_n5465 & 2_n6783;
assign 2_n11067 = ~(2_n2877 ^ 2_n7973);
assign 2_n23 = 2_n1519 & 2_n564;
assign 2_n801 = ~(2_n1207 ^ 2_n10696);
assign 2_n842 = ~(2_n8998 ^ 2_n8575);
assign 2_n10028 = ~(2_n1516 ^ 2_n2181);
assign 2_n10546 = 2_n12023 & 2_n7734;
assign 2_n5356 = ~(2_n12282 ^ 2_n4631);
assign 2_n2547 = ~(2_n12728 ^ 2_n340);
assign 2_n1276 = 2_n636 | 2_n10854;
assign 2_n4033 = ~(2_n10921 | 2_n7522);
assign 2_n240 = 2_n2217 | 2_n9078;
assign 2_n3397 = ~2_n7735;
assign 2_n12626 = 2_n7283 | 2_n6389;
assign 2_n1605 = 2_n8228 | 2_n956;
assign 2_n5053 = 2_n8336 & 2_n7946;
assign 2_n8017 = ~(2_n5280 | 2_n1801);
assign 2_n10009 = ~(2_n3313 ^ 2_n11809);
assign 2_n5209 = 2_n1349 | 2_n8258;
assign 2_n6614 = ~(2_n451 ^ 2_n9502);
assign 2_n8223 = ~(2_n5148 | 2_n6675);
assign 2_n5934 = ~(2_n917 ^ 2_n7262);
assign 2_n12359 = 2_n8074 & 2_n735;
assign 2_n1327 = 2_n6674 & 2_n7075;
assign 2_n5052 = ~(2_n12667 ^ 2_n11737);
assign 2_n2662 = ~(2_n1792 ^ 2_n8636);
assign 2_n7035 = 2_n12503 | 2_n795;
assign 2_n7153 = 2_n8764 | 2_n8918;
assign 2_n9581 = 2_n11473 & 2_n6925;
assign 2_n7201 = ~(2_n4863 ^ 2_n7145);
assign 2_n11269 = ~(2_n9746 | 2_n6586);
assign 2_n2540 = ~(2_n9791 ^ 2_n7905);
assign 2_n3791 = 2_n10142 | 2_n7246;
assign 2_n12421 = 2_n77 & 2_n8056;
assign 2_n5955 = 2_n3605 & 2_n9888;
assign 2_n4315 = ~(2_n2586 ^ 2_n2486);
assign 2_n9219 = 2_n1076 | 2_n3439;
assign 2_n3982 = ~(2_n6597 ^ 2_n6845);
assign 2_n10883 = 2_n2031 & 2_n650;
assign 2_n10950 = ~(2_n9656 ^ 2_n12411);
assign 2_n10282 = 2_n5769 | 2_n7239;
assign 2_n1555 = ~(2_n7838 ^ 2_n9135);
assign 2_n9100 = 2_n11697 | 2_n2985;
assign 2_n6718 = ~2_n8384;
assign 2_n6829 = ~(2_n9508 | 2_n146);
assign 2_n183 = 2_n11958 | 2_n7395;
assign 2_n8825 = ~(2_n6330 ^ 2_n6996);
assign 2_n8813 = 2_n7376 | 2_n7465;
assign 2_n6544 = 2_n9373 | 2_n795;
assign 2_n3798 = ~(2_n12789 | 2_n2355);
assign 2_n1879 = 2_n11433 | 2_n5012;
assign 2_n8687 = ~2_n5857;
assign 2_n9156 = ~(2_n3944 ^ 2_n1719);
assign 2_n3052 = ~(2_n11079 | 2_n3847);
assign 2_n3501 = ~2_n927;
assign 2_n5708 = ~(2_n290 ^ 2_n4551);
assign 2_n8522 = 2_n7778 & 2_n7276;
assign 2_n8837 = ~2_n2921;
assign 2_n7015 = ~2_n6891;
assign 2_n7195 = 2_n10966 | 2_n7447;
assign 2_n9015 = ~2_n5846;
assign 2_n8113 = ~2_n8556;
assign 2_n7799 = ~(2_n10912 ^ 2_n6143);
assign 2_n10555 = 2_n2217 | 2_n11698;
assign 2_n10820 = 2_n4778 | 2_n12080;
assign 2_n9724 = ~2_n6343;
assign 2_n4077 = ~(2_n852 | 2_n8335);
assign 2_n563 = ~2_n8927;
assign 2_n1648 = 2_n3478 & 2_n1104;
assign 2_n10700 = ~(2_n1307 ^ 2_n3239);
assign 2_n9209 = ~(2_n11544 ^ 2_n5944);
assign 2_n855 = 2_n7116 | 2_n9741;
assign 2_n3072 = 2_n636 | 2_n8655;
assign 2_n12387 = ~(2_n4416 ^ 2_n4253);
assign 2_n6197 = ~2_n8595;
assign 2_n7344 = 2_n9066 & 2_n11894;
assign 2_n7365 = 2_n636 | 2_n7928;
assign 2_n9427 = ~(2_n3222 | 2_n12228);
assign 2_n749 = ~(2_n7253 | 2_n12848);
assign 2_n11645 = ~2_n5808;
assign 2_n9374 = 2_n11433 | 2_n995;
assign 2_n10226 = ~2_n8851;
assign 2_n8467 = 2_n8410 | 2_n6101;
assign 2_n10233 = ~(2_n4759 | 2_n1569);
assign 2_n7364 = 2_n6559 & 2_n2977;
assign 2_n785 = 2_n3665 & 2_n2452;
assign 2_n4402 = ~(2_n11591 | 2_n9841);
assign 2_n2987 = 2_n10847 | 2_n12626;
assign 2_n2702 = ~(2_n8381 | 2_n3163);
assign 2_n4273 = ~(2_n10529 ^ 2_n626);
assign 2_n12210 = 2_n5081 & 2_n3953;
assign 2_n10257 = ~2_n3795;
assign 2_n1407 = 2_n4247 & 2_n554;
assign 2_n8082 = ~2_n1408;
assign 2_n10921 = 2_n10947 & 2_n11800;
assign 2_n7618 = 2_n8209 | 2_n160;
assign 2_n9969 = ~(2_n5129 | 2_n11770);
assign 2_n4062 = 2_n6115 & 2_n1566;
assign 2_n11737 = ~(2_n10306 ^ 2_n1042);
assign 2_n5514 = 2_n4296 | 2_n11865;
assign 2_n4494 = ~(2_n5567 ^ 2_n4959);
assign 2_n7156 = 2_n338 | 2_n11885;
assign 2_n8935 = ~(2_n333 ^ 2_n2955);
assign 2_n12001 = 2_n3627 & 2_n9956;
assign 2_n7047 = ~(2_n1726 ^ 2_n3718);
assign 2_n6109 = 2_n7487 & 2_n7752;
assign 2_n8014 = ~(2_n8628 ^ 2_n12625);
assign 2_n12537 = ~(2_n1837 ^ 2_n5565);
assign 2_n12846 = 2_n1699 | 2_n6513;
assign 2_n4999 = ~(2_n1588 ^ 2_n12677);
assign 2_n1853 = ~(2_n3576 ^ 2_n6403);
assign 2_n12196 = ~(2_n3516 | 2_n11845);
assign 2_n889 = ~2_n4697;
assign 2_n7588 = 2_n7758 | 2_n1861;
assign 2_n1721 = ~(2_n6229 ^ 2_n3473);
assign 2_n1723 = 2_n3445 & 2_n10261;
assign 2_n11489 = 2_n10661 & 2_n5276;
assign 2_n12109 = ~(2_n9989 | 2_n10408);
assign 2_n4950 = 2_n7071 | 2_n8338;
assign 2_n8131 = ~(2_n11242 ^ 2_n3597);
assign 2_n2057 = ~(2_n5987 ^ 2_n8723);
assign 2_n10181 = 2_n12335 & 2_n9743;
assign 2_n10804 = 2_n9584 | 2_n4527;
assign 2_n2361 = ~(2_n4564 | 2_n4487);
assign 2_n6931 = 2_n5765 | 2_n3606;
assign 2_n12154 = ~(2_n11219 ^ 2_n4800);
assign 2_n6459 = ~(2_n7267 ^ 2_n11797);
assign 2_n8664 = ~(2_n2855 ^ 2_n8874);
assign 2_n9509 = ~(2_n8208 ^ 2_n5512);
assign 2_n9486 = ~2_n6423;
assign 2_n8630 = 2_n2600 & 2_n12332;
assign 2_n8799 = 2_n9838 & 2_n11645;
assign 2_n11027 = 2_n8489 & 2_n5696;
assign 2_n4287 = 2_n7638 | 2_n7419;
assign 2_n2158 = ~(2_n6896 ^ 2_n7636);
assign 2_n412 = 2_n8584 | 2_n12605;
assign 2_n10165 = ~(2_n6116 ^ 2_n4188);
assign 2_n9010 = 2_n3992 & 2_n6611;
assign 2_n2711 = 2_n12443 | 2_n1734;
assign 2_n12632 = 2_n7397 & 2_n11166;
assign 2_n3823 = 2_n7577 | 2_n5796;
assign 2_n7117 = 2_n6373 | 2_n12771;
assign 2_n4404 = ~(2_n928 ^ 2_n3650);
assign 2_n4135 = 2_n5778 & 2_n1591;
assign 2_n10037 = ~(2_n12057 ^ 2_n654);
assign 2_n404 = 2_n373 | 2_n10191;
assign 2_n11945 = ~(2_n12854 ^ 2_n7589);
assign 2_n8558 = 2_n5951 | 2_n5678;
assign 2_n9272 = ~2_n604;
assign 2_n12357 = ~2_n4190;
assign 2_n3132 = ~(2_n10864 ^ 2_n4198);
assign 2_n4283 = 2_n8428 | 2_n995;
assign 2_n11250 = 2_n8428 | 2_n3468;
assign 2_n8374 = ~(2_n12692 ^ 2_n11882);
assign 2_n2397 = ~(2_n6561 ^ 2_n10705);
assign 2_n3685 = 2_n7393 & 2_n12362;
assign 2_n1728 = 2_n9792 & 2_n7554;
assign 2_n12012 = 2_n740 & 2_n406;
assign 2_n2978 = 2_n5809 | 2_n8740;
assign 2_n972 = 2_n10928 & 2_n3719;
assign 2_n12159 = ~(2_n6405 ^ 2_n7440);
assign 2_n5170 = 2_n3544 & 2_n4715;
assign 2_n10652 = 2_n6718 | 2_n1509;
assign 2_n10896 = 2_n5765 | 2_n1509;
assign 2_n10432 = ~(2_n7457 | 2_n872);
assign 2_n2482 = 2_n12119 | 2_n10311;
assign 2_n1845 = 2_n713 & 2_n96;
assign 2_n8667 = ~(2_n650 ^ 2_n2031);
assign 2_n10376 = ~2_n12880;
assign 2_n11529 = ~(2_n10199 ^ 2_n7637);
assign 2_n3202 = 2_n10750 | 2_n7928;
assign 2_n4931 = 2_n8189 | 2_n5797;
assign 2_n11359 = ~(2_n9697 | 2_n1778);
assign 2_n2745 = ~(2_n5219 ^ 2_n3461);
assign 2_n11135 = ~2_n8467;
assign 2_n6284 = 2_n2659 | 2_n3186;
assign 2_n7023 = 2_n3401 & 2_n1996;
assign 2_n9845 = ~(2_n12760 | 2_n2199);
assign 2_n6447 = ~(2_n7866 ^ 2_n2115);
assign 2_n9966 = ~(2_n9068 ^ 2_n9871);
assign 2_n5936 = 2_n12584 & 2_n5733;
assign 2_n12341 = 2_n8789 & 2_n1733;
assign 2_n10131 = ~(2_n2172 ^ 2_n11897);
assign 2_n11910 = 2_n10750 | 2_n10854;
assign 2_n8986 = ~(2_n8896 | 2_n4710);
assign 2_n5111 = 2_n697 | 2_n1109;
assign 2_n5110 = 2_n12380 & 2_n4985;
assign 2_n931 = ~(2_n269 | 2_n10924);
assign 2_n4104 = ~2_n5652;
assign 2_n5921 = ~(2_n8469 ^ 2_n2617);
assign 2_n8677 = ~(2_n11578 ^ 2_n975);
assign 2_n4399 = ~(2_n12266 ^ 2_n2438);
assign 2_n10771 = 2_n11552 | 2_n4527;
assign 2_n2896 = 2_n9262 | 2_n2020;
assign 2_n5183 = 2_n1339 | 2_n8940;
assign 2_n3213 = ~2_n7993;
assign 2_n10336 = 2_n6358 & 2_n11791;
assign 2_n9778 = 2_n7993 & 2_n5845;
assign 2_n12788 = ~(2_n1520 ^ 2_n8247);
assign 2_n7074 = 2_n7236 & 2_n10848;
assign 2_n6922 = ~2_n12247;
assign 2_n9836 = 2_n5575 | 2_n3421;
assign 2_n1770 = ~(2_n8079 ^ 2_n741);
assign 2_n1453 = ~(2_n9555 ^ 2_n10550);
assign 2_n4791 = 2_n7283 | 2_n7703;
assign 2_n12676 = ~(2_n11287 ^ 2_n11954);
assign 2_n10565 = 2_n6373 | 2_n9160;
assign 2_n6051 = ~(2_n12718 ^ 2_n234);
assign 2_n11072 = ~2_n11783;
assign 2_n11406 = 2_n12361 | 2_n11775;
assign 2_n2682 = 2_n3141 & 2_n4721;
assign 2_n1206 = ~(2_n902 ^ 2_n5829);
assign 2_n8672 = 2_n2941 & 2_n1567;
assign 2_n10765 = ~(2_n11445 ^ 2_n247);
assign 2_n3936 = 2_n11026 | 2_n5502;
assign 2_n6700 = 2_n11607 | 2_n10719;
assign 2_n6423 = ~(2_n7206 ^ 2_n11655);
assign 2_n6918 = ~(2_n6628 ^ 2_n1424);
assign 2_n5197 = ~(2_n8996 ^ 2_n4053);
assign 2_n10103 = 2_n4791 | 2_n5762;
assign 2_n9382 = 2_n4411 & 2_n10007;
assign 2_n3850 = ~(2_n409 ^ 2_n12094);
assign 2_n9031 = 2_n12842 & 2_n5654;
assign 2_n8652 = ~(2_n8979 ^ 2_n4334);
assign 2_n3081 = 2_n6695 | 2_n6006;
assign 2_n1559 = ~2_n2752;
assign 2_n8012 = ~(2_n11366 | 2_n7237);
assign 2_n5672 = ~(2_n12024 | 2_n8821);
assign 2_n8602 = ~(2_n4385 ^ 2_n7266);
assign 2_n1773 = 2_n7540 | 2_n3055;
assign 2_n12730 = 2_n11887 | 2_n7382;
assign 2_n612 = ~(2_n11369 | 2_n2990);
assign 2_n1171 = ~2_n10788;
assign 2_n7624 = ~(2_n5898 | 2_n633);
assign 2_n10396 = ~2_n3579;
assign 2_n7141 = 2_n1784 | 2_n11355;
assign 2_n3570 = 2_n5575 | 2_n3356;
assign 2_n532 = ~(2_n1912 ^ 2_n2546);
assign 2_n5044 = ~2_n1397;
assign 2_n960 = 2_n2987 & 2_n6214;
assign 2_n4924 = ~2_n2180;
assign 2_n12796 = 2_n7316 & 2_n9090;
assign 2_n17 = ~2_n4923;
assign 2_n7332 = ~(2_n225 ^ 2_n8039);
assign 2_n12903 = ~(2_n5441 ^ 2_n1862);
assign 2_n4536 = 2_n2456 | 2_n4818;
assign 2_n1632 = 2_n2532 & 2_n4802;
assign 2_n12884 = ~(2_n5799 ^ 2_n801);
assign 2_n5202 = 2_n6577 | 2_n11410;
assign 2_n12144 = 2_n5530 | 2_n1932;
assign 2_n4815 = 2_n9878 | 2_n9188;
assign 2_n10004 = 2_n10282 & 2_n3409;
assign 2_n12657 = ~(2_n9029 ^ 2_n3500);
assign 2_n2746 = ~(2_n7516 ^ 2_n3809);
assign 2_n11040 = 2_n9241 & 2_n6703;
assign 2_n6981 = 2_n5765 | 2_n11698;
assign 2_n3631 = 2_n4343 | 2_n826;
assign 2_n4911 = ~2_n12705;
assign 2_n3443 = ~(2_n11348 ^ 2_n472);
assign 2_n3286 = 2_n10365 & 2_n10723;
assign 2_n2677 = 2_n5575 | 2_n7425;
assign 2_n9737 = 2_n3325 & 2_n1386;
assign 2_n432 = 2_n2217 | 2_n4875;
assign 2_n8882 = 2_n5915 | 2_n10854;
assign 2_n4316 = ~(2_n1256 | 2_n3254);
assign 2_n12551 = 2_n1403 & 2_n765;
assign 2_n12319 = ~(2_n5965 ^ 2_n169);
assign 2_n12501 = ~2_n2111;
assign 2_n10438 = 2_n7197 | 2_n8069;
assign 2_n12640 = ~2_n3732;
assign 2_n69 = 2_n1438 | 2_n2409;
assign 2_n7961 = 2_n4716 | 2_n7;
assign 2_n9423 = ~(2_n11838 ^ 2_n7344);
assign 2_n3810 = 2_n12237 | 2_n7382;
assign 2_n7945 = 2_n7807 & 2_n1412;
assign 2_n1612 = ~2_n2519;
assign 2_n10356 = 2_n595 | 2_n9449;
assign 2_n12053 = 2_n4059 | 2_n7341;
assign 2_n8452 = 2_n6373 | 2_n9568;
assign 2_n11325 = ~(2_n4771 ^ 2_n5082);
assign 2_n4765 = ~(2_n11961 | 2_n1090);
assign 2_n3967 = 2_n8552 | 2_n826;
assign 2_n1595 = 2_n10180 & 2_n4234;
assign 2_n12130 = ~2_n6725;
assign 2_n964 = 2_n8687 | 2_n9160;
assign 2_n12825 = 2_n11282 | 2_n3517;
assign 2_n6541 = 2_n1018 & 2_n6093;
assign 2_n12713 = ~(2_n9115 ^ 2_n11924);
assign 2_n1202 = ~(2_n8857 ^ 2_n7842);
assign 2_n7660 = ~(2_n4819 | 2_n10515);
assign 2_n9264 = ~(2_n3198 ^ 2_n7596);
assign 2_n9142 = ~2_n7027;
assign 2_n7859 = 2_n5971 | 2_n8824;
assign 2_n3149 = ~(2_n4535 ^ 2_n501);
assign 2_n1609 = ~(2_n2109 ^ 2_n859);
assign 2_n9327 = ~2_n3990;
assign 2_n3231 = 2_n6130 & 2_n6708;
assign 2_n10429 = 2_n10673 & 2_n8926;
assign 2_n12950 = 2_n12210 & 2_n601;
assign 2_n1874 = 2_n5765 | 2_n4864;
assign 2_n3148 = ~(2_n10798 ^ 2_n10707);
assign 2_n616 = 2_n7284 | 2_n10144;
assign 2_n671 = ~(2_n10853 ^ 2_n11300);
assign 2_n2086 = ~(2_n553 ^ 2_n4133);
assign 2_n5024 = 2_n11026 | 2_n4474;
assign 2_n11107 = ~(2_n202 | 2_n9086);
assign 2_n6869 = 2_n5110 | 2_n2795;
assign 2_n7584 = 2_n9304 | 2_n8148;
assign 2_n315 = 2_n5664 | 2_n2145;
assign 2_n1401 = 2_n2154 | 2_n6459;
assign 2_n9243 = ~2_n11225;
assign 2_n3861 = 2_n1891 | 2_n11920;
assign 2_n1212 = 2_n1960 | 2_n1019;
assign 2_n3297 = 2_n9370 | 2_n6402;
assign 2_n3300 = 2_n8405 | 2_n9188;
assign 2_n12046 = 2_n8870 | 2_n8648;
assign 2_n9496 = 2_n8687 | 2_n4474;
assign 2_n6471 = 2_n11598 | 2_n5096;
assign 2_n9681 = 2_n5348 | 2_n581;
assign 2_n4006 = ~(2_n2937 ^ 2_n1297);
assign 2_n9338 = ~(2_n11968 ^ 2_n6);
assign 2_n5893 = 2_n6221 | 2_n9851;
assign 2_n3578 = ~2_n3003;
assign 2_n12745 = ~2_n9381;
assign 2_n10475 = ~2_n10394;
assign 2_n856 = 2_n6977 | 2_n10919;
assign 2_n12524 = 2_n3617 | 2_n6513;
assign 2_n3777 = 2_n11032 | 2_n12830;
assign 2_n9834 = 2_n1937 | 2_n11820;
assign 2_n6502 = ~(2_n11937 ^ 2_n1547);
assign 2_n6989 = ~(2_n100 ^ 2_n12100);
assign 2_n4632 = 2_n3494 & 2_n2646;
assign 2_n8749 = ~2_n1304;
assign 2_n11275 = 2_n9858 & 2_n10972;
assign 2_n12554 = 2_n5602 | 2_n2463;
assign 2_n4247 = 2_n7449 | 2_n8830;
assign 2_n5965 = ~(2_n1010 ^ 2_n5187);
assign 2_n8509 = ~2_n2533;
assign 2_n10224 = 2_n4535 | 2_n501;
assign 2_n9119 = 2_n12324 | 2_n2736;
assign 2_n8402 = ~(2_n730 ^ 2_n4345);
assign 2_n499 = 2_n9093 & 2_n5682;
assign 2_n7520 = 2_n9886 & 2_n3370;
assign 2_n155 = ~(2_n2826 ^ 2_n758);
assign 2_n7515 = ~(2_n6365 ^ 2_n9702);
assign 2_n9034 = ~(2_n6512 | 2_n12681);
assign 2_n4643 = ~2_n8580;
assign 2_n9096 = ~(2_n946 ^ 2_n3258);
assign 2_n6187 = ~(2_n8339 ^ 2_n9540);
assign 2_n225 = ~(2_n8448 ^ 2_n10161);
assign 2_n1700 = ~2_n3531;
assign 2_n2099 = ~2_n5331;
assign 2_n4100 = ~2_n12582;
assign 2_n4853 = ~2_n8324;
assign 2_n4009 = ~(2_n6813 ^ 2_n4156);
assign 2_n10504 = 2_n5575 | 2_n7395;
assign 2_n2525 = 2_n12361 | 2_n12816;
assign 2_n9048 = 2_n7116 | 2_n7952;
assign 2_n9907 = 2_n8750 & 2_n10537;
assign 2_n3115 = ~2_n1017;
assign 2_n5151 = 2_n10118 | 2_n5887;
assign 2_n7448 = ~(2_n8044 | 2_n8319);
assign 2_n6453 = ~(2_n10008 ^ 2_n8494);
assign 2_n3989 = ~2_n11563;
assign 2_n7642 = 2_n2407 | 2_n12137;
assign 2_n5270 = ~(2_n7953 ^ 2_n12148);
assign 2_n5078 = ~(2_n7531 ^ 2_n9259);
assign 2_n7414 = 2_n10677 | 2_n5079;
assign 2_n12390 = 2_n1169 | 2_n4891;
assign 2_n6062 = 2_n7984 | 2_n1541;
assign 2_n1414 = ~(2_n5260 ^ 2_n1108);
assign 2_n2996 = ~(2_n2120 ^ 2_n12885);
assign 2_n5538 = ~2_n4141;
assign 2_n11698 = ~2_n4903;
assign 2_n6460 = 2_n1534 & 2_n8112;
assign 2_n8951 = ~2_n1646;
assign 2_n4434 = ~2_n12723;
assign 2_n4728 = 2_n5575 | 2_n7558;
assign 2_n5354 = 2_n4568 | 2_n12558;
assign 2_n11527 = ~(2_n1456 ^ 2_n8842);
assign 2_n3938 = 2_n12633 | 2_n6508;
assign 2_n326 = 2_n5989 | 2_n6704;
assign 2_n6828 = ~(2_n12430 | 2_n6281);
assign 2_n8698 = 2_n4422 | 2_n12809;
assign 2_n11688 = 2_n5619 & 2_n7308;
assign 2_n7048 = ~(2_n7474 ^ 2_n7654);
assign 2_n12364 = ~(2_n2536 ^ 2_n2670);
assign 2_n2420 = 2_n2011 & 2_n4899;
assign 2_n11659 = 2_n8304 & 2_n10469;
assign 2_n6239 = 2_n11958 | 2_n6455;
assign 2_n6399 = ~(2_n8781 | 2_n4330);
assign 2_n3254 = 2_n2506 & 2_n11807;
assign 2_n3583 = 2_n7384 | 2_n2005;
assign 2_n11976 = ~2_n6303;
assign 2_n105 = 2_n11037 & 2_n10573;
assign 2_n7795 = 2_n8510 & 2_n8274;
assign 2_n11420 = 2_n10202 & 2_n9729;
assign 2_n3834 = 2_n5419 & 2_n11619;
assign 2_n11656 = 2_n3176 & 2_n8167;
assign 2_n6357 = ~(2_n9414 ^ 2_n2038);
assign 2_n7319 = 2_n9081 | 2_n6258;
assign 2_n12450 = ~(2_n8304 ^ 2_n190);
assign 2_n7780 = 2_n10761 | 2_n3234;
assign 2_n4585 = 2_n4725 | 2_n12396;
assign 2_n6924 = 2_n10750 | 2_n7382;
assign 2_n1344 = ~2_n165;
assign 2_n10221 = ~(2_n8436 ^ 2_n86);
assign 2_n4150 = 2_n11694 | 2_n4377;
assign 2_n12927 = ~(2_n6566 | 2_n4542);
assign 2_n483 = 2_n9621 | 2_n1490;
assign 2_n652 = ~(2_n4962 ^ 2_n10016);
assign 2_n642 = ~(2_n296 ^ 2_n6837);
assign 2_n952 = ~(2_n9134 ^ 2_n5775);
assign 2_n7066 = ~(2_n6659 ^ 2_n7524);
assign 2_n10687 = ~(2_n9445 ^ 2_n4567);
assign 2_n6400 = ~(2_n474 ^ 2_n1556);
assign 2_n3230 = ~(2_n12359 ^ 2_n94);
assign 2_n2231 = 2_n8730 & 2_n5588;
assign 2_n7988 = ~(2_n5881 ^ 2_n9979);
assign 2_n4169 = ~2_n11628;
assign 2_n6295 = 2_n8838 | 2_n8029;
assign 2_n7770 = 2_n5600 | 2_n2793;
assign 2_n984 = ~(2_n6076 | 2_n5169);
assign 2_n3712 = ~2_n5495;
assign 2_n4571 = 2_n955 | 2_n5442;
assign 2_n1828 = 2_n4956 & 2_n5000;
assign 2_n6352 = 2_n6290 | 2_n11439;
assign 2_n3454 = ~(2_n12422 | 2_n8568);
assign 2_n9128 = ~(2_n2532 | 2_n4802);
assign 2_n10895 = 2_n3065 & 2_n577;
assign 2_n2137 = 2_n11417 | 2_n1314;
assign 2_n11597 = 2_n10101 | 2_n2218;
assign 2_n1858 = ~(2_n9969 ^ 2_n7604);
assign 2_n2815 = ~2_n7946;
assign 2_n5332 = ~(2_n3608 ^ 2_n11467);
assign 2_n10626 = 2_n11037 | 2_n10573;
assign 2_n4548 = 2_n10564 | 2_n9733;
assign 2_n4560 = 2_n11390 | 2_n3431;
assign 2_n9409 = ~(2_n4536 ^ 2_n4220);
assign 2_n7329 = 2_n7404 & 2_n11438;
assign 2_n3841 = 2_n5913 | 2_n2751;
assign 2_n11393 = ~(2_n9942 ^ 2_n2477);
assign 2_n3788 = ~(2_n8557 | 2_n7653);
assign 2_n5763 = ~2_n12115;
assign 2_n1122 = ~2_n2413;
assign 2_n1862 = 2_n1699 | 2_n8740;
assign 2_n2768 = 2_n11621 & 2_n11956;
assign 2_n1739 = ~2_n6431;
assign 2_n4996 = ~(2_n1960 ^ 2_n1019);
assign 2_n3355 = ~(2_n11992 | 2_n1293);
assign 2_n2410 = ~(2_n195 ^ 2_n12049);
assign 2_n12878 = ~2_n2038;
assign 2_n131 = 2_n11601 | 2_n10724;
assign 2_n4482 = 2_n7474 & 2_n1681;
assign 2_n4398 = 2_n3549 & 2_n98;
assign 2_n6733 = ~(2_n1804 ^ 2_n1105);
assign 2_n8381 = ~(2_n5202 ^ 2_n12240);
assign 2_n4423 = ~2_n302;
assign 2_n3714 = ~2_n1716;
assign 2_n4126 = 2_n11958 | 2_n10919;
assign 2_n5410 = ~2_n8940;
assign 2_n12702 = ~(2_n8864 ^ 2_n8788);
assign 2_n3908 = 2_n3891 | 2_n8409;
assign 2_n11517 = 2_n11958 | 2_n12357;
assign 2_n2762 = ~2_n11553;
assign 2_n10149 = ~(2_n7248 | 2_n12159);
assign 2_n77 = 2_n8227 | 2_n10209;
assign 2_n4282 = 2_n12195 & 2_n4622;
assign 2_n1430 = ~(2_n4910 ^ 2_n4361);
assign 2_n2182 = 2_n994 | 2_n2076;
assign 2_n12015 = 2_n686 | 2_n5012;
assign 2_n4532 = 2_n2078 | 2_n10596;
assign 2_n7843 = 2_n12632 | 2_n10244;
assign 2_n7202 = 2_n2626 | 2_n4041;
assign 2_n6034 = 2_n2288 & 2_n1145;
assign 2_n10859 = ~(2_n9744 ^ 2_n3963);
assign 2_n8203 = 2_n9748 & 2_n10395;
assign 2_n4563 = ~(2_n3463 | 2_n8178);
assign 2_n7756 = 2_n4498 | 2_n1851;
assign 2_n10277 = ~(2_n8277 | 2_n12370);
assign 2_n7168 = 2_n6595 | 2_n6639;
assign 2_n364 = ~(2_n3551 ^ 2_n12205);
assign 2_n4227 = ~(2_n3210 ^ 2_n11192);
assign 2_n5123 = ~(2_n2155 ^ 2_n5786);
assign 2_n8311 = 2_n4768 | 2_n9619;
assign 2_n2206 = ~(2_n5618 ^ 2_n1430);
assign 2_n5762 = ~(2_n12913 ^ 2_n12239);
assign 2_n11817 = ~(2_n3106 | 2_n11945);
assign 2_n8807 = ~2_n3465;
assign 2_n5023 = 2_n674 & 2_n10606;
assign 2_n401 = 2_n10852 | 2_n12019;
assign 2_n10162 = 2_n2756 | 2_n327;
assign 2_n11990 = 2_n8984 & 2_n12268;
assign 2_n4216 = ~2_n4275;
assign 2_n2041 = 2_n12157 | 2_n11197;
assign 2_n10514 = ~2_n10711;
assign 2_n7764 = 2_n12503 | 2_n4654;
assign 2_n7305 = 2_n6242 & 2_n8791;
assign 2_n8679 = 2_n2526 | 2_n8491;
assign 2_n10193 = 2_n705 & 2_n1310;
assign 2_n10558 = ~(2_n12880 ^ 2_n2690);
assign 2_n7848 = ~(2_n8713 | 2_n6850);
assign 2_n5792 = 2_n4932 & 2_n12548;
assign 2_n2567 = ~(2_n2686 ^ 2_n10618);
assign 2_n8252 = ~(2_n8011 ^ 2_n10518);
assign 2_n1488 = ~2_n11227;
assign 2_n8435 = 2_n4637 & 2_n11288;
assign 2_n2748 = ~2_n5916;
assign 2_n6449 = ~(2_n5177 | 2_n10438);
assign 2_n10775 = 2_n677 & 2_n7811;
assign 2_n8491 = ~(2_n6258 ^ 2_n12412);
assign 2_n9787 = 2_n11026 | 2_n2020;
assign 2_n2235 = ~(2_n9109 ^ 2_n6207);
assign 2_n9084 = ~(2_n1961 ^ 2_n6791);
assign 2_n8796 = ~2_n3179;
assign 2_n1920 = 2_n1266 | 2_n2090;
assign 2_n8261 = 2_n3126 & 2_n188;
assign 2_n12905 = 2_n7998 & 2_n4153;
assign 2_n8722 = ~2_n9541;
assign 2_n8593 = ~(2_n5024 ^ 2_n5255);
assign 2_n1489 = 2_n3050 & 2_n11524;
assign 2_n11566 = ~(2_n7572 ^ 2_n7394);
assign 2_n5954 = ~2_n5967;
assign 2_n11030 = ~(2_n7761 ^ 2_n3259);
assign 2_n2011 = 2_n4628 | 2_n12754;
assign 2_n5685 = 2_n3743 | 2_n9144;
assign 2_n8083 = 2_n1471 & 2_n8433;
assign 2_n638 = 2_n12119 | 2_n530;
assign 2_n991 = 2_n5530 | 2_n7382;
assign 2_n4829 = ~(2_n7148 ^ 2_n8106);
assign 2_n12781 = 2_n5575 | 2_n12274;
assign 2_n4380 = 2_n10142 | 2_n7703;
assign 2_n913 = 2_n6977 | 2_n11122;
assign 2_n9121 = ~(2_n597 ^ 2_n1289);
assign 2_n12879 = 2_n1051 | 2_n11820;
assign 2_n4064 = 2_n6534 & 2_n10826;
assign 2_n11024 = 2_n8127 | 2_n4400;
assign 2_n12561 = 2_n12669 | 2_n6360;
assign 2_n12946 = ~2_n8353;
assign 2_n12712 = 2_n996 & 2_n11791;
assign 2_n10033 = 2_n1727 & 2_n12514;
assign 2_n796 = 2_n5341 & 2_n11947;
assign 2_n3550 = 2_n1153 | 2_n55;
assign 2_n869 = ~(2_n3440 | 2_n5755);
assign 2_n2998 = ~(2_n436 | 2_n3299);
assign 2_n6342 = ~(2_n6293 ^ 2_n9157);
assign 2_n1655 = 2_n12110 & 2_n1133;
assign 2_n2497 = 2_n7864 & 2_n8099;
assign 2_n5487 = ~(2_n8299 ^ 2_n10860);
assign 2_n5028 = ~(2_n9719 ^ 2_n11529);
assign 2_n1382 = 2_n12622 | 2_n3919;
assign 2_n11584 = ~(2_n6813 | 2_n10871);
assign 2_n2309 = 2_n12200 & 2_n6975;
assign 2_n10029 = ~(2_n12765 ^ 2_n8664);
assign 2_n12674 = ~(2_n205 ^ 2_n11965);
assign 2_n10869 = 2_n6373 | 2_n28;
assign 2_n8536 = 2_n191 | 2_n8970;
assign 2_n8136 = 2_n8423 & 2_n7315;
assign 2_n5890 = 2_n9222 | 2_n342;
assign 2_n5009 = ~(2_n9480 ^ 2_n6956);
assign 2_n4650 = 2_n11887 | 2_n3224;
assign 2_n7491 = 2_n12119 | 2_n7136;
assign 2_n12636 = 2_n4266 & 2_n3626;
assign 2_n3462 = 2_n7495 | 2_n1162;
assign 2_n9426 = 2_n1808 & 2_n2210;
assign 2_n7404 = 2_n8348 | 2_n12282;
assign 2_n543 = ~2_n7530;
assign 2_n3620 = 2_n4059 | 2_n1079;
assign 2_n11869 = 2_n383 | 2_n10621;
assign 2_n3671 = 2_n10339 | 2_n10854;
assign 2_n10915 = 2_n6461 | 2_n3148;
assign 2_n6221 = ~2_n4868;
assign 2_n5223 = ~2_n2629;
assign 2_n10058 = ~(2_n1061 | 2_n12022);
assign 2_n1296 = ~(2_n4986 ^ 2_n4810);
assign 2_n12138 = ~2_n6816;
assign 2_n6716 = ~(2_n6894 ^ 2_n1616);
assign 2_n11859 = ~(2_n4389 | 2_n6680);
assign 2_n7521 = ~(2_n5644 | 2_n7220);
assign 2_n1782 = ~2_n12764;
assign 2_n1405 = 2_n3285 | 2_n2738;
assign 2_n9298 = ~(2_n3374 ^ 2_n11789);
assign 2_n8247 = 2_n4953 & 2_n8301;
assign 2_n2925 = 2_n11689 | 2_n11058;
assign 2_n12747 = 2_n3743 | 2_n4654;
assign 2_n2475 = 2_n7504 & 2_n224;
assign 2_n5822 = ~(2_n10402 ^ 2_n3249);
assign 2_n12616 = 2_n11556 & 2_n6173;
assign 2_n963 = ~(2_n2893 ^ 2_n1014);
assign 2_n8619 = 2_n3804 | 2_n1700;
assign 2_n10886 = 2_n5945 | 2_n3903;
assign 2_n4017 = ~(2_n10839 ^ 2_n600);
assign 2_n10893 = 2_n6717 | 2_n5867;
assign 2_n8059 = ~2_n4700;
assign 2_n3188 = ~(2_n12734 ^ 2_n1283);
assign 2_n8489 = 2_n9570 | 2_n12050;
assign 2_n2148 = ~(2_n688 | 2_n7853);
assign 2_n11557 = 2_n5355 | 2_n1455;
assign 2_n6198 = ~(2_n5234 | 2_n9597);
assign 2_n2380 = ~2_n3083;
assign 2_n6612 = ~(2_n7312 ^ 2_n8718);
assign 2_n1606 = 2_n636 | 2_n8259;
assign 2_n3728 = 2_n1511 | 2_n7602;
assign 2_n6980 = ~(2_n3005 ^ 2_n9251);
assign 2_n2114 = ~(2_n3201 | 2_n10782);
assign 2_n8246 = ~2_n9454;
assign 2_n12433 = 2_n12503 | 2_n12771;
assign 2_n4570 = ~(2_n10481 ^ 2_n6480);
assign 2_n11006 = ~(2_n5064 ^ 2_n8974);
assign 2_n3482 = ~2_n2871;
assign 2_n3076 = 2_n12361 | 2_n7876;
assign 2_n4757 = ~(2_n8573 ^ 2_n9691);
assign 2_n10076 = ~(2_n5364 | 2_n9781);
assign 2_n12586 = 2_n2597 & 2_n934;
assign 2_n11270 = ~(2_n6242 ^ 2_n2469);
assign 2_n149 = ~2_n2913;
assign 2_n160 = 2_n5710 & 2_n12926;
assign 2_n576 = ~2_n7726;
assign 2_n9706 = ~(2_n4427 ^ 2_n1110);
assign 2_n7932 = 2_n8545 | 2_n12783;
assign 2_n9585 = 2_n7662 & 2_n1800;
assign 2_n330 = 2_n7919 & 2_n5872;
assign 2_n9976 = 2_n12237 | 2_n6513;
assign 2_n2714 = 2_n6977 | 2_n11896;
assign 2_n4618 = 2_n8348 & 2_n12282;
assign 2_n11782 = 2_n7449 | 2_n5258;
assign 2_n4518 = ~2_n11623;
assign 2_n7754 = 2_n3746 | 2_n6114;
assign 2_n12410 = ~(2_n10401 | 2_n8771);
assign 2_n90 = ~(2_n5995 | 2_n769);
assign 2_n4872 = 2_n2089 | 2_n7962;
assign 2_n3264 = 2_n12025 & 2_n9956;
assign 2_n4345 = ~(2_n5503 ^ 2_n12844);
assign 2_n5596 = 2_n4958 & 2_n5514;
assign 2_n7112 = 2_n4498 | 2_n3911;
assign 2_n1803 = 2_n10142 | 2_n11430;
assign 2_n2250 = ~(2_n6702 ^ 2_n9901);
assign 2_n3203 = ~(2_n6582 ^ 2_n10121);
assign 2_n9288 = 2_n11294 & 2_n7507;
assign 2_n8125 = 2_n5377 & 2_n6701;
assign 2_n1431 = ~(2_n6994 ^ 2_n1538);
assign 2_n7742 = ~2_n2094;
assign 2_n11261 = ~(2_n9165 | 2_n2729);
assign 2_n11581 = 2_n11433 | 2_n3903;
assign 2_n11738 = ~(2_n9699 ^ 2_n2084);
assign 2_n9679 = ~(2_n6137 ^ 2_n3901);
assign 2_n11000 = ~(2_n1177 | 2_n5354);
assign 2_n2752 = ~(2_n10480 ^ 2_n1173);
assign 2_n12198 = 2_n7685 & 2_n3179;
assign 2_n7007 = ~2_n4241;
assign 2_n3221 = 2_n5355 | 2_n8859;
assign 2_n3234 = 2_n348 & 2_n5667;
assign 2_n4925 = ~2_n9390;
assign 2_n3330 = 2_n9070 & 2_n9786;
assign 2_n4488 = 2_n8291 & 2_n3104;
assign 2_n453 = 2_n8674 | 2_n5642;
assign 2_n769 = 2_n6718 | 2_n1476;
assign 2_n8876 = ~(2_n10443 ^ 2_n5544);
assign 2_n4905 = ~(2_n10568 ^ 2_n133);
assign 2_n10736 = ~2_n3294;
assign 2_n6135 = ~(2_n12428 ^ 2_n7210);
assign 2_n11558 = ~(2_n3684 ^ 2_n12333);
assign 2_n8109 = ~2_n7159;
assign 2_n6179 = ~(2_n4468 ^ 2_n3034);
assign 2_n6378 = ~2_n4953;
assign 2_n6256 = 2_n4628 | 2_n1163;
assign 2_n6773 = ~(2_n6688 ^ 2_n6255);
assign 2_n3693 = 2_n8692 & 2_n2421;
assign 2_n2210 = 2_n2786 & 2_n9009;
assign 2_n9140 = 2_n2584 & 2_n9258;
assign 2_n6262 = ~(2_n5018 ^ 2_n12593);
assign 2_n11649 = 2_n9825 & 2_n8469;
assign 2_n10766 = 2_n5209 ^ 2_n7241;
assign 2_n1167 = ~(2_n11864 ^ 2_n11458);
assign 2_n9615 = 2_n857 & 2_n6691;
assign 2_n11176 = 2_n4059 | 2_n7246;
assign 2_n2469 = 2_n1397 & 2_n8359;
assign 2_n11483 = ~2_n9351;
assign 2_n6801 = 2_n11958 | 2_n9971;
assign 2_n5086 = ~2_n12511;
assign 2_n9292 = 2_n3567 | 2_n11440;
assign 2_n4954 = ~(2_n7906 ^ 2_n4338);
assign 2_n4183 = 2_n3746 | 2_n5540;
assign 2_n5466 = 2_n2099 | 2_n4818;
assign 2_n7573 = ~2_n9838;
assign 2_n9361 = ~(2_n24 ^ 2_n7334);
assign 2_n2864 = 2_n5743 | 2_n7840;
assign 2_n6837 = 2_n7709 | 2_n28;
assign 2_n2683 = ~2_n544;
assign 2_n3826 = 2_n2137 & 2_n4335;
assign 2_n3475 = ~(2_n0 ^ 2_n2127);
assign 2_n12050 = 2_n1212 & 2_n3039;
assign 2_n10782 = 2_n5899 & 2_n2928;
assign 2_n10116 = ~(2_n6935 ^ 2_n12438);
assign 2_n5062 = ~(2_n11642 ^ 2_n8562);
assign 2_n289 = ~(2_n2714 ^ 2_n7125);
assign 2_n8818 = 2_n7084 | 2_n9091;
assign 2_n2673 = ~(2_n6301 ^ 2_n2823);
assign 2_n539 = 2_n4769 & 2_n8956;
assign 2_n2058 = 2_n3014 & 2_n9939;
assign 2_n5975 = 2_n9036 & 2_n8225;
assign 2_n5728 = ~(2_n496 ^ 2_n2939);
assign 2_n56 = ~(2_n8342 ^ 2_n5900);
assign 2_n11183 = 2_n1054 | 2_n12657;
assign 2_n324 = 2_n5378 & 2_n8697;
assign 2_n10323 = 2_n8959 | 2_n1413;
assign 2_n2912 = ~(2_n12478 ^ 2_n7759);
assign 2_n5250 = 2_n8847 | 2_n9356;
assign 2_n5931 = 2_n5291 & 2_n11040;
assign 2_n12306 = 2_n1051 | 2_n5540;
assign 2_n9761 = ~2_n2742;
assign 2_n6666 = 2_n5456 | 2_n87;
assign 2_n12597 = 2_n12361 | 2_n8768;
assign 2_n8574 = 2_n969 | 2_n5046;
assign 2_n251 = ~(2_n11285 ^ 2_n33);
assign 2_n1620 = 2_n686 | 2_n9741;
assign 2_n11691 = 2_n9082 | 2_n10865;
assign 2_n6496 = ~(2_n12318 | 2_n6900);
assign 2_n11088 = ~2_n4145;
assign 2_n1251 = 2_n10392 & 2_n10911;
assign 2_n9870 = 2_n1642 & 2_n12325;
assign 2_n5828 = 2_n5355 | 2_n1915;
assign 2_n12824 = ~(2_n1418 ^ 2_n8941);
assign 2_n7883 = 2_n9370 | 2_n4400;
assign 2_n11635 = ~(2_n12479 | 2_n8174);
assign 2_n994 = ~2_n1333;
assign 2_n11092 = ~(2_n5368 | 2_n2221);
assign 2_n8943 = 2_n5394 & 2_n5152;
assign 2_n5904 = ~(2_n6149 | 2_n3454);
assign 2_n6419 = ~(2_n3930 ^ 2_n4483);
assign 2_n4116 = 2_n6977 | 2_n3903;
assign 2_n10352 = 2_n8738 | 2_n1509;
assign 2_n3461 = 2_n4628 | 2_n10854;
assign 2_n9628 = ~(2_n4857 ^ 2_n2310);
assign 2_n6820 = 2_n636 | 2_n12754;
assign 2_n5055 = 2_n8187 | 2_n11746;
assign 2_n11986 = ~(2_n1657 ^ 2_n9030);
assign 2_n6598 = ~(2_n2783 | 2_n1531);
assign 2_n7412 = ~(2_n7221 ^ 2_n10500);
assign 2_n5296 = ~2_n6188;
assign 2_n11344 = 2_n10953 | 2_n9999;
assign 2_n9275 = 2_n7431 & 2_n1175;
assign 2_n1063 = ~(2_n9834 ^ 2_n11043);
assign 2_n5188 = 2_n12053 & 2_n4464;
assign 2_n7789 = ~2_n9311;
assign 2_n3644 = ~2_n11908;
assign 2_n8030 = ~(2_n5805 ^ 2_n11447);
assign 2_n1814 = ~(2_n8084 ^ 2_n11976);
assign 2_n924 = ~(2_n4272 ^ 2_n11833);
assign 2_n8132 = 2_n2472 | 2_n11952;
assign 2_n3956 = 2_n504 & 2_n3873;
assign 2_n6270 = ~2_n12537;
assign 2_n10871 = ~2_n1385;
assign 2_n562 = 2_n5982 | 2_n9166;
assign 2_n6206 = ~2_n6748;
assign 2_n10680 = ~(2_n9134 | 2_n10397);
assign 2_n10912 = 2_n2217 | 2_n10916;
assign 2_n4091 = 2_n3552 & 2_n7061;
assign 2_n8474 = 2_n1699 | 2_n8648;
assign 2_n5043 = ~(2_n8917 ^ 2_n5487);
assign 2_n12082 = ~(2_n10432 | 2_n154);
assign 2_n10052 = 2_n7050 & 2_n2106;
assign 2_n3677 = ~(2_n4720 ^ 2_n11918);
assign 2_n7712 = 2_n8308 & 2_n6581;
assign 2_n2944 = ~(2_n384 | 2_n5972);
assign 2_n9802 = 2_n7493 & 2_n8551;
assign 2_n5768 = ~(2_n5972 ^ 2_n384);
assign 2_n4753 = ~2_n4960;
assign 2_n4979 = ~(2_n6951 | 2_n12081);
assign 2_n7857 = ~(2_n10104 ^ 2_n4835);
assign 2_n12113 = ~(2_n12456 ^ 2_n12743);
assign 2_n11039 = ~(2_n11351 ^ 2_n6023);
assign 2_n1225 = 2_n7551 | 2_n10825;
assign 2_n640 = 2_n12177 & 2_n12386;
assign 2_n9727 = 2_n4628 | 2_n9188;
assign 2_n9122 = 2_n12119 | 2_n8655;
assign 2_n4755 = 2_n5530 | 2_n10311;
assign 2_n5530 = ~2_n12069;
assign 2_n497 = 2_n7266 | 2_n4385;
assign 2_n12282 = ~(2_n3967 ^ 2_n5927);
assign 2_n2717 = 2_n3096 | 2_n5012;
assign 2_n7361 = ~(2_n107 ^ 2_n11005);
assign 2_n7368 = ~(2_n9274 ^ 2_n12513);
assign 2_n5546 = 2_n3642 | 2_n10963;
assign 2_n12813 = ~2_n3258;
assign 2_n3629 = 2_n276 | 2_n3507;
assign 2_n6746 = 2_n7191 | 2_n942;
assign 2_n3613 = ~(2_n3747 ^ 2_n1561);
assign 2_n8190 = ~(2_n5202 | 2_n9513);
assign 2_n6972 = ~(2_n6788 | 2_n1214);
assign 2_n1398 = 2_n8738 | 2_n4875;
assign 2_n12487 = 2_n507 & 2_n2797;
assign 2_n3707 = 2_n8390 & 2_n2744;
assign 2_n6547 = ~2_n10531;
assign 2_n12945 = 2_n10750 | 2_n12124;
assign 2_n7389 = ~2_n9583;
assign 2_n7140 = 2_n9268 | 2_n11706;
assign 2_n4336 = 2_n686 | 2_n11820;
assign 2_n5627 = 2_n4529 & 2_n8749;
assign 2_n3392 = 2_n9170 | 2_n1546;
assign 2_n11855 = 2_n11390 & 2_n3431;
assign 2_n1999 = ~(2_n9931 ^ 2_n7926);
assign 2_n1937 = ~2_n11311;
assign 2_n5678 = ~(2_n6208 | 2_n5878);
assign 2_n8494 = ~(2_n2056 ^ 2_n2595);
assign 2_n8235 = ~(2_n10421 ^ 2_n11367);
assign 2_n5008 = ~2_n555;
assign 2_n700 = ~(2_n1202 ^ 2_n10115);
assign 2_n1006 = ~(2_n6442 | 2_n10619);
assign 2_n2088 = ~(2_n3810 ^ 2_n3181);
assign 2_n11449 = 2_n4304 | 2_n1117;
assign 2_n5640 = ~(2_n8296 ^ 2_n1427);
assign 2_n7928 = ~2_n6016;
assign 2_n8504 = 2_n2530 & 2_n7610;
assign 2_n4309 = ~(2_n11039 ^ 2_n6641);
assign 2_n8000 = 2_n1699 | 2_n2964;
assign 2_n6977 = ~2_n6986;
assign 2_n6535 = 2_n393 & 2_n7260;
assign 2_n10388 = ~(2_n7890 | 2_n9162);
assign 2_n12864 = 2_n5016 & 2_n12202;
assign 2_n8040 = ~2_n308;
assign 2_n6960 = 2_n5505 & 2_n5009;
assign 2_n10655 = ~2_n8538;
assign 2_n5681 = 2_n5809 | 2_n8655;
assign 2_n1919 = 2_n6373 | 2_n9078;
assign 2_n2609 = ~(2_n4415 ^ 2_n8175);
assign 2_n2488 = 2_n7283 | 2_n10419;
assign 2_n2474 = 2_n10827 & 2_n10944;
assign 2_n6550 = 2_n453 & 2_n9013;
assign 2_n5549 = 2_n4911 | 2_n7703;
assign 2_n12049 = ~2_n12256;
assign 2_n1716 = 2_n6354 & 2_n10952;
assign 2_n12575 = ~(2_n7850 ^ 2_n3394);
assign 2_n9033 = ~2_n12001;
assign 2_n7518 = ~(2_n2003 ^ 2_n12762);
assign 2_n10586 = ~(2_n10701 | 2_n7148);
assign 2_n10897 = ~2_n4657;
assign 2_n2658 = ~2_n5274;
assign 2_n2016 = ~2_n3064;
assign 2_n10394 = 2_n3992 & 2_n7270;
assign 2_n726 = 2_n8452 | 2_n8978;
assign 2_n2833 = 2_n2050 | 2_n4736;
assign 2_n1734 = 2_n9370 | 2_n6389;
assign 2_n2423 = ~(2_n10290 | 2_n12640);
assign 2_n4318 = ~(2_n432 ^ 2_n10882);
assign 2_n4322 = 2_n10142 | 2_n1738;
assign 2_n12133 = 2_n12391 & 2_n4970;
assign 2_n12124 = ~2_n2347;
assign 2_n4099 = 2_n3912 & 2_n10030;
assign 2_n11142 = 2_n7449 | 2_n4642;
assign 2_n2331 = ~(2_n10272 ^ 2_n3390);
assign 2_n660 = ~2_n6624;
assign 2_n6574 = 2_n12596 | 2_n3288;
assign 2_n182 = 2_n5809 | 2_n826;
assign 2_n1979 = 2_n10298 | 2_n9596;
assign 2_n12658 = ~(2_n6465 ^ 2_n8843);
assign 2_n10534 = ~2_n6007;
assign 2_n6608 = 2_n12454 | 2_n1029;
assign 2_n9547 = 2_n4498 | 2_n6389;
assign 2_n7502 = 2_n12853 | 2_n9586;
assign 2_n12444 = ~(2_n6913 ^ 2_n11383);
assign 2_n622 = ~(2_n5366 ^ 2_n6476);
assign 2_n2161 = 2_n7319 & 2_n2521;
assign 2_n8889 = ~2_n8373;
assign 2_n529 = 2_n2887 & 2_n6963;
assign 2_n10588 = 2_n7407 & 2_n10662;
assign 2_n5690 = 2_n11923 | 2_n9144;
assign 2_n5602 = 2_n8135 & 2_n2229;
assign 2_n8184 = ~(2_n7072 ^ 2_n12449);
assign 2_n4656 = ~(2_n6814 ^ 2_n2929);
assign 2_n2594 = 2_n9082 & 2_n10865;
assign 2_n10180 = 2_n191 | 2_n7881;
assign 2_n1410 = ~(2_n8804 ^ 2_n8391);
assign 2_n12373 = ~(2_n12713 | 2_n10027);
assign 2_n2985 = ~(2_n2550 | 2_n2422);
assign 2_n11223 = ~(2_n3226 ^ 2_n5066);
assign 2_n2440 = ~(2_n2569 ^ 2_n9855);
assign 2_n10010 = 2_n12262 & 2_n8253;
assign 2_n9387 = ~(2_n739 ^ 2_n1318);
assign 2_n6585 = ~(2_n4075 ^ 2_n3385);
assign 2_n2415 = 2_n2363 & 2_n229;
assign 2_n5007 = 2_n10351 & 2_n3629;
assign 2_n8994 = ~(2_n8550 | 2_n10934);
assign 2_n6953 = 2_n1466 | 2_n7055;
assign 2_n2403 = 2_n9190 | 2_n8079;
assign 2_n2513 = ~2_n9124;
assign 2_n6026 = ~(2_n11037 ^ 2_n1883);
assign 2_n10887 = 2_n5945 | 2_n1413;
assign 2_n5511 = 2_n9297 | 2_n10020;
assign 2_n1718 = 2_n8428 | 2_n3356;
assign 2_n10399 = ~(2_n2744 ^ 2_n1553);
assign 2_n3339 = ~(2_n2412 ^ 2_n7991);
assign 2_n6576 = ~(2_n1544 ^ 2_n9558);
assign 2_n6402 = ~2_n2585;
assign 2_n4893 = 2_n9389 | 2_n510;
assign 2_n7638 = ~(2_n7882 | 2_n8454);
assign 2_n8267 = 2_n636 | 2_n7382;
assign 2_n5401 = 2_n9732 & 2_n3404;
assign 2_n12096 = 2_n114 | 2_n1413;
assign 2_n398 = 2_n928 | 2_n6381;
assign 2_n3169 = 2_n11041 | 2_n7423;
assign 2_n3713 = ~2_n10497;
assign 2_n6191 = 2_n11415 | 2_n12606;
assign 2_n8582 = 2_n11425 & 2_n6025;
assign 2_n8860 = 2_n8582 | 2_n772;
assign 2_n9571 = ~(2_n767 ^ 2_n9686);
assign 2_n7830 = ~2_n11055;
assign 2_n4846 = 2_n10835 | 2_n7921;
assign 2_n4588 = ~(2_n5681 | 2_n10646);
assign 2_n4525 = ~(2_n546 ^ 2_n7011);
assign 2_n1315 = 2_n5530 | 2_n12686;
assign 2_n3018 = ~(2_n7740 ^ 2_n12724);
assign 2_n7461 = 2_n3131 | 2_n10813;
assign 2_n3421 = ~2_n12145;
assign 2_n3748 = 2_n5438 & 2_n11986;
assign 2_n9828 = 2_n5543 & 2_n3485;
assign 2_n6905 = 2_n7690 & 2_n12925;
assign 2_n8563 = ~(2_n11784 ^ 2_n5536);
assign 2_n12276 = ~(2_n858 ^ 2_n7757);
assign 2_n9926 = ~(2_n5982 ^ 2_n3923);
assign 2_n993 = 2_n11887 | 2_n12535;
assign 2_n12477 = 2_n6407 | 2_n2208;
assign 2_n3227 = ~2_n1091;
assign 2_n5004 = 2_n4647 & 2_n11236;
assign 2_n12027 = 2_n7283 | 2_n11430;
assign 2_n6899 = 2_n5575 | 2_n5540;
assign 2_n10743 = ~(2_n11620 ^ 2_n3100);
assign 2_n2002 = ~2_n11541;
assign 2_n6594 = ~(2_n400 | 2_n4034);
assign 2_n5861 = 2_n4911 | 2_n11827;
assign 2_n8806 = 2_n4617 & 2_n9736;
assign 2_n3838 = ~(2_n4349 | 2_n3580);
assign 2_n4529 = 2_n8247 & 2_n3868;
assign 2_n6879 = 2_n5666 & 2_n8134;
assign 2_n10300 = ~(2_n1990 ^ 2_n8207);
assign 2_n9526 = 2_n10502 & 2_n6189;
assign 2_n6967 = 2_n2633 | 2_n11339;
assign 2_n6615 = ~2_n5282;
assign 2_n4579 = 2_n4561 & 2_n10280;
assign 2_n7892 = 2_n11127 | 2_n9555;
assign 2_n810 = ~2_n8537;
assign 2_n3343 = 2_n5312 | 2_n2886;
assign 2_n3472 = 2_n11478 & 2_n2558;
assign 2_n9125 = ~(2_n34 ^ 2_n11214);
assign 2_n12346 = 2_n2599 | 2_n10681;
assign 2_n9549 = 2_n11923 | 2_n9521;
assign 2_n8650 = 2_n1990 & 2_n7635;
assign 2_n7896 = 2_n4508 & 2_n6184;
assign 2_n11541 = 2_n7449 | 2_n1476;
assign 2_n9612 = ~2_n7081;
assign 2_n12529 = ~(2_n12582 ^ 2_n3893);
assign 2_n7992 = 2_n752 | 2_n7558;
assign 2_n9708 = ~(2_n9293 ^ 2_n4664);
assign 2_n8139 = 2_n8187 | 2_n10419;
assign 2_n10890 = ~(2_n6228 ^ 2_n9525);
assign 2_n1680 = ~(2_n11505 ^ 2_n520);
assign 2_n12464 = ~2_n6709;
assign 2_n5953 = 2_n11719 | 2_n6389;
assign 2_n552 = 2_n5361 & 2_n6282;
assign 2_n2026 = ~2_n3834;
assign 2_n10589 = ~(2_n6997 ^ 2_n5692);
assign 2_n3939 = 2_n2700 | 2_n3268;
assign 2_n4768 = ~(2_n2504 | 2_n3814);
assign 2_n7272 = ~(2_n6914 ^ 2_n4447);
assign 2_n1250 = 2_n2147 | 2_n10329;
assign 2_n2150 = 2_n8505 & 2_n11731;
assign 2_n5586 = ~(2_n11181 ^ 2_n9803);
assign 2_n11110 = 2_n4644 | 2_n11624;
assign 2_n12320 = ~(2_n11851 ^ 2_n9255);
assign 2_n1989 = ~2_n9358;
assign 2_n10267 = ~2_n3953;
assign 2_n11334 = 2_n2197 | 2_n11855;
assign 2_n4907 = 2_n989 | 2_n8859;
assign 2_n9173 = ~(2_n7812 ^ 2_n559);
assign 2_n7137 = 2_n2456 | 2_n8644;
assign 2_n12249 = ~(2_n7753 ^ 2_n11771);
assign 2_n4531 = 2_n5441 | 2_n1862;
assign 2_n7762 = 2_n8462 & 2_n736;
assign 2_n7924 = 2_n1811 & 2_n829;
assign 2_n2184 = 2_n9744 & 2_n3963;
assign 2_n7068 = ~(2_n1310 ^ 2_n7818);
assign 2_n3200 = ~(2_n3056 ^ 2_n3367);
assign 2_n4392 = 2_n11958 | 2_n2589;
assign 2_n973 = ~2_n10228;
assign 2_n1590 = ~(2_n7700 ^ 2_n9132);
assign 2_n10051 = 2_n6687 & 2_n2509;
assign 2_n1271 = 2_n2605 & 2_n11921;
assign 2_n5926 = 2_n807 | 2_n5540;
assign 2_n2391 = ~(2_n387 | 2_n11859);
assign 2_n2175 = 2_n11317 | 2_n1265;
assign 2_n1546 = ~2_n3842;
assign 2_n5719 = ~(2_n10973 ^ 2_n4399);
assign 2_n2399 = ~(2_n11711 | 2_n4833);
assign 2_n5148 = ~(2_n1392 | 2_n2337);
assign 2_n656 = 2_n9246 & 2_n3017;
assign 2_n8493 = ~(2_n7643 ^ 2_n8232);
assign 2_n5875 = ~(2_n12551 | 2_n8647);
assign 2_n252 = 2_n8187 | 2_n1162;
assign 2_n11149 = ~(2_n5075 ^ 2_n9434);
assign 2_n8062 = ~2_n10640;
assign 2_n9332 = 2_n2494 | 2_n10775;
assign 2_n3594 = 2_n11782 | 2_n5114;
assign 2_n5382 = ~(2_n12375 | 2_n7444);
assign 2_n6650 = 2_n7116 | 2_n5540;
assign 2_n7563 = ~(2_n3027 ^ 2_n8459);
assign 2_n12917 = ~(2_n10502 ^ 2_n6189);
assign 2_n10809 = ~(2_n10260 ^ 2_n9975);
assign 2_n2872 = ~2_n10174;
assign 2_n8638 = ~(2_n11744 ^ 2_n499);
assign 2_n10784 = ~(2_n3126 ^ 2_n188);
assign 2_n12553 = ~(2_n3679 ^ 2_n4494);
assign 2_n10274 = 2_n1259 | 2_n3778;
assign 2_n7832 = 2_n41 | 2_n1255;
assign 2_n5288 = 2_n12617 & 2_n1648;
assign 2_n895 = ~2_n4422;
assign 2_n11104 = 2_n688 & 2_n7853;
assign 2_n2340 = 2_n5530 | 2_n8957;
assign 2_n12889 = 2_n2919 | 2_n6319;
assign 2_n1808 = 2_n10750 | 2_n4818;
assign 2_n11719 = ~2_n11257;
assign 2_n4601 = ~(2_n8352 ^ 2_n9879);
assign 2_n9565 = ~(2_n3585 ^ 2_n3554);
assign 2_n1062 = ~(2_n11295 ^ 2_n6155);
assign 2_n3917 = ~2_n6621;
assign 2_n4200 = 2_n164 & 2_n10881;
assign 2_n9304 = 2_n8552 | 2_n6513;
assign 2_n9056 = ~2_n12031;
assign 2_n9981 = ~(2_n2828 ^ 2_n12623);
assign 2_n11507 = 2_n10750 | 2_n8644;
assign 2_n1895 = 2_n1827 & 2_n11479;
assign 2_n9152 = ~(2_n1892 ^ 2_n481);
assign 2_n4302 = 2_n1384 | 2_n9194;
assign 2_n12136 = ~(2_n6322 | 2_n8035);
assign 2_n12915 = 2_n10928 & 2_n6703;
assign 2_n5584 = ~(2_n4767 | 2_n4987);
assign 2_n11661 = ~(2_n8329 | 2_n11063);
assign 2_n10768 = 2_n994 | 2_n7389;
assign 2_n3806 = ~(2_n9163 ^ 2_n402);
assign 2_n7208 = 2_n3561 | 2_n8312;
assign 2_n9439 = ~(2_n12084 ^ 2_n6502);
assign 2_n5925 = 2_n12330 & 2_n3980;
assign 2_n3916 = 2_n4796 | 2_n9493;
assign 2_n565 = ~(2_n10842 ^ 2_n2123);
assign 2_n5036 = 2_n12033 & 2_n6781;
assign 2_n1092 = ~2_n3988;
assign 2_n11535 = 2_n1271 | 2_n12528;
assign 2_n6209 = 2_n4173 & 2_n7858;
assign 2_n7664 = 2_n12512 & 2_n7414;
assign 2_n8792 = 2_n6252 & 2_n7089;
assign 2_n4582 = 2_n8313 | 2_n879;
assign 2_n11277 = ~2_n5526;
assign 2_n7056 = ~(2_n10776 | 2_n5683);
assign 2_n9754 = 2_n4121 & 2_n11975;
assign 2_n11007 = 2_n5783 & 2_n12915;
assign 2_n3398 = ~(2_n11332 ^ 2_n2772);
assign 2_n742 = ~(2_n8927 ^ 2_n9071);
assign 2_n12454 = 2_n4777 & 2_n7475;
assign 2_n1616 = 2_n12503 | 2_n1509;
assign 2_n3964 = 2_n5355 | 2_n7389;
assign 2_n10292 = 2_n12503 | 2_n9144;
assign 2_n6279 = ~(2_n4207 | 2_n3371);
assign 2_n6950 = ~(2_n10379 ^ 2_n964);
assign 2_n1339 = ~(2_n6807 ^ 2_n10465);
assign 2_n6968 = ~2_n6430;
assign 2_n1683 = 2_n5739 & 2_n10241;
assign 2_n4831 = 2_n4510 | 2_n6410;
assign 2_n12036 = ~(2_n7766 | 2_n12898);
assign 2_n1809 = 2_n12237 | 2_n8655;
assign 2_n1702 = 2_n10750 | 2_n6513;
assign 2_n8502 = 2_n7718 | 2_n5884;
assign 2_n8422 = 2_n332 | 2_n3703;
assign 2_n822 = 2_n5362 & 2_n7725;
assign 2_n9091 = 2_n11602 & 2_n7707;
assign 2_n3191 = ~(2_n1755 | 2_n6913);
assign 2_n4720 = ~2_n9332;
assign 2_n5101 = 2_n10797 & 2_n7954;
assign 2_n8516 = 2_n1141 | 2_n1192;
assign 2_n9495 = ~(2_n7317 | 2_n11492);
assign 2_n2303 = ~(2_n11885 ^ 2_n9804);
assign 2_n8389 = 2_n11150 & 2_n6726;
assign 2_n2356 = ~2_n6786;
assign 2_n5392 = 2_n8882 | 2_n12435;
assign 2_n280 = ~(2_n1335 ^ 2_n10027);
assign 2_n2392 = 2_n149 & 2_n368;
assign 2_n6309 = ~2_n7458;
assign 2_n3817 = ~(2_n3247 ^ 2_n5028);
assign 2_n2091 = ~(2_n5904 ^ 2_n1379);
assign 2_n2964 = ~2_n5798;
assign 2_n12714 = ~(2_n2312 ^ 2_n3899);
assign 2_n10672 = 2_n3638 | 2_n7528;
assign 2_n2534 = ~(2_n11468 ^ 2_n7789);
assign 2_n4364 = ~2_n8544;
assign 2_n8147 = ~(2_n12277 ^ 2_n1769);
assign 2_n5610 = ~(2_n7405 ^ 2_n11066);
assign 2_n6249 = 2_n6881 & 2_n6489;
assign 2_n9051 = 2_n12561 & 2_n1586;
assign 2_n9728 = 2_n1471 & 2_n9763;
assign 2_n4522 = 2_n3734 | 2_n12508;
assign 2_n12890 = ~(2_n4292 | 2_n3690);
assign 2_n763 = ~2_n5128;
assign 2_n194 = ~(2_n5281 ^ 2_n8777);
assign 2_n4780 = 2_n1937 | 2_n2232;
assign 2_n6637 = ~(2_n8719 | 2_n2637);
assign 2_n3352 = ~2_n9341;
assign 2_n9252 = 2_n708 & 2_n2032;
assign 2_n4241 = ~(2_n11561 ^ 2_n4067);
assign 2_n595 = 2_n9248 & 2_n6592;
assign 2_n10018 = 2_n2456 | 2_n12686;
assign 2_n7317 = 2_n8026 | 2_n7395;
assign 2_n10951 = 2_n5554 & 2_n11625;
assign 2_n3259 = ~(2_n5828 ^ 2_n5186);
assign 2_n11502 = 2_n9943 & 2_n9035;
assign 2_n6282 = ~(2_n10604 ^ 2_n7356);
assign 2_n3831 = 2_n8276 & 2_n11728;
assign 2_n9930 = ~(2_n1392 ^ 2_n1992);
assign 2_n2193 = ~(2_n5345 ^ 2_n2614);
assign 2_n6264 = ~(2_n5922 ^ 2_n9614);
assign 2_n7343 = ~2_n11155;
assign 2_n2335 = 2_n9370 | 2_n4775;
assign 2_n8458 = 2_n9370 | 2_n7341;
assign 2_n6825 = ~(2_n9861 | 2_n6047);
assign 2_n2968 = 2_n1963 & 2_n11769;
assign 2_n8041 = 2_n1003 & 2_n6517;
assign 2_n5529 = 2_n4302 & 2_n4927;
assign 2_n1133 = ~2_n9197;
assign 2_n5396 = ~2_n3208;
assign 2_n2001 = 2_n1170 | 2_n6748;
assign 2_n1870 = ~2_n6745;
assign 2_n8745 = ~2_n10022;
assign 2_n741 = ~(2_n9190 ^ 2_n7901);
assign 2_n4752 = ~(2_n7350 ^ 2_n454);
assign 2_n4328 = 2_n8405 | 2_n12535;
assign 2_n8263 = ~(2_n9676 | 2_n1451);
assign 2_n4685 = 2_n7641 & 2_n9910;
assign 2_n10865 = ~(2_n9651 ^ 2_n12543);
assign 2_n8508 = 2_n5486 | 2_n3557;
assign 2_n6328 = 2_n962 | 2_n2020;
assign 2_n8461 = 2_n12284 & 2_n663;
assign 2_n6020 = 2_n3211 | 2_n8653;
assign 2_n4290 = 2_n1051 | 2_n6455;
assign 2_n12847 = 2_n4363 | 2_n6321;
assign 2_n10080 = 2_n6977 | 2_n7558;
assign 2_n10250 = 2_n1123 & 2_n396;
assign 2_n7085 = ~(2_n11905 ^ 2_n6715);
assign 2_n7759 = ~2_n9102;
assign 2_n3922 = ~2_n4462;
assign 2_n9718 = ~(2_n11306 ^ 2_n5381);
assign 2_n6467 = ~(2_n8350 ^ 2_n4455);
assign 2_n8032 = ~(2_n6754 ^ 2_n6573);
assign 2_n10281 = 2_n10912 | 2_n6143;
assign 2_n11914 = ~2_n11679;
assign 2_n226 = ~(2_n5350 ^ 2_n5175);
assign 2_n5119 = 2_n4256 | 2_n4467;
assign 2_n2563 = 2_n2108 & 2_n5590;
assign 2_n6651 = 2_n2285 & 2_n2525;
assign 2_n12670 = 2_n1445 & 2_n5727;
assign 2_n6363 = 2_n4356 & 2_n6210;
assign 2_n9064 = 2_n2413 & 2_n10802;
assign 2_n10311 = ~2_n4436;
assign 2_n747 = ~(2_n7772 ^ 2_n5421);
assign 2_n10133 = 2_n11266 & 2_n8286;
assign 2_n9945 = ~(2_n12951 ^ 2_n12840);
assign 2_n9035 = ~(2_n10413 ^ 2_n12254);
assign 2_n11459 = 2_n7690 & 2_n1564;
assign 2_n1282 = 2_n6696 | 2_n1938;
assign 2_n9042 = ~(2_n9328 ^ 2_n11826);
assign 2_n11057 = 2_n1903 | 2_n3332;
assign 2_n12839 = 2_n2893 | 2_n1014;
assign 2_n4677 = ~2_n1500;
assign 2_n6788 = 2_n6373 | 2_n7506;
assign 2_n1330 = 2_n10349 | 2_n7328;
assign 2_n721 = ~(2_n11099 ^ 2_n3288);
assign 2_n11622 = ~(2_n12088 | 2_n3490);
assign 2_n6946 = 2_n2456 | 2_n530;
assign 2_n2151 = ~(2_n4365 | 2_n4323);
assign 2_n9606 = ~(2_n6816 ^ 2_n7132);
assign 2_n4355 = 2_n5445 | 2_n9215;
assign 2_n7597 = ~(2_n9250 ^ 2_n12117);
assign 2_n201 = ~2_n6239;
assign 2_n444 = 2_n9122 | 2_n4460;
assign 2_n8654 = ~(2_n7306 ^ 2_n10584);
assign 2_n10791 = 2_n8810 | 2_n318;
assign 2_n8688 = 2_n5101 & 2_n9206;
assign 2_n1978 = 2_n7686 | 2_n6074;
assign 2_n10825 = 2_n7100 & 2_n9714;
assign 2_n2606 = 2_n7083 | 2_n672;
assign 2_n1375 = 2_n2285 | 2_n2525;
assign 2_n3236 = 2_n752 | 2_n3903;
assign 2_n10609 = 2_n724 | 2_n8022;
assign 2_n8788 = ~(2_n983 ^ 2_n4109);
assign 2_n12365 = 2_n3746 | 2_n3903;
assign 2_n8907 = 2_n2613 & 2_n3826;
assign 2_n2123 = 2_n8870 | 2_n8740;
assign 2_n6693 = 2_n9364 & 2_n1458;
assign 2_n1473 = 2_n9170 | 2_n4242;
assign 2_n3604 = 2_n7862 & 2_n3932;
assign 2_n10007 = ~2_n7616;
assign 2_n2504 = ~2_n11754;
assign 2_n5666 = ~2_n11184;
assign 2_n1354 = 2_n5765 | 2_n9078;
assign 2_n6367 = ~(2_n7019 ^ 2_n9666);
assign 2_n791 = 2_n3618 ^ 2_n11585;
assign 2_n988 = 2_n11531 | 2_n10295;
assign 2_n10905 = 2_n9021 | 2_n4170;
assign 2_n7587 = 2_n7283 | 2_n1915;
assign 2_n4391 = ~2_n6905;
assign 2_n1733 = 2_n4426 & 2_n1225;
assign 2_n12515 = ~(2_n9179 ^ 2_n4217);
assign 2_n6339 = 2_n4059 | 2_n10066;
assign 2_n8607 = ~2_n8634;
assign 2_n12243 = 2_n10169 | 2_n1411;
assign 2_n2018 = 2_n7306 | 2_n10584;
assign 2_n2248 = ~(2_n161 | 2_n550);
assign 2_n12892 = 2_n1814 | 2_n739;
assign 2_n7547 = ~(2_n6551 ^ 2_n8243);
assign 2_n5553 = ~(2_n7569 ^ 2_n12207);
assign 2_n2554 = ~(2_n8262 ^ 2_n11093);
assign 2_n704 = ~(2_n9201 ^ 2_n5911);
assign 2_n1345 = ~2_n3166;
assign 2_n4592 = 2_n1539 | 2_n4400;
assign 2_n1522 = ~(2_n10417 ^ 2_n3660);
assign 2_n6936 = ~(2_n5181 ^ 2_n3410);
assign 2_n3097 = ~(2_n8983 | 2_n4172);
assign 2_n1584 = 2_n2650 & 2_n9728;
assign 2_n10427 = ~(2_n4384 ^ 2_n6587);
assign 2_n974 = 2_n7221 & 2_n6453;
assign 2_n3913 = 2_n1183 | 2_n5468;
assign 2_n2934 = 2_n1936 & 2_n6723;
assign 2_n5858 = ~2_n10547;
assign 2_n12360 = ~(2_n3460 ^ 2_n12229);
assign 2_n3380 = ~(2_n5533 | 2_n7726);
assign 2_n799 = ~2_n10964;
assign 2_n7651 = 2_n7391 | 2_n12328;
assign 2_n1172 = 2_n7992 | 2_n8569;
assign 2_n6151 = 2_n5994 & 2_n8722;
assign 2_n8322 = 2_n10309 | 2_n11180;
assign 2_n11015 = 2_n11674 | 2_n2726;
assign 2_n1529 = 2_n4071 | 2_n5612;
assign 2_n537 = 2_n1937 | 2_n11122;
assign 2_n9631 = 2_n7564 & 2_n1363;
assign 2_n7006 = 2_n5596 | 2_n6829;
assign 2_n10829 = 2_n9791 | 2_n10393;
assign 2_n5380 = 2_n8026 | 2_n6169;
assign 2_n5692 = ~(2_n4806 ^ 2_n6236);
assign 2_n8800 = 2_n8020 & 2_n1644;
assign 2_n12200 = 2_n5507 & 2_n5045;
assign 2_n10099 = ~(2_n12423 ^ 2_n7303);
assign 2_n8960 = ~(2_n12597 ^ 2_n5313);
assign 2_n8869 = 2_n1941 | 2_n6169;
assign 2_n629 = ~2_n11913;
assign 2_n10884 = ~(2_n6830 ^ 2_n9316);
assign 2_n3222 = ~(2_n12353 ^ 2_n2350);
assign 2_n11177 = 2_n6718 | 2_n2020;
assign 2_n10362 = ~(2_n6989 ^ 2_n4836);
assign 2_n8515 = 2_n7678 & 2_n1526;
assign 2_n12415 = ~(2_n12466 ^ 2_n8960);
assign 2_n1832 = 2_n5120 | 2_n174;
assign 2_n12328 = ~2_n9195;
assign 2_n5637 = 2_n3453 | 2_n2809;
assign 2_n3995 = 2_n998 & 2_n4129;
assign 2_n11330 = 2_n5031 | 2_n6798;
assign 2_n11682 = ~(2_n3058 | 2_n5901);
assign 2_n11615 = ~(2_n4061 | 2_n10437);
assign 2_n8816 = 2_n1937 | 2_n11896;
assign 2_n3699 = 2_n4131 | 2_n10190;
assign 2_n6452 = ~(2_n605 | 2_n9288);
assign 2_n9490 = ~2_n9544;
assign 2_n2051 = ~(2_n8839 ^ 2_n5774);
assign 2_n3318 = 2_n855 | 2_n10699;
assign 2_n12503 = ~2_n5319;
assign 2_n5444 = ~(2_n8315 ^ 2_n2789);
assign 2_n7118 = ~(2_n6244 | 2_n8180);
assign 2_n1777 = 2_n5013 & 2_n3588;
assign 2_n8787 = ~2_n10116;
assign 2_n9618 = ~2_n3762;
assign 2_n729 = ~(2_n11409 ^ 2_n9032);
assign 2_n1681 = ~(2_n7458 ^ 2_n11748);
assign 2_n7181 = 2_n1249 | 2_n7963;
assign 2_n547 = ~(2_n2684 ^ 2_n5103);
assign 2_n3695 = 2_n4798 | 2_n4368;
assign 2_n2572 = 2_n4286 & 2_n8472;
assign 2_n7379 = ~2_n8225;
assign 2_n7576 = ~(2_n8184 ^ 2_n10655);
assign 2_n9296 = ~(2_n5338 | 2_n8933);
assign 2_n10119 = 2_n4911 | 2_n2358;
assign 2_n12899 = ~2_n10391;
assign 2_n1294 = ~(2_n6392 ^ 2_n4090);
assign 2_n10601 = ~(2_n6946 ^ 2_n9104);
assign 2_n2550 = 2_n12819 & 2_n3379;
assign 2_n7098 = ~(2_n5097 | 2_n9773);
assign 2_n7291 = ~(2_n2148 | 2_n5275);
assign 2_n9501 = ~(2_n9365 ^ 2_n3307);
assign 2_n2900 = 2_n7802 & 2_n7141;
assign 2_n3756 = 2_n10502 | 2_n6189;
assign 2_n11938 = ~(2_n11545 ^ 2_n5067);
assign 2_n4067 = ~(2_n8072 ^ 2_n11527);
assign 2_n8400 = ~(2_n7271 ^ 2_n11263);
assign 2_n1020 = 2_n2177 ^ 2_n1150;
assign 2_n9226 = 2_n7116 | 2_n2232;
assign 2_n2222 = ~(2_n7286 ^ 2_n7443);
assign 2_n8718 = ~2_n2408;
assign 2_n448 = 2_n11543 & 2_n3378;
assign 2_n2052 = ~2_n1105;
assign 2_n11322 = 2_n8118 & 2_n9965;
assign 2_n8351 = ~(2_n7071 ^ 2_n8338);
assign 2_n162 = ~(2_n8835 ^ 2_n8793);
assign 2_n4590 = ~(2_n2448 ^ 2_n12070);
assign 2_n3077 = ~(2_n11828 ^ 2_n5133);
assign 2_n9161 = ~2_n9416;
assign 2_n7575 = 2_n7133 & 2_n2395;
assign 2_n5991 = ~2_n7826;
assign 2_n11756 = 2_n6352 & 2_n1533;
assign 2_n7177 = 2_n5767 & 2_n5760;
assign 2_n10285 = ~(2_n8714 ^ 2_n10468);
assign 2_n12453 = ~2_n458;
assign 2_n9185 = ~2_n10604;
assign 2_n8723 = ~(2_n6933 ^ 2_n3994);
assign 2_n12772 = ~2_n8323;
assign 2_n6112 = ~(2_n2180 ^ 2_n927);
assign 2_n6971 = ~(2_n6121 | 2_n5946);
assign 2_n3862 = ~2_n9099;
assign 2_n2094 = ~(2_n10922 ^ 2_n11650);
assign 2_n3376 = 2_n580 & 2_n2469;
assign 2_n8116 = 2_n8583 | 2_n1476;
assign 2_n6393 = ~(2_n4892 | 2_n583);
assign 2_n6433 = ~2_n535;
assign 2_n7819 = ~(2_n11875 | 2_n1408);
assign 2_n6561 = 2_n8870 | 2_n9188;
assign 2_n4246 = 2_n4628 | 2_n12883;
assign 2_n11528 = 2_n4561 | 2_n10280;
assign 2_n2960 = ~(2_n2909 ^ 2_n6280);
assign 2_n6948 = 2_n2630 | 2_n5324;
assign 2_n9337 = ~(2_n2405 ^ 2_n10090);
assign 2_n719 = 2_n7862 & 2_n4921;
assign 2_n11062 = ~(2_n5166 ^ 2_n4285);
assign 2_n9489 = 2_n2653 & 2_n12359;
assign 2_n872 = 2_n5915 | 2_n8648;
assign 2_n10689 = 2_n2293 & 2_n10956;
assign 2_n706 = 2_n12594 | 2_n5469;
assign 2_n2142 = ~(2_n8473 | 2_n2442);
assign 2_n8823 = 2_n7578 & 2_n3644;
assign 2_n9344 = ~2_n2047;
assign 2_n456 = ~(2_n3262 ^ 2_n4072);
assign 2_n5307 = ~2_n9443;
assign 2_n528 = ~(2_n4379 ^ 2_n11693);
assign 2_n4426 = 2_n7100 | 2_n9714;
assign 2_n3480 = 2_n2830 | 2_n4405;
assign 2_n6709 = 2_n9920 & 2_n5212;
assign 2_n4415 = 2_n11026 | 2_n9160;
assign 2_n7192 = ~(2_n5695 | 2_n6745);
assign 2_n11059 = ~(2_n10996 | 2_n8292);
assign 2_n3910 = ~(2_n12630 ^ 2_n5074);
assign 2_n6670 = 2_n4393 & 2_n4829;
assign 2_n3825 = 2_n1581 & 2_n437;
assign 2_n349 = 2_n1699 | 2_n12080;
assign 2_n3943 = ~2_n7831;
assign 2_n7362 = ~(2_n4019 ^ 2_n2027);
assign 2_n12949 = ~(2_n10034 ^ 2_n5413);
assign 2_n430 = 2_n2456 | 2_n10854;
assign 2_n1424 = 2_n1714 & 2_n2592;
assign 2_n7099 = 2_n3746 | 2_n3356;
assign 2_n8271 = ~(2_n8166 ^ 2_n3253);
assign 2_n5980 = ~(2_n2416 ^ 2_n9088);
assign 2_n7078 = 2_n6577 | 2_n7876;
assign 2_n6044 = 2_n7487 | 2_n7752;
assign 2_n7043 = 2_n5860 & 2_n9111;
assign 2_n2624 = ~(2_n651 ^ 2_n10687);
assign 2_n4280 = ~2_n10178;
assign 2_n11532 = 2_n1941 | 2_n12816;
assign 2_n3596 = ~(2_n10228 | 2_n11971);
assign 2_n6677 = 2_n10057 | 2_n5822;
assign 2_n2963 = 2_n5765 | 2_n12771;
assign 2_n8773 = 2_n12243 & 2_n11331;
assign 2_n11523 = ~(2_n3000 ^ 2_n6639);
assign 2_n5876 = ~2_n7377;
assign 2_n1781 = ~2_n4522;
assign 2_n94 = ~(2_n10686 ^ 2_n8935);
assign 2_n369 = ~(2_n6066 ^ 2_n8814);
assign 2_n7585 = ~(2_n4107 ^ 2_n11695);
assign 2_n10305 = 2_n2670 | 2_n10220;
assign 2_n7985 = ~(2_n2216 ^ 2_n2810);
assign 2_n10073 = 2_n3433 & 2_n1722;
assign 2_n508 = 2_n7862 & 2_n11407;
assign 2_n7359 = ~(2_n10210 ^ 2_n8366);
assign 2_n4047 = 2_n10926 | 2_n11396;
assign 2_n12123 = ~(2_n12379 ^ 2_n1429);
assign 2_n9676 = ~(2_n494 ^ 2_n2070);
assign 2_n12775 = 2_n4059 | 2_n7424;
assign 2_n475 = ~(2_n9413 ^ 2_n9022);
assign 2_n9546 = ~(2_n11788 ^ 2_n3641);
assign 2_n8004 = 2_n744 | 2_n11432;
assign 2_n2890 = 2_n12503 | 2_n9521;
assign 2_n7658 = 2_n648 & 2_n6769;
assign 2_n5102 = 2_n10530 | 2_n1038;
assign 2_n2104 = ~(2_n10461 ^ 2_n12523);
assign 2_n7554 = 2_n2575 & 2_n175;
assign 2_n423 = ~2_n7023;
assign 2_n9781 = 2_n3954 & 2_n8955;
assign 2_n4930 = ~(2_n4893 ^ 2_n5085);
assign 2_n6787 = 2_n3961 & 2_n9219;
assign 2_n2995 = 2_n8129 | 2_n12603;
assign 2_n8202 = ~(2_n3296 ^ 2_n5557);
assign 2_n2794 = ~(2_n3297 | 2_n12424);
assign 2_n6288 = ~2_n1190;
assign 2_n12556 = ~(2_n2702 | 2_n449);
assign 2_n8362 = ~(2_n3128 ^ 2_n12381);
assign 2_n1637 = ~(2_n10023 ^ 2_n11085);
assign 2_n3545 = ~(2_n8142 | 2_n6308);
assign 2_n2578 = ~2_n9216;
assign 2_n11983 = ~(2_n3991 ^ 2_n12154);
assign 2_n7036 = ~(2_n4904 ^ 2_n5493);
assign 2_n1591 = 2_n10262 | 2_n5630;
assign 2_n12287 = ~(2_n6544 ^ 2_n6435);
assign 2_n1370 = 2_n7839 | 2_n1413;
assign 2_n3559 = ~(2_n4114 ^ 2_n7336);
assign 2_n10348 = 2_n905 & 2_n11505;
assign 2_n1316 = 2_n2619 & 2_n4978;
assign 2_n1073 = 2_n8789 | 2_n1733;
assign 2_n2977 = ~2_n9683;
assign 2_n2582 = ~2_n8763;
assign 2_n10370 = 2_n2911 | 2_n4530;
assign 2_n4809 = ~(2_n11534 ^ 2_n9184);
assign 2_n10385 = 2_n8814 | 2_n6278;
assign 2_n3847 = ~(2_n7157 | 2_n6746);
assign 2_n5112 = ~(2_n5578 ^ 2_n780);
assign 2_n8284 = 2_n6386 & 2_n3841;
assign 2_n1015 = ~(2_n4566 ^ 2_n10370);
assign 2_n5175 = ~(2_n382 ^ 2_n1060);
assign 2_n8163 = ~(2_n8239 ^ 2_n11857);
assign 2_n12572 = ~(2_n6650 ^ 2_n305);
assign 2_n2583 = ~(2_n10269 ^ 2_n5295);
assign 2_n7441 = 2_n1051 | 2_n7952;
assign 2_n3994 = ~(2_n10092 | 2_n1666);
assign 2_n3796 = 2_n12552 | 2_n6989;
assign 2_n6635 = 2_n8187 | 2_n7341;
assign 2_n1299 = ~(2_n3244 | 2_n6024);
assign 2_n3409 = 2_n5450 | 2_n6694;
assign 2_n3720 = ~(2_n10761 ^ 2_n3234);
assign 2_n12505 = ~(2_n9572 ^ 2_n6711);
assign 2_n7824 = ~(2_n4259 ^ 2_n10003);
assign 2_n5434 = ~2_n8347;
assign 2_n10459 = ~(2_n6570 ^ 2_n8478);
assign 2_n3554 = ~(2_n7441 ^ 2_n3009);
assign 2_n1350 = 2_n9677 & 2_n12869;
assign 2_n9238 = ~(2_n4788 ^ 2_n2787);
assign 2_n10529 = 2_n4059 | 2_n6402;
assign 2_n4684 = 2_n9299 & 2_n11158;
assign 2_n7850 = 2_n6002 & 2_n9590;
assign 2_n1948 = ~(2_n816 ^ 2_n7530);
assign 2_n579 = ~(2_n2856 ^ 2_n3165);
assign 2_n6894 = 2_n11552 | 2_n1047;
assign 2_n9967 = ~(2_n3895 ^ 2_n1729);
assign 2_n6641 = ~(2_n6488 ^ 2_n5731);
assign 2_n5469 = 2_n2249 & 2_n1676;
assign 2_n8897 = ~(2_n12399 | 2_n4889);
assign 2_n8312 = 2_n12098 & 2_n5499;
assign 2_n11497 = ~2_n4089;
assign 2_n34 = ~(2_n64 | 2_n5143);
assign 2_n11185 = ~(2_n10575 ^ 2_n3187);
assign 2_n8613 = 2_n11616 & 2_n3023;
assign 2_n2400 = 2_n5355 | 2_n12328;
assign 2_n5451 = ~(2_n4562 ^ 2_n12689);
assign 2_n8468 = ~(2_n4237 ^ 2_n12852);
assign 2_n7721 = ~(2_n3858 ^ 2_n9738);
assign 2_n6323 = ~2_n525;
assign 2_n4265 = 2_n5915 | 2_n8644;
assign 2_n9816 = 2_n8206 | 2_n3195;
assign 2_n5067 = 2_n2816 & 2_n9378;
assign 2_n5321 = 2_n254 | 2_n7775;
assign 2_n5484 = 2_n180 | 2_n285;
assign 2_n655 = ~(2_n6045 ^ 2_n6432);
assign 2_n4593 = ~2_n2485;
assign 2_n7736 = 2_n8835 & 2_n9595;
assign 2_n6898 = 2_n2308 & 2_n11133;
assign 2_n176 = ~(2_n4620 ^ 2_n9912);
assign 2_n9594 = ~(2_n1712 ^ 2_n11632);
assign 2_n1667 = ~2_n8319;
assign 2_n12578 = 2_n7111 | 2_n11131;
assign 2_n8836 = ~(2_n11395 ^ 2_n4735);
assign 2_n11690 = 2_n1051 | 2_n7558;
assign 2_n9407 = ~(2_n8692 ^ 2_n2421);
assign 2_n1255 = ~(2_n5808 ^ 2_n7573);
assign 2_n11342 = ~(2_n6018 ^ 2_n5892);
assign 2_n9900 = ~(2_n2492 ^ 2_n12099);
assign 2_n2844 = ~2_n10013;
assign 2_n7403 = ~(2_n2332 ^ 2_n6034);
assign 2_n7050 = ~2_n2602;
assign 2_n8539 = ~2_n1420;
assign 2_n7703 = ~2_n2508;
assign 2_n4245 = ~(2_n10838 ^ 2_n3060);
assign 2_n5670 = ~(2_n5649 ^ 2_n3004);
assign 2_n6819 = ~(2_n2073 | 2_n12028);
assign 2_n4881 = 2_n8705 | 2_n12336;
assign 2_n1300 = 2_n398 & 2_n2322;
assign 2_n10344 = 2_n1442 & 2_n3668;
assign 2_n12514 = 2_n12840 | 2_n12951;
assign 2_n1764 = ~(2_n6612 | 2_n4896);
assign 2_n4477 = ~(2_n2943 ^ 2_n11097);
assign 2_n1014 = 2_n7283 | 2_n12843;
assign 2_n2591 = 2_n5786 | 2_n9464;
assign 2_n6337 = ~(2_n4438 ^ 2_n12498);
assign 2_n3837 = ~(2_n7507 ^ 2_n7658);
assign 2_n7938 = ~2_n11526;
assign 2_n5186 = 2_n10739 & 2_n3938;
assign 2_n3551 = ~(2_n10249 ^ 2_n12082);
assign 2_n1419 = ~(2_n3565 ^ 2_n1894);
assign 2_n12379 = 2_n9696 | 2_n6394;
assign 2_n1516 = 2_n9953 & 2_n6396;
assign 2_n3060 = 2_n7964 & 2_n9329;
assign 2_n2573 = 2_n6251 | 2_n3403;
assign 2_n11766 = ~(2_n2531 ^ 2_n9945);
assign 2_n1314 = 2_n2511 & 2_n926;
assign 2_n9943 = ~(2_n11541 ^ 2_n4936);
assign 2_n2503 = 2_n12503 | 2_n1047;
assign 2_n7949 = ~2_n2467;
assign 2_n9460 = ~(2_n5 ^ 2_n3720);
assign 2_n6768 = 2_n7965 & 2_n11876;
assign 2_n3804 = 2_n2437 & 2_n2085;
assign 2_n11809 = ~(2_n6424 ^ 2_n1332);
assign 2_n7867 = ~(2_n11408 ^ 2_n12450);
assign 2_n2605 = ~(2_n7956 ^ 2_n11251);
assign 2_n4645 = ~2_n8843;
assign 2_n1638 = 2_n8267 & 2_n11939;
assign 2_n9714 = 2_n8428 | 2_n5540;
assign 2_n9983 = ~(2_n7659 ^ 2_n117);
assign 2_n1928 = 2_n2267 | 2_n1096;
assign 2_n10381 = 2_n2456 | 2_n2964;
assign 2_n2470 = 2_n5305 & 2_n3932;
assign 2_n570 = ~(2_n10071 | 2_n1604);
assign 2_n12724 = ~2_n3728;
assign 2_n3253 = 2_n8026 | 2_n12899;
assign 2_n3054 = ~(2_n11715 ^ 2_n12575);
assign 2_n10552 = ~(2_n4739 | 2_n1846);
assign 2_n59 = ~(2_n5598 ^ 2_n11672);
assign 2_n11034 = 2_n7914 & 2_n4351;
assign 2_n4408 = ~(2_n12513 | 2_n12690);
assign 2_n10948 = ~(2_n9250 | 2_n10453);
assign 2_n2831 = ~(2_n6381 ^ 2_n4404);
assign 2_n4401 = 2_n6660 & 2_n5406;
assign 2_n10347 = 2_n6977 | 2_n11820;
assign 2_n10172 = 2_n8552 | 2_n7928;
assign 2_n646 = 2_n3743 | 2_n6138;
assign 2_n7060 = 2_n12155 & 2_n6473;
assign 2_n11196 = 2_n10500 | 2_n974;
assign 2_n2265 = ~(2_n1006 | 2_n9217);
assign 2_n3639 = ~(2_n8029 ^ 2_n9423);
assign 2_n9052 = 2_n3604 & 2_n4421;
assign 2_n3503 = ~(2_n5936 | 2_n2998);
assign 2_n3311 = 2_n4092 | 2_n5907;
assign 2_n10780 = ~2_n12623;
assign 2_n3771 = ~(2_n1776 ^ 2_n9452);
assign 2_n12281 = 2_n2099 | 2_n10311;
assign 2_n5467 = ~(2_n9860 ^ 2_n9100);
assign 2_n1594 = 2_n2393 & 2_n11791;
assign 2_n11993 = 2_n6303 | 2_n8084;
assign 2_n2638 = 2_n11380 | 2_n11115;
assign 2_n7493 = ~(2_n4171 ^ 2_n10077);
assign 2_n7720 = 2_n5961 & 2_n2804;
assign 2_n9428 = 2_n191 | 2_n7246;
assign 2_n7929 = ~(2_n1240 ^ 2_n10183);
assign 2_n11137 = ~2_n11777;
assign 2_n8417 = ~(2_n8824 ^ 2_n7272);
assign 2_n3783 = ~(2_n4718 ^ 2_n11260);
assign 2_n6925 = ~2_n3633;
assign 2_n3883 = ~(2_n12291 ^ 2_n923);
assign 2_n8355 = 2_n10222 & 2_n3828;
assign 2_n6003 = 2_n1937 | 2_n3903;
assign 2_n9987 = ~(2_n2618 | 2_n1654);
assign 2_n2757 = ~(2_n10057 ^ 2_n5399);
assign 2_n156 = ~2_n9010;
assign 2_n12250 = ~(2_n7595 ^ 2_n4709);
assign 2_n2308 = 2_n2548 | 2_n8435;
assign 2_n3003 = 2_n186 & 2_n3435;
assign 2_n12381 = ~(2_n2852 ^ 2_n1789);
assign 2_n4106 = ~(2_n11684 ^ 2_n10731);
assign 2_n2581 = ~(2_n3945 ^ 2_n7259);
assign 2_n4708 = ~(2_n12841 ^ 2_n6563);
assign 2_n7800 = ~2_n8779;
assign 2_n10261 = 2_n4185 | 2_n4965;
assign 2_n5237 = 2_n10079 | 2_n10538;
assign 2_n743 = ~(2_n4211 | 2_n6259);
assign 2_n7732 = ~2_n7814;
assign 2_n9905 = 2_n10835 | 2_n9568;
assign 2_n9918 = 2_n4628 | 2_n4913;
assign 2_n3001 = ~(2_n5872 ^ 2_n9018);
assign 2_n10275 = ~2_n4034;
assign 2_n1337 = 2_n1223 | 2_n2892;
assign 2_n2311 = ~(2_n4899 ^ 2_n4329);
assign 2_n2499 = ~2_n613;
assign 2_n3035 = ~(2_n6771 ^ 2_n9662);
assign 2_n3114 = 2_n10605 | 2_n3388;
assign 2_n8721 = ~(2_n70 ^ 2_n11210);
assign 2_n10726 = 2_n5809 | 2_n12686;
assign 2_n5813 = 2_n8822 | 2_n4472;
assign 2_n2634 = 2_n12708 & 2_n9745;
assign 2_n12767 = 2_n196 | 2_n11477;
assign 2_n6246 = ~(2_n12074 ^ 2_n1540);
assign 2_n11087 = ~(2_n9810 | 2_n11696);
assign 2_n5604 = ~(2_n11281 ^ 2_n4629);
assign 2_n12066 = ~(2_n8919 | 2_n1582);
assign 2_n828 = ~(2_n7400 ^ 2_n10089);
assign 2_n7557 = 2_n114 | 2_n11775;
assign 2_n11946 = ~(2_n3420 ^ 2_n594);
assign 2_n10187 = 2_n10088 & 2_n3295;
assign 2_n3249 = ~2_n6884;
assign 2_n7484 = ~(2_n4630 ^ 2_n7722);
assign 2_n11735 = 2_n2042 & 2_n10305;
assign 2_n96 = 2_n4502 | 2_n9610;
assign 2_n1627 = 2_n2424 | 2_n12846;
assign 2_n11452 = 2_n10355 | 2_n5863;
assign 2_n11130 = ~(2_n8017 ^ 2_n3364);
assign 2_n2666 = ~(2_n5756 ^ 2_n11913);
assign 2_n9548 = ~2_n11934;
assign 2_n10448 = 2_n10879 | 2_n3911;
assign 2_n12797 = ~2_n7523;
assign 2_n7263 = ~(2_n6812 ^ 2_n12018);
assign 2_n3624 = ~2_n933;
assign 2_n11758 = 2_n8961 & 2_n3193;
assign 2_n10499 = 2_n2262 & 2_n2066;
assign 2_n6892 = ~(2_n11289 ^ 2_n11024);
assign 2_n2042 = 2_n2536 | 2_n12112;
assign 2_n8503 = ~(2_n7393 | 2_n12362);
assign 2_n9650 = ~2_n1;
assign 2_n1913 = 2_n5859 & 2_n11824;
assign 2_n8130 = ~(2_n12409 ^ 2_n11258);
assign 2_n5969 = 2_n9878 | 2_n1932;
assign 2_n733 = ~(2_n5167 ^ 2_n11781);
assign 2_n768 = ~(2_n5852 ^ 2_n4095);
assign 2_n9992 = ~(2_n683 ^ 2_n12953);
assign 2_n3892 = ~(2_n5594 | 2_n11095);
assign 2_n4501 = 2_n1699 | 2_n10422;
assign 2_n5725 = ~2_n11141;
assign 2_n8196 = ~(2_n3115 ^ 2_n4853);
assign 2_n7204 = 2_n114 | 2_n2232;
assign 2_n299 = ~2_n3874;
assign 2_n11078 = 2_n10194 | 2_n9928;
assign 2_n2576 = ~(2_n1995 | 2_n464);
assign 2_n4084 = ~2_n6174;
assign 2_n12548 = ~(2_n6272 ^ 2_n2126);
assign 2_n12347 = 2_n1122 & 2_n12427;
assign 2_n10304 = ~2_n2924;
assign 2_n7589 = ~(2_n2871 ^ 2_n6415);
assign 2_n10002 = 2_n962 | 2_n3606;
assign 2_n11668 = 2_n5394 | 2_n5152;
assign 2_n5225 = ~(2_n3420 | 2_n7634);
assign 2_n669 = 2_n6462 & 2_n7742;
assign 2_n5871 = ~2_n3479;
assign 2_n12829 = 2_n430 | 2_n10085;
assign 2_n2671 = 2_n6256 & 2_n7489;
assign 2_n2730 = ~2_n10061;
assign 2_n311 = ~2_n399;
assign 2_n6962 = ~(2_n7594 | 2_n4902);
assign 2_n12801 = ~2_n3087;
assign 2_n10971 = ~(2_n4697 ^ 2_n6430);
assign 2_n10296 = 2_n11449 & 2_n1365;
assign 2_n5095 = 2_n1809 & 2_n882;
assign 2_n165 = 2_n10142 | 2_n3911;
assign 2_n11594 = 2_n12662 | 2_n10491;
assign 2_n7212 = ~2_n5758;
assign 2_n2354 = 2_n9787 | 2_n7619;
assign 2_n2068 = 2_n1561 | 2_n12817;
assign 2_n1671 = ~(2_n8227 ^ 2_n10209);
assign 2_n38 = ~(2_n12426 ^ 2_n12085);
assign 2_n8114 = ~2_n2307;
assign 2_n7094 = 2_n3413 | 2_n4877;
assign 2_n11157 = ~(2_n10541 ^ 2_n8852);
assign 2_n5961 = ~2_n12746;
assign 2_n10431 = ~(2_n9570 ^ 2_n12050);
assign 2_n1418 = 2_n7593 & 2_n3377;
assign 2_n10719 = 2_n9929 & 2_n4842;
assign 2_n3985 = ~(2_n6727 ^ 2_n9439);
assign 2_n5788 = ~2_n7667;
assign 2_n853 = ~(2_n6773 ^ 2_n9419);
assign 2_n9984 = ~(2_n2947 ^ 2_n6033);
assign 2_n122 = ~(2_n6825 ^ 2_n6100);
assign 2_n10800 = ~(2_n4637 ^ 2_n4454);
assign 2_n1404 = 2_n7749 & 2_n8602;
assign 2_n8622 = ~2_n7820;
assign 2_n5437 = ~(2_n10433 | 2_n4485);
assign 2_n3178 = 2_n8678 & 2_n10154;
assign 2_n12602 = ~2_n11942;
assign 2_n12476 = 2_n4698 & 2_n3815;
assign 2_n12784 = 2_n1319 | 2_n3417;
assign 2_n7459 = ~(2_n6788 ^ 2_n4495);
assign 2_n9477 = ~(2_n6896 | 2_n9856);
assign 2_n374 = 2_n1111 | 2_n11177;
assign 2_n12723 = 2_n9373 | 2_n10916;
assign 2_n10437 = 2_n3116 & 2_n9931;
assign 2_n6832 = 2_n5816 & 2_n6522;
assign 2_n7722 = ~(2_n1415 ^ 2_n4431);
assign 2_n9521 = ~2_n8433;
assign 2_n110 = ~(2_n7792 ^ 2_n12048);
assign 2_n2152 = ~(2_n8329 ^ 2_n6434);
assign 2_n5775 = ~(2_n8896 ^ 2_n4710);
assign 2_n7611 = 2_n4380 & 2_n5245;
assign 2_n4669 = ~(2_n9898 ^ 2_n1513);
assign 2_n2425 = ~(2_n85 ^ 2_n2884);
assign 2_n6567 = ~(2_n3784 | 2_n3317);
assign 2_n7339 = 2_n6909 & 2_n845;
assign 2_n6022 = ~(2_n11752 | 2_n11781);
assign 2_n3562 = ~(2_n5396 | 2_n6757);
assign 2_n8968 = ~(2_n356 ^ 2_n3398);
assign 2_n4389 = 2_n989 | 2_n1738;
assign 2_n7900 = 2_n3820 | 2_n10916;
assign 2_n8268 = 2_n114 | 2_n6455;
assign 2_n8368 = 2_n7112 | 2_n7795;
assign 2_n9350 = ~2_n6947;
assign 2_n9741 = ~2_n6429;
assign 2_n9591 = 2_n6317 & 2_n12929;
assign 2_n5306 = 2_n4059 | 2_n12843;
assign 2_n5612 = 2_n11801 & 2_n10413;
assign 2_n6329 = 2_n8598 | 2_n5581;
assign 2_n1226 = 2_n11867 | 2_n6075;
assign 2_n6120 = ~(2_n2541 ^ 2_n10427);
assign 2_n7864 = 2_n4628 | 2_n5326;
assign 2_n11165 = ~2_n8973;
assign 2_n10795 = 2_n5250 & 2_n2214;
assign 2_n3854 = ~(2_n8765 ^ 2_n29);
assign 2_n3958 = ~2_n5041;
assign 2_n1045 = ~(2_n2700 ^ 2_n566);
assign 2_n7109 = 2_n11652 | 2_n5939;
assign 2_n8401 = 2_n8687 | 2_n1509;
assign 2_n5787 = ~2_n528;
assign 2_n1236 = 2_n6294 & 2_n1067;
assign 2_n9832 = ~(2_n5576 ^ 2_n4353);
assign 2_n510 = ~2_n11662;
assign 2_n10755 = ~2_n2233;
assign 2_n11603 = 2_n2123 | 2_n11101;
assign 2_n1742 = ~(2_n9753 | 2_n12671);
assign 2_n1237 = ~(2_n12584 ^ 2_n436);
assign 2_n3242 = ~2_n11936;
assign 2_n6838 = ~(2_n8475 ^ 2_n12600);
assign 2_n5298 = ~(2_n9341 ^ 2_n1765);
assign 2_n5544 = ~(2_n1334 ^ 2_n5566);
assign 2_n9995 = 2_n1183 | 2_n12080;
assign 2_n3800 = 2_n9530 | 2_n7879;
assign 2_n3591 = ~2_n11875;
assign 2_n2191 = 2_n4984 | 2_n9153;
assign 2_n11770 = ~(2_n3729 | 2_n10250);
assign 2_n3084 = 2_n1092 | 2_n3175;
assign 2_n7649 = ~2_n3089;
assign 2_n2155 = 2_n5355 | 2_n7881;
assign 2_n9222 = 2_n10196 | 2_n795;
assign 2_n12156 = 2_n4059 | 2_n11430;
assign 2_n3770 = ~(2_n5174 ^ 2_n6068);
assign 2_n1381 = ~(2_n12536 | 2_n883);
assign 2_n3174 = 2_n8262 | 2_n3085;
assign 2_n5432 = 2_n5575 | 2_n6455;
assign 2_n3518 = 2_n4325 | 2_n628;
assign 2_n4314 = 2_n137 & 2_n11922;
assign 2_n12226 = ~(2_n3863 ^ 2_n3293);
assign 2_n7517 = 2_n5087 & 2_n5357;
assign 2_n6528 = ~(2_n6662 ^ 2_n8311);
assign 2_n8153 = 2_n10844 | 2_n5699;
assign 2_n10271 = ~(2_n6834 ^ 2_n2996);
assign 2_n9556 = ~(2_n10605 ^ 2_n1964);
assign 2_n2476 = 2_n10545 & 2_n2498;
assign 2_n915 = ~(2_n3221 ^ 2_n7846);
assign 2_n5372 = ~2_n6361;
assign 2_n7758 = ~(2_n7909 ^ 2_n4432);
assign 2_n11861 = ~(2_n10666 ^ 2_n10431);
assign 2_n6640 = 2_n3699 & 2_n2733;
assign 2_n2271 = 2_n9131 & 2_n12463;
assign 2_n2286 = ~(2_n12235 | 2_n12154);
assign 2_n6873 = ~(2_n4057 ^ 2_n908);
assign 2_n10059 = 2_n3053 & 2_n7943;
assign 2_n6590 = 2_n994 | 2_n1851;
assign 2_n11436 = ~(2_n952 | 2_n9828);
assign 2_n9818 = ~2_n6440;
assign 2_n12471 = ~(2_n4602 ^ 2_n6980);
assign 2_n11650 = ~(2_n78 ^ 2_n1934);
assign 2_n5766 = ~2_n173;
assign 2_n12883 = ~2_n12044;
assign 2_n7004 = 2_n11417 & 2_n1314;
assign 2_n3341 = ~(2_n11523 | 2_n7973);
assign 2_n10701 = 2_n8113 & 2_n8626;
assign 2_n9877 = ~2_n10253;
assign 2_n10870 = 2_n800 & 2_n2468;
assign 2_n7286 = 2_n8738 | 2_n4527;
assign 2_n462 = ~(2_n9453 ^ 2_n9646);
assign 2_n9267 = ~(2_n5958 | 2_n4765);
assign 2_n4597 = 2_n5271 | 2_n2006;
assign 2_n1180 = 2_n11552 | 2_n5258;
assign 2_n8712 = ~(2_n3093 ^ 2_n6690);
assign 2_n7861 = ~2_n10378;
assign 2_n12074 = ~(2_n8751 ^ 2_n523);
assign 2_n7973 = ~2_n572;
assign 2_n9224 = ~(2_n7084 ^ 2_n9091);
assign 2_n5474 = ~2_n3931;
assign 2_n12530 = 2_n3743 | 2_n8285;
assign 2_n4638 = 2_n4546 | 2_n7545;
assign 2_n4691 = ~(2_n3088 ^ 2_n853);
assign 2_n6890 = 2_n9878 | 2_n4818;
assign 2_n12388 = ~2_n12099;
assign 2_n5839 = 2_n573 & 2_n11044;
assign 2_n2751 = 2_n10744 & 2_n2240;
assign 2_n6415 = ~(2_n4993 ^ 2_n6099);
assign 2_n6864 = 2_n9432 & 2_n7226;
assign 2_n7105 = 2_n7709 | 2_n795;
assign 2_n12736 = ~(2_n6145 ^ 2_n12101);
assign 2_n8259 = ~2_n12826;
assign 2_n4393 = 2_n351 | 2_n10275;
assign 2_n3161 = ~(2_n7019 | 2_n3782);
assign 2_n3150 = 2_n1051 | 2_n6169;
assign 2_n4514 = 2_n4858 & 2_n2243;
assign 2_n3246 = ~(2_n7652 ^ 2_n4830);
assign 2_n2457 = ~(2_n9935 ^ 2_n9488);
assign 2_n9101 = ~(2_n8911 ^ 2_n2734);
assign 2_n4473 = ~(2_n9900 ^ 2_n5063);
assign 2_n12135 = 2_n1768 | 2_n206;
assign 2_n5324 = ~(2_n5572 ^ 2_n12908);
assign 2_n4063 = ~(2_n6210 ^ 2_n6112);
assign 2_n5074 = ~(2_n8758 ^ 2_n12027);
assign 2_n1793 = ~(2_n3236 ^ 2_n1057);
assign 2_n10255 = 2_n6336 | 2_n4077;
assign 2_n8009 = ~(2_n7078 ^ 2_n838);
assign 2_n3904 = 2_n5314 & 2_n217;
assign 2_n5143 = ~(2_n6260 | 2_n2770);
assign 2_n6831 = 2_n8981 & 2_n4379;
assign 2_n3768 = ~2_n5368;
assign 2_n279 = 2_n5026 | 2_n9139;
assign 2_n9693 = ~(2_n12555 | 2_n9947);
assign 2_n2197 = 2_n6977 | 2_n12816;
assign 2_n7997 = 2_n8855 & 2_n10760;
assign 2_n6101 = ~(2_n5980 ^ 2_n3532);
assign 2_n4300 = ~(2_n9734 ^ 2_n2857);
assign 2_n10204 = ~(2_n8633 | 2_n5713);
assign 2_n219 = ~(2_n12832 | 2_n4271);
assign 2_n12414 = 2_n274 | 2_n11815;
assign 2_n9464 = 2_n2155 & 2_n11112;
assign 2_n9376 = 2_n8850 | 2_n10805;
assign 2_n7937 = ~(2_n8492 | 2_n6188);
assign 2_n3972 = ~(2_n8682 ^ 2_n6736);
assign 2_n807 = ~2_n7320;
assign 2_n7170 = ~2_n7526;
assign 2_n607 = 2_n5859 | 2_n11824;
assign 2_n6688 = ~(2_n354 ^ 2_n12793);
assign 2_n11329 = 2_n5204 & 2_n283;
assign 2_n7825 = 2_n5036 | 2_n2991;
assign 2_n3244 = 2_n12012 & 2_n11889;
assign 2_n2856 = ~(2_n8101 | 2_n10885);
assign 2_n11416 = ~(2_n866 ^ 2_n1580);
assign 2_n2502 = 2_n12361 | 2_n7395;
assign 2_n10787 = 2_n1867 & 2_n7371;
assign 2_n9349 = 2_n4465 | 2_n12916;
assign 2_n8868 = 2_n11074 & 2_n3652;
assign 2_n12904 = 2_n3256 & 2_n1081;
assign 2_n1901 = 2_n3210 & 2_n10527;
assign 2_n9473 = ~(2_n10927 ^ 2_n2051);
assign 2_n5710 = 2_n10117 | 2_n5140;
assign 2_n10748 = 2_n3816 & 2_n5228;
assign 2_n10469 = ~2_n190;
assign 2_n8217 = ~2_n2699;
assign 2_n6085 = ~(2_n1009 ^ 2_n1639);
assign 2_n215 = 2_n8941 & 2_n1418;
assign 2_n12820 = ~(2_n8308 ^ 2_n5607);
assign 2_n273 = 2_n7480 | 2_n1080;
assign 2_n9977 = ~(2_n4914 | 2_n4364);
assign 2_n4449 = ~2_n1229;
assign 2_n11677 = 2_n6185 & 2_n5017;
assign 2_n1537 = ~(2_n1809 | 2_n882);
assign 2_n5780 = 2_n5355 | 2_n2358;
assign 2_n740 = ~2_n11802;
assign 2_n5573 = 2_n5247 | 2_n9020;
assign 2_n10922 = 2_n636 | 2_n9188;
assign 2_n9685 = 2_n6579 | 2_n3093;
assign 2_n1446 = 2_n3698 & 2_n2394;
assign 2_n12581 = ~(2_n11867 ^ 2_n6475);
assign 2_n7847 = 2_n11678 | 2_n5805;
assign 2_n288 = 2_n11923 | 2_n1047;
assign 2_n4751 = ~(2_n1296 ^ 2_n12948);
assign 2_n6257 = ~2_n7869;
assign 2_n12380 = 2_n10435 | 2_n4895;
assign 2_n4223 = ~2_n11955;
assign 2_n12937 = ~(2_n2880 ^ 2_n792);
assign 2_n3348 = 2_n6666 & 2_n8991;
assign 2_n2039 = 2_n5959 & 2_n8534;
assign 2_n7631 = 2_n11577 & 2_n8053;
assign 2_n4621 = ~(2_n2275 ^ 2_n4543);
assign 2_n1508 = 2_n6191 & 2_n8895;
assign 2_n6211 = ~(2_n7396 | 2_n5885);
assign 2_n185 = ~(2_n6204 ^ 2_n11735);
assign 2_n2126 = ~(2_n1465 ^ 2_n848);
assign 2_n11077 = ~2_n150;
assign 2_n1890 = ~(2_n755 ^ 2_n3080);
assign 2_n8820 = ~(2_n8087 ^ 2_n10371);
assign 2_n11538 = 2_n752 | 2_n7425;
assign 2_n1961 = ~(2_n6454 ^ 2_n177);
assign 2_n3383 = ~2_n7459;
assign 2_n6662 = ~(2_n3359 | 2_n10047);
assign 2_n12361 = ~2_n12299;
assign 2_n6676 = ~(2_n11305 ^ 2_n10501);
assign 2_n9217 = ~(2_n3462 | 2_n7240);
assign 2_n5299 = 2_n825 | 2_n10284;
assign 2_n5580 = 2_n11221 & 2_n3260;
assign 2_n384 = ~(2_n10252 ^ 2_n8932);
assign 2_n748 = ~2_n9265;
assign 2_n12291 = ~(2_n2204 ^ 2_n751);
assign 2_n9953 = ~2_n6068;
assign 2_n1763 = ~(2_n1645 | 2_n11000);
assign 2_n262 = ~(2_n3723 ^ 2_n712);
assign 2_n6673 = 2_n5915 | 2_n10422;
assign 2_n1965 = ~(2_n929 | 2_n11453);
assign 2_n5040 = 2_n945 | 2_n4521;
assign 2_n2566 = ~(2_n804 ^ 2_n1716);
assign 2_n1230 = 2_n835 | 2_n7979;
assign 2_n4957 = 2_n8181 | 2_n8485;
assign 2_n7396 = 2_n1941 | 2_n7952;
assign 2_n33 = ~(2_n12365 ^ 2_n11406);
assign 2_n6577 = ~2_n2464;
assign 2_n2975 = ~(2_n5762 ^ 2_n6217);
assign 2_n5716 = ~(2_n11138 | 2_n10218);
assign 2_n864 = 2_n3996 | 2_n1046;
assign 2_n708 = 2_n8367 | 2_n388;
assign 2_n12286 = 2_n9843 & 2_n1066;
assign 2_n868 = ~(2_n9345 ^ 2_n3167);
assign 2_n1217 = 2_n2384 & 2_n3852;
assign 2_n3612 = 2_n3682 & 2_n8958;
assign 2_n5322 = ~(2_n6010 ^ 2_n2117);
assign 2_n12368 = ~(2_n9785 | 2_n574);
assign 2_n3109 = ~(2_n9187 ^ 2_n12113);
assign 2_n8594 = 2_n3743 | 2_n5759;
assign 2_n12071 = 2_n4773 & 2_n403;
assign 2_n3083 = 2_n938 & 2_n3311;
assign 2_n238 = ~(2_n4799 | 2_n7147);
assign 2_n11154 = 2_n11878 | 2_n10215;
assign 2_n12901 = ~(2_n5848 | 2_n3913);
assign 2_n12656 = ~(2_n4119 | 2_n378);
assign 2_n5635 = ~(2_n3667 ^ 2_n3090);
assign 2_n7826 = 2_n6877 & 2_n7354;
assign 2_n8770 = ~(2_n12271 | 2_n12707);
assign 2_n5077 = 2_n3791 | 2_n11806;
assign 2_n3386 = 2_n5530 | 2_n12446;
assign 2_n2580 = 2_n10682 | 2_n4011;
assign 2_n6383 = 2_n7441 & 2_n3009;
assign 2_n5745 = 2_n10239 & 2_n9325;
assign 2_n11189 = 2_n6877 & 2_n9640;
assign 2_n10879 = ~2_n3627;
assign 2_n10268 = ~(2_n6554 ^ 2_n5201);
assign 2_n6274 = ~2_n11439;
assign 2_n949 = 2_n638 | 2_n7227;
assign 2_n2724 = 2_n10955 | 2_n6744;
assign 2_n1838 = 2_n4683 & 2_n2732;
assign 2_n11205 = ~(2_n9123 | 2_n3969);
assign 2_n7628 = ~(2_n12520 ^ 2_n12664);
assign 2_n10019 = ~(2_n144 | 2_n7137);
assign 2_n8244 = ~2_n2398;
assign 2_n12298 = 2_n7116 | 2_n5538;
assign 2_n3235 = 2_n1297 & 2_n1391;
assign 2_n5873 = ~(2_n5553 ^ 2_n2765);
assign 2_n12679 = 2_n3076 | 2_n10868;
assign 2_n8149 = ~2_n874;
assign 2_n394 = ~(2_n8235 ^ 2_n10175);
assign 2_n11958 = ~2_n8336;
assign 2_n2562 = 2_n3015 | 2_n2294;
assign 2_n3133 = 2_n12093 & 2_n10939;
assign 2_n1969 = ~(2_n10874 ^ 2_n1300);
assign 2_n12672 = ~(2_n6270 ^ 2_n11978);
assign 2_n5264 = ~2_n12133;
assign 2_n11520 = ~2_n11983;
assign 2_n1272 = 2_n4562 | 2_n12689;
assign 2_n5241 = ~(2_n353 ^ 2_n10828);
assign 2_n775 = 2_n752 | 2_n12357;
assign 2_n5071 = 2_n3533 | 2_n5660;
assign 2_n8566 = ~(2_n6399 ^ 2_n1740);
assign 2_n1610 = ~(2_n12129 ^ 2_n5165);
assign 2_n11049 = 2_n10340 & 2_n1460;
assign 2_n3005 = ~(2_n11081 ^ 2_n3086);
assign 2_n6077 = 2_n7850 | 2_n3566;
assign 2_n6259 = ~(2_n4357 | 2_n3103);
assign 2_n8124 = 2_n12940 & 2_n4297;
assign 2_n4506 = 2_n8583 | 2_n2020;
assign 2_n2742 = 2_n5964 & 2_n6038;
assign 2_n7667 = ~(2_n4501 ^ 2_n6334);
assign 2_n7806 = 2_n10142 | 2_n130;
assign 2_n907 = 2_n4528 | 2_n6187;
assign 2_n3718 = 2_n989 | 2_n11746;
assign 2_n866 = 2_n2456 | 2_n10422;
assign 2_n6163 = 2_n9262 | 2_n9521;
assign 2_n3255 = 2_n2099 | 2_n8109;
assign 2_n4031 = ~(2_n7316 ^ 2_n9090);
assign 2_n6403 = ~(2_n10601 ^ 2_n1802);
assign 2_n10833 = 2_n5828 & 2_n5186;
assign 2_n5879 = ~(2_n1688 ^ 2_n8703);
assign 2_n5852 = ~(2_n6663 ^ 2_n8456);
assign 2_n2918 = ~(2_n672 ^ 2_n11454);
assign 2_n4185 = 2_n4582 & 2_n3955;
assign 2_n3633 = ~(2_n9139 ^ 2_n2200);
assign 2_n10186 = 2_n6293 | 2_n11194;
assign 2_n4922 = 2_n8831 ^ 2_n6406;
assign 2_n6365 = 2_n8959 | 2_n3903;
assign 2_n5015 = ~(2_n11027 ^ 2_n3611);
assign 2_n12085 = ~(2_n58 ^ 2_n6146);
assign 2_n8798 = 2_n1375 & 2_n3527;
assign 2_n10892 = 2_n6283 & 2_n3543;
assign 2_n8559 = 2_n6554 | 2_n5201;
assign 2_n9514 = 2_n8951 & 2_n11022;
assign 2_n10732 = ~2_n8960;
assign 2_n2169 = ~2_n5635;
assign 2_n6921 = 2_n1583 & 2_n7077;
assign 2_n4351 = 2_n4101 & 2_n9349;
assign 2_n10207 = ~2_n6326;
assign 2_n12256 = 2_n1078 | 2_n5983;
assign 2_n9852 = 2_n2696 & 2_n10412;
assign 2_n3637 = ~(2_n1044 ^ 2_n5602);
assign 2_n5022 = ~(2_n8826 | 2_n631);
assign 2_n9170 = ~2_n9920;
assign 2_n11241 = 2_n4038 & 2_n8589;
assign 2_n5436 = 2_n9000 | 2_n5391;
assign 2_n9979 = ~(2_n10218 ^ 2_n11393);
assign 2_n12520 = 2_n1185 & 2_n7755;
assign 2_n9065 = ~(2_n3452 ^ 2_n1370);
assign 2_n7031 = ~(2_n4195 ^ 2_n12121);
assign 2_n8309 = ~2_n12904;
assign 2_n2381 = ~(2_n6777 ^ 2_n2908);
assign 2_n4504 = 2_n4511 & 2_n8863;
assign 2_n7522 = ~(2_n3593 | 2_n12291);
assign 2_n8552 = ~2_n12648;
assign 2_n7340 = ~(2_n6337 ^ 2_n9447);
assign 2_n6425 = ~2_n12539;
assign 2_n11940 = 2_n5915 | 2_n8740;
assign 2_n5644 = ~(2_n1415 | 2_n4630);
assign 2_n8099 = 2_n10725 & 2_n5111;
assign 2_n2066 = ~2_n10959;
assign 2_n7617 = 2_n11744 | 2_n2222;
assign 2_n3293 = ~(2_n3625 ^ 2_n9031);
assign 2_n10781 = 2_n7405 | 2_n1148;
assign 2_n12956 = 2_n7427 & 2_n11868;
assign 2_n6884 = 2_n2515 & 2_n12925;
assign 2_n6050 = 2_n10157 | 2_n7506;
assign 2_n12348 = 2_n12119 | 2_n9188;
assign 2_n6523 = ~2_n5001;
assign 2_n7555 = ~2_n8083;
assign 2_n9005 = 2_n2213 & 2_n1443;
assign 2_n5284 = ~(2_n9973 ^ 2_n7180);
assign 2_n5695 = ~2_n4023;
assign 2_n9894 = ~(2_n6661 ^ 2_n4493);
assign 2_n7267 = 2_n4770 & 2_n560;
assign 2_n8822 = 2_n2456 | 2_n8109;
assign 2_n253 = 2_n10142 | 2_n1455;
assign 2_n9837 = 2_n8187 | 2_n1455;
assign 2_n7833 = ~(2_n10975 ^ 2_n2152);
assign 2_n4485 = ~(2_n3469 | 2_n12326);
assign 2_n2592 = 2_n10283 | 2_n4947;
assign 2_n3875 = 2_n11552 | 2_n2020;
assign 2_n4672 = ~(2_n12625 | 2_n9963);
assign 2_n2109 = ~(2_n1218 ^ 2_n4600);
assign 2_n5901 = 2_n8967 & 2_n1673;
assign 2_n2295 = 2_n10216 & 2_n2238;
assign 2_n2797 = 2_n4 | 2_n3283;
assign 2_n1523 = ~(2_n2262 ^ 2_n3564);
assign 2_n1050 = ~(2_n1706 ^ 2_n313);
assign 2_n10671 = 2_n2228 | 2_n5286;
assign 2_n12941 = ~2_n4619;
assign 2_n3401 = 2_n5767 & 2_n10848;
assign 2_n3000 = 2_n11732 & 2_n5506;
assign 2_n7854 = ~2_n2488;
assign 2_n6822 = ~(2_n7030 ^ 2_n10271);
assign 2_n5758 = 2_n11958 | 2_n5012;
assign 2_n2081 = 2_n5416 & 2_n7347;
assign 2_n3248 = 2_n11462 & 2_n11148;
assign 2_n9798 = 2_n3820 | 2_n4527;
assign 2_n5222 = ~(2_n7082 | 2_n10579);
assign 2_n5405 = ~(2_n9549 ^ 2_n4318);
assign 2_n8671 = 2_n5240 & 2_n3932;
assign 2_n8936 = ~(2_n2731 ^ 2_n5702);
assign 2_n5157 = 2_n4785 & 2_n6869;
assign 2_n8398 = ~(2_n7997 ^ 2_n3092);
assign 2_n4758 = ~2_n564;
assign 2_n12738 = 2_n9388 | 2_n10302;
assign 2_n11229 = 2_n12569 | 2_n9067;
assign 2_n610 = 2_n4983 & 2_n9636;
assign 2_n12953 = 2_n1747 & 2_n8610;
assign 2_n8315 = ~(2_n6961 ^ 2_n9019);
assign 2_n9202 = ~2_n9036;
assign 2_n12802 = ~(2_n9527 | 2_n8050);
assign 2_n8005 = 2_n10587 & 2_n10140;
assign 2_n12865 = ~(2_n236 ^ 2_n3770);
assign 2_n11003 = 2_n4415 & 2_n325;
assign 2_n9696 = ~(2_n5474 | 2_n11287);
assign 2_n6727 = ~(2_n2372 ^ 2_n1032);
assign 2_n12697 = ~(2_n288 ^ 2_n11386);
assign 2_n3292 = ~2_n9277;
assign 2_n8150 = ~(2_n5518 ^ 2_n9327);
assign 2_n7221 = ~(2_n904 ^ 2_n7464);
assign 2_n7572 = 2_n7449 | 2_n5759;
assign 2_n5818 = 2_n8907 | 2_n10483;
assign 2_n4960 = 2_n6353 & 2_n3601;
assign 2_n9346 = ~2_n5140;
assign 2_n4307 = 2_n7891 & 2_n521;
assign 2_n7064 = 2_n686 | 2_n7876;
assign 2_n8682 = 2_n2832 | 2_n4400;
assign 2_n4012 = 2_n8870 | 2_n3224;
assign 2_n3305 = 2_n12853 | 2_n8648;
assign 2_n8701 = 2_n5025 & 2_n56;
assign 2_n5869 = ~(2_n2525 ^ 2_n7174);
assign 2_n9160 = ~2_n10898;
assign 2_n477 = 2_n12797 | 2_n6455;
assign 2_n3710 = 2_n8738 | 2_n9521;
assign 2_n835 = 2_n5355 | 2_n4242;
assign 2_n8662 = ~(2_n9564 | 2_n706);
assign 2_n12815 = 2_n925 | 2_n1958;
assign 2_n9017 = 2_n4628 | 2_n8644;
assign 2_n1384 = ~2_n4349;
assign 2_n10836 = ~(2_n2048 | 2_n8939);
assign 2_n10408 = 2_n4222 & 2_n11724;
assign 2_n9774 = ~(2_n2820 ^ 2_n9672);
assign 2_n6411 = 2_n3251 | 2_n1274;
assign 2_n11125 = 2_n12635 | 2_n4988;
assign 2_n111 = 2_n10849 & 2_n6284;
assign 2_n1833 = 2_n5181 & 2_n3410;
assign 2_n5945 = ~2_n9241;
assign 2_n12455 = 2_n11923 | 2_n5258;
assign 2_n900 = ~(2_n7796 | 2_n4348);
assign 2_n3047 = ~(2_n4162 ^ 2_n10406);
assign 2_n11448 = ~(2_n2201 ^ 2_n12725);
assign 2_n6381 = 2_n636 | 2_n826;
assign 2_n8678 = ~2_n5955;
assign 2_n6269 = ~(2_n2055 ^ 2_n9941);
assign 2_n3977 = 2_n2921 | 2_n5604;
assign 2_n8521 = 2_n3797 & 2_n10816;
assign 2_n11664 = ~(2_n6835 ^ 2_n11469);
assign 2_n5201 = ~(2_n1671 ^ 2_n5862);
assign 2_n10662 = 2_n4628 | 2_n8109;
assign 2_n2773 = ~(2_n6211 | 2_n2576);
assign 2_n7407 = 2_n2099 | 2_n7382;
assign 2_n3935 = ~(2_n9967 ^ 2_n1893);
assign 2_n5524 = 2_n1937 | 2_n2815;
assign 2_n848 = 2_n4046 & 2_n12171;
assign 2_n3820 = ~2_n5198;
assign 2_n1498 = ~2_n993;
assign 2_n2192 = ~(2_n10555 | 2_n7791);
assign 2_n9892 = 2_n11552 | 2_n10916;
assign 2_n7537 = 2_n4015 & 2_n4740;
assign 2_n6407 = 2_n5575 | 2_n3903;
assign 2_n2450 = ~2_n6772;
assign 2_n6202 = ~(2_n4892 ^ 2_n4591);
assign 2_n6542 = 2_n5793 | 2_n798;
assign 2_n2756 = ~2_n2885;
assign 2_n814 = ~(2_n6496 | 2_n8190);
assign 2_n1888 = ~(2_n7082 ^ 2_n7845);
assign 2_n8442 = 2_n2300 & 2_n4130;
assign 2_n10048 = ~(2_n11569 ^ 2_n7880);
assign 2_n4366 = 2_n10750 | 2_n12735;
assign 2_n9675 = ~(2_n3934 ^ 2_n8888);
assign 2_n3566 = ~2_n3394;
assign 2_n1896 = 2_n4536 & 2_n4220;
assign 2_n8780 = ~(2_n4451 ^ 2_n1852);
assign 2_n5805 = ~(2_n5889 ^ 2_n7103);
assign 2_n6368 = 2_n1699 | 2_n7382;
assign 2_n6840 = ~(2_n7207 ^ 2_n12674);
assign 2_n12296 = 2_n11026 | 2_n9078;
assign 2_n6231 = 2_n752 | 2_n5538;
assign 2_n1699 = ~2_n5283;
assign 2_n9529 = 2_n3743 | 2_n8643;
assign 2_n5866 = 2_n1982 | 2_n7621;
assign 2_n202 = 2_n2382 & 2_n948;
assign 2_n3745 = ~(2_n6705 ^ 2_n5909);
assign 2_n3603 = ~2_n5544;
assign 2_n11988 = 2_n10879 | 2_n7881;
assign 2_n3331 = ~(2_n7462 ^ 2_n2105);
assign 2_n2817 = 2_n4498 | 2_n10066;
assign 2_n1089 = 2_n1024 | 2_n7498;
assign 2_n3836 = ~2_n2565;
assign 2_n4622 = 2_n12361 | 2_n5012;
assign 2_n7429 = ~(2_n5453 ^ 2_n5550);
assign 2_n9245 = 2_n2872 | 2_n7876;
assign 2_n1193 = ~(2_n515 ^ 2_n5941);
assign 2_n429 = ~(2_n6629 ^ 2_n8667);
assign 2_n2030 = 2_n7961 & 2_n10969;
assign 2_n10761 = 2_n10835 | 2_n5502;
assign 2_n11066 = ~(2_n8937 ^ 2_n534);
assign 2_n9733 = ~(2_n422 ^ 2_n12482);
assign 2_n11844 = ~(2_n2760 ^ 2_n1555);
assign 2_n4406 = ~(2_n12122 ^ 2_n11191);
assign 2_n5933 = ~(2_n4501 | 2_n8630);
assign 2_n1569 = 2_n10108 | 2_n1455;
assign 2_n12004 = ~(2_n5633 ^ 2_n9424);
assign 2_n7829 = ~2_n4409;
assign 2_n9063 = ~(2_n621 | 2_n6844);
assign 2_n3675 = ~2_n6251;
assign 2_n1836 = ~2_n10783;
assign 2_n1356 = ~(2_n12838 ^ 2_n3450);
assign 2_n10844 = ~(2_n7309 ^ 2_n9083);
assign 2_n5349 = ~(2_n90 | 2_n12732);
assign 2_n2232 = ~2_n11728;
assign 2_n1007 = 2_n989 | 2_n7246;
assign 2_n8573 = 2_n1944 & 2_n782;
assign 2_n1279 = 2_n4849 | 2_n1935;
assign 2_n300 = ~(2_n12487 | 2_n1857);
assign 2_n8732 = 2_n7449 | 2_n795;
assign 2_n11885 = ~(2_n8848 ^ 2_n5651);
assign 2_n53 = ~(2_n7227 ^ 2_n10494);
assign 2_n1023 = ~(2_n1034 ^ 2_n5722);
assign 2_n4578 = 2_n6241 & 2_n9948;
assign 2_n6461 = 2_n5765 | 2_n8643;
assign 2_n8997 = ~(2_n5415 | 2_n389);
assign 2_n5039 = 2_n10679 | 2_n6409;
assign 2_n7126 = 2_n5575 | 2_n5311;
assign 2_n1328 = ~(2_n5822 ^ 2_n2757);
assign 2_n12741 = ~2_n9246;
assign 2_n11901 = ~2_n6521;
assign 2_n10663 = ~2_n6889;
assign 2_n681 = 2_n2215 | 2_n6729;
assign 2_n7034 = ~(2_n12960 | 2_n10487);
assign 2_n6563 = 2_n127 & 2_n12679;
assign 2_n1570 = ~(2_n10720 ^ 2_n8088);
assign 2_n10690 = ~(2_n7032 | 2_n10895);
assign 2_n2956 = 2_n9607 | 2_n4429;
assign 2_n227 = ~(2_n8205 ^ 2_n6820);
assign 2_n1035 = ~(2_n5397 ^ 2_n6346);
assign 2_n3479 = 2_n4441 & 2_n4854;
assign 2_n12533 = ~(2_n12701 ^ 2_n5309);
assign 2_n470 = ~(2_n6975 ^ 2_n11853);
assign 2_n8088 = ~(2_n5643 ^ 2_n9173);
assign 2_n1556 = 2_n2367 | 2_n9521;
assign 2_n11616 = 2_n10983 | 2_n2817;
assign 2_n8421 = ~2_n2831;
assign 2_n474 = 2_n10835 | 2_n3451;
assign 2_n10444 = ~(2_n41 ^ 2_n383);
assign 2_n2156 = 2_n10518 | 2_n2916;
assign 2_n874 = ~(2_n2571 ^ 2_n11342);
assign 2_n7765 = ~2_n10096;
assign 2_n2010 = 2_n9943 | 2_n9035;
assign 2_n9771 = ~(2_n8612 ^ 2_n2335);
assign 2_n3407 = ~(2_n4619 | 2_n2719);
assign 2_n3918 = 2_n7937 | 2_n11145;
assign 2_n6804 = ~(2_n8003 | 2_n11638);
assign 2_n7648 = ~(2_n3645 ^ 2_n3493);
assign 2_n6926 = ~2_n508;
assign 2_n6571 = 2_n5915 | 2_n4913;
assign 2_n1352 = 2_n752 | 2_n2754;
assign 2_n10816 = ~2_n6467;
assign 2_n12193 = ~(2_n7045 ^ 2_n10937);
assign 2_n8492 = ~2_n12910;
assign 2_n3952 = 2_n4514 & 2_n9659;
assign 2_n7455 = ~(2_n1665 ^ 2_n5196);
assign 2_n522 = 2_n8738 | 2_n1047;
assign 2_n7087 = ~(2_n6801 | 2_n6011);
assign 2_n11079 = 2_n760 ^ 2_n12835;
assign 2_n1155 = 2_n6053 & 2_n5830;
assign 2_n1899 = 2_n9170 | 2_n3911;
assign 2_n7207 = ~(2_n7288 ^ 2_n4845);
assign 2_n9055 = 2_n7527 & 2_n9772;
assign 2_n10744 = 2_n5575 | 2_n11122;
assign 2_n11866 = ~2_n11022;
assign 2_n1903 = ~(2_n5544 | 2_n10443);
assign 2_n4298 = 2_n2832 | 2_n11827;
assign 2_n1982 = 2_n11984 & 2_n6460;
assign 2_n4167 = 2_n3127 | 2_n7881;
assign 2_n1086 = ~(2_n8776 | 2_n11526);
assign 2_n9447 = ~(2_n12270 ^ 2_n11676);
assign 2_n12139 = ~(2_n7549 ^ 2_n8096);
assign 2_n10906 = ~2_n9414;
assign 2_n3574 = 2_n7629 & 2_n2112;
assign 2_n2832 = ~2_n4516;
assign 2_n7381 = ~(2_n9028 | 2_n3945);
assign 2_n9860 = ~(2_n3276 | 2_n10787);
assign 2_n6025 = 2_n10818 & 2_n9949;
assign 2_n541 = 2_n4131 & 2_n10190;
assign 2_n4878 = 2_n683 & 2_n12834;
assign 2_n2883 = 2_n2834 & 2_n10526;
assign 2_n8855 = ~2_n11557;
assign 2_n46 = 2_n10776 & 2_n5683;
assign 2_n5837 = ~2_n6855;
assign 2_n9186 = 2_n12878 & 2_n10906;
assign 2_n1280 = ~2_n8241;
assign 2_n5114 = 2_n2168 & 2_n2354;
assign 2_n9281 = 2_n379 | 2_n5193;
assign 2_n1132 = ~(2_n2659 ^ 2_n6419);
assign 2_n6136 = 2_n124 & 2_n11883;
assign 2_n7899 = 2_n7449 | 2_n9144;
assign 2_n10597 = ~(2_n37 ^ 2_n11920);
assign 2_n7578 = 2_n11055 & 2_n12958;
assign 2_n6874 = ~(2_n10488 | 2_n6039);
assign 2_n12633 = 2_n7283 | 2_n11746;
assign 2_n2635 = ~(2_n1866 ^ 2_n10603);
assign 2_n6566 = 2_n12957 & 2_n71;
assign 2_n5107 = 2_n12237 | 2_n3924;
assign 2_n10603 = ~(2_n9271 ^ 2_n4185);
assign 2_n8154 = ~2_n1765;
assign 2_n9959 = ~2_n8455;
assign 2_n2216 = ~(2_n8288 | 2_n3999);
assign 2_n4410 = ~(2_n420 ^ 2_n10308);
assign 2_n11970 = ~2_n8122;
assign 2_n11969 = 2_n9887 | 2_n9226;
assign 2_n1656 = 2_n5902 | 2_n1455;
assign 2_n8345 = ~2_n1232;
assign 2_n3270 = ~(2_n5720 ^ 2_n6565);
assign 2_n8359 = 2_n7690 & 2_n12489;
assign 2_n4022 = 2_n5491 | 2_n7743;
assign 2_n5855 = 2_n1072 | 2_n2975;
assign 2_n7608 = 2_n3743 | 2_n1739;
assign 2_n9364 = ~2_n2345;
assign 2_n1649 = 2_n1231 | 2_n10446;
assign 2_n7316 = 2_n1051 | 2_n3903;
assign 2_n4358 = 2_n191 | 2_n8524;
assign 2_n7427 = 2_n2470 & 2_n1994;
assign 2_n9596 = ~(2_n2653 | 2_n12359);
assign 2_n12891 = ~(2_n7894 | 2_n1693);
assign 2_n3586 = ~(2_n8829 | 2_n8979);
assign 2_n7881 = ~2_n11877;
assign 2_n4268 = ~(2_n10929 ^ 2_n6328);
assign 2_n118 = 2_n8481 | 2_n1048;
assign 2_n2598 = ~2_n12644;
assign 2_n2170 = 2_n10846 | 2_n5525;
assign 2_n7942 = ~(2_n10405 ^ 2_n11004);
assign 2_n2877 = ~2_n11523;
assign 2_n8912 = 2_n994 | 2_n11827;
assign 2_n1640 = 2_n3196 & 2_n2274;
assign 2_n10097 = 2_n4929 & 2_n6833;
assign 2_n4056 = 2_n10051 & 2_n1836;
assign 2_n3946 = ~(2_n11069 | 2_n10056);
assign 2_n8999 = ~(2_n9604 | 2_n1743);
assign 2_n5874 = ~(2_n11265 ^ 2_n957);
assign 2_n7716 = 2_n7731 & 2_n3472;
assign 2_n11132 = 2_n4973 & 2_n12687;
assign 2_n3251 = 2_n8870 | 2_n1932;
assign 2_n2876 = 2_n4539 | 2_n893;
assign 2_n10541 = 2_n10157 | 2_n6138;
assign 2_n12057 = ~(2_n8404 ^ 2_n11739);
assign 2_n6437 = 2_n11341 | 2_n8484;
assign 2_n4294 = ~(2_n12788 | 2_n11907);
assign 2_n9517 = ~2_n1820;
assign 2_n2793 = 2_n10926 & 2_n11396;
assign 2_n10159 = 2_n10377 & 2_n6673;
assign 2_n11537 = ~(2_n9283 ^ 2_n9623);
assign 2_n128 = 2_n12119 | 2_n4818;
assign 2_n12288 = 2_n5915 | 2_n2964;
assign 2_n11235 = ~2_n2537;
assign 2_n1231 = 2_n3222 & 2_n12228;
assign 2_n4661 = ~2_n7720;
assign 2_n10702 = 2_n7965 & 2_n10990;
assign 2_n7827 = 2_n9389 | 2_n7703;
assign 2_n498 = ~(2_n6944 ^ 2_n3897);
assign 2_n5759 = ~2_n11296;
assign 2_n978 = ~(2_n8386 ^ 2_n5136);
assign 2_n9656 = 2_n10750 | 2_n12686;
assign 2_n12955 = 2_n12858 | 2_n8742;
assign 2_n5373 = 2_n3324 | 2_n9160;
assign 2_n4967 = 2_n2515 & 2_n5645;
assign 2_n9036 = 2_n6358 & 2_n2749;
assign 2_n9024 = ~(2_n2979 | 2_n4298);
assign 2_n6292 = 2_n2287 & 2_n12313;
assign 2_n2238 = ~(2_n6810 ^ 2_n635);
assign 2_n3703 = 2_n6836 & 2_n2004;
assign 2_n3878 = 2_n3072 | 2_n8111;
assign 2_n3744 = ~(2_n9240 ^ 2_n11671);
assign 2_n9623 = ~(2_n9884 ^ 2_n3411);
assign 2_n4852 = ~(2_n370 ^ 2_n2780);
assign 2_n4711 = ~(2_n7322 ^ 2_n256);
assign 2_n8604 = ~(2_n11526 ^ 2_n7175);
assign 2_n9339 = 2_n11887 | 2_n3924;
assign 2_n3856 = ~2_n1994;
assign 2_n9363 = ~(2_n4563 ^ 2_n8007);
assign 2_n12896 = ~(2_n2981 | 2_n6444);
assign 2_n71 = ~2_n1412;
assign 2_n4191 = ~(2_n7848 ^ 2_n10574);
assign 2_n3460 = ~(2_n9326 ^ 2_n4920);
assign 2_n4608 = 2_n1896 | 2_n1135;
assign 2_n3219 = 2_n6358 & 2_n7294;
assign 2_n24 = 2_n7283 | 2_n1079;
assign 2_n8815 = 2_n4613 & 2_n4098;
assign 2_n11820 = ~2_n3022;
assign 2_n970 = 2_n8295 | 2_n5242;
assign 2_n5919 = 2_n10417 & 2_n10146;
assign 2_n11685 = 2_n12468 & 2_n1749;
assign 2_n6440 = 2_n11038 & 2_n12451;
assign 2_n9043 = 2_n636 | 2_n12080;
assign 2_n2272 = 2_n11958 | 2_n11896;
assign 2_n6935 = ~(2_n7409 ^ 2_n10099);
assign 2_n11432 = ~(2_n4468 | 2_n7508);
assign 2_n10001 = 2_n1407 | 2_n4886;
assign 2_n3020 = 2_n137 & 2_n521;
assign 2_n7488 = ~(2_n6937 ^ 2_n12257);
assign 2_n6757 = ~(2_n12374 ^ 2_n7179);
assign 2_n7444 = ~(2_n9776 | 2_n11649);
assign 2_n12447 = 2_n1937 | 2_n5540;
assign 2_n9829 = 2_n5631 & 2_n5068;
assign 2_n12262 = 2_n8428 | 2_n10903;
assign 2_n4481 = ~2_n5732;
assign 2_n961 = 2_n953 & 2_n10528;
assign 2_n1504 = ~2_n8184;
assign 2_n9359 = ~(2_n7539 ^ 2_n2078);
assign 2_n11403 = ~2_n7168;
assign 2_n189 = 2_n1937 | 2_n8768;
assign 2_n7001 = 2_n1470 & 2_n1917;
assign 2_n3296 = 2_n4168 & 2_n4572;
assign 2_n7214 = 2_n6924 & 2_n12527;
assign 2_n11201 = 2_n1097 & 2_n3842;
assign 2_n10919 = ~2_n12221;
assign 2_n5268 = ~(2_n12781 ^ 2_n3843);
assign 2_n1460 = ~(2_n8341 ^ 2_n8747);
assign 2_n7665 = ~(2_n1462 ^ 2_n10617);
assign 2_n1312 = ~(2_n11589 ^ 2_n9892);
assign 2_n3635 = ~(2_n9346 ^ 2_n12926);
assign 2_n3897 = ~2_n8783;
assign 2_n468 = 2_n10097 | 2_n2415;
assign 2_n7641 = 2_n9982 | 2_n2386;
assign 2_n9398 = ~(2_n2449 ^ 2_n5721);
assign 2_n12105 = 2_n8164 & 2_n4762;
assign 2_n8394 = 2_n10196 | 2_n10916;
assign 2_n8085 = 2_n114 | 2_n2815;
assign 2_n5838 = 2_n10281 & 2_n9087;
assign 2_n3142 = ~2_n9089;
assign 2_n1883 = 2_n636 | 2_n1932;
assign 2_n10783 = 2_n989 | 2_n10066;
assign 2_n8115 = 2_n6391 & 2_n5824;
assign 2_n8106 = ~(2_n12794 ^ 2_n8113);
assign 2_n1310 = ~(2_n2203 ^ 2_n6915);
assign 2_n9749 = 2_n3127 | 2_n12328;
assign 2_n589 = 2_n10142 | 2_n1546;
assign 2_n9968 = ~(2_n5043 ^ 2_n2237);
assign 2_n12013 = ~2_n5742;
assign 2_n8915 = 2_n8026 | 2_n8414;
assign 2_n1188 = ~(2_n7528 ^ 2_n12216);
assign 2_n5729 = 2_n349 & 2_n3520;
assign 2_n2054 = ~(2_n6843 ^ 2_n12156);
assign 2_n5789 = 2_n2324 & 2_n3730;
assign 2_n11488 = ~2_n11577;
assign 2_n9085 = 2_n5172 | 2_n3111;
assign 2_n8369 = 2_n9370 | 2_n3911;
assign 2_n6638 = ~(2_n12098 ^ 2_n3561);
assign 2_n11590 = ~(2_n1157 ^ 2_n12418);
assign 2_n8967 = 2_n4213 | 2_n6233;
assign 2_n7093 = ~(2_n10060 ^ 2_n11229);
assign 2_n366 = ~(2_n7378 ^ 2_n2914);
assign 2_n9087 = 2_n3607 | 2_n4794;
assign 2_n3725 = 2_n6561 | 2_n8008;
assign 2_n11797 = ~(2_n9842 ^ 2_n7080);
assign 2_n2167 = 2_n10091 | 2_n100;
assign 2_n11207 = ~2_n6990;
assign 2_n6286 = ~2_n12516;
assign 2_n387 = ~(2_n12223 | 2_n7114);
assign 2_n2108 = 2_n7160 & 2_n7610;
assign 2_n1624 = 2_n5053 & 2_n12655;
assign 2_n3481 = ~(2_n2710 | 2_n4982);
assign 2_n9734 = 2_n6538 & 2_n10035;
assign 2_n11493 = ~2_n9342;
assign 2_n11549 = ~(2_n2036 ^ 2_n2853);
assign 2_n6207 = ~(2_n6426 ^ 2_n11009);
assign 2_n7297 = ~(2_n12857 ^ 2_n2212);
assign 2_n2731 = ~(2_n10544 ^ 2_n3315);
assign 2_n148 = 2_n10569 | 2_n3479;
assign 2_n8304 = 2_n8870 | 2_n12735;
assign 2_n4179 = ~2_n4799;
assign 2_n2080 = 2_n284 & 2_n10693;
assign 2_n12696 = 2_n7757 | 2_n858;
assign 2_n11123 = 2_n8959 | 2_n11410;
assign 2_n7620 = 2_n4498 | 2_n7881;
assign 2_n12330 = 2_n4206 | 2_n4303;
assign 2_n10932 = ~(2_n7415 ^ 2_n1499);
assign 2_n2895 = ~(2_n11373 ^ 2_n9883);
assign 2_n9922 = 2_n191 | 2_n9397;
assign 2_n5582 = 2_n11958 | 2_n11775;
assign 2_n3016 = 2_n10404 & 2_n8624;
assign 2_n9117 = ~(2_n6930 | 2_n8873);
assign 2_n4224 = 2_n4287 & 2_n12376;
assign 2_n10240 = ~(2_n1783 ^ 2_n906);
assign 2_n4895 = 2_n3688 & 2_n12045;
assign 2_n4559 = ~(2_n12309 | 2_n4593);
assign 2_n11204 = 2_n58 | 2_n12426;
assign 2_n11314 = ~(2_n11861 ^ 2_n4410);
assign 2_n5799 = ~(2_n10420 ^ 2_n1875);
assign 2_n8387 = 2_n191 | 2_n7341;
assign 2_n7741 = 2_n6996 & 2_n1137;
assign 2_n4969 = ~(2_n4508 ^ 2_n8495);
assign 2_n8663 = 2_n380 & 2_n12540;
assign 2_n7300 = 2_n8367 & 2_n388;
assign 2_n10203 = ~(2_n6137 | 2_n9404);
assign 2_n11349 = 2_n11433 | 2_n11820;
assign 2_n3521 = 2_n1824 & 2_n5011;
assign 2_n11305 = 2_n10835 | 2_n7506;
assign 2_n10460 = ~(2_n8002 ^ 2_n1494);
assign 2_n9891 = ~(2_n2799 ^ 2_n7711);
assign 2_n8581 = ~(2_n12296 ^ 2_n12877);
assign 2_n10148 = 2_n3820 | 2_n4875;
assign 2_n119 = ~(2_n5563 | 2_n5749);
assign 2_n2479 = 2_n1222 & 2_n9417;
assign 2_n3990 = ~(2_n2235 ^ 2_n5763);
assign 2_n11061 = 2_n5109 & 2_n12295;
assign 2_n6213 = 2_n9504 & 2_n11910;
assign 2_n3657 = ~(2_n12642 ^ 2_n1589);
assign 2_n3287 = ~(2_n6443 ^ 2_n8820);
assign 2_n1500 = 2_n3743 | 2_n2020;
assign 2_n9633 = 2_n6827 & 2_n10221;
assign 2_n7592 = ~(2_n7893 ^ 2_n6344);
assign 2_n7828 = ~(2_n11068 | 2_n7813);
assign 2_n3204 = ~(2_n6792 ^ 2_n6315);
assign 2_n10649 = ~2_n1088;
assign 2_n12871 = ~2_n223;
assign 2_n5536 = ~(2_n6165 ^ 2_n3663);
assign 2_n10853 = ~(2_n10819 ^ 2_n2776);
assign 2_n450 = ~(2_n1797 | 2_n8525);
assign 2_n10249 = ~(2_n5139 | 2_n5385);
assign 2_n5239 = ~2_n7428;
assign 2_n12637 = ~(2_n7042 ^ 2_n10717);
assign 2_n647 = ~(2_n12315 ^ 2_n1277);
assign 2_n6617 = ~2_n10163;
assign 2_n1128 = ~2_n4199;
assign 2_n11481 = ~2_n6688;
assign 2_n10867 = 2_n11867 & 2_n6075;
assign 2_n11271 = 2_n8114 | 2_n12902;
assign 2_n12020 = ~(2_n467 ^ 2_n10549);
assign 2_n5872 = ~(2_n7308 ^ 2_n12751);
assign 2_n6679 = ~(2_n3010 | 2_n3702);
assign 2_n1912 = ~(2_n4980 ^ 2_n6139);
assign 2_n3335 = 2_n6577 | 2_n5538;
assign 2_n4470 = ~(2_n4880 ^ 2_n7931);
assign 2_n1261 = ~2_n9592;
assign 2_n8358 = ~(2_n10740 ^ 2_n4444);
assign 2_n11548 = ~(2_n10615 | 2_n4699);
assign 2_n1022 = ~2_n10643;
assign 2_n2083 = 2_n3862 & 2_n57;
assign 2_n10173 = 2_n7078 | 2_n12905;
assign 2_n7804 = 2_n12878 | 2_n10906;
assign 2_n3519 = 2_n5125 & 2_n7598;
assign 2_n2234 = ~(2_n4278 | 2_n9769);
assign 2_n12119 = ~2_n4805;
assign 2_n3123 = 2_n10339 | 2_n8109;
assign 2_n9644 = ~2_n9482;
assign 2_n1070 = ~2_n2968;
assign 2_n11217 = ~(2_n4613 ^ 2_n10352);
assign 2_n6088 = 2_n11193 | 2_n5636;
assign 2_n2822 = 2_n6036 | 2_n707;
assign 2_n9664 = 2_n11849 | 2_n7971;
assign 2_n5957 = 2_n784 | 2_n4440;
assign 2_n8385 = ~(2_n9810 ^ 2_n7183);
assign 2_n5152 = 2_n1699 | 2_n5468;
assign 2_n12372 = 2_n852 ^ 2_n9711;
assign 2_n10 = ~2_n10987;
assign 2_n2537 = 2_n4828 & 2_n1512;
assign 2_n4343 = ~2_n4938;
assign 2_n4850 = 2_n12241 & 2_n9235;
assign 2_n8786 = 2_n12119 | 2_n12441;
assign 2_n10071 = ~(2_n10377 | 2_n6673);
assign 2_n7872 = 2_n6486 | 2_n1464;
assign 2_n2681 = 2_n5010 | 2_n2080;
assign 2_n3370 = ~2_n12106;
assign 2_n12301 = 2_n529 | 2_n8272;
assign 2_n3698 = 2_n5181 | 2_n3410;
assign 2_n2886 = ~(2_n2997 | 2_n6848);
assign 2_n4737 = ~(2_n547 | 2_n2487);
assign 2_n1762 = 2_n889 & 2_n6430;
assign 2_n953 = 2_n2564 & 2_n11662;
assign 2_n8982 = ~2_n3517;
assign 2_n3506 = 2_n386 | 2_n9354;
assign 2_n7102 = ~(2_n7769 ^ 2_n1970);
assign 2_n4269 = ~(2_n10139 ^ 2_n3615);
assign 2_n4838 = 2_n9010 & 2_n10988;
assign 2_n5236 = 2_n6877 & 2_n2024;
assign 2_n1820 = 2_n9372 & 2_n3358;
assign 2_n4814 = 2_n8512 | 2_n3286;
assign 2_n4508 = 2_n18 | 2_n9599;
assign 2_n737 = 2_n10196 | 2_n3606;
assign 2_n3807 = 2_n2217 | 2_n4474;
assign 2_n6133 = 2_n10750 | 2_n7136;
assign 2_n1297 = ~2_n12280;
assign 2_n927 = ~(2_n6673 ^ 2_n12863);
assign 2_n12821 = ~2_n8487;
assign 2_n5458 = 2_n252 | 2_n3957;
assign 2_n2020 = ~2_n10990;
assign 2_n403 = ~2_n7748;
assign 2_n3138 = ~(2_n8548 | 2_n6380);
assign 2_n10996 = ~2_n9263;
assign 2_n8450 = 2_n890 & 2_n2327;
assign 2_n2160 = ~(2_n9699 | 2_n4684);
assign 2_n9655 = ~(2_n5207 ^ 2_n7367);
assign 2_n1834 = ~2_n5614;
assign 2_n12604 = 2_n3743 | 2_n3599;
assign 2_n11450 = 2_n8870 | 2_n7928;
assign 2_n7737 = ~(2_n9922 ^ 2_n7669);
assign 2_n4790 = 2_n4778 | 2_n1932;
assign 2_n6652 = 2_n11433 | 2_n11775;
assign 2_n4575 = ~(2_n12949 | 2_n8289);
assign 2_n12579 = ~2_n9711;
assign 2_n10955 = 2_n7116 | 2_n6169;
assign 2_n10060 = ~(2_n12663 | 2_n593);
assign 2_n7469 = 2_n3127 | 2_n2358;
assign 2_n2903 = ~(2_n8542 ^ 2_n8434);
assign 2_n12562 = ~(2_n8862 ^ 2_n6630);
assign 2_n12722 = 2_n1177 & 2_n5354;
assign 2_n4325 = ~(2_n1596 ^ 2_n2450);
assign 2_n10112 = 2_n12303 & 2_n1394;
assign 2_n12517 = ~(2_n10552 ^ 2_n11925);
assign 2_n7419 = ~(2_n4511 ^ 2_n2623);
assign 2_n11022 = 2_n684 & 2_n11483;
assign 2_n11181 = 2_n9373 | 2_n3606;
assign 2_n2334 = ~2_n2851;
assign 2_n3071 = 2_n12746 ^ 2_n742;
assign 2_n944 = ~(2_n1708 ^ 2_n8882);
assign 2_n10937 = 2_n1323 | 2_n11688;
assign 2_n3651 = 2_n147 & 2_n12571;
assign 2_n3687 = 2_n9917 | 2_n9958;
assign 2_n10931 = 2_n1449 & 2_n1174;
assign 2_n9059 = 2_n6672 & 2_n1529;
assign 2_n12033 = 2_n989 | 2_n4242;
assign 2_n6789 = 2_n8613 | 2_n5943;
assign 2_n6992 = ~(2_n10697 ^ 2_n3995);
assign 2_n7371 = ~2_n8734;
assign 2_n11044 = 2_n989 | 2_n12843;
assign 2_n5903 = ~(2_n8605 | 2_n2161);
assign 2_n11618 = 2_n7485 & 2_n6576;
assign 2_n611 = ~(2_n11109 | 2_n80);
assign 2_n9919 = ~(2_n12448 ^ 2_n4930);
assign 2_n9108 = 2_n994 | 2_n1915;
assign 2_n4863 = 2_n3127 | 2_n6402;
assign 2_n9415 = ~(2_n8361 ^ 2_n9641);
assign 2_n4543 = ~(2_n8147 ^ 2_n5270);
assign 2_n5677 = 2_n7526 | 2_n790;
assign 2_n6082 = ~(2_n4738 | 2_n2794);
assign 2_n2106 = 2_n8600 & 2_n2445;
assign 2_n3830 = 2_n4995 & 2_n1652;
assign 2_n7296 = ~(2_n5967 ^ 2_n7486);
assign 2_n9242 = ~(2_n301 ^ 2_n10285);
assign 2_n11121 = 2_n10822 | 2_n4711;
assign 2_n8176 = 2_n5434 & 2_n11354;
assign 2_n4382 = 2_n1867 | 2_n7371;
assign 2_n4262 = ~2_n2387;
assign 2_n2258 = 2_n365 | 2_n5457;
assign 2_n11810 = 2_n6313 & 2_n4816;
assign 2_n11767 = 2_n7299 | 2_n2239;
assign 2_n6984 = ~(2_n4147 | 2_n9011);
assign 2_n6306 = ~2_n2116;
assign 2_n10293 = 2_n7978 & 2_n9566;
assign 2_n6771 = ~(2_n10526 ^ 2_n3458);
assign 2_n5769 = 2_n10835 | 2_n4864;
assign 2_n5025 = ~2_n6070;
assign 2_n11025 = ~(2_n7098 ^ 2_n2391);
assign 2_n2813 = ~2_n7244;
assign 2_n9800 = 2_n12417 | 2_n11590;
assign 2_n1673 = 2_n986 | 2_n11426;
assign 2_n6300 = ~(2_n6408 ^ 2_n528);
assign 2_n2539 = 2_n2099 | 2_n12754;
assign 2_n6486 = 2_n7449 | 2_n10916;
assign 2_n9172 = ~2_n11672;
assign 2_n7226 = 2_n11384 & 2_n668;
assign 2_n12271 = 2_n5355 | 2_n2076;
assign 2_n1588 = ~(2_n7600 ^ 2_n8463);
assign 2_n9467 = ~(2_n8593 ^ 2_n6511);
assign 2_n5569 = 2_n8870 | 2_n530;
assign 2_n11736 = ~2_n2402;
assign 2_n693 = 2_n897 | 2_n4850;
assign 2_n9488 = ~(2_n2563 | 2_n2196);
assign 2_n4054 = 2_n9500 | 2_n9964;
assign 2_n10580 = ~(2_n10221 ^ 2_n5461);
assign 2_n10398 = 2_n6078 | 2_n2672;
assign 2_n4854 = 2_n4979 | 2_n8884;
assign 2_n2153 = ~(2_n6731 ^ 2_n2283);
assign 2_n8726 = ~(2_n12248 ^ 2_n1573);
assign 2_n11426 = 2_n4213 & 2_n6233;
assign 2_n12131 = 2_n95 & 2_n6792;
assign 2_n3363 = ~(2_n981 | 2_n3296);
assign 2_n9630 = ~(2_n6560 ^ 2_n3741);
assign 2_n875 = 2_n7874 & 2_n12918;
assign 2_n1463 = 2_n5183 & 2_n6299;
assign 2_n2195 = 2_n9648 | 2_n5802;
assign 2_n485 = ~(2_n12670 | 2_n8341);
assign 2_n3373 = ~(2_n7919 | 2_n5872);
assign 2_n10500 = 2_n11580 & 2_n3823;
assign 2_n2329 = 2_n2456 | 2_n12124;
assign 2_n9276 = ~2_n662;
assign 2_n7686 = 2_n9389 | 2_n7881;
assign 2_n303 = 2_n1404 | 2_n10558;
assign 2_n5698 = 2_n10771 | 2_n11045;
assign 2_n8170 = ~(2_n2161 ^ 2_n8605);
assign 2_n3416 = ~(2_n10288 ^ 2_n7900);
assign 2_n8719 = ~(2_n1152 ^ 2_n10123);
assign 2_n10618 = ~(2_n12319 ^ 2_n2030);
assign 2_n5808 = 2_n686 | 2_n2815;
assign 2_n3812 = ~(2_n9026 ^ 2_n4683);
assign 2_n6835 = ~(2_n9229 ^ 2_n6762);
assign 2_n5408 = 2_n3743 | 2_n9521;
assign 2_n5608 = 2_n2167 & 2_n8413;
assign 2_n4137 = ~(2_n5254 ^ 2_n8264);
assign 2_n5887 = 2_n8583 | 2_n4527;
assign 2_n11927 = 2_n10915 & 2_n6020;
assign 2_n11194 = 2_n2976 & 2_n11495;
assign 2_n12498 = ~(2_n11450 ^ 2_n10908);
assign 2_n1105 = 2_n5134 & 2_n5477;
assign 2_n5566 = ~(2_n3964 ^ 2_n2981);
assign 2_n10819 = ~(2_n2119 ^ 2_n2264);
assign 2_n795 = ~2_n8028;
assign 2_n5802 = 2_n8959 | 2_n11775;
assign 2_n2859 = ~(2_n9204 ^ 2_n8693);
assign 2_n762 = 2_n2456 | 2_n1932;
assign 2_n7188 = 2_n3096 | 2_n6455;
assign 2_n6203 = 2_n4059 | 2_n4242;
assign 2_n8285 = ~2_n6441;
assign 2_n3727 = ~(2_n2029 ^ 2_n8500);
assign 2_n1544 = ~(2_n10128 ^ 2_n2451);
assign 2_n1909 = 2_n9656 | 2_n12411;
assign 2_n12880 = 2_n9812 | 2_n10836;
assign 2_n10740 = 2_n4662 | 2_n8987;
assign 2_n304 = ~2_n4484;
assign 2_n4317 = 2_n4547 & 2_n7335;
assign 2_n8390 = ~(2_n7200 ^ 2_n7499);
assign 2_n8526 = 2_n4772 & 2_n9470;
assign 2_n8908 = 2_n12361 | 2_n10919;
assign 2_n6624 = ~(2_n7365 ^ 2_n1753);
assign 2_n1861 = ~2_n4439;
assign 2_n10624 = 2_n12344 & 2_n815;
assign 2_n9682 = 2_n2367 | 2_n795;
assign 2_n7688 = 2_n4628 | 2_n12686;
assign 2_n8859 = ~2_n1835;
assign 2_n10216 = 2_n8159 | 2_n5299;
assign 2_n82 = ~(2_n12348 ^ 2_n9399);
assign 2_n746 = ~(2_n3437 ^ 2_n12075);
assign 2_n2775 = ~(2_n12052 ^ 2_n6440);
assign 2_n7308 = ~(2_n1631 ^ 2_n7296);
assign 2_n9531 = 2_n10157 | 2_n4654;
assign 2_n4147 = ~(2_n9369 | 2_n2952);
assign 2_n11588 = ~(2_n11262 ^ 2_n9056);
assign 2_n7244 = 2_n11552 | 2_n4654;
assign 2_n8120 = 2_n5504 | 2_n9925;
assign 2_n3186 = 2_n3930 & 2_n4483;
assign 2_n12024 = 2_n9827 & 2_n11599;
assign 2_n657 = ~(2_n7662 ^ 2_n1800);
assign 2_n9856 = ~2_n1050;
assign 2_n5854 = ~(2_n6472 | 2_n2174);
assign 2_n2629 = 2_n5945 | 2_n6455;
assign 2_n3384 = ~(2_n7520 ^ 2_n9133);
assign 2_n8391 = ~(2_n1151 ^ 2_n6998);
assign 2_n5662 = 2_n9498 | 2_n3880;
assign 2_n2449 = ~(2_n9155 ^ 2_n3395);
assign 2_n6591 = ~(2_n7790 ^ 2_n6416);
assign 2_n2251 = 2_n6667 | 2_n604;
assign 2_n3839 = ~(2_n12443 ^ 2_n1734);
assign 2_n4896 = ~2_n4850;
assign 2_n4211 = ~(2_n7916 | 2_n2642);
assign 2_n12199 = ~2_n1456;
assign 2_n4036 = ~(2_n4588 | 2_n7660);
assign 2_n9136 = ~(2_n1228 ^ 2_n7560);
assign 2_n10338 = 2_n2217 | 2_n8643;
assign 2_n3997 = 2_n5809 | 2_n4818;
assign 2_n9722 = ~(2_n8617 ^ 2_n2375);
assign 2_n2159 = 2_n6924 | 2_n12527;
assign 2_n1052 = 2_n7024 | 2_n4661;
assign 2_n2994 = ~2_n3734;
assign 2_n1696 = 2_n8583 | 2_n4474;
assign 2_n5509 = ~(2_n1624 ^ 2_n6194);
assign 2_n1954 = ~(2_n5825 ^ 2_n12620);
assign 2_n4085 = ~2_n8760;
assign 2_n9061 = 2_n11714 | 2_n5551;
assign 2_n9772 = ~2_n5344;
assign 2_n11704 = 2_n191 | 2_n130;
assign 2_n11193 = ~2_n7416;
assign 2_n5285 = 2_n8416 | 2_n2933;
assign 2_n8790 = 2_n752 | 2_n2232;
assign 2_n1790 = ~2_n8204;
assign 2_n9072 = ~(2_n12287 ^ 2_n241);
assign 2_n10779 = ~(2_n10038 ^ 2_n9451);
assign 2_n6627 = ~2_n8094;
assign 2_n9150 = 2_n6577 | 2_n12816;
assign 2_n7683 = ~2_n11243;
assign 2_n8045 = 2_n5575 | 2_n12357;
assign 2_n3761 = 2_n3127 | 2_n12843;
assign 2_n2149 = 2_n4679 & 2_n1668;
assign 2_n4486 = ~(2_n12611 ^ 2_n10753);
assign 2_n10479 = ~2_n10402;
assign 2_n11931 = 2_n9171 | 2_n9221;
assign 2_n2365 = ~(2_n4991 ^ 2_n7427);
assign 2_n9810 = ~(2_n8275 ^ 2_n9052);
assign 2_n12552 = ~(2_n5948 ^ 2_n233);
assign 2_n7979 = 2_n11255 & 2_n2591;
assign 2_n5742 = ~(2_n4465 ^ 2_n475);
assign 2_n8350 = ~(2_n5486 ^ 2_n3662);
assign 2_n11878 = 2_n10611 | 2_n7249;
assign 2_n4546 = 2_n7116 | 2_n5012;
assign 2_n1301 = ~(2_n262 ^ 2_n5634);
assign 2_n4057 = 2_n5233 & 2_n11201;
assign 2_n11687 = 2_n989 | 2_n8524;
assign 2_n12041 = 2_n6042 | 2_n576;
assign 2_n635 = 2_n3018 ^ 2_n11831;
assign 2_n7158 = 2_n3976 & 2_n12059;
assign 2_n3195 = ~(2_n4908 | 2_n6596);
assign 2_n7605 = ~(2_n6153 ^ 2_n9374);
assign 2_n7273 = ~2_n3020;
assign 2_n12398 = 2_n7420 | 2_n12475;
assign 2_n1492 = ~(2_n12324 ^ 2_n2736);
assign 2_n12911 = ~(2_n4148 ^ 2_n8399);
assign 2_n2871 = 2_n9634 & 2_n1250;
assign 2_n1641 = ~2_n633;
assign 2_n8332 = 2_n7052 | 2_n1864;
assign 2_n8363 = ~2_n9757;
assign 2_n7253 = 2_n1951 ^ 2_n3432;
assign 2_n2270 = 2_n6516 | 2_n4321;
assign 2_n360 = ~(2_n178 ^ 2_n5387);
assign 2_n4624 = ~2_n1826;
assign 2_n1706 = 2_n2217 | 2_n28;
assign 2_n2384 = ~2_n6661;
assign 2_n11991 = ~(2_n4595 | 2_n5624);
assign 2_n6058 = 2_n6977 | 2_n3468;
assign 2_n3029 = 2_n8354 | 2_n4913;
assign 2_n36 = 2_n4387 & 2_n4162;
assign 2_n5600 = 2_n7391 | 2_n11746;
assign 2_n8036 = ~(2_n4906 | 2_n9830);
assign 2_n4527 = ~2_n11876;
assign 2_n7877 = ~(2_n4283 ^ 2_n10925);
assign 2_n2274 = 2_n6017 | 2_n7056;
assign 2_n9567 = ~(2_n9203 ^ 2_n66);
assign 2_n5693 = ~(2_n6640 ^ 2_n9463);
assign 2_n6783 = 2_n10749 | 2_n7229;
assign 2_n4327 = ~2_n6129;
assign 2_n6745 = 2_n6369 & 2_n3522;
assign 2_n3365 = ~(2_n8194 | 2_n4035);
assign 2_n207 = ~(2_n1811 ^ 2_n829);
assign 2_n9123 = 2_n294 & 2_n7023;
assign 2_n11209 = ~(2_n1809 ^ 2_n8290);
assign 2_n593 = ~(2_n3441 | 2_n2121);
assign 2_n12921 = ~(2_n7189 ^ 2_n3107);
assign 2_n8901 = 2_n1472 | 2_n5;
assign 2_n1322 = 2_n5425 & 2_n2245;
assign 2_n10956 = 2_n525 | 2_n8058;
assign 2_n12500 = ~(2_n9014 | 2_n10933);
assign 2_n7972 = ~(2_n9708 | 2_n3779);
assign 2_n9933 = 2_n8267 | 2_n11939;
assign 2_n5388 = ~2_n2166;
assign 2_n7089 = 2_n5919 | 2_n9242;
assign 2_n8189 = 2_n994 | 2_n7424;
assign 2_n1027 = ~(2_n9307 ^ 2_n1948);
assign 2_n5041 = ~(2_n6704 ^ 2_n6428);
assign 2_n2032 = ~(2_n8647 ^ 2_n8408);
assign 2_n8376 = 2_n5205 & 2_n1662;
assign 2_n8715 = ~(2_n9469 ^ 2_n10314);
assign 2_n8300 = ~(2_n5323 ^ 2_n9025);
assign 2_n8914 = ~(2_n10483 ^ 2_n7852);
assign 2_n1275 = 2_n7495 | 2_n11827;
assign 2_n4705 = ~(2_n5279 ^ 2_n2147);
assign 2_n9710 = ~2_n12089;
assign 2_n751 = ~(2_n4301 ^ 2_n11741);
assign 2_n11813 = 2_n5614 & 2_n12895;
assign 2_n7462 = 2_n2099 | 2_n12735;
assign 2_n7251 = 2_n8026 | 2_n995;
assign 2_n7084 = 2_n752 | 2_n11896;
assign 2_n6067 = 2_n7233 & 2_n10059;
assign 2_n3615 = 2_n1514 & 2_n1149;
assign 2_n7919 = 2_n2002 & 2_n12342;
assign 2_n2836 = ~(2_n196 ^ 2_n11477);
assign 2_n1923 = ~2_n7342;
assign 2_n7256 = 2_n9110 | 2_n10628;
assign 2_n5381 = ~(2_n2142 ^ 2_n6216);
assign 2_n518 = ~2_n2630;
assign 2_n6009 = ~(2_n885 | 2_n5836);
assign 2_n8692 = 2_n5765 | 2_n8830;
assign 2_n7071 = 2_n10142 | 2_n6402;
assign 2_n2986 = 2_n2982 & 2_n4319;
assign 2_n1260 = 2_n7495 | 2_n7341;
assign 2_n8865 = 2_n8295 & 2_n5242;
assign 2_n8706 = ~(2_n9450 ^ 2_n11002);
assign 2_n11533 = 2_n10750 | 2_n9586;
assign 2_n8978 = 2_n11026 | 2_n12771;
assign 2_n6251 = 2_n2171 | 2_n10445;
assign 2_n7661 = 2_n1598 | 2_n5564;
assign 2_n2112 = 2_n12116 | 2_n6938;
assign 2_n7255 = ~(2_n9595 ^ 2_n162);
assign 2_n6427 = ~(2_n9785 ^ 2_n7764);
assign 2_n1479 = ~(2_n2542 ^ 2_n12206);
assign 2_n4883 = 2_n7388 & 2_n11876;
assign 2_n1748 = 2_n639 & 2_n1669;
assign 2_n7868 = ~(2_n5508 ^ 2_n3349);
assign 2_n11971 = 2_n3032 & 2_n281;
assign 2_n5323 = 2_n1764 | 2_n3495;
assign 2_n3157 = 2_n1705 & 2_n12251;
assign 2_n11446 = 2_n11416 & 2_n2535;
assign 2_n2189 = ~2_n2181;
assign 2_n8286 = 2_n8583 | 2_n4654;
assign 2_n9988 = ~(2_n3706 | 2_n10461);
assign 2_n4193 = ~2_n2858;
assign 2_n1710 = 2_n505 & 2_n12592;
assign 2_n883 = ~(2_n12210 | 2_n601);
assign 2_n11160 = ~(2_n1988 ^ 2_n4194);
assign 2_n1040 = ~(2_n6782 ^ 2_n1503);
assign 2_n1003 = ~(2_n8347 ^ 2_n8488);
assign 2_n5203 = 2_n10697 | 2_n4968;
assign 2_n3488 = ~2_n11467;
assign 2_n7905 = 2_n5663 & 2_n11387;
assign 2_n9883 = 2_n2466 & 2_n10806;
assign 2_n3451 = ~2_n1357;
assign 2_n10371 = ~(2_n10563 ^ 2_n7222);
assign 2_n12349 = ~2_n11040;
assign 2_n5622 = 2_n11478 & 2_n12925;
assign 2_n9076 = 2_n12227 | 2_n11940;
assign 2_n8305 = ~2_n8044;
assign 2_n11731 = ~2_n1750;
assign 2_n8866 = 2_n282 | 2_n7494;
assign 2_n10713 = ~(2_n10381 ^ 2_n2837);
assign 2_n1106 = 2_n12552 & 2_n6989;
assign 2_n8778 = 2_n8583 | 2_n9568;
assign 2_n6847 = ~2_n9450;
assign 2_n4573 = ~2_n6998;
assign 2_n2299 = ~(2_n1223 ^ 2_n9500);
assign 2_n12028 = ~2_n8420;
assign 2_n2242 = ~2_n12915;
assign 2_n10201 = ~(2_n9476 | 2_n10602);
assign 2_n9201 = ~(2_n1321 ^ 2_n10886);
assign 2_n7524 = ~(2_n1921 ^ 2_n12402);
assign 2_n10038 = 2_n191 | 2_n6524;
assign 2_n2747 = ~(2_n10318 | 2_n10110);
assign 2_n5286 = ~(2_n7616 ^ 2_n1723);
assign 2_n10025 = 2_n8310 & 2_n2912;
assign 2_n8456 = 2_n5858 | 2_n3911;
assign 2_n184 = ~2_n11423;
assign 2_n9438 = ~(2_n2305 ^ 2_n10643);
assign 2_n9557 = ~(2_n4174 ^ 2_n4470);
assign 2_n8063 = 2_n1699 | 2_n8259;
assign 2_n8772 = 2_n10928 & 2_n7946;
assign 2_n933 = ~(2_n11413 ^ 2_n5653);
assign 2_n3805 = ~(2_n11637 ^ 2_n11738);
assign 2_n12671 = ~(2_n7311 ^ 2_n10151);
assign 2_n1332 = ~(2_n2842 ^ 2_n6260);
assign 2_n12007 = ~(2_n4154 | 2_n5746);
assign 2_n11495 = 2_n989 | 2_n6389;
assign 2_n7995 = 2_n6943 & 2_n7182;
assign 2_n3608 = 2_n8622 & 2_n6200;
assign 2_n4050 = ~2_n1021;
assign 2_n554 = 2_n10774 & 2_n6765;
assign 2_n9353 = 2_n10750 | 2_n3224;
assign 2_n7246 = ~2_n4005;
assign 2_n7496 = ~(2_n551 ^ 2_n7975);
assign 2_n9735 = 2_n4628 | 2_n6071;
assign 2_n9487 = ~(2_n12619 ^ 2_n10166);
assign 2_n4603 = ~(2_n2878 ^ 2_n10786);
assign 2_n3864 = ~2_n4678;
assign 2_n5711 = 2_n6740 & 2_n9524;
assign 2_n9784 = ~(2_n7331 ^ 2_n1865);
assign 2_n7149 = ~2_n6954;
assign 2_n5574 = ~2_n7520;
assign 2_n3784 = ~(2_n3659 | 2_n4993);
assign 2_n11307 = 2_n1882 | 2_n2043;
assign 2_n1887 = 2_n4647 | 2_n11236;
assign 2_n11811 = ~2_n7289;
assign 2_n10495 = ~(2_n255 ^ 2_n6879);
assign 2_n3494 = 2_n7662 | 2_n1800;
assign 2_n9827 = 2_n10780 & 2_n12942;
assign 2_n7914 = 2_n11958 | 2_n7558;
assign 2_n2514 = ~(2_n11664 ^ 2_n8314);
assign 2_n966 = 2_n994 | 2_n12843;
assign 2_n5282 = 2_n11433 | 2_n2815;
assign 2_n11332 = ~(2_n8376 | 2_n1378);
assign 2_n5076 = 2_n11451 & 2_n6466;
assign 2_n824 = ~2_n6322;
assign 2_n8472 = ~(2_n6730 ^ 2_n7510);
assign 2_n4435 = ~(2_n9263 ^ 2_n8292);
assign 2_n865 = ~(2_n10191 ^ 2_n9654);
assign 2_n8983 = 2_n12871 & 2_n5649;
assign 2_n7384 = 2_n7462 & 2_n2105;
assign 2_n5360 = 2_n10381 & 2_n6177;
assign 2_n11696 = ~2_n10857;
assign 2_n1960 = 2_n989 | 2_n1851;
assign 2_n5568 = ~(2_n7020 ^ 2_n5668);
assign 2_n9341 = 2_n3127 | 2_n1915;
assign 2_n5942 = ~(2_n11488 ^ 2_n192);
assign 2_n891 = 2_n3820 | 2_n4474;
assign 2_n2430 = 2_n12361 | 2_n5540;
assign 2_n10798 = 2_n11552 | 2_n9521;
assign 2_n2363 = 2_n191 | 2_n12328;
assign 2_n11867 = 2_n9389 | 2_n7341;
assign 2_n2328 = ~(2_n8592 | 2_n5609);
assign 2_n1915 = ~2_n7456;
assign 2_n1249 = 2_n191 | 2_n4242;
assign 2_n7602 = ~(2_n8333 ^ 2_n5446);
assign 2_n3011 = 2_n4805 & 2_n1067;
assign 2_n6708 = ~(2_n5035 ^ 2_n4003);
assign 2_n5922 = 2_n11958 | 2_n12274;
assign 2_n8258 = 2_n11534 & 2_n483;
assign 2_n9013 = 2_n10389 | 2_n9041;
assign 2_n840 = ~(2_n11086 ^ 2_n5120);
assign 2_n4320 = ~2_n12733;
assign 2_n8713 = ~(2_n9849 | 2_n8268);
assign 2_n9372 = 2_n2312 | 2_n3899;
assign 2_n9232 = 2_n12715 | 2_n7065;
assign 2_n5907 = ~(2_n4491 ^ 2_n235);
assign 2_n5083 = ~(2_n7899 ^ 2_n10565);
assign 2_n2637 = ~2_n11758;
assign 2_n8899 = ~(2_n5894 ^ 2_n9436);
assign 2_n2359 = 2_n12503 | 2_n9160;
assign 2_n11170 = 2_n3464 & 2_n8805;
assign 2_n3456 = ~(2_n8160 ^ 2_n7692);
assign 2_n9742 = 2_n6758 | 2_n3387;
assign 2_n7983 = 2_n2456 | 2_n9586;
assign 2_n10519 = ~(2_n5888 ^ 2_n12923);
assign 2_n4127 = 2_n10960 | 2_n10315;
assign 2_n2969 = ~2_n2;
assign 2_n2230 = 2_n994 | 2_n561;
assign 2_n4277 = 2_n5510 | 2_n6609;
assign 2_n10611 = ~2_n5606;
assign 2_n2915 = 2_n4674 | 2_n12535;
assign 2_n10357 = ~(2_n6012 ^ 2_n5440);
assign 2_n3095 = ~2_n11594;
assign 2_n12876 = ~(2_n6009 | 2_n1613);
assign 2_n8195 = 2_n11887 | 2_n8109;
assign 2_n912 = ~(2_n10768 ^ 2_n328);
assign 2_n1033 = ~(2_n8146 ^ 2_n5613);
assign 2_n1753 = ~(2_n4576 ^ 2_n8052);
assign 2_n6162 = 2_n3724 | 2_n53;
assign 2_n7994 = 2_n11850 & 2_n5458;
assign 2_n9835 = ~2_n250;
assign 2_n8081 = ~(2_n622 ^ 2_n7987);
assign 2_n774 = ~(2_n6316 ^ 2_n210);
assign 2_n2176 = ~(2_n2635 ^ 2_n1232);
assign 2_n9946 = 2_n1699 | 2_n8644;
assign 2_n8774 = ~2_n6867;
assign 2_n7026 = ~(2_n10052 | 2_n7353);
assign 2_n9303 = 2_n6373 | 2_n4864;
assign 2_n1234 = ~(2_n5067 | 2_n12236);
assign 2_n11304 = ~2_n12573;
assign 2_n11203 = 2_n994 | 2_n4775;
assign 2_n7151 = ~(2_n8634 ^ 2_n11370);
assign 2_n2891 = ~(2_n5873 ^ 2_n8867);
assign 2_n2034 = ~2_n7983;
assign 2_n6862 = ~(2_n7845 | 2_n5222);
assign 2_n7184 = 2_n12244 | 2_n9425;
assign 2_n4081 = ~(2_n6919 | 2_n4935);
assign 2_n3496 = ~(2_n3585 | 2_n6383);
assign 2_n5491 = 2_n7116 | 2_n995;
assign 2_n9441 = 2_n8920 | 2_n8547;
assign 2_n857 = 2_n6331 | 2_n9550;
assign 2_n2135 = ~2_n531;
assign 2_n3241 = ~(2_n4806 | 2_n10449);
assign 2_n4740 = 2_n10798 | 2_n10133;
assign 2_n12924 = ~2_n12266;
assign 2_n4230 = ~(2_n5447 ^ 2_n4621);
assign 2_n11421 = ~2_n1810;
assign 2_n2927 = ~2_n10834;
assign 2_n9578 = ~(2_n1669 ^ 2_n5142);
assign 2_n10345 = ~(2_n12204 ^ 2_n1858);
assign 2_n10301 = ~2_n2321;
assign 2_n35 = ~(2_n5570 ^ 2_n8963);
assign 2_n3408 = 2_n8601 | 2_n2737;
assign 2_n3514 = ~(2_n2190 ^ 2_n2663);
assign 2_n9491 = ~(2_n12377 ^ 2_n8881);
assign 2_n9511 = ~(2_n10830 | 2_n1631);
assign 2_n9785 = 2_n11552 | 2_n4875;
assign 2_n6583 = 2_n9751 | 2_n10758;
assign 2_n1124 = ~(2_n1826 ^ 2_n8280);
assign 2_n10648 = 2_n2380 & 2_n8177;
assign 2_n10717 = 2_n10163 | 2_n10321;
assign 2_n9694 = ~2_n5845;
assign 2_n11316 = ~2_n5978;
assign 2_n9109 = ~(2_n1715 ^ 2_n2961);
assign 2_n12655 = ~2_n7442;
assign 2_n2029 = ~(2_n3180 ^ 2_n10086);
assign 2_n11082 = ~2_n167;
assign 2_n6186 = 2_n8480 & 2_n5865;
assign 2_n9901 = ~(2_n4948 ^ 2_n11275);
assign 2_n6230 = 2_n10424 | 2_n7245;
assign 2_n834 = ~2_n990;
assign 2_n8694 = 2_n7449 | 2_n5502;
assign 2_n7185 = 2_n12119 | 2_n8259;
assign 2_n3573 = ~(2_n2 | 2_n11783);
assign 2_n10818 = 2_n12263 | 2_n9203;
assign 2_n12919 = ~(2_n2570 ^ 2_n5038);
assign 2_n7535 = ~(2_n12286 ^ 2_n11836);
assign 2_n10191 = 2_n9730 & 2_n3306;
assign 2_n6580 = ~(2_n10324 ^ 2_n7333);
assign 2_n6790 = 2_n12341 | 2_n3075;
assign 2_n2739 = 2_n12199 & 2_n4028;
assign 2_n8750 = 2_n10762 & 2_n11365;
assign 2_n630 = 2_n8598 & 2_n5581;
assign 2_n10790 = 2_n1183 | 2_n3224;
assign 2_n10280 = 2_n3066 & 2_n8669;
assign 2_n8549 = 2_n2791 | 2_n278;
assign 2_n12396 = 2_n11245 & 2_n2673;
assign 2_n3560 = 2_n3905 & 2_n2270;
assign 2_n7655 = 2_n10157 | 2_n4864;
assign 2_n8143 = 2_n4916 | 2_n1263;
assign 2_n5 = ~(2_n11790 ^ 2_n2280);
assign 2_n11324 = 2_n8026 | 2_n7558;
assign 2_n6661 = 2_n1941 | 2_n5540;
assign 2_n6704 = 2_n6373 | 2_n9521;
assign 2_n6749 = 2_n58 & 2_n12426;
assign 2_n12224 = ~(2_n11721 ^ 2_n4146);
assign 2_n3056 = 2_n5990 & 2_n11078;
assign 2_n3340 = 2_n11026 | 2_n1476;
assign 2_n5781 = ~2_n1353;
assign 2_n5048 = 2_n10360 & 2_n12013;
assign 2_n6170 = ~2_n1306;
assign 2_n11655 = ~2_n12219;
assign 2_n5773 = ~2_n12520;
assign 2_n4948 = 2_n8870 | 2_n5326;
assign 2_n12384 = ~2_n11884;
assign 2_n5974 = ~2_n7778;
assign 2_n11387 = 2_n9426 | 2_n5790;
assign 2_n651 = ~2_n8048;
assign 2_n8608 = ~2_n7151;
assign 2_n10993 = 2_n6671 | 2_n4526;
assign 2_n6188 = ~(2_n8013 ^ 2_n1075);
assign 2_n8037 = ~(2_n8162 | 2_n9845);
assign 2_n3679 = ~2_n7187;
assign 2_n12023 = 2_n752 | 2_n3421;
assign 2_n11997 = 2_n1796 & 2_n10623;
assign 2_n12445 = ~(2_n3794 ^ 2_n12285);
assign 2_n8342 = 2_n2052 & 2_n1367;
assign 2_n4288 = ~2_n6879;
assign 2_n3957 = 2_n6738 & 2_n11179;
assign 2_n5968 = ~(2_n11182 ^ 2_n4200);
assign 2_n12061 = 2_n1699 | 2_n8109;
assign 2_n2471 = ~(2_n1991 ^ 2_n6692);
assign 2_n3281 = ~(2_n8602 ^ 2_n5897);
assign 2_n2569 = 2_n11511 & 2_n6885;
assign 2_n1645 = 2_n12647 ^ 2_n10665;
assign 2_n7229 = ~(2_n12742 ^ 2_n11768);
assign 2_n12353 = ~(2_n8515 ^ 2_n6760);
assign 2_n5564 = 2_n3892 | 2_n10358;
assign 2_n1502 = 2_n11528 & 2_n2654;
assign 2_n12309 = ~(2_n11908 ^ 2_n7578);
assign 2_n6927 = ~(2_n8155 | 2_n4408);
assign 2_n12751 = ~(2_n9059 ^ 2_n6865);
assign 2_n11267 = 2_n4056 & 2_n2169;
assign 2_n11585 = ~(2_n3837 ^ 2_n9096);
assign 2_n11840 = 2_n10670 & 2_n5488;
assign 2_n4596 = 2_n1100 | 2_n7763;
assign 2_n11785 = 2_n7688 & 2_n11465;
assign 2_n11567 = 2_n7587 | 2_n2343;
assign 2_n12830 = 2_n2697 & 2_n11348;
assign 2_n11411 = ~2_n2470;
assign 2_n11073 = ~(2_n1782 ^ 2_n12598);
assign 2_n12172 = ~2_n6660;
assign 2_n3225 = ~(2_n10909 | 2_n3496);
assign 2_n9577 = ~(2_n1956 ^ 2_n8570);
assign 2_n3907 = 2_n1993 | 2_n5090;
assign 2_n11747 = 2_n5840 | 2_n6614;
assign 2_n5134 = 2_n11036 | 2_n8030;
assign 2_n11210 = ~(2_n4489 ^ 2_n7013);
assign 2_n12598 = ~2_n4834;
assign 2_n11037 = 2_n8870 | 2_n4913;
assign 2_n2811 = 2_n1653 & 2_n10896;
assign 2_n12030 = ~2_n4999;
assign 2_n12324 = 2_n11958 | 2_n8768;
assign 2_n5973 = 2_n7889 & 2_n11993;
assign 2_n5421 = ~(2_n9764 ^ 2_n3997);
assign 2_n555 = 2_n3011 & 2_n8660;
assign 2_n10054 = ~(2_n3369 | 2_n9471);
assign 2_n7422 = ~2_n10009;
assign 2_n3308 = 2_n7251 & 2_n4264;
assign 2_n12417 = 2_n2045 & 2_n11274;
assign 2_n1521 = 2_n4696 | 2_n2475;
assign 2_n6048 = ~2_n3824;
assign 2_n2729 = ~(2_n9522 ^ 2_n2205);
assign 2_n1021 = 2_n11283 | 2_n12773;
assign 2_n4205 = 2_n1941 | 2_n7876;
assign 2_n11167 = ~(2_n10560 ^ 2_n2889);
assign 2_n7018 = ~(2_n4942 ^ 2_n7580);
assign 2_n1746 = 2_n10835 | 2_n8285;
assign 2_n4834 = 2_n2530 & 2_n2802;
assign 2_n5523 = ~2_n5291;
assign 2_n5786 = 2_n7283 | 2_n5497;
assign 2_n8696 = ~(2_n11029 ^ 2_n10800);
assign 2_n8590 = 2_n8687 | 2_n28;
assign 2_n1163 = ~2_n11922;
assign 2_n10298 = ~(2_n9489 | 2_n8935);
assign 2_n4295 = 2_n167 | 2_n408;
assign 2_n6592 = 2_n2025 | 2_n5322;
assign 2_n6115 = 2_n12262 | 2_n8253;
assign 2_n3025 = ~2_n5728;
assign 2_n3759 = ~2_n2714;
assign 2_n12819 = 2_n8949 | 2_n6724;
assign 2_n12297 = ~2_n7331;
assign 2_n2214 = 2_n8332 | 2_n10866;
assign 2_n7014 = 2_n11550 | 2_n7051;
assign 2_n5494 = ~(2_n10257 | 2_n8868);
assign 2_n4049 = ~(2_n4212 ^ 2_n1485);
assign 2_n4769 = 2_n4176 | 2_n3948;
assign 2_n11442 = ~(2_n6464 ^ 2_n9143);
assign 2_n7473 = 2_n8848 | 2_n1008;
assign 2_n9322 = 2_n6718 | 2_n4474;
assign 2_n794 = 2_n2950 & 2_n1164;
assign 2_n11555 = ~(2_n12445 ^ 2_n1351);
assign 2_n8842 = ~2_n4028;
assign 2_n375 = ~2_n11834;
assign 2_n2127 = 2_n10157 | 2_n12771;
assign 2_n3556 = ~2_n625;
assign 2_n336 = ~(2_n7978 ^ 2_n4997);
assign 2_n7954 = 2_n5283 & 2_n521;
assign 2_n950 = ~(2_n6221 ^ 2_n11379);
assign 2_n11184 = 2_n3096 | 2_n1413;
assign 2_n43 = 2_n925 & 2_n1958;
assign 2_n10902 = 2_n9655 | 2_n12580;
assign 2_n6526 = ~2_n10243;
assign 2_n11923 = ~2_n5314;
assign 2_n3548 = ~2_n1822;
assign 2_n12541 = 2_n9400 & 2_n10439;
assign 2_n10527 = 2_n3324 | 2_n4527;
assign 2_n8949 = 2_n5575 | 2_n3468;
assign 2_n1535 = ~(2_n6954 ^ 2_n3812);
assign 2_n8110 = ~(2_n3079 ^ 2_n9237);
assign 2_n1600 = ~2_n1294;
assign 2_n11856 = 2_n8428 | 2_n9741;
assign 2_n8101 = 2_n1760 & 2_n2859;
assign 2_n11188 = ~(2_n5277 ^ 2_n6240);
assign 2_n3723 = ~(2_n12354 ^ 2_n7165);
assign 2_n3873 = 2_n6977 | 2_n5538;
assign 2_n11225 = 2_n12069 & 2_n1512;
assign 2_n102 = 2_n4734 & 2_n11489;
assign 2_n6318 = 2_n1941 | 2_n1413;
assign 2_n8993 = ~(2_n10945 ^ 2_n5348);
assign 2_n5631 = ~2_n2030;
assign 2_n10443 = 2_n4150 & 2_n4627;
assign 2_n11903 = ~(2_n11831 | 2_n12798);
assign 2_n1253 = ~2_n812;
assign 2_n11146 = ~(2_n12935 ^ 2_n9808);
assign 2_n8455 = 2_n6411 & 2_n4132;
assign 2_n2905 = 2_n8026 | 2_n6114;
assign 2_n7072 = ~(2_n2726 ^ 2_n3289);
assign 2_n12862 = 2_n10712 | 2_n5583;
assign 2_n9193 = 2_n1226 & 2_n2750;
assign 2_n1962 = 2_n10135 | 2_n9854;
assign 2_n11321 = 2_n4120 & 2_n2805;
assign 2_n9674 = 2_n191 | 2_n1738;
assign 2_n7132 = ~(2_n3387 ^ 2_n12334);
assign 2_n8174 = ~(2_n2567 ^ 2_n2455);
assign 2_n3371 = ~(2_n2928 ^ 2_n12650);
assign 2_n11619 = ~2_n11017;
assign 2_n1391 = ~2_n2937;
assign 2_n11230 = 2_n10772 & 2_n10793;
assign 2_n10273 = ~(2_n10997 ^ 2_n10940);
assign 2_n6500 = ~(2_n3936 ^ 2_n1946);
assign 2_n10264 = ~(2_n8176 ^ 2_n324);
assign 2_n3802 = ~(2_n10722 ^ 2_n5535);
assign 2_n2633 = 2_n7084 & 2_n9091;
assign 2_n10929 = 2_n3820 | 2_n28;
assign 2_n4581 = 2_n3316 & 2_n7888;
assign 2_n11255 = 2_n2155 | 2_n11112;
assign 2_n4204 = ~2_n3247;
assign 2_n9038 = 2_n2718 & 2_n4611;
assign 2_n577 = 2_n8354 | 2_n826;
assign 2_n103 = ~(2_n3130 ^ 2_n7555);
assign 2_n4365 = ~2_n5263;
assign 2_n10778 = 2_n4383 | 2_n6297;
assign 2_n4812 = 2_n10590 | 2_n7821;
assign 2_n1829 = 2_n6373 | 2_n7921;
assign 2_n1517 = ~(2_n3970 ^ 2_n7091);
assign 2_n12663 = ~(2_n11080 | 2_n12597);
assign 2_n11473 = ~2_n3825;
assign 2_n12957 = ~2_n7807;
assign 2_n1208 = ~(2_n4788 | 2_n9620);
assign 2_n5987 = ~(2_n5492 ^ 2_n10072);
assign 2_n6495 = ~(2_n5921 ^ 2_n7360);
assign 2_n7476 = ~2_n6527;
assign 2_n9074 = ~2_n5582;
assign 2_n7934 = ~(2_n2993 ^ 2_n6468);
assign 2_n12539 = 2_n7116 | 2_n11896;
assign 2_n4163 = ~(2_n9926 ^ 2_n1969);
assign 2_n7372 = ~(2_n9305 | 2_n6205);
assign 2_n5233 = 2_n5964 & 2_n2577;
assign 2_n3659 = 2_n5575 | 2_n6114;
assign 2_n11228 = ~2_n2443;
assign 2_n12070 = 2_n6893 & 2_n1068;
assign 2_n6240 = ~(2_n5087 ^ 2_n5357);
assign 2_n8779 = 2_n8026 | 2_n12816;
assign 2_n11445 = ~(2_n9613 ^ 2_n4425);
assign 2_n9465 = 2_n4312 & 2_n7456;
assign 2_n9413 = 2_n11958 | 2_n995;
assign 2_n1203 = ~(2_n10703 ^ 2_n12311);
assign 2_n7197 = ~(2_n9438 | 2_n8982);
assign 2_n4076 = ~(2_n12176 ^ 2_n7150);
assign 2_n11392 = 2_n6718 | 2_n5502;
assign 2_n12852 = ~(2_n9043 ^ 2_n10840);
assign 2_n6729 = 2_n3848 & 2_n4974;
assign 2_n7769 = ~(2_n9643 | 2_n10076);
assign 2_n8054 = 2_n1937 | 2_n6169;
assign 2_n10868 = 2_n5832 & 2_n6531;
assign 2_n6815 = ~(2_n6341 ^ 2_n4419);
assign 2_n6463 = 2_n3007 | 2_n8561;
assign 2_n60 = 2_n11958 | 2_n6084;
assign 2_n478 = 2_n8337 & 2_n5622;
assign 2_n2884 = ~(2_n10918 ^ 2_n6420);
assign 2_n8361 = ~(2_n9392 ^ 2_n7263);
assign 2_n9964 = 2_n1223 & 2_n2892;
assign 2_n11638 = ~2_n12564;
assign 2_n4699 = 2_n11572 | 2_n3192;
assign 2_n10518 = 2_n6718 | 2_n9160;
assign 2_n7687 = ~2_n2643;
assign 2_n692 = ~2_n8694;
assign 2_n5402 = ~2_n1481;
assign 2_n12079 = ~2_n649;
assign 2_n6853 = 2_n962 | 2_n28;
assign 2_n9589 = ~2_n9725;
assign 2_n5797 = 2_n9370 | 2_n1162;
assign 2_n5971 = 2_n6914 & 2_n4447;
assign 2_n1056 = ~(2_n2763 ^ 2_n12633);
assign 2_n11456 = 2_n3617 | 2_n10854;
assign 2_n2685 = ~(2_n12960 ^ 2_n10487);
assign 2_n3680 = ~(2_n9722 ^ 2_n3739);
assign 2_n8156 = 2_n9360 & 2_n7633;
assign 2_n2247 = 2_n4859 & 2_n2263;
assign 2_n7565 = ~(2_n10615 ^ 2_n4523);
assign 2_n9331 = 2_n7872 & 2_n9468;
assign 2_n2846 = 2_n2099 | 2_n4249;
assign 2_n2461 = 2_n8737 & 2_n5874;
assign 2_n12715 = ~(2_n10866 ^ 2_n8332);
assign 2_n10760 = ~2_n12360;
assign 2_n6330 = ~(2_n12533 ^ 2_n9996);
assign 2_n7556 = ~(2_n1642 ^ 2_n6707);
assign 2_n3334 = ~(2_n5301 | 2_n8701);
assign 2_n1553 = ~(2_n8390 ^ 2_n757);
assign 2_n6636 = ~2_n11844;
assign 2_n4196 = 2_n12146 & 2_n10609;
assign 2_n1615 = ~(2_n9130 ^ 2_n9279);
assign 2_n10467 = 2_n4628 | 2_n12124;
assign 2_n10272 = ~(2_n10769 ^ 2_n2241);
assign 2_n7886 = 2_n10108 | 2_n11746;
assign 2_n3055 = ~(2_n8111 ^ 2_n9012);
assign 2_n10000 = ~(2_n6466 ^ 2_n6079);
assign 2_n12078 = ~2_n8913;
assign 2_n12442 = ~2_n10560;
assign 2_n348 = 2_n5589 | 2_n11291;
assign 2_n6766 = 2_n12256 | 2_n195;
assign 2_n6406 = 2_n2968 ^ 2_n4306;
assign 2_n3540 = ~2_n382;
assign 2_n9913 = 2_n636 | 2_n6071;
assign 2_n5398 = 2_n3389 & 2_n10001;
assign 2_n11281 = 2_n12119 | 2_n12754;
assign 2_n7998 = 2_n5575 | 2_n11820;
assign 2_n12267 = 2_n9705 & 2_n971;
assign 2_n11410 = ~2_n10451;
assign 2_n5676 = ~(2_n4500 ^ 2_n3469);
assign 2_n10245 = ~(2_n1331 ^ 2_n12919);
assign 2_n4020 = ~(2_n8920 ^ 2_n295);
assign 2_n12459 = ~(2_n7176 ^ 2_n506);
assign 2_n10156 = 2_n7986 | 2_n968;
assign 2_n234 = ~(2_n8778 ^ 2_n955);
assign 2_n8010 = ~2_n83;
assign 2_n4000 = ~(2_n10808 ^ 2_n2529);
assign 2_n2055 = 2_n5876 & 2_n5307;
assign 2_n10406 = ~(2_n4387 ^ 2_n4894);
assign 2_n7689 = ~(2_n84 | 2_n9350);
assign 2_n5900 = ~(2_n1364 ^ 2_n1517);
assign 2_n9747 = ~(2_n885 ^ 2_n5836);
assign 2_n2028 = ~(2_n7672 ^ 2_n220);
assign 2_n792 = 2_n7090 | 2_n7255;
assign 2_n7104 = ~(2_n1863 | 2_n11916);
assign 2_n8657 = ~(2_n10143 ^ 2_n909);
assign 2_n3879 = ~(2_n5736 ^ 2_n9955);
assign 2_n9493 = ~(2_n7088 ^ 2_n2926);
assign 2_n8076 = ~(2_n7775 ^ 2_n8490);
assign 2_n12483 = ~(2_n774 | 2_n5608);
assign 2_n12599 = 2_n9389 | 2_n7246;
assign 2_n6607 = ~2_n12611;
assign 2_n2244 = 2_n1144 & 2_n5210;
assign 2_n4773 = ~2_n4390;
assign 2_n12766 = 2_n7169 & 2_n1238;
assign 2_n1026 = 2_n1215 | 2_n5055;
assign 2_n11599 = ~2_n12893;
assign 2_n2040 = 2_n6073 | 2_n8947;
assign 2_n894 = 2_n7449 | 2_n9160;
assign 2_n4680 = ~(2_n7355 ^ 2_n5444);
assign 2_n12233 = ~(2_n324 | 2_n5686);
assign 2_n6606 = 2_n12361 | 2_n8414;
assign 2_n3277 = 2_n11241 | 2_n7689;
assign 2_n2824 = 2_n4805 & 2_n5645;
assign 2_n6517 = ~(2_n11268 ^ 2_n3525);
assign 2_n6443 = ~(2_n4570 ^ 2_n9874);
assign 2_n9593 = 2_n6231 & 2_n3444;
assign 2_n4835 = ~2_n7784;
assign 2_n174 = ~(2_n6575 | 2_n9458);
assign 2_n12146 = 2_n1803 | 2_n6421;
assign 2_n2424 = 2_n12119 | 2_n7382;
assign 2_n5315 = ~(2_n1315 ^ 2_n2211);
assign 2_n12838 = ~(2_n7112 ^ 2_n12654);
assign 2_n6564 = 2_n3743 | 2_n8745;
assign 2_n7936 = ~(2_n4409 ^ 2_n11220);
assign 2_n10458 = 2_n994 | 2_n11746;
assign 2_n1563 = 2_n9519 & 2_n9023;
assign 2_n2453 = 2_n4737 | 2_n5932;
assign 2_n1698 = ~(2_n1653 ^ 2_n10896);
assign 2_n11363 = 2_n2072 & 2_n3908;
assign 2_n10426 = ~2_n12452;
assign 2_n9476 = 2_n10879 | 2_n6389;
assign 2_n8380 = 2_n4697 & 2_n6968;
assign 2_n5032 = 2_n6418 | 2_n729;
assign 2_n1711 = ~(2_n11056 | 2_n1535);
assign 2_n10999 = ~(2_n5194 | 2_n8710);
assign 2_n11843 = ~2_n12052;
assign 2_n804 = 2_n1937 | 2_n10903;
assign 2_n4463 = 2_n5964 & 2_n9956;
assign 2_n9780 = 2_n3995 | 2_n482;
assign 2_n8523 = ~2_n5353;
assign 2_n1455 = ~2_n9956;
assign 2_n4456 = ~2_n758;
assign 2_n5754 = 2_n6307 & 2_n4636;
assign 2_n9324 = ~(2_n11836 | 2_n12286);
assign 2_n1390 = ~(2_n10307 ^ 2_n999);
assign 2_n1235 = 2_n4892 & 2_n583;
assign 2_n11108 = ~(2_n2640 ^ 2_n12181);
assign 2_n7878 = ~(2_n7130 ^ 2_n11464);
assign 2_n8325 = 2_n3820 | 2_n8830;
assign 2_n5648 = ~(2_n386 ^ 2_n9354);
assign 2_n386 = 2_n8026 | 2_n7952;
assign 2_n3646 = 2_n1701 & 2_n3338;
assign 2_n11431 = 2_n9180 | 2_n11564;
assign 2_n236 = 2_n5530 | 2_n6071;
assign 2_n5498 = ~(2_n5608 ^ 2_n774);
assign 2_n11915 = ~(2_n2363 ^ 2_n10097);
assign 2_n6408 = 2_n9644 & 2_n4925;
assign 2_n10372 = ~(2_n12737 | 2_n1742);
assign 2_n946 = ~(2_n4808 ^ 2_n2166);
assign 2_n2851 = 2_n5283 & 2_n6254;
assign 2_n621 = 2_n9878 | 2_n8655;
assign 2_n4977 = 2_n7203 & 2_n3304;
assign 2_n83 = 2_n6706 & 2_n10702;
assign 2_n5506 = ~2_n11972;
assign 2_n8425 = ~(2_n3203 ^ 2_n9601);
assign 2_n10543 = ~(2_n3733 | 2_n8200);
assign 2_n4947 = 2_n12610 & 2_n7794;
assign 2_n9328 = 2_n10879 | 2_n1851;
assign 2_n561 = ~2_n10327;
assign 2_n9116 = ~(2_n1082 ^ 2_n11336);
assign 2_n10206 = 2_n12616 | 2_n10627;
assign 2_n7981 = ~(2_n11730 ^ 2_n6215);
assign 2_n12362 = 2_n636 | 2_n8648;
assign 2_n844 = ~(2_n2607 ^ 2_n5472);
assign 2_n10584 = 2_n5211 & 2_n9287;
assign 2_n7434 = 2_n2456 | 2_n12446;
assign 2_n327 = ~(2_n788 ^ 2_n12009);
assign 2_n10334 = 2_n12496 & 2_n10286;
assign 2_n8454 = ~2_n10870;
assign 2_n292 = ~(2_n433 ^ 2_n11705);
assign 2_n658 = ~(2_n10146 ^ 2_n1522);
assign 2_n1248 = ~(2_n5382 ^ 2_n2905);
assign 2_n8066 = 2_n4498 | 2_n4400;
assign 2_n6470 = 2_n5530 | 2_n12735;
assign 2_n5104 = ~(2_n2922 | 2_n5244);
assign 2_n1942 = ~(2_n9124 ^ 2_n11629);
assign 2_n6324 = ~(2_n3145 ^ 2_n1267);
assign 2_n114 = ~2_n12753;
assign 2_n9445 = ~2_n12562;
assign 2_n2907 = 2_n12061 | 2_n10900;
assign 2_n5849 = ~(2_n7762 ^ 2_n1213);
assign 2_n10405 = ~(2_n643 | 2_n11979);
assign 2_n11579 = 2_n2313 | 2_n2669;
assign 2_n5578 = ~(2_n5021 ^ 2_n1414);
assign 2_n10660 = 2_n3947 | 2_n172;
assign 2_n9041 = ~(2_n891 ^ 2_n4598);
assign 2_n1839 = 2_n11245 | 2_n2673;
assign 2_n1776 = 2_n9370 | 2_n7703;
assign 2_n12470 = 2_n1941 | 2_n10903;
assign 2_n8880 = 2_n10139 | 2_n3615;
assign 2_n7714 = ~2_n8160;
assign 2_n10731 = 2_n7337 | 2_n3400;
assign 2_n12569 = 2_n9365 & 2_n3307;
assign 2_n439 = 2_n596 | 2_n5716;
assign 2_n9551 = 2_n5503 & 2_n730;
assign 2_n7644 = ~(2_n5214 ^ 2_n2616);
assign 2_n3852 = 2_n4203 & 2_n7354;
assign 2_n5468 = ~2_n2498;
assign 2_n7562 = 2_n6003 | 2_n11614;
assign 2_n4940 = 2_n6385 | 2_n8468;
assign 2_n10030 = 2_n9112 | 2_n8186;
assign 2_n11472 = ~2_n7531;
assign 2_n12422 = 2_n1082 & 2_n919;
assign 2_n11600 = ~(2_n1662 ^ 2_n6713);
assign 2_n433 = ~(2_n5217 ^ 2_n9200);
assign 2_n932 = ~(2_n5039 ^ 2_n12358);
assign 2_n2688 = ~(2_n11714 ^ 2_n4251);
assign 2_n11831 = 2_n6101 ^ 2_n2023;
assign 2_n11569 = 2_n7391 | 2_n1455;
assign 2_n7472 = ~(2_n6584 ^ 2_n12702);
assign 2_n11427 = ~(2_n5685 ^ 2_n5658);
assign 2_n7838 = ~(2_n5761 ^ 2_n5831);
assign 2_n5199 = ~2_n2436;
assign 2_n8457 = ~(2_n161 ^ 2_n550);
assign 2_n6891 = ~(2_n12362 ^ 2_n9811);
assign 2_n7409 = 2_n1699 | 2_n3224;
assign 2_n11550 = ~(2_n6060 ^ 2_n299);
assign 2_n12609 = ~(2_n11633 ^ 2_n9647);
assign 2_n5738 = ~2_n8906;
assign 2_n3970 = 2_n5462 & 2_n4080;
assign 2_n7923 = ~(2_n9698 ^ 2_n12540);
assign 2_n12742 = 2_n5530 | 2_n8644;
assign 2_n9311 = 2_n3992 & 2_n159;
assign 2_n9002 = ~(2_n5899 | 2_n2928);
assign 2_n2935 = ~2_n2943;
assign 2_n6061 = ~(2_n1750 ^ 2_n2500);
assign 2_n4877 = 2_n4872 & 2_n12374;
assign 2_n12773 = 2_n947 & 2_n6533;
assign 2_n2416 = ~(2_n2933 ^ 2_n9760);
assign 2_n12428 = ~(2_n1309 ^ 2_n9602);
assign 2_n9357 = 2_n11626 | 2_n12763;
assign 2_n10979 = 2_n12495 & 2_n4729;
assign 2_n7761 = ~(2_n5525 ^ 2_n5552);
assign 2_n7458 = 2_n5945 | 2_n12816;
assign 2_n1548 = 2_n5355 | 2_n3911;
assign 2_n11710 = 2_n807 | 2_n1413;
assign 2_n12099 = 2_n3872 & 2_n2814;
assign 2_n11980 = ~2_n4314;
assign 2_n3547 = ~(2_n3790 ^ 2_n4106);
assign 2_n1412 = 2_n6091 & 2_n6855;
assign 2_n11094 = ~(2_n10493 ^ 2_n9947);
assign 2_n4616 = ~(2_n9943 ^ 2_n4488);
assign 2_n5701 = 2_n9190 & 2_n8079;
assign 2_n7250 = 2_n6525 | 2_n2860;
assign 2_n9182 = 2_n1990 | 2_n7635;
assign 2_n11168 = ~2_n3401;
assign 2_n8343 = 2_n9373 | 2_n1476;
assign 2_n12732 = ~(2_n8594 | 2_n10081);
assign 2_n9846 = 2_n5355 | 2_n8735;
assign 2_n12302 = 2_n7709 | 2_n4474;
assign 2_n9499 = 2_n6876 & 2_n6818;
assign 2_n6515 = 2_n8187 | 2_n510;
assign 2_n12284 = 2_n2099 | 2_n10422;
assign 2_n11933 = 2_n3974 & 2_n2041;
assign 2_n7817 = ~(2_n3210 | 2_n10527);
assign 2_n11846 = 2_n7449 | 2_n9568;
assign 2_n10194 = 2_n910 & 2_n9852;
assign 2_n4225 = 2_n9002 | 2_n2114;
assign 2_n2383 = ~(2_n8811 ^ 2_n9774);
assign 2_n3735 = ~2_n8235;
assign 2_n12462 = 2_n4911 | 2_n1546;
assign 2_n7065 = ~(2_n1878 | 2_n11494);
assign 2_n6196 = 2_n12447 | 2_n4665;
assign 2_n6706 = 2_n5331 & 2_n12489;
assign 2_n1265 = 2_n10542 & 2_n5178;
assign 2_n11519 = ~2_n12505;
assign 2_n12108 = ~(2_n2482 ^ 2_n2163);
assign 2_n6313 = 2_n11808 | 2_n1838;
assign 2_n6154 = ~2_n12448;
assign 2_n1215 = 2_n9389 | 2_n1851;
assign 2_n9789 = ~(2_n12368 | 2_n7583);
assign 2_n6969 = ~2_n11173;
assign 2_n12404 = 2_n11375 & 2_n6144;
assign 2_n3813 = ~2_n233;
assign 2_n8862 = ~(2_n4002 ^ 2_n6061);
assign 2_n2385 = ~(2_n613 ^ 2_n836);
assign 2_n11545 = ~(2_n5164 ^ 2_n513);
assign 2_n8166 = ~(2_n434 | 2_n11871);
assign 2_n10532 = 2_n5724 | 2_n8890;
assign 2_n11842 = 2_n5530 | 2_n10854;
assign 2_n3940 = 2_n12289 | 2_n9253;
assign 2_n4493 = ~2_n3852;
assign 2_n10474 = 2_n9803 | 2_n6160;
assign 2_n2697 = 2_n2761 | 2_n6288;
assign 2_n3690 = ~2_n12480;
assign 2_n10102 = 2_n6249 | 2_n251;
assign 2_n2350 = 2_n9208 & 2_n12696;
assign 2_n7659 = ~2_n10450;
assign 2_n11793 = ~2_n10845;
assign 2_n9790 = ~(2_n11335 ^ 2_n12278);
assign 2_n732 = ~2_n49;
assign 2_n1192 = 2_n12661 & 2_n2753;
assign 2_n3590 = ~2_n6974;
assign 2_n7751 = ~(2_n3176 ^ 2_n10322);
assign 2_n152 = ~(2_n7446 ^ 2_n1023);
assign 2_n12118 = 2_n5915 | 2_n12735;
assign 2_n11784 = ~(2_n11482 ^ 2_n10635);
assign 2_n7045 = ~(2_n12607 | 2_n10204);
assign 2_n515 = 2_n4628 | 2_n4818;
assign 2_n8963 = 2_n6577 | 2_n7425;
assign 2_n10169 = 2_n10835 | 2_n12120;
assign 2_n6275 = 2_n8103 | 2_n5741;
assign 2_n6647 = ~(2_n8550 ^ 2_n10934);
assign 2_n4744 = 2_n11189 & 2_n7922;
assign 2_n2538 = ~2_n12122;
assign 2_n6731 = ~(2_n7059 ^ 2_n3835);
assign 2_n734 = ~2_n10972;
assign 2_n7682 = 2_n3188 & 2_n689;
assign 2_n8944 = ~2_n3904;
assign 2_n12577 = ~2_n1275;
assign 2_n7790 = 2_n2217 | 2_n2020;
assign 2_n1692 = ~(2_n6231 ^ 2_n12103);
assign 2_n5120 = ~(2_n10773 ^ 2_n490);
assign 2_n12828 = ~(2_n3795 ^ 2_n8868);
assign 2_n2834 = ~(2_n6539 ^ 2_n47);
assign 2_n12420 = ~(2_n3301 ^ 2_n691);
assign 2_n7784 = ~(2_n12933 ^ 2_n8989);
assign 2_n6503 = ~(2_n3544 ^ 2_n3414);
assign 2_n10337 = ~2_n1124;
assign 2_n11539 = 2_n5231 | 2_n5217;
assign 2_n9865 = ~(2_n8869 ^ 2_n12806);
assign 2_n12614 = ~2_n2305;
assign 2_n12627 = ~(2_n2005 ^ 2_n3331);
assign 2_n11171 = 2_n3096 | 2_n7425;
assign 2_n3495 = 2_n693 & 2_n3069;
assign 2_n3439 = 2_n240 & 2_n983;
assign 2_n3780 = 2_n9098 | 2_n2812;
assign 2_n3914 = ~(2_n9198 ^ 2_n8640);
assign 2_n4917 = ~(2_n9479 ^ 2_n12515);
assign 2_n3906 = 2_n191 | 2_n5851;
assign 2_n4139 = ~(2_n9042 ^ 2_n11399);
assign 2_n4637 = 2_n5225 | 2_n1625;
assign 2_n4201 = 2_n12284 | 2_n663;
assign 2_n685 = ~2_n6002;
assign 2_n5659 = 2_n11060 & 2_n11247;
assign 2_n9075 = ~(2_n11842 ^ 2_n7027);
assign 2_n12461 = 2_n148 & 2_n3927;
assign 2_n2467 = ~(2_n772 ^ 2_n2645);
assign 2_n6870 = ~(2_n6800 | 2_n8436);
assign 2_n393 = 2_n719 & 2_n6314;
assign 2_n10129 = ~(2_n8015 | 2_n12716);
assign 2_n6435 = ~(2_n2136 ^ 2_n10652);
assign 2_n12800 = ~(2_n8444 | 2_n6693);
assign 2_n6545 = ~(2_n6805 ^ 2_n869);
assign 2_n5615 = ~(2_n7122 ^ 2_n746);
assign 2_n3980 = 2_n1126 | 2_n4143;
assign 2_n5118 = ~(2_n11240 | 2_n3993);
assign 2_n6260 = 2_n10829 & 2_n3589;
assign 2_n3523 = 2_n10835 | 2_n3599;
assign 2_n4385 = ~(2_n6939 ^ 2_n208);
assign 2_n10676 = ~(2_n203 ^ 2_n8447);
assign 2_n531 = ~(2_n6453 ^ 2_n7412);
assign 2_n120 = ~2_n8093;
assign 2_n7907 = ~(2_n7567 ^ 2_n11794);
assign 2_n604 = 2_n19 & 2_n4533;
assign 2_n11145 = 2_n2014 & 2_n9821;
assign 2_n11601 = 2_n4223 | 2_n1819;
assign 2_n2760 = 2_n8459 & 2_n11573;
assign 2_n4644 = 2_n3743 | 2_n4875;
assign 2_n10098 = ~2_n12047;
assign 2_n7467 = ~(2_n6318 ^ 2_n7064);
assign 2_n4982 = ~(2_n11514 | 2_n3012);
assign 2_n9198 = 2_n12485 | 2_n7670;
assign 2_n6554 = ~(2_n8231 ^ 2_n11135);
assign 2_n945 = 2_n11195 & 2_n9292;
assign 2_n8317 = 2_n9584 | 2_n2020;
assign 2_n3256 = 2_n4846 | 2_n11562;
assign 2_n4736 = ~2_n578;
assign 2_n11408 = ~(2_n12524 ^ 2_n2088);
assign 2_n9542 = ~(2_n12309 ^ 2_n10651);
assign 2_n10511 = 2_n2170 & 2_n1897;
assign 2_n5712 = 2_n11433 | 2_n9741;
assign 2_n672 = ~(2_n1346 ^ 2_n5163);
assign 2_n9940 = 2_n10879 | 2_n1162;
assign 2_n11559 = ~(2_n10693 ^ 2_n8709);
assign 2_n11929 = ~(2_n9897 ^ 2_n979);
assign 2_n11476 = ~(2_n9486 | 2_n1264);
assign 2_n8449 = 2_n8026 | 2_n8768;
assign 2_n10959 = ~(2_n7075 ^ 2_n4746);
assign 2_n6713 = ~(2_n5205 ^ 2_n3949);
assign 2_n6599 = 2_n9389 | 2_n1546;
assign 2_n1878 = 2_n11560 | 2_n9658;
assign 2_n12528 = 2_n5516 & 2_n6719;
assign 2_n7978 = ~(2_n3283 ^ 2_n2849);
assign 2_n6125 = ~(2_n709 | 2_n1568);
assign 2_n2374 = 2_n2832 | 2_n5497;
assign 2_n12668 = 2_n7449 | 2_n5914;
assign 2_n9102 = 2_n7690 & 2_n2558;
assign 2_n6397 = ~(2_n1028 | 2_n5924);
assign 2_n7345 = 2_n8256 & 2_n2373;
assign 2_n11798 = ~(2_n11669 ^ 2_n652);
assign 2_n8436 = ~(2_n5532 ^ 2_n8501);
assign 2_n8647 = ~(2_n11514 ^ 2_n7727);
assign 2_n10144 = 2_n12853 | 2_n12535;
assign 2_n9990 = 2_n1475 | 2_n4986;
assign 2_n5094 = ~(2_n11491 ^ 2_n12222);
assign 2_n8294 = 2_n11958 | 2_n184;
assign 2_n4132 = 2_n6134 | 2_n12401;
assign 2_n6685 = ~(2_n3354 | 2_n7607);
assign 2_n7841 = ~2_n7631;
assign 2_n5824 = 2_n12864 | 2_n9456;
assign 2_n3524 = 2_n11968 & 2_n6;
assign 2_n7200 = 2_n989 | 2_n12328;
assign 2_n12727 = 2_n10398 & 2_n1601;
assign 2_n11636 = ~(2_n722 ^ 2_n10325);
assign 2_n10556 = ~(2_n5079 ^ 2_n10084);
assign 2_n11598 = 2_n7449 | 2_n28;
assign 2_n4028 = 2_n2464 & 2_n5105;
assign 2_n2839 = 2_n6782 & 2_n7054;
assign 2_n9815 = ~2_n820;
assign 2_n4507 = ~(2_n688 ^ 2_n7853);
assign 2_n6253 = ~(2_n4907 ^ 2_n8766);
assign 2_n581 = 2_n10945 & 2_n7318;
assign 2_n9909 = 2_n9382 & 2_n3760;
assign 2_n9307 = 2_n752 | 2_n6169;
assign 2_n10847 = 2_n5355 | 2_n1079;
assign 2_n1324 = 2_n8476 & 2_n1564;
assign 2_n4889 = ~(2_n6861 | 2_n10985);
assign 2_n4804 = 2_n9313 & 2_n190;
assign 2_n4397 = 2_n165 ^ 2_n6990;
assign 2_n9266 = 2_n4628 | 2_n12080;
assign 2_n12215 = ~(2_n12603 ^ 2_n8696);
assign 2_n1677 = 2_n8996 | 2_n9518;
assign 2_n923 = ~(2_n11800 ^ 2_n7358);
assign 2_n3279 = 2_n12365 | 2_n11406;
assign 2_n3599 = ~2_n1906;
assign 2_n11402 = 2_n11493 | 2_n8122;
assign 2_n1589 = ~(2_n9391 ^ 2_n5302);
assign 2_n7194 = ~(2_n9114 ^ 2_n11581);
assign 2_n8245 = ~(2_n1205 ^ 2_n5617);
assign 2_n10284 = 2_n11740 & 2_n4969;
assign 2_n5730 = ~(2_n3202 ^ 2_n8683);
assign 2_n8598 = ~(2_n2440 ^ 2_n9261);
assign 2_n11310 = 2_n3243 & 2_n5880;
assign 2_n10963 = 2_n1282 & 2_n12458;
assign 2_n1586 = ~(2_n8840 ^ 2_n11315);
assign 2_n7884 = 2_n6656 | 2_n9548;
assign 2_n3504 = 2_n7398 & 2_n12219;
assign 2_n12246 = 2_n8738 | 2_n9160;
assign 2_n2212 = ~(2_n10112 | 2_n12547);
assign 2_n11746 = ~2_n3932;
assign 2_n2171 = ~2_n8521;
assign 2_n9001 = ~(2_n418 ^ 2_n207);
assign 2_n11808 = ~(2_n6954 | 2_n4912);
assign 2_n9261 = 2_n12194 & 2_n2351;
assign 2_n5650 = 2_n10835 | 2_n6138;
assign 2_n7387 = ~(2_n8737 ^ 2_n6644);
assign 2_n6522 = 2_n6271 | 2_n11420;
assign 2_n5387 = 2_n5858 | 2_n4400;
assign 2_n10211 = 2_n10387 & 2_n3019;
assign 2_n10756 = 2_n2010 & 2_n2261;
assign 2_n9929 = ~(2_n3694 ^ 2_n1849);
assign 2_n7815 = ~(2_n12071 ^ 2_n11230);
assign 2_n9257 = ~(2_n12177 ^ 2_n2430);
assign 2_n8592 = ~2_n6584;
assign 2_n6490 = ~2_n5093;
assign 2_n1095 = 2_n12701 | 2_n6897;
assign 2_n10208 = 2_n11547 & 2_n6832;
assign 2_n8910 = 2_n6686 & 2_n5407;
assign 2_n2118 = 2_n11162 & 2_n1302;
assign 2_n9403 = 2_n11936 & 2_n3346;
assign 2_n8281 = 2_n11478 & 2_n1564;
assign 2_n1109 = 2_n9266 & 2_n8711;
assign 2_n8233 = 2_n2319 & 2_n10252;
assign 2_n12166 = 2_n4950 & 2_n2596;
assign 2_n11872 = ~(2_n8892 ^ 2_n8906);
assign 2_n7673 = ~2_n9348;
assign 2_n6587 = 2_n4741 ^ 2_n7253;
assign 2_n1147 = 2_n12438 & 2_n8185;
assign 2_n10989 = ~(2_n10880 ^ 2_n7361);
assign 2_n12519 = ~(2_n7248 ^ 2_n12159);
assign 2_n3134 = 2_n8516 ^ 2_n4682;
assign 2_n2571 = 2_n7166 & 2_n11163;
assign 2_n5422 = 2_n8010 | 2_n12089;
assign 2_n7607 = ~2_n4427;
assign 2_n413 = 2_n3381 | 2_n10811;
assign 2_n12427 = ~2_n10802;
assign 2_n3643 = 2_n8816 & 2_n1084;
assign 2_n12142 = 2_n2456 | 2_n7382;
assign 2_n3508 = 2_n5575 | 2_n2589;
assign 2_n1174 = 2_n8959 | 2_n5012;
assign 2_n7507 = ~(2_n8389 ^ 2_n10747);
assign 2_n5628 = ~(2_n6008 ^ 2_n4581);
assign 2_n677 = 2_n7452 | 2_n8615;
assign 2_n12729 = 2_n443 & 2_n10200;
assign 2_n10508 = 2_n7911 & 2_n5323;
assign 2_n3860 = ~(2_n23 | 2_n7844);
assign 2_n8591 = ~(2_n1438 ^ 2_n6778);
assign 2_n3843 = 2_n114 | 2_n5012;
assign 2_n5375 = ~(2_n7230 | 2_n11019);
assign 2_n4092 = 2_n10354 & 2_n1502;
assign 2_n3520 = 2_n12853 | 2_n5468;
assign 2_n9164 = 2_n4778 | 2_n5468;
assign 2_n6844 = 2_n11887 | 2_n10854;
assign 2_n673 = ~2_n1317;
assign 2_n8937 = 2_n12220 & 2_n6388;
assign 2_n4346 = 2_n1941 | 2_n6197;
assign 2_n1444 = 2_n11851 | 2_n9255;
assign 2_n11346 = ~2_n12355;
assign 2_n5097 = ~(2_n2411 | 2_n8486);
assign 2_n11759 = ~2_n4930;
assign 2_n7590 = 2_n6971 | 2_n7178;
assign 2_n8872 = ~(2_n6581 ^ 2_n12820);
assign 2_n9663 = ~(2_n11988 ^ 2_n2374);
assign 2_n1797 = ~(2_n8938 | 2_n578);
assign 2_n7423 = 2_n4457 & 2_n622;
assign 2_n8921 = ~2_n2760;
assign 2_n5894 = ~(2_n3481 ^ 2_n575);
assign 2_n4611 = ~2_n6838;
assign 2_n1012 = 2_n191 | 2_n6402;
assign 2_n12923 = ~(2_n2019 ^ 2_n462);
assign 2_n193 = ~(2_n8452 ^ 2_n8978);
assign 2_n4219 = 2_n1449 | 2_n1174;
assign 2_n5184 = ~(2_n11442 ^ 2_n728);
assign 2_n7325 = 2_n9373 | 2_n9078;
assign 2_n11995 = ~(2_n6594 | 2_n6670);
assign 2_n1411 = ~(2_n1924 ^ 2_n10014);
assign 2_n5075 = ~(2_n9718 ^ 2_n3738);
assign 2_n7559 = ~(2_n7325 ^ 2_n8325);
assign 2_n11671 = 2_n3594 & 2_n7156;
assign 2_n7016 = ~(2_n3483 ^ 2_n12894);
assign 2_n10659 = 2_n9421 & 2_n1885;
assign 2_n437 = 2_n10429 | 2_n7158;
assign 2_n1802 = 2_n10064 & 2_n10905;
assign 2_n7445 = 2_n7537 | 2_n4803;
assign 2_n2421 = 2_n5800 & 2_n738;
assign 2_n10227 = ~(2_n12198 ^ 2_n4024);
assign 2_n5570 = 2_n8428 | 2_n11122;
assign 2_n8740 = ~2_n1067;
assign 2_n11714 = 2_n8870 | 2_n12535;
assign 2_n6738 = 2_n9389 | 2_n7424;
assign 2_n3065 = 2_n5809 | 2_n3924;
assign 2_n11755 = ~(2_n5327 ^ 2_n11912);
assign 2_n6494 = ~(2_n12895 ^ 2_n1834);
assign 2_n1882 = 2_n3717 | 2_n1894;
assign 2_n4764 = ~2_n9072;
assign 2_n703 = ~(2_n5049 ^ 2_n958);
assign 2_n11315 = ~(2_n3346 ^ 2_n3242);
assign 2_n6072 = 2_n6718 | 2_n9568;
assign 2_n1740 = 2_n8428 | 2_n6114;
assign 2_n12141 = 2_n10512 & 2_n2742;
assign 2_n10986 = ~2_n9805;
assign 2_n9939 = 2_n6136 | 2_n5835;
assign 2_n4326 = ~(2_n5978 ^ 2_n10597);
assign 2_n7809 = 2_n3628 | 2_n894;
assign 2_n3782 = 2_n2608 & 2_n4615;
assign 2_n12383 = ~(2_n9258 ^ 2_n2584);
assign 2_n12615 = ~(2_n11490 ^ 2_n10318);
assign 2_n6493 = ~2_n9467;
assign 2_n12080 = ~2_n5579;
assign 2_n10330 = ~2_n1984;
assign 2_n9508 = ~(2_n11208 ^ 2_n1911);
assign 2_n8532 = 2_n1371 & 2_n6392;
assign 2_n10061 = ~(2_n11955 ^ 2_n1819);
assign 2_n4242 = ~2_n4370;
assign 2_n7398 = ~2_n7206;
assign 2_n4195 = 2_n12186 | 2_n6455;
assign 2_n11563 = 2_n10835 | 2_n4654;
assign 2_n362 = ~2_n3715;
assign 2_n754 = ~(2_n10582 | 2_n6998);
assign 2_n1837 = 2_n7773 & 2_n1633;
assign 2_n6754 = ~(2_n3711 ^ 2_n912);
assign 2_n12875 = 2_n3240 & 2_n8801;
assign 2_n11221 = 2_n10142 | 2_n7424;
assign 2_n4156 = ~(2_n1021 ^ 2_n3502);
assign 2_n6555 = ~(2_n1258 ^ 2_n7250);
assign 2_n12266 = 2_n9739 & 2_n7224;
assign 2_n10725 = 2_n9266 | 2_n8711;
assign 2_n1806 = 2_n7839 | 2_n5012;
assign 2_n1796 = ~2_n6370;
assign 2_n11863 = ~2_n12292;
assign 2_n2869 = ~(2_n11575 ^ 2_n9057);
assign 2_n1783 = 2_n12891 | 2_n11506;
assign 2_n2763 = 2_n5355 | 2_n1851;
assign 2_n5311 = ~2_n783;
assign 2_n11857 = ~2_n11271;
assign 2_n271 = 2_n9389 | 2_n12843;
assign 2_n8055 = 2_n191 | 2_n10419;
assign 2_n3180 = 2_n10879 | 2_n7341;
assign 2_n11787 = 2_n12525 & 2_n3298;
assign 2_n4851 = 2_n8327 & 2_n2701;
assign 2_n9454 = 2_n4600 & 2_n410;
assign 2_n5397 = 2_n5809 | 2_n6513;
assign 2_n10047 = 2_n8720 & 2_n12064;
assign 2_n10126 = ~(2_n7653 ^ 2_n4688);
assign 2_n12661 = 2_n914 | 2_n2429;
assign 2_n12951 = ~(2_n2539 ^ 2_n5910);
assign 2_n4953 = 2_n5305 & 2_n5212;
assign 2_n6007 = 2_n12051 & 2_n3091;
assign 2_n10899 = 2_n5501 | 2_n4792;
assign 2_n3422 = 2_n12070 | 2_n2621;
assign 2_n1988 = 2_n6158 | 2_n3052;
assign 2_n3896 = 2_n9081 & 2_n6258;
assign 2_n998 = 2_n11324 | 2_n12756;
assign 2_n11372 = ~(2_n7793 ^ 2_n536);
assign 2_n12840 = 2_n7865 | 2_n12338;
assign 2_n319 = ~(2_n9455 | 2_n513);
assign 2_n7990 = ~(2_n2058 ^ 2_n4218);
assign 2_n7699 = 2_n12063 & 2_n12149;
assign 2_n10328 = ~(2_n1810 ^ 2_n7990);
assign 2_n6996 = ~(2_n10404 ^ 2_n1132);
assign 2_n2588 = ~(2_n9270 ^ 2_n6356);
assign 2_n1524 = 2_n1516 & 2_n2189;
assign 2_n4090 = ~(2_n1371 ^ 2_n690);
assign 2_n10629 = ~2_n6760;
assign 2_n10316 = ~2_n3094;
assign 2_n6695 = 2_n3746 | 2_n5012;
assign 2_n9757 = 2_n12936 & 2_n6796;
assign 2_n1603 = ~(2_n9492 ^ 2_n4546);
assign 2_n6999 = ~2_n9167;
assign 2_n9709 = ~2_n2089;
assign 2_n6056 = ~(2_n1947 ^ 2_n3151);
assign 2_n12716 = 2_n10093 | 2_n12105;
assign 2_n4840 = ~(2_n12198 | 2_n1562);
assign 2_n2324 = 2_n6767 | 2_n6250;
assign 2_n7744 = ~(2_n6853 | 2_n5076);
assign 2_n12482 = ~(2_n9443 ^ 2_n7377);
assign 2_n2626 = 2_n8428 | 2_n11820;
assign 2_n1864 = ~(2_n5907 ^ 2_n5343);
assign 2_n10070 = ~2_n10844;
assign 2_n4266 = 2_n1549 | 2_n10856;
assign 2_n9163 = ~(2_n3135 ^ 2_n11057);
assign 2_n8728 = ~(2_n2071 ^ 2_n10323);
assign 2_n12278 = 2_n10157 | 2_n7921;
assign 2_n12115 = 2_n9707 & 2_n6526;
assign 2_n11658 = 2_n1779 | 2_n4685;
assign 2_n4497 = ~(2_n5661 ^ 2_n7164);
assign 2_n390 = 2_n10962 & 2_n9333;
assign 2_n2178 = 2_n1341 & 2_n9522;
assign 2_n9809 = ~(2_n11069 ^ 2_n11128);
assign 2_n9505 = ~2_n1240;
assign 2_n12743 = 2_n7709 | 2_n4654;
assign 2_n1493 = 2_n9370 | 2_n2358;
assign 2_n867 = ~(2_n12269 | 2_n7003);
assign 2_n3347 = ~2_n10648;
assign 2_n12045 = 2_n8369 | 2_n4108;
assign 2_n9518 = 2_n1699 | 2_n826;
assign 2_n793 = ~(2_n935 ^ 2_n606);
assign 2_n820 = 2_n994 | 2_n4400;
assign 2_n11778 = 2_n4237 | 2_n10229;
assign 2_n3167 = ~(2_n11339 ^ 2_n9224);
assign 2_n2067 = ~2_n20;
assign 2_n4255 = 2_n9037 | 2_n448;
assign 2_n11451 = 2_n3820 | 2_n3606;
assign 2_n7594 = ~(2_n7756 | 2_n4681);
assign 2_n5205 = 2_n8755 & 2_n6648;
assign 2_n11921 = ~(2_n12226 ^ 2_n6340);
assign 2_n11365 = 2_n11892 & 2_n7294;
assign 2_n2651 = ~(2_n3353 | 2_n5545);
assign 2_n1994 = 2_n5964 & 2_n1798;
assign 2_n10703 = ~(2_n11704 ^ 2_n2368);
assign 2_n9917 = ~2_n10488;
assign 2_n4743 = ~(2_n8828 ^ 2_n4123);
assign 2_n4261 = 2_n4911 | 2_n4242;
assign 2_n7356 = ~2_n3250;
assign 2_n7421 = 2_n4360 | 2_n8396;
assign 2_n7925 = 2_n2186 & 2_n12453;
assign 2_n10043 = ~(2_n63 ^ 2_n11595);
assign 2_n12681 = 2_n3480 & 2_n2611;
assign 2_n12756 = 2_n1107 & 2_n5287;
assign 2_n3288 = ~(2_n3136 ^ 2_n8886);
assign 2_n107 = 2_n12119 | 2_n12080;
assign 2_n7146 = 2_n10520 & 2_n543;
assign 2_n8775 = ~(2_n7929 ^ 2_n5588);
assign 2_n10523 = ~(2_n2934 | 2_n2353);
assign 2_n4870 = 2_n420 | 2_n10308;
assign 2_n7763 = ~(2_n11593 ^ 2_n4128);
assign 2_n9484 = ~2_n12934;
assign 2_n4419 = ~(2_n7034 | 2_n10058);
assign 2_n1079 = ~2_n10223;
assign 2_n2910 = 2_n1465 & 2_n6272;
assign 2_n12592 = ~(2_n10231 ^ 2_n993);
assign 2_n4257 = 2_n1246 & 2_n4355;
assign 2_n10920 = 2_n7383 & 2_n4893;
assign 2_n9068 = 2_n5765 | 2_n5759;
assign 2_n11717 = 2_n6365 | 2_n6285;
assign 2_n4655 = ~(2_n9684 ^ 2_n6936);
assign 2_n12437 = ~2_n3011;
assign 2_n9880 = 2_n12208 | 2_n10017;
assign 2_n12550 = 2_n2456 | 2_n12883;
assign 2_n12116 = 2_n3984 & 2_n3902;
assign 2_n8295 = 2_n5915 | 2_n1932;
assign 2_n3468 = ~2_n8717;
assign 2_n3890 = 2_n6707 | 2_n9870;
assign 2_n8104 = ~(2_n7348 ^ 2_n1806);
assign 2_n8833 = ~(2_n2773 ^ 2_n1718);
assign 2_n12178 = 2_n7391 | 2_n1546;
assign 2_n7871 = 2_n3127 | 2_n510;
assign 2_n2483 = ~2_n3742;
assign 2_n8716 = ~(2_n4804 | 2_n9957);
assign 2_n1725 = ~(2_n8903 ^ 2_n5834);
assign 2_n1403 = ~2_n4734;
assign 2_n1800 = 2_n8583 | 2_n28;
assign 2_n12378 = ~(2_n23 ^ 2_n1830);
assign 2_n5668 = ~(2_n3676 ^ 2_n3173);
assign 2_n12929 = ~2_n38;
assign 2_n3664 = 2_n11546 & 2_n4638;
assign 2_n32 = ~(2_n7559 ^ 2_n4712);
assign 2_n6010 = 2_n1406 | 2_n12168;
assign 2_n2173 = ~(2_n445 ^ 2_n9866);
assign 2_n7836 = ~(2_n1111 ^ 2_n7959);
assign 2_n4987 = ~(2_n4976 | 2_n5657);
assign 2_n1704 = ~2_n8270;
assign 2_n1149 = 2_n11147 | 2_n12290;
assign 2_n10889 = ~(2_n9965 ^ 2_n6803);
assign 2_n4683 = ~(2_n21 ^ 2_n3705);
assign 2_n7963 = 2_n9600 & 2_n7860;
assign 2_n6854 = 2_n3837 & 2_n9096;
assign 2_n7807 = 2_n6770 & 2_n4634;
assign 2_n10536 = ~(2_n8445 | 2_n8754);
assign 2_n1892 = ~(2_n12770 | 2_n8877);
assign 2_n3387 = ~(2_n3215 ^ 2_n567);
assign 2_n11707 = ~(2_n6942 ^ 2_n10303);
assign 2_n6569 = 2_n7839 | 2_n6455;
assign 2_n11491 = 2_n8153 & 2_n10266;
assign 2_n7574 = 2_n3820 | 2_n4642;
assign 2_n8229 = 2_n10750 | 2_n8655;
assign 2_n7583 = ~(2_n7764 | 2_n6710);
assign 2_n10947 = 2_n4312 & 2_n4634;
assign 2_n3153 = 2_n10750 | 2_n4913;
assign 2_n8626 = ~2_n12794;
assign 2_n2541 = ~(2_n298 ^ 2_n4919);
assign 2_n10686 = ~(2_n12506 ^ 2_n2489);
assign 2_n1774 = ~(2_n9269 | 2_n9169);
assign 2_n2974 = ~2_n10993;
assign 2_n5364 = 2_n3617 | 2_n3224;
assign 2_n10053 = 2_n3667 | 2_n5580;
assign 2_n6169 = ~2_n7354;
assign 2_n4796 = 2_n6470 & 2_n7392;
assign 2_n5898 = ~(2_n5869 ^ 2_n7231);
assign 2_n1363 = ~(2_n6895 ^ 2_n414);
assign 2_n9003 = 2_n3818 | 2_n10716;
assign 2_n6920 = ~(2_n3268 ^ 2_n1045);
assign 2_n3023 = 2_n91 | 2_n3162;
assign 2_n2847 = 2_n630 | 2_n12394;
assign 2_n3859 = ~2_n8573;
assign 2_n1505 = 2_n10781 & 2_n4941;
assign 2_n8803 = ~2_n8477;
assign 2_n10694 = ~(2_n8161 ^ 2_n8218);
assign 2_n1536 = ~(2_n10984 ^ 2_n11643);
assign 2_n5481 = ~(2_n3984 ^ 2_n3902);
assign 2_n3628 = 2_n10835 | 2_n9144;
assign 2_n10712 = ~2_n8605;
assign 2_n25 = ~2_n12201;
assign 2_n1533 = 2_n4479 | 2_n859;
assign 2_n3962 = ~2_n7309;
assign 2_n231 = 2_n10049 & 2_n1521;
assign 2_n12167 = 2_n7283 | 2_n4775;
assign 2_n1715 = 2_n11026 | 2_n795;
assign 2_n636 = ~2_n7891;
assign 2_n6596 = ~2_n2296;
assign 2_n10577 = ~(2_n5928 | 2_n3511);
assign 2_n9233 = ~2_n3255;
assign 2_n12325 = ~(2_n4696 ^ 2_n416);
assign 2_n1815 = 2_n9657 & 2_n1807;
assign 2_n7124 = ~2_n3202;
assign 2_n124 = 2_n10055 | 2_n12613;
assign 2_n10602 = 2_n2979 & 2_n4298;
assign 2_n8475 = 2_n752 | 2_n7876;
assign 2_n11726 = 2_n9179 & 2_n9479;
assign 2_n10735 = 2_n10142 | 2_n1915;
assign 2_n2559 = 2_n4193 | 2_n12637;
assign 2_n9289 = 2_n6797 & 2_n5645;
assign 2_n11434 = 2_n2677 & 2_n9579;
assign 2_n12311 = ~(2_n8036 ^ 2_n10094);
assign 2_n10512 = 2_n5305 & 2_n2509;
assign 2_n9167 = 2_n11923 | 2_n8830;
assign 2_n3974 = 2_n12775 | 2_n12913;
assign 2_n4182 = 2_n5858 | 2_n11827;
assign 2_n2721 = 2_n5575 | 2_n12816;
assign 2_n8676 = 2_n4741 & 2_n4384;
assign 2_n4110 = 2_n11597 & 2_n9573;
assign 2_n7727 = ~(2_n392 ^ 2_n9940);
assign 2_n5723 = ~(2_n9553 ^ 2_n1771);
assign 2_n232 = 2_n5848 & 2_n3913;
assign 2_n3307 = ~(2_n10473 ^ 2_n10167);
assign 2_n2505 = 2_n11013 | 2_n1346;
assign 2_n6232 = ~(2_n6053 ^ 2_n2118);
assign 2_n11837 = ~(2_n10562 ^ 2_n8250);
assign 2_n8239 = ~(2_n1363 ^ 2_n6438);
assign 2_n8512 = 2_n1026 & 2_n11169;
assign 2_n2687 = 2_n183 | 2_n10638;
assign 2_n11826 = 2_n2832 | 2_n11746;
assign 2_n5669 = ~(2_n7029 ^ 2_n9249);
assign 2_n790 = ~2_n9038;
assign 2_n5508 = ~(2_n6384 | 2_n12233);
assign 2_n6785 = ~2_n6148;
assign 2_n12701 = 2_n6373 | 2_n4527;
assign 2_n1108 = ~(2_n12668 ^ 2_n10462);
assign 2_n10027 = ~2_n1440;
assign 2_n11233 = ~2_n7057;
assign 2_n6099 = ~(2_n3659 ^ 2_n11250);
assign 2_n12376 = 2_n8954 | 2_n10870;
assign 2_n1127 = ~(2_n4202 | 2_n9496);
assign 2_n10294 = ~2_n8868;
assign 2_n12081 = 2_n9106 & 2_n1488;
assign 2_n8086 = ~(2_n1024 ^ 2_n7498);
assign 2_n1 = 2_n2346 | 2_n6228;
assign 2_n8465 = ~(2_n8181 ^ 2_n8485);
assign 2_n10503 = ~(2_n6534 ^ 2_n10826);
assign 2_n7179 = ~(2_n2089 ^ 2_n2015);
assign 2_n10416 = ~(2_n2199 ^ 2_n10954);
assign 2_n11572 = ~(2_n3921 | 2_n3199);
assign 2_n2924 = 2_n8476 & 2_n6016;
assign 2_n9912 = ~(2_n5274 ^ 2_n2418);
assign 2_n10815 = ~(2_n4205 ^ 2_n8931);
assign 2_n4767 = 2_n8117 & 2_n745;
assign 2_n9213 = ~(2_n2144 | 2_n2392);
assign 2_n4208 = ~(2_n2479 ^ 2_n8144);
assign 2_n12107 = 2_n12186 | 2_n12816;
assign 2_n10516 = 2_n6577 | 2_n10919;
assign 2_n427 = 2_n4338 | 2_n10237;
assign 2_n11912 = ~(2_n10378 ^ 2_n7279);
assign 2_n8996 = 2_n12119 | 2_n3924;
assign 2_n5809 = ~2_n10545;
assign 2_n8738 = ~2_n3986;
assign 2_n8810 = 2_n5765 | 2_n4875;
assign 2_n5146 = 2_n3328 & 2_n10633;
assign 2_n3358 = 2_n10637 | 2_n3057;
assign 2_n9760 = ~(2_n8416 ^ 2_n5562);
assign 2_n12861 = ~(2_n7521 ^ 2_n4244);
assign 2_n7505 = 2_n12312 & 2_n7063;
assign 2_n84 = ~(2_n6535 ^ 2_n1482);
assign 2_n10077 = ~2_n3772;
assign 2_n1447 = 2_n4301 & 2_n2204;
assign 2_n12708 = 2_n5383 | 2_n10553;
assign 2_n3909 = 2_n11401 | 2_n2666;
assign 2_n578 = 2_n11539 & 2_n7445;
assign 2_n5976 = 2_n10095 & 2_n6546;
assign 2_n11046 = ~(2_n6064 | 2_n7069);
assign 2_n8748 = 2_n10365 | 2_n10723;
assign 2_n602 = 2_n752 | 2_n8414;
assign 2_n2019 = 2_n10162 & 2_n1558;
assign 2_n12189 = 2_n12503 | 2_n9568;
assign 2_n8013 = ~(2_n4373 ^ 2_n5628);
assign 2_n11331 = 2_n2473 | 2_n7782;
assign 2_n4652 = 2_n3072 & 2_n8111;
assign 2_n29 = ~(2_n7490 ^ 2_n10974);
assign 2_n4443 = 2_n8964 | 2_n5839;
assign 2_n6343 = ~(2_n3726 ^ 2_n277);
assign 2_n8902 = ~(2_n2962 | 2_n6955);
assign 2_n3625 = 2_n3743 | 2_n10916;
assign 2_n11490 = 2_n10835 | 2_n11698;
assign 2_n6104 = 2_n2656 | 2_n5536;
assign 2_n5671 = ~2_n11178;
assign 2_n648 = 2_n11712 | 2_n9574;
assign 2_n2674 = ~(2_n6041 | 2_n6923);
assign 2_n1738 = ~2_n9637;
assign 2_n4121 = 2_n2456 | 2_n5326;
assign 2_n8793 = 2_n3261 & 2_n11673;
assign 2_n7083 = ~(2_n5652 ^ 2_n12768);
assign 2_n720 = 2_n5452 & 2_n6117;
assign 2_n3317 = ~(2_n11250 | 2_n5379);
assign 2_n705 = 2_n2217 | 2_n7506;
assign 2_n5776 = ~(2_n8133 ^ 2_n10317);
assign 2_n3600 = 2_n2001 & 2_n8698;
assign 2_n10343 = 2_n5530 | 2_n12754;
assign 2_n2657 = 2_n6186 | 2_n4998;
assign 2_n7709 = ~2_n9457;
assign 2_n2418 = ~(2_n3314 ^ 2_n915);
assign 2_n4760 = 2_n4366 | 2_n10752;
assign 2_n7355 = ~(2_n361 ^ 2_n7728);
assign 2_n2981 = 2_n7283 | 2_n561;
assign 2_n12065 = 2_n4498 | 2_n1546;
assign 2_n609 = ~2_n5153;
assign 2_n6928 = ~2_n2141;
assign 2_n9666 = ~(2_n2608 ^ 2_n4615);
assign 2_n1935 = 2_n2893 & 2_n1014;
assign 2_n7835 = 2_n4808 & 2_n5388;
assign 2_n9580 = ~(2_n7311 | 2_n2344);
assign 2_n2919 = 2_n9058 & 2_n4197;
assign 2_n7203 = 2_n6270 | 2_n3877;
assign 2_n11112 = 2_n4059 | 2_n4400;
assign 2_n8051 = 2_n1685 | 2_n11030;
assign 2_n6774 = 2_n4674 | 2_n3224;
assign 2_n9416 = 2_n4702 & 2_n3750;
assign 2_n296 = 2_n12503 | 2_n3606;
assign 2_n8175 = 2_n6373 | 2_n9144;
assign 2_n1170 = ~(2_n895 | 2_n290);
assign 2_n12194 = 2_n7185 | 2_n2895;
assign 2_n10777 = 2_n4628 | 2_n10422;
assign 2_n9225 = ~2_n7976;
assign 2_n4495 = ~(2_n5650 ^ 2_n11675);
assign 2_n9707 = 2_n8241 & 2_n8962;
assign 2_n1997 = ~2_n12163;
assign 2_n11038 = 2_n9920 & 2_n3932;
assign 2_n3886 = 2_n8216 & 2_n10480;
assign 2_n12315 = 2_n12163 & 2_n8684;
assign 2_n5265 = 2_n9734 | 2_n900;
assign 2_n3141 = 2_n8026 | 2_n11820;
assign 2_n1058 = ~2_n2918;
assign 2_n459 = ~(2_n1495 ^ 2_n1506);
assign 2_n6540 = 2_n3310 | 2_n2706;
assign 2_n2923 = 2_n10434 | 2_n9894;
assign 2_n5210 = ~2_n7499;
assign 2_n9904 = ~(2_n5690 ^ 2_n1607);
assign 2_n12565 = ~(2_n6356 | 2_n9270);
assign 2_n3044 = ~(2_n9398 ^ 2_n446);
assign 2_n1159 = ~(2_n2583 ^ 2_n954);
assign 2_n6643 = 2_n8428 | 2_n10919;
assign 2_n4483 = 2_n4628 | 2_n8740;
assign 2_n9262 = ~2_n4722;
assign 2_n4861 = ~(2_n6283 ^ 2_n5838);
assign 2_n6242 = 2_n8552 | 2_n12735;
assign 2_n550 = 2_n8428 | 2_n6084;
assign 2_n920 = 2_n2056 & 2_n10008;
assign 2_n4430 = ~(2_n9267 ^ 2_n9044);
assign 2_n12750 = 2_n8070 | 2_n473;
assign 2_n8415 = 2_n8920 & 2_n8547;
assign 2_n8323 = 2_n936 | 2_n5520;
assign 2_n9300 = ~(2_n4852 ^ 2_n7868);
assign 2_n50 = 2_n9389 | 2_n4775;
assign 2_n9137 = ~(2_n12081 ^ 2_n153);
assign 2_n6514 = 2_n962 | 2_n9144;
assign 2_n10006 = ~(2_n4084 | 2_n2120);
assign 2_n2976 = 2_n10142 | 2_n1079;
assign 2_n12063 = 2_n2838 | 2_n6164;
assign 2_n11240 = ~(2_n9647 | 2_n11633);
assign 2_n10832 = 2_n8458 | 2_n3761;
assign 2_n1635 = ~(2_n7275 | 2_n3788);
assign 2_n2718 = ~2_n1548;
assign 2_n2047 = 2_n5082 & 2_n8365;
assign 2_n11285 = 2_n8959 | 2_n6455;
assign 2_n3425 = ~2_n8776;
assign 2_n3889 = ~(2_n11507 | 2_n3685);
assign 2_n12121 = 2_n6940 | 2_n7615;
assign 2_n6387 = ~(2_n12703 ^ 2_n8033);
assign 2_n3489 = ~2_n5078;
assign 2_n5744 = 2_n6377 & 2_n12854;
assign 2_n1572 = ~(2_n7824 | 2_n12880);
assign 2_n2338 = 2_n8687 | 2_n4654;
assign 2_n4490 = 2_n1839 & 2_n4585;
assign 2_n10015 = ~(2_n12556 ^ 2_n997);
assign 2_n4381 = ~2_n11189;
assign 2_n8990 = ~(2_n820 ^ 2_n12499);
assign 2_n3866 = 2_n3414 | 2_n5170;
assign 2_n218 = ~(2_n4112 ^ 2_n2282);
assign 2_n8209 = ~(2_n4766 | 2_n9346);
assign 2_n12412 = ~(2_n9081 ^ 2_n3026);
assign 2_n5050 = 2_n10211 | 2_n8355;
assign 2_n3089 = ~(2_n2197 ^ 2_n2281);
assign 2_n694 = 2_n2191 & 2_n3550;
assign 2_n1205 = 2_n8959 | 2_n2815;
assign 2_n9274 = 2_n10835 | 2_n5914;
assign 2_n8811 = ~(2_n11149 ^ 2_n7385);
assign 2_n12255 = ~(2_n12550 ^ 2_n9946);
assign 2_n10035 = 2_n2639 | 2_n6420;
assign 2_n8817 = ~2_n5059;
assign 2_n12544 = ~(2_n2271 | 2_n2399);
assign 2_n6867 = 2_n6776 & 2_n10439;
assign 2_n2401 = 2_n989 | 2_n9589;
assign 2_n2511 = 2_n6740 | 2_n9524;
assign 2_n2852 = 2_n12853 | 2_n10422;
assign 2_n4667 = 2_n6570 | 2_n11756;
assign 2_n5867 = ~2_n11840;
assign 2_n6451 = 2_n8959 | 2_n5540;
assign 2_n3116 = 2_n5530 | 2_n7136;
assign 2_n538 = ~(2_n5386 ^ 2_n12572);
assign 2_n1868 = 2_n12423 & 2_n7303;
assign 2_n8756 = ~2_n8784;
assign 2_n2116 = 2_n8959 | 2_n7425;
assign 2_n3441 = 2_n3746 | 2_n6084;
assign 2_n8331 = ~(2_n7 ^ 2_n4663);
assign 2_n4783 = 2_n3242 & 2_n6957;
assign 2_n2889 = ~(2_n8551 ^ 2_n12230);
assign 2_n12439 = ~2_n10841;
assign 2_n11360 = ~(2_n12040 ^ 2_n11349);
assign 2_n717 = 2_n9077 & 2_n5332;
assign 2_n11692 = ~(2_n758 | 2_n2826);
assign 2_n882 = 2_n3617 | 2_n12535;
assign 2_n3874 = 2_n11653 | 2_n4524;
assign 2_n10031 = ~(2_n6037 ^ 2_n5347);
assign 2_n8758 = 2_n5355 | 2_n9589;
assign 2_n9516 = ~(2_n7602 ^ 2_n1841);
assign 2_n3008 = ~(2_n7115 ^ 2_n2330);
assign 2_n11506 = ~(2_n11460 | 2_n12888);
assign 2_n11962 = 2_n8220 | 2_n7838;
assign 2_n12222 = ~(2_n3579 ^ 2_n8300);
assign 2_n5163 = ~(2_n11013 ^ 2_n2022);
assign 2_n3500 = ~(2_n8149 ^ 2_n109);
assign 2_n6027 = 2_n660 | 2_n2927;
assign 2_n7856 = ~2_n953;
assign 2_n7918 = ~(2_n9606 | 2_n679);
assign 2_n9131 = ~(2_n666 ^ 2_n10519);
assign 2_n4492 = 2_n7854 & 2_n4952;
assign 2_n596 = ~(2_n5881 | 2_n10150);
assign 2_n8556 = 2_n2393 & 2_n7294;
assign 2_n12478 = ~2_n2476;
assign 2_n5176 = ~(2_n5660 ^ 2_n6107);
assign 2_n1221 = ~(2_n5898 ^ 2_n3139);
assign 2_n702 = ~(2_n8458 ^ 2_n3761);
assign 2_n6796 = 2_n5369 | 2_n4259;
assign 2_n7299 = ~(2_n1864 ^ 2_n10145);
assign 2_n5171 = ~(2_n3910 | 2_n6548);
assign 2_n11308 = ~(2_n8914 ^ 2_n11802);
assign 2_n1705 = 2_n5355 | 2_n7424;
assign 2_n1426 = 2_n1848 & 2_n1374;
assign 2_n3372 = ~(2_n5635 ^ 2_n4056);
assign 2_n10723 = ~(2_n10448 ^ 2_n6747);
assign 2_n10668 = 2_n6681 & 2_n10894;
assign 2_n10933 = 2_n7765 & 2_n4208;
assign 2_n1751 = ~(2_n2459 ^ 2_n4594);
assign 2_n7499 = 2_n9389 | 2_n2358;
assign 2_n6988 = 2_n5283 & 2_n7610;
assign 2_n12229 = ~2_n12241;
assign 2_n8871 = 2_n8429 | 2_n10376;
assign 2_n5404 = 2_n8187 | 2_n7881;
assign 2_n9957 = ~(2_n11659 | 2_n11408);
assign 2_n11605 = 2_n5765 | 2_n6922;
assign 2_n12211 = ~2_n7850;
assign 2_n8330 = ~2_n10689;
assign 2_n9120 = 2_n9702 | 2_n4844;
assign 2_n5352 = ~(2_n12539 ^ 2_n10409);
assign 2_n9325 = 2_n2133 | 2_n11530;
assign 2_n767 = ~2_n9882;
assign 2_n2653 = ~2_n10686;
assign 2_n10840 = 2_n8870 | 2_n5468;
assign 2_n9279 = ~2_n7668;
assign 2_n5518 = ~2_n721;
assign 2_n1476 = ~2_n6611;
assign 2_n7903 = 2_n5366 | 2_n5004;
assign 2_n8640 = 2_n5108 ^ 2_n8939;
assign 2_n7111 = 2_n6373 | 2_n4654;
assign 2_n4324 = 2_n6098 | 2_n1845;
assign 2_n11613 = 2_n3820 | 2_n1047;
assign 2_n8207 = 2_n9687 & 2_n11344;
assign 2_n5443 = ~(2_n7012 ^ 2_n3834);
assign 2_n6510 = ~2_n7929;
assign 2_n9239 = 2_n7268 | 2_n1767;
assign 2_n10942 = ~2_n10214;
assign 2_n282 = 2_n9389 | 2_n6389;
assign 2_n4207 = ~2_n11323;
assign 2_n1977 = ~(2_n10834 ^ 2_n6624);
assign 2_n8562 = ~(2_n9404 ^ 2_n9679);
assign 2_n8655 = ~2_n4826;
assign 2_n10484 = ~(2_n7284 ^ 2_n365);
assign 2_n10881 = 2_n11998 | 2_n11648;
assign 2_n2888 = ~(2_n4023 ^ 2_n7696);
assign 2_n6073 = 2_n10142 | 2_n4242;
assign 2_n5657 = ~(2_n8117 | 2_n745);
assign 2_n5906 = ~(2_n9627 ^ 2_n833);
assign 2_n5525 = 2_n7391 | 2_n3911;
assign 2_n11199 = ~2_n7370;
assign 2_n11776 = ~(2_n11754 ^ 2_n3814);
assign 2_n7890 = 2_n10531 & 2_n1467;
assign 2_n4995 = 2_n10065 | 2_n198;
assign 2_n9788 = ~(2_n7666 ^ 2_n11010);
assign 2_n10576 = 2_n5495 | 2_n10986;
assign 2_n11640 = ~(2_n12500 ^ 2_n2829);
assign 2_n10623 = ~2_n5408;
assign 2_n11693 = ~(2_n5059 ^ 2_n4099);
assign 2_n2390 = 2_n1064 | 2_n4813;
assign 2_n1030 = ~(2_n3381 ^ 2_n10811);
assign 2_n5470 = ~(2_n120 | 2_n65);
assign 2_n487 = ~(2_n12939 | 2_n6858);
assign 2_n443 = 2_n6368 | 2_n1309;
assign 2_n6721 = ~(2_n7680 | 2_n8662);
assign 2_n12003 = ~(2_n822 ^ 2_n7162);
assign 2_n8905 = 2_n12237 | 2_n12735;
assign 2_n11500 = 2_n2997 & 2_n6848;
assign 2_n8145 = 2_n9373 | 2_n7506;
assign 2_n7735 = 2_n5331 & 2_n1512;
assign 2_n6218 = 2_n8011 | 2_n4866;
assign 2_n9843 = 2_n8310 | 2_n2912;
assign 2_n3155 = 2_n357 | 2_n5306;
assign 2_n395 = ~(2_n7635 ^ 2_n10300);
assign 2_n1799 = ~2_n4914;
assign 2_n1182 = 2_n62 | 2_n377;
assign 2_n12673 = 2_n5361 | 2_n6282;
assign 2_n12137 = ~(2_n10514 | 2_n11187);
assign 2_n12434 = ~(2_n4779 | 2_n4890);
assign 2_n7122 = ~(2_n7622 ^ 2_n10067);
assign 2_n4253 = ~(2_n7675 ^ 2_n6828);
assign 2_n2941 = 2_n3962 & 2_n4463;
assign 2_n780 = ~(2_n5707 ^ 2_n9944);
assign 2_n6161 = 2_n989 | 2_n2076;
assign 2_n3827 = ~(2_n6882 ^ 2_n6622);
assign 2_n10055 = ~2_n6773;
assign 2_n11870 = ~(2_n6660 ^ 2_n7096);
assign 2_n3402 = ~(2_n2443 | 2_n3859);
assign 2_n142 = 2_n5621 & 2_n4075;
assign 2_n6413 = 2_n12133 & 2_n6866;
assign 2_n4256 = 2_n5893 & 2_n6088;
assign 2_n5565 = ~(2_n1046 ^ 2_n3683);
assign 2_n919 = ~2_n11336;
assign 2_n5278 = 2_n5527 & 2_n1217;
assign 2_n11518 = 2_n8273 | 2_n4909;
assign 2_n526 = ~2_n4292;
assign 2_n9570 = 2_n989 | 2_n1915;
assign 2_n261 = ~2_n8035;
assign 2_n7531 = ~(2_n7614 ^ 2_n471);
assign 2_n8674 = 2_n10157 | 2_n10916;
assign 2_n2500 = 2_n4870 & 2_n500;
assign 2_n5030 = ~(2_n4323 ^ 2_n7426);
assign 2_n11187 = 2_n2520 & 2_n1745;
assign 2_n10235 = ~(2_n8596 | 2_n3584);
assign 2_n3086 = ~(2_n720 ^ 2_n12516);
assign 2_n2343 = ~(2_n11396 ^ 2_n4847);
assign 2_n6630 = ~2_n6059;
assign 2_n11789 = ~(2_n1461 ^ 2_n7491);
assign 2_n2865 = ~(2_n5715 | 2_n7720);
assign 2_n2607 = 2_n1469 | 2_n10489;
assign 2_n4777 = 2_n3743 | 2_n5258;
assign 2_n8112 = 2_n966 | 2_n11943;
assign 2_n5982 = 2_n8870 | 2_n826;
assign 2_n54 = 2_n12361 | 2_n6084;
assign 2_n12898 = ~(2_n4511 | 2_n8863);
assign 2_n11224 = ~(2_n8267 ^ 2_n11939);
assign 2_n6991 = ~2_n12215;
assign 2_n11370 = 2_n989 | 2_n3911;
assign 2_n12858 = 2_n3743 | 2_n609;
assign 2_n9115 = ~(2_n4289 ^ 2_n3035);
assign 2_n9941 = ~(2_n601 ^ 2_n3269);
assign 2_n1884 = ~(2_n577 ^ 2_n8482);
assign 2_n12560 = 2_n4263 & 2_n8131;
assign 2_n9539 = ~(2_n8293 ^ 2_n12519);
assign 2_n7996 = 2_n962 | 2_n4654;
assign 2_n6029 = 2_n12443 & 2_n1734;
assign 2_n7564 = 2_n10142 | 2_n12328;
assign 2_n7186 = ~2_n3313;
assign 2_n5082 = 2_n173 & 2_n3686;
assign 2_n1034 = ~(2_n10031 ^ 2_n5467);
assign 2_n5532 = 2_n8687 | 2_n2020;
assign 2_n12235 = ~2_n3991;
assign 2_n2282 = 2_n11923 | 2_n12771;
assign 2_n8848 = 2_n10196 | 2_n2020;
assign 2_n12913 = 2_n4911 | 2_n10066;
assign 2_n10517 = 2_n11311 & 2_n2522;
assign 2_n530 = ~2_n4970;
assign 2_n3432 = ~(2_n2033 ^ 2_n8014);
assign 2_n3593 = 2_n7358 & 2_n466;
assign 2_n4542 = ~(2_n4298 ^ 2_n1001);
assign 2_n2722 = 2_n12423 | 2_n7303;
assign 2_n6243 = 2_n1415 & 2_n4630;
assign 2_n7138 = ~2_n6121;
assign 2_n1346 = ~(2_n4449 ^ 2_n4391);
assign 2_n6860 = ~(2_n12693 ^ 2_n10616);
assign 2_n5172 = 2_n3533 & 2_n5660;
assign 2_n8031 = ~2_n4417;
assign 2_n1697 = 2_n5855 & 2_n3487;
assign 2_n3474 = 2_n114 | 2_n7876;
assign 2_n4267 = ~2_n3807;
assign 2_n3487 = 2_n11051 | 2_n9731;
assign 2_n2524 = 2_n3611 | 2_n11027;
assign 2_n7242 = ~(2_n3305 ^ 2_n6890);
assign 2_n8399 = ~(2_n10873 ^ 2_n1950);
assign 2_n6509 = 2_n8480 | 2_n5865;
assign 2_n11565 = ~(2_n4442 ^ 2_n11248);
assign 2_n1157 = 2_n1941 | 2_n6455;
assign 2_n10878 = 2_n5363 & 2_n3006;
assign 2_n8605 = ~(2_n10814 ^ 2_n7368);
assign 2_n8423 = 2_n11958 | 2_n6197;
assign 2_n4045 = 2_n8557 & 2_n7653;
assign 2_n3641 = ~(2_n2061 ^ 2_n1158);
assign 2_n2855 = ~(2_n4755 ^ 2_n11338);
assign 2_n8615 = ~2_n9737;
assign 2_n10464 = ~2_n9326;
assign 2_n6653 = ~(2_n7480 ^ 2_n1080);
assign 2_n8044 = ~(2_n12526 ^ 2_n5750);
assign 2_n2858 = 2_n6298 | 2_n6721;
assign 2_n10872 = 2_n6077 & 2_n11715;
assign 2_n6111 = 2_n3106 & 2_n11945;
assign 2_n2803 = ~(2_n2284 ^ 2_n11102);
assign 2_n7220 = ~(2_n4431 | 2_n6243);
assign 2_n11026 = ~2_n2393;
assign 2_n2961 = ~(2_n5204 ^ 2_n283);
assign 2_n9804 = ~(2_n11782 ^ 2_n5114);
assign 2_n12218 = ~2_n12747;
assign 2_n7558 = ~2_n2522;
assign 2_n11425 = 2_n2217 | 2_n5258;
assign 2_n4614 = ~(2_n8503 | 2_n3889);
assign 2_n5733 = ~(2_n10452 ^ 2_n10676);
assign 2_n11192 = 2_n962 | 2_n9160;
assign 2_n9133 = ~(2_n11945 ^ 2_n6487);
assign 2_n8714 = ~2_n4603;
assign 2_n2931 = ~2_n7490;
assign 2_n7693 = ~(2_n129 ^ 2_n9330);
assign 2_n9702 = 2_n2195 & 2_n1101;
assign 2_n6525 = ~(2_n391 | 2_n1821);
assign 2_n10914 = ~(2_n1644 ^ 2_n11612);
assign 2_n9183 = ~(2_n5503 | 2_n730);
assign 2_n7970 = ~2_n9727;
assign 2_n679 = ~2_n7647;
assign 2_n8333 = ~(2_n4866 ^ 2_n8252);
assign 2_n7739 = ~2_n11575;
assign 2_n4880 = ~(2_n12305 ^ 2_n3223);
assign 2_n3700 = 2_n1872 | 2_n3556;
assign 2_n11352 = 2_n5575 | 2_n7876;
assign 2_n6235 = 2_n4053 | 2_n10130;
assign 2_n1578 = ~(2_n1879 | 2_n142);
assign 2_n358 = 2_n8959 | 2_n2232;
assign 2_n7090 = ~2_n12790;
assign 2_n2625 = 2_n10157 | 2_n609;
assign 2_n1032 = ~(2_n4690 ^ 2_n8965);
assign 2_n3163 = 2_n7432 & 2_n5058;
assign 2_n11300 = ~(2_n9557 ^ 2_n4574);
assign 2_n3692 = 2_n11475 & 2_n7800;
assign 2_n3463 = ~(2_n737 | 2_n6132);
assign 2_n7734 = 2_n1172 & 2_n3669;
assign 2_n3818 = ~2_n9508;
assign 2_n8360 = ~(2_n11588 ^ 2_n9112);
assign 2_n5389 = ~2_n1062;
assign 2_n9050 = 2_n11542 & 2_n6333;
assign 2_n7755 = ~2_n8533;
assign 2_n5010 = 2_n10594 & 2_n6540;
assign 2_n1158 = ~(2_n7297 ^ 2_n7935);
assign 2_n6224 = 2_n10108 | 2_n12843;
assign 2_n12659 = 2_n3743 | 2_n5502;
assign 2_n8215 = 2_n11753 | 2_n3341;
assign 2_n2204 = 2_n11719 | 2_n11827;
assign 2_n7321 = 2_n8430 & 2_n1452;
assign 2_n1148 = ~2_n8460;
assign 2_n7967 = 2_n12023 | 2_n7734;
assign 2_n3857 = ~(2_n2881 | 2_n7744);
assign 2_n4799 = 2_n6437 & 2_n12847;
assign 2_n5587 = ~(2_n1355 ^ 2_n7273);
assign 2_n5944 = 2_n6718 | 2_n4864;
assign 2_n345 = ~(2_n6931 ^ 2_n1197);
assign 2_n9058 = 2_n2427 | 2_n1157;
assign 2_n9248 = 2_n7586 | 2_n1505;
assign 2_n211 = ~2_n3536;
assign 2_n11414 = ~(2_n1784 ^ 2_n11686);
assign 2_n3611 = ~(2_n7856 ^ 2_n2798);
assign 2_n1393 = 2_n7381 | 2_n865;
assign 2_n12806 = ~(2_n320 ^ 2_n12447);
assign 2_n7917 = ~(2_n11360 ^ 2_n2803);
assign 2_n1338 = 2_n2101 & 2_n3422;
assign 2_n11056 = ~(2_n5269 | 2_n12488);
assign 2_n1066 = 2_n8450 | 2_n10025;
assign 2_n1843 = ~2_n7652;
assign 2_n5445 = 2_n664 & 2_n9991;
assign 2_n6312 = 2_n1699 | 2_n4913;
assign 2_n9884 = 2_n994 | 2_n7703;
assign 2_n3145 = 2_n5575 | 2_n995;
assign 2_n126 = ~2_n5789;
assign 2_n3139 = ~(2_n849 ^ 2_n329);
assign 2_n12908 = ~(2_n3265 ^ 2_n1454);
assign 2_n11592 = 2_n5393 | 2_n6733;
assign 2_n8609 = ~(2_n10516 ^ 2_n778);
assign 2_n5485 = 2_n11026 | 2_n4527;
assign 2_n11264 = ~(2_n2673 ^ 2_n2648);
assign 2_n8278 = ~(2_n9616 ^ 2_n5262);
assign 2_n6030 = 2_n3544 | 2_n4715;
assign 2_n6852 = ~2_n7419;
assign 2_n12318 = 2_n5575 | 2_n184;
assign 2_n5619 = 2_n6171 | 2_n7351;
assign 2_n9654 = ~(2_n3921 ^ 2_n429);
assign 2_n4344 = ~(2_n2503 ^ 2_n5908);
assign 2_n2264 = ~(2_n8023 ^ 2_n9300);
assign 2_n11761 = ~(2_n2162 | 2_n7307);
assign 2_n2079 = ~2_n11633;
assign 2_n4882 = 2_n4791 & 2_n5762;
assign 2_n2386 = ~2_n10923;
assign 2_n3130 = 2_n3820 | 2_n4654;
assign 2_n147 = 2_n12648 & 2_n2802;
assign 2_n7700 = ~(2_n10958 ^ 2_n540);
assign 2_n6982 = 2_n12144 & 2_n5251;
assign 2_n5290 = ~(2_n2309 | 2_n3798);
assign 2_n7621 = ~(2_n10992 ^ 2_n14);
assign 2_n9840 = ~(2_n248 ^ 2_n11837);
assign 2_n6200 = ~2_n10457;
assign 2_n1160 = ~2_n822;
assign 2_n5705 = ~(2_n9481 ^ 2_n12507);
assign 2_n63 = ~(2_n12095 | 2_n1578);
assign 2_n6428 = ~(2_n5989 ^ 2_n3457);
assign 2_n3674 = ~2_n10877;
assign 2_n11762 = 2_n7329 | 2_n8461;
assign 2_n9016 = 2_n12119 | 2_n8109;
assign 2_n606 = ~(2_n6121 ^ 2_n2158);
assign 2_n1420 = ~(2_n7278 ^ 2_n598);
assign 2_n8611 = ~2_n12628;
assign 2_n1374 = 2_n8019 | 2_n9631;
assign 2_n12497 = 2_n209 | 2_n4050;
assign 2_n3773 = 2_n10309 & 2_n11180;
assign 2_n9504 = 2_n5530 | 2_n8655;
assign 2_n7960 = 2_n810 & 2_n2058;
assign 2_n4983 = ~2_n7612;
assign 2_n2966 = 2_n11892 & 2_n806;
assign 2_n1178 = 2_n4097 & 2_n11394;
assign 2_n9830 = 2_n6478 & 2_n3855;
assign 2_n4112 = 2_n5765 | 2_n9568;
assign 2_n10091 = 2_n7116 | 2_n11820;
assign 2_n1905 = ~(2_n2858 ^ 2_n5772);
assign 2_n1277 = ~2_n2784;
assign 2_n10861 = ~(2_n12715 ^ 2_n11494);
assign 2_n9751 = ~2_n5688;
assign 2_n5502 = ~2_n159;
assign 2_n257 = 2_n11594 | 2_n272;
assign 2_n10688 = 2_n5700 | 2_n2958;
assign 2_n2412 = ~2_n628;
assign 2_n614 = 2_n573 | 2_n11044;
assign 2_n10802 = 2_n5479 & 2_n8519;
assign 2_n1860 = ~(2_n8070 ^ 2_n473);
assign 2_n6767 = ~(2_n8774 ^ 2_n3152);
assign 2_n6705 = ~(2_n10407 ^ 2_n2755);
assign 2_n10864 = ~(2_n11734 | 2_n6862);
assign 2_n11251 = ~2_n9007;
assign 2_n12279 = ~(2_n5361 ^ 2_n12729);
assign 2_n5507 = ~2_n904;
assign 2_n5658 = 2_n10157 | 2_n9160;
assign 2_n1039 = 2_n1518 & 2_n211;
assign 2_n5718 = 2_n7391 | 2_n6389;
assign 2_n11279 = ~(2_n12782 ^ 2_n2379);
assign 2_n1707 = ~(2_n6536 ^ 2_n6532);
assign 2_n2999 = 2_n255 & 2_n4288;
assign 2_n1123 = 2_n752 | 2_n9971;
assign 2_n9256 = 2_n3348 | 2_n67;
assign 2_n8881 = 2_n5620 | 2_n9864;
assign 2_n11032 = ~(2_n2574 | 2_n1190);
assign 2_n4545 = 2_n4214 & 2_n7650;
assign 2_n7879 = 2_n8452 & 2_n8978;
assign 2_n4448 = ~2_n3914;
assign 2_n962 = ~2_n1471;
assign 2_n4454 = ~(2_n5856 ^ 2_n10890);
assign 2_n2288 = 2_n4112 | 2_n2282;
assign 2_n11134 = ~(2_n5554 ^ 2_n12161);
assign 2_n4873 = ~2_n12939;
assign 2_n9299 = 2_n3160 | 2_n1116;
assign 2_n5090 = ~(2_n8103 ^ 2_n5741);
assign 2_n2601 = ~(2_n3235 | 2_n407);
assign 2_n6214 = 2_n11413 | 2_n937;
assign 2_n1037 = ~(2_n6987 ^ 2_n3200);
assign 2_n6521 = 2_n5195 & 2_n4478;
assign 2_n4766 = ~2_n10117;
assign 2_n4331 = 2_n9185 & 2_n3250;
assign 2_n1036 = 2_n8453 & 2_n4625;
assign 2_n343 = ~(2_n11119 ^ 2_n7274);
assign 2_n942 = 2_n1947 & 2_n11587;
assign 2_n7245 = 2_n11073 & 2_n5965;
assign 2_n11323 = ~(2_n10096 ^ 2_n4208);
assign 2_n2100 = 2_n9878 | 2_n4913;
assign 2_n7604 = 2_n6854 | 2_n2439;
assign 2_n10050 = 2_n612 | 2_n9775;
assign 2_n10521 = 2_n10242 & 2_n12660;
assign 2_n6937 = ~(2_n1483 ^ 2_n5676);
assign 2_n1131 = 2_n2456 | 2_n7928;
assign 2_n800 = 2_n3361 | 2_n1243;
assign 2_n6610 = ~(2_n12739 ^ 2_n6652);
assign 2_n11823 = ~2_n4435;
assign 2_n12018 = ~(2_n9899 | 2_n3737);
assign 2_n9127 = ~(2_n10738 ^ 2_n6451);
assign 2_n3686 = ~2_n11498;
assign 2_n10817 = 2_n12622 & 2_n3919;
assign 2_n9744 = 2_n191 | 2_n8859;
assign 2_n5567 = ~2_n2376;
assign 2_n12147 = ~2_n10918;
assign 2_n2190 = 2_n6977 | 2_n6084;
assign 2_n2823 = ~2_n1210;
assign 2_n4374 = ~(2_n6557 ^ 2_n11804);
assign 2_n7793 = ~(2_n8872 ^ 2_n11270);
assign 2_n2025 = ~(2_n3372 | 2_n6124);
assign 2_n2929 = ~(2_n3633 ^ 2_n3825);
assign 2_n5289 = 2_n9448 | 2_n4181;
assign 2_n9848 = ~(2_n11727 ^ 2_n1119);
assign 2_n7055 = ~(2_n9342 | 2_n11970);
assign 2_n5477 = 2_n5252 | 2_n3309;
assign 2_n10750 = ~2_n12391;
assign 2_n68 = ~(2_n7016 ^ 2_n11437);
assign 2_n11845 = ~(2_n656 | 2_n10580);
assign 2_n5478 = ~(2_n5243 ^ 2_n11640);
assign 2_n7511 = 2_n8549 & 2_n2493;
assign 2_n11743 = 2_n9054 | 2_n10082;
assign 2_n9855 = ~(2_n2859 ^ 2_n2949);
assign 2_n11689 = 2_n9370 | 2_n5497;
assign 2_n4375 = 2_n2254 & 2_n10227;
assign 2_n7211 = ~(2_n4759 ^ 2_n929);
assign 2_n9871 = 2_n11923 | 2_n9280;
assign 2_n1973 = 2_n11958 | 2_n2232;
assign 2_n3377 = 2_n591 | 2_n11790;
assign 2_n6315 = ~(2_n95 ^ 2_n5882);
assign 2_n6809 = ~(2_n6700 ^ 2_n6120);
assign 2_n3779 = ~(2_n6212 ^ 2_n10328);
assign 2_n1362 = 2_n12721 & 2_n6196;
assign 2_n12931 = ~(2_n8294 | 2_n6316);
assign 2_n6897 = 2_n3628 & 2_n894;
assign 2_n12430 = ~(2_n4613 | 2_n4098);
assign 2_n10468 = ~2_n9608;
assign 2_n2942 = ~(2_n8816 ^ 2_n1217);
assign 2_n5189 = 2_n8928 ^ 2_n2974;
assign 2_n3544 = 2_n11958 | 2_n3421;
assign 2_n11486 = ~(2_n9161 | 2_n2531);
assign 2_n6665 = 2_n3998 & 2_n608;
assign 2_n1211 = ~(2_n2598 ^ 2_n265);
assign 2_n3329 = ~(2_n6782 | 2_n7054);
assign 2_n567 = ~(2_n3141 ^ 2_n4721);
assign 2_n10232 = ~(2_n6738 ^ 2_n252);
assign 2_n4458 = 2_n12853 | 2_n6513;
assign 2_n3385 = ~(2_n5621 ^ 2_n1879);
assign 2_n4700 = 2_n2923 & 2_n7999;
assign 2_n8641 = 2_n1642 | 2_n12325;
assign 2_n2958 = ~(2_n5863 ^ 2_n3149);
assign 2_n11477 = 2_n12758 & 2_n7584;
assign 2_n7811 = ~(2_n6750 ^ 2_n3701);
assign 2_n5727 = ~2_n3815;
assign 2_n7443 = ~2_n6364;
assign 2_n7052 = 2_n9007 | 2_n7956;
assign 2_n8140 = 2_n9105 & 2_n1981;
assign 2_n12573 = 2_n7128 & 2_n6684;
assign 2_n4359 = ~(2_n12117 | 2_n143);
assign 2_n274 = 2_n9453 & 2_n9646;
assign 2_n5180 = 2_n7694 & 2_n12015;
assign 2_n4460 = 2_n1699 | 2_n12535;
assign 2_n3108 = 2_n807 | 2_n6455;
assign 2_n7366 = ~(2_n10619 ^ 2_n11819);
assign 2_n9833 = 2_n3105 & 2_n358;
assign 2_n5699 = ~2_n7997;
assign 2_n239 = ~2_n8864;
assign 2_n6488 = ~(2_n5080 ^ 2_n7917);
assign 2_n6912 = ~(2_n11677 ^ 2_n1025);
assign 2_n697 = 2_n8552 | 2_n9188;
assign 2_n2107 = ~2_n1113;
assign 2_n8221 = 2_n12853 | 2_n1932;
assign 2_n8970 = ~2_n11536;
assign 2_n344 = 2_n204 & 2_n6608;
assign 2_n4428 = 2_n3110 & 2_n4940;
assign 2_n3211 = 2_n10791 & 2_n8508;
assign 2_n4602 = 2_n8858 & 2_n4452;
assign 2_n347 = 2_n5685 | 2_n5658;
assign 2_n3513 = 2_n5950 & 2_n5359;
assign 2_n10248 = ~2_n4181;
assign 2_n1486 = ~2_n3326;
assign 2_n9066 = 2_n7468 | 2_n271;
assign 2_n10093 = ~(2_n6085 | 2_n12029);
assign 2_n2933 = 2_n9878 | 2_n826;
assign 2_n4175 = 2_n1024 & 2_n7498;
assign 2_n1482 = ~(2_n7621 ^ 2_n8614);
assign 2_n5937 = ~2_n11136;
assign 2_n12780 = 2_n1089 & 2_n10310;
assign 2_n4016 = 2_n6637 | 2_n461;
assign 2_n11673 = 2_n6739 | 2_n9109;
assign 2_n10846 = 2_n7283 | 2_n1851;
assign 2_n2622 = ~(2_n9290 ^ 2_n6049);
assign 2_n2437 = ~2_n6539;
assign 2_n8410 = 2_n8702 | 2_n8911;
assign 2_n2357 = 2_n2176 & 2_n8516;
assign 2_n1416 = 2_n5158 & 2_n7751;
assign 2_n6122 = 2_n6577 | 2_n6084;
assign 2_n5563 = ~(2_n6447 ^ 2_n11891);
assign 2_n7927 = 2_n5671 | 2_n1134;
assign 2_n10607 = ~2_n8445;
assign 2_n9180 = 2_n3611 & 2_n11027;
assign 2_n9285 = 2_n10148 & 2_n7996;
assign 2_n4649 = ~(2_n7493 | 2_n8551);
assign 2_n10069 = ~(2_n6470 ^ 2_n7392);
assign 2_n5221 = ~(2_n4981 ^ 2_n12209);
assign 2_n1334 = 2_n4059 | 2_n510;
assign 2_n4843 = ~2_n11388;
assign 2_n10130 = 2_n8996 & 2_n9518;
assign 2_n5825 = ~(2_n12545 ^ 2_n1180);
assign 2_n9008 = ~(2_n10225 | 2_n3598);
assign 2_n10422 = ~2_n2551;
assign 2_n10213 = ~(2_n11205 ^ 2_n11622);
assign 2_n8094 = 2_n6439 | 2_n6447;
assign 2_n3530 = ~2_n3170;
assign 2_n9371 = ~(2_n7380 ^ 2_n11427);
assign 2_n1668 = 2_n3740 | 2_n10116;
assign 2_n9951 = ~(2_n8879 | 2_n7199);
assign 2_n7647 = 2_n5330 & 2_n1401;
assign 2_n3941 = 2_n11709 & 2_n831;
assign 2_n3926 = 2_n11181 | 2_n4268;
assign 2_n9503 = ~(2_n10598 | 2_n2601);
assign 2_n11239 = 2_n1409 & 2_n12780;
assign 2_n5557 = ~(2_n1629 ^ 2_n5509);
assign 2_n98 = ~(2_n7910 ^ 2_n8706);
assign 2_n6674 = ~2_n4746;
assign 2_n6952 = 2_n10142 | 2_n6524;
assign 2_n8781 = ~(2_n1341 | 2_n9522);
assign 2_n2194 = ~(2_n7433 | 2_n1884);
assign 2_n4424 = 2_n6718 | 2_n9280;
assign 2_n9247 = ~2_n10742;
assign 2_n9558 = ~(2_n12723 ^ 2_n1584);
assign 2_n11674 = 2_n7449 | 2_n4875;
assign 2_n803 = ~(2_n3925 | 2_n4797);
assign 2_n10158 = ~(2_n11844 | 2_n6991);
assign 2_n11577 = 2_n8276 & 2_n2024;
assign 2_n5927 = ~(2_n12227 ^ 2_n11940);
assign 2_n1950 = ~(2_n1530 ^ 2_n1115);
assign 2_n337 = 2_n4628 | 2_n7382;
assign 2_n8335 = 2_n12579 & 2_n6506;
assign 2_n9993 = 2_n7231 & 2_n6505;
assign 2_n11935 = 2_n11923 | 2_n7506;
assign 2_n9069 = ~(2_n9848 ^ 2_n2568);
assign 2_n2520 = 2_n2730 | 2_n3094;
assign 2_n2490 = 2_n4343 | 2_n9188;
assign 2_n5155 = ~(2_n7318 ^ 2_n8993);
assign 2_n1525 = 2_n9369 & 2_n2952;
assign 2_n12734 = 2_n6577 | 2_n7558;
assign 2_n2660 = 2_n6181 | 2_n10334;
assign 2_n744 = ~(2_n9353 ^ 2_n9243);
assign 2_n11098 = 2_n961 & 2_n9553;
assign 2_n7019 = 2_n6373 | 2_n5502;
assign 2_n1772 = ~(2_n9735 | 2_n12481);
assign 2_n325 = 2_n10196 | 2_n4527;
assign 2_n8764 = 2_n9277 | 2_n9473;
assign 2_n11075 = ~(2_n11783 ^ 2_n2);
assign 2_n9811 = ~(2_n7393 ^ 2_n11507);
assign 2_n1925 = ~(2_n10169 ^ 2_n2473);
assign 2_n9333 = ~2_n6507;
assign 2_n12179 = 2_n885 & 2_n5836;
assign 2_n618 = ~(2_n5773 | 2_n12664);
assign 2_n5992 = ~(2_n8417 ^ 2_n9857);
assign 2_n7771 = 2_n12150 | 2_n538;
assign 2_n12664 = 2_n10763 & 2_n11582;
assign 2_n4813 = 2_n2516 & 2_n11559;
assign 2_n8746 = ~2_n4919;
assign 2_n8314 = ~(2_n675 ^ 2_n2290);
assign 2_n1653 = 2_n2217 | 2_n1047;
assign 2_n2496 = 2_n2252 | 2_n8340;
assign 2_n11111 = ~2_n10702;
assign 2_n2901 = 2_n515 | 2_n5941;
assign 2_n8517 = ~(2_n2605 ^ 2_n11921);
assign 2_n317 = 2_n5355 | 2_n8970;
assign 2_n5244 = ~(2_n7054 ^ 2_n1040);
assign 2_n210 = ~(2_n8294 ^ 2_n7317);
assign 2_n11749 = 2_n7512 | 2_n12181;
assign 2_n12534 = ~(2_n302 ^ 2_n12214);
assign 2_n11560 = 2_n7299 & 2_n2239;
assign 2_n8338 = 2_n4029 & 2_n8834;
assign 2_n11643 = ~(2_n11212 ^ 2_n12002);
assign 2_n8069 = 2_n12825 & 2_n8744;
assign 2_n3192 = 2_n404 & 2_n429;
assign 2_n10056 = 2_n807 | 2_n6169;
assign 2_n12356 = ~2_n8823;
assign 2_n690 = 2_n7947 & 2_n493;
assign 2_n1078 = ~2_n9347;
assign 2_n7051 = 2_n6602 | 2_n2951;
assign 2_n1991 = ~(2_n10254 ^ 2_n8833);
assign 2_n4236 = ~(2_n3330 ^ 2_n7693);
assign 2_n2983 = 2_n5915 | 2_n6071;
assign 2_n10927 = ~(2_n9456 ^ 2_n3101);
assign 2_n2466 = 2_n1409 | 2_n12780;
assign 2_n5238 = ~(2_n8380 | 2_n1786);
assign 2_n1506 = 2_n686 | 2_n995;
assign 2_n8220 = 2_n1249 & 2_n7963;
assign 2_n2777 = ~(2_n4007 ^ 2_n7095);
assign 2_n1678 = 2_n4643 | 2_n8913;
assign 2_n5679 = 2_n2217 | 2_n9568;
assign 2_n7959 = 2_n10157 | 2_n28;
assign 2_n8146 = ~(2_n8741 ^ 2_n2942);
assign 2_n2838 = 2_n5575 | 2_n5538;
assign 2_n4293 = ~(2_n11317 ^ 2_n916);
assign 2_n4321 = 2_n10347 & 2_n12182;
assign 2_n10414 = 2_n7449 | 2_n12120;
assign 2_n11348 = ~(2_n532 ^ 2_n480);
assign 2_n410 = ~2_n1218;
assign 2_n9399 = ~2_n8529;
assign 2_n5207 = 2_n994 | 2_n3911;
assign 2_n9849 = 2_n1941 | 2_n3903;
assign 2_n6035 = ~(2_n9141 ^ 2_n901);
assign 2_n3226 = 2_n586 & 2_n6172;
assign 2_n1417 = ~(2_n372 | 2_n1060);
assign 2_n12678 = 2_n12471 & 2_n6433;
assign 2_n8087 = ~(2_n3044 ^ 2_n7066);
assign 2_n7420 = ~2_n478;
assign 2_n12490 = ~(2_n2277 ^ 2_n4865);
assign 2_n2358 = ~2_n4634;
assign 2_n8858 = ~2_n5157;
assign 2_n8702 = 2_n5008 | 2_n6841;
assign 2_n5035 = ~(2_n8085 ^ 2_n11814);
assign 2_n9411 = 2_n12870 & 2_n10107;
assign 2_n10106 = ~(2_n3105 ^ 2_n358);
assign 2_n8733 = ~2_n6483;
assign 2_n2904 = 2_n3457 | 2_n3786;
assign 2_n4184 = 2_n4457 | 2_n622;
assign 2_n1659 = 2_n4001 & 2_n592;
assign 2_n10613 = 2_n2217 | 2_n1739;
assign 2_n3473 = ~(2_n7373 | 2_n1340);
assign 2_n7875 = ~2_n12653;
assign 2_n1916 = ~(2_n8992 ^ 2_n5106);
assign 2_n5497 = ~2_n5212;
assign 2_n6648 = ~2_n6599;
assign 2_n1636 = ~2_n4406;
assign 2_n10772 = 2_n722 | 2_n3987;
assign 2_n3183 = ~(2_n5208 | 2_n4917);
assign 2_n3887 = 2_n7462 | 2_n2105;
assign 2_n1519 = ~2_n8449;
assign 2_n12208 = 2_n2456 | 2_n1163;
assign 2_n3007 = 2_n3127 | 2_n7341;
assign 2_n8760 = 2_n11293 & 2_n6013;
assign 2_n8218 = ~(2_n5288 | 2_n3040);
assign 2_n115 = ~2_n9512;
assign 2_n5271 = ~(2_n331 | 2_n11840);
assign 2_n12389 = ~(2_n11798 ^ 2_n11143);
assign 2_n10793 = 2_n10325 | 2_n10127;
assign 2_n5248 = 2_n3906 & 2_n11203;
assign 2_n2819 = ~(2_n9551 | 2_n4044);
assign 2_n582 = 2_n10750 | 2_n12080;
assign 2_n7935 = ~(2_n9559 ^ 2_n5050);
assign 2_n3953 = 2_n1097 & 2_n7456;
assign 2_n12754 = ~2_n447;
assign 2_n10342 = 2_n11812 & 2_n6879;
assign 2_n5267 = ~(2_n135 | 2_n11786);
assign 2_n4095 = ~(2_n3045 ^ 2_n8558);
assign 2_n10549 = ~(2_n10551 ^ 2_n7988);
assign 2_n145 = ~(2_n9519 ^ 2_n1648);
assign 2_n10645 = 2_n2455 | 2_n2567;
assign 2_n2700 = 2_n8959 | 2_n7952;
assign 2_n1881 = ~2_n6415;
assign 2_n1041 = 2_n10277 | 2_n6343;
assign 2_n4690 = ~(2_n11113 ^ 2_n1005);
assign 2_n7131 = 2_n686 | 2_n6455;
assign 2_n7569 = ~(2_n5437 ^ 2_n7104);
assign 2_n7548 = ~(2_n8757 ^ 2_n5031);
assign 2_n9897 = ~(2_n10948 | 2_n4359);
assign 2_n10612 = ~(2_n11050 ^ 2_n1336);
assign 2_n8877 = ~(2_n7091 | 2_n5427);
assign 2_n8888 = ~(2_n6880 ^ 2_n12440);
assign 2_n11141 = 2_n2515 & 2_n12489;
assign 2_n11326 = 2_n3722 ^ 2_n11793;
assign 2_n3403 = ~(2_n10590 ^ 2_n7821);
assign 2_n2089 = 2_n692 & 2_n8763;
assign 2_n3649 = ~(2_n4956 ^ 2_n10521);
assign 2_n3934 = ~(2_n12470 ^ 2_n4336);
assign 2_n6558 = ~(2_n7791 ^ 2_n1227);
assign 2_n7003 = ~(2_n3335 | 2_n5740);
assign 2_n3961 = 2_n240 | 2_n983;
assign 2_n11827 = ~2_n7265;
assign 2_n4670 = ~2_n438;
assign 2_n513 = ~(2_n5130 ^ 2_n9831);
assign 2_n1936 = ~2_n7469;
assign 2_n1886 = 2_n9050 | 2_n2873;
assign 2_n6511 = ~(2_n9797 ^ 2_n2900);
assign 2_n5810 = 2_n1012 & 2_n11537;
assign 2_n3440 = 2_n1543 & 2_n1600;
assign 2_n2103 = 2_n1752 | 2_n2688;
assign 2_n7898 = ~(2_n11683 ^ 2_n7110);
assign 2_n12002 = 2_n5915 | 2_n12754;
assign 2_n10943 = 2_n7625 | 2_n2709;
assign 2_n11338 = 2_n8405 | 2_n6513;
assign 2_n2917 = 2_n6977 | 2_n6455;
assign 2_n5000 = ~(2_n1135 ^ 2_n9409);
assign 2_n8984 = 2_n12611 | 2_n1437;
assign 2_n4060 = ~(2_n9806 | 2_n8579);
assign 2_n1526 = ~2_n5475;
assign 2_n5882 = 2_n6979 & 2_n6404;
assign 2_n6089 = ~(2_n7301 ^ 2_n3237);
assign 2_n7534 = ~2_n9647;
assign 2_n9857 = ~(2_n5179 ^ 2_n529);
assign 2_n10410 = 2_n8596 & 2_n3584;
assign 2_n8205 = 2_n10750 | 2_n5781;
assign 2_n11752 = ~2_n5167;
assign 2_n5038 = ~(2_n7869 ^ 2_n12455);
assign 2_n4962 = ~(2_n11690 ^ 2_n1914);
assign 2_n2798 = ~2_n10528;
assign 2_n12526 = 2_n6577 | 2_n3421;
assign 2_n7870 = ~(2_n11174 | 2_n2863);
assign 2_n9093 = 2_n4415 | 2_n325;
assign 2_n8288 = ~(2_n12879 | 2_n7792);
assign 2_n7058 = 2_n9107 | 2_n2986;
assign 2_n11919 = ~(2_n7081 ^ 2_n1713);
assign 2_n11014 = 2_n636 | 2_n5468;
assign 2_n10794 = 2_n9531 | 2_n1436;
assign 2_n2279 = ~(2_n4235 | 2_n7828);
assign 2_n4073 = ~2_n1821;
assign 2_n2377 = 2_n4167 & 2_n6892;
assign 2_n4120 = ~(2_n9733 ^ 2_n10564);
assign 2_n6331 = ~2_n1361;
assign 2_n7418 = ~(2_n2146 ^ 2_n2636);
assign 2_n9838 = 2_n4187 & 2_n2024;
assign 2_n10630 = ~(2_n1626 ^ 2_n1376);
assign 2_n7380 = 2_n6718 | 2_n4527;
assign 2_n135 = 2_n10831 & 2_n10959;
assign 2_n5493 = 2_n428 & 2_n244;
assign 2_n3978 = 2_n10727 & 2_n5662;
assign 2_n12624 = 2_n1335 | 2_n1440;
assign 2_n6698 = 2_n7138 | 2_n935;
assign 2_n1115 = 2_n8263 | 2_n4545;
assign 2_n2761 = 2_n2034 & 2_n2851;
assign 2_n10369 = ~2_n2966;
assign 2_n5252 = 2_n8641 & 2_n3890;
assign 2_n6728 = ~(2_n12831 ^ 2_n2915);
assign 2_n1367 = ~2_n1804;
assign 2_n5160 = 2_n9884 & 2_n3411;
assign 2_n4567 = ~(2_n10963 ^ 2_n465);
assign 2_n11716 = ~2_n6159;
assign 2_n9179 = 2_n5809 | 2_n1932;
assign 2_n2548 = 2_n5856 & 2_n10890;
assign 2_n7069 = ~(2_n8555 | 2_n11568);
assign 2_n9037 = 2_n4272 & 2_n11833;
assign 2_n9079 = 2_n752 | 2_n995;
assign 2_n12940 = 2_n10607 | 2_n341;
assign 2_n8708 = ~(2_n7005 | 2_n1291);
assign 2_n1875 = ~(2_n6903 | 2_n8419);
assign 2_n2448 = 2_n5530 | 2_n10422;
assign 2_n5391 = 2_n6373 | 2_n2020;
assign 2_n10125 = ~(2_n11834 ^ 2_n6459);
assign 2_n3801 = 2_n3078 & 2_n6895;
assign 2_n1402 = 2_n11984 | 2_n6460;
assign 2_n10571 = ~(2_n4217 | 2_n11726);
assign 2_n298 = ~(2_n9827 ^ 2_n12893);
assign 2_n1110 = ~(2_n3354 ^ 2_n8604);
assign 2_n9025 = ~(2_n7911 ^ 2_n6753);
assign 2_n11019 = 2_n808 & 2_n9934;
assign 2_n4039 = ~(2_n6291 | 2_n5035);
assign 2_n2826 = 2_n7745 & 2_n11854;
assign 2_n1074 = 2_n9881 & 2_n9474;
assign 2_n3655 = 2_n9437 & 2_n7908;
assign 2_n9282 = ~(2_n504 | 2_n3873);
assign 2_n8334 = ~2_n8159;
assign 2_n12329 = 2_n5915 | 2_n8109;
assign 2_n2517 = ~(2_n6133 ^ 2_n9913);
assign 2_n12197 = 2_n4358 | 2_n10165;
assign 2_n10877 = 2_n752 | 2_n2815;
assign 2_n3835 = ~(2_n12476 | 2_n485);
assign 2_n2678 = ~2_n7790;
assign 2_n3156 = 2_n7009 | 2_n4534;
assign 2_n8529 = 2_n7236 & 2_n9763;
assign 2_n11195 = 2_n2124 | 2_n3553;
assign 2_n12643 = 2_n4859 | 2_n2263;
assign 2_n7154 = 2_n8187 | 2_n7424;
assign 2_n301 = 2_n7232 | 2_n1013;
assign 2_n1966 = 2_n10104 & 2_n10498;
assign 2_n11333 = ~(2_n3876 ^ 2_n10111);
assign 2_n4229 = ~2_n3017;
assign 2_n196 = 2_n4628 | 2_n12735;
assign 2_n6856 = ~(2_n5107 ^ 2_n258);
assign 2_n9221 = ~(2_n1816 | 2_n5037);
assign 2_n10463 = 2_n3622 | 2_n7803;
assign 2_n6722 = ~(2_n5099 ^ 2_n570);
assign 2_n5342 = 2_n5902 | 2_n10066;
assign 2_n6002 = 2_n6776 & 2_n10451;
assign 2_n4464 = 2_n7391 | 2_n12843;
assign 2_n10797 = ~2_n1131;
assign 2_n527 = 2_n5655 | 2_n2296;
assign 2_n11458 = ~(2_n5394 ^ 2_n5152);
assign 2_n2053 = 2_n9914 | 2_n1573;
assign 2_n9755 = ~(2_n843 | 2_n717);
assign 2_n7966 = ~(2_n5615 ^ 2_n5717);
assign 2_n7302 = 2_n6374 & 2_n5757;
assign 2_n11623 = 2_n3691 | 2_n4315;
assign 2_n8879 = ~(2_n3464 | 2_n8805);
assign 2_n1459 = 2_n3571 & 2_n4869;
assign 2_n2743 = 2_n11846 | 2_n7117;
assign 2_n4888 = 2_n636 | 2_n8644;
assign 2_n12191 = ~2_n9590;
assign 2_n7447 = ~2_n5206;
assign 2_n2287 = 2_n7663 | 2_n11886;
assign 2_n8957 = ~2_n10685;
assign 2_n4354 = ~(2_n1160 | 2_n7162);
assign 2_n12333 = 2_n9170 | 2_n7703;
assign 2_n725 = 2_n4327 | 2_n8059;
assign 2_n295 = 2_n1303 & 2_n4754;
assign 2_n12188 = 2_n6286 | 2_n424;
assign 2_n6902 = 2_n5562 | 2_n4550;
assign 2_n3175 = ~2_n5039;
assign 2_n4004 = 2_n8977 & 2_n5040;
assign 2_n12201 = ~(2_n7519 ^ 2_n9371);
assign 2_n7955 = 2_n3038 | 2_n11124;
assign 2_n11679 = 2_n5530 | 2_n8109;
assign 2_n8947 = 2_n9685 & 2_n1926;
assign 2_n12237 = ~2_n4828;
assign 2_n12317 = 2_n1883 | 2_n105;
assign 2_n1162 = ~2_n2509;
assign 2_n8537 = ~(2_n9440 ^ 2_n7068);
assign 2_n4787 = 2_n10750 | 2_n1163;
assign 2_n9867 = ~(2_n7100 ^ 2_n9714);
assign 2_n208 = ~(2_n10399 ^ 2_n1426);
assign 2_n11095 = 2_n4549 & 2_n8215;
assign 2_n4904 = ~(2_n1131 ^ 2_n11159);
assign 2_n8927 = ~(2_n8171 ^ 2_n11111);
assign 2_n4521 = 2_n9784 & 2_n6920;
assign 2_n5108 = ~(2_n12405 ^ 2_n3415);
assign 2_n11396 = 2_n4911 | 2_n3911;
assign 2_n4275 = 2_n1333 & 2_n9195;
assign 2_n11262 = ~2_n12541;
assign 2_n861 = ~(2_n51 ^ 2_n3764);
assign 2_n3894 = ~(2_n6591 ^ 2_n10653);
assign 2_n99 = ~(2_n4658 | 2_n2723);
assign 2_n12808 = 2_n7620 & 2_n1724;
assign 2_n9107 = 2_n2099 | 2_n5326;
assign 2_n10430 = ~(2_n10135 ^ 2_n4632);
assign 2_n2990 = 2_n2848 & 2_n3695;
assign 2_n6813 = ~(2_n5500 ^ 2_n393);
assign 2_n10209 = ~(2_n10556 ^ 2_n7390);
assign 2_n4673 = ~(2_n1807 ^ 2_n6477);
assign 2_n9624 = 2_n2544 | 2_n9477;
assign 2_n9550 = 2_n12026 & 2_n6104;
assign 2_n8024 = 2_n10135 & 2_n9854;
assign 2_n1244 = ~(2_n2097 ^ 2_n8794);
assign 2_n8318 = 2_n6819 | 2_n3191;
assign 2_n8709 = ~(2_n284 ^ 2_n5010);
assign 2_n8038 = 2_n4403 | 2_n8198;
assign 2_n11779 = 2_n9632 & 2_n9210;
assign 2_n3789 = ~(2_n5189 | 2_n7960);
assign 2_n9999 = ~(2_n9729 ^ 2_n1690);
assign 2_n1119 = 2_n7839 | 2_n5540;
assign 2_n11214 = 2_n2774 | 2_n1617;
assign 2_n10620 = 2_n5328 | 2_n7647;
assign 2_n7330 = 2_n9352 & 2_n11275;
assign 2_n6907 = ~(2_n10592 ^ 2_n216);
assign 2_n9893 = ~(2_n1672 | 2_n8513);
assign 2_n8117 = 2_n3833 & 2_n11418;
assign 2_n9791 = ~(2_n6086 ^ 2_n2356);
assign 2_n6842 = ~(2_n10387 ^ 2_n3019);
assign 2_n5621 = 2_n3096 | 2_n995;
assign 2_n8160 = 2_n1344 & 2_n11207;
assign 2_n4212 = 2_n9536 & 2_n6755;
assign 2_n10151 = ~(2_n621 ^ 2_n6844);
assign 2_n2229 = 2_n1560 | 2_n12132;
assign 2_n258 = 2_n1183 | 2_n8740;
assign 2_n9617 = 2_n7914 | 2_n4351;
assign 2_n10440 = 2_n12729 | 2_n552;
assign 2_n3484 = ~(2_n4644 ^ 2_n9531);
assign 2_n7956 = ~(2_n1167 ^ 2_n8971);
assign 2_n5131 = ~2_n461;
assign 2_n3947 = 2_n5014 & 2_n11938;
assign 2_n4019 = ~(2_n7808 ^ 2_n2306);
assign 2_n10409 = 2_n10122 & 2_n11428;
assign 2_n150 = 2_n11153 & 2_n9763;
assign 2_n7382 = ~2_n12777;
assign 2_n8546 = 2_n5809 | 2_n1163;
assign 2_n980 = ~(2_n4932 ^ 2_n6550);
assign 2_n2446 = ~2_n5363;
assign 2_n9480 = ~(2_n1313 ^ 2_n5117);
assign 2_n5385 = 2_n7927 & 2_n5358;
assign 2_n9683 = ~(2_n7718 ^ 2_n1933);
assign 2_n1210 = 2_n3986 & 2_n10990;
assign 2_n7312 = 2_n3746 | 2_n6455;
assign 2_n9451 = 2_n5902 | 2_n4400;
assign 2_n7082 = 2_n6257 & 2_n8845;
assign 2_n11150 = ~2_n9284;
assign 2_n5427 = ~(2_n3970 | 2_n1364);
assign 2_n11672 = ~(2_n11109 ^ 2_n11391);
assign 2_n11069 = 2_n3096 | 2_n7952;
assign 2_n11151 = ~(2_n2129 ^ 2_n7529);
assign 2_n339 = 2_n10339 | 2_n4913;
assign 2_n8366 = 2_n8354 | 2_n8109;
assign 2_n157 = 2_n2160 | 2_n8725;
assign 2_n4778 = ~2_n7690;
assign 2_n2260 = ~2_n7783;
assign 2_n5084 = 2_n7310 | 2_n11202;
assign 2_n12252 = ~(2_n5014 | 2_n11938);
assign 2_n12264 = ~(2_n12010 ^ 2_n7886);
assign 2_n10854 = ~2_n7733;
assign 2_n7969 = 2_n3174 & 2_n12043;
assign 2_n7490 = 2_n2099 | 2_n10854;
assign 2_n11596 = 2_n4778 | 2_n3924;
assign 2_n9740 = 2_n5159 | 2_n2304;
assign 2_n8179 = ~(2_n9206 ^ 2_n293);
assign 2_n2084 = ~(2_n5516 ^ 2_n8517);
assign 2_n2845 = ~2_n5909;
assign 2_n4471 = ~2_n7276;
assign 2_n10434 = 2_n1937 | 2_n7952;
assign 2_n6575 = 2_n8040 & 2_n4677;
assign 2_n12778 = 2_n8560 & 2_n4532;
assign 2_n4642 = ~2_n2749;
assign 2_n9691 = ~(2_n2443 ^ 2_n3391);
assign 2_n4666 = 2_n10838 & 2_n3060;
assign 2_n849 = 2_n5422 & 2_n7885;
assign 2_n1908 = 2_n991 | 2_n354;
assign 2_n1497 = ~(2_n6452 ^ 2_n8226);
assign 2_n11090 = 2_n7474 | 2_n1681;
assign 2_n4665 = 2_n320 & 2_n8869;
assign 2_n6482 = 2_n10504 | 2_n6682;
assign 2_n5889 = 2_n3096 | 2_n12816;
assign 2_n11729 = 2_n5945 | 2_n11820;
assign 2_n3452 = 2_n752 | 2_n2589;
assign 2_n8584 = 2_n4911 | 2_n4400;
assign 2_n6725 = ~(2_n5639 ^ 2_n11146);
assign 2_n1580 = 2_n1699 | 2_n1163;
assign 2_n1811 = 2_n5915 | 2_n12080;
assign 2_n6930 = ~(2_n9744 | 2_n3963);
assign 2_n8673 = ~2_n9199;
assign 2_n76 = 2_n6669 | 2_n3568;
assign 2_n321 = 2_n8692 | 2_n2421;
assign 2_n12077 = ~(2_n3559 ^ 2_n11725);
assign 2_n5941 = 2_n12752 & 2_n1425;
assign 2_n5193 = 2_n4660 & 2_n4399;
assign 2_n10287 = ~(2_n2526 ^ 2_n9331);
assign 2_n9699 = ~2_n11108;
assign 2_n3669 = 2_n2157 | 2_n8245;
assign 2_n9078 = ~2_n12704;
assign 2_n1185 = 2_n5964 & 2_n2585;
assign 2_n3013 = ~2_n2771;
assign 2_n7401 = 2_n12119 | 2_n5468;
assign 2_n10812 = ~(2_n6415 | 2_n2871);
assign 2_n10745 = 2_n8959 | 2_n11820;
assign 2_n1107 = 2_n7251 | 2_n4264;
assign 2_n12559 = ~2_n9353;
assign 2_n9997 = 2_n989 | 2_n5497;
assign 2_n10496 = ~(2_n12463 ^ 2_n3197);
assign 2_n6189 = 2_n6718 | 2_n12771;
assign 2_n6549 = ~(2_n3334 ^ 2_n2580);
assign 2_n6138 = ~2_n11999;
assign 2_n955 = 2_n2727 & 2_n2735;
assign 2_n7704 = ~2_n384;
assign 2_n941 = ~(2_n289 ^ 2_n11681);
assign 2_n6081 = ~(2_n8213 ^ 2_n12073);
assign 2_n7530 = 2_n10835 | 2_n795;
assign 2_n9552 = ~(2_n11702 ^ 2_n4296);
assign 2_n5623 = ~(2_n11362 | 2_n2314);
assign 2_n7439 = 2_n3620 | 2_n5718;
assign 2_n1904 = ~(2_n2326 ^ 2_n10869);
assign 2_n476 = ~2_n12466;
assign 2_n5452 = 2_n5438 | 2_n11986;
assign 2_n6516 = 2_n3096 | 2_n7876;
assign 2_n7513 = 2_n4498 | 2_n2358;
assign 2_n1088 = 2_n8574 & 2_n8739;
assign 2_n1940 = ~(2_n5830 ^ 2_n6232);
assign 2_n11215 = ~(2_n3844 ^ 2_n3360);
assign 2_n12510 = ~2_n11395;
assign 2_n1752 = 2_n1315 & 2_n2211;
assign 2_n10167 = 2_n10671 & 2_n4295;
assign 2_n5338 = 2_n1686 & 2_n2898;
assign 2_n10583 = ~(2_n8117 ^ 2_n4976);
assign 2_n4635 = 2_n3820 | 2_n9568;
assign 2_n2619 = ~(2_n8357 ^ 2_n3670);
assign 2_n3502 = ~(2_n7936 ^ 2_n8298);
assign 2_n7619 = 2_n2326 & 2_n10869;
assign 2_n3306 = ~2_n12265;
assign 2_n2640 = 2_n5558 & 2_n316;
assign 2_n10507 = ~(2_n1815 | 2_n6225);
assign 2_n1098 = ~(2_n3780 ^ 2_n11357);
assign 2_n1880 = ~(2_n3170 ^ 2_n11583);
assign 2_n2117 = ~(2_n4756 ^ 2_n2323);
assign 2_n9524 = 2_n12361 | 2_n1413;
assign 2_n632 = 2_n3771 | 2_n3302;
assign 2_n9270 = 2_n3318 & 2_n2675;
assign 2_n6422 = 2_n2136 & 2_n10652;
assign 2_n1932 = ~2_n533;
assign 2_n9639 = ~2_n5317;
assign 2_n2485 = 2_n12786 & 2_n5687;
assign 2_n8471 = ~(2_n4850 ^ 2_n8016);
assign 2_n1501 = ~(2_n9385 ^ 2_n12529);
assign 2_n11540 = 2_n10157 | 2_n8285;
assign 2_n5279 = 2_n1937 | 2_n9741;
assign 2_n11158 = 2_n1434 | 2_n4887;
assign 2_n4066 = ~(2_n4753 | 2_n4851);
assign 2_n4259 = ~(2_n4126 ^ 2_n12608);
assign 2_n1822 = 2_n10344 & 2_n8541;
assign 2_n3605 = 2_n5605 | 2_n3745;
assign 2_n2143 = ~(2_n5880 ^ 2_n3243);
assign 2_n5255 = ~(2_n11846 ^ 2_n7117);
assign 2_n4641 = 2_n12322 | 2_n10872;
assign 2_n12631 = ~2_n585;
assign 2_n12493 = 2_n4692 & 2_n4977;
assign 2_n1252 = 2_n1646 & 2_n11866;
assign 2_n4496 = ~(2_n7408 ^ 2_n3547);
assign 2_n6691 = 2_n10991 | 2_n6056;
assign 2_n11100 = ~(2_n4783 | 2_n8840);
assign 2_n12038 = 2_n3822 & 2_n1071;
assign 2_n3928 = ~(2_n4320 ^ 2_n1840);
assign 2_n863 = ~(2_n2514 ^ 2_n12097);
assign 2_n2275 = ~(2_n768 ^ 2_n10131);
assign 2_n12521 = 2_n8251 | 2_n6109;
assign 2_n1068 = 2_n2649 | 2_n9926;
assign 2_n2140 = ~(2_n1317 ^ 2_n4386);
assign 2_n1341 = 2_n1941 | 2_n9741;
assign 2_n4387 = 2_n752 | 2_n8768;
assign 2_n1011 = 2_n589 | 2_n12321;
assign 2_n827 = ~2_n7672;
assign 2_n6956 = ~(2_n10802 ^ 2_n1122);
assign 2_n7740 = ~(2_n2958 ^ 2_n11663);
assign 2_n12675 = 2_n9544 | 2_n9882;
assign 2_n5741 = ~(2_n6917 ^ 2_n990);
assign 2_n6536 = ~(2_n7806 ^ 2_n519);
assign 2_n10554 = ~(2_n10548 ^ 2_n1579);
assign 2_n7723 = ~2_n6665;
assign 2_n6717 = ~(2_n9591 ^ 2_n10044);
assign 2_n6446 = ~(2_n2248 | 2_n5854);
assign 2_n5949 = 2_n10338 | 2_n6123;
assign 2_n11564 = ~(2_n10723 ^ 2_n10858);
assign 2_n11909 = ~(2_n7291 ^ 2_n9523);
assign 2_n10733 = 2_n4219 & 2_n1817;
assign 2_n7586 = ~2_n3372;
assign 2_n4580 = 2_n3534 & 2_n11350;
assign 2_n8547 = ~(2_n9547 ^ 2_n3194);
assign 2_n7357 = ~2_n4554;
assign 2_n7453 = 2_n6231 | 2_n3444;
assign 2_n5583 = ~2_n2161;
assign 2_n9385 = 2_n2827 & 2_n6170;
assign 2_n1475 = 2_n9389 | 2_n1162;
assign 2_n7860 = 2_n7883 | 2_n1595;
assign 2_n6732 = 2_n11087 | 2_n7183;
assign 2_n9435 = ~(2_n6178 ^ 2_n6494);
assign 2_n2 = ~(2_n548 ^ 2_n10859);
assign 2_n8388 = 2_n2022 | 2_n514;
assign 2_n4217 = 2_n4778 | 2_n4913;
assign 2_n4586 = 2_n11307 | 2_n1550;
assign 2_n5951 = ~(2_n8853 | 2_n9941);
assign 2_n12225 = 2_n347 & 2_n5560;
assign 2_n5158 = ~2_n6872;
assign 2_n9141 = 2_n752 | 2_n3356;
assign 2_n8791 = ~2_n2469;
assign 2_n10395 = 2_n3345 & 2_n2925;
assign 2_n3243 = ~(2_n1493 ^ 2_n4216);
assign 2_n6098 = 2_n11958 | 2_n5538;
assign 2_n2164 = 2_n12237 | 2_n1163;
assign 2_n11806 = ~(2_n11198 ^ 2_n12166);
assign 2_n11404 = ~(2_n9652 ^ 2_n1766);
assign 2_n7581 = ~(2_n1036 | 2_n11520);
assign 2_n1222 = ~2_n1251;
assign 2_n11504 = ~(2_n7434 ^ 2_n8063);
assign 2_n8187 = ~2_n6770;
assign 2_n3730 = 2_n1508 | 2_n9862;
assign 2_n511 = ~2_n2128;
assign 2_n9703 = ~(2_n11512 ^ 2_n5065);
assign 2_n4679 = ~(2_n718 ^ 2_n7454);
assign 2_n4083 = ~(2_n7171 ^ 2_n1999);
assign 2_n12484 = 2_n1955 & 2_n7008;
assign 2_n9408 = 2_n10506 | 2_n7060;
assign 2_n10154 = ~(2_n3920 ^ 2_n11164);
assign 2_n12067 = ~2_n866;
assign 2_n10346 = ~(2_n6995 | 2_n2405);
assign 2_n1945 = 2_n11097 & 2_n2935;
assign 2_n9661 = 2_n4838 | 2_n12102;
assign 2_n8008 = 2_n582 & 2_n11014;
assign 2_n6686 = 2_n10196 | 2_n4875;
assign 2_n8157 = 2_n5235 & 2_n433;
assign 2_n2699 = 2_n8583 | 2_n10916;
assign 2_n3147 = 2_n4632 | 2_n8024;
assign 2_n9927 = ~(2_n6167 | 2_n8883);
assign 2_n9584 = ~2_n4817;
assign 2_n9513 = 2_n12318 & 2_n6900;
assign 2_n3289 = ~(2_n11674 ^ 2_n7111);
assign 2_n11439 = 2_n1186 & 2_n12849;
assign 2_n7542 = ~(2_n3964 | 2_n1334);
assign 2_n10368 = ~(2_n4362 ^ 2_n5115);
assign 2_n9483 = 2_n12395 | 2_n11818;
assign 2_n958 = 2_n1539 | 2_n3911;
assign 2_n3168 = 2_n8127 | 2_n6389;
assign 2_n9254 = ~(2_n12262 ^ 2_n8253);
assign 2_n1422 = ~2_n9891;
assign 2_n9825 = 2_n3096 | 2_n9741;
assign 2_n3607 = 2_n10912 & 2_n6143;
assign 2_n10540 = ~(2_n9379 ^ 2_n5110);
assign 2_n11992 = ~(2_n7383 | 2_n4893);
assign 2_n5833 = 2_n8026 | 2_n3356;
assign 2_n11937 = ~(2_n5318 | 2_n1327);
assign 2_n1096 = 2_n2064 & 2_n5122;
assign 2_n9854 = ~(2_n2695 ^ 2_n9302);
assign 2_n9022 = 2_n8026 | 2_n5012;
assign 2_n525 = 2_n8966 | 2_n3960;
assign 2_n1789 = 2_n9878 | 2_n1163;
assign 2_n9030 = ~2_n9485;
assign 2_n11354 = 2_n5283 & 2_n2802;
assign 2_n9463 = ~(2_n7342 ^ 2_n9839);
assign 2_n6031 = ~2_n1655;
assign 2_n10669 = ~(2_n9849 ^ 2_n2664);
assign 2_n7726 = 2_n1962 & 2_n3147;
assign 2_n7289 = ~(2_n6339 ^ 2_n10539);
assign 2_n9007 = 2_n7933 | 2_n10989;
assign 2_n4042 = 2_n12503 | 2_n28;
assign 2_n11949 = ~2_n5598;
assign 2_n3091 = 2_n8344 | 2_n1756;
assign 2_n11724 = ~(2_n7592 ^ 2_n2775);
assign 2_n1278 = ~2_n7685;
assign 2_n2165 = 2_n2862 | 2_n8865;
assign 2_n11106 = 2_n9370 | 2_n7246;
assign 2_n12458 = 2_n12642 | 2_n12185;
assign 2_n9250 = 2_n9170 | 2_n7341;
assign 2_n10415 = ~(2_n2619 ^ 2_n4978);
assign 2_n3661 = ~(2_n7051 ^ 2_n12323);
assign 2_n3891 = 2_n8880 & 2_n12629;
assign 2_n481 = 2_n12797 | 2_n12816;
assign 2_n5724 = ~2_n8381;
assign 2_n352 = ~(2_n3534 ^ 2_n10914);
assign 2_n12907 = ~(2_n8562 | 2_n11642);
assign 2_n12841 = 2_n752 | 2_n10903;
assign 2_n7876 = ~2_n6703;
assign 2_n4858 = 2_n2031 | 2_n650;
assign 2_n11317 = ~(2_n1304 ^ 2_n7767);
assign 2_n5515 = ~2_n1139;
assign 2_n7399 = ~(2_n526 ^ 2_n3690);
assign 2_n4123 = ~(2_n9317 ^ 2_n12645);
assign 2_n1759 = 2_n5599 & 2_n7256;
assign 2_n1617 = ~(2_n10647 | 2_n7422);
assign 2_n11744 = 2_n11026 | 2_n9144;
assign 2_n4746 = 2_n76 & 2_n9323;
assign 2_n6150 = 2_n200 & 2_n6906;
assign 2_n4949 = ~(2_n701 ^ 2_n7036);
assign 2_n8634 = 2_n10142 | 2_n11746;
assign 2_n2349 = ~2_n10762;
assign 2_n5979 = ~2_n12657;
assign 2_n12263 = 2_n2217 | 2_n3606;
assign 2_n2130 = 2_n12186 | 2_n6169;
assign 2_n7079 = ~(2_n8606 ^ 2_n170);
assign 2_n4918 = ~(2_n882 ^ 2_n11209);
assign 2_n1810 = ~(2_n4701 ^ 2_n6811);
assign 2_n188 = 2_n11015 & 2_n12578;
assign 2_n6941 = ~2_n12712;
assign 2_n8426 = ~2_n3722;
assign 2_n263 = ~(2_n3503 ^ 2_n11139);
assign 2_n4901 = 2_n131 | 2_n1228;
assign 2_n11202 = 2_n636 | 2_n8740;
assign 2_n11163 = ~2_n7878;
assign 2_n2452 = ~(2_n5595 ^ 2_n8170);
assign 2_n10351 = 2_n1695 | 2_n8066;
assign 2_n3067 = 2_n12361 | 2_n6455;
assign 2_n821 = ~(2_n4257 ^ 2_n20);
assign 2_n12153 = ~(2_n2730 ^ 2_n10316);
assign 2_n2181 = ~(2_n11956 ^ 2_n1168);
assign 2_n4153 = 2_n8428 | 2_n1413;
assign 2_n765 = ~2_n11489;
assign 2_n3726 = 2_n7410 | 2_n3763;
assign 2_n12570 = ~(2_n144 ^ 2_n7137);
assign 2_n10088 = 2_n7899 | 2_n5485;
assign 2_n2694 = 2_n4498 | 2_n4242;
assign 2_n10353 = 2_n749 | 2_n8676;
assign 2_n4721 = 2_n6977 | 2_n1413;
assign 2_n4166 = 2_n7391 | 2_n10419;
assign 2_n5293 = ~(2_n1322 ^ 2_n2565);
assign 2_n5910 = ~(2_n7428 ^ 2_n1113);
assign 2_n10318 = 2_n7449 | 2_n7921;
assign 2_n7405 = ~(2_n10783 ^ 2_n12039);
assign 2_n3614 = ~2_n557;
assign 2_n1025 = ~2_n10336;
assign 2_n5258 = ~2_n11791;
assign 2_n4101 = 2_n9413 | 2_n9022;
assign 2_n5575 = ~2_n6877;
assign 2_n3539 = ~(2_n1945 | 2_n3972);
assign 2_n11115 = ~2_n5459;
assign 2_n2800 = 2_n182 | 2_n6267;
assign 2_n2246 = ~(2_n797 ^ 2_n12169);
assign 2_n5863 = ~(2_n9798 ^ 2_n11404);
assign 2_n10375 = ~(2_n5681 ^ 2_n4819);
assign 2_n5377 = 2_n8527 | 2_n11948;
assign 2_n1867 = ~(2_n3384 ^ 2_n2550);
assign 2_n1480 = ~(2_n10172 ^ 2_n8119);
assign 2_n7516 = ~(2_n3752 ^ 2_n2920);
assign 2_n3870 = 2_n2834 | 2_n10526;
assign 2_n7880 = ~(2_n357 ^ 2_n5306);
assign 2_n8660 = 2_n11478 & 2_n5645;
assign 2_n9240 = ~(2_n12741 ^ 2_n4229);
assign 2_n10739 = 2_n2763 | 2_n789;
assign 2_n2736 = 2_n8514 & 2_n7406;
assign 2_n12375 = ~(2_n9825 | 2_n8469);
assign 2_n4209 = 2_n10511 | 2_n484;
assign 2_n10393 = ~(2_n1274 ^ 2_n6492);
assign 2_n200 = ~2_n10265;
assign 2_n8347 = 2_n2456 | 2_n8648;
assign 2_n12523 = ~(2_n3706 ^ 2_n2625);
assign 2_n3344 = ~2_n6575;
assign 2_n2218 = ~(2_n1751 ^ 2_n4178);
assign 2_n1238 = 2_n11446 | 2_n9084;
assign 2_n2767 = ~(2_n12266 | 2_n10337);
assign 2_n12910 = ~(2_n3492 ^ 2_n698);
assign 2_n1817 = 2_n9228 | 2_n10931;
assign 2_n1992 = 2_n8026 | 2_n6084;
assign 2_n1513 = ~(2_n1675 ^ 2_n344);
assign 2_n12300 = ~(2_n10033 | 2_n11823);
assign 2_n4500 = 2_n4911 | 2_n1851;
assign 2_n4583 = 2_n1052 & 2_n266;
assign 2_n5653 = ~(2_n10847 ^ 2_n12626);
assign 2_n11335 = 2_n3743 | 2_n11698;
assign 2_n5816 = 2_n10202 | 2_n9729;
assign 2_n8479 = ~2_n6766;
assign 2_n9963 = ~2_n8628;
assign 2_n8198 = ~(2_n7777 ^ 2_n11872);
assign 2_n5843 = ~(2_n12516 | 2_n720);
assign 2_n4660 = 2_n2552 | 2_n6974;
assign 2_n9766 = ~(2_n8567 ^ 2_n341);
assign 2_n9720 = 2_n12755 | 2_n9954;
assign 2_n7931 = ~(2_n3046 ^ 2_n7201);
assign 2_n4468 = 2_n4414 & 2_n3781;
assign 2_n9898 = ~(2_n5155 ^ 2_n1860);
assign 2_n424 = ~2_n720;
assign 2_n2552 = ~2_n10973;
assign 2_n9130 = 2_n8629 & 2_n1498;
assign 2_n465 = ~(2_n3642 ^ 2_n7601);
assign 2_n5085 = ~(2_n7383 ^ 2_n12914);
assign 2_n4040 = ~2_n390;
assign 2_n11256 = ~(2_n2110 ^ 2_n11776);
assign 2_n620 = ~(2_n3442 ^ 2_n2694);
assign 2_n11013 = 2_n8552 | 2_n8655;
assign 2_n8580 = 2_n3303 & 2_n1744;
assign 2_n8955 = 2_n1183 | 2_n4913;
assign 2_n8802 = ~(2_n1123 ^ 2_n3729);
assign 2_n10506 = 2_n9373 | 2_n4654;
assign 2_n9166 = 2_n7310 & 2_n11202;
assign 2_n12128 = ~(2_n7554 ^ 2_n9792);
assign 2_n12488 = 2_n9977 | 2_n4375;
assign 2_n9779 = 2_n11825 & 2_n10592;
assign 2_n7053 = 2_n11902 & 2_n6883;
assign 2_n818 = ~(2_n4401 | 2_n9629);
assign 2_n9259 = ~2_n8418;
assign 2_n10419 = ~2_n5320;
assign 2_n6070 = 2_n11592 & 2_n12419;
assign 2_n3208 = 2_n9625 & 2_n5937;
assign 2_n6247 = 2_n5423 | 2_n1528;
assign 2_n979 = ~(2_n7940 | 2_n818);
assign 2_n7773 = 2_n2499 & 2_n5418;
assign 2_n4561 = 2_n12119 | 2_n5326;
assign 2_n3497 = 2_n4694 | 2_n2768;
assign 2_n1859 = 2_n7839 | 2_n12816;
assign 2_n7314 = ~(2_n10850 | 2_n9605);
assign 2_n722 = ~(2_n4390 ^ 2_n7748);
assign 2_n3601 = 2_n2464 & 2_n11023;
assign 2_n7218 = 2_n6636 | 2_n12215;
assign 2_n11297 = 2_n107 & 2_n10880;
assign 2_n4845 = 2_n4354 | 2_n11639;
assign 2_n11854 = 2_n3082 | 2_n2875;
assign 2_n3509 = 2_n527 & 2_n9816;
assign 2_n8931 = ~(2_n12622 ^ 2_n3919);
assign 2_n4886 = ~(2_n9222 ^ 2_n5162);
assign 2_n6546 = 2_n1086 | 2_n123;
assign 2_n6848 = 2_n2236 & 2_n3277;
assign 2_n5607 = 2_n4778 | 2_n8109;
assign 2_n2848 = 2_n7774 | 2_n7127;
assign 2_n383 = 2_n1887 & 2_n7903;
assign 2_n7190 = ~2_n4612;
assign 2_n9669 = 2_n656 & 2_n10580;
assign 2_n4631 = ~(2_n8348 ^ 2_n111);
assign 2_n678 = 2_n3243 | 2_n5880;
assign 2_n9194 = 2_n6621 & 2_n10910;
assign 2_n4433 = 2_n284 | 2_n10693;
assign 2_n3094 = ~(2_n8577 ^ 2_n8249);
assign 2_n12 = 2_n8412 & 2_n3521;
assign 2_n723 = ~(2_n4821 ^ 2_n48);
assign 2_n12336 = ~(2_n3232 ^ 2_n5997);
assign 2_n12134 = ~(2_n7305 | 2_n8872);
assign 2_n125 = ~2_n1948;
assign 2_n3663 = ~(2_n10116 ^ 2_n4679);
assign 2_n8768 = ~2_n10439;
assign 2_n764 = ~(2_n634 ^ 2_n11178);
assign 2_n4707 = 2_n3772 | 2_n4171;
assign 2_n10321 = ~(2_n3799 ^ 2_n4590);
assign 2_n9928 = ~(2_n8584 ^ 2_n7644);
assign 2_n9406 = ~(2_n11839 ^ 2_n12876);
assign 2_n5905 = ~(2_n8455 ^ 2_n6891);
assign 2_n7962 = ~2_n2015;
assign 2_n2930 = 2_n9428 | 2_n9981;
assign 2_n3042 = 2_n11182 & 2_n4200;
assign 2_n3697 = ~(2_n2819 ^ 2_n11830);
assign 2_n2723 = ~(2_n2787 | 2_n1208);
assign 2_n1972 = 2_n11281 | 2_n4629;
assign 2_n5345 = 2_n8959 | 2_n7876;
assign 2_n12405 = ~(2_n4715 ^ 2_n6503);
assign 2_n6683 = 2_n1471 & 2_n11876;
assign 2_n6934 = 2_n10738 | 2_n3150;
assign 2_n4926 = 2_n5915 | 2_n12535;
assign 2_n12314 = 2_n9564 ^ 2_n7680;
assign 2_n2125 = 2_n6697 | 2_n12225;
assign 2_n9157 = ~(2_n2976 ^ 2_n11495);
assign 2_n2473 = 2_n2188 & 2_n8006;
assign 2_n5064 = 2_n11958 | 2_n11820;
assign 2_n12768 = ~2_n8504;
assign 2_n7383 = 2_n10142 | 2_n7389;
assign 2_n5139 = ~(2_n11178 | 2_n634);
assign 2_n1153 = 2_n9273 & 2_n11048;
assign 2_n12605 = 2_n5214 & 2_n2616;
assign 2_n7695 = ~(2_n12144 ^ 2_n3153);
assign 2_n7561 = 2_n11165 & 2_n352;
assign 2_n10786 = ~(2_n12325 ^ 2_n7556);
assign 2_n3345 = 2_n8704 | 2_n5761;
assign 2_n10143 = ~(2_n5412 ^ 2_n12255);
assign 2_n10200 = 2_n12416 | 2_n9961;
assign 2_n6106 = ~2_n3499;
assign 2_n879 = 2_n326 & 2_n2904;
assign 2_n9923 = ~(2_n10788 ^ 2_n8523);
assign 2_n4323 = 2_n4667 & 2_n6199;
assign 2_n8379 = ~(2_n4984 ^ 2_n1153);
assign 2_n223 = ~(2_n5627 ^ 2_n1770);
assign 2_n11226 = ~2_n2418;
assign 2_n6100 = ~(2_n11378 | 2_n11991);
assign 2_n441 = 2_n12267 | 2_n12890;
assign 2_n1585 = ~(2_n3386 | 2_n129);
assign 2_n9853 = ~2_n6618;
assign 2_n3691 = 2_n8699 | 2_n228;
assign 2_n7328 = 2_n6219 & 2_n4959;
assign 2_n10197 = 2_n1539 | 2_n10066;
assign 2_n9027 = ~(2_n10777 ^ 2_n10171);
assign 2_n3769 = ~(2_n6250 ^ 2_n93);
assign 2_n10452 = ~(2_n3972 ^ 2_n4477);
assign 2_n10803 = 2_n4911 | 2_n1915;
assign 2_n9419 = ~(2_n9567 ^ 2_n5754);
assign 2_n8548 = 2_n10265 & 2_n11132;
assign 2_n6432 = ~(2_n12618 ^ 2_n10353);
assign 2_n8129 = ~(2_n5606 ^ 2_n7249);
assign 2_n0 = 2_n3743 | 2_n9568;
assign 2_n6484 = 2_n5815 | 2_n6018;
assign 2_n11083 = 2_n1474 | 2_n9633;
assign 2_n1081 = 2_n792 | 2_n2880;
assign 2_n12618 = ~(2_n10917 | 2_n6238);
assign 2_n4441 = 2_n2385 | 2_n5803;
assign 2_n4356 = 2_n3501 | 2_n4924;
assign 2_n6524 = ~2_n6604;
assign 2_n2422 = ~2_n3384;
assign 2_n4867 = 2_n12494 | 2_n12719;
assign 2_n10625 = ~2_n2104;
assign 2_n5369 = 2_n773 | 2_n12405;
assign 2_n8025 = 2_n12733 & 2_n5820;
assign 2_n3140 = 2_n191 | 2_n2076;
assign 2_n11302 = 2_n7918 | 2_n544;
assign 2_n434 = ~(2_n12739 | 2_n3108);
assign 2_n11375 = 2_n12946 & 2_n8265;
assign 2_n4140 = ~2_n6591;
assign 2_n1688 = 2_n10835 | 2_n28;
assign 2_n6255 = 2_n11914 & 2_n6839;
assign 2_n9134 = 2_n636 | 2_n9586;
assign 2_n5014 = ~(2_n12564 ^ 2_n8003);
assign 2_n426 = 2_n3118 | 2_n2203;
assign 2_n6388 = ~2_n11062;
assign 2_n5632 = ~(2_n8442 ^ 2_n4745);
assign 2_n3912 = 2_n11588 | 2_n5476;
assign 2_n3252 = 2_n6095 & 2_n781;
assign 2_n8043 = ~(2_n6981 ^ 2_n9149);
assign 2_n1046 = ~(2_n9837 ^ 2_n12126);
assign 2_n4260 = ~(2_n2746 ^ 2_n7887);
assign 2_n356 = ~(2_n12882 ^ 2_n11249);
assign 2_n12335 = ~2_n1577;
assign 2_n11739 = 2_n11433 | 2_n7952;
assign 2_n10962 = ~2_n2978;
assign 2_n9452 = ~2_n3833;
assign 2_n6001 = 2_n3821 | 2_n4701;
assign 2_n6078 = 2_n5915 | 2_n7382;
assign 2_n4438 = ~(2_n9995 ^ 2_n10754);
assign 2_n9148 = ~2_n3726;
assign 2_n11862 = 2_n2071 & 2_n10323;
assign 2_n272 = ~(2_n377 ^ 2_n1492);
assign 2_n5496 = ~2_n9016;
assign 2_n2878 = 2_n3692 & 2_n7649;
assign 2_n12620 = ~(2_n61 ^ 2_n8393);
assign 2_n4306 = ~(2_n1543 ^ 2_n1294);
assign 2_n4617 = ~2_n2665;
assign 2_n3968 = 2_n11090 & 2_n7010;
assign 2_n6468 = 2_n4396 | 2_n10296;
assign 2_n8432 = ~2_n5756;
assign 2_n6347 = 2_n11958 | 2_n10903;
assign 2_n4712 = ~(2_n5812 ^ 2_n5984);
assign 2_n12653 = 2_n4433 & 2_n2681;
assign 2_n8053 = 2_n9241 & 2_n7946;
assign 2_n5958 = ~(2_n158 | 2_n9260);
assign 2_n7386 = ~(2_n407 ^ 2_n4006);
assign 2_n5414 = 2_n989 | 2_n7424;
assign 2_n5490 = ~(2_n855 ^ 2_n5190);
assign 2_n2322 = 2_n3650 | 2_n1285;
assign 2_n8495 = ~(2_n9101 ^ 2_n9516);
assign 2_n1877 = 2_n12237 | 2_n12686;
assign 2_n8686 = 2_n5748 | 2_n5639;
assign 2_n3558 = 2_n5563 & 2_n5749;
assign 2_n4554 = 2_n4111 & 2_n4215;
assign 2_n5169 = ~(2_n11095 ^ 2_n10087);
assign 2_n5415 = ~2_n5504;
assign 2_n9342 = 2_n8851 & 2_n6768;
assign 2_n9146 = ~(2_n1039 | 2_n5611);
assign 2_n8545 = ~(2_n7338 ^ 2_n10267);
assign 2_n1077 = ~2_n9281;
assign 2_n10557 = ~(2_n10230 ^ 2_n10273);
assign 2_n3747 = 2_n5530 | 2_n9586;
assign 2_n11020 = ~(2_n4254 ^ 2_n5926);
assign 2_n5847 = ~(2_n8509 | 2_n3099);
assign 2_n5431 = ~2_n6917;
assign 2_n1055 = 2_n4270 ^ 2_n7579;
assign 2_n10789 = ~(2_n3343 ^ 2_n7849);
assign 2_n2771 = 2_n7364 & 2_n1843;
assign 2_n1325 = 2_n4707 | 2_n495;
assign 2_n9831 = ~(2_n4838 ^ 2_n5901);
assign 2_n9284 = 2_n7768 & 2_n2631;
assign 2_n4725 = 2_n11773 & 2_n7473;
assign 2_n2396 = ~(2_n3050 ^ 2_n11524);
assign 2_n4517 = ~(2_n4577 ^ 2_n4887);
assign 2_n436 = 2_n1664 & 2_n6851;
assign 2_n6055 = ~2_n4806;
assign 2_n1016 = ~(2_n3419 ^ 2_n4610);
assign 2_n10578 = 2_n2081 | 2_n4068;
assign 2_n11471 = 2_n9170 | 2_n1915;
assign 2_n7497 = 2_n4124 & 2_n11935;
assign 2_n2318 = 2_n11779 & 2_n2256;
assign 2_n10160 = ~(2_n555 ^ 2_n6841);
assign 2_n7752 = 2_n9170 | 2_n11827;
assign 2_n4600 = 2_n8607 & 2_n371;
assign 2_n789 = 2_n4059 | 2_n3911;
assign 2_n12143 = ~(2_n1651 | 2_n12695);
assign 2_n10650 = ~(2_n8277 ^ 2_n9724);
assign 2_n8543 = ~2_n2954;
assign 2_n5300 = ~(2_n12293 ^ 2_n5833);
assign 2_n6913 = 2_n11470 & 2_n7264;
assign 2_n333 = 2_n1099 & 2_n11183;
assign 2_n5688 = 2_n1619 & 2_n3477;
assign 2_n8739 = 2_n9366 | 2_n3709;
assign 2_n11580 = 2_n4787 | 2_n1889;
assign 2_n5234 = 2_n6151 & 2_n11219;
assign 2_n11362 = 2_n2446 & 2_n11631;
assign 2_n7952 = ~2_n1209;
assign 2_n6049 = 2_n4059 | 2_n1738;
assign 2_n8707 = ~(2_n6628 | 2_n11372);
assign 2_n1474 = ~(2_n7459 | 2_n4490);
assign 2_n11033 = 2_n7777 | 2_n11872;
assign 2_n6424 = ~(2_n7182 ^ 2_n5905);
assign 2_n3776 = 2_n7041 | 2_n2932;
assign 2_n6987 = ~(2_n10865 ^ 2_n8849);
assign 2_n11058 = 2_n8704 & 2_n5761;
assign 2_n9801 = 2_n1937 | 2_n11775;
assign 2_n1801 = ~(2_n12027 | 2_n10176);
assign 2_n2044 = 2_n11846 & 2_n7117;
assign 2_n1257 = 2_n4552 | 2_n12184;
assign 2_n3332 = 2_n2946 & 2_n7488;
assign 2_n11464 = ~(2_n5089 ^ 2_n10823);
assign 2_n7545 = 2_n9492 & 2_n4420;
assign 2_n2075 = ~(2_n5650 | 2_n11675);
assign 2_n136 = ~(2_n8140 | 2_n9877);
assign 2_n1427 = ~(2_n8531 ^ 2_n11985);
assign 2_n3963 = 2_n994 | 2_n1738;
assign 2_n4263 = ~(2_n3971 ^ 2_n10897);
assign 2_n1136 = ~(2_n4587 ^ 2_n4975);
assign 2_n6947 = ~(2_n11115 ^ 2_n3320);
assign 2_n1597 = ~(2_n11052 ^ 2_n7719);
assign 2_n12120 = ~2_n7270;
assign 2_n3902 = 2_n2040 & 2_n1605;
assign 2_n1792 = ~(2_n7609 ^ 2_n7907);
assign 2_n12638 = 2_n1728 | 2_n7627;
assign 2_n7338 = ~2_n5081;
assign 2_n4383 = ~(2_n8714 | 2_n9608);
assign 2_n4732 = ~(2_n8491 ^ 2_n10287);
assign 2_n7498 = 2_n1677 & 2_n6235;
assign 2_n7337 = 2_n10566 & 2_n6730;
assign 2_n5266 = ~2_n2650;
assign 2_n1386 = 2_n5448 | 2_n932;
assign 2_n11750 = ~2_n5233;
assign 2_n9271 = 2_n10835 | 2_n1476;
assign 2_n2720 = 2_n8354 | 2_n10854;
assign 2_n4420 = 2_n3096 | 2_n2815;
assign 2_n8224 = ~(2_n237 | 2_n4556);
assign 2_n4329 = ~(2_n2011 ^ 2_n6268);
assign 2_n11742 = ~2_n2571;
assign 2_n2323 = ~(2_n4552 ^ 2_n12011);
assign 2_n12209 = ~(2_n9695 ^ 2_n10708);
assign 2_n302 = 2_n967 & 2_n6615;
assign 2_n4484 = ~(2_n5391 ^ 2_n11320);
assign 2_n5691 = ~2_n1878;
assign 2_n8554 = ~2_n3070;
assign 2_n2821 = ~(2_n8124 | 2_n5367);
assign 2_n12522 = 2_n7709 | 2_n4527;
assign 2_n6765 = 2_n1715 | 2_n11329;
assign 2_n1574 = 2_n2071 | 2_n10323;
assign 2_n6075 = 2_n9170 | 2_n1455;
assign 2_n6290 = ~2_n2109;
assign 2_n10679 = ~(2_n9967 | 2_n7357);
assign 2_n5056 = ~(2_n9598 | 2_n4395);
assign 2_n10992 = 2_n3127 | 2_n1455;
assign 2_n2481 = ~(2_n12112 ^ 2_n12364);
assign 2_n6140 = 2_n12216 & 2_n10672;
assign 2_n7747 = 2_n4728 | 2_n10505;
assign 2_n12337 = 2_n12271 & 2_n12707;
assign 2_n831 = 2_n6685 | 2_n8604;
assign 2_n7508 = ~2_n8018;
assign 2_n9443 = ~(2_n12783 ^ 2_n12943);
assign 2_n772 = ~(2_n4506 ^ 2_n345);
assign 2_n10476 = ~(2_n12573 ^ 2_n1610);
assign 2_n7013 = ~(2_n2641 ^ 2_n11574);
assign 2_n665 = ~2_n12540;
assign 2_n7248 = ~(2_n12338 ^ 2_n2528);
assign 2_n8206 = ~(2_n10178 ^ 2_n9727);
assign 2_n10013 = 2_n587 & 2_n12665;
assign 2_n3901 = 2_n994 | 2_n11430;
assign 2_n11138 = ~2_n11393;
assign 2_n8755 = ~2_n11687;
assign 2_n12700 = 2_n11433 | 2_n6455;
assign 2_n2553 = ~(2_n7590 ^ 2_n10490);
assign 2_n569 = ~2_n1037;
assign 2_n5476 = ~(2_n11614 ^ 2_n7152);
assign 2_n8934 = ~(2_n3319 ^ 2_n516);
assign 2_n5141 = 2_n4873 | 2_n11880;
assign 2_n12564 = ~(2_n10181 ^ 2_n10126);
assign 2_n7855 = 2_n10471 | 2_n9765;
assign 2_n4069 = ~(2_n11001 ^ 2_n6528);
assign 2_n1927 = ~(2_n4367 | 2_n119);
assign 2_n6697 = 2_n3743 | 2_n4642;
assign 2_n10960 = 2_n6373 | 2_n1047;
assign 2_n2015 = 2_n4466 & 2_n9793;
assign 2_n8155 = ~(2_n9274 | 2_n10814);
assign 2_n7486 = 2_n2260 & 2_n2454;
assign 2_n10994 = ~(2_n11879 ^ 2_n7655);
assign 2_n662 = ~(2_n6725 ^ 2_n9344);
assign 2_n7939 = 2_n2456 | 2_n5781;
assign 2_n5200 = 2_n8552 | 2_n1932;
assign 2_n10998 = 2_n12025 & 2_n11407;
assign 2_n9455 = ~2_n5164;
assign 2_n3414 = 2_n9617 & 2_n139;
assign 2_n11524 = 2_n7449 | 2_n1509;
assign 2_n5333 = ~(2_n60 ^ 2_n11213);
assign 2_n8127 = ~2_n11821;
assign 2_n2413 = 2_n137 & 2_n2802;
assign 2_n926 = 2_n5345 | 2_n5711;
assign 2_n7849 = ~(2_n1890 ^ 2_n6436);
assign 2_n10930 = ~(2_n4855 | 2_n6753);
assign 2_n8675 = 2_n6551 & 2_n2086;
assign 2_n1383 = ~2_n6056;
assign 2_n6609 = ~(2_n12716 ^ 2_n10524);
assign 2_n9629 = ~(2_n10453 ^ 2_n7597);
assign 2_n1509 = ~2_n10848;
assign 2_n8843 = ~(2_n10579 ^ 2_n1888);
assign 2_n4750 = 2_n8870 | 2_n10854;
assign 2_n10564 = 2_n8051 | 2_n3966;
assign 2_n9885 = ~2_n3194;
assign 2_n1952 = 2_n3512 | 2_n10293;
assign 2_n12793 = ~(2_n991 ^ 2_n5664);
assign 2_n9961 = 2_n6368 & 2_n1309;
assign 2_n9635 = ~(2_n9231 ^ 2_n6395);
assign 2_n3557 = 2_n8810 & 2_n318;
assign 2_n9424 = ~(2_n4337 ^ 2_n6558);
assign 2_n2529 = 2_n9878 | 2_n5326;
assign 2_n2628 = ~(2_n10756 | 2_n3373);
assign 2_n10120 = ~(2_n573 ^ 2_n11044);
assign 2_n9609 = ~(2_n12234 | 2_n7292);
assign 2_n12590 = ~(2_n3810 | 2_n3181);
assign 2_n10882 = 2_n5765 | 2_n4654;
assign 2_n3949 = 2_n11571 & 2_n5511;
assign 2_n4539 = 2_n6227 & 2_n11129;
assign 2_n12011 = ~(2_n1637 ^ 2_n11325);
assign 2_n8600 = 2_n12705 & 2_n2509;
assign 2_n12406 = ~2_n2108;
assign 2_n5005 = ~(2_n680 | 2_n2996);
assign 2_n10046 = ~(2_n5903 | 2_n7119);
assign 2_n12757 = 2_n8476 & 2_n11967;
assign 2_n1831 = ~2_n12588;
assign 2_n400 = ~(2_n1919 ^ 2_n12615);
assign 2_n6157 = 2_n4365 & 2_n4323;
assign 2_n6174 = ~(2_n4165 ^ 2_n6878);
assign 2_n10856 = ~2_n11642;
assign 2_n5411 = ~(2_n604 ^ 2_n1329);
assign 2_n4308 = ~2_n11365;
assign 2_n2166 = ~(2_n2452 ^ 2_n11298);
assign 2_n342 = 2_n10960 & 2_n10315;
assign 2_n8002 = 2_n752 | 2_n11410;
assign 2_n4221 = ~2_n2364;
assign 2_n6751 = ~(2_n769 ^ 2_n3129);
assign 2_n4808 = 2_n4841 & 2_n6456;
assign 2_n6537 = 2_n12365 & 2_n11406;
assign 2_n9434 = ~(2_n5640 ^ 2_n6840);
assign 2_n6015 = 2_n6718 | 2_n8830;
assign 2_n11725 = ~(2_n5410 ^ 2_n460);
assign 2_n8049 = 2_n12666 & 2_n3624;
assign 2_n4647 = 2_n6577 | 2_n995;
assign 2_n9258 = 2_n11518 & 2_n878;
assign 2_n6634 = ~2_n12533;
assign 2_n10455 = 2_n3687 & 2_n532;
assign 2_n12354 = ~(2_n450 ^ 2_n11516);
assign 2_n5226 = 2_n7630 & 2_n5736;
assign 2_n12646 = 2_n8405 | 2_n3224;
assign 2_n1873 = ~(2_n10637 ^ 2_n12714);
assign 2_n12886 = 2_n4167 | 2_n6892;
assign 2_n248 = ~(2_n8104 ^ 2_n7934);
assign 2_n1189 = ~2_n4707;
assign 2_n8898 = 2_n3810 & 2_n3181;
assign 2_n284 = 2_n7116 | 2_n3903;
assign 2_n6872 = 2_n11033 & 2_n8038;
assign 2_n975 = 2_n11719 | 2_n5497;
assign 2_n5521 = ~(2_n4120 ^ 2_n10032);
assign 2_n11968 = 2_n8428 | 2_n7952;
assign 2_n6737 = 2_n3773 | 2_n12287;
assign 2_n10489 = 2_n6436 & 2_n7645;
assign 2_n10531 = 2_n1937 | 2_n6197;
assign 2_n10441 = ~(2_n12303 ^ 2_n6904);
assign 2_n285 = ~(2_n3015 ^ 2_n2294);
assign 2_n8377 = 2_n4283 | 2_n5524;
assign 2_n11632 = ~(2_n11501 ^ 2_n11188);
assign 2_n9053 = ~(2_n1503 | 2_n2839);
assign 2_n3855 = ~2_n5973;
assign 2_n11625 = 2_n5794 | 2_n4340;
assign 2_n11705 = ~(2_n5235 ^ 2_n11927);
assign 2_n7568 = ~(2_n1952 ^ 2_n2092);
assign 2_n7009 = 2_n9311 & 2_n9534;
assign 2_n11614 = ~(2_n7131 ^ 2_n8807);
assign 2_n12304 = ~2_n8952;
assign 2_n4310 = ~2_n8486;
assign 2_n2144 = 2_n1571 & 2_n1422;
assign 2_n8928 = ~(2_n12249 ^ 2_n3613);
assign 2_n8644 = ~2_n5069;
assign 2_n6584 = ~(2_n3125 ^ 2_n11199);
assign 2_n9730 = ~2_n11352;
assign 2_n5684 = 2_n8759 & 2_n12709;
assign 2_n10122 = ~2_n12692;
assign 2_n10127 = 2_n722 & 2_n3987;
assign 2_n4113 = ~2_n1639;
assign 2_n3525 = ~(2_n8221 ^ 2_n5445);
assign 2_n1850 = ~(2_n667 ^ 2_n10978);
assign 2_n6321 = ~(2_n6222 | 2_n3323);
assign 2_n6880 = 2_n6577 | 2_n7395;
assign 2_n7805 = ~(2_n3163 ^ 2_n8381);
assign 2_n8262 = ~(2_n1241 ^ 2_n492);
assign 2_n5709 = ~(2_n10381 | 2_n6177);
assign 2_n3009 = 2_n5945 | 2_n5540;
assign 2_n2627 = ~(2_n5776 ^ 2_n10454);
assign 2_n9470 = ~2_n6799;
assign 2_n8924 = 2_n9262 | 2_n4527;
assign 2_n11429 = ~2_n10512;
assign 2_n12695 = ~(2_n12167 | 2_n4774);
assign 2_n7713 = 2_n10750 | 2_n1932;
assign 2_n10502 = 2_n10157 | 2_n9568;
assign 2_n5947 = ~(2_n5992 ^ 2_n12384);
assign 2_n1464 = 2_n2743 & 2_n8597;
assign 2_n1933 = ~(2_n5679 ^ 2_n2963);
assign 2_n1938 = ~2_n5302;
assign 2_n10095 = 2_n3425 | 2_n7938;
assign 2_n7323 = 2_n3681 | 2_n7492;
assign 2_n10944 = ~2_n10059;
assign 2_n10852 = ~(2_n7665 ^ 2_n4557);
assign 2_n488 = ~2_n8015;
assign 2_n11700 = 2_n1183 | 2_n8655;
assign 2_n2459 = 2_n2217 | 2_n7921;
assign 2_n11096 = ~(2_n4923 ^ 2_n2693);
assign 2_n9649 = ~(2_n6649 | 2_n542);
assign 2_n7360 = ~(2_n11132 ^ 2_n200);
assign 2_n2664 = 2_n686 | 2_n11775;
assign 2_n7454 = ~(2_n5292 ^ 2_n369);
assign 2_n9149 = 2_n11923 | 2_n7921;
assign 2_n5629 = ~(2_n12590 | 2_n11035);
assign 2_n7503 = ~(2_n3808 | 2_n8460);
assign 2_n5823 = 2_n12237 | 2_n826;
assign 2_n6772 = 2_n2766 | 2_n1770;
assign 2_n3201 = 2_n10290 ^ 2_n3732;
assign 2_n10973 = ~(2_n6899 ^ 2_n8856);
assign 2_n2033 = ~(2_n9712 ^ 2_n7511);
assign 2_n507 = 2_n4322 | 2_n512;
assign 2_n5012 = ~2_n2024;
assign 2_n2432 = ~(2_n12530 ^ 2_n12779);
assign 2_n2382 = ~(2_n6478 ^ 2_n5973);
assign 2_n2543 = ~(2_n8307 | 2_n3539);
assign 2_n431 = 2_n8552 | 2_n10422;
assign 2_n12181 = ~(2_n10505 ^ 2_n11441);
assign 2_n10493 = 2_n11944 & 2_n5389;
assign 2_n2706 = 2_n4116 & 2_n7188;
assign 2_n12725 = 2_n1937 | 2_n5538;
assign 2_n9004 = ~(2_n1987 | 2_n3049);
assign 2_n3490 = ~(2_n1616 | 2_n1002);
assign 2_n7600 = ~(2_n2978 ^ 2_n6507);
assign 2_n9520 = 2_n11120 | 2_n12373;
assign 2_n4623 = ~2_n10409;
assign 2_n8320 = 2_n3617 | 2_n9188;
assign 2_n738 = 2_n3653 | 2_n5764;
assign 2_n1755 = 2_n2073 & 2_n12028;
assign 2_n3353 = ~2_n7925;
assign 2_n6299 = ~(2_n7292 ^ 2_n4786);
assign 2_n6472 = 2_n6577 | 2_n8768;
assign 2_n4717 = 2_n11552 | 2_n9568;
assign 2_n8524 = ~2_n2577;
assign 2_n1347 = 2_n5809 | 2_n12535;
assign 2_n12060 = ~(2_n9663 ^ 2_n6623);
assign 2_n10283 = 2_n12767 & 2_n6780;
assign 2_n6492 = ~(2_n3251 ^ 2_n6134);
assign 2_n5915 = ~2_n2530;
assign 2_n9305 = 2_n11887 | 2_n5468;
assign 2_n3455 = 2_n1708 | 2_n12114;
assign 2_n5801 = 2_n1183 | 2_n7382;
assign 2_n11836 = ~(2_n9223 ^ 2_n9747);
assign 2_n2604 = 2_n737 & 2_n6132;
assign 2_n11174 = ~(2_n8308 | 2_n6581);
assign 2_n3223 = ~(2_n2182 ^ 2_n11106);
assign 2_n3039 = 2_n9196 | 2_n8349;
assign 2_n1093 = 2_n6398 & 2_n9442;
assign 2_n3144 = ~2_n7327;
assign 2_n192 = ~2_n8053;
assign 2_n11050 = 2_n5496 & 2_n9603;
assign 2_n1242 = 2_n7283 | 2_n4400;
assign 2_n4738 = ~(2_n3140 | 2_n3447);
assign 2_n8623 = 2_n7293 | 2_n1641;
assign 2_n4943 = 2_n6098 & 2_n1845;
assign 2_n2737 = 2_n3767 & 2_n7600;
assign 2_n9626 = ~(2_n2759 ^ 2_n16);
assign 2_n8121 = ~(2_n6653 ^ 2_n2956);
assign 2_n11849 = 2_n1737 & 2_n11299;
assign 2_n9569 = ~(2_n8483 ^ 2_n2495);
assign 2_n3549 = 2_n7704 | 2_n9671;
assign 2_n8643 = ~2_n217;
assign 2_n5093 = 2_n5314 & 2_n2749;
assign 2_n6457 = ~2_n2788;
assign 2_n2841 = ~(2_n9024 | 2_n10201);
assign 2_n10834 = 2_n12173 & 2_n1405;
assign 2_n11628 = ~(2_n308 ^ 2_n1500);
assign 2_n331 = ~2_n6717;
assign 2_n4097 = 2_n4904 | 2_n701;
assign 2_n7276 = 2_n5439 & 2_n8083;
assign 2_n9255 = 2_n3672 & 2_n8255;
assign 2_n11880 = ~2_n6858;
assign 2_n11071 = 2_n7839 | 2_n11775;
assign 2_n9955 = 2_n10005 ^ 2_n791;
assign 2_n1125 = ~(2_n6974 ^ 2_n5719);
assign 2_n3996 = 2_n589 & 2_n12321;
assign 2_n2177 = ~(2_n7442 ^ 2_n568);
assign 2_n12568 = ~2_n4257;
assign 2_n9538 = 2_n7116 | 2_n6455;
assign 2_n12834 = ~(2_n5522 ^ 2_n115);
assign 2_n5743 = ~(2_n2418 | 2_n5274);
assign 2_n6978 = ~(2_n2516 ^ 2_n1064);
assign 2_n7292 = 2_n627 | 2_n11964;
assign 2_n12223 = 2_n10142 | 2_n8859;
assign 2_n1685 = ~2_n12956;
assign 2_n1963 = 2_n4373 | 2_n5628;
assign 2_n9653 = ~2_n12198;
assign 2_n897 = ~2_n6612;
assign 2_n7410 = 2_n12234 & 2_n7292;
assign 2_n8853 = ~2_n2055;
assign 2_n10520 = ~2_n816;
assign 2_n4779 = 2_n1453 ^ 2_n1000;
assign 2_n8181 = 2_n8026 | 2_n11896;
assign 2_n5051 = ~(2_n4914 ^ 2_n10227);
assign 2_n9677 = 2_n12853 | 2_n12735;
assign 2_n7180 = ~2_n10642;
assign 2_n30 = ~(2_n12089 ^ 2_n5879);
assign 2_n3258 = 2_n273 & 2_n9126;
assign 2_n7171 = 2_n6677 & 2_n12175;
assign 2_n10738 = 2_n12361 | 2_n7952;
assign 2_n4726 = 2_n2872 | 2_n12816;
assign 2_n4609 = ~(2_n2699 ^ 2_n10941);
assign 2_n108 = 2_n12062 | 2_n73;
assign 2_n12394 = 2_n3780 & 2_n6329;
assign 2_n2207 = 2_n2740 | 2_n2844;
assign 2_n2555 = ~(2_n12866 ^ 2_n194);
assign 2_n22 = ~2_n5947;
assign 2_n10111 = ~(2_n3448 ^ 2_n12744);
assign 2_n10147 = 2_n9108 & 2_n3983;
assign 2_n7783 = 2_n10196 | 2_n4654;
assign 2_n4806 = ~(2_n7289 ^ 2_n12141);
assign 2_n7639 = ~2_n8359;
assign 2_n10242 = 2_n128 | 2_n5460;
assign 2_n10212 = 2_n2332 | 2_n6034;
assign 2_n7976 = ~(2_n5867 ^ 2_n11522);
assign 2_n3668 = ~2_n4432;
assign 2_n2676 = ~2_n6980;
assign 2_n6626 = ~(2_n1147 ^ 2_n729);
assign 2_n7375 = ~(2_n11309 ^ 2_n7738);
assign 2_n3973 = ~(2_n2578 ^ 2_n5842);
assign 2_n7885 = 2_n5879 | 2_n2940;
assign 2_n12293 = ~(2_n3946 | 2_n7724);
assign 2_n3099 = ~(2_n11117 ^ 2_n7628);
assign 2_n4338 = 2_n12853 | 2_n10854;
assign 2_n5827 = ~(2_n814 ^ 2_n2847);
assign 2_n10505 = ~(2_n5524 ^ 2_n7877);
assign 2_n7802 = 2_n9905 | 2_n10792;
assign 2_n10276 = ~(2_n5539 ^ 2_n7430);
assign 2_n10488 = ~(2_n1061 ^ 2_n2685);
assign 2_n10413 = ~(2_n7783 ^ 2_n3710);
assign 2_n8835 = 2_n10835 | 2_n9078;
assign 2_n2463 = 2_n1044 & 2_n6668;
assign 2_n346 = 2_n11958 | 2_n8414;
assign 2_n5243 = ~(2_n12109 ^ 2_n3355);
assign 2_n948 = 2_n4900 | 2_n2219;
assign 2_n3299 = ~(2_n12584 | 2_n5733);
assign 2_n2442 = ~(2_n8085 | 2_n5180);
assign 2_n5461 = ~(2_n4490 ^ 2_n7459);
assign 2_n8364 = ~2_n11024;
assign 2_n10826 = 2_n6977 | 2_n11775;
assign 2_n2097 = 2_n2099 | 2_n7928;
assign 2_n5065 = ~(2_n7651 ^ 2_n10119);
assign 2_n2431 = ~(2_n7618 ^ 2_n12836);
assign 2_n1291 = ~2_n11094;
assign 2_n1306 = ~(2_n7327 ^ 2_n2971);
assign 2_n10683 = 2_n11415 & 2_n12606;
assign 2_n2102 = ~(2_n6462 ^ 2_n2094);
assign 2_n1060 = ~(2_n4633 ^ 2_n2255);
assign 2_n10604 = 2_n9878 | 2_n8109;
assign 2_n10107 = ~(2_n1652 ^ 2_n5498);
assign 2_n6248 = ~(2_n1524 | 2_n8540);
assign 2_n4990 = 2_n5964 & 2_n7265;
assign 2_n2920 = ~(2_n2116 ^ 2_n12452);
assign 2_n3210 = 2_n3820 | 2_n9144;
assign 2_n9915 = 2_n6373 | 2_n1476;
assign 2_n9088 = ~(2_n12208 ^ 2_n10017);
assign 2_n10326 = ~2_n9060;
assign 2_n12313 = 2_n7591 | 2_n1787;
assign 2_n5080 = ~(2_n10630 ^ 2_n12861);
assign 2_n7097 = 2_n11884 | 2_n5992;
assign 2_n233 = 2_n6977 | 2_n10903;
assign 2_n11357 = ~(2_n8598 ^ 2_n5581);
assign 2_n3316 = 2_n6283 | 2_n3543;
assign 2_n9190 = 2_n5355 | 2_n10419;
assign 2_n2641 = ~(2_n6734 | 2_n9049);
assign 2_n3933 = 2_n6534 | 2_n10826;
assign 2_n1709 = 2_n7552 | 2_n12553;
assign 2_n8480 = ~(2_n1790 ^ 2_n2016);
assign 2_n8891 = 2_n6162 | 2_n12432;
assign 2_n3298 = 2_n8552 | 2_n3224;
assign 2_n5066 = ~(2_n6015 ^ 2_n8673);
assign 2_n8386 = 2_n1183 | 2_n3924;
assign 2_n6621 = 2_n6877 & 2_n7946;
assign 2_n10616 = ~(2_n8990 ^ 2_n11496);
assign 2_n7172 = 2_n7804 & 2_n10341;
assign 2_n10799 = ~2_n1672;
assign 2_n2587 = 2_n3324 | 2_n28;
assign 2_n3350 = ~(2_n8585 ^ 2_n12187);
assign 2_n9980 = 2_n1459 & 2_n10330;
assign 2_n256 = ~(2_n10245 ^ 2_n8760);
assign 2_n4792 = 2_n1011 & 2_n864;
assign 2_n7678 = ~2_n1395;
assign 2_n2528 = ~2_n7865;
assign 2_n5664 = 2_n10750 | 2_n8109;
assign 2_n4528 = 2_n2332 & 2_n6034;
assign 2_n1207 = 2_n989 | 2_n7389;
assign 2_n9178 = 2_n7509 | 2_n3117;
assign 2_n5182 = 2_n6504 | 2_n3863;
assign 2_n7489 = 2_n9076 & 2_n4032;
assign 2_n3467 = ~(2_n6824 ^ 2_n6614);
assign 2_n3326 = 2_n5331 & 2_n1067;
assign 2_n10880 = 2_n1699 | 2_n9188;
assign 2_n377 = ~(2_n4440 ^ 2_n6083);
assign 2_n6818 = 2_n11337 | 2_n11092;
assign 2_n9280 = ~2_n6359;
assign 2_n870 = 2_n5638 | 2_n10767;
assign 2_n5962 = 2_n343 & 2_n7278;
assign 2_n6102 = 2_n2330 & 2_n6450;
assign 2_n1183 = ~2_n2515;
assign 2_n11587 = 2_n6626 | 2_n6106;
assign 2_n3027 = ~(2_n7883 ^ 2_n4341);
assign 2_n7216 = ~(2_n5850 ^ 2_n3218);
assign 2_n11435 = ~(2_n3491 ^ 2_n2954);
assign 2_n4188 = ~(2_n5341 ^ 2_n11947);
assign 2_n6171 = ~2_n6865;
assign 2_n2728 = 2_n289 & 2_n11772;
assign 2_n4909 = 2_n3282 & 2_n2907;
assign 2_n5247 = ~(2_n7463 ^ 2_n5146);
assign 2_n7715 = 2_n2689 | 2_n10649;
assign 2_n11526 = 2_n12392 | 2_n2231;
assign 2_n1676 = 2_n10450 | 2_n117;
assign 2_n8095 = 2_n5329 | 2_n9898;
assign 2_n6376 = ~2_n3574;
assign 2_n11085 = 2_n11225 & 2_n12559;
assign 2_n1378 = ~(2_n3949 | 2_n5935);
assign 2_n1465 = 2_n9373 | 2_n9568;
assign 2_n3325 = 2_n10350 | 2_n7081;
assign 2_n2031 = ~(2_n12437 ^ 2_n11238);
assign 2_n6586 = 2_n3386 & 2_n129;
assign 2_n8636 = ~(2_n3159 ^ 2_n3459);
assign 2_n7506 = ~2_n12947;
assign 2_n1599 = 2_n11923 | 2_n9568;
assign 2_n11961 = 2_n7495 | 2_n5497;
assign 2_n766 = 2_n3944 & 2_n334;
assign 2_n4797 = 2_n2496 & 2_n10452;
assign 2_n9888 = 2_n5337 | 2_n3492;
assign 2_n8339 = 2_n11552 | 2_n4474;
assign 2_n3606 = ~2_n1478;
assign 2_n4759 = 2_n4498 | 2_n7341;
assign 2_n11715 = ~(2_n7008 ^ 2_n155);
assign 2_n12625 = 2_n3909 & 2_n6105;
assign 2_n11175 = ~2_n12895;
assign 2_n12277 = ~(2_n3217 ^ 2_n5669);
assign 2_n2402 = 2_n2403 & 2_n6763;
assign 2_n3477 = ~2_n8975;
assign 2_n4715 = ~(2_n9113 ^ 2_n12032);
assign 2_n3261 = 2_n6426 | 2_n11009;
assign 2_n6045 = ~(2_n12016 ^ 2_n6082);
assign 2_n4234 = 2_n994 | 2_n5497;
assign 2_n2881 = ~(2_n11451 | 2_n6466);
assign 2_n901 = 2_n3746 | 2_n8414;
assign 2_n7413 = ~2_n9651;
assign 2_n1644 = ~(2_n7374 ^ 2_n7805);
assign 2_n12835 = ~2_n5032;
assign 2_n8832 = ~2_n3691;
assign 2_n910 = 2_n7283 | 2_n4242;
assign 2_n2434 = ~(2_n1507 ^ 2_n12153);
assign 2_n1651 = ~(2_n4972 | 2_n2542);
assign 2_n329 = ~(2_n12949 ^ 2_n8289);
assign 2_n10113 = 2_n9648 & 2_n5802;
assign 2_n9181 = ~(2_n9094 ^ 2_n5113);
assign 2_n667 = ~(2_n11608 ^ 2_n3839);
assign 2_n4698 = ~2_n1445;
assign 2_n6724 = ~(2_n12106 ^ 2_n8284);
assign 2_n2665 = 2_n7436 & 2_n11023;
assign 2_n10670 = 2_n8969 | 2_n10961;
assign 2_n12916 = 2_n9413 & 2_n9022;
assign 2_n11509 = ~(2_n3059 | 2_n10126);
assign 2_n5003 = 2_n994 | 2_n510;
assign 2_n7571 = ~2_n186;
assign 2_n684 = ~2_n12306;
assign 2_n7774 = ~(2_n5003 ^ 2_n892);
assign 2_n4915 = ~(2_n8486 ^ 2_n2411);
assign 2_n8469 = 2_n807 | 2_n12816;
assign 2_n8875 = 2_n9383 & 2_n8195;
assign 2_n9731 = 2_n1072 & 2_n2975;
assign 2_n501 = 2_n6218 & 2_n2156;
assign 2_n12331 = ~(2_n5350 | 2_n3540);
assign 2_n1791 = ~2_n7527;
assign 2_n5181 = 2_n12119 | 2_n12686;
assign 2_n3828 = 2_n10387 | 2_n3019;
assign 2_n4989 = 2_n718 & 2_n1643;
assign 2_n12629 = 2_n7951 | 2_n7215;
assign 2_n1369 = ~(2_n4166 ^ 2_n4261);
assign 2_n3764 = 2_n10108 | 2_n6389;
assign 2_n3396 = 2_n3096 | 2_n11775;
assign 2_n11701 = ~2_n7321;
assign 2_n12411 = 2_n2187 & 2_n9061;
assign 2_n2940 = ~(2_n83 | 2_n9710);
assign 2_n12894 = ~(2_n3109 ^ 2_n1103);
assign 2_n8254 = ~2_n11796;
assign 2_n1675 = 2_n3743 | 2_n7506;
assign 2_n9291 = ~2_n719;
assign 2_n1042 = 2_n9411 | 2_n12408;
assign 2_n8831 = ~(2_n10154 ^ 2_n5955);
assign 2_n6507 = 2_n4778 | 2_n826;
assign 2_n132 = ~(2_n4026 | 2_n12410);
assign 2_n5649 = 2_n2175 & 2_n1709;
assign 2_n451 = ~(2_n1126 ^ 2_n6970);
assign 2_n1541 = ~(2_n10222 ^ 2_n6842);
assign 2_n7237 = ~(2_n9055 | 2_n8077);
assign 2_n9697 = ~(2_n3906 | 2_n11203);
assign 2_n1240 = 2_n3746 | 2_n2815;
assign 2_n11461 = ~(2_n4131 ^ 2_n3973);
assign 2_n10916 = ~2_n806;
assign 2_n7640 = 2_n6373 | 2_n795;
assign 2_n1075 = 2_n3013 | 2_n10567;
assign 2_n8234 = ~(2_n4692 | 2_n4977);
assign 2_n7609 = ~(2_n12604 ^ 2_n11118);
assign 2_n564 = 2_n6986 & 2_n8595;
assign 2_n12175 = 2_n5399 | 2_n5400;
assign 2_n2451 = ~(2_n4635 ^ 2_n12369);
assign 2_n3240 = ~2_n6558;
assign 2_n11272 = 2_n12530 | 2_n12779;
assign 2_n4340 = ~(2_n6859 ^ 2_n10268);
assign 2_n11955 = 2_n3504 & 2_n524;
assign 2_n9214 = ~2_n1580;
assign 2_n8128 = ~(2_n2124 ^ 2_n3553);
assign 2_n11063 = 2_n4207 & 2_n3371;
assign 2_n9071 = ~2_n5684;
assign 2_n11875 = ~(2_n3297 ^ 2_n10757);
assign 2_n9313 = ~2_n8304;
assign 2_n4933 = ~2_n11677;
assign 2_n556 = 2_n5200 | 2_n1010;
assign 2_n7541 = ~2_n3724;
assign 2_n5275 = ~(2_n10730 | 2_n11104);
assign 2_n3381 = 2_n191 | 2_n1079;
assign 2_n520 = ~(2_n905 ^ 2_n3168);
assign 2_n4252 = 2_n12041 & 2_n10416;
assign 2_n5423 = 2_n9373 | 2_n9144;
assign 2_n7986 = ~(2_n3347 | 2_n8179);
assign 2_n4082 = ~(2_n1820 ^ 2_n3206);
assign 2_n4125 = ~(2_n2202 | 2_n8402);
assign 2_n1258 = ~(2_n11503 | 2_n10388);
assign 2_n11956 = ~(2_n11479 ^ 2_n4083);
assign 2_n3493 = 2_n5519 | 2_n1441;
assign 2_n1914 = 2_n5945 | 2_n995;
assign 2_n5667 = 2_n11455 | 2_n7614;
assign 2_n3125 = ~(2_n12959 ^ 2_n6355);
assign 2_n12269 = ~(2_n3570 | 2_n9972);
assign 2_n12127 = 2_n9079 | 2_n6414;
assign 2_n10903 = ~2_n11023;
assign 2_n9608 = ~(2_n5929 ^ 2_n8196);
assign 2_n829 = 2_n8552 | 2_n5468;
assign 2_n11116 = ~(2_n12056 | 2_n12678);
assign 2_n1998 = 2_n7534 | 2_n2079;
assign 2_n2366 = ~2_n7957;
assign 2_n11963 = ~2_n7463;
assign 2_n12507 = 2_n5915 | 2_n8259;
assign 2_n6478 = ~(2_n1220 ^ 2_n1410);
assign 2_n10228 = ~(2_n3873 ^ 2_n9320);
assign 2_n8074 = 2_n8836 | 2_n3941;
assign 2_n4830 = ~2_n7364;
assign 2_n12305 = ~(2_n1468 ^ 2_n9097);
assign 2_n2013 = 2_n4151 & 2_n3840;
assign 2_n6689 = ~(2_n7720 ^ 2_n1732);
assign 2_n6629 = 2_n2824 & 2_n10042;
assign 2_n5643 = ~(2_n6983 ^ 2_n10037);
assign 2_n12574 = ~2_n4989;
assign 2_n9124 = 2_n5684 & 2_n563;
assign 2_n2799 = ~(2_n98 ^ 2_n5768);
assign 2_n1152 = ~(2_n5393 ^ 2_n6733);
assign 2_n8553 = ~(2_n12932 ^ 2_n2320);
assign 2_n5503 = 2_n12776 & 2_n12587;
assign 2_n2240 = ~(2_n2965 ^ 2_n5968);
assign 2_n12694 = 2_n3025 | 2_n6054;
assign 2_n8648 = ~2_n6806;
assign 2_n10762 = 2_n7388 & 2_n12704;
assign 2_n4102 = ~(2_n12003 ^ 2_n10876);
assign 2_n10595 = 2_n7959 | 2_n2725;
assign 2_n12467 = ~2_n6356;
assign 2_n10596 = 2_n7539 & 2_n1328;
assign 2_n3929 = 2_n6137 & 2_n9404;
assign 2_n9756 = ~(2_n3479 ^ 2_n4505);
assign 2_n8413 = 2_n3560 | 2_n3505;
assign 2_n3453 = ~(2_n7739 | 2_n9057);
assign 2_n6958 = ~(2_n4316 ^ 2_n943);
assign 2_n10841 = ~(2_n11147 ^ 2_n12850);
assign 2_n6769 = 2_n1156 | 2_n871;
assign 2_n7999 = 2_n1362 | 2_n8878;
assign 2_n6454 = ~2_n1236;
assign 2_n6366 = ~(2_n11172 ^ 2_n4832);
assign 2_n9850 = ~(2_n4250 ^ 2_n7101);
assign 2_n11097 = ~2_n10522;
assign 2_n8867 = ~(2_n12785 ^ 2_n3806);
assign 2_n1930 = ~(2_n7366 ^ 2_n10062);
assign 2_n549 = ~(2_n337 ^ 2_n12329);
assign 2_n896 = ~2_n4119;
assign 2_n5337 = 2_n8373 | 2_n1940;
assign 2_n11745 = ~2_n1419;
assign 2_n10823 = 2_n4628 | 2_n5468;
assign 2_n5079 = ~(2_n1528 ^ 2_n2273);
assign 2_n8046 = 2_n9308 & 2_n9562;
assign 2_n2290 = ~(2_n3132 ^ 2_n435);
assign 2_n8850 = ~(2_n7632 ^ 2_n4518);
assign 2_n7254 = ~(2_n7697 ^ 2_n8566);
assign 2_n1604 = ~(2_n11 | 2_n10159);
assign 2_n10190 = ~2_n3973;
assign 2_n6348 = ~(2_n8235 | 2_n4597);
assign 2_n571 = ~(2_n6654 ^ 2_n3765);
assign 2_n10023 = ~(2_n5251 ^ 2_n7695);
assign 2_n2645 = ~(2_n11425 ^ 2_n6025);
assign 2_n3435 = ~2_n6195;
assign 2_n5492 = ~(2_n2944 | 2_n4398);
assign 2_n713 = 2_n2272 | 2_n10258;
assign 2_n2518 = ~(2_n6180 ^ 2_n3678);
assign 2_n8216 = 2_n752 | 2_n7952;
assign 2_n12334 = ~(2_n6347 ^ 2_n9890);
assign 2_n8656 = 2_n12069 & 2_n5645;
assign 2_n971 = 2_n4671 | 2_n8300;
assign 2_n3542 = ~(2_n8831 | 2_n3918);
assign 2_n11941 = ~2_n11836;
assign 2_n67 = 2_n4856 & 2_n10610;
assign 2_n1065 = 2_n10517 & 2_n8799;
assign 2_n9973 = ~(2_n3802 ^ 2_n8151);
assign 2_n10100 = 2_n1923 & 2_n6640;
assign 2_n9544 = ~(2_n456 ^ 2_n779);
assign 2_n3881 = ~(2_n3121 ^ 2_n2436);
assign 2_n2875 = 2_n10745 & 2_n12072;
assign 2_n954 = ~(2_n7914 ^ 2_n4351);
assign 2_n5450 = 2_n11716 | 2_n9460;
assign 2_n1452 = 2_n848 | 2_n2910;
assign 2_n3824 = ~(2_n6553 ^ 2_n11062);
assign 2_n11586 = 2_n12327 & 2_n1660;
assign 2_n7613 = ~2_n2890;
assign 2_n1631 = ~(2_n5407 ^ 2_n5390);
assign 2_n6019 = ~(2_n1515 | 2_n4832);
assign 2_n6750 = 2_n3084 & 2_n2801;
assign 2_n3609 = 2_n11851 & 2_n9255;
assign 2_n3965 = ~2_n6413;
assign 2_n3647 = 2_n3959 & 2_n2008;
assign 2_n2818 = ~(2_n6745 ^ 2_n2888);
assign 2_n7148 = ~(2_n4098 ^ 2_n11217);
assign 2_n5714 = ~(2_n1140 ^ 2_n10543);
assign 2_n4832 = ~2_n2218;
assign 2_n1135 = ~(2_n334 ^ 2_n9156);
assign 2_n12717 = ~(2_n8688 | 2_n7086);
assign 2_n1318 = ~(2_n1814 ^ 2_n5708);
assign 2_n1084 = ~2_n1217;
assign 2_n10901 = ~(2_n1072 ^ 2_n11051);
assign 2_n6215 = ~(2_n2532 ^ 2_n1880);
assign 2_n5717 = ~(2_n9546 ^ 2_n5184);
assign 2_n10314 = ~(2_n5456 ^ 2_n87);
assign 2_n12684 = ~(2_n6296 ^ 2_n10197);
assign 2_n7239 = ~(2_n11136 ^ 2_n8370);
assign 2_n10482 = 2_n3682 | 2_n8958;
assign 2_n7241 = ~(2_n2593 ^ 2_n8497);
assign 2_n7474 = 2_n8959 | 2_n9741;
assign 2_n332 = 2_n5949 & 2_n661;
assign 2_n11319 = ~2_n2411;
assign 2_n6394 = 2_n11805 & 2_n8047;
assign 2_n2857 = ~(2_n6036 ^ 2_n4348);
assign 2_n1558 = 2_n12855 | 2_n9717;
assign 2_n6966 = ~(2_n8736 | 2_n12526);
assign 2_n12525 = 2_n4628 | 2_n1932;
assign 2_n12073 = ~(2_n8225 ^ 2_n9202);
assign 2_n359 = ~(2_n11656 | 2_n1416);
assign 2_n10758 = ~(2_n8245 ^ 2_n8464);
assign 2_n4626 = ~(2_n5596 ^ 2_n9906);
assign 2_n1114 = ~2_n4897;
assign 2_n3120 = ~2_n7908;
assign 2_n2735 = 2_n8339 | 2_n4450;
assign 2_n5230 = 2_n9151 | 2_n951;
assign 2_n2096 = ~(2_n9038 ^ 2_n7623);
assign 2_n6845 = ~(2_n1585 | 2_n11269);
assign 2_n9869 = 2_n5355 | 2_n6389;
assign 2_n8105 = ~(2_n8320 | 2_n232);
assign 2_n1415 = 2_n3096 | 2_n11820;
assign 2_n2527 = ~(2_n4290 ^ 2_n12634);
assign 2_n3291 = 2_n12935 | 2_n9808;
assign 2_n4286 = ~(2_n197 ^ 2_n10689);
assign 2_n553 = ~(2_n8077 ^ 2_n3575);
assign 2_n11612 = ~(2_n4960 ^ 2_n4851);
assign 2_n4088 = ~(2_n2485 ^ 2_n9542);
assign 2_n11712 = 2_n2099 | 2_n2964;
assign 2_n4011 = ~(2_n2790 | 2_n666);
assign 2_n12355 = 2_n8642 | 2_n259;
assign 2_n8599 = ~2_n7286;
assign 2_n10222 = 2_n11635 | 2_n3037;
assign 2_n12446 = ~2_n4094;
assign 2_n8003 = 2_n6542 & 2_n8891;
assign 2_n1307 = ~(2_n4087 ^ 2_n5451);
assign 2_n4371 = 2_n6458 & 2_n9204;
assign 2_n6158 = 2_n7157 & 2_n6746;
assign 2_n11981 = ~(2_n6643 | 2_n9092);
assign 2_n3478 = 2_n5240 & 2_n4921;
assign 2_n2301 = ~(2_n1663 ^ 2_n7833);
assign 2_n1176 = ~(2_n12246 | 2_n287);
assign 2_n2035 = ~(2_n11060 ^ 2_n11247);
assign 2_n1985 = 2_n3236 | 2_n3067;
assign 2_n9092 = 2_n8736 & 2_n12526;
assign 2_n10628 = 2_n35 & 2_n887;
assign 2_n12086 = 2_n4728 & 2_n10505;
assign 2_n151 = ~2_n10790;
assign 2_n8067 = ~2_n11002;
assign 2_n5820 = 2_n11153 & 2_n8433;
assign 2_n8735 = ~2_n615;
assign 2_n6346 = ~(2_n6078 ^ 2_n2672);
assign 2_n2698 = ~(2_n9186 | 2_n7172);
assign 2_n11741 = 2_n7495 | 2_n6389;
assign 2_n2129 = ~(2_n1191 ^ 2_n9630);
assign 2_n12339 = ~(2_n8945 ^ 2_n11068);
assign 2_n6194 = ~(2_n4619 ^ 2_n9932);
assign 2_n9397 = ~2_n753;
assign 2_n3849 = ~(2_n1265 ^ 2_n4293);
assign 2_n12669 = ~2_n7693;
assign 2_n12112 = 2_n9370 | 2_n10066;
assign 2_n4899 = 2_n5915 | 2_n9586;
assign 2_n11727 = 2_n752 | 2_n5311;
assign 2_n957 = ~2_n10770;
assign 2_n12960 = 2_n12119 | 2_n5781;
assign 2_n6271 = 2_n6718 | 2_n4654;
assign 2_n9559 = ~(2_n2972 | 2_n10888);
assign 2_n12782 = ~(2_n12131 | 2_n11647);
assign 2_n12811 = 2_n1731 & 2_n2068;
assign 2_n5442 = 2_n8778 & 2_n12718;
assign 2_n8026 = ~2_n10928;
assign 2_n1090 = 2_n158 & 2_n9260;
assign 2_n5103 = ~(2_n5963 ^ 2_n4102);
assign 2_n3177 = ~(2_n9355 | 2_n2065);
assign 2_n6530 = ~2_n9345;
assign 2_n9528 = 2_n2739 & 2_n1033;
assign 2_n4703 = ~(2_n4232 ^ 2_n12549);
assign 2_n9700 = 2_n4540 | 2_n4448;
assign 2_n3068 = ~(2_n11318 ^ 2_n8924);
assign 2_n1902 = ~(2_n10507 ^ 2_n1484);
assign 2_n2786 = 2_n7713 | 2_n4012;
assign 2_n6258 = ~(2_n4612 ^ 2_n2417);
assign 2_n11485 = 2_n12586 | 2_n1320;
assign 2_n8777 = 2_n3630 | 2_n6831;
assign 2_n2783 = ~(2_n2311 | 2_n5206);
assign 2_n2224 = 2_n1494 | 2_n7198;
assign 2_n11626 = ~(2_n791 | 2_n5226);
assign 2_n11361 = 2_n11327 & 2_n599;
assign 2_n5272 = ~(2_n9122 ^ 2_n430);
assign 2_n5593 = 2_n2036 | 2_n2853;
assign 2_n4745 = ~(2_n5014 ^ 2_n11938);
assign 2_n9527 = 2_n8515 & 2_n10629;
assign 2_n12922 = ~(2_n3519 ^ 2_n6751);
assign 2_n8642 = ~(2_n12582 | 2_n10891);
assign 2_n1470 = 2_n10364 | 2_n5156;
assign 2_n986 = 2_n12845 & 2_n260;
assign 2_n7510 = 2_n10566 ^ 2_n2183;
assign 2_n2642 = 2_n989 | 2_n11430;
assign 2_n1664 = 2_n6131 | 2_n2060;
assign 2_n7495 = ~2_n12025;
assign 2_n5263 = ~(2_n11388 ^ 2_n11314);
assign 2_n9931 = 2_n636 | 2_n530;
assign 2_n28 = ~2_n5760;
assign 2_n3282 = 2_n12142 | 2_n4458;
assign 2_n9723 = 2_n11538 & 2_n8798;
assign 2_n5543 = 2_n6654 | 2_n8578;
assign 2_n4646 = 2_n2207 & 2_n5795;
assign 2_n391 = ~(2_n6472 ^ 2_n8457);
assign 2_n6916 = ~(2_n6310 ^ 2_n1606);
assign 2_n9715 = ~(2_n12855 ^ 2_n11989);
assign 2_n10302 = 2_n3007 & 2_n8561;
assign 2_n1974 = ~(2_n8986 | 2_n10680);
assign 2_n4368 = ~(2_n11986 ^ 2_n11644);
assign 2_n3051 = ~(2_n4756 | 2_n6010);
assign 2_n1775 = ~(2_n4202 ^ 2_n9497);
assign 2_n7313 = ~(2_n10098 | 2_n4004);
assign 2_n11457 = ~2_n9778;
assign 2_n10196 = ~2_n5860;
assign 2_n4932 = ~(2_n10475 ^ 2_n748);
assign 2_n5361 = 2_n12853 | 2_n7382;
assign 2_n847 = ~(2_n9150 ^ 2_n5308);
assign 2_n3959 = 2_n3746 | 2_n9741;
assign 2_n7987 = ~(2_n4457 ^ 2_n11041);
assign 2_n5878 = ~2_n6269;
assign 2_n4361 = ~(2_n4601 ^ 2_n7093);
assign 2_n7106 = ~(2_n10531 ^ 2_n670);
assign 2_n2472 = ~2_n952;
assign 2_n8633 = 2_n10835 | 2_n5759;
assign 2_n2186 = ~2_n2992;
assign 2_n4844 = 2_n6365 & 2_n6285;
assign 2_n250 = 2_n5353 & 2_n1171;
assign 2_n1139 = 2_n3820 | 2_n9160;
assign 2_n7637 = 2_n2523 & 2_n5753;
assign 2_n10168 = ~(2_n1999 | 2_n7171);
assign 2_n2269 = 2_n3367 & 2_n3056;
assign 2_n3715 = 2_n8564 | 2_n12226;
assign 2_n4181 = ~(2_n6148 ^ 2_n2748);
assign 2_n9906 = ~(2_n9508 ^ 2_n146);
assign 2_n4972 = 2_n5355 | 2_n5851;
assign 2_n902 = ~(2_n3596 | 2_n7345);
assign 2_n7760 = 2_n7271 & 2_n11263;
assign 2_n7155 = ~(2_n4286 ^ 2_n8472);
assign 2_n8057 = 2_n12227 & 2_n11940;
assign 2_n10631 = ~(2_n4513 ^ 2_n2331);
assign 2_n7746 = ~(2_n2057 ^ 2_n1431);
assign 2_n9729 = 2_n9373 | 2_n9521;
assign 2_n3666 = ~2_n9440;
assign 2_n1657 = ~2_n8671;
assign 2_n2174 = 2_n161 & 2_n550;
assign 2_n5001 = ~(2_n2892 ^ 2_n2299);
assign 2_n8177 = ~2_n4949;
assign 2_n8601 = 2_n5593 & 2_n2800;
assign 2_n1008 = 2_n6857 & 2_n4544;
assign 2_n9614 = 2_n807 | 2_n5012;
assign 2_n12872 = 2_n8556 & 2_n12794;
assign 2_n5726 = ~(2_n6374 ^ 2_n2230);
assign 2_n6508 = 2_n2763 & 2_n789;
assign 2_n6532 = ~(2_n5420 ^ 2_n7855);
assign 2_n9599 = ~(2_n25 | 2_n3952);
assign 2_n1894 = ~(2_n7085 ^ 2_n1725);
assign 2_n6139 = ~(2_n9383 ^ 2_n8195);
assign 2_n4892 = 2_n2217 | 2_n5914;
assign 2_n6849 = ~2_n2878;
assign 2_n5347 = 2_n12907 | 2_n12636;
assign 2_n5806 = ~(2_n1686 ^ 2_n860);
assign 2_n5063 = ~(2_n4255 ^ 2_n9501);
assign 2_n6603 = ~(2_n3133 ^ 2_n6541);
assign 2_n12536 = 2_n7932 & 2_n6065;
assign 2_n12408 = ~(2_n440 | 2_n5986);
assign 2_n4377 = 2_n4047 & 2_n7770;
assign 2_n27 = ~2_n6896;
assign 2_n12254 = ~(2_n11801 ^ 2_n4071);
assign 2_n8834 = 2_n7611 | 2_n1296;
assign 2_n1929 = ~2_n12309;
assign 2_n4572 = ~2_n2177;
assign 2_n12535 = ~2_n12925;
assign 2_n3795 = 2_n10394 & 2_n9265;
assign 2_n6238 = 2_n11011 & 2_n3869;
assign 2_n6418 = ~2_n1147;
assign 2_n11048 = 2_n796 | 2_n6116;
assign 2_n20 = ~(2_n8474 ^ 2_n12570);
assign 2_n229 = ~(2_n10627 ^ 2_n3656);
assign 2_n1409 = 2_n12119 | 2_n10422;
assign 2_n11514 = 2_n2832 | 2_n10066;
assign 2_n10145 = ~2_n7052;
assign 2_n9642 = ~2_n8892;
assign 2_n6087 = ~(2_n3047 ^ 2_n11403);
assign 2_n5794 = ~(2_n1550 ^ 2_n7129);
assign 2_n4961 = 2_n8026 | 2_n7425;
assign 2_n5019 = 2_n4904 & 2_n701;
assign 2_n6645 = ~(2_n10525 ^ 2_n1245);
assign 2_n10339 = ~2_n3146;
assign 2_n11925 = 2_n8428 | 2_n184;
assign 2_n8704 = 2_n994 | 2_n7881;
assign 2_n4710 = 2_n10750 | 2_n12754;
assign 2_n5636 = ~(2_n4868 | 2_n11379);
assign 2_n5191 = 2_n2342 ^ 2_n6926;
assign 2_n8248 = ~(2_n10529 | 2_n12337);
assign 2_n1392 = 2_n11958 | 2_n12899;
assign 2_n10229 = 2_n9043 & 2_n10840;
assign 2_n3632 = 2_n12208 & 2_n10017;
assign 2_n11440 = ~(2_n3150 ^ 2_n9127);
assign 2_n11178 = ~(2_n872 ^ 2_n230);
assign 2_n11942 = 2_n7705 & 2_n11863;
assign 2_n2892 = ~(2_n6668 ^ 2_n3637);
assign 2_n10792 = 2_n7449 | 2_n12771;
assign 2_n6462 = 2_n10987 & 2_n5526;
assign 2_n1924 = ~(2_n9530 ^ 2_n193);
assign 2_n6350 = ~(2_n7105 ^ 2_n6716);
assign 2_n12630 = 2_n4059 | 2_n10419;
assign 2_n10918 = ~(2_n6342 ^ 2_n3655);
assign 2_n7666 = ~(2_n9041 ^ 2_n6276);
assign 2_n6442 = 2_n4911 | 2_n7424;
assign 2_n8809 = 2_n5563 ^ 2_n4367;
assign 2_n8846 = ~(2_n8555 ^ 2_n6064);
assign 2_n2744 = ~(2_n1958 ^ 2_n5232);
assign 2_n551 = ~(2_n3982 ^ 2_n6005);
assign 2_n6012 = ~(2_n10368 ^ 2_n7269);
assign 2_n172 = ~(2_n8442 | 2_n12252);
assign 2_n10698 = 2_n12098 | 2_n5499;
assign 2_n8396 = 2_n8458 & 2_n3761;
assign 2_n5618 = ~(2_n2153 ^ 2_n704);
assign 2_n5977 = ~2_n804;
assign 2_n4946 = ~2_n12315;
assign 2_n3127 = ~2_n11757;
assign 2_n3073 = ~2_n3814;
assign 2_n3528 = ~(2_n10235 | 2_n3427);
assign 2_n308 = 2_n12119 | 2_n6513;
assign 2_n7580 = ~(2_n4374 ^ 2_n3595);
assign 2_n951 = ~(2_n695 ^ 2_n2389);
assign 2_n5386 = 2_n3096 | 2_n6169;
assign 2_n12382 = ~(2_n2999 | 2_n7484);
assign 2_n3069 = ~(2_n8102 ^ 2_n3854);
assign 2_n2208 = 2_n8428 | 2_n11775;
assign 2_n11173 = ~(2_n9275 ^ 2_n8402);
assign 2_n12322 = ~(2_n12211 | 2_n3394);
assign 2_n1303 = 2_n12327 | 2_n1660;
assign 2_n12399 = 2_n9701 & 2_n2799;
assign 2_n12868 = ~2_n9728;
assign 2_n2314 = ~(2_n6305 ^ 2_n4761);
assign 2_n11571 = 2_n1031 | 2_n8378;
assign 2_n11907 = ~2_n4583;
assign 2_n7125 = ~2_n8091;
assign 2_n778 = 2_n1937 | 2_n3421;
assign 2_n594 = ~(2_n3881 ^ 2_n10612);
assign 2_n10153 = ~(2_n6911 ^ 2_n52);
assign 2_n8849 = ~(2_n9082 ^ 2_n7944);
assign 2_n982 = 2_n12053 | 2_n4464;
assign 2_n7061 = 2_n2268 | 2_n3351;
assign 2_n11814 = ~(2_n7694 ^ 2_n12015);
assign 2_n3753 = ~(2_n4849 ^ 2_n963);
assign 2_n6404 = 2_n11681 | 2_n2728;
assign 2_n3390 = ~(2_n7737 ^ 2_n2000);
assign 2_n10425 = 2_n7461 & 2_n7892;
assign 2_n4955 = 2_n3221 & 2_n3314;
assign 2_n2394 = 2_n1833 | 2_n9684;
assign 2_n7706 = 2_n10585 | 2_n11862;
assign 2_n6762 = ~(2_n6058 ^ 2_n10182);
assign 2_n3526 = ~(2_n3036 ^ 2_n6549);
assign 2_n12948 = ~(2_n4380 ^ 2_n5245);
assign 2_n3499 = ~(2_n9072 ^ 2_n12574);
assign 2_n3198 = ~2_n868;
assign 2_n2648 = ~(2_n11245 ^ 2_n4725);
assign 2_n4860 = ~(2_n2846 ^ 2_n7904);
assign 2_n1827 = 2_n10478 | 2_n4055;
assign 2_n12257 = ~(2_n3003 ^ 2_n2843);
assign 2_n5634 = ~(2_n11156 ^ 2_n11906);
assign 2_n4537 = 2_n8618 | 2_n2247;
assign 2_n4935 = ~(2_n7655 | 2_n9410);
assign 2_n1567 = ~2_n3753;
assign 2_n5952 = ~(2_n12525 ^ 2_n6571);
assign 2_n1054 = ~(2_n5128 | 2_n5018);
assign 2_n5812 = 2_n10157 | 2_n11698;
assign 2_n1934 = 2_n10750 | 2_n5468;
assign 2_n12818 = 2_n6261 & 2_n6732;
assign 2_n3582 = 2_n8959 | 2_n5538;
assign 2_n3561 = 2_n11026 | 2_n4654;
assign 2_n2063 = ~(2_n7087 | 2_n611);
assign 2_n1449 = 2_n12361 | 2_n995;
assign 2_n4388 = ~(2_n3399 ^ 2_n4328);
assign 2_n1984 = ~(2_n9594 ^ 2_n2370);
assign 2_n2542 = 2_n4059 | 2_n12328;
assign 2_n6276 = ~(2_n8674 ^ 2_n5642);
assign 2_n7283 = ~2_n5964;
assign 2_n9354 = 2_n6977 | 2_n5540;
assign 2_n2124 = 2_n3746 | 2_n11896;
assign 2_n2647 = ~(2_n2661 | 2_n9511);
assign 2_n4775 = ~2_n2253;
assign 2_n414 = ~(2_n3078 ^ 2_n6032);
assign 2_n10661 = ~2_n6096;
assign 2_n6616 = 2_n9027 | 2_n1588;
assign 2_n10256 = 2_n7912 & 2_n4136;
assign 2_n11029 = ~2_n8129;
assign 2_n1395 = 2_n168 & 2_n6761;
assign 2_n11484 = ~2_n10747;
assign 2_n5073 = ~(2_n10932 ^ 2_n8425);
assign 2_n8646 = 2_n5977 & 2_n1716;
assign 2_n7315 = 2_n8813 & 2_n9401;
assign 2_n3732 = ~(2_n11777 ^ 2_n470);
assign 2_n11139 = 2_n9713 | 2_n9873;
assign 2_n7915 = ~(2_n9260 ^ 2_n3981);
assign 2_n9540 = ~(2_n1599 ^ 2_n11816);
assign 2_n11503 = 2_n6547 & 2_n670;
assign 2_n187 = 2_n12299 & 2_n8595;
assign 2_n5966 = 2_n2790 & 2_n666;
assign 2_n5034 = ~(2_n6390 ^ 2_n322);
assign 2_n1744 = 2_n29 | 2_n4027;
assign 2_n3650 = 2_n5530 | 2_n3924;
assign 2_n2198 = ~(2_n4279 ^ 2_n3446);
assign 2_n8632 = 2_n8132 & 2_n7867;
assign 2_n7011 = ~(2_n5482 | 2_n6960);
assign 2_n8544 = 2_n201 & 2_n8695;
assign 2_n2713 = 2_n2843 & 2_n3578;
assign 2_n5985 = ~2_n1355;
assign 2_n10757 = ~(2_n3140 ^ 2_n3447);
assign 2_n6417 = ~2_n2827;
assign 2_n95 = 2_n8091 & 2_n3759;
assign 2_n11889 = ~2_n3054;
assign 2_n6973 = 2_n9921 | 2_n10533;
assign 2_n6910 = ~(2_n871 ^ 2_n2769);
assign 2_n9563 = ~2_n3420;
assign 2_n6932 = ~(2_n5259 ^ 2_n828);
assign 2_n6327 = ~2_n8392;
assign 2_n12214 = ~2_n8844;
assign 2_n1944 = 2_n6423 | 2_n7786;
assign 2_n1100 = 2_n6204 & 2_n11735;
assign 2_n8019 = 2_n5429 & 2_n7702;
assign 2_n4794 = ~(2_n1696 ^ 2_n218);
assign 2_n2701 = 2_n4062 | 2_n5962;
assign 2_n5130 = ~(2_n8956 ^ 2_n12922);
assign 2_n1613 = ~(2_n9223 | 2_n12179);
assign 2_n6305 = 2_n8687 | 2_n4527;
assign 2_n12345 = ~(2_n2296 ^ 2_n8206);
assign 2_n12792 = 2_n11527 | 2_n8072;
assign 2_n4304 = 2_n8204 & 2_n3064;
assign 2_n8383 = 2_n4066 | 2_n8800;
assign 2_n10759 = 2_n1475 & 2_n4986;
assign 2_n959 = 2_n8070 & 2_n473;
assign 2_n7480 = 2_n10835 | 2_n609;
assign 2_n4729 = 2_n10709 | 2_n4822;
assign 2_n11630 = ~(2_n335 | 2_n6702);
assign 2_n4788 = 2_n5088 & 2_n3636;
assign 2_n2419 = 2_n4343 | 2_n12535;
assign 2_n5147 = 2_n7495 | 2_n1851;
assign 2_n1658 = ~(2_n11966 ^ 2_n9847);
assign 2_n11120 = 2_n4519 & 2_n7109;
assign 2_n10952 = ~2_n7064;
assign 2_n6543 = 2_n3820 | 2_n795;
assign 2_n7115 = ~2_n1016;
assign 2_n12473 = ~(2_n5499 ^ 2_n6638);
assign 2_n12170 = ~2_n11971;
assign 2_n6434 = ~(2_n3371 ^ 2_n11323);
assign 2_n11231 = ~(2_n3639 ^ 2_n6499);
assign 2_n10814 = 2_n6373 | 2_n12120;
assign 2_n2203 = ~(2_n3875 ^ 2_n657);
assign 2_n5273 = ~(2_n8770 | 2_n8248);
assign 2_n4111 = ~2_n8475;
assign 2_n13 = 2_n2832 | 2_n1162;
assign 2_n666 = 2_n4016 & 2_n9314;
assign 2_n7533 = 2_n6864 | 2_n451;
assign 2_n4093 = ~(2_n4042 | 2_n11666);
assign 2_n11895 = ~(2_n8145 ^ 2_n3449);
assign 2_n9110 = 2_n5844 & 2_n5938;
assign 2_n5002 = ~2_n4752;
assign 2_n8932 = ~(2_n2319 ^ 2_n1874);
assign 2_n2615 = 2_n874 | 2_n109;
assign 2_n7086 = ~(2_n1178 | 2_n3563);
assign 2_n9211 = 2_n8262 & 2_n3085;
assign 2_n9533 = ~(2_n10347 ^ 2_n12182);
assign 2_n675 = ~(2_n5556 ^ 2_n642);
assign 2_n4007 = ~(2_n8068 ^ 2_n11566);
assign 2_n11390 = 2_n11958 | 2_n9741;
assign 2_n7238 = 2_n3324 | 2_n4654;
assign 2_n6272 = ~(2_n5266 ^ 2_n12868);
assign 2_n12426 = 2_n6977 | 2_n6169;
assign 2_n3160 = ~2_n4577;
assign 2_n7219 = ~(2_n3901 | 2_n3929);
assign 2_n10026 = ~2_n9603;
assign 2_n5029 = 2_n6600 | 2_n2074;
assign 2_n6644 = 2_n4127 & 2_n5890;
assign 2_n7889 = 2_n12203 | 2_n10593;
assign 2_n4220 = 2_n1812 & 2_n10855;
assign 2_n9568 = ~2_n3342;
assign 2_n10987 = 2_n12069 & 2_n2498;
assign 2_n259 = 2_n7352 & 2_n3893;
assign 2_n5224 = 2_n835 & 2_n7979;
assign 2_n5689 = 2_n5518 | 2_n3990;
assign 2_n943 = 2_n1165 | 2_n1640;
assign 2_n11607 = ~(2_n4138 | 2_n4587);
assign 2_n9396 = ~(2_n2401 ^ 2_n11973);
assign 2_n750 = ~(2_n8936 ^ 2_n10192);
assign 2_n1298 = 2_n10735 & 2_n4091;
assign 2_n6185 = ~2_n10929;
assign 2_n4551 = ~(2_n895 ^ 2_n6206);
assign 2_n3424 = 2_n6718 | 2_n5258;
assign 2_n12207 = ~(2_n12920 ^ 2_n2113);
assign 2_n1283 = ~2_n5895;
assign 2_n5886 = 2_n3735 | 2_n2325;
assign 2_n1587 = 2_n3530 & 2_n11583;
assign 2_n6252 = 2_n10417 | 2_n10146;
assign 2_n4378 = ~(2_n12787 ^ 2_n2960);
assign 2_n6682 = ~(2_n1420 ^ 2_n557);
assign 2_n1371 = 2_n8477 & 2_n8952;
assign 2_n8316 = 2_n5064 & 2_n8974;
assign 2_n8219 = ~(2_n181 | 2_n5375);
assign 2_n8144 = ~(2_n10107 ^ 2_n6156);
assign 2_n573 = 2_n10142 | 2_n7341;
assign 2_n6121 = ~(2_n1973 ^ 2_n8779);
assign 2_n9380 = 2_n3728 | 2_n7740;
assign 2_n10198 = 2_n699 | 2_n7085;
assign 2_n5764 = 2_n3757 & 2_n10363;
assign 2_n1481 = 2_n827 & 2_n3264;
assign 2_n838 = ~(2_n7998 ^ 2_n4153);
assign 2_n1830 = 2_n9158 & 2_n2390;
assign 2_n8027 = 2_n10635 & 2_n8078;
assign 2_n8337 = ~2_n8585;
assign 2_n11960 = 2_n8127 | 2_n7424;
assign 2_n6311 = 2_n12275 | 2_n12086;
assign 2_n8341 = ~(2_n6569 ^ 2_n4031);
assign 2_n6658 = ~(2_n961 | 2_n9553);
assign 2_n1592 = 2_n2526 & 2_n8491;
assign 2_n2000 = ~(2_n11116 ^ 2_n10050);
assign 2_n9199 = 2_n3992 & 2_n12704;
assign 2_n1396 = 2_n6808 | 2_n9124;
assign 2_n11280 = 2_n11402 & 2_n6953;
assign 2_n2643 = 2_n4989 & 2_n4764;
assign 2_n12799 = 2_n1051 | 2_n11896;
assign 2_n1669 = 2_n3033 & 2_n1049;
assign 2_n12882 = 2_n10142 | 2_n8970;
assign 2_n8409 = 2_n97 & 2_n2129;
assign 2_n10574 = 2_n8428 | 2_n12899;
assign 2_n12842 = 2_n0 | 2_n9322;
assign 2_n3215 = 2_n7116 | 2_n7876;
assign 2_n11401 = 2_n12119 | 2_n8644;
assign 2_n4162 = ~(2_n2527 ^ 2_n7257);
assign 2_n3833 = 2_n1333 & 2_n2585;
assign 2_n9998 = ~(2_n6407 ^ 2_n2208);
assign 2_n2263 = ~(2_n1035 ^ 2_n2836);
assign 2_n5280 = ~(2_n8758 | 2_n12630);
assign 2_n7285 = 2_n11552 | 2_n9160;
assign 2_n8344 = 2_n7181 & 2_n11962;
assign 2_n2069 = 2_n191 | 2_n1851;
assign 2_n5140 = ~(2_n4656 ^ 2_n1781);
assign 2_n10682 = ~(2_n12923 | 2_n5966);
assign 2_n9692 = ~2_n7758;
assign 2_n12125 = ~(2_n6448 ^ 2_n7570);
assign 2_n5448 = ~(2_n2365 | 2_n9612);
assign 2_n7341 = ~2_n11917;
assign 2_n854 = 2_n5449 & 2_n427;
assign 2_n1607 = 2_n8583 | 2_n9160;
assign 2_n5609 = 2_n4154 & 2_n5746;
assign 2_n1826 = 2_n12119 | 2_n4913;
assign 2_n1351 = ~(2_n12316 ^ 2_n8576);
assign 2_n5713 = 2_n6993 & 2_n9915;
assign 2_n1173 = ~(2_n8216 ^ 2_n4183);
assign 2_n5440 = ~(2_n9415 ^ 2_n9968);
assign 2_n87 = 2_n12477 & 2_n9178;
assign 2_n12959 = ~(2_n5790 ^ 2_n12174);
assign 2_n4874 = 2_n3706 & 2_n10461;
assign 2_n10215 = ~(2_n2240 ^ 2_n6127);
assign 2_n4800 = ~(2_n6151 ^ 2_n694);
assign 2_n6316 = 2_n6977 | 2_n11410;
assign 2_n4694 = ~(2_n3965 | 2_n12778);
assign 2_n9890 = 2_n7282 & 2_n11604;
assign 2_n10246 = ~(2_n1003 ^ 2_n6265);
assign 2_n10608 = ~(2_n2917 ^ 2_n2426);
assign 2_n3062 = ~2_n5783;
assign 2_n3368 = 2_n8583 | 2_n5502;
assign 2_n6613 = 2_n2599 & 2_n10681;
assign 2_n9673 = ~(2_n4787 ^ 2_n1889);
assign 2_n11570 = ~(2_n132 ^ 2_n5637);
assign 2_n7235 = 2_n9048 & 2_n5993;
assign 2_n8533 = 2_n4059 | 2_n7703;
assign 2_n3187 = ~(2_n4339 ^ 2_n5246);
assign 2_n11939 = 2_n8870 | 2_n8109;
assign 2_n3429 = ~2_n3805;
assign 2_n5832 = 2_n752 | 2_n11820;
assign 2_n6149 = 2_n6182 & 2_n11336;
assign 2_n9704 = ~(2_n10718 | 2_n6585);
assign 2_n5779 = 2_n6881 | 2_n6489;
assign 2_n3314 = 2_n4059 | 2_n8524;
assign 2_n6632 = 2_n5548 | 2_n9768;
assign 2_n9143 = ~(2_n6387 ^ 2_n1487);
assign 2_n9782 = ~2_n5229;
assign 2_n4598 = ~(2_n6072 ^ 2_n5473);
assign 2_n8980 = ~(2_n6881 ^ 2_n6489);
assign 2_n9386 = ~(2_n10002 ^ 2_n2587);
assign 2_n7633 = ~2_n4260;
assign 2_n9176 = ~(2_n10304 ^ 2_n6928);
assign 2_n4533 = 2_n4951 | 2_n11496;
assign 2_n5412 = ~(2_n10137 ^ 2_n2179);
assign 2_n5227 = 2_n4648 & 2_n10473;
assign 2_n5590 = 2_n10479 & 2_n6884;
assign 2_n6301 = ~2_n10692;
assign 2_n10360 = 2_n7212 & 2_n8772;
assign 2_n4053 = 2_n2456 | 2_n8740;
assign 2_n7953 = ~(2_n6562 ^ 2_n8861);
assign 2_n4332 = 2_n5691 | 2_n6338;
assign 2_n11576 = 2_n9335 | 2_n11031;
assign 2_n4515 = 2_n9172 | 2_n11949;
assign 2_n7538 = 2_n11864 | 2_n8943;
assign 2_n5072 = ~(2_n710 ^ 2_n12851);
assign 2_n922 = ~(2_n3643 | 2_n8741);
assign 2_n8497 = ~(2_n5752 ^ 2_n5930);
assign 2_n5626 = ~(2_n7688 ^ 2_n11465);
assign 2_n10032 = ~2_n3975;
assign 2_n1735 = ~(2_n5146 | 2_n11963);
assign 2_n8460 = 2_n3498 & 2_n6048;
assign 2_n9018 = ~(2_n7919 ^ 2_n10756);
assign 2_n3012 = 2_n392 & 2_n9940;
assign 2_n11101 = 2_n10842 & 2_n5823;
assign 2_n8725 = 2_n10485 & 2_n2084;
assign 2_n739 = 2_n5005 | 2_n1968;
assign 2_n12164 = 2_n305 | 2_n3321;
assign 2_n10975 = ~(2_n1373 ^ 2_n1074);
assign 2_n10483 = ~(2_n12072 ^ 2_n6263);
assign 2_n12413 = 2_n5981 | 2_n5661;
assign 2_n10657 = 2_n420 & 2_n10308;
assign 2_n8231 = ~(2_n7185 ^ 2_n2895);
assign 2_n2561 = ~(2_n4124 | 2_n11935);
assign 2_n1440 = ~(2_n9161 ^ 2_n11766);
assign 2_n8612 = 2_n994 | 2_n5851;
assign 2_n4681 = 2_n8127 | 2_n11746;
assign 2_n852 = 2_n12790 ^ 2_n7255;
assign 2_n12418 = ~(2_n2427 ^ 2_n9801);
assign 2_n12699 = ~2_n1009;
assign 2_n5920 = ~(2_n10566 | 2_n6730);
assign 2_n11288 = 2_n5856 | 2_n10890;
assign 2_n10407 = ~(2_n3285 ^ 2_n5513);
assign 2_n12494 = ~(2_n1575 | 2_n6521);
assign 2_n8372 = ~(2_n10820 ^ 2_n10737);
assign 2_n467 = 2_n1290 | 2_n7002;
assign 2_n8918 = ~(2_n183 ^ 2_n10638);
assign 2_n11009 = 2_n9588 & 2_n3832;
assign 2_n2043 = ~(2_n10681 ^ 2_n5433);
assign 2_n8018 = ~(2_n11498 ^ 2_n5766);
assign 2_n5471 = 2_n1766 | 2_n1532;
assign 2_n2595 = 2_n6103 & 2_n11603;
assign 2_n7290 = ~(2_n4286 | 2_n8472);
assign 2_n12881 = 2_n9782 | 2_n7875;
assign 2_n3767 = 2_n8552 | 2_n3924;
assign 2_n1893 = ~(2_n9342 ^ 2_n6052);
assign 2_n3552 = 2_n1726 | 2_n3718;
assign 2_n283 = 2_n6373 | 2_n1509;
assign 2_n10946 = ~(2_n83 ^ 2_n30);
assign 2_n2646 = 2_n3875 | 2_n9585;
assign 2_n12812 = ~(2_n6095 ^ 2_n781);
assign 2_n4158 = ~(2_n11016 | 2_n3968);
assign 2_n7691 = ~2_n11702;
assign 2_n2754 = ~2_n1198;
assign 2_n8808 = ~(2_n1278 ^ 2_n8796);
assign 2_n6618 = 2_n5767 & 2_n9111;
assign 2_n3059 = ~2_n10181;
assign 2_n2228 = 2_n10835 | 2_n9280;
assign 2_n7874 = 2_n989 | 2_n7881;
assign 2_n12093 = ~2_n6050;
assign 2_n4762 = ~(2_n6575 ^ 2_n840);
assign 2_n9841 = 2_n5969 & 2_n1313;
assign 2_n10289 = ~(2_n6113 | 2_n4646);
assign 2_n7144 = 2_n10157 | 2_n5914;
assign 2_n37 = ~(2_n9444 ^ 2_n9291);
assign 2_n9062 = ~(2_n3570 ^ 2_n9972);
assign 2_n8510 = 2_n9370 | 2_n1851;
assign 2_n2313 = 2_n8428 | 2_n2232;
assign 2_n5460 = 2_n2722 & 2_n10136;
assign 2_n9012 = ~(2_n3072 ^ 2_n4750);
assign 2_n1343 = ~(2_n4591 | 2_n1235);
assign 2_n9204 = ~(2_n5624 ^ 2_n1450);
assign 2_n1844 = 2_n10514 & 2_n11187;
assign 2_n1514 = 2_n9368 | 2_n809;
assign 2_n7425 = ~2_n8819;
assign 2_n8514 = 2_n8423 | 2_n7315;
assign 2_n10908 = 2_n12237 | 2_n5326;
assign 2_n6338 = ~(2_n4871 ^ 2_n12090);
assign 2_n8103 = 2_n5575 | 2_n10919;
assign 2_n4037 = ~(2_n8596 ^ 2_n1007);
assign 2_n9321 = 2_n10142 | 2_n10066;
assign 2_n9991 = 2_n1719 | 2_n766;
assign 2_n7526 = ~(2_n11411 ^ 2_n3856);
assign 2_n583 = 2_n11923 | 2_n12120;
assign 2_n9462 = 2_n757 | 2_n3707;
assign 2_n1204 = ~(2_n8223 ^ 2_n988);
assign 2_n1628 = 2_n3407 | 2_n1087;
assign 2_n422 = 2_n5355 | 2_n561;
assign 2_n6990 = ~(2_n1306 ^ 2_n6417);
assign 2_n5924 = ~(2_n12278 | 2_n3853);
assign 2_n8841 = ~(2_n11547 ^ 2_n6832);
assign 2_n4130 = 2_n3680 | 2_n777;
assign 2_n4574 = ~(2_n2471 ^ 2_n2662);
assign 2_n7166 = 2_n4280 & 2_n7970;
assign 2_n7038 = 2_n12047 | 2_n3803;
assign 2_n10764 = ~(2_n759 ^ 2_n10907);
assign 2_n241 = ~(2_n10309 ^ 2_n11180);
assign 2_n3399 = 2_n5530 | 2_n12441;
assign 2_n862 = ~2_n6910;
assign 2_n6277 = 2_n8510 | 2_n8274;
assign 2_n9564 = ~(2_n10321 ^ 2_n6617);
assign 2_n7909 = 2_n10142 | 2_n5497;
assign 2_n9006 = ~(2_n9627 | 2_n833);
assign 2_n5174 = ~(2_n1328 ^ 2_n9359);
assign 2_n5326 = ~2_n521;
assign 2_n4981 = ~(2_n11703 ^ 2_n7648);
assign 2_n5881 = 2_n9520 & 2_n12624;
assign 2_n2536 = 2_n191 | 2_n7424;
assign 2_n10297 = 2_n4628 | 2_n7136;
assign 2_n2741 = 2_n1372 | 2_n1873;
assign 2_n1756 = 2_n8055 & 2_n3802;
assign 2_n6208 = 2_n11487 & 2_n4548;
assign 2_n10236 = 2_n12188 & 2_n11081;
assign 2_n10640 = 2_n8276 & 2_n3602;
assign 2_n4936 = ~2_n12342;
assign 2_n9713 = ~(2_n3098 | 2_n6711);
assign 2_n3438 = 2_n5561 | 2_n7682;
assign 2_n7304 = 2_n4498 | 2_n1162;
assign 2_n771 = 2_n7449 | 2_n11698;
assign 2_n5409 = 2_n5858 | 2_n10066;
assign 2_n7475 = 2_n374 & 2_n10595;
assign 2_n9175 = 2_n10530 & 2_n1038;
assign 2_n5981 = 2_n989 | 2_n1079;
assign 2_n2368 = 2_n5902 | 2_n11827;
assign 2_n7930 = 2_n2430 | 2_n640;
assign 2_n9384 = ~(2_n6256 ^ 2_n7489);
assign 2_n2602 = 2_n7391 | 2_n7703;
assign 2_n846 = ~2_n1956;
assign 2_n97 = 2_n2217 | 2_n5502;
assign 2_n2954 = 2_n7413 & 2_n10998;
assign 2_n9960 = 2_n12562 | 2_n8048;
assign 2_n3129 = ~(2_n5995 ^ 2_n8594);
assign 2_n12593 = ~(2_n763 ^ 2_n5979);
assign 2_n12432 = ~(2_n5793 ^ 2_n798);
assign 2_n5599 = 2_n35 | 2_n887;
assign 2_n3262 = 2_n191 | 2_n11430;
assign 2_n7394 = 2_n6373 | 2_n9280;
assign 2_n12089 = ~(2_n3255 ^ 2_n2398);
assign 2_n6833 = 2_n1683 | 2_n667;
assign 2_n10569 = ~2_n4210;
assign 2_n389 = ~2_n9925;
assign 2_n3553 = 2_n4509 & 2_n7930;
assign 2_n11118 = 2_n9262 | 2_n795;
assign 2_n1150 = ~2_n4168;
assign 2_n12853 = ~2_n137;
assign 2_n7264 = 2_n3975 | 2_n11321;
assign 2_n5752 = ~(2_n11779 ^ 2_n2007);
assign 2_n11900 = 2_n1572 | 2_n12710;
assign 2_n11890 = 2_n4059 | 2_n11746;
assign 2_n8253 = 2_n7202 & 2_n4103;
assign 2_n9393 = 2_n6750 | 2_n8346;
assign 2_n752 = ~2_n8759;
assign 2_n12472 = ~2_n12343;
assign 2_n1284 = ~2_n3111;
assign 2_n3642 = ~(2_n8918 ^ 2_n8764);
assign 2_n4138 = ~2_n9136;
assign 2_n2953 = 2_n2870 & 2_n6700;
assign 2_n11652 = ~2_n1330;
assign 2_n6095 = ~(2_n1940 ^ 2_n8889);
assign 2_n12744 = ~(2_n6655 ^ 2_n5827);
assign 2_n4923 = ~(2_n10989 ^ 2_n7716);
assign 2_n10063 = ~2_n2897;
assign 2_n3366 = ~(2_n12066 ^ 2_n10179);
assign 2_n8974 = 2_n8026 | 2_n1413;
assign 2_n3066 = 2_n107 | 2_n10880;
assign 2_n8142 = 2_n12539 & 2_n4623;
assign 2_n9842 = ~(2_n10841 ^ 2_n9560);
assign 2_n4239 = 2_n8570 & 2_n846;
assign 2_n12822 = 2_n7088 | 2_n7214;
assign 2_n11242 = ~(2_n11401 ^ 2_n2666);
assign 2_n40 = 2_n12691 & 2_n6543;
assign 2_n12787 = ~(2_n152 ^ 2_n9181);
assign 2_n6123 = 2_n12261 & 2_n3190;
assign 2_n2887 = 2_n11538 | 2_n8798;
assign 2_n12280 = 2_n12648 & 2_n7610;
assign 2_n3362 = 2_n686 | 2_n2232;
assign 2_n808 = ~(2_n1886 ^ 2_n12641);
assign 2_n5425 = 2_n3845 | 2_n10733;
assign 2_n11286 = ~(2_n5861 ^ 2_n9994);
assign 2_n12803 = 2_n12520 | 2_n12307;
assign 2_n8534 = ~(2_n2343 ^ 2_n8930);
assign 2_n3981 = ~(2_n158 ^ 2_n11961);
assign 2_n4547 = 2_n6678 | 2_n3267;
assign 2_n3323 = ~2_n8484;
assign 2_n10003 = ~2_n5369;
assign 2_n1104 = 2_n11821 & 2_n9956;
assign 2_n2289 = 2_n2677 | 2_n9579;
assign 2_n5630 = ~(2_n11997 | 2_n9582);
assign 2_n4148 = ~(2_n11895 ^ 2_n11157);
assign 2_n5896 = ~(2_n3817 | 2_n9276);
assign 2_n3858 = ~(2_n11772 ^ 2_n941);
assign 2_n6699 = ~(2_n9504 ^ 2_n11910);
assign 2_n11790 = ~(2_n325 ^ 2_n2609);
assign 2_n9343 = 2_n636 | 2_n4913;
assign 2_n11295 = ~(2_n8578 ^ 2_n571);
assign 2_n11005 = 2_n2456 | 2_n5468;
assign 2_n10591 = ~(2_n6606 ^ 2_n3582);
assign 2_n11291 = 2_n7809 & 2_n1095;
assign 2_n11841 = 2_n639 | 2_n1669;
assign 2_n9414 = 2_n11829 & 2_n4571;
assign 2_n9721 = 2_n9834 & 2_n7467;
assign 2_n990 = 2_n7107 & 2_n12400;
assign 2_n9089 = 2_n1236 & 2_n9289;
assign 2_n5132 = ~(2_n4833 ^ 2_n10496);
assign 2_n9404 = 2_n9370 | 2_n10419;
assign 2_n6995 = 2_n9878 | 2_n12080;
assign 2_n3529 = ~(2_n5988 | 2_n10706);
assign 2_n5845 = 2_n3992 & 2_n9763;
assign 2_n16 = ~(2_n10292 ^ 2_n11368);
assign 2_n8167 = ~2_n10322;
assign 2_n5303 = 2_n1012 | 2_n11537;
assign 2_n1503 = 2_n8127 | 2_n1162;
assign 2_n8531 = 2_n962 | 2_n9568;
assign 2_n1618 = ~2_n10941;
assign 2_n1376 = ~(2_n10342 | 2_n12382);
assign 2_n9566 = 2_n7025 | 2_n8234;
assign 2_n2991 = ~(2_n6074 ^ 2_n1400);
assign 2_n12104 = ~(2_n10694 ^ 2_n11012);
assign 2_n3792 = ~(2_n9001 ^ 2_n1650);
assign 2_n10548 = 2_n2456 | 2_n7136;
assign 2_n6181 = ~(2_n3864 | 2_n3246);
assign 2_n10445 = ~(2_n2004 ^ 2_n11398);
assign 2_n10538 = 2_n7686 & 2_n6074;
assign 2_n11989 = ~2_n327;
assign 2_n7487 = 2_n9389 | 2_n1079;
assign 2_n6353 = 2_n9400 & 2_n10451;
assign 2_n6743 = 2_n9416 | 2_n12276;
assign 2_n12403 = ~(2_n6681 ^ 2_n10894);
assign 2_n11064 = ~(2_n3845 ^ 2_n10733);
assign 2_n5499 = 2_n10196 | 2_n9521;
assign 2_n850 = 2_n7080 & 2_n10509;
assign 2_n8689 = ~(2_n1358 ^ 2_n12462);
assign 2_n10466 = 2_n12069 & 2_n12489;
assign 2_n664 = 2_n3944 | 2_n334;
assign 2_n10972 = 2_n2515 & 2_n2558;
assign 2_n4291 = 2_n10846 & 2_n5525;
assign 2_n731 = ~(2_n9308 ^ 2_n9562);
assign 2_n3498 = ~2_n9321;
assign 2_n361 = ~(2_n12684 ^ 2_n3697);
assign 2_n3036 = ~(2_n803 ^ 2_n743);
assign 2_n3876 = ~(2_n72 ^ 2_n9675);
assign 2_n6131 = ~(2_n3205 ^ 2_n12472);
assign 2_n12932 = ~(2_n3423 ^ 2_n8948);
assign 2_n328 = 2_n9370 | 2_n561;
assign 2_n701 = ~(2_n12834 ^ 2_n9992);
assign 2_n10074 = 2_n4480 & 2_n7866;
assign 2_n12431 = 2_n9791 & 2_n10393;
assign 2_n12460 = ~(2_n7369 ^ 2_n4867);
assign 2_n10581 = ~2_n11601;
assign 2_n11800 = 2_n2680 & 2_n12577;
assign 2_n4480 = 2_n5530 | 2_n530;
assign 2_n934 = 2_n11785 | 2_n11284;
assign 2_n4357 = 2_n9389 | 2_n10419;
assign 2_n3733 = 2_n2665 & 2_n5931;
assign 2_n4386 = 2_n5765 | 2_n4527;
assign 2_n2885 = 2_n4820 | 2_n3789;
assign 2_n12424 = 2_n3140 & 2_n3447;
assign 2_n6622 = 2_n1788 | 2_n11990;
assign 2_n12677 = ~(2_n9027 ^ 2_n2081);
assign 2_n11818 = 2_n5200 & 2_n1010;
assign 2_n8052 = 2_n10750 | 2_n2964;
assign 2_n9383 = 2_n9878 | 2_n7382;
assign 2_n4862 = 2_n695 | 2_n2389;
assign 2_n8092 = ~2_n11380;
assign 2_n237 = ~(2_n3206 | 2_n1820);
assign 2_n5918 = 2_n128 & 2_n5460;
assign 2_n4339 = ~(2_n10168 | 2_n1895);
assign 2_n2549 = 2_n7469 & 2_n12465;
assign 2_n8439 = ~(2_n2841 ^ 2_n7582);
assign 2_n10575 = 2_n12583 | 2_n10333;
assign 2_n213 = 2_n1 | 2_n4669;
assign 2_n11830 = 2_n4125 | 2_n2655;
assign 2_n8572 = 2_n2447 | 2_n9150;
assign 2_n1364 = ~(2_n6495 ^ 2_n2588);
assign 2_n10138 = ~(2_n8964 ^ 2_n10120);
assign 2_n2725 = 2_n1111 & 2_n11177;
assign 2_n5245 = 2_n11881 & 2_n10053;
assign 2_n7478 = ~(2_n9529 ^ 2_n7950);
assign 2_n3119 = 2_n7157 ^ 2_n11079;
assign 2_n139 = 2_n11034 | 2_n2583;
assign 2_n10072 = ~(2_n6752 | 2_n12017);
assign 2_n1812 = 2_n762 | 2_n6312;
assign 2_n6882 = ~(2_n794 | 2_n2083);
assign 2_n10664 = ~2_n5603;
assign 2_n7206 = 2_n191 | 2_n1162;
assign 2_n686 = ~2_n4203;
assign 2_n6379 = ~(2_n1655 ^ 2_n3787);
assign 2_n7161 = ~2_n8102;
assign 2_n7615 = 2_n2984 & 2_n7350;
assign 2_n6736 = ~(2_n9369 ^ 2_n2952);
assign 2_n11045 = 2_n5690 & 2_n1607;
assign 2_n9019 = ~(2_n12139 ^ 2_n8043);
assign 2_n8588 = 2_n5945 | 2_n9741;
assign 2_n3232 = ~(2_n7304 ^ 2_n11017);
assign 2_n9678 = ~(2_n182 ^ 2_n11549);
assign 2_n11462 = ~(2_n2349 ^ 2_n4308);
assign 2_n8805 = 2_n3746 | 2_n3468;
assign 2_n2829 = 2_n11661 | 2_n6279;
assign 2_n11574 = 2_n6921 | 2_n8812;
assign 2_n9978 = ~2_n12506;
assign 2_n12906 = 2_n10879 | 2_n1079;
assign 2_n11444 = ~(2_n8156 | 2_n6908);
assign 2_n1197 = 2_n11923 | 2_n28;
assign 2_n287 = 2_n10361 & 2_n6305;
assign 2_n4117 = 2_n5007 | 2_n2377;
assign 2_n5216 = ~(2_n11873 | 2_n1758);
assign 2_n1423 = 2_n9652 | 2_n9798;
assign 2_n5972 = 2_n5102 & 2_n10400;
assign 2_n9601 = ~(2_n6446 ^ 2_n10660);
assign 2_n5262 = 2_n2491 & 2_n3725;
assign 2_n3799 = ~(2_n5796 ^ 2_n9673);
assign 2_n10457 = ~(2_n6920 ^ 2_n1262);
assign 2_n1630 = ~2_n3478;
assign 2_n8173 = ~2_n7012;
assign 2_n674 = ~2_n10777;
assign 2_n9873 = ~(2_n4196 | 2_n11519);
assign 2_n3445 = 2_n9271 | 2_n1866;
assign 2_n5142 = ~(2_n639 ^ 2_n88);
assign 2_n12707 = 2_n7283 | 2_n7246;
assign 2_n728 = ~(2_n9069 ^ 2_n5785);
assign 2_n5996 = 2_n1802 | 2_n1869;
assign 2_n12457 = ~(2_n3528 ^ 2_n4944);
assign 2_n10551 = ~(2_n733 ^ 2_n682);
assign 2_n7167 = ~2_n9942;
assign 2_n12855 = ~(2_n4711 ^ 2_n10822);
assign 2_n11654 = 2_n9140 | 2_n3592;
assign 2_n4934 = ~2_n11164;
assign 2_n11367 = ~2_n10862;
assign 2_n12596 = ~2_n11099;
assign 2_n7464 = 2_n636 | 2_n1163;
assign 2_n4292 = ~(2_n8672 ^ 2_n4538);
assign 2_n5149 = 2_n12361 | 2_n5538;
assign 2_n4913 = ~2_n1512;
assign 2_n452 = 2_n5530 | 2_n2259;
assign 2_n8056 = 2_n9380 | 2_n1671;
assign 2_n3517 = 2_n5042 & 2_n125;
assign 2_n4786 = 2_n12234 ^ 2_n9814;
assign 2_n8753 = ~2_n5930;
assign 2_n4218 = 2_n5189 ^ 2_n8537;
assign 2_n6 = 2_n6577 | 2_n5540;
assign 2_n4431 = 2_n11433 | 2_n1413;
assign 2_n5751 = ~2_n12370;
assign 2_n1432 = ~2_n9499;
assign 2_n2997 = ~2_n3559;
assign 2_n7670 = 2_n11931 & 2_n10576;
assign 2_n9039 = ~(2_n12284 ^ 2_n7329);
assign 2_n8485 = 2_n3506 & 2_n2724;
assign 2_n12026 = 2_n12585 | 2_n1077;
assign 2_n2049 = ~2_n1850;
assign 2_n8627 = ~(2_n3708 ^ 2_n11253);
assign 2_n8922 = ~(2_n9611 | 2_n6178);
assign 2_n3915 = ~(2_n8321 ^ 2_n13);
assign 2_n4566 = ~(2_n9282 | 2_n5464);
assign 2_n5796 = ~(2_n5823 ^ 2_n565);
assign 2_n5187 = ~(2_n5200 ^ 2_n12395);
assign 2_n1647 = ~(2_n9806 ^ 2_n9164);
assign 2_n6906 = ~2_n11132;
assign 2_n6280 = ~(2_n7018 ^ 2_n6735);
assign 2_n11848 = ~(2_n9497 | 2_n10472);
assign 2_n9768 = 2_n8619 & 2_n2746;
assign 2_n8954 = ~2_n7882;
assign 2_n379 = ~(2_n10973 | 2_n3590);
assign 2_n10155 = ~(2_n3087 ^ 2_n511);
assign 2_n4143 = 2_n4206 & 2_n4303;
assign 2_n12040 = 2_n3096 | 2_n10903;
assign 2_n7374 = ~(2_n9605 ^ 2_n2566);
assign 2_n3930 = 2_n2099 | 2_n3924;
assign 2_n12692 = 2_n3096 | 2_n5540;
assign 2_n3446 = ~(2_n12108 ^ 2_n1818);
assign 2_n3778 = ~(2_n11926 | 2_n6362);
assign 2_n10894 = 2_n3290 & 2_n2989;
assign 2_n8428 = ~2_n9400;
assign 2_n5914 = ~2_n2507;
assign 2_n735 = 2_n11699 | 2_n6262;
assign 2_n1458 = 2_n9085 & 2_n5071;
assign 2_n4487 = 2_n2618 & 2_n1654;
assign 2_n4541 = ~(2_n6891 | 2_n8455);
assign 2_n5428 = ~(2_n8762 | 2_n12509);
assign 2_n7450 = 2_n7154 & 2_n10837;
assign 2_n471 = ~(2_n5589 ^ 2_n11291);
assign 2_n2337 = 2_n6977 | 2_n8768;
assign 2_n12436 = ~(2_n9840 ^ 2_n3238);
assign 2_n8021 = 2_n78 & 2_n1934;
assign 2_n2406 = ~2_n7285;
assign 2_n11920 = ~(2_n11942 ^ 2_n11765);
assign 2_n6146 = 2_n8026 | 2_n5540;
assign 2_n12516 = ~(2_n5757 ^ 2_n5726);
assign 2_n7310 = 2_n10750 | 2_n3924;
assign 2_n4968 = ~(2_n7743 ^ 2_n10967);
assign 2_n11996 = 2_n4515 & 2_n6220;
assign 2_n4155 = 2_n2209 ^ 2_n7039;
assign 2_n8039 = ~(2_n2279 ^ 2_n7754);
assign 2_n11511 = ~2_n9883;
assign 2_n3126 = 2_n7449 | 2_n8643;
assign 2_n5790 = ~(2_n10573 ^ 2_n6026);
assign 2_n3336 = 2_n2116 & 2_n10426;
assign 2_n9899 = ~(2_n10148 | 2_n7996);
assign 2_n8033 = 2_n11719 | 2_n1162;
assign 2_n7539 = ~(2_n5264 ^ 2_n11803);
assign 2_n11604 = 2_n6175 | 2_n8316;
assign 2_n11351 = ~(2_n5052 ^ 2_n5478);
assign 2_n4427 = 2_n5817 & 2_n2053;
assign 2_n11047 = 2_n5959 | 2_n8534;
assign 2_n1413 = ~2_n9640;
assign 2_n9587 = ~(2_n4241 ^ 2_n7699);
assign 2_n294 = ~2_n6945;
assign 2_n10728 = ~(2_n8343 ^ 2_n5706);
assign 2_n5211 = 2_n11968 | 2_n6;
assign 2_n11374 = ~2_n12734;
assign 2_n3447 = 2_n994 | 2_n7246;
assign 2_n1083 = 2_n2936 & 2_n10198;
assign 2_n9468 = 2_n11898 | 2_n1924;
assign 2_n1018 = 2_n4151 | 2_n3840;
assign 2_n3312 = ~(2_n390 ^ 2_n2483);
assign 2_n7073 = ~(2_n5714 ^ 2_n7985);
assign 2_n10610 = ~(2_n11590 ^ 2_n2778);
assign 2_n3171 = 2_n2128 & 2_n12801;
assign 2_n509 = 2_n6066 | 2_n5292;
assign 2_n9627 = ~(2_n3960 ^ 2_n6775);
assign 2_n4871 = ~(2_n12858 ^ 2_n8742);
assign 2_n8557 = 2_n2134 & 2_n6988;
assign 2_n5686 = ~(2_n8176 | 2_n2388);
assign 2_n7165 = ~(2_n8012 ^ 2_n9789);
assign 2_n617 = ~(2_n2739 ^ 2_n3369);
assign 2_n7598 = 2_n103 | 2_n7134;
assign 2_n9144 = ~2_n3754;
assign 2_n10824 = ~(2_n641 | 2_n11230);
assign 2_n8829 = 2_n2111 & 2_n7841;
assign 2_n5343 = ~(2_n10354 ^ 2_n1502);
assign 2_n3921 = ~(2_n4381 ^ 2_n26);
assign 2_n9746 = 2_n10750 | 2_n8259;
assign 2_n277 = ~(2_n3680 ^ 2_n8031);
assign 2_n2614 = ~(2_n6740 ^ 2_n9524);
assign 2_n10428 = ~(2_n505 ^ 2_n854);
assign 2_n9378 = 2_n3739 | 2_n9722;
assign 2_n3324 = ~2_n7646;
assign 2_n12351 = ~(2_n2265 ^ 2_n7026);
assign 2_n11148 = ~(2_n5874 ^ 2_n7387);
assign 2_n9610 = ~(2_n10955 ^ 2_n5648);
assign 2_n6553 = 2_n11958 | 2_n6169;
assign 2_n4916 = ~(2_n6128 | 2_n8784);
assign 2_n9391 = ~(2_n9473 ^ 2_n3292);
assign 2_n10011 = 2_n8839 & 2_n10927;
assign 2_n5647 = 2_n5203 & 2_n9780;
assign 2_n3411 = 2_n4931 & 2_n4459;
assign 2_n965 = ~2_n6008;
assign 2_n5394 = 2_n2456 | 2_n12080;
assign 2_n10691 = ~2_n12716;
assign 2_n9334 = ~(2_n8767 ^ 2_n1974);
assign 2_n178 = 2_n5355 | 2_n6524;
assign 2_n6410 = 2_n8108 & 2_n101;
assign 2_n4839 = ~2_n5159;
assign 2_n4956 = 2_n12119 | 2_n8648;
assign 2_n11556 = 2_n994 | 2_n2358;
assign 2_n11070 = ~2_n5570;
assign 2_n5312 = ~(2_n11500 | 2_n11725);
assign 2_n6265 = 2_n12217 & 2_n4608;
assign 2_n7630 = ~2_n10005;
assign 2_n4215 = ~2_n12600;
assign 2_n6761 = 2_n7729 | 2_n2303;
assign 2_n10525 = 2_n5249 & 2_n10356;
assign 2_n3037 = ~(2_n12937 | 2_n2339);
assign 2_n7519 = 2_n2336 & 2_n3775;
assign 2_n363 = ~(2_n8224 ^ 2_n6397);
assign 2_n10684 = 2_n7097 | 2_n9115;
assign 2_n559 = ~(2_n1015 ^ 2_n10240);
assign 2_n8731 = 2_n1665 & 2_n10889;
assign 2_n8070 = 2_n10157 | 2_n5258;
assign 2_n9336 = ~(2_n2565 | 2_n1322);
assign 2_n1824 = 2_n1929 | 2_n2485;
assign 2_n12897 = ~(2_n9448 ^ 2_n10248);
assign 2_n9365 = ~(2_n57 ^ 2_n9099);
assign 2_n10171 = 2_n5915 | 2_n1163;
assign 2_n2239 = ~(2_n9788 ^ 2_n362);
assign 2_n3781 = ~2_n5166;
assign 2_n10039 = ~(2_n10812 | 2_n5744);
assign 2_n3313 = 2_n8611 & 2_n9015;
assign 2_n9903 = ~(2_n9177 ^ 2_n9386);
assign 2_n8488 = ~2_n11354;
assign 2_n12259 = ~(2_n8492 ^ 2_n5296);
assign 2_n2245 = 2_n5942 | 2_n8925;
assign 2_n1273 = ~(2_n9688 ^ 2_n8446);
assign 2_n12608 = ~(2_n7957 ^ 2_n9592);
assign 2_n10390 = ~2_n6629;
assign 2_n9562 = 2_n11722 & 2_n10186;
assign 2_n1304 = ~(2_n3851 ^ 2_n11091);
assign 2_n8192 = 2_n7287 & 2_n8860;
assign 2_n6320 = 2_n5720 & 2_n6565;
assign 2_n7435 = ~2_n6583;
assign 2_n11313 = 2_n8197 | 2_n1098;
assign 2_n6876 = 2_n3768 | 2_n1611;
assign 2_n2937 = 2_n1229 & 2_n6905;
assign 2_n8161 = ~(2_n10233 | 2_n1965);
assign 2_n421 = 2_n9893 | 2_n2553;
assign 2_n3444 = ~(2_n11440 ^ 2_n8128);
assign 2_n9474 = 2_n6059 | 2_n8862;
assign 2_n3567 = 2_n2124 & 2_n3553;
assign 2_n11152 = 2_n3612 | 2_n12676;
assign 2_n5464 = ~(2_n8915 | 2_n3956);
assign 2_n8992 = ~(2_n7126 ^ 2_n5154);
assign 2_n8291 = 2_n3126 | 2_n188;
assign 2_n5294 = ~(2_n9435 ^ 2_n7535);
assign 2_n12805 = 2_n6028 & 2_n9435;
assign 2_n8164 = 2_n2866 | 2_n4742;
assign 2_n6675 = ~(2_n1992 | 2_n12212);
assign 2_n3245 = ~(2_n9301 ^ 2_n12244);
assign 2_n12083 = 2_n1083 | 2_n6613;
assign 2_n2939 = ~(2_n5559 ^ 2_n9735);
assign 2_n10325 = 2_n1444 & 2_n3951;
assign 2_n11733 = ~2_n5450;
assign 2_n10239 = 2_n2400 | 2_n2705;
assign 2_n12952 = 2_n7298 & 2_n1325;
assign 2_n153 = ~(2_n2385 ^ 2_n8884);
assign 2_n11799 = 2_n5679 | 2_n2963;
assign 2_n3660 = ~2_n9242;
assign 2_n4210 = ~(2_n10138 ^ 2_n7773);
assign 2_n627 = 2_n8535 & 2_n2410;
assign 2_n3010 = ~(2_n1461 | 2_n3374);
assign 2_n10885 = ~(2_n12766 | 2_n4704);
assign 2_n9191 = ~2_n5276;
assign 2_n11516 = ~(2_n8994 | 2_n3041);
assign 2_n8126 = ~(2_n785 | 2_n3177);
assign 2_n5256 = ~(2_n11130 ^ 2_n3871);
assign 2_n7922 = 2_n9400 & 2_n6703;
assign 2_n5054 = ~2_n4010;
assign 2_n4335 = 2_n7004 | 2_n3319;
assign 2_n10707 = ~(2_n11266 ^ 2_n8286);
assign 2_n10837 = ~(2_n6096 ^ 2_n9191);
assign 2_n65 = ~(2_n2388 ^ 2_n10264);
assign 2_n12647 = 2_n10951 | 2_n9916;
assign 2_n2411 = ~(2_n7114 ^ 2_n44);
assign 2_n11954 = ~(2_n3931 ^ 2_n8047);
assign 2_n10380 = ~(2_n12302 ^ 2_n2462);
assign 2_n4222 = 2_n11759 | 2_n6154;
assign 2_n817 = 2_n7391 | 2_n11827;
assign 2_n930 = ~(2_n3350 ^ 2_n10262);
assign 2_n9362 = ~(2_n6198 ^ 2_n12567);
assign 2_n787 = ~(2_n9689 ^ 2_n7040);
assign 2_n9418 = ~(2_n9364 | 2_n1458);
assign 2_n8939 = 2_n2660 ^ 2_n12812;
assign 2_n8230 = 2_n7378 | 2_n5188;
assign 2_n12532 = 2_n1941 | 2_n7425;
assign 2_n11424 = 2_n7192 | 2_n7696;
assign 2_n598 = ~(2_n343 ^ 2_n4062);
assign 2_n12006 = 2_n7495 | 2_n1079;
assign 2_n3919 = 2_n1937 | 2_n1413;
assign 2_n7049 = ~(2_n2560 | 2_n6965);
assign 2_n10984 = ~(2_n7870 ^ 2_n2341);
assign 2_n502 = 2_n8287 | 2_n1196;
assign 2_n4706 = 2_n11743 & 2_n12004;
assign 2_n2284 = 2_n6977 | 2_n7395;
assign 2_n1921 = ~(2_n12281 ^ 2_n4939);
assign 2_n6014 = 2_n1177 ^ 2_n1645;
assign 2_n619 = ~2_n147;
assign 2_n2501 = ~(2_n910 ^ 2_n9852);
assign 2_n1766 = 2_n9373 | 2_n9160;
assign 2_n8885 = 2_n12813 & 2_n946;
assign 2_n11415 = 2_n3746 | 2_n6197;
assign 2_n7280 = ~(2_n7225 ^ 2_n5070);
assign 2_n4633 = 2_n5168 | 2_n8997;
assign 2_n3638 = ~2_n3509;
assign 2_n2456 = ~2_n11478;
assign 2_n12204 = ~(2_n8126 ^ 2_n2692);
assign 2_n3431 = 2_n8026 | 2_n2232;
assign 2_n8416 = 2_n1699 | 2_n3924;
assign 2_n11713 = ~(2_n5843 | 2_n10236);
assign 2_n623 = ~(2_n4368 ^ 2_n7543);
assign 2_n11965 = 2_n714 | 2_n3537;
assign 2_n8923 = 2_n5219 & 2_n4926;
assign 2_n4114 = ~(2_n10165 ^ 2_n2276);
assign 2_n8895 = 2_n10683 | 2_n2527;
assign 2_n12645 = ~(2_n5290 ^ 2_n11551);
assign 2_n8661 = ~(2_n10852 ^ 2_n11134);
assign 2_n4041 = 2_n6577 | 2_n1413;
assign 2_n5540 = ~2_n7500;
assign 2_n7438 = 2_n10717 | 2_n7042;
assign 2_n11932 = ~(2_n6473 ^ 2_n1194);
assign 2_n2494 = ~(2_n140 | 2_n9737);
assign 2_n2596 = 2_n12366 | 2_n1366;
assign 2_n8597 = 2_n5024 | 2_n2044;
assign 2_n981 = ~2_n1629;
assign 2_n9611 = 2_n1834 & 2_n11175;
assign 2_n12752 = 2_n12525 | 2_n3298;
assign 2_n2444 = ~(2_n10361 | 2_n6305);
assign 2_n10260 = ~(2_n163 | 2_n1093);
assign 2_n7460 = ~(2_n1821 ^ 2_n391);
assign 2_n12232 = ~(2_n3430 ^ 2_n579);
assign 2_n645 = 2_n6847 & 2_n11002;
assign 2_n8171 = ~2_n6706;
assign 2_n3469 = 2_n7495 | 2_n11746;
assign 2_n7350 = ~(2_n1460 ^ 2_n12415);
assign 2_n8162 = 2_n12712 & 2_n9872;
assign 2_n2608 = 2_n10835 | 2_n6922;
assign 2_n11911 = 2_n4283 & 2_n5524;
assign 2_n7792 = 2_n7839 | 2_n7876;
assign 2_n4549 = 2_n2877 | 2_n572;
assign 2_n11318 = 2_n3743 | 2_n5086;
assign 2_n2136 = 2_n10157 | 2_n1047;
assign 2_n7010 = 2_n7654 | 2_n4482;
assign 2_n11339 = ~(2_n12386 ^ 2_n9257);
assign 2_n797 = ~(2_n12557 ^ 2_n1270);
assign 2_n1336 = ~(2_n12846 ^ 2_n7514);
assign 2_n5128 = ~(2_n5688 ^ 2_n10758);
assign 2_n3955 = 2_n1805 | 2_n7072;
assign 2_n12566 = ~(2_n4281 | 2_n10380);
assign 2_n5417 = 2_n4717 & 2_n12302;
assign 2_n10721 = 2_n3141 | 2_n4721;
assign 2_n1309 = 2_n9878 | 2_n6513;
assign 2_n12101 = ~(2_n3959 ^ 2_n2008);
assign 2_n5049 = 2_n10142 | 2_n9397;
assign 2_n7685 = 2_n12069 & 2_n12925;
assign 2_n8747 = ~(2_n1445 ^ 2_n3815);
assign 2_n2325 = ~2_n4597;
assign 2_n31 = ~(2_n7469 ^ 2_n6723);
assign 2_n9767 = ~(2_n12420 ^ 2_n4309);
assign 2_n11881 = 2_n11221 | 2_n3260;
assign 2_n9223 = 2_n5915 | 2_n7928;
assign 2_n4051 = ~2_n5900;
assign 2_n3430 = ~(2_n10936 ^ 2_n3631);
assign 2_n9231 = ~(2_n8803 ^ 2_n12304);
assign 2_n7582 = ~(2_n7945 | 2_n12927);
assign 2_n4455 = ~(2_n10338 ^ 2_n6123);
assign 2_n2495 = ~(2_n9951 ^ 2_n1649);
assign 2_n12726 = ~(2_n5278 | 2_n922);
assign 2_n659 = ~(2_n6157 | 2_n3657);
assign 2_n12463 = ~(2_n12505 ^ 2_n4196);
assign 2_n939 = ~(2_n2222 ^ 2_n8638);
assign 2_n12367 = ~2_n312;
assign 2_n7470 = ~2_n7248;
assign 2_n6744 = 2_n386 & 2_n9354;
assign 2_n11582 = 2_n5196 | 2_n8731;
assign 2_n716 = ~(2_n12548 ^ 2_n980);
assign 2_n8473 = ~(2_n7694 | 2_n12015);
assign 2_n8287 = ~(2_n951 ^ 2_n9151);
assign 2_n605 = 2_n8389 & 2_n11484;
assign 2_n1918 = 2_n4250 & 2_n7101;
assign 2_n3104 = 2_n8261 | 2_n12473;
assign 2_n11754 = 2_n12764 & 2_n4834;
assign 2_n4160 = 2_n3617 | 2_n8109;
assign 2_n1051 = ~2_n8276;
assign 2_n1550 = ~(2_n10504 ^ 2_n6682);
assign 2_n7593 = 2_n11142 | 2_n10187;
assign 2_n11783 = 2_n6463 & 2_n12738;
assign 2_n7133 = 2_n2099 | 2_n1932;
assign 2_n2059 = 2_n12103 | 2_n9593;
assign 2_n6620 = ~(2_n2835 ^ 2_n4033);
assign 2_n6456 = ~2_n4732;
assign 2_n4412 = ~(2_n3222 ^ 2_n12228);
assign 2_n1017 = ~(2_n10976 ^ 2_n4526);
assign 2_n3028 = ~2_n7486;
assign 2_n7017 = ~(2_n4161 ^ 2_n4888);
assign 2_n3057 = 2_n2312 & 2_n3899;
assign 2_n12103 = 2_n8818 & 2_n6967;
assign 2_n5939 = ~(2_n5947 | 2_n9539);
assign 2_n8134 = 2_n10678 & 2_n6703;
assign 2_n10491 = ~(2_n4879 ^ 2_n4157);
assign 2_n7579 = 2_n3918 ^ 2_n4922;
assign 2_n58 = 2_n11958 | 2_n7952;
assign 2_n12217 = 2_n4536 | 2_n4220;
assign 2_n12619 = 2_n21 & 2_n10600;
assign 2_n3137 = 2_n5269 & 2_n12488;
assign 2_n3654 = ~(2_n1570 ^ 2_n4680);
assign 2_n8078 = ~2_n11482;
assign 2_n3634 = 2_n8733 & 2_n5632;
assign 2_n2297 = ~2_n4490;
assign 2_n1462 = 2_n191 | 2_n561;
assign 2_n318 = 2_n11923 | 2_n4654;
assign 2_n2610 = 2_n994 | 2_n8524;
assign 2_n5154 = 2_n114 | 2_n5540;
assign 2_n5892 = ~(2_n9107 ^ 2_n2986);
assign 2_n10178 = 2_n2099 | 2_n5468;
assign 2_n6086 = 2_n636 | 2_n4818;
assign 2_n5655 = ~2_n4908;
assign 2_n10763 = 2_n1665 | 2_n10889;
assign 2_n3790 = ~(2_n7094 ^ 2_n3900);
assign 2_n1689 = 2_n12237 | 2_n8740;
assign 2_n12248 = ~(2_n9869 ^ 2_n11852);
assign 2_n11765 = ~(2_n5213 ^ 2_n6533);
assign 2_n12587 = ~2_n7827;
assign 2_n914 = ~(2_n8580 | 2_n12078);
assign 2_n2906 = 2_n636 | 2_n12535;
assign 2_n7492 = 2_n7014 & 2_n5176;
assign 2_n6671 = ~2_n10976;
assign 2_n12440 = 2_n1937 | 2_n11410;
assign 2_n5089 = 2_n2099 | 2_n12080;
assign 2_n6040 = 2_n1988 & 2_n10674;
assign 2_n2837 = 2_n12119 | 2_n12124;
assign 2_n4115 = 2_n357 & 2_n5306;
assign 2_n2661 = 2_n5954 & 2_n7486;
assign 2_n5891 = 2_n5861 | 2_n9506;
assign 2_n1313 = 2_n10339 | 2_n3224;
assign 2_n8583 = ~2_n996;
assign 2_n10021 = 2_n616 & 2_n2258;
assign 2_n6180 = 2_n5765 | 2_n5914;
assign 2_n9522 = 2_n114 | 2_n12816;
assign 2_n6513 = ~2_n12489;
assign 2_n3667 = 2_n9389 | 2_n10066;
assign 2_n3096 = ~2_n1094;
assign 2_n1761 = ~2_n2235;
assign 2_n5145 = 2_n3959 | 2_n2008;
assign 2_n9425 = 2_n9301 & 2_n2028;
assign 2_n5785 = ~(2_n3535 ^ 2_n11795);
assign 2_n3742 = 2_n12648 & 2_n11922;
assign 2_n2926 = ~(2_n6924 ^ 2_n12527);
assign 2_n6573 = ~(2_n12264 ^ 2_n11385);
assign 2_n420 = 2_n10142 | 2_n510;
assign 2_n2992 = 2_n8782 & 2_n4555;
assign 2_n12206 = ~(2_n4972 ^ 2_n12167);
assign 2_n7485 = 2_n10625 | 2_n11701;
assign 2_n10241 = 2_n413 & 2_n7955;
assign 2_n10976 = 2_n6255 & 2_n11481;
assign 2_n11180 = 2_n509 & 2_n10385;
assign 2_n6267 = 2_n2036 & 2_n2853;
assign 2_n3576 = ~(2_n12592 ^ 2_n10428);
assign 2_n3845 = 2_n8959 | 2_n995;
assign 2_n2755 = ~(2_n5730 ^ 2_n4428);
assign 2_n8568 = ~(2_n9496 ^ 2_n1775);
assign 2_n2266 = ~(2_n2104 | 2_n7321);
assign 2_n3588 = 2_n7388 & 2_n10990;
assign 2_n7749 = 2_n8397 & 2_n9700;
assign 2_n2868 = ~(2_n6759 | 2_n3694);
assign 2_n7845 = 2_n385 & 2_n6108;
assign 2_n714 = 2_n5963 & 2_n4102;
assign 2_n4664 = 2_n1822 & 2_n8375;
assign 2_n12711 = ~2_n9712;
assign 2_n11898 = 2_n6486 & 2_n1464;
assign 2_n9118 = ~(2_n11192 | 2_n1901);
assign 2_n10524 = ~(2_n8015 ^ 2_n11946);
assign 2_n3464 = 2_n752 | 2_n6114;
assign 2_n10969 = 2_n7053 | 2_n7346;
assign 2_n121 = ~(2_n11515 ^ 2_n8271);
assign 2_n8072 = 2_n2018 & 2_n10383;
assign 2_n1951 = 2_n12560 | 2_n6040;
assign 2_n1805 = 2_n8313 & 2_n879;
assign 2_n5363 = 2_n2393 & 2_n2749;
assign 2_n631 = ~(2_n7846 | 2_n4955);
assign 2_n624 = 2_n8988 & 2_n8804;
assign 2_n11699 = 2_n8836 & 2_n3941;
assign 2_n9429 = 2_n5974 & 2_n4471;
assign 2_n568 = ~2_n5053;
assign 2_n11186 = 2_n2626 & 2_n4041;
assign 2_n1554 = ~2_n11747;
assign 2_n4026 = 2_n5023 & 2_n4063;
assign 2_n9461 = ~(2_n927 | 2_n2180);
assign 2_n1869 = 2_n10601 & 2_n3576;
assign 2_n4214 = 2_n11144 | 2_n2139;
assign 2_n3179 = 2_n11222 & 2_n8433;
assign 2_n10322 = ~(2_n1365 ^ 2_n7787);
assign 2_n776 = ~(2_n1449 ^ 2_n1174);
assign 2_n1143 = 2_n8687 | 2_n12771;
assign 2_n6152 = 2_n8405 | 2_n826;
assign 2_n1219 = ~(2_n3133 | 2_n10313);
assign 2_n371 = ~2_n11370;
assign 2_n10478 = ~2_n1999;
assign 2_n7044 = 2_n9240 | 2_n11264;
assign 2_n12393 = ~(2_n5185 | 2_n5410);
assign 2_n7529 = ~(2_n97 ^ 2_n3891);
assign 2_n222 = 2_n6347 | 2_n9890;
assign 2_n3136 = ~(2_n3298 ^ 2_n5952);
assign 2_n6018 = ~(2_n697 ^ 2_n1295);
assign 2_n5674 = 2_n8757 | 2_n3021;
assign 2_n9671 = ~2_n5972;
assign 2_n1665 = ~(2_n8533 ^ 2_n6193);
assign 2_n12076 = ~(2_n8958 ^ 2_n1551);
assign 2_n3346 = 2_n1129 & 2_n4967;
assign 2_n8941 = ~(2_n8694 ^ 2_n2582);
assign 2_n5680 = ~2_n12242;
assign 2_n11513 = ~(2_n4213 ^ 2_n986);
assign 2_n7662 = 2_n11923 | 2_n3606;
assign 2_n6380 = ~(2_n6150 | 2_n5921);
assign 2_n9561 = ~2_n7146;
assign 2_n6816 = 2_n11007 & 2_n1253;
assign 2_n7858 = 2_n11623 | 2_n7632;
assign 2_n10230 = ~(2_n12906 ^ 2_n9889);
assign 2_n10244 = ~2_n2990;
assign 2_n12039 = ~2_n10051;
assign 2_n11453 = 2_n4759 & 2_n1569;
assign 2_n8518 = ~2_n2244;
assign 2_n4008 = ~(2_n3712 ^ 2_n10986);
assign 2_n7675 = ~(2_n12872 | 2_n10586);
assign 2_n3247 = 2_n11085 & 2_n486;
assign 2_n7025 = ~(2_n12493 | 2_n3785);
assign 2_n11617 = ~(2_n10863 ^ 2_n4245);
assign 2_n1543 = 2_n1399 & 2_n965;
assign 2_n293 = ~(2_n5101 ^ 2_n1178);
assign 2_n4985 = 2_n3623 | 2_n8591;
assign 2_n3694 = ~2_n10805;
assign 2_n6778 = ~(2_n6590 ^ 2_n11930);
assign 2_n6593 = ~(2_n1682 ^ 2_n9303);
assign 2_n4171 = ~(2_n3444 ^ 2_n1692);
assign 2_n6519 = 2_n7391 | 2_n6402;
assign 2_n12496 = 2_n238 | 2_n1813;
assign 2_n11155 = ~(2_n9556 ^ 2_n3043);
assign 2_n8767 = ~(2_n11436 | 2_n8632);
assign 2_n10807 = ~(2_n4116 ^ 2_n3310);
assign 2_n12163 = 2_n4187 & 2_n11728;
assign 2_n1571 = 2_n8201 & 2_n3922;
assign 2_n9813 = ~2_n1493;
assign 2_n6091 = ~2_n10012;
assign 2_n7258 = 2_n10587 | 2_n10140;
assign 2_n10150 = 2_n11138 & 2_n10218;
assign 2_n9971 = ~2_n10217;
assign 2_n6090 = 2_n11923 | 2_n795;
assign 2_n2312 = 2_n9373 | 2_n1047;
assign 2_n4301 = 2_n4911 | 2_n1079;
assign 2_n249 = 2_n7747 & 2_n6311;
assign 2_n9099 = 2_n3940 & 2_n9740;
assign 2_n6466 = 2_n3324 | 2_n2020;
assign 2_n2131 = ~(2_n6848 ^ 2_n12077);
assign 2_n8616 = ~(2_n10141 ^ 2_n2223);
assign 2_n12037 = ~(2_n10366 ^ 2_n11185);
assign 2_n2439 = 2_n3618 & 2_n3793;
assign 2_n758 = ~(2_n7234 ^ 2_n9234);
assign 2_n6374 = 2_n191 | 2_n7389;
assign 2_n2346 = 2_n5199 | 2_n3121;
assign 2_n4865 = ~(2_n9403 | 2_n11100);
assign 2_n12395 = 2_n970 & 2_n2165;
assign 2_n9698 = 2_n8870 | 2_n4818;
assign 2_n7471 = 2_n3220 & 2_n9239;
assign 2_n407 = ~(2_n10646 ^ 2_n10375);
assign 2_n6057 = ~2_n12463;
assign 2_n9290 = 2_n7283 | 2_n8859;
assign 2_n4742 = 2_n6491 & 2_n4169;
assign 2_n2304 = ~(2_n12289 ^ 2_n9253);
assign 2_n6957 = ~2_n3346;
assign 2_n2850 = 2_n5456 & 2_n87;
assign 2_n3196 = ~(2_n11807 ^ 2_n6092);
assign 2_n8913 = ~(2_n6799 ^ 2_n4772);
assign 2_n11952 = ~2_n9828;
assign 2_n9896 = 2_n7862 & 2_n5212;
assign 2_n5100 = ~(2_n2435 ^ 2_n10995);
assign 2_n1765 = 2_n8671 & 2_n9485;
assign 2_n9098 = 2_n6554 & 2_n5201;
assign 2_n12161 = ~(2_n5794 ^ 2_n4340);
assign 2_n6216 = 2_n8428 | 2_n9971;
assign 2_n8699 = ~2_n8027;
assign 2_n11670 = 2_n5601 | 2_n8237;
assign 2_n11018 = ~2_n8134;
assign 2_n4552 = 2_n7750 & 2_n8004;
assign 2_n736 = 2_n779 | 2_n456;
assign 2_n11578 = 2_n7495 | 2_n7881;
endmodule
