module top( n9 , n22 , n103 , n124 , n134 , n201 , n211 , n287 , n353 , n358 , n370 , n389 , n396 , n401 , n411 , n443 , n460 , n469 , n497 , n499 , n510 , n537 , n573 , n603 , n728 , n758 , n761 , n762 , n767 , n772 , n777 , n800 , n817 , n831 , n834 , n846 , n854 , n922 , n927 , n937 , n951 , n985 , n1007 , n1084 , n1097 , n1112 , n1165 , n1181 , n1198 , n1231 , n1302 , n1307 , n1364 , n1392 , n1401 , n1487 , n1561 , n1636 , n1650 , n1709 , n1724 , n1757 , n1806 , n1860 , n1912 , n1916 , n1937 , n1982 , n2057 , n2061 , n2068 , n2174 , n2190 , n2235 , n2252 , n2295 , n2339 , n2341 , n2458 , n2482 , n2498 , n2549 , n2590 , n2592 , n2666 , n2709 , n2737 , n2758 , n2771 , n2777 , n2805 , n2882 , n2904 , n2934 , n3006 , n3076 , n3085 , n3112 , n3130 , n3178 , n3262 , n3311 , n3323 , n3362 , n3409 , n3591 , n3641 , n3669 , n3677 , n3748 , n3769 , n3790 , n3815 , n3832 , n3946 , n4006 , n4059 , n4075 , n4114 , n4122 , n4141 , n4202 , n4330 , n4335 , n4357 , n4382 , n4419 , n4452 , n4470 , n4553 , n4743 , n4748 , n4777 , n4824 , n4862 , n4864 , n4964 , n4998 , n5003 , n5031 , n5060 , n5065 , n5167 , n5189 , n5214 , n5320 , n5356 , n5364 , n5427 , n5470 , n5536 , n5548 , n5549 , n5557 , n5568 , n5586 , n5609 , n5671 , n5684 , n5715 , n5729 , n5758 , n5801 , n5882 , n5884 , n5920 , n5962 , n5969 , n6019 , n6023 , n6085 , n6103 , n6109 , n6149 , n6168 , n6297 , n6301 , n6333 , n6392 , n6409 , n6434 , n6586 , n6655 , n6668 , n6683 , n6818 , n6826 , n6843 , n6862 , n6937 , n7034 , n7061 , n7111 , n7113 , n7132 , n7161 , n7241 , n7374 , n7411 , n7529 , n7553 , n7582 , n7659 , n7687 , n7715 , n7720 , n7729 , n7755 , n7772 , n7790 , n7812 , n7858 , n7860 , n7968 , n7974 , n8139 , n8163 , n8172 , n8183 , n8219 , n8228 , n8230 , n8233 , n8265 , n8290 , n8308 , n8332 , n8336 , n8466 , n8468 , n8506 , n8516 , n8522 , n8701 , n8716 , n8768 , n8820 , n8859 , n8860 , n8940 , n9041 , n9093 , n9100 , n9187 , n9216 , n9300 , n9329 , n9353 , n9475 , n9528 , n9531 , n9570 , n9591 , n9620 , n9669 , n9732 , n9747 , n9846 , n9866 , n9872 , n9887 , n9906 , n9915 , n10063 , n10101 , n10113 , n10122 , n10142 , n10162 , n10168 , n10243 , n10408 , n10416 , n10451 , n10453 , n10522 , n10524 , n10560 , n10594 , n10606 , n10628 , n10642 , n10657 , n10736 , n10770 , n10797 , n10805 , n10866 , n10874 , n10908 , n11030 , n11057 , n11058 , n11061 , n11077 , n11109 , n11111 , n11140 , n11147 , n11180 , n11222 , n11236 , n11252 , n11264 , n11324 , n11350 , n11396 , n11411 , n11429 , n11484 , n11488 , n11537 , n11574 , n11634 , n11665 , n11667 , n11732 , n11734 , n11778 , n11792 , n11835 , n11879 , n11882 , n11891 , n11895 , n12003 , n12059 , n12065 , n12067 , n12187 , n12263 , n12284 , n12289 , n12306 , n12334 , n12348 , n12352 , n12372 , n12406 , n12408 , n12463 , n12482 , n12503 , n12515 , n12579 , n12592 , n12605 , n12616 , n12651 , n12693 , n12750 , n12839 , n12853 , n12912 , n12965 , n12968 , n13002 , n13035 , n13058 , n13060 , n13201 );
    input n9 , n22 , n103 , n124 , n287 , n353 , n389 , n401 , n411 , n443 , n469 , n497 , n499 , n510 , n603 , n761 , n767 , n772 , n817 , n834 , n854 , n937 , n951 , n1007 , n1084 , n1165 , n1198 , n1231 , n1302 , n1307 , n1364 , n1392 , n1636 , n1650 , n1709 , n1724 , n1757 , n1912 , n1916 , n1982 , n2057 , n2068 , n2174 , n2252 , n2295 , n2339 , n2341 , n2458 , n2482 , n2498 , n2590 , n2592 , n2666 , n2737 , n2758 , n2771 , n2777 , n2882 , n3006 , n3076 , n3085 , n3112 , n3130 , n3178 , n3311 , n3409 , n3591 , n3641 , n3669 , n3677 , n3769 , n3815 , n3832 , n4006 , n4075 , n4114 , n4122 , n4141 , n4330 , n4335 , n4357 , n4382 , n4419 , n4452 , n4470 , n4743 , n4748 , n4862 , n4964 , n4998 , n5031 , n5065 , n5167 , n5189 , n5214 , n5320 , n5356 , n5427 , n5470 , n5536 , n5548 , n5568 , n5586 , n5671 , n5684 , n5715 , n5729 , n5758 , n5801 , n5884 , n5920 , n5962 , n5969 , n6023 , n6085 , n6149 , n6168 , n6333 , n6392 , n6409 , n6655 , n6668 , n6818 , n6826 , n6843 , n6937 , n7061 , n7113 , n7161 , n7374 , n7411 , n7529 , n7659 , n7715 , n7720 , n7729 , n7772 , n7812 , n7974 , n8139 , n8163 , n8183 , n8228 , n8230 , n8233 , n8290 , n8308 , n8332 , n8466 , n8468 , n8506 , n8522 , n8716 , n8768 , n8820 , n8859 , n8860 , n8940 , n9041 , n9093 , n9187 , n9216 , n9300 , n9353 , n9475 , n9528 , n9531 , n9570 , n9591 , n9620 , n9669 , n9732 , n9747 , n9846 , n9887 , n9906 , n9915 , n10063 , n10113 , n10122 , n10142 , n10162 , n10168 , n10408 , n10416 , n10451 , n10522 , n10560 , n10594 , n10606 , n10642 , n10657 , n10770 , n10805 , n10866 , n10874 , n10908 , n11030 , n11058 , n11061 , n11109 , n11111 , n11180 , n11222 , n11236 , n11324 , n11350 , n11396 , n11411 , n11429 , n11488 , n11537 , n11574 , n11634 , n11665 , n11734 , n11835 , n11891 , n12003 , n12065 , n12263 , n12284 , n12289 , n12306 , n12348 , n12352 , n12372 , n12408 , n12482 , n12579 , n12592 , n12605 , n12651 , n12693 , n12750 , n12853 , n12912 , n12965 , n13058 , n13060 , n13201 ;
    output n134 , n201 , n211 , n358 , n370 , n396 , n460 , n537 , n573 , n728 , n758 , n762 , n777 , n800 , n831 , n846 , n922 , n927 , n985 , n1097 , n1112 , n1181 , n1401 , n1487 , n1561 , n1806 , n1860 , n1937 , n2061 , n2190 , n2235 , n2549 , n2709 , n2805 , n2904 , n2934 , n3262 , n3323 , n3362 , n3748 , n3790 , n3946 , n4059 , n4202 , n4553 , n4777 , n4824 , n4864 , n5003 , n5060 , n5364 , n5549 , n5557 , n5609 , n5882 , n6019 , n6103 , n6109 , n6297 , n6301 , n6434 , n6586 , n6683 , n6862 , n7034 , n7111 , n7132 , n7241 , n7553 , n7582 , n7687 , n7755 , n7790 , n7858 , n7860 , n7968 , n8172 , n8219 , n8265 , n8336 , n8516 , n8701 , n9100 , n9329 , n9866 , n9872 , n10101 , n10243 , n10453 , n10524 , n10628 , n10736 , n10797 , n11057 , n11077 , n11140 , n11147 , n11252 , n11264 , n11484 , n11667 , n11732 , n11778 , n11792 , n11879 , n11882 , n11895 , n12059 , n12067 , n12187 , n12334 , n12406 , n12463 , n12503 , n12515 , n12616 , n12839 , n12968 , n13002 , n13035 ;
    wire n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n354 , n355 , n356 , n357 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n390 , n391 , n392 , n393 , n394 , n395 , n397 , n398 , n399 , n400 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n498 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n759 , n760 , n763 , n764 , n765 , n766 , n768 , n769 , n770 , n771 , n773 , n774 , n775 , n776 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n832 , n833 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n923 , n924 , n925 , n926 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1303 , n1304 , n1305 , n1306 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1913 , n1914 , n1915 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2058 , n2059 , n2060 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2340 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2591 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2772 , n2773 , n2774 , n2775 , n2776 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4331 , n4332 , n4333 , n4334 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4744 , n4745 , n4746 , n4747 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4863 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4999 , n5000 , n5001 , n5002 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5061 , n5062 , n5063 , n5064 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5883 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6020 , n6021 , n6022 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6104 , n6105 , n6106 , n6107 , n6108 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6298 , n6299 , n6300 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7112 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7716 , n7717 , n7718 , n7719 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7859 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7969 , n7970 , n7971 , n7972 , n7973 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8229 , n8231 , n8232 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8333 , n8334 , n8335 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8467 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8517 , n8518 , n8519 , n8520 , n8521 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9529 , n9530 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9867 , n9868 , n9869 , n9870 , n9871 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10163 , n10164 , n10165 , n10166 , n10167 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , n10452 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10523 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11059 , n11060 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11110 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11485 , n11486 , n11487 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11666 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11733 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11791 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11880 , n11881 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11892 , n11893 , n11894 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12060 , n12061 , n12062 , n12063 , n12064 , n12066 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12285 , n12286 , n12287 , n12288 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12349 , n12350 , n12351 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12407 , n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , n12481 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , n12516 , n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , n12591 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , n12606 , n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , n12851 , n12852 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , n12911 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , n12929 , n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , n12947 , n12948 , n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , n12960 , n12961 , n12962 , n12963 , n12964 , n12966 , n12967 , n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , n12988 , n12989 , n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , n12999 , n13000 , n13001 , n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , n13009 , n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , n13036 , n13037 , n13038 , n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , n13049 , n13050 , n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , n13057 , n13059 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , n13109 , n13110 , n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , n13117 , n13118 , n13119 , n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , n13130 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , n13199 , n13200 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , n13219 , n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , n13240 , n13241 , n13242 , n13243 ;
assign n3523 = n7151 & n6767;
assign n1818 = ~(n11618 ^ n10125);
assign n6666 = n1354 | n6635;
assign n13003 = n10781 | n8348;
assign n8017 = n995 | n12970;
assign n9879 = n4074 & n12255;
assign n849 = ~(n1713 ^ n1158);
assign n837 = ~(n3701 | n2651);
assign n3470 = ~(n12726 ^ n4668);
assign n6673 = ~(n2914 ^ n655);
assign n8353 = ~(n3258 ^ n2954);
assign n1644 = n7660 | n10173;
assign n4458 = ~(n11074 ^ n9291);
assign n4154 = n12552 | n10871;
assign n5448 = ~n13203;
assign n938 = n2711 | n11144;
assign n9174 = ~n72;
assign n6954 = n3044 | n11894;
assign n224 = ~(n10835 ^ n2683);
assign n7171 = ~n2309;
assign n1343 = ~(n8789 | n7265);
assign n3099 = ~n5324;
assign n12128 = ~n5568;
assign n12514 = ~(n5673 | n13166);
assign n5497 = n10761 | n6732;
assign n6006 = n3747 & n4857;
assign n8827 = ~(n6431 ^ n7145);
assign n9763 = n7126 & n2227;
assign n11908 = n4316 | n2924;
assign n2161 = ~(n11270 ^ n1874);
assign n618 = ~(n7815 ^ n4460);
assign n1422 = ~n12965;
assign n9158 = ~(n601 ^ n9373);
assign n9135 = n1550 | n2209;
assign n12910 = n1958 & n4654;
assign n13069 = n10439 | n12388;
assign n13000 = ~(n4381 ^ n10298);
assign n12582 = ~(n1459 ^ n1950);
assign n1273 = ~(n8182 ^ n8861);
assign n11174 = ~n485;
assign n5045 = ~n5586;
assign n7486 = n6079 | n4448;
assign n9434 = n6006 | n9735;
assign n6268 = n7700 | n1026;
assign n11498 = n6991 | n11644;
assign n1005 = ~n10373;
assign n10206 = ~n6964;
assign n746 = ~(n4418 ^ n496);
assign n12707 = n7675 | n1144;
assign n11383 = n5865 | n5242;
assign n12636 = ~n9701;
assign n6506 = ~n3311;
assign n5217 = n7939 | n1337;
assign n6028 = ~n12482;
assign n7328 = ~(n6204 ^ n12282);
assign n3430 = n12568 | n12847;
assign n13217 = ~(n8937 ^ n9105);
assign n7035 = ~(n3487 ^ n1164);
assign n11295 = n10032 | n7254;
assign n734 = ~n11411;
assign n11278 = ~(n9811 ^ n9427);
assign n10946 = ~(n12215 ^ n3738);
assign n610 = ~(n10055 ^ n774);
assign n10496 = ~(n10728 ^ n13055);
assign n12601 = ~(n3959 ^ n9631);
assign n10620 = n6939 | n9159;
assign n5216 = ~n1426;
assign n3802 = ~(n596 ^ n1088);
assign n12895 = n13027 | n10662;
assign n11521 = ~n9732;
assign n4884 = ~n3670;
assign n9741 = ~n8078;
assign n1826 = n6083 ^ n7616;
assign n3658 = ~(n12111 ^ n4323);
assign n6851 = n11030 & n12289;
assign n10227 = ~(n10752 ^ n594);
assign n11559 = n6226 ^ n4888;
assign n127 = n10882 | n11551;
assign n8256 = n7819 | n10043;
assign n10029 = n8852;
assign n4473 = ~n2295;
assign n10956 = ~n5729;
assign n3456 = ~n11682;
assign n9718 = ~n6670;
assign n7609 = n8188 | n4490;
assign n10187 = ~(n330 | n12782);
assign n5538 = n4081 & n9186;
assign n1464 = ~(n520 ^ n7499);
assign n9928 = ~(n4616 ^ n9260);
assign n1570 = n12471;
assign n1525 = ~(n8885 ^ n10490);
assign n3435 = n3669 & n834;
assign n11902 = n2848 | n12501;
assign n2414 = n4258 | n10106;
assign n252 = n10338 & n6627;
assign n9289 = n1168 | n7723;
assign n12010 = n5480 | n2796;
assign n13046 = ~(n6622 ^ n10271);
assign n12280 = n683 | n9080;
assign n7727 = n7912 | n13118;
assign n8096 = ~(n8582 ^ n10826);
assign n9186 = n5455 | n4724;
assign n4933 = ~(n5944 ^ n5560);
assign n7994 = ~(n2528 ^ n8607);
assign n10128 = ~n11891;
assign n1597 = n3186 | n3500;
assign n12870 = ~(n1824 | n10842);
assign n11470 = n1782 & n10313;
assign n5626 = ~n7556;
assign n5131 = ~(n7739 ^ n3051);
assign n425 = n1907 & n9672;
assign n7539 = ~(n9415 ^ n9935);
assign n3425 = n10761 | n8702;
assign n8270 = ~(n465 ^ n727);
assign n12783 = n7695 & n9404;
assign n3269 = ~(n6985 ^ n12644);
assign n12026 = n3006 & n6149;
assign n12042 = ~n10925;
assign n9682 = ~n11324;
assign n10094 = n4795 & n8792;
assign n8499 = ~n10451;
assign n12046 = n10812 | n2937;
assign n2932 = ~(n4047 ^ n10504);
assign n3026 = n3135 & n5808;
assign n12849 = n8207 & n1545;
assign n4076 = ~(n12132 ^ n965);
assign n7769 = n7041 | n12695;
assign n11615 = ~(n1868 ^ n639);
assign n12282 = ~(n6713 ^ n6848);
assign n4146 = n8868 | n2958;
assign n12518 = ~n2646;
assign n4928 = n2430 & n13186;
assign n2372 = ~(n8740 ^ n9673);
assign n1964 = ~(n12106 ^ n11044);
assign n2158 = n5607 | n9431;
assign n12165 = n12737 | n5956;
assign n9096 = n11398 & n5467;
assign n6181 = n5378 & n7277;
assign n10765 = ~(n5090 ^ n5825);
assign n10235 = n7933 | n7244;
assign n10691 = n4755 | n10289;
assign n11500 = ~(n7563 ^ n3718);
assign n2741 = ~(n10187 ^ n4817);
assign n12881 = ~n4470;
assign n8882 = n48 | n4947;
assign n12252 = n5759 & n664;
assign n11017 = ~(n5932 ^ n284);
assign n8688 = n2580 | n7533;
assign n6625 = n7931 | n11255;
assign n7215 = n11183 | n7859;
assign n10018 = ~n8468;
assign n3622 = n8063 & n3371;
assign n11049 = ~(n2108 ^ n7715);
assign n7369 = ~(n2074 | n6239);
assign n7264 = ~(n3499 ^ n5493);
assign n15 = ~(n2867 | n11302);
assign n6977 = n7625 & n3577;
assign n1657 = ~(n1414 ^ n11594);
assign n8071 = n11471 & n3006;
assign n8822 = n2106 & n10607;
assign n8482 = ~(n8706 ^ n9916);
assign n6836 = n6039 & n5862;
assign n8910 = ~(n745 | n1899);
assign n6581 = ~n12682;
assign n4969 = n264 & n10423;
assign n4875 = ~n1198;
assign n7723 = n10879;
assign n4889 = n10680 & n4121;
assign n1511 = ~n12263;
assign n10200 = n5671 & n8233;
assign n9518 = n6162 & n8361;
assign n3167 = ~n2840;
assign n12055 = n9429 | n12501;
assign n3747 = ~(n8035 ^ n9201);
assign n1459 = ~(n1525 ^ n4142);
assign n7157 = ~(n2593 ^ n8114);
assign n2025 = n4595 | n11343;
assign n8315 = ~n772;
assign n5117 = n8183 & n10606;
assign n10969 = ~(n2741 ^ n7724);
assign n9023 = n1365 | n11162;
assign n11207 = ~(n4982 ^ n12583);
assign n8844 = ~(n9406 ^ n3154);
assign n5897 = ~(n405 ^ n1808);
assign n9959 = n5670 | n10135;
assign n5651 = ~(n3346 ^ n1154);
assign n2272 = n965 | n7619;
assign n12545 = ~(n6303 ^ n2855);
assign n6019 = ~(n1466 ^ n5895);
assign n7748 = ~n772;
assign n1773 = n5605 | n5868;
assign n5741 = ~(n123 ^ n5069);
assign n8776 = ~n401;
assign n6970 = n7597 | n6265;
assign n7467 = ~(n2424 ^ n5326);
assign n1797 = n11535 & n8925;
assign n663 = ~n12379;
assign n3064 = ~(n4914 ^ n10942);
assign n3127 = ~n6818;
assign n5021 = n11125 | n998;
assign n7406 = ~(n13149 ^ n9556);
assign n7055 = ~n10418;
assign n5403 = ~(n9797 ^ n1532);
assign n8895 = ~(n4557 ^ n11784);
assign n12945 = ~(n681 | n8347);
assign n6336 = n6743 | n4936;
assign n9803 = n59 | n5406;
assign n8253 = n10998 & n11890;
assign n1039 = ~n224;
assign n12475 = n7125 & n12365;
assign n1123 = ~(n11737 ^ n2953);
assign n4878 = n3122 | n10100;
assign n12483 = ~n12853;
assign n11066 = ~(n9898 ^ n2);
assign n9060 = n454 | n2192;
assign n6801 = ~(n2647 ^ n58);
assign n11464 = n4808 | n2133;
assign n56 = ~n12893;
assign n3394 = n2109 | n2232;
assign n8591 = ~(n5698 ^ n3242);
assign n12397 = n2986 & n1262;
assign n5936 = n11482 | n8822;
assign n12536 = n3346 | n10828;
assign n182 = n7840 & n12178;
assign n5374 = n8977 | n6404;
assign n5665 = n5260 | n7302;
assign n6797 = n1329 | n12847;
assign n11384 = n10300 & n5027;
assign n544 = ~n7328;
assign n9948 = n13239 & n826;
assign n7302 = ~(n972 | n10692);
assign n12985 = ~(n12564 ^ n295);
assign n6934 = n4842 | n1686;
assign n10213 = ~n11488;
assign n4065 = ~(n9986 ^ n9694);
assign n4118 = ~(n4117 | n3250);
assign n548 = ~(n3150 ^ n6695);
assign n11717 = n850 | n6339;
assign n10634 = ~(n641 ^ n12418);
assign n2885 = ~(n8464 ^ n9392);
assign n7889 = n6250 | n479;
assign n10884 = n5639 & n7441;
assign n4336 = n6699 | n9784;
assign n7686 = ~(n4311 ^ n7280);
assign n4585 = n6714 & n12135;
assign n5941 = ~(n7983 ^ n10957);
assign n2699 = ~(n2064 ^ n6719);
assign n1667 = n12621 | n12695;
assign n1128 = n5597 | n5846;
assign n7241 = ~(n1858 ^ n8884);
assign n4706 = n7207 | n6789;
assign n12100 = ~(n8789 ^ n11047);
assign n1720 = ~n854;
assign n1727 = n7903 | n12768;
assign n2694 = n3859 & n10391;
assign n11269 = n10950 | n7723;
assign n12665 = n3311 & n854;
assign n9038 = ~(n4915 ^ n11245);
assign n7103 = n8280 ^ n7205;
assign n11224 = ~(n1700 ^ n6224);
assign n10194 = ~(n7726 ^ n9611);
assign n8063 = n7571 | n9749;
assign n9003 = n1986 | n5515;
assign n2603 = ~(n11198 ^ n9001);
assign n12041 = ~(n12652 | n12699);
assign n10243 = ~(n9664 ^ n5837);
assign n8126 = ~(n3976 | n3723);
assign n509 = ~(n11533 ^ n8434);
assign n926 = ~(n10067 | n11759);
assign n3428 = ~n772;
assign n6790 = n10770 & n8290;
assign n7120 = ~(n10782 ^ n12379);
assign n1432 = n10770 & n8506;
assign n3993 = ~(n3936 | n4810);
assign n8434 = n10287 | n4724;
assign n10369 = n2036 & n2434;
assign n2820 = ~(n5750 ^ n5873);
assign n11906 = ~(n11583 ^ n11939);
assign n10844 = ~(n6507 | n5848);
assign n5991 = ~(n11605 ^ n3565);
assign n3182 = ~(n12290 ^ n207);
assign n1127 = n6084 & n8061;
assign n8535 = ~(n7139 ^ n886);
assign n6715 = n8625 & n9970;
assign n12405 = ~(n9026 ^ n1435);
assign n12489 = n869 & n11564;
assign n10275 = n12829 | n6461;
assign n6766 = ~(n10996 | n12420);
assign n895 = n11793 | n4354;
assign n6200 = ~(n1966 ^ n3658);
assign n5125 = n7216 | n4947;
assign n8232 = n2916 & n4466;
assign n3698 = ~n3085;
assign n9623 = n4884 & n1116;
assign n5759 = ~(n11271 ^ n1944);
assign n7298 = n12955 | n8360;
assign n13065 = ~(n11051 ^ n5718);
assign n4814 = n3158 | n2133;
assign n12076 = n10448 | n11101;
assign n3499 = n9170 & n4661;
assign n7258 = ~n966;
assign n5466 = ~n9831;
assign n9354 = n6964 | n1211;
assign n684 = n156 & n2342;
assign n13035 = ~(n680 ^ n2364);
assign n1952 = n10369 | n12854;
assign n7505 = n9975 & n5700;
assign n1378 = ~(n7408 ^ n893);
assign n3432 = ~(n4910 | n2820);
assign n7681 = n11391 & n516;
assign n1009 = ~(n4594 ^ n11293);
assign n11528 = ~(n12916 ^ n2735);
assign n5451 = n3049 | n11137;
assign n870 = ~(n5330 ^ n8870);
assign n11889 = n11092 | n8712;
assign n274 = ~(n10086 | n1322);
assign n1816 = ~(n5099 | n364);
assign n8711 = n3488 & n5835;
assign n8045 = ~(n11306 ^ n1909);
assign n5854 = ~n9654;
assign n4148 = n6718 & n8567;
assign n6276 = ~n7969;
assign n2215 = ~n10264;
assign n10363 = n2785 | n10802;
assign n3736 = n4029 | n12800;
assign n392 = ~n10805;
assign n1523 = ~(n8333 ^ n2906);
assign n5909 = n11344 | n9480;
assign n9058 = ~(n7915 ^ n4106);
assign n6101 = ~n6080;
assign n4479 = n1320 | n4237;
assign n1323 = ~n9887;
assign n2727 = n7455 | n7734;
assign n3146 = n1527 & n6961;
assign n8865 = ~(n4591 | n1885);
assign n3829 = ~n6124;
assign n3233 = ~(n11991 ^ n7273);
assign n8698 = ~(n11223 ^ n9998);
assign n11480 = ~(n9789 ^ n5206);
assign n4666 = n8675 | n7127;
assign n6098 = n7657 | n11608;
assign n3812 = n1475 | n1714;
assign n10472 = ~(n13151 ^ n5156);
assign n2397 = ~(n8743 ^ n408);
assign n4537 = ~n10866;
assign n7474 = n5126 & n7225;
assign n7175 = ~(n4591 ^ n9284);
assign n10810 = n17 & n11460;
assign n6935 = ~(n3991 ^ n12749);
assign n2867 = ~(n8207 | n1545);
assign n12294 = n560 | n7530;
assign n5141 = n10109 | n62;
assign n5614 = n8289 & n5294;
assign n11789 = ~(n996 ^ n11902);
assign n8977 = ~n1650;
assign n8289 = ~(n4193 ^ n12634);
assign n230 = n7395 | n8535;
assign n3147 = ~(n10089 ^ n6641);
assign n3582 = n8074 | n7668;
assign n3248 = n8976 & n13179;
assign n5393 = ~(n513 ^ n651);
assign n4574 = n6295 | n12188;
assign n12391 = ~n6155;
assign n533 = ~(n6504 | n9459);
assign n51 = n3260 | n10823;
assign n10044 = n6949 | n7524;
assign n8003 = ~(n8072 ^ n4549);
assign n2402 = ~(n10052 ^ n10264);
assign n1561 = ~(n11576 ^ n12742);
assign n2185 = n11102 ^ n12014;
assign n8205 = ~(n5664 ^ n3556);
assign n5438 = n694 | n6635;
assign n11137 = ~n9475;
assign n4718 = ~(n7818 ^ n7274);
assign n2290 = n10375 & n1128;
assign n9296 = ~n5770;
assign n2386 = ~n5136;
assign n1843 = n2767 & n10584;
assign n9720 = ~n7330;
assign n855 = ~n11473;
assign n332 = n67 & n2774;
assign n10445 = n13234 & n2257;
assign n1752 = ~(n10102 ^ n11894);
assign n12259 = n4272 | n12847;
assign n429 = ~(n13177 ^ n2844);
assign n9627 = ~(n9654 | n11323);
assign n3695 = n13082 | n12273;
assign n2591 = n7718 | n5242;
assign n90 = n8339 & n8542;
assign n1663 = ~n8137;
assign n8095 = ~(n12747 | n10337);
assign n7881 = ~(n12896 | n3312);
assign n10569 = ~(n12468 ^ n1255);
assign n7775 = ~(n1632 | n12013);
assign n1531 = ~(n13132 | n3777);
assign n9569 = ~n4712;
assign n6228 = n761 & n834;
assign n3946 = ~(n11968 ^ n12523);
assign n9352 = n4745 & n12411;
assign n2675 = n5045;
assign n9577 = n2486 ^ n11084;
assign n6099 = ~n287;
assign n4341 = ~(n4533 ^ n12320);
assign n1594 = n3613 | n9130;
assign n8671 = ~n5800;
assign n6873 = n10501 | n12959;
assign n178 = n10343 | n9182;
assign n13113 = n3453 & n5335;
assign n11699 = ~(n9176 ^ n3054);
assign n6311 = ~(n3400 ^ n1203);
assign n11801 = n1406 | n8534;
assign n7251 = n4994 & n10077;
assign n12189 = n2853 & n2854;
assign n5069 = n2850 & n8526;
assign n1955 = n3068 | n6732;
assign n5377 = ~n10405;
assign n4152 = ~n3918;
assign n6769 = n9272;
assign n5399 = n3607 & n8996;
assign n2997 = ~(n4593 | n6096);
assign n10914 = n3415 & n11558;
assign n2496 = ~(n5094 ^ n7517);
assign n11981 = n7543 & n931;
assign n739 = n9793 | n12789;
assign n3519 = n2107 & n8548;
assign n1193 = ~n11325;
assign n12300 = n1213 | n7682;
assign n5727 = ~(n11867 ^ n421);
assign n11662 = n1735 | n10674;
assign n11301 = ~(n6653 | n7490);
assign n7195 = n4016 | n4095;
assign n1514 = n1090 | n1292;
assign n2389 = ~(n2023 ^ n5824);
assign n2911 = ~(n10278 | n1441);
assign n8704 = n2615 | n2871;
assign n5375 = ~n7877;
assign n2898 = ~(n4861 ^ n8377);
assign n4381 = ~(n3291 ^ n3601);
assign n7605 = n12568 | n12273;
assign n4105 = n4539 | n11234;
assign n3697 = ~(n7549 | n2597);
assign n463 = ~(n3247 ^ n3560);
assign n2596 = n8613 | n7312;
assign n2478 = ~n11468;
assign n13056 = n6489 ^ n2342;
assign n2996 = n1375 & n12097;
assign n9031 = ~(n377 ^ n10083);
assign n3689 = ~(n5030 | n12908);
assign n4506 = n4044 | n12672;
assign n1419 = n3534 | n4947;
assign n8101 = n2609 & n5342;
assign n3043 = ~(n6049 ^ n8427);
assign n5126 = ~(n10506 ^ n10151);
assign n3081 = ~(n12492 ^ n7263);
assign n11804 = ~(n7304 | n11649);
assign n3982 = n9882 | n4373;
assign n2457 = n4001 ^ n9692;
assign n3511 = ~(n10667 ^ n11474);
assign n4502 = ~(n7870 | n5043);
assign n1971 = n6668 & n12853;
assign n399 = n3544 | n1702;
assign n9564 = n7095 & n4211;
assign n6266 = ~(n10405 | n608);
assign n12834 = ~n5758;
assign n9321 = ~n5094;
assign n5198 = ~(n2237 | n9953);
assign n12272 = ~n983;
assign n7857 = n4004 | n9549;
assign n7666 = ~(n3916 ^ n4907);
assign n1115 = ~(n5410 ^ n2779);
assign n5408 = ~(n3985 ^ n885);
assign n10498 = n10013 ^ n12578;
assign n6375 = ~n469;
assign n3083 = n10188 | n3963;
assign n10718 = ~(n10888 ^ n4826);
assign n8854 = ~(n11573 ^ n9844);
assign n210 = n1934 & n1234;
assign n11453 = n4467 | n12142;
assign n11636 = n6355 | n3890;
assign n10322 = n4382 & n1636;
assign n292 = n13229 & n7849;
assign n9220 = n5005 & n13110;
assign n1930 = ~n7374;
assign n9271 = ~(n1880 ^ n6551);
assign n4672 = ~(n10482 ^ n4254);
assign n2409 = n8661 & n5568;
assign n10371 = ~(n10940 ^ n5821);
assign n9032 = n78 & n116;
assign n7027 = ~(n11092 ^ n8712);
assign n7525 = ~(n5996 ^ n6844);
assign n6474 = n1514 & n8318;
assign n7432 = n241 | n9070;
assign n10678 = n3299 | n7741;
assign n2549 = ~(n4889 ^ n1122);
assign n2497 = ~(n2176 ^ n10951);
assign n6026 = ~(n12553 ^ n4350);
assign n6046 = ~n11830;
assign n1271 = ~n972;
assign n3381 = ~(n10378 | n4249);
assign n11526 = ~(n11658 ^ n5101);
assign n5339 = ~(n6859 ^ n4823);
assign n933 = n2263 & n1443;
assign n10111 = n12972 & n3927;
assign n3969 = ~(n988 ^ n4873);
assign n3765 = ~(n3214 ^ n7173);
assign n2361 = n1175 & n8084;
assign n4052 = ~(n10931 ^ n13164);
assign n6662 = ~(n6515 ^ n8755);
assign n765 = ~n9;
assign n6541 = n13109 & n12435;
assign n9259 = n5545 & n2025;
assign n9554 = ~(n2044 ^ n13048);
assign n11395 = n11331 & n2881;
assign n11489 = n5440 | n2244;
assign n8091 = n3047 | n12273;
assign n8203 = ~(n5798 ^ n6252);
assign n6681 = ~(n3205 ^ n9751);
assign n8349 = n8206 | n2059;
assign n7052 = ~n8253;
assign n7594 = ~(n3504 | n13045);
assign n12464 = ~(n12628 | n5484);
assign n5388 = ~(n9095 | n3813);
assign n4931 = ~(n12021 ^ n6893);
assign n10179 = n2623;
assign n2164 = ~(n228 ^ n6127);
assign n7297 = n12050 | n4899;
assign n2307 = ~n3496;
assign n1474 = n2247 & n12928;
assign n12274 = n3099 | n3074;
assign n4948 = ~(n5561 ^ n2060);
assign n9880 = n9722 | n9974;
assign n8188 = ~n761;
assign n1910 = n2425 & n2380;
assign n1330 = ~(n4977 ^ n1221);
assign n6567 = ~(n2732 | n11081);
assign n5706 = ~(n3305 ^ n9368);
assign n8665 = ~n4743;
assign n6879 = n1059 & n6856;
assign n5417 = ~(n4427 | n5663);
assign n2569 = n11617 & n11630;
assign n150 = n10943 | n6511;
assign n5642 = ~(n1143 ^ n6994);
assign n2342 = n1364 & n3815;
assign n10507 = n7669 | n9101;
assign n5389 = n10253 ^ n12182;
assign n13198 = ~n4337;
assign n8336 = ~(n7491 ^ n1362);
assign n11164 = n4625 & n9331;
assign n9237 = n8386 | n615;
assign n6491 = n9702 | n1571;
assign n8204 = n228 & n2829;
assign n1520 = n1270 | n6903;
assign n11777 = ~(n13180 ^ n3624);
assign n2242 = ~(n2014 ^ n13224);
assign n11936 = ~(n9678 ^ n9999);
assign n3480 = n2156 & n7971;
assign n3327 = n8653 & n2808;
assign n986 = ~(n6761 | n2571);
assign n649 = n1769 & n12117;
assign n10528 = ~(n5421 | n9376);
assign n5825 = ~(n7638 ^ n3728);
assign n7667 = n12246 & n888;
assign n5062 = ~(n10288 ^ n1014);
assign n809 = n10434 | n12723;
assign n2516 = n12930 | n1144;
assign n12791 = n10558 | n12273;
assign n5917 = ~n1707;
assign n10134 = n11635 & n2482;
assign n3524 = ~n4574;
assign n4204 = n5842 | n10761;
assign n10913 = ~(n8382 ^ n4813);
assign n9727 = n4275 | n9842;
assign n501 = ~(n11461 ^ n2444);
assign n3544 = n13218 & n9420;
assign n3000 = n10097 & n12071;
assign n379 = ~n5536;
assign n12648 = ~n1982;
assign n107 = ~n10537;
assign n11887 = ~n4479;
assign n1666 = ~(n10902 ^ n12198);
assign n9122 = n12324 | n2133;
assign n3828 = n8077 & n9720;
assign n2725 = ~n4688;
assign n3496 = ~(n5593 ^ n5055);
assign n10149 = n12832 ^ n1174;
assign n5725 = n3352 ^ n3435;
assign n8495 = n12643 & n11888;
assign n10348 = ~(n535 ^ n7178);
assign n1388 = ~n9428;
assign n5130 = n3928 | n1985;
assign n2031 = ~(n11266 ^ n3774);
assign n5562 = ~n10408;
assign n3645 = n10416 & n12306;
assign n12119 = n9323 | n1797;
assign n3302 = n1919 | n4373;
assign n10622 = ~(n10688 ^ n9990);
assign n6263 = ~(n2363 ^ n11420);
assign n39 = ~n4240;
assign n2081 = ~n9794;
assign n3477 = n12563 | n4949;
assign n4950 = n7457 & n3117;
assign n1220 = n5583 | n6017;
assign n1176 = n10037 | n4373;
assign n502 = ~(n4486 ^ n8345);
assign n5047 = n1208 & n7264;
assign n45 = ~n1084;
assign n9656 = n5297 | n11619;
assign n5033 = n3752 & n6153;
assign n2712 = n2849 | n2793;
assign n11275 = n5058 & n1922;
assign n13171 = ~(n9972 ^ n9555);
assign n672 = ~n192;
assign n9274 = ~(n8133 ^ n3302);
assign n11590 = ~(n11954 ^ n12210);
assign n11495 = n60 & n5230;
assign n2905 = ~(n5034 | n4222);
assign n5159 = ~(n1062 ^ n3947);
assign n9641 = ~n988;
assign n7598 = n11987 | n3019;
assign n2616 = ~(n5929 | n10215);
assign n188 = n9059 | n4089;
assign n9469 = ~(n5736 ^ n3986);
assign n6938 = n2024 & n6508;
assign n1448 = n1263 | n4058;
assign n3772 = n10189 & n7743;
assign n11589 = ~(n87 ^ n7373);
assign n1943 = n6583 & n7231;
assign n12342 = n6816 | n4551;
assign n10636 = ~n7845;
assign n5678 = ~(n2644 ^ n6709);
assign n4456 = n11449 | n8348;
assign n4644 = n10603 & n6540;
assign n7554 = ~(n7099 ^ n2620);
assign n459 = ~(n9851 ^ n5144);
assign n7349 = ~(n7484 | n3848);
assign n11018 = ~n4006;
assign n12926 = ~n12867;
assign n7704 = n7232 & n8733;
assign n6699 = ~n5189;
assign n3956 = n2289 | n3538;
assign n10422 = n2457 | n8964;
assign n4266 = ~(n12250 | n8692);
assign n3169 = ~n10908;
assign n6909 = n518 & n7776;
assign n10542 = ~(n5695 ^ n7339);
assign n1094 = ~n5244;
assign n4697 = ~(n12184 | n10030);
assign n9731 = n1360 | n3972;
assign n12155 = n6177 & n5857;
assign n594 = ~(n13187 ^ n12641);
assign n10143 = ~n9570;
assign n11515 = n2246 | n6145;
assign n3713 = ~(n6058 ^ n2976);
assign n13109 = n1131 | n1153;
assign n2260 = ~(n3272 | n12869);
assign n6139 = n12485 | n9192;
assign n8594 = n4515 | n10681;
assign n1229 = n599 & n876;
assign n8019 = ~n8410;
assign n11928 = ~n6826;
assign n2766 = n1438 | n1985;
assign n6868 = ~(n3260 ^ n1913);
assign n8169 = ~(n3448 | n8317);
assign n2393 = n2458 & n3409;
assign n3007 = n9450 | n12623;
assign n5048 = ~n3085;
assign n9266 = n6254 | n8326;
assign n4453 = ~n951;
assign n10011 = n4088 & n7043;
assign n10056 = n8108 | n10179;
assign n6860 = ~(n4528 | n12906);
assign n3010 = ~(n3366 ^ n570);
assign n11130 = ~n180;
assign n1338 = ~(n8368 | n9441);
assign n2371 = ~(n7879 ^ n6997);
assign n3974 = ~(n4113 ^ n1707);
assign n10043 = ~n3085;
assign n6331 = n1936 & n4383;
assign n8636 = n4148 | n900;
assign n3218 = ~(n8042 | n2533);
assign n6755 = ~n8768;
assign n1336 = ~(n11262 ^ n5379);
assign n954 = n11355 & n7774;
assign n8211 = n8843 | n4640;
assign n3813 = ~n5073;
assign n5895 = ~(n11448 ^ n9226);
assign n644 = ~n3669;
assign n10737 = ~(n10735 ^ n5276);
assign n11979 = ~(n129 ^ n2929);
assign n4557 = n428 & n5117;
assign n9241 = ~(n798 ^ n7603);
assign n1227 = n3965 | n5460;
assign n12060 = n11203 | n3926;
assign n3483 = n1712 | n12784;
assign n279 = ~(n1801 | n2477);
assign n10673 = ~n6956;
assign n6206 = ~(n8926 ^ n9469);
assign n9026 = n4980 | n2875;
assign n6117 = ~(n91 | n7641);
assign n8847 = n53 | n10761;
assign n9255 = n2973 | n5646;
assign n27 = ~(n9633 ^ n12887);
assign n11775 = n6140 & n3031;
assign n3768 = n5922 | n7874;
assign n9249 = n11591 | n10319;
assign n741 = n3077 & n2687;
assign n9369 = n12262 & n3227;
assign n7999 = n5401 | n13039;
assign n3665 = n9392 | n8464;
assign n5046 = ~(n12899 ^ n6899);
assign n5929 = ~(n10865 ^ n3010);
assign n11044 = ~(n7929 ^ n7735);
assign n1542 = n6606 | n8504;
assign n12327 = n12798 | n12240;
assign n8181 = ~(n9059 ^ n4089);
assign n5402 = ~n7841;
assign n1298 = ~(n9307 ^ n9097);
assign n7463 = n7296 & n8914;
assign n8970 = ~(n2205 ^ n2654);
assign n985 = ~(n6362 ^ n7772);
assign n393 = ~(n576 ^ n3757);
assign n7286 = ~n6347;
assign n12809 = n5806 | n121;
assign n8944 = ~(n7786 | n9562);
assign n1592 = n7086 & n666;
assign n11884 = ~(n9047 | n12231);
assign n11342 = n11842 & n10197;
assign n722 = ~(n10007 ^ n9337);
assign n357 = n9927 | n10493;
assign n9798 = ~(n4930 ^ n3070);
assign n6461 = ~(n9610 ^ n6456);
assign n9210 = ~(n13150 ^ n2396);
assign n2113 = ~(n5699 ^ n3604);
assign n209 = ~n7888;
assign n7931 = n10043 | n2675;
assign n616 = ~(n4263 | n1649);
assign n4758 = n4382 & n12284;
assign n7029 = n11311 | n5712;
assign n5960 = ~(n1041 ^ n10910);
assign n3749 = n6220 | n894;
assign n7186 = ~(n600 | n12425);
assign n12746 = n860 ^ n5393;
assign n10843 = n9513 & n1400;
assign n8782 = ~(n11589 ^ n6312);
assign n6356 = ~(n9025 | n11374);
assign n3705 = ~(n7320 ^ n8267);
assign n569 = ~n2758;
assign n7199 = ~n2787;
assign n946 = ~n5427;
assign n6939 = ~n4330;
assign n10464 = ~(n5537 ^ n11629);
assign n11596 = n8801 | n4644;
assign n7728 = n875 & n4509;
assign n3797 = n10757 & n467;
assign n623 = n6326 | n12543;
assign n1940 = n2048 | n9682;
assign n5287 = n778 & n10704;
assign n7446 = n10472 & n12172;
assign n7434 = n4037 | n7495;
assign n4168 = ~(n13163 ^ n5143);
assign n4197 = ~(n12455 | n12161);
assign n12162 = n6721 | n5076;
assign n592 = ~(n3541 ^ n2587);
assign n7031 = n12362 | n3987;
assign n4268 = n10780 | n8268;
assign n3629 = ~(n2739 | n9232);
assign n5038 = n11640 ^ n3830;
assign n11553 = n338 | n2544;
assign n8402 = n9238 | n12166;
assign n12856 = ~n1369;
assign n439 = ~(n8815 ^ n7622);
assign n3532 = n2899 | n1570;
assign n11799 = ~n10033;
assign n4101 = ~(n7181 ^ n13103);
assign n5414 = ~n10770;
assign n2998 = ~(n9022 | n10038);
assign n10067 = ~(n4695 ^ n9504);
assign n10513 = n1436 | n9159;
assign n3707 = ~(n2149 ^ n2085);
assign n2620 = ~(n108 ^ n2892);
assign n6561 = ~(n4513 ^ n9267);
assign n8476 = ~(n11321 ^ n748);
assign n13184 = n1258 & n4971;
assign n8721 = n1025 ^ n8760;
assign n455 = ~(n1904 ^ n6974);
assign n6788 = ~(n631 ^ n11724);
assign n1487 = n8253 ^ n7584;
assign n10920 = n13170 | n6404;
assign n10261 = n13012 | n1985;
assign n7017 = n860 | n8371;
assign n921 = n13194 | n4947;
assign n6257 = n8894 & n5898;
assign n12770 = n1892 | n1679;
assign n44 = ~n11109;
assign n2761 = ~(n4153 ^ n7032);
assign n2359 = n808 | n4621;
assign n9541 = ~(n10571 ^ n3798);
assign n6212 = n6182 | n2059;
assign n7045 = ~n6610;
assign n2344 = ~(n7705 | n5239);
assign n11714 = n1883 | n6404;
assign n2076 = n1451 | n2059;
assign n9848 = n234 | n3843;
assign n7843 = n6768 | n4455;
assign n4258 = ~n499;
assign n1175 = ~n5845;
assign n7911 = n2238 | n9586;
assign n11948 = ~(n2301 ^ n7524);
assign n11444 = ~(n7797 ^ n7525);
assign n12081 = ~(n12230 ^ n9542);
assign n11587 = ~(n5640 ^ n9746);
assign n12317 = ~(n550 | n6594);
assign n11406 = ~(n8758 ^ n2629);
assign n9771 = ~(n2820 ^ n4646);
assign n12520 = n7591 & n4547;
assign n431 = n4782 & n12793;
assign n4665 = ~n5884;
assign n574 = ~(n1759 | n11382);
assign n3652 = ~n3203;
assign n4946 = ~(n3251 ^ n8686);
assign n12676 = n6166 | n9195;
assign n5868 = ~(n7317 ^ n3261);
assign n9319 = n3914 & n8017;
assign n1335 = ~n5969;
assign n9597 = n11087 | n542;
assign n2668 = n66 & n4111;
assign n4119 = ~(n4814 ^ n2891);
assign n12135 = n4741 | n177;
assign n3140 = ~(n12399 ^ n10706);
assign n3867 = ~n11647;
assign n5886 = ~(n296 ^ n1083);
assign n1481 = ~(n11909 ^ n4125);
assign n3944 = n1897 | n1832;
assign n6015 = ~n11482;
assign n10292 = ~n3358;
assign n7905 = ~(n12486 ^ n892);
assign n6297 = ~(n3000 ^ n5751);
assign n13095 = ~(n6517 ^ n6493);
assign n8981 = n448 & n10345;
assign n2636 = ~n4460;
assign n9491 = ~(n3271 | n10677);
assign n4124 = ~(n9437 | n779);
assign n3165 = ~n2569;
assign n3315 = n6224 | n7186;
assign n4087 = ~n3251;
assign n3795 = n11505 | n2367;
assign n12386 = ~(n5687 ^ n3300);
assign n1632 = ~n8222;
assign n9548 = ~(n5220 | n11636);
assign n12899 = ~n6783;
assign n12255 = n2592 & n8860;
assign n4863 = n1737 | n8534;
assign n9893 = ~n42;
assign n65 = n4598 & n5843;
assign n7806 = ~(n2834 ^ n5298);
assign n8065 = ~n7309;
assign n10998 = ~n9087;
assign n11147 = ~(n4315 ^ n12278);
assign n6253 = n558 & n9294;
assign n668 = n6419 | n8030;
assign n3628 = ~(n6771 ^ n7268);
assign n6746 = n6919 & n1559;
assign n1805 = n5401 | n617;
assign n2052 = ~(n13128 ^ n12609);
assign n12371 = ~n6312;
assign n6800 = n5323 & n4094;
assign n1019 = n8058 & n2285;
assign n7622 = n1571 | n2675;
assign n2461 = ~(n4332 | n11200);
assign n8025 = n2475 & n6513;
assign n4717 = n2352 | n7049;
assign n4362 = n9711 | n9195;
assign n8301 = ~n5729;
assign n7442 = n4428 & n786;
assign n476 = n12653 | n3884;
assign n2980 = n8306 | n8563;
assign n11793 = n11920 | n8348;
assign n4855 = ~n443;
assign n4029 = n10991 | n7723;
assign n11544 = ~n12115;
assign n6661 = ~(n2986 ^ n7744);
assign n12612 = n8940 & n7720;
assign n7327 = n13031 & n9399;
assign n8088 = n11150 | n2034;
assign n2256 = ~(n3430 ^ n7557);
assign n5810 = ~(n1213 ^ n8886);
assign n8667 = ~(n11958 ^ n3469);
assign n10025 = n5243 & n10234;
assign n6804 = ~(n8930 | n8103);
assign n4576 = n6333 & n2295;
assign n1897 = ~n3964;
assign n9980 = n5448 | n5487;
assign n3410 = ~(n4050 ^ n5305);
assign n1185 = n12671 | n5242;
assign n914 = n11854 & n8644;
assign n12154 = ~(n7646 ^ n1464);
assign n4175 = n2771 & n2758;
assign n11370 = ~n3591;
assign n6088 = n3157 | n10471;
assign n7272 = ~n9336;
assign n2764 = n4792 | n10573;
assign n48 = ~n12284;
assign n8840 = ~n10622;
assign n4833 = ~(n11838 ^ n9296);
assign n3951 = n3062 | n6769;
assign n4582 = n9129 | n3459;
assign n5336 = n4363 & n12888;
assign n11391 = n12964 | n2679;
assign n2533 = n10465 | n4949;
assign n8781 = ~(n10743 | n3399);
assign n577 = ~(n1787 ^ n10399);
assign n5081 = ~(n5993 ^ n1298);
assign n4445 = n11612 | n12328;
assign n9511 = ~n287;
assign n8214 = ~(n11382 ^ n1759);
assign n2612 = ~(n11909 | n10595);
assign n12920 = n2729 | n76;
assign n811 = ~(n3540 ^ n7909);
assign n11753 = n5966 & n8257;
assign n11982 = ~n3130;
assign n6482 = ~n170;
assign n8273 = ~(n13139 ^ n4318);
assign n5435 = n9891 | n6973;
assign n4698 = ~n948;
assign n6151 = n1674 & n5274;
assign n6663 = n8211 & n6111;
assign n10505 = ~(n302 ^ n2300);
assign n9142 = ~(n12457 ^ n3449);
assign n2975 = ~n446;
assign n2493 = ~n12219;
assign n9441 = n1887 | n6635;
assign n4275 = n3537 | n8490;
assign n11100 = n3344 | n6635;
assign n5950 = ~(n5738 | n11403);
assign n8580 = ~n10276;
assign n5823 = n12581 | n5836;
assign n3384 = ~n2798;
assign n1223 = n6758 & n5930;
assign n8748 = ~(n502 | n3319);
assign n7202 = n13051 | n8383;
assign n9337 = ~(n9388 | n7520);
assign n5636 = n7798 | n2133;
assign n12971 = n6841 | n11609;
assign n311 = n4927 | n11100;
assign n5400 = ~n10504;
assign n11468 = ~n1742;
assign n5905 = ~n5083;
assign n7981 = ~(n2081 | n12810);
assign n12019 = ~n9585;
assign n5795 = n5713 | n1463;
assign n6122 = ~(n5300 ^ n3125);
assign n7079 = ~(n6605 ^ n6020);
assign n1792 = n1677 & n9814;
assign n9239 = n11061 & n287;
assign n5915 = ~n9833;
assign n7050 = ~(n10420 ^ n7466);
assign n2600 = ~n1254;
assign n1857 = ~n1110;
assign n6280 = n12213 & n6045;
assign n7814 = ~n7537;
assign n7210 = n10400 | n4724;
assign n7109 = n11262 | n2992;
assign n3801 = ~(n5805 | n9786);
assign n3841 = ~(n7153 ^ n13166);
assign n9501 = ~(n8369 | n3286);
assign n5429 = ~(n7085 ^ n1266);
assign n11233 = ~(n13236 ^ n4734);
assign n5053 = ~(n7938 | n11204);
assign n11035 = n12052 | n4253;
assign n2216 = ~(n7183 ^ n6604);
assign n4847 = n1498 ^ n9623;
assign n2972 = n1135 | n5264;
assign n9490 = ~n6892;
assign n11025 = ~(n3273 ^ n1780);
assign n2507 = n6603 | n362;
assign n6508 = n8646 | n6732;
assign n3426 = ~(n7210 ^ n12499);
assign n12768 = ~n3085;
assign n1457 = n4022 | n4936;
assign n11 = n4041 | n12404;
assign n12724 = n6684 & n2971;
assign n3916 = n7522 | n3703;
assign n407 = ~n7294;
assign n1001 = n5503 | n1452;
assign n10966 = ~n6085;
assign n11904 = ~(n7271 ^ n8618);
assign n8086 = ~(n3765 | n10734);
assign n4956 = ~(n3278 | n12385);
assign n12303 = ~n1195;
assign n8871 = n8995 | n7863;
assign n4596 = ~(n9058 ^ n4687);
assign n6920 = n10770 & n8233;
assign n902 = ~n8230;
assign n1945 = ~n10671;
assign n6537 = n7076 | n9223;
assign n12553 = ~(n12168 ^ n904);
assign n4519 = n12481 & n8750;
assign n5607 = ~n3357;
assign n5900 = n11629 | n7768;
assign n4995 = n1451 | n121;
assign n8832 = n10714 | n10474;
assign n8325 = ~n4122;
assign n9404 = ~(n13240 ^ n7285);
assign n12071 = n2646 | n9381;
assign n12557 = n542 | n8702;
assign n1374 = ~(n3931 ^ n1790);
assign n6651 = n69 | n8534;
assign n9788 = ~n12692;
assign n11421 = n4403 & n1828;
assign n7499 = ~(n11478 ^ n12208);
assign n12800 = n4334 & n1777;
assign n9786 = ~n5868;
assign n3023 = n10845 & n200;
assign n10296 = ~(n6615 | n450);
assign n10547 = n6120 & n4783;
assign n376 = n12099 & n11866;
assign n7910 = ~(n8161 ^ n38);
assign n3637 = n2109 | n2726;
assign n3500 = n11849 & n3778;
assign n12777 = n9400 | n11107;
assign n7507 = ~(n6445 | n3845);
assign n5692 = ~n6068;
assign n8255 = n5535 | n9847;
assign n4917 = ~(n9487 ^ n4870);
assign n9793 = ~n11734;
assign n255 = n7473 | n196;
assign n10386 = n2710 | n1871;
assign n3734 = ~(n5961 ^ n8190);
assign n5739 = n7484 & n3848;
assign n1619 = ~(n3193 ^ n5803);
assign n6194 = ~n9343;
assign n3380 = ~n2597;
assign n1243 = ~(n3150 | n6839);
assign n1276 = ~(n7592 ^ n11299);
assign n12399 = ~(n2103 | n12325);
assign n174 = n9588 | n10708;
assign n4113 = n9736 & n10667;
assign n11483 = ~(n11233 | n12498);
assign n5633 = n11235 | n6113;
assign n894 = ~n12853;
assign n3541 = ~(n1839 ^ n11409);
assign n2884 = ~n497;
assign n3030 = n2484 | n8383;
assign n9831 = n9283 & n7220;
assign n4522 = ~n11434;
assign n12418 = n4028 & n6851;
assign n1517 = ~(n13185 | n10309);
assign n9526 = ~(n6898 | n6027);
assign n3846 = n7827 & n10549;
assign n2816 = ~n10642;
assign n4301 = ~n6639;
assign n12936 = ~(n10593 ^ n5576);
assign n12828 = n1982 & n11488;
assign n11428 = ~(n4995 ^ n7551);
assign n12860 = ~(n4711 | n10787);
assign n6470 = ~(n7745 ^ n3844);
assign n705 = n564 & n9596;
assign n900 = ~(n8947 | n12176);
assign n13123 = n12432 | n3417;
assign n8632 = ~n6668;
assign n4575 = n9426 | n3053;
assign n6653 = n798 & n8331;
assign n12240 = ~n3472;
assign n216 = n1472 ^ n2652;
assign n8809 = ~n10126;
assign n5902 = ~(n6401 ^ n9798);
assign n6376 = n6131 | n9757;
assign n4317 = n13154 | n12273;
assign n10110 = n2183 | n6635;
assign n2815 = ~(n6248 | n8968);
assign n10293 = ~n6536;
assign n10975 = ~n9616;
assign n5570 = ~(n3002 ^ n8698);
assign n712 = ~n865;
assign n9582 = n8502 & n5720;
assign n2434 = n1447 | n206;
assign n10165 = n6847 & n8994;
assign n6992 = n8169 | n10407;
assign n12209 = ~(n10110 ^ n11195);
assign n2384 = ~(n5013 ^ n12238);
assign n8662 = n8280 | n11016;
assign n2046 = n10421 | n7935;
assign n11967 = n10469 | n4404;
assign n1754 = n9424 & n6619;
assign n11677 = ~n6765;
assign n6791 = n8236 & n3184;
assign n13147 = n6668 & n5729;
assign n11892 = ~(n8316 ^ n12353);
assign n100 = n444 | n3383;
assign n6056 = ~n10142;
assign n12635 = n8436 | n1155;
assign n6038 = n4513 & n3309;
assign n12540 = ~(n6354 ^ n8707);
assign n5742 = ~n4348;
assign n10124 = ~(n4048 ^ n827);
assign n11670 = n3304 & n4916;
assign n3590 = ~(n11925 | n11342);
assign n161 = ~n7974;
assign n4510 = ~(n2036 ^ n5925);
assign n6918 = n8294 | n10685;
assign n2523 = n5105 | n11772;
assign n1908 = ~n11454;
assign n12854 = n4975 & n10520;
assign n10854 = ~(n10933 | n10799);
assign n3451 = ~(n10405 ^ n7393);
assign n2738 = ~n3815;
assign n10795 = ~n10002;
assign n12737 = n11810 | n8268;
assign n6849 = ~(n10356 | n8809);
assign n1688 = ~n8522;
assign n2521 = ~(n2826 | n10965);
assign n1242 = n7907 & n10108;
assign n9993 = n1364 & n124;
assign n3943 = ~(n10273 | n5198);
assign n8547 = n6399 | n5063;
assign n12032 = ~n817;
assign n6278 = n3926 & n11203;
assign n1814 = n8707 & n6354;
assign n8460 = n11457 | n5349;
assign n9766 = ~(n9881 ^ n1740);
assign n9262 = ~(n12181 ^ n12130);
assign n11838 = ~n4312;
assign n4245 = n2763 & n9366;
assign n8953 = ~(n2465 ^ n11615);
assign n8796 = ~(n4685 | n1045);
assign n13073 = ~n7982;
assign n12196 = n4731 | n210;
assign n1425 = ~(n10857 ^ n4577);
assign n5553 = ~(n9895 ^ n384);
assign n8421 = n8450 | n5669;
assign n8329 = ~n6843;
assign n2772 = ~n6822;
assign n11089 = ~(n7901 ^ n8955);
assign n7048 = ~(n1766 | n1358);
assign n9639 = n13201 & n5548;
assign n9294 = ~(n6636 ^ n1660);
assign n8842 = ~(n7842 ^ n6147);
assign n11847 = n6229 | n1417;
assign n6267 = ~n1203;
assign n3300 = n4612 | n3949;
assign n12597 = n8356 | n8918;
assign n8136 = ~(n6535 ^ n4064);
assign n8226 = n240 & n8734;
assign n9057 = ~(n6478 | n11678);
assign n8823 = ~(n4571 ^ n3823);
assign n5910 = ~(n3561 | n12830);
assign n652 = ~n9093;
assign n9375 = ~n3876;
assign n8297 = ~n10728;
assign n3272 = ~(n11570 | n4239);
assign n348 = ~(n8539 ^ n2293);
assign n64 = ~n6087;
assign n9303 = n10113 & n10451;
assign n2122 = ~n8399;
assign n9010 = ~n469;
assign n4858 = ~(n9959 ^ n8896);
assign n688 = ~(n10327 | n6711);
assign n10215 = n9748 & n12895;
assign n1182 = ~(n7934 ^ n289);
assign n110 = n9273 | n9686;
assign n10072 = ~(n11930 | n3924);
assign n4770 = n10872 & n12308;
assign n7208 = n828 ^ n5483;
assign n1190 = n1952 & n2601;
assign n9273 = n2496 & n4988;
assign n5802 = ~n1874;
assign n12370 = ~n6897;
assign n4525 = n9917 | n10049;
assign n1562 = n7794 | n7563;
assign n10532 = n626 & n7887;
assign n6306 = ~n2590;
assign n9182 = ~n11280;
assign n1823 = n10984 & n3404;
assign n118 = ~n13192;
assign n12029 = n1259 & n297;
assign n6058 = n2604 & n12358;
assign n5180 = n7146 | n5076;
assign n2454 = ~(n1517 ^ n430);
assign n3237 = ~(n10643 | n3633);
assign n2794 = n9788 & n9989;
assign n12410 = ~(n3321 ^ n10190);
assign n8058 = ~n5304;
assign n851 = n5491 & n10171;
assign n6579 = ~n6226;
assign n7339 = n4608 & n1918;
assign n12170 = ~n7813;
assign n5004 = n1436 | n4640;
assign n11900 = n12033 | n4416;
assign n1833 = n13112 & n12851;
assign n9840 = ~(n12528 ^ n2694);
assign n11760 = n2003 & n9237;
assign n12880 = ~(n1896 | n11005);
assign n6754 = ~(n8272 ^ n11062);
assign n701 = n3682 | n7013;
assign n7402 = ~(n10444 | n8586);
assign n4171 = n7969 ^ n6433;
assign n12463 = ~(n1192 ^ n13029);
assign n3283 = ~(n9067 ^ n7341);
assign n11560 = n7247 | n2228;
assign n11740 = ~n8358;
assign n11431 = ~n12428;
assign n10893 = ~n2758;
assign n7502 = n11322 & n11662;
assign n6486 = ~n1231;
assign n4225 = n6051 | n11998;
assign n8980 = n7052 & n2219;
assign n4957 = n2540 ^ n9013;
assign n4999 = ~(n3909 ^ n698);
assign n12995 = ~n441;
assign n1729 = n12551 | n5781;
assign n4334 = n12997 | n2133;
assign n8641 = ~(n9734 | n8523);
assign n4446 = n3416 | n4474;
assign n2399 = ~(n668 | n6663);
assign n3539 = n5656 | n11538;
assign n3671 = ~n5684;
assign n11869 = ~n6515;
assign n699 = ~(n11859 ^ n6877);
assign n7421 = ~n4572;
assign n7071 = ~(n374 | n5225);
assign n12454 = ~(n5509 | n12875);
assign n1008 = ~n8932;
assign n10648 = ~(n2973 ^ n5646);
assign n12656 = n559 | n4947;
assign n11197 = n12602 | n3902;
assign n7111 = ~(n2212 ^ n9768);
assign n13182 = ~n9669;
assign n10052 = n9172 & n4231;
assign n3294 = n6744 & n347;
assign n8398 = ~(n5530 ^ n2138);
assign n1568 = ~(n5636 ^ n152);
assign n1489 = ~(n1657 ^ n2828);
assign n9336 = ~(n1465 ^ n12973);
assign n2237 = ~(n12897 ^ n10216);
assign n11565 = n10908 & n854;
assign n12320 = n5964 & n2270;
assign n4191 = n2937 & n10812;
assign n11632 = n10809 & n4342;
assign n5701 = ~(n2474 ^ n12017);
assign n7465 = ~(n3024 ^ n2119);
assign n368 = ~(n12410 ^ n1027);
assign n259 = n2806 & n2189;
assign n2479 = n4792 | n3454;
assign n3875 = ~(n12269 ^ n1519);
assign n12554 = ~(n10450 ^ n5201);
assign n2550 = ~n471;
assign n5281 = ~(n10806 ^ n5977);
assign n11448 = ~(n282 ^ n8916);
assign n4125 = ~(n3869 ^ n8717);
assign n7537 = n4370 | n6635;
assign n346 = n1647 & n4402;
assign n12705 = n3024 | n2119;
assign n12070 = n9968 | n9850;
assign n10912 = n628 | n10106;
assign n4010 = n11664 | n9795;
assign n4235 = n12093 | n12847;
assign n5623 = n7538 & n2782;
assign n6811 = ~n4387;
assign n8734 = n4251 | n3079;
assign n10183 = n8053 | n2675;
assign n10051 = ~n3298;
assign n8338 = ~(n1375 | n12097);
assign n1372 = n6904 | n5915;
assign n3555 = ~n9188;
assign n4492 = n11318 & n8880;
assign n12900 = n5252 & n2573;
assign n7599 = ~(n11193 ^ n6705);
assign n8415 = ~(n9790 | n10831);
assign n7722 = n6333 & n834;
assign n9622 = ~n6392;
assign n728 = ~(n3271 ^ n1776);
assign n5129 = n8969 | n9141;
assign n228 = ~(n5725 ^ n5928);
assign n10763 = ~(n149 ^ n6773);
assign n6784 = ~(n4359 ^ n12775);
assign n4104 = n1567 | n12400;
assign n1048 = n9675 | n6265;
assign n12199 = ~(n8891 ^ n3182);
assign n1158 = n3225 | n6265;
assign n9537 = ~n11324;
assign n2388 = n4732 | n4230;
assign n12173 = ~(n4000 ^ n8477);
assign n7542 = n11087 | n2449;
assign n7184 = ~n12579;
assign n5589 = n7085 | n1781;
assign n587 = ~(n6572 ^ n6546);
assign n11452 = ~n5174;
assign n9366 = n11335 | n2123;
assign n13087 = n13243 & n7003;
assign n9572 = n12877 & n12288;
assign n7548 = ~(n10477 | n8965);
assign n2449 = n10240;
assign n5386 = ~(n6887 ^ n13024);
assign n4108 = n13117 | n10871;
assign n9905 = n420 & n1798;
assign n575 = n8067 & n10817;
assign n11909 = n334 | n12948;
assign n8972 = n10761 | n1570;
assign n9203 = n4099 & n10691;
assign n5526 = n2195 | n3523;
assign n11135 = ~(n6195 | n1900);
assign n9610 = ~(n2992 ^ n1336);
assign n6377 = n8688 & n548;
assign n8453 = ~n7165;
assign n13138 = n10756 | n9195;
assign n10001 = ~(n3822 ^ n1613);
assign n2092 = n7339 & n5695;
assign n11644 = ~(n11881 | n9535);
assign n7968 = n9705 ^ n12101;
assign n10341 = n1113 | n1144;
assign n5609 = ~(n5914 ^ n12729);
assign n10239 = ~(n279 | n11338);
assign n4694 = ~n1543;
assign n3653 = n6188 & n12922;
assign n1996 = n5711 & n5085;
assign n301 = ~(n1617 ^ n5596);
assign n5404 = ~(n528 ^ n5870);
assign n10356 = ~(n1553 ^ n7964);
assign n4589 = ~n6601;
assign n1095 = ~(n4197 | n4697);
assign n3443 = n11608 & n7657;
assign n1637 = ~(n2242 ^ n9073);
assign n9733 = n1983 | n6255;
assign n9228 = ~n10162;
assign n10757 = ~n2703;
assign n8410 = n9622 | n4420;
assign n2288 = ~(n6902 ^ n10750);
assign n2534 = n7981 | n6089;
assign n8801 = n2919 | n12388;
assign n9590 = n6423 & n593;
assign n12689 = n6206 | n11097;
assign n6313 = ~n11993;
assign n7917 = n5949 | n6635;
assign n10198 = ~n9943;
assign n929 = n4334 | n1777;
assign n2355 = n8994 | n6847;
assign n5155 = n4418 | n6926;
assign n12841 = ~n9475;
assign n3019 = n2162 & n4678;
assign n7936 = ~(n12085 ^ n2071);
assign n6428 = n4809 | n3632;
assign n8967 = ~(n3625 ^ n6871);
assign n6527 = ~(n11743 | n12727);
assign n12622 = n2266 & n3743;
assign n2993 = n11120 | n5885;
assign n7708 = ~n7585;
assign n8345 = ~(n1735 ^ n10164);
assign n12548 = n12141 | n10513;
assign n4394 = ~(n5445 ^ n5681);
assign n4380 = ~(n10186 ^ n8151);
assign n3468 = ~n10150;
assign n8803 = n7128 ^ n4078;
assign n9027 = ~(n3833 ^ n3754);
assign n298 = n3821 | n12755;
assign n4223 = n5510 & n5795;
assign n4271 = ~(n5762 ^ n2501);
assign n9209 = ~n9843;
assign n5315 = n8668 & n8381;
assign n6536 = ~(n9831 ^ n11025);
assign n9900 = n2613 | n12233;
assign n10031 = ~(n4713 | n11441);
assign n10431 = ~(n2167 | n7535);
assign n949 = n7675 | n9195;
assign n10045 = ~n3076;
assign n2683 = ~(n1400 ^ n9513);
assign n7976 = ~(n11131 | n1137);
assign n6162 = n5867 & n8088;
assign n2907 = n8816 & n11999;
assign n3587 = ~n1084;
assign n3138 = ~(n1009 ^ n3678);
assign n5190 = n2903 & n8803;
assign n4703 = n11324 & n1724;
assign n11865 = ~(n8551 ^ n1249);
assign n7338 = ~(n11095 | n6390);
assign n2895 = ~(n1975 ^ n356);
assign n5989 = n644 | n542;
assign n12820 = n8600 ^ n3137;
assign n1643 = ~(n2817 | n1299);
assign n3004 = n4313 | n3487;
assign n4012 = ~(n1223 | n7673);
assign n63 = ~n9531;
assign n13093 = n7276 & n3106;
assign n4866 = ~n2038;
assign n5791 = n5371 & n3097;
assign n3503 = ~(n1607 ^ n2745);
assign n5863 = n3408 | n11086;
assign n12718 = ~n11537;
assign n1210 = n1072 | n2851;
assign n4940 = n11269 | n8196;
assign n4205 = n4612 | n8563;
assign n10572 = ~(n12419 ^ n3196);
assign n5416 = n4668 | n12726;
assign n2968 = ~(n374 ^ n11992);
assign n4185 = ~n9887;
assign n10712 = n1571 | n6265;
assign n3673 = ~(n1752 | n11106);
assign n7001 = ~n8273;
assign n11185 = ~n1278;
assign n4296 = ~(n6118 ^ n1229);
assign n9230 = ~(n10412 ^ n4031);
assign n8990 = ~(n3874 | n7198);
assign n3729 = ~n7238;
assign n8501 = ~(n8289 ^ n1502);
assign n1418 = n9942 & n890;
assign n7621 = ~(n8632 | n9913);
assign n7774 = ~(n5642 ^ n4422);
assign n6372 = n10761 | n6404;
assign n8685 = n4878 & n10141;
assign n1704 = n519 & n11896;
assign n9856 = ~(n5093 ^ n2506);
assign n11922 = ~n1923;
assign n3710 = ~(n4192 ^ n7114);
assign n6373 = ~(n7101 ^ n1132);
assign n11415 = n470 & n8370;
assign n8174 = ~n11835;
assign n8604 = ~(n99 ^ n10416);
assign n309 = n11876 & n1657;
assign n9781 = n3478 | n5537;
assign n9829 = ~n3894;
assign n12175 = n8757 | n6404;
assign n4673 = n1184 & n11188;
assign n4252 = n959 ^ n4758;
assign n8448 = n10448 | n5076;
assign n8625 = n4208 | n1144;
assign n10396 = ~(n6651 ^ n9657);
assign n9128 = ~(n7581 ^ n9973);
assign n896 = n9225 | n3023;
assign n7095 = n5019 | n6141;
assign n4966 = ~(n1549 | n5753);
assign n472 = ~(n12133 ^ n7595);
assign n3848 = n4272 | n5797;
assign n3806 = ~(n1178 ^ n10489);
assign n3592 = n3096 | n542;
assign n6667 = n1968 | n12745;
assign n2732 = n1160 & n2446;
assign n7894 = n9911 | n1843;
assign n1954 = ~n10398;
assign n12148 = ~(n12172 ^ n5223);
assign n11582 = n12904 & n12427;
assign n1139 = n9901 & n11801;
assign n10129 = n7934 | n289;
assign n11227 = ~n6868;
assign n6161 = ~(n7978 ^ n1129);
assign n3376 = n8873 & n4804;
assign n10085 = ~n5969;
assign n4110 = n2223 & n4706;
assign n10425 = ~n727;
assign n4707 = n9776 ^ n4037;
assign n10637 = n2463 | n10871;
assign n5016 = ~n10563;
assign n5328 = ~n9747;
assign n9168 = n5671 & n3769;
assign n1265 = n13170 | n12388;
assign n7242 = ~n6195;
assign n1660 = ~(n11272 ^ n10087);
assign n10479 = n12673 & n7761;
assign n8083 = n3647 & n5098;
assign n8147 = ~(n12389 ^ n6138);
assign n7426 = ~(n12817 ^ n12872);
assign n155 = n652 | n2544;
assign n5887 = ~(n6425 | n13091);
assign n12502 = ~(n11392 ^ n9760);
assign n2229 = n7715 & n12306;
assign n10927 = ~n5334;
assign n10548 = ~(n9270 ^ n2422);
assign n6204 = n8040 & n7464;
assign n12805 = n10641 | n11152;
assign n8587 = n5601 & n10265;
assign n4401 = n6304 | n539;
assign n10819 = n7609 & n11924;
assign n2648 = n9464 & n9191;
assign n6158 = ~(n3526 ^ n350);
assign n6833 = n5517 & n12559;
assign n303 = n2091 | n3597;
assign n9079 = ~(n7406 ^ n1182);
assign n13240 = n698 & n3909;
assign n6289 = ~(n6893 | n948);
assign n13230 = ~(n10496 ^ n5159);
assign n2425 = n9089 | n7760;
assign n9305 = ~n5189;
assign n11592 = ~(n3105 ^ n6410);
assign n3093 = ~(n7438 ^ n3732);
assign n10887 = ~(n7448 ^ n194);
assign n1024 = n2057 & n834;
assign n8542 = n8228 & n411;
assign n8951 = ~n486;
assign n2532 = ~(n293 | n7150);
assign n11806 = ~n9376;
assign n11243 = ~(n9365 ^ n636);
assign n9666 = n7208 ^ n11846;
assign n4288 = n3000 | n9971;
assign n12875 = n4725 & n2265;
assign n10607 = n8922 | n5389;
assign n2054 = ~(n8990 ^ n3675);
assign n11509 = ~n4441;
assign n798 = ~(n217 ^ n3889);
assign n4091 = n953 & n8107;
assign n10007 = ~(n1564 | n512);
assign n8729 = ~n7411;
assign n6808 = ~n323;
assign n12757 = ~(n9958 | n3719);
assign n9022 = ~(n12974 | n11587);
assign n2004 = ~(n3484 | n13189);
assign n8611 = ~(n11383 ^ n8396);
assign n4316 = n5461 | n2449;
assign n648 = ~(n10568 ^ n12520);
assign n9438 = n11370 | n5797;
assign n4521 = n7626 | n5340;
assign n7522 = ~n2737;
assign n13001 = n5218 | n496;
assign n12721 = ~n3130;
assign n12455 = n18 | n11668;
assign n790 = n7537 ^ n3211;
assign n9394 = ~(n9364 ^ n10058);
assign n5699 = ~(n11312 ^ n7812);
assign n11501 = n11037 | n2059;
assign n5350 = n12150 | n4145;
assign n13004 = ~(n5720 ^ n8502);
assign n4806 = ~(n9894 ^ n5210);
assign n3161 = ~(n4834 ^ n11934);
assign n2309 = ~(n8362 ^ n4011);
assign n4019 = ~(n4941 ^ n2628);
assign n9044 = n6003 | n10579;
assign n9651 = ~n10709;
assign n5373 = n3557 & n6742;
assign n11923 = ~(n5778 ^ n2381);
assign n11508 = n4398 & n8997;
assign n8894 = ~(n6273 ^ n12144);
assign n1576 = ~(n10620 ^ n1569);
assign n4144 = ~n4470;
assign n3775 = n9888 & n6394;
assign n9103 = ~(n7012 ^ n1160);
assign n12059 = ~(n7324 ^ n7996);
assign n10755 = ~n6196;
assign n12701 = n2268 & n3245;
assign n8992 = n1871 & n2710;
assign n10729 = ~(n8922 ^ n11759);
assign n6919 = n5212 & n6802;
assign n4991 = ~(n10766 ^ n2078);
assign n13025 = ~n443;
assign n227 = ~n8290;
assign n9330 = n1340 | n8435;
assign n3220 = ~(n10344 | n266);
assign n10433 = ~n9620;
assign n2208 = ~(n3218 | n6437);
assign n6394 = n8940 & n6392;
assign n9358 = ~(n5479 ^ n2951);
assign n5094 = n6680 | n7306;
assign n10335 = n7184 | n8268;
assign n8191 = ~(n6499 ^ n7343);
assign n4299 = ~(n5941 ^ n4972);
assign n2143 = ~(n5585 ^ n8092);
assign n4902 = ~(n1454 ^ n9185);
assign n3636 = n569 | n9195;
assign n12699 = n10830 | n6732;
assign n10764 = ~n10408;
assign n10644 = ~n12550;
assign n4214 = ~(n6898 ^ n10146);
assign n5149 = n9980 & n11424;
assign n8319 = n9217 & n3688;
assign n2621 = n7240 & n1528;
assign n2112 = n190 & n12063;
assign n9297 = n10781 | n8268;
assign n5573 = ~(n4550 | n3968);
assign n13127 = n9476 | n3772;
assign n5608 = n2802 | n12410;
assign n558 = ~n212;
assign n11654 = n584 | n10029;
assign n9947 = ~(n1393 ^ n5442);
assign n3230 = n12976 & n4533;
assign n1586 = n8480 | n10012;
assign n4803 = ~(n5358 ^ n7027);
assign n10377 = ~(n10115 | n9799);
assign n12248 = ~(n8842 ^ n5984);
assign n7571 = n4657 | n10179;
assign n760 = n9878 & n3030;
assign n5443 = ~(n7454 | n7099);
assign n2261 = n13012 | n11107;
assign n5507 = ~(n12593 | n350);
assign n10211 = ~n12356;
assign n911 = ~(n8135 | n6822);
assign n6258 = ~(n7460 | n4450);
assign n2060 = ~(n1864 ^ n10712);
assign n4840 = n12378 & n11059;
assign n12125 = ~(n8284 ^ n4543);
assign n11932 = ~(n9206 ^ n2645);
assign n8379 = ~(n9948 ^ n6288);
assign n816 = ~n8071;
assign n3939 = n9710 & n11846;
assign n2326 = n11492 | n8711;
assign n8413 = ~n7376;
assign n8674 = ~(n2442 ^ n8634);
assign n12799 = n3003 | n4662;
assign n4352 = ~n6085;
assign n5574 = ~(n2786 ^ n669);
assign n1490 = n2556 | n4230;
assign n10592 = ~(n1131 ^ n8192);
assign n324 = ~(n6396 | n11425);
assign n13044 = n9966 & n4720;
assign n10503 = n5847 | n7515;
assign n9568 = n5921 & n8571;
assign n8655 = ~n1626;
assign n5973 = ~n12284;
assign n5708 = n6580 & n8942;
assign n6519 = ~n2339;
assign n7592 = ~(n1763 ^ n5132);
assign n9516 = ~(n8979 ^ n10320);
assign n9757 = n2427 & n2178;
assign n4530 = ~n832;
assign n11311 = n2736 & n2659;
assign n2346 = ~n12579;
assign n10756 = ~n3409;
assign n614 = n1553 | n7964;
assign n9381 = n9468 & n11919;
assign n11929 = ~n9906;
assign n12122 = n7805 | n2059;
assign n11496 = ~(n7114 | n4192);
assign n8209 = n5275 & n3109;
assign n4702 = ~(n7693 | n5977);
assign n4851 = n11587 & n12974;
assign n199 = n7026 & n10964;
assign n943 = n3109 | n5275;
assign n1719 = n11498 & n458;
assign n3798 = n12788 & n6900;
assign n3603 = ~(n7958 ^ n2682);
assign n5308 = ~(n10538 | n5650);
assign n2210 = ~(n7345 | n11613);
assign n4918 = ~(n5110 ^ n1217);
assign n8730 = n794 & n2980;
assign n7647 = ~(n10666 | n10752);
assign n7408 = ~(n12728 ^ n9139);
assign n1130 = n2104 & n10808;
assign n1966 = ~(n6545 ^ n4131);
assign n4483 = ~(n3007 ^ n8847);
assign n12691 = ~(n998 ^ n1399);
assign n8288 = ~(n7938 ^ n12966);
assign n2924 = n7152 | n1570;
assign n9834 = n2204 | n1546;
assign n11477 = ~(n4181 ^ n11013);
assign n867 = n8850 | n9907;
assign n1401 = n66 ^ n4111;
assign n818 = n13173 & n1388;
assign n2018 = ~n10866;
assign n2759 = n10662 & n13027;
assign n9256 = n1474 | n5450;
assign n8038 = ~n2771;
assign n11816 = ~(n10961 ^ n6552);
assign n1527 = n6063 | n2544;
assign n2652 = n5586 & n12263;
assign n2219 = ~(n4574 ^ n12340);
assign n12752 = ~n6032;
assign n8300 = ~(n4648 ^ n11155);
assign n8862 = n321 | n3981;
assign n7871 = n11827 & n9395;
assign n7929 = n11231 & n9202;
assign n6125 = n2641 | n6404;
assign n2539 = n10099 & n10275;
assign n12402 = n9910 | n9741;
assign n10545 = n7915 & n5395;
assign n10046 = ~(n3238 | n9242);
assign n7602 = ~n8822;
assign n9253 = n4876 | n769;
assign n10135 = ~n2758;
assign n4541 = ~(n1928 ^ n8089);
assign n4344 = ~(n3585 | n5779);
assign n7196 = n5477 | n5174;
assign n6621 = ~(n8976 ^ n13179);
assign n11901 = n3892 | n7935;
assign n8857 = ~n7116;
assign n9447 = ~(n791 ^ n2376);
assign n3556 = n2848 | n479;
assign n5076 = n218;
assign n2554 = ~(n8272 | n3337);
assign n8197 = ~(n364 ^ n5178);
assign n8496 = n9519 | n6541;
assign n1199 = ~n12289;
assign n12487 = ~(n4797 | n1405);
assign n6563 = ~n5284;
assign n10676 = n11562 | n7335;
assign n9778 = n12220 & n2100;
assign n11285 = ~(n5945 ^ n13199);
assign n111 = ~n11433;
assign n3584 = ~n4630;
assign n11114 = ~n10594;
assign n8117 = ~(n7680 ^ n12818);
assign n9408 = n10427 & n3424;
assign n5931 = ~(n8631 | n9752);
assign n12894 = ~(n3819 ^ n10295);
assign n7262 = ~n4682;
assign n6975 = n7216 | n8563;
assign n4639 = n334 | n3225;
assign n2964 = ~(n4475 ^ n6999);
assign n166 = ~(n7639 ^ n4327);
assign n9229 = n5227 & n6391;
assign n10578 = n9701 & n10457;
assign n12925 = ~(n12777 ^ n13210);
assign n5270 = n1757 & n9669;
assign n94 = ~(n6549 ^ n9167);
assign n6321 = n7595 & n12133;
assign n11465 = n5308 | n9379;
assign n6521 = ~(n3322 | n4913);
assign n83 = ~(n7376 ^ n1567);
assign n589 = n11635 & n3006;
assign n6910 = ~(n6471 | n4955);
assign n9602 = ~(n5345 | n11727);
assign n2271 = ~n1646;
assign n10401 = ~(n5380 ^ n7417);
assign n7920 = ~(n197 | n8785);
assign n12560 = n4366 | n6635;
assign n6848 = ~(n9700 ^ n4652);
assign n6764 = ~n564;
assign n3497 = n1739 & n11462;
assign n3472 = ~(n11280 ^ n8000);
assign n1012 = ~n11488;
assign n4973 = ~(n2258 ^ n4017);
assign n1153 = n6970 & n4445;
assign n1973 = ~n9032;
assign n5737 = n9310 | n6040;
assign n8753 = n6004 | n12443;
assign n462 = n5261 | n5242;
assign n8545 = n9809 | n1094;
assign n1161 = n8305 & n9695;
assign n4137 = n2027 | n6728;
assign n7307 = n685 & n8068;
assign n144 = n2381 | n5778;
assign n12593 = ~(n3526 | n12933);
assign n5987 = ~(n6531 ^ n1717);
assign n3945 = n12376 | n6081;
assign n694 = ~n772;
assign n2681 = ~n5735;
assign n3513 = n11419 & n943;
assign n5332 = ~(n3209 ^ n8721);
assign n6608 = ~n1972;
assign n3406 = ~(n12431 ^ n3782);
assign n12584 = n8463 | n7306;
assign n11136 = ~(n11935 ^ n3811);
assign n8141 = n13159 | n3981;
assign n7331 = n1398 | n11616;
assign n12641 = n162 & n8051;
assign n1157 = n5459 & n5474;
assign n5952 = ~(n8521 ^ n2577);
assign n3676 = ~n937;
assign n8893 = ~(n11379 ^ n11995);
assign n5162 = n484 & n7618;
assign n13156 = ~(n10583 | n5241);
assign n6246 = ~(n1225 ^ n8583);
assign n11262 = n160 ^ n6585;
assign n5988 = n12776 | n11603;
assign n5264 = ~n411;
assign n11576 = n2624 & n5135;
assign n1283 = ~(n10658 ^ n11579);
assign n721 = n667 & n5693;
assign n4017 = n8239 & n12500;
assign n6552 = ~(n8394 ^ n5310);
assign n9785 = ~(n4717 ^ n5115);
assign n11409 = ~(n6189 ^ n5685);
assign n6113 = n10772 | n4947;
assign n12219 = n10044 & n1376;
assign n5476 = ~(n12885 | n2629);
assign n10943 = n10761 | n12328;
assign n8477 = ~(n5795 ^ n5510);
assign n12001 = n6359 | n6014;
assign n7306 = ~n5920;
assign n7483 = n8609 | n12174;
assign n6838 = n4186 & n1269;
assign n2221 = ~n6392;
assign n3613 = n1002 & n5390;
assign n11388 = ~(n6811 ^ n11364);
assign n12904 = n10279 | n9754;
assign n4292 = ~(n9584 ^ n7948);
assign n11485 = ~n5784;
assign n6420 = ~n959;
assign n12261 = ~(n10313 ^ n1782);
assign n5584 = n4269 & n8293;
assign n9397 = n995 & n12970;
assign n12730 = ~(n11669 ^ n7936);
assign n3805 = ~n9915;
assign n1896 = n12955 | n488;
assign n4184 = n3963 | n9492;
assign n1041 = ~n9508;
assign n10973 = n9277 ^ n6269;
assign n5809 = n3575 & n2700;
assign n9386 = ~(n7426 | n5080);
assign n6022 = ~(n3530 ^ n5676);
assign n4442 = ~n6668;
assign n9363 = ~(n10703 | n4905);
assign n6189 = n1971 & n939;
assign n7557 = n10426 & n2098;
assign n11727 = ~(n1294 | n12975);
assign n942 = ~(n3721 ^ n4053);
assign n12430 = n12535 & n2271;
assign n5726 = n8592 & n8579;
assign n8789 = n2744 & n12424;
assign n12885 = ~n8758;
assign n5322 = ~(n5603 ^ n1176);
assign n12787 = n5054 & n1574;
assign n1696 = ~n761;
assign n12009 = ~n7729;
assign n11053 = n6451 | n8032;
assign n7591 = n12767 | n10445;
assign n2814 = ~(n12286 ^ n113);
assign n11818 = n7317 | n3261;
assign n7358 = ~n3669;
assign n5488 = ~(n6156 ^ n12403);
assign n7132 = ~(n8822 ^ n1162);
assign n1755 = ~(n2928 ^ n3228);
assign n2108 = ~(n11228 ^ n7529);
assign n9698 = ~n11930;
assign n13208 = ~(n9164 ^ n3256);
assign n1545 = n10437 | n2544;
assign n7454 = ~(n108 | n2892);
assign n306 = n3070 & n4930;
assign n3510 = ~n3974;
assign n3005 = ~(n11718 ^ n5081);
assign n1211 = ~n10186;
assign n3098 = ~(n6813 ^ n3284);
assign n1676 = n377 & n6930;
assign n6863 = n4433 & n9964;
assign n6247 = n3512 & n5794;
assign n10244 = ~n1974;
assign n11504 = n7033 | n10213;
assign n11564 = n11192 | n9199;
assign n12245 = ~(n11657 ^ n10176);
assign n5821 = n5455 | n4373;
assign n10148 = ~(n6525 | n12730);
assign n7091 = ~n6763;
assign n4905 = ~(n8442 ^ n221);
assign n6360 = ~n11584;
assign n12109 = ~n1165;
assign n11682 = ~(n1090 ^ n7835);
assign n7877 = ~n7281;
assign n8494 = ~n7844;
assign n9050 = ~(n4898 ^ n3028);
assign n4008 = ~(n4496 ^ n3370);
assign n3329 = n7156 & n1932;
assign n3834 = n10883 | n10319;
assign n1390 = ~n4135;
assign n5644 = n1139 | n6216;
assign n3321 = n6295 | n2637;
assign n8533 = ~n3439;
assign n354 = n9579 & n5233;
assign n5119 = ~n7734;
assign n6444 = n3958 | n2846;
assign n1737 = ~n8290;
assign n1014 = ~(n3893 ^ n1993);
assign n6385 = n2673 & n5726;
assign n2298 = n3928 | n10871;
assign n12466 = ~(n12864 | n2110);
assign n1248 = ~(n8308 | n5214);
assign n13101 = n1941 | n4640;
assign n12578 = n8308 & n9669;
assign n1293 = ~(n6738 ^ n9486);
assign n2276 = ~n8183;
assign n2470 = ~(n3654 ^ n12070);
assign n7038 = ~(n2764 ^ n4123);
assign n1508 = ~n6471;
assign n2176 = ~(n8659 ^ n9755);
assign n6419 = ~n7113;
assign n682 = ~(n3695 | n5723);
assign n830 = n4153 | n10973;
assign n3240 = n12851 | n13112;
assign n5539 = ~(n114 | n10866);
assign n7259 = ~(n13000 ^ n9753);
assign n8059 = ~(n10326 ^ n7793);
assign n4082 = ~(n540 ^ n8760);
assign n2212 = n7662 & n1006;
assign n1981 = ~(n10564 | n7521);
assign n2151 = n11840 & n12036;
assign n2007 = ~(n12716 | n7785);
assign n12585 = n6801 | n4062;
assign n192 = ~n4821;
assign n5877 = n9159 | n5076;
assign n2398 = n4456 & n5353;
assign n6740 = ~(n2310 ^ n7605);
assign n6389 = n7154 & n8898;
assign n416 = ~(n6104 ^ n9053);
assign n846 = ~(n7779 ^ n2482);
assign n11591 = ~n854;
assign n6042 = ~(n3061 | n13192);
assign n1212 = n5168 | n10029;
assign n10780 = ~n3112;
assign n10947 = n6303 | n10601;
assign n11577 = ~(n12756 | n8557);
assign n5804 = ~(n8919 ^ n167);
assign n4741 = ~n11634;
assign n3413 = ~n684;
assign n2427 = n2357 | n11857;
assign n7919 = ~(n7467 ^ n1476);
assign n2731 = n9721 & n7606;
assign n1148 = n11225 | n4373;
assign n12412 = n7172 | n11978;
assign n5074 = n12256 & n10353;
assign n7065 = ~(n4458 ^ n11083);
assign n5406 = n11195 & n10110;
assign n6381 = ~n9906;
assign n4920 = n5279 & n10305;
assign n9373 = ~(n4507 ^ n1342);
assign n2075 = ~(n8420 ^ n12064);
assign n9688 = ~(n656 ^ n3685);
assign n1975 = n7707 | n121;
assign n6185 = ~(n9728 ^ n11555);
assign n8532 = ~n4335;
assign n11524 = ~(n1225 | n6716);
assign n2428 = n7889 | n2685;
assign n3547 = n3520 | n6377;
assign n424 = n10256 | n10871;
assign n11423 = n1571 | n6404;
assign n218 = ~n7715;
assign n4656 = ~(n4491 ^ n7733);
assign n5201 = ~(n9462 ^ n11795);
assign n11209 = n2236 & n5774;
assign n6108 = n4310 & n13205;
assign n5807 = n9479 | n8883;
assign n8792 = n10712 | n1864;
assign n10298 = ~(n8288 ^ n10442);
assign n9338 = ~(n8497 | n7400);
assign n1861 = ~(n9227 | n9207);
assign n3196 = ~(n790 ^ n7528);
assign n10365 = ~(n12157 ^ n6070);
assign n1732 = ~n7617;
assign n5731 = ~(n11681 ^ n13065);
assign n4061 = n3132 | n5286;
assign n4165 = n2589 & n12806;
assign n7413 = n3898 | n3981;
assign n4735 = ~(n749 | n7756);
assign n9291 = ~(n4685 ^ n12443);
assign n11201 = ~(n10070 ^ n10663);
assign n6703 = ~(n13220 | n3232);
assign n8736 = n13149 | n13113;
assign n12287 = n2281 & n973;
assign n6097 = ~n1718;
assign n988 = ~(n2169 ^ n8624);
assign n4781 = ~(n3153 ^ n3806);
assign n7256 = ~(n6523 ^ n9241);
assign n641 = n6939 | n9195;
assign n1163 = ~(n2090 ^ n11305);
assign n9212 = n677 & n5703;
assign n2094 = ~(n11655 | n870);
assign n6021 = ~(n8908 ^ n8376);
assign n1074 = ~(n1746 | n262);
assign n3466 = n4857 | n3747;
assign n6749 = ~n103;
assign n737 = ~n8163;
assign n9968 = n3746 & n10913;
assign n5401 = ~n4998;
assign n6464 = ~n9705;
assign n7564 = n2861 | n206;
assign n5146 = ~n603;
assign n3931 = ~n7455;
assign n217 = ~(n2476 ^ n10707);
assign n10710 = n5035 | n859;
assign n11446 = ~n411;
assign n6485 = ~(n3888 ^ n7828);
assign n12031 = ~n344;
assign n6380 = ~n4773;
assign n11782 = ~(n9640 ^ n12158);
assign n2456 = ~(n6366 | n6871);
assign n12529 = n1941 | n10106;
assign n7351 = n8329 | n4724;
assign n7895 = n5772 & n7899;
assign n5551 = ~(n7426 ^ n635);
assign n1902 = ~(n7401 ^ n5852);
assign n12323 = n6259 | n3461;
assign n9860 = n3630 | n2675;
assign n4227 = ~n502;
assign n12389 = ~(n10608 ^ n12898);
assign n2248 = n9679 | n11137;
assign n3378 = ~(n7354 ^ n501);
assign n861 = n6388 | n8461;
assign n2961 = n6568 | n6290;
assign n2680 = n4128 | n9982;
assign n12260 = ~(n11685 ^ n6124);
assign n222 = n3816 | n4682;
assign n1706 = ~n10167;
assign n3012 = n3901 & n12326;
assign n4543 = n2318 & n12046;
assign n104 = n9769 | n6044;
assign n12194 = ~(n11918 | n6962);
assign n10842 = n4105 & n9354;
assign n12407 = ~(n10513 ^ n1550);
assign n5946 = n4988 | n2496;
assign n9963 = ~(n7811 ^ n6179);
assign n1441 = n9040 & n4381;
assign n3197 = n5018 | n4477;
assign n11946 = n12394 | n8367;
assign n9145 = ~n1641;
assign n3888 = n7780 | n10871;
assign n9484 = n628 | n9195;
assign n461 = ~(n10132 ^ n1779);
assign n1813 = ~n6661;
assign n5723 = n12812 & n602;
assign n213 = ~(n6043 ^ n12423);
assign n2077 = ~(n11261 | n4216);
assign n11844 = ~(n7882 | n1923);
assign n10521 = n6591 & n11385;
assign n6304 = ~(n11937 | n2920);
assign n1118 = ~(n7933 ^ n7244);
assign n10161 = ~n2164;
assign n4274 = n7414 | n8845;
assign n8138 = n4201 | n2059;
assign n6064 = n2482 & n6149;
assign n9138 = ~(n2024 ^ n12006);
assign n13016 = n3783 | n10818;
assign n692 = n8062 | n99;
assign n4410 = ~(n10476 ^ n8809);
assign n8647 = n3282 & n7196;
assign n3601 = ~(n1766 ^ n976);
assign n4002 = n4506 & n3617;
assign n10476 = ~n10356;
assign n9380 = ~n12820;
assign n3069 = n1733 | n7079;
assign n8079 = ~n9620;
assign n168 = ~n6386;
assign n4089 = n11661 & n9525;
assign n6693 = ~(n8048 ^ n11210);
assign n3038 = ~n5572;
assign n5925 = ~(n2434 ^ n12854);
assign n8312 = ~(n9347 ^ n10933);
assign n2199 = ~n5336;
assign n3465 = ~(n492 ^ n5894);
assign n3778 = n4432 | n6119;
assign n6037 = ~(n13226 | n13064);
assign n8772 = ~(n9877 ^ n7777);
assign n191 = n8065 & n2157;
assign n1469 = n4982 & n3652;
assign n8855 = ~n1192;
assign n1348 = ~(n3771 ^ n158);
assign n7020 = n1504 & n11669;
assign n12141 = n7291 | n2287;
assign n3985 = n12620 & n6170;
assign n9996 = n8486 & n3141;
assign n9165 = ~(n10941 ^ n7407);
assign n11588 = ~(n7307 ^ n1818);
assign n852 = n11869 & n8755;
assign n11876 = n1377 | n6760;
assign n5050 = n10923 | n804;
assign n2281 = n6625 & n9346;
assign n9630 = ~(n7225 | n5126);
assign n559 = ~n5920;
assign n1294 = n1051 | n1144;
assign n2435 = ~(n942 ^ n2084);
assign n6762 = ~(n12124 ^ n12205);
assign n9842 = ~(n7177 ^ n12265);
assign n5672 = n6365 ^ n872;
assign n2542 = ~n6668;
assign n4443 = n11427 & n2021;
assign n4170 = ~(n7714 | n7338);
assign n12304 = ~n5951;
assign n525 = n8637 | n3686;
assign n11880 = n5694 | n10319;
assign n2791 = ~n9358;
assign n7382 = ~(n3033 ^ n11207);
assign n9364 = ~(n6202 ^ n8897);
assign n10653 = ~(n11248 ^ n5179);
assign n5063 = ~(n4242 | n598);
assign n6035 = n2338 | n10319;
assign n1476 = ~(n3780 ^ n8685);
assign n9692 = ~(n7051 ^ n9380);
assign n8546 = n13159 | n10319;
assign n1557 = n3791 | n10008;
assign n6398 = ~(n226 | n12075);
assign n9095 = ~n8330;
assign n3320 = n1959 & n11139;
assign n9861 = n8585 | n5076;
assign n5169 = ~n2771;
assign n5606 = ~(n419 | n6577);
assign n7711 = ~(n50 ^ n11782);
assign n9075 = n16;
assign n8920 = ~(n6804 ^ n8372);
assign n6460 = ~(n699 ^ n6798);
assign n7021 = ~(n1123 ^ n7967);
assign n5152 = ~n9093;
assign n13008 = ~(n7797 | n5996);
assign n12882 = ~n1307;
assign n6633 = n5017 & n1019;
assign n8425 = n434 | n3787;
assign n10449 = ~(n1840 ^ n8844);
assign n9525 = n10566 | n11877;
assign n6573 = ~(n12041 | n2635);
assign n3290 = ~(n4749 ^ n9044);
assign n6631 = ~(n3288 ^ n5291);
assign n11516 = ~(n1568 ^ n11043);
assign n2103 = ~(n5799 | n9645);
assign n2866 = ~(n299 ^ n10773);
assign n3830 = n5031 & n8233;
assign n6179 = n5634 | n3981;
assign n4598 = n8976 | n13179;
assign n13185 = n1728 & n5551;
assign n6586 = ~(n9381 ^ n10192);
assign n3325 = n7393 | n6266;
assign n4106 = ~(n5395 ^ n11639);
assign n5799 = n6332 | n6404;
assign n2701 = ~n10451;
assign n1915 = n7149 & n6098;
assign n5278 = n8095 | n4932;
assign n1488 = ~(n243 ^ n4863);
assign n12893 = ~(n4802 ^ n1149);
assign n7596 = ~(n931 ^ n7543);
assign n2537 = ~(n8357 ^ n6865);
assign n7041 = ~n2339;
assign n2486 = n1671 & n11642;
assign n10752 = ~(n10651 ^ n6876);
assign n2744 = ~n11096;
assign n12027 = n9048 | n3635;
assign n13223 = ~(n8407 ^ n4247);
assign n3333 = n9962 | n9195;
assign n1668 = n5799 & n9645;
assign n550 = n4086 & n6064;
assign n4529 = ~(n2908 | n6060);
assign n1478 = ~(n4244 | n5961);
assign n10477 = ~(n1507 ^ n7097);
assign n11778 = ~(n8560 ^ n5672);
assign n7977 = ~n8970;
assign n13042 = ~(n2164 ^ n7090);
assign n4441 = n6056 | n12164;
assign n1150 = n8556 | n10871;
assign n11435 = ~(n9559 ^ n9704);
assign n4436 = ~(n11526 ^ n12347);
assign n11721 = n10603 | n6540;
assign n6680 = ~n9732;
assign n4820 = ~(n1185 ^ n5059);
assign n8928 = n11379 | n8841;
assign n11159 = ~(n294 ^ n6648);
assign n2538 = ~n10408;
assign n4040 = n1635 | n1572;
assign n2987 = n6487 ^ n826;
assign n7371 = ~n11872;
assign n11837 = ~(n6385 ^ n2836);
assign n10583 = ~(n12790 | n9807);
assign n12927 = ~(n6933 | n7562);
assign n11823 = ~n1176;
assign n1486 = n4822 & n830;
assign n5454 = n2965 ^ n6704;
assign n3301 = ~n2962;
assign n10203 = ~n11201;
assign n9349 = n2799 | n2451;
assign n4872 = ~(n1351 ^ n4205);
assign n9997 = n8720 | n3703;
assign n1671 = ~n10547;
assign n5600 = n11729 | n8348;
assign n8116 = n265 & n6657;
assign n438 = ~n1007;
assign n5398 = ~(n9432 ^ n9263);
assign n13110 = n333 | n2222;
assign n1516 = n1962 & n3685;
assign n6876 = ~(n11070 ^ n3503);
assign n5582 = n11094 | n8490;
assign n6948 = ~(n2418 ^ n2139);
assign n7794 = n5923 | n7935;
assign n9302 = ~(n12719 | n10778);
assign n7110 = ~n6574;
assign n6750 = ~n2734;
assign n4971 = n4257 & n12988;
assign n1566 = n12510 & n619;
assign n10871 = n4517;
assign n5578 = ~(n10683 ^ n12393);
assign n9702 = ~n5758;
assign n3476 = ~(n7549 ^ n3380);
assign n1313 = n5303 | n2032;
assign n7032 = n11797 & n12311;
assign n5370 = n12052 | n6635;
assign n4020 = n10716 & n9813;
assign n2246 = n5010 & n8943;
assign n9494 = n1353 | n1144;
assign n77 = ~(n4007 ^ n6665);
assign n10174 = n39 | n3103;
assign n2028 = ~n7273;
assign n11424 = n4558 | n1811;
assign n8110 = ~(n10713 ^ n1692);
assign n1748 = ~(n12030 ^ n6748);
assign n7102 = ~n12683;
assign n4497 = n4157 | n4326;
assign n3031 = ~n12953;
assign n240 = n4496 | n1247;
assign n6195 = ~(n3037 ^ n11390);
assign n11377 = ~(n12633 ^ n8309);
assign n4677 = n2598 | n13151;
assign n12902 = n4372 | n1678;
assign n11170 = n4719 & n1096;
assign n12432 = n79 | n4640;
assign n4650 = ~(n4624 | n11495);
assign n9551 = ~(n7975 ^ n7523);
assign n4415 = n12004 & n7738;
assign n3549 = n12848 & n9466;
assign n1595 = n8115 & n11041;
assign n1363 = ~(n7225 ^ n12359);
assign n6822 = n367 | n12566;
assign n8960 = n6402 & n9918;
assign n10164 = ~(n10674 ^ n6837);
assign n13216 = n12054 | n5392;
assign n1494 = n10383 | n7723;
assign n7792 = n333 | n10956;
assign n8987 = ~n5989;
assign n3267 = ~(n4444 ^ n8589);
assign n7273 = n13174 & n1596;
assign n13165 = n5568 & n10451;
assign n1207 = n11466 | n10106;
assign n12308 = ~n7035;
assign n3298 = n8971 & n8936;
assign n7767 = ~(n11828 | n3452);
assign n2713 = n4291 | n2562;
assign n12686 = ~n9124;
assign n9029 = n2250 | n10701;
assign n6127 = ~(n2829 ^ n8128);
assign n12586 = ~(n1098 | n2311);
assign n2323 = ~n10134;
assign n8912 = ~n11061;
assign n4313 = n7419 ^ n9619;
assign n515 = ~(n4673 | n292);
assign n3048 = n10026 & n4542;
assign n897 = n5037 & n9651;
assign n6299 = ~(n8271 ^ n10626);
assign n12296 = n9310 | n1571;
assign n4478 = n13077 | n4640;
assign n5058 = ~n11850;
assign n2930 = ~n4426;
assign n8775 = ~n3365;
assign n6318 = n4693 | n814;
assign n5111 = n9614 | n1581;
assign n8416 = n10476 | n10126;
assign n10591 = ~n7720;
assign n10355 = n1887 | n8348;
assign n7827 = ~n3693;
assign n10615 = n4206 & n9023;
assign n7878 = ~n7659;
assign n6320 = n2377 | n6860;
assign n6350 = ~(n11705 ^ n4662);
assign n7576 = ~(n966 ^ n7336);
assign n4852 = n1096 | n4719;
assign n8221 = n8487 | n11822;
assign n159 = ~n8150;
assign n2289 = n8904 | n8030;
assign n5086 = ~n103;
assign n12220 = n10591 | n8534;
assign n115 = ~n499;
assign n10567 = ~(n7147 ^ n397);
assign n11911 = ~(n5185 | n1734);
assign n11080 = n2872 | n10029;
assign n6156 = ~n3042;
assign n10303 = ~(n13081 ^ n11263);
assign n9063 = ~(n9188 ^ n1815);
assign n3715 = n10783 & n125;
assign n4816 = ~n4285;
assign n2720 = n7493 & n2553;
assign n903 = ~(n8402 ^ n2783);
assign n7314 = ~(n11486 ^ n9410);
assign n11256 = n8161 & n6651;
assign n3139 = n3572 | n10352;
assign n2475 = ~(n1523 ^ n6197);
assign n11420 = n3225 | n6732;
assign n8902 = ~(n1411 ^ n476);
assign n11294 = n13201 & n11058;
assign n7595 = n5031 & n287;
assign n7820 = n6005 & n1150;
assign n8799 = n7730 | n650;
assign n11145 = ~(n11423 ^ n3408);
assign n9483 = n2321 | n3999;
assign n12753 = ~(n7958 | n5864);
assign n9701 = n9510 & n11525;
assign n6917 = ~n745;
assign n422 = n3284 | n6813;
assign n10395 = ~(n10026 ^ n9802);
assign n8487 = n8744 | n4179;
assign n6109 = ~(n2112 ^ n8501);
assign n5662 = n10127 & n6645;
assign n13013 = ~n937;
assign n8879 = n11333 | n2942;
assign n9975 = ~(n7702 ^ n5989);
assign n13191 = ~n6948;
assign n727 = n8406 & n6076;
assign n11814 = n10304 & n9517;
assign n6199 = ~(n3481 | n9338);
assign n10284 = n2095 | n11810;
assign n11334 = ~(n12696 ^ n648);
assign n10979 = n7119 | n12328;
assign n9328 = n6125 | n9608;
assign n10845 = n7550 | n9518;
assign n653 = n2280 & n11102;
assign n172 = n8843 | n12501;
assign n2750 = ~(n10889 ^ n4425);
assign n4921 = n7011 | n7117;
assign n12262 = n2296 | n10029;
assign n11593 = ~n6650;
assign n71 = n784 & n2433;
assign n12840 = n6355 | n1696;
assign n7364 = ~(n10625 | n10160);
assign n6103 = ~(n4023 ^ n474);
assign n1380 = ~(n2016 | n2050);
assign n11148 = ~n4382;
assign n1107 = ~(n1798 ^ n420);
assign n10786 = ~n8675;
assign n5483 = n3178 & n5548;
assign n7961 = ~n1364;
assign n7403 = n6245 | n3698;
assign n3562 = ~(n8156 ^ n10170);
assign n10060 = n6309 | n6037;
assign n945 = ~(n5269 ^ n4939);
assign n563 = n7102 & n1054;
assign n8556 = ~n12306;
assign n8267 = ~(n5942 ^ n7334);
assign n24 = n11536 | n911;
assign n11657 = ~(n11407 ^ n9550);
assign n6884 = ~(n1854 ^ n1273);
assign n9647 = n9557 | n4686;
assign n2000 = ~(n7840 ^ n9435);
assign n9374 = ~(n5230 ^ n9636);
assign n12512 = n998 & n11125;
assign n562 = ~(n3929 | n1853);
assign n11206 = ~(n3057 ^ n10863);
assign n10541 = n6225 | n5414;
assign n2969 = n7429 & n9567;
assign n11393 = ~(n12143 | n3793);
assign n8176 = ~n8768;
assign n6050 = ~(n12451 ^ n2402);
assign n1701 = n1278 | n3712;
assign n11029 = ~n1876;
assign n8663 = ~n10697;
assign n3789 = ~(n502 ^ n11588);
assign n9091 = n1584 & n11572;
assign n11879 = ~(n9418 ^ n1057);
assign n12568 = ~n497;
assign n9383 = ~n5356;
assign n13202 = ~(n6021 | n1186);
assign n9576 = ~(n4239 ^ n11570);
assign n759 = ~n2939;
assign n7892 = ~(n4731 ^ n5790);
assign n4606 = ~n12488;
assign n10858 = ~n12609;
assign n1841 = n2148 | n1043;
assign n5700 = n10017 | n12388;
assign n2239 = ~(n6799 ^ n7826);
assign n2913 = ~(n8356 ^ n456);
assign n10065 = n2677 | n10912;
assign n604 = ~(n6015 | n7602);
assign n3352 = n3225 | n10900;
assign n7639 = ~(n11791 ^ n269);
assign n1810 = ~(n9951 ^ n3495);
assign n4646 = ~(n10537 ^ n5049);
assign n549 = ~n1254;
assign n4372 = n7821 & n5039;
assign n6399 = n13000 & n8981;
assign n5972 = ~(n3958 ^ n2846);
assign n11940 = ~n8466;
assign n4062 = ~(n10004 | n3358);
assign n381 = ~(n6657 ^ n265);
assign n2168 = n7467 | n2249;
assign n3538 = n12432 & n3417;
assign n435 = n5767 | n6589;
assign n1162 = ~(n6015 ^ n1529);
assign n1067 = ~n7613;
assign n8732 = n476 & n1411;
assign n3045 = n2232 | n6814;
assign n11291 = ~n9300;
assign n11831 = ~(n214 | n4378);
assign n2790 = n1212 & n13061;
assign n10980 = n11130 & n5208;
assign n6459 = ~(n9567 ^ n7429);
assign n7392 = ~(n2337 ^ n8277);
assign n5852 = ~(n11343 ^ n4595);
assign n3278 = n10582 & n11887;
assign n2029 = ~(n1310 ^ n5632);
assign n3260 = n12948 | n6265;
assign n8597 = n11706 & n1379;
assign n5020 = n10366 & n10328;
assign n2127 = n10566 & n11877;
assign n4704 = n8998 | n12132;
assign n12538 = ~(n13203 ^ n5487);
assign n10639 = ~(n12313 ^ n522);
assign n1247 = n3079 & n4251;
assign n9119 = ~n11059;
assign n7344 = n4668 & n12726;
assign n12339 = n10860 & n1347;
assign n12265 = ~(n147 ^ n10094);
assign n3654 = ~(n6082 | n12542);
assign n6802 = n5164 | n7412;
assign n5185 = ~(n4971 ^ n6597);
assign n5800 = ~(n13184 ^ n6891);
assign n2970 = ~n10642;
assign n2167 = n11643 & n7378;
assign n345 = ~(n4157 ^ n2317);
assign n2551 = ~n9929;
assign n12581 = n10530 & n12938;
assign n2259 = n3940 | n2637;
assign n2868 = n941 & n12599;
assign n9552 = n1241 | n11817;
assign n7424 = ~n4141;
assign n935 = ~n287;
assign n8677 = n4478 & n1599;
assign n6756 = ~n4597;
assign n4157 = n4077 | n9638;
assign n7998 = ~n9475;
assign n6959 = n12790 & n9807;
assign n3309 = ~(n12567 ^ n8465);
assign n4134 = n1125 | n4606;
assign n8637 = n6739 & n9279;
assign n5668 = n12592 & n3076;
assign n3389 = ~(n8031 ^ n4450);
assign n8032 = n7324 & n6682;
assign n631 = ~(n7298 ^ n8266);
assign n5983 = n7195 & n311;
assign n5766 = ~n9856;
assign n3774 = n6407 | n6732;
assign n10207 = ~(n8208 ^ n3873);
assign n2564 = n13201 & n9915;
assign n9725 = n11347 | n824;
assign n6763 = ~(n2335 ^ n12892);
assign n1416 = ~n5320;
assign n1672 = ~n5780;
assign n480 = ~(n6701 ^ n7844);
assign n11440 = ~(n6427 ^ n5886);
assign n781 = n7247 | n10059;
assign n12614 = n1571 | n2718;
assign n9643 = ~(n96 | n10390);
assign n11020 = n1790 | n11686;
assign n4839 = ~(n5552 ^ n7367);
assign n260 = ~(n11874 | n2716);
assign n6511 = n12795 | n8490;
assign n8551 = ~(n1940 ^ n11880);
assign n6599 = ~(n1862 | n6180);
assign n11733 = ~(n12833 ^ n4005);
assign n11039 = n2254 | n8534;
assign n7357 = n1587 | n3890;
assign n7503 = n6724 | n7221;
assign n5226 = ~n2498;
assign n2477 = ~(n4572 ^ n981);
assign n9588 = n3553 | n4640;
assign n11738 = ~n4847;
assign n12465 = ~n5189;
assign n3239 = ~n11390;
assign n12013 = n12104 & n12018;
assign n12191 = n2338 | n13148;
assign n10195 = ~n9684;
assign n966 = ~(n11095 ^ n11243);
assign n11271 = ~(n232 ^ n1870);
assign n13180 = ~(n9082 ^ n9687);
assign n4327 = ~(n10672 ^ n11442);
assign n11116 = ~(n6899 | n7214);
assign n3948 = ~(n8361 ^ n6162);
assign n9768 = ~(n1988 ^ n6143);
assign n4242 = ~(n8981 | n13000);
assign n4678 = n9195 | n1144;
assign n202 = ~n12306;
assign n8787 = n4727 | n13196;
assign n7028 = ~(n1727 ^ n4060);
assign n10878 = n1370 | n4640;
assign n1616 = n10527 | n12188;
assign n1980 = ~(n7313 ^ n3500);
assign n12157 = ~(n2020 | n5267);
assign n10236 = ~(n10081 ^ n7282);
assign n8187 = n8182 | n3716;
assign n11317 = ~(n8770 ^ n2284);
assign n12205 = n8938 & n8164;
assign n2314 = n7667 ^ n12961;
assign n10746 = n4149 & n7147;
assign n3061 = ~(n11530 ^ n9589);
assign n4455 = ~n2771;
assign n4540 = ~n7113;
assign n1633 = ~(n1826 | n9871);
assign n7762 = n11780 & n5869;
assign n1859 = ~(n6345 ^ n8879);
assign n9499 = n12730 & n6525;
assign n7228 = ~(n1540 | n8150);
assign n1602 = n11800 & n5424;
assign n7318 = n5865 | n4947;
assign n2770 = ~(n1578 ^ n8597);
assign n4431 = ~(n7480 | n11052);
assign n5492 = ~(n4066 | n12622);
assign n11735 = n10123 & n10822;
assign n2649 = n13097 & n1577;
assign n12550 = n3130 & n12284;
assign n81 = n11581 | n3328;
assign n541 = n10947 & n2862;
assign n6556 = n6283 | n11173;
assign n7683 = ~n5889;
assign n282 = n13165 & n8322;
assign n4978 = n5845 ^ n8084;
assign n3053 = n12051 & n2086;
assign n11546 = n11682 ^ n5355;
assign n6741 = n8803 | n2903;
assign n856 = n3646 | n12273;
assign n8113 = n10973 & n4153;
assign n1076 = n10447 | n4979;
assign n2362 = n6024 | n4915;
assign n9871 = ~n10627;
assign n4025 = n2028 & n5468;
assign n1662 = n693 & n11453;
assign n9890 = ~(n8648 ^ n8774);
assign n3114 = n9832 & n3683;
assign n12373 = ~(n7437 ^ n6762);
assign n12954 = ~n5801;
assign n6230 = ~(n12698 | n2051);
assign n10976 = ~(n11944 ^ n4299);
assign n6114 = ~(n10505 ^ n6161);
assign n5926 = n8863 | n4640;
assign n3319 = n11554 | n1156;
assign n11310 = n5431 & n440;
assign n4432 = n4464 | n4640;
assign n1056 = n6914 | n9615;
assign n3682 = n9017 | n7723;
assign n6013 = ~(n10820 ^ n10763);
assign n12951 = ~(n11327 | n394);
assign n13197 = ~(n1891 ^ n10084);
assign n804 = n1644 & n12646;
assign n97 = ~n9887;
assign n4439 = ~(n12511 ^ n2966);
assign n7363 = ~(n4659 ^ n11507);
assign n9894 = n7135 | n7075;
assign n10230 = ~n10294;
assign n12477 = ~(n4231 ^ n2073);
assign n10114 = ~n39;
assign n1760 = ~(n2426 ^ n9912);
assign n8333 = ~(n5912 ^ n1982);
assign n6870 = n7084 | n2675;
assign n9222 = ~(n9925 ^ n6361);
assign n1808 = ~(n1394 ^ n3233);
assign n8673 = n425 & n6205;
assign n1994 = ~(n1286 ^ n2617);
assign n4022 = ~n12693;
assign n11154 = n5031 & n1916;
assign n5157 = ~n1364;
assign n8010 = n464 | n1466;
assign n13064 = ~(n4560 ^ n12923);
assign n2662 = n3434 & n4021;
assign n10250 = ~n9535;
assign n999 = ~(n4857 ^ n9735);
assign n9705 = n8225 | n1985;
assign n2338 = ~n9906;
assign n6629 = ~n3641;
assign n3405 = ~(n5151 | n7843);
assign n10931 = n9428 ^ n13173;
assign n11248 = n5569 | n4373;
assign n404 = ~(n704 ^ n11516);
assign n977 = n8174 | n9075;
assign n6412 = n9581 | n4230;
assign n8681 = ~n7374;
assign n9001 = n115 | n10871;
assign n7587 = ~(n2794 | n1467);
assign n13186 = ~n12121;
assign n10409 = ~(n11274 ^ n10559);
assign n4201 = ~n3677;
assign n10632 = ~(n4879 ^ n563);
assign n6690 = n8492 & n6120;
assign n7216 = ~n1724;
assign n1921 = n8453 & n4825;
assign n5832 = ~n6873;
assign n7493 = n9909 | n7803;
assign n11856 = ~(n4211 | n7095);
assign n1571 = n438;
assign n4685 = n8173 | n121;
assign n5475 = ~(n5647 ^ n1837);
assign n12075 = ~(n8080 | n10140);
assign n9004 = ~(n3106 ^ n7276);
assign n10885 = n2685 & n7889;
assign n10581 = n6984 & n1297;
assign n808 = ~n5320;
assign n8472 = ~n4862;
assign n12983 = ~(n9082 | n13074);
assign n3604 = ~(n8949 ^ n6637);
assign n8375 = n8401 & n337;
assign n8062 = ~(n10416 | n11030);
assign n2593 = ~(n5833 ^ n10370);
assign n12661 = n1938 ^ n12932;
assign n5227 = n3563 | n11870;
assign n1978 = n2449 | n8702;
assign n12616 = ~(n3372 ^ n7577);
assign n10389 = n2493 & n4203;
assign n5479 = ~n3894;
assign n12798 = ~n10019;
assign n3475 = ~(n10247 ^ n2756);
assign n11643 = ~n7516;
assign n10945 = ~(n2389 ^ n2051);
assign n2842 = n12224 | n1144;
assign n10103 = ~n61;
assign n3454 = ~n8230;
assign n5073 = n8978 & n9733;
assign n9070 = ~n3192;
assign n9399 = n5871 ^ n8974;
assign n492 = n2015 & n1701;
assign n9054 = n13073 | n3426;
assign n1031 = ~(n529 ^ n8705);
assign n10251 = ~(n9375 ^ n10204);
assign n12966 = n10512 ^ n5827;
assign n4562 = n1998 & n5357;
assign n4773 = n5214 & n4330;
assign n1317 = ~(n6418 | n1738);
assign n295 = n7219 & n7222;
assign n2608 = n172 | n4973;
assign n4003 = n11227 & n2676;
assign n5354 = n3078 & n6952;
assign n12395 = ~n8183;
assign n484 = n9810 | n542;
assign n3089 = ~(n605 | n11395);
assign n4769 = ~(n710 ^ n3376);
assign n9758 = ~(n3117 ^ n7457);
assign n304 = ~(n6144 | n11621);
assign n4368 = ~(n6643 ^ n2845);
assign n2084 = ~(n6465 ^ n9647);
assign n3363 = n8621 | n9935;
assign n6824 = ~(n11824 | n10658);
assign n2401 = n8173 | n12395;
assign n326 = ~(n1988 | n10035);
assign n2128 = ~(n4937 ^ n6192);
assign n3960 = n5231 & n7227;
assign n3002 = ~(n10456 ^ n7664);
assign n7117 = n3293 | n947;
assign n470 = n7354 | n5743;
assign n7459 = n1718 | n7567;
assign n6316 = n3407 | n1026;
assign n7888 = ~n11123;
assign n7221 = n11940;
assign n7313 = n9729 ^ n6758;
assign n7918 = n10005 | n10117;
assign n9234 = n10465 | n1463;
assign n6284 = n723 & n10506;
assign n8390 = n5683 | n12721;
assign n7906 = n121 | n1869;
assign n3635 = ~(n7328 | n6025);
assign n7469 = n11420 | n2363;
assign n1404 = n9760 & n11392;
assign n780 = ~(n4742 ^ n3837);
assign n12696 = ~(n10344 ^ n70);
assign n233 = n621 | n3246;
assign n2481 = n4400 & n12285;
assign n545 = ~n5594;
assign n3291 = ~(n1901 ^ n11874);
assign n1953 = n8466 & n8233;
assign n6899 = n7906;
assign n4801 = ~(n7131 ^ n11136);
assign n8524 = n5748 & n11221;
assign n200 = n8361 | n6162;
assign n2871 = n9949 & n11889;
assign n12547 = ~(n386 ^ n3369);
assign n2570 = n12836 | n1819;
assign n409 = ~(n10613 | n10711);
assign n511 = n2872 | n9159;
assign n4682 = n10981 & n5187;
assign n3724 = ~n11953;
assign n10850 = ~(n6717 ^ n291);
assign n5826 = n12490 | n2059;
assign n1237 = n2018 & n854;
assign n5828 = n2329 | n1026;
assign n5100 = ~(n3914 ^ n8503);
assign n5424 = n5905 & n6727;
assign n8271 = n11537 & n9915;
assign n6895 = ~(n7774 ^ n11355);
assign n3929 = ~(n12270 | n12076);
assign n10077 = n8306 | n11982;
assign n10354 = n5913 & n6412;
assign n7006 = n10908 & n8468;
assign n2282 = n845 | n8563;
assign n11568 = ~(n10850 ^ n1486);
assign n5293 = ~(n8674 ^ n1403);
assign n3467 = n12357 | n13133;
assign n11599 = n3281 | n3981;
assign n7572 = n4267 & n6152;
assign n9018 = ~n11906;
assign n6355 = ~n817;
assign n2643 = n11871 | n3225;
assign n8193 = n6481 | n3651;
assign n8777 = ~n5962;
assign n3229 = n5004 & n4314;
assign n6016 = n11542 | n12695;
assign n940 = n712 | n9136;
assign n10385 = n8210 & n10310;
assign n13108 = ~n761;
assign n196 = ~n8134;
assign n3936 = n5086 | n1741;
assign n6906 = ~n4687;
assign n879 = n1823 | n7704;
assign n758 = ~(n3715 ^ n8831);
assign n2650 = ~(n2196 ^ n1295);
assign n4910 = ~n6244;
assign n4272 = ~n11350;
assign n11620 = n10317 | n12361;
assign n12138 = n10752 & n10666;
assign n10540 = ~(n1219 | n4567);
assign n8890 = n5694 | n5242;
assign n752 = n3428 | n12695;
assign n3625 = ~(n40 ^ n7873);
assign n350 = n1588 & n12536;
assign n2664 = ~(n8328 ^ n10434);
assign n4602 = n1335 | n1089;
assign n8100 = ~(n2911 ^ n11506);
assign n8440 = n12294 | n7435;
assign n7611 = n2443 & n11641;
assign n403 = ~(n6892 ^ n9952);
assign n10981 = n8495 | n8929;
assign n4064 = n9104 & n4852;
assign n2244 = ~(n862 ^ n7895);
assign n2232 = ~n4862;
assign n10456 = ~(n8080 ^ n1576);
assign n909 = n1757 & n3409;
assign n3917 = ~(n10242 | n10050);
assign n11309 = ~(n8683 ^ n10208);
assign n10915 = ~(n5690 | n4032);
assign n10171 = n6412 | n5913;
assign n5070 = n379 | n12273;
assign n6542 = ~(n11063 ^ n8862);
assign n9931 = ~n12482;
assign n6705 = ~(n13054 ^ n12084);
assign n12604 = ~n9620;
assign n11381 = n7160 & n4374;
assign n10099 = n7688 | n12524;
assign n6776 = n3115 | n597;
assign n5290 = n10032 | n8030;
assign n7864 = ~n2072;
assign n10833 = ~(n3001 ^ n12179);
assign n5115 = n5146 | n3981;
assign n4460 = n12274 & n5111;
assign n918 = ~(n2900 ^ n6793);
assign n10309 = ~(n1655 | n1482);
assign n7438 = n44 | n3981;
assign n5937 = ~(n3730 ^ n9932);
assign n2030 = n4943 & n2124;
assign n1744 = ~n8203;
assign n5027 = n89 & n1813;
assign n1822 = ~(n1481 | n7848);
assign n4667 = ~(n11490 ^ n6282);
assign n11748 = n7658 & n8512;
assign n4539 = n12560 ^ n7854;
assign n11071 = ~(n472 ^ n5260);
assign n7691 = n13024 & n6887;
assign n2734 = ~(n11663 ^ n8269);
assign n2556 = ~n8506;
assign n23 = ~(n4629 ^ n2643);
assign n5824 = ~(n2874 ^ n8635);
assign n8391 = ~n2501;
assign n12734 = ~n5371;
assign n6760 = ~n13076;
assign n9226 = ~(n6822 ^ n10776);
assign n1580 = ~(n12130 | n12181);
assign n9609 = n19 & n3549;
assign n9687 = ~(n4074 ^ n6232);
assign n9691 = n2165 | n5409;
assign n12972 = n1943 | n12519;
assign n6123 = n1052 | n8563;
assign n8040 = ~n4933;
assign n12759 = n6454 & n1975;
assign n1901 = ~n10459;
assign n9799 = ~(n4934 | n5084);
assign n7684 = n5163 | n5242;
assign n1049 = ~(n2260 ^ n4446);
assign n447 = n6671 & n6441;
assign n5269 = ~(n5213 | n12687);
assign n8586 = n3687 & n1800;
assign n9204 = n3157 | n8206;
assign n2844 = n3705 ^ n5938;
assign n7366 = n6629 | n1985;
assign n8128 = n7649 & n7031;
assign n3264 = n4114 & n11222;
assign n10323 = ~(n2187 | n2612);
assign n2948 = n5562 | n3981;
assign n11153 = n10018 | n121;
assign n588 = ~n1393;
assign n10487 = ~(n5020 | n1512);
assign n11772 = ~n8230;
assign n1733 = ~n12627;
assign n522 = ~(n2193 ^ n4167);
assign n5268 = ~n1160;
assign n1006 = n235 | n4285;
assign n13229 = ~n5543;
assign n12234 = ~n7336;
assign n13227 = ~(n9161 ^ n1726);
assign n4638 = n1361 | n6910;
assign n9695 = n5890 | n4373;
assign n7552 = ~(n10731 ^ n7540);
assign n2728 = n11722 | n7502;
assign n4054 = n6526 | n1951;
assign n55 = ~(n1223 ^ n8189);
assign n6529 = ~(n10479 ^ n4522);
assign n10597 = ~n6654;
assign n5840 = n2834 | n5298;
assign n1867 = n11303 | n4990;
assign n9802 = ~(n4542 ^ n12259);
assign n646 = ~(n7696 ^ n13230);
assign n4825 = n9889 & n4841;
assign n6193 = ~n8716;
assign n9895 = n5974 & n3655;
assign n8595 = ~(n1306 | n1682);
assign n2041 = ~n5729;
assign n4990 = ~(n4789 | n8467);
assign n13034 = ~(n9158 ^ n2288);
assign n7304 = n4338 & n13093;
assign n7484 = n11542 | n4373;
assign n5777 = ~(n1489 ^ n5281);
assign n8819 = n9284 & n11660;
assign n1178 = n9702 | n3225;
assign n11124 = n12473 | n2530;
assign n9109 = n8758 | n10285;
assign n1475 = ~(n8590 ^ n3035);
assign n2624 = n2111 | n3162;
assign n8343 = ~(n6042 | n6829);
assign n6322 = ~(n1074 ^ n4893);
assign n6979 = n1268 | n6885;
assign n9965 = n3514 & n8191;
assign n12673 = ~n3040;
assign n10961 = n6979 & n57;
assign n11703 = n9389 | n5061;
assign n8962 = ~(n5385 ^ n8636);
assign n2227 = n2542 | n2287;
assign n7512 = ~(n6947 ^ n4511);
assign n1360 = ~n4998;
assign n9615 = n534 & n5416;
assign n11051 = ~(n7782 ^ n13038);
assign n11845 = ~(n12861 ^ n6440);
assign n12678 = ~(n10296 ^ n5145);
assign n4709 = n1252 ^ n13165;
assign n7661 = ~n2882;
assign n5247 = n7856 | n9873;
assign n5172 = n12772 | n4991;
assign n6431 = ~(n61 ^ n9896);
assign n7326 = ~(n4392 ^ n12893);
assign n2915 = ~n7515;
assign n9696 = ~(n591 | n7554);
assign n10984 = ~(n11862 ^ n4129);
assign n10562 = ~(n6235 ^ n8802);
assign n5873 = ~(n7162 ^ n3672);
assign n10628 = ~(n8071 ^ n7799);
assign n6142 = ~n10799;
assign n3659 = ~(n6530 ^ n9758);
assign n7963 = ~n1497;
assign n1440 = n8724 | n12064;
assign n2894 = ~(n6855 ^ n8832);
assign n11394 = ~(n3175 ^ n10769);
assign n5079 = ~n9187;
assign n878 = n26 & n1239;
assign n3738 = ~(n10220 ^ n5387);
assign n11897 = ~(n6349 ^ n11309);
assign n802 = ~(n12457 | n2810);
assign n7677 = ~(n7573 ^ n9219);
assign n11595 = n4986 | n4694;
assign n6709 = ~(n3657 ^ n7650);
assign n8330 = n11049 ^ n4320;
assign n12190 = n1286 | n12736;
assign n11040 = ~n5705;
assign n12485 = ~(n9969 ^ n6249);
assign n7907 = ~n4909;
assign n939 = n8230 & n9531;
assign n10996 = ~(n8396 | n11383);
assign n6978 = n8871 & n7139;
assign n5490 = ~n11190;
assign n12364 = ~(n524 ^ n5617);
assign n12785 = n1285 & n12055;
assign n11550 = n2678 | n5076;
assign n12769 = ~(n13107 ^ n5619);
assign n7970 = n7501 ^ n9063;
assign n4282 = ~(n509 ^ n4882);
assign n11977 = ~(n8099 ^ n12766);
assign n25 = ~(n4879 ^ n8760);
assign n4891 = ~n9738;
assign n11364 = ~n726;
assign n12886 = ~n1900;
assign n7651 = ~(n11118 ^ n6214);
assign n60 = ~n9636;
assign n8747 = ~(n2835 | n6833);
assign n11621 = ~n362;
assign n3379 = ~(n12574 ^ n5951);
assign n3965 = ~n12605;
assign n8579 = n1908 & n11279;
assign n6767 = n9144 | n6870;
assign n4764 = ~(n8772 ^ n506);
assign n814 = n9140 & n174;
assign n387 = ~(n1060 ^ n10159);
assign n704 = ~(n463 ^ n9961);
assign n10245 = ~n4828;
assign n5461 = ~n11537;
assign n9703 = ~(n10051 | n1140);
assign n13164 = ~(n1903 ^ n8375);
assign n7334 = ~(n5892 ^ n2030);
assign n3017 = ~n8715;
assign n10020 = n8510 | n12718;
assign n8915 = n11472 | n6882;
assign n11503 = n5360 ^ n7970;
assign n1433 = n9482 & n12323;
assign n9978 = n4109 | n964;
assign n11839 = ~(n2034 ^ n11150);
assign n9125 = ~n11673;
assign n12577 = ~(n7688 ^ n12524);
assign n8108 = ~n1165;
assign n12943 = n12595 & n1881;
assign n5395 = ~(n8846 ^ n4440);
assign n10918 = n3126 | n2958;
assign n783 = ~n8841;
assign n11921 = ~(n2432 ^ n3521);
assign n2587 = ~(n3964 ^ n6879);
assign n5128 = ~(n3568 ^ n5641);
assign n220 = ~(n3679 ^ n7600);
assign n11189 = ~(n8157 ^ n9576);
assign n742 = ~(n11012 | n3674);
assign n12700 = n4397 & n8165;
assign n12814 = ~n4862;
assign n11098 = ~(n7795 | n3803);
assign n12924 = ~(n10114 | n11332);
assign n11360 = n9316 | n10072;
assign n7291 = ~n5729;
assign n6913 = ~n5185;
assign n11554 = ~(n12661 | n10321);
assign n6229 = n6407 | n6404;
assign n11759 = ~n5389;
assign n5613 = n9289 | n7831;
assign n11542 = ~n9846;
assign n7170 = n321 | n10319;
assign n1863 = ~(n10183 | n1949);
assign n8516 = ~(n7959 ^ n2529);
assign n10314 = ~n2737;
assign n10302 = ~(n11645 | n2);
assign n8351 = ~n1764;
assign n8449 = n10914 | n7185;
assign n2940 = ~(n7862 ^ n7166);
assign n13224 = ~(n678 ^ n166);
assign n7150 = ~(n612 | n9986);
assign n7890 = ~n5470;
assign n6780 = ~(n2962 ^ n1415);
assign n89 = ~n6675;
assign n8381 = n5445 | n5681;
assign n6628 = ~(n12843 ^ n8988);
assign n6138 = ~n7539;
assign n5619 = ~(n5280 | n8439);
assign n8976 = ~(n1418 ^ n10875);
assign n5383 = ~n8887;
assign n7741 = ~n12853;
assign n5880 = ~(n11715 ^ n2968);
assign n7047 = ~(n10120 | n346);
assign n8828 = ~(n2550 | n9472);
assign n10267 = ~(n6754 | n8094);
assign n6024 = n2449 | n6404;
assign n2383 = n3532 | n9190;
assign n8376 = n11957 & n4958;
assign n10347 = ~(n10817 ^ n8067);
assign n2433 = n11851 | n157;
assign n2851 = ~(n12545 ^ n6631);
assign n2568 = ~(n8124 | n4262);
assign n11068 = n8987 & n3508;
assign n3552 = ~n1503;
assign n11382 = n1688 | n1463;
assign n1225 = ~(n7611 ^ n6570);
assign n12048 = ~(n8714 | n11853);
assign n8465 = ~(n6336 ^ n8752);
assign n4609 = ~(n695 | n7483);
assign n8619 = n8599 | n6468;
assign n12332 = n6875 | n4373;
assign n10593 = n12914 | n5917;
assign n7939 = ~n9138;
assign n7249 = ~n6385;
assign n5194 = n7135 | n9195;
assign n3979 = ~(n7064 | n4250);
assign n6454 = ~(n1598 ^ n2273);
assign n8363 = ~n3321;
assign n273 = ~(n11674 ^ n7092);
assign n8052 = n12412 & n4174;
assign n5495 = ~(n1764 | n2213);
assign n8469 = n1594 & n7337;
assign n2236 = n7880 | n4230;
assign n11027 = n12225 | n9012;
assign n6301 = ~(n11452 ^ n6815);
assign n3722 = n2057 & n2882;
assign n1941 = ~n6149;
assign n11307 = n10499 | n6893;
assign n1649 = ~n11816;
assign n12779 = ~(n8882 ^ n1850);
assign n1670 = ~(n1240 ^ n12630);
assign n3935 = n2581 | n13108;
assign n1605 = ~n951;
assign n3886 = ~(n8229 | n4633);
assign n1807 = ~n10548;
assign n3490 = n6488 | n12388;
assign n11251 = n8179 | n7140;
assign n7856 = n8400 | n5242;
assign n3029 = n1325 | n5423;
assign n2 = n4365 & n2507;
assign n3271 = n3932 & n7015;
assign n13075 = n6132 | n8783;
assign n3558 = n6378 & n9325;
assign n11131 = n2386 & n6899;
assign n5767 = n11274 & n12993;
assign n2853 = n6928 & n1711;
assign n5012 = ~(n12976 ^ n4341);
assign n7243 = ~n8288;
assign n8626 = ~n12916;
assign n8186 = n7376 | n2455;
assign n1880 = ~(n8565 ^ n4938);
assign n5618 = ~(n13093 ^ n2436);
assign n12496 = n5611 | n2544;
assign n7957 = n2963 & n8010;
assign n4234 = ~(n3496 ^ n12862);
assign n157 = n9854 & n11193;
assign n3349 = ~(n3594 ^ n4632);
assign n5746 = ~n6904;
assign n7902 = n10045 | n7935;
assign n12704 = n9905 & n173;
assign n871 = ~n12085;
assign n2136 = ~n1130;
assign n6337 = n9730 | n11479;
assign n5066 = ~n7710;
assign n12239 = ~(n12162 ^ n511);
assign n12484 = ~n5408;
assign n836 = n10279 ^ n9447;
assign n3819 = ~n10563;
assign n9587 = ~(n1284 ^ n12369);
assign n5698 = ~(n10073 ^ n731);
assign n12892 = ~(n2913 ^ n10747);
assign n9676 = ~(n3307 ^ n11326);
assign n6364 = ~n11488;
assign n1951 = ~(n2937 ^ n7764);
assign n8599 = n5949 | n4230;
assign n5351 = n6883 | n4947;
assign n11003 = ~n3264;
assign n193 = ~n2220;
assign n6604 = n81 & n9884;
assign n3764 = ~n9898;
assign n5234 = n9430 & n2579;
assign n9824 = ~(n1866 ^ n2075);
assign n5179 = n10780 | n8348;
assign n7008 = n7862 & n9861;
assign n4248 = n2418 & n9945;
assign n12385 = ~(n729 | n4700);
assign n1423 = ~(n6280 ^ n8121);
assign n11617 = n10901 | n10687;
assign n2303 = ~(n8489 ^ n7853);
assign n6068 = n10587 | n10871;
assign n3663 = ~(n11997 ^ n10062);
assign n12285 = n6129 | n9075;
assign n8948 = ~n7895;
assign n8798 = ~(n2433 ^ n5064);
assign n6922 = ~n11350;
assign n2145 = ~n938;
assign n10695 = ~(n5131 ^ n10397);
assign n8358 = n7950 | n4936;
assign n7835 = ~(n8957 ^ n581);
assign n7951 = n1207 | n7008;
assign n11708 = n9161 & n6372;
assign n4397 = n7372 | n4107;
assign n284 = ~(n11283 ^ n349);
assign n8770 = n12249 | n5242;
assign n2936 = ~(n3027 | n3717);
assign n4210 = ~(n484 ^ n960);
assign n1129 = ~(n2776 ^ n6201);
assign n3751 = ~(n1682 ^ n4347);
assign n7776 = n12434 | n479;
assign n5099 = ~n3354;
assign n11754 = n895 & n1639;
assign n1312 = n1296 | n4936;
assign n4021 = n4540 | n1463;
assign n992 = n10230 | n8283;
assign n8576 = n2264 | n11144;
assign n1771 = n8139 & n6826;
assign n5864 = n8693 & n709;
assign n11357 = n12528 | n2694;
assign n13038 = ~(n11915 ^ n4133);
assign n8539 = n1416 | n8868;
assign n2837 = ~(n5503 ^ n1452);
assign n2855 = ~(n2842 ^ n9484);
assign n681 = ~(n1173 | n3628);
assign n6252 = ~(n2016 ^ n9685);
assign n9473 = ~(n10811 ^ n10008);
assign n10557 = ~(n3045 | n8577);
assign n6840 = n1729 & n6745;
assign n7447 = ~(n8671 ^ n1624);
assign n3667 = ~(n4681 ^ n11979);
assign n797 = n10527 | n1463;
assign n8231 = ~n346;
assign n7093 = n9967 & n1442;
assign n815 = n313 & n4212;
assign n11994 = n569 | n2544;
assign n3293 = ~n9475;
assign n9742 = ~(n2585 ^ n11238);
assign n7287 = n971 | n5242;
assign n2682 = ~(n5307 ^ n709);
assign n8490 = n2557;
assign n5597 = n9069 | n8534;
assign n5482 = ~(n6165 | n2448);
assign n9810 = ~n401;
assign n3274 = ~(n8223 ^ n6520);
assign n5718 = ~(n7953 ^ n2871);
assign n6144 = ~n6603;
assign n12045 = ~n1771;
assign n3338 = ~n4043;
assign n12618 = ~(n11924 ^ n7609);
assign n5874 = n4209 | n7846;
assign n3448 = n4043 ^ n1171;
assign n9694 = ~(n1620 ^ n2743);
assign n11570 = n4722 | n8563;
assign n7816 = ~(n9731 ^ n674);
assign n4151 = ~(n8675 ^ n6429);
assign n9141 = n12674 & n1001;
assign n12202 = ~(n11084 | n4931);
assign n10886 = ~n11324;
assign n2349 = ~(n12218 ^ n10283);
assign n4133 = n9266 & n5822;
assign n4659 = n9808 | n542;
assign n12228 = ~(n7982 ^ n3426);
assign n7 = n6033 | n13242;
assign n1866 = ~(n2496 ^ n6696);
assign n6593 = ~(n12662 ^ n6691);
assign n436 = ~n10048;
assign n8134 = n10958 | n792;
assign n2625 = ~n13014;
assign n7482 = ~(n5700 ^ n8278);
assign n4147 = ~(n11281 | n4702);
assign n9083 = n2129 | n12062;
assign n11184 = ~(n10001 ^ n6673);
assign n5707 = ~n4885;
assign n7575 = n9924 ^ n5668;
assign n4572 = ~(n3797 ^ n4705);
assign n7082 = ~n4249;
assign n1393 = ~(n8924 ^ n3439);
assign n1250 = n9767 | n9195;
assign n1195 = ~(n11717 ^ n8608);
assign n11193 = n7422 | n9178;
assign n10524 = ~(n5253 ^ n4860);
assign n4081 = n6638 | n6635;
assign n10412 = n9511 | n8348;
assign n4202 = ~(n170 ^ n12547);
assign n7380 = ~(n5354 | n1831);
assign n1567 = ~(n1683 ^ n12557);
assign n11978 = ~(n299 | n967);
assign n13128 = n11284 | n1043;
assign n5816 = ~(n7747 ^ n1183);
assign n12351 = ~(n2568 | n1608);
assign n9806 = n11114 | n12188;
assign n5595 = ~n8332;
assign n4083 = ~(n10847 ^ n10061);
assign n7693 = ~(n10806 | n1489);
assign n11878 = n11861 | n8016;
assign n5425 = n5146 | n5242;
assign n11419 = n10859 | n8209;
assign n5314 = n5935 | n4854;
assign n12334 = ~(n6248 ^ n1016);
assign n12093 = ~n9887;
assign n9650 = ~n1734;
assign n5108 = n2971 | n6684;
assign n10050 = ~(n7850 | n3329);
assign n11380 = n5163 | n9223;
assign n6583 = ~(n7028 ^ n10542);
assign n10332 = ~n4439;
assign n11791 = ~(n7497 | n3386);
assign n8355 = n8629 | n1161;
assign n6450 = ~(n6750 ^ n7653);
assign n10361 = ~n1758;
assign n12960 = ~(n12703 ^ n13046);
assign n7451 = ~(n11714 ^ n1772);
assign n8659 = n12155 | n10362;
assign n3337 = n3382 & n10640;
assign n5545 = n7401 | n7855;
assign n2321 = ~n3311;
assign n11094 = ~n12372;
assign n266 = n5787 & n735;
assign n7476 = ~(n12619 ^ n6115);
assign n6217 = n533 | n1287;
assign n9163 = ~(n10153 ^ n9183);
assign n163 = ~(n7463 | n11884);
assign n8397 = n790 | n12419;
assign n1066 = ~(n2227 ^ n7126);
assign n5405 = ~(n4757 ^ n11450);
assign n26 = ~n4747;
assign n3512 = ~(n6299 ^ n1882);
assign n5158 = ~n2343;
assign n5297 = ~(n5380 | n6524);
assign n6091 = n12656 & n10807;
assign n10801 = ~(n11698 ^ n7492);
assign n9426 = n12495 & n4772;
assign n3078 = ~n8149;
assign n62 = ~(n9334 ^ n8456);
assign n11675 = ~(n4614 ^ n8014);
assign n5015 = n1989 | n7377;
assign n9693 = ~n8689;
assign n1641 = ~(n1939 ^ n381);
assign n9822 = n12665 & n11091;
assign n5289 = ~n2731;
assign n4612 = ~n12065;
assign n922 = ~(n7957 ^ n9566);
assign n6005 = n6858 & n3665;
assign n4254 = ~(n5998 ^ n724);
assign n12723 = ~(n8328 | n12508);
assign n11368 = ~(n4651 | n10210);
assign n4377 = n8661 & n7529;
assign n11385 = n12462 | n5092;
assign n131 = ~(n12237 ^ n9506);
assign n4914 = ~(n10348 ^ n7590);
assign n1375 = n13036 | n10871;
assign n1016 = ~(n120 ^ n12028);
assign n6029 = n8412 | n273;
assign n6830 = n2002 | n2308;
assign n3976 = ~(n1984 ^ n4483);
assign n4457 = n9706 & n412;
assign n685 = n5038 | n11368;
assign n9935 = ~(n4128 ^ n9982);
assign n10078 = n7715 & n3409;
assign n3585 = ~(n10774 | n11777);
assign n2983 = ~(n10238 ^ n6286);
assign n7848 = n343 & n9750;
assign n4997 = ~(n6835 ^ n3476);
assign n2641 = ~n10805;
assign n3068 = ~n2341;
assign n285 = ~(n12632 | n3990);
assign n7478 = ~(n9970 ^ n8625);
assign n9654 = n7087 ^ n3008;
assign n5138 = n13231 | n6128;
assign n11450 = n1695 | n6635;
assign n6987 = n11213 & n11241;
assign n5018 = n7925 | n5242;
assign n5879 = ~(n6455 ^ n2724);
assign n1299 = ~(n10799 ^ n4097);
assign n13077 = ~n9093;
assign n9035 = n11184 & n7503;
assign n12126 = ~n9531;
assign n9356 = n11933 | n8702;
assign n121 = n12335;
assign n8891 = n3498 | n905;
assign n8041 = n2961 & n9142;
assign n3714 = n12732 | n9075;
assign n4465 = ~n287;
assign n10701 = n11065 & n8708;
assign n269 = ~(n12505 | n9787);
assign n9193 = ~(n1265 ^ n8804);
assign n7535 = ~(n1628 | n3202);
assign n2445 = n2469 & n2383;
assign n6982 = n6850 & n4229;
assign n4775 = ~(n7235 ^ n7703);
assign n1428 = n2670 | n546;
assign n2395 = ~(n3942 ^ n3089);
assign n621 = n1040 & n5564;
assign n8078 = n609 & n4677;
assign n6140 = n10168 & n12263;
assign n7714 = ~(n636 | n9365);
assign n6559 = ~n11134;
assign n11562 = n493 | n1144;
assign n5341 = ~n7036;
assign n13059 = n5120 & n8474;
assign n8294 = ~(n8052 ^ n11038);
assign n9116 = ~(n8422 | n7407);
assign n7360 = ~(n6311 ^ n11568);
assign n9084 = n6710 | n1197;
assign n10440 = ~n3438;
assign n1692 = n5957 & n8808;
assign n6578 = ~n12186;
assign n6966 = ~n9258;
assign n3913 = n8637 ^ n10569;
assign n10397 = ~(n2079 ^ n11153);
assign n2830 = ~(n7580 ^ n4985);
assign n3446 = ~(n786 ^ n5484);
assign n13172 = n9340 & n142;
assign n2078 = ~(n1742 ^ n6893);
assign n1241 = n12410 & n2802;
assign n11070 = ~(n1443 ^ n6496);
assign n1858 = ~n4636;
assign n7470 = n12575 | n5623;
assign n13195 = n7481 & n10644;
assign n1111 = n7686 & n4508;
assign n4166 = ~n1198;
assign n3536 = n9245 & n12866;
assign n6943 = n406 | n11446;
assign n10279 = n9628 & n7459;
assign n4555 = n2512 & n12237;
assign n5330 = ~(n1481 ^ n11848);
assign n5805 = ~n5605;
assign n11128 = ~(n7601 | n3779);
assign n10804 = n5540 & n1917;
assign n6512 = n1056 & n3582;
assign n9782 = n10281 | n2675;
assign n9589 = ~(n2492 ^ n250);
assign n8076 = ~(n6763 | n10440);
assign n1236 = ~n7378;
assign n645 = ~n4570;
assign n12434 = ~n8522;
assign n9006 = ~(n2072 ^ n12283);
assign n4404 = ~(n8970 ^ n12701);
assign n3299 = ~n7061;
assign n5140 = ~(n2912 ^ n4900);
assign n2831 = n7707 | n4947;
assign n7197 = n9712 & n1592;
assign n5082 = ~n8794;
assign n3033 = n8081 & n13191;
assign n4974 = ~n6655;
assign n5641 = ~(n13169 ^ n3083);
assign n9013 = n8940 & n287;
assign n8263 = n8039 | n360;
assign n9221 = n10586 | n1199;
assign n10144 = n2720 | n4160;
assign n1327 = n11076 ^ n412;
assign n12629 = ~n1198;
assign n9509 = n11736 | n2695;
assign n5663 = ~(n141 | n13195);
assign n10265 = n13116 | n3709;
assign n1796 = n4654 | n1958;
assign n3822 = n3972 | n11152;
assign n8695 = n5220 & n11636;
assign n4079 = n2437 | n6652;
assign n2035 = ~(n3270 ^ n13143);
assign n5183 = ~(n11374 ^ n9025);
assign n10609 = n7900 | n8030;
assign n12492 = ~(n5553 ^ n3);
assign n365 = n9397 | n9319;
assign n10922 = ~(n8803 ^ n12787);
assign n7589 = n6343 | n10788;
assign n10832 = n1732 & n10502;
assign n2558 = ~(n8760 | n3209);
assign n12594 = ~(n2262 ^ n4535);
assign n8883 = n6271 | n7723;
assign n7746 = ~(n3285 | n7381);
assign n7944 = ~(n12252 | n5573);
assign n9533 = ~(n10318 | n530);
assign n12307 = ~(n12681 ^ n6685);
assign n1827 = n694 | n12717;
assign n11032 = n7244 & n7933;
assign n8779 = n737 | n6404;
assign n1962 = n3713 | n7962;
assign n6658 = ~n6023;
assign n355 = ~(n12168 | n1890);
assign n1718 = n3431 ^ n9717;
assign n4308 = n8254 | n11107;
assign n3054 = n9131 | n8030;
assign n12006 = ~(n6508 ^ n4199);
assign n3879 = n7265 & n8789;
assign n7699 = n7742 | n5076;
assign n5811 = n3809 | n2290;
assign n5519 = ~(n9817 ^ n4014);
assign n9604 = ~(n4130 | n1627);
assign n7441 = n1779 | n10132;
assign n10137 = ~n11222;
assign n1572 = ~(n6990 | n974);
assign n11255 = n3425 & n1028;
assign n11974 = ~n25;
assign n7022 = n3419 | n2035;
assign n2274 = ~(n12867 ^ n11079);
assign n7879 = ~(n9819 ^ n10555);
assign n9085 = n9693 | n4325;
assign n4239 = n12009 | n9223;
assign n7793 = ~(n11050 ^ n11401);
assign n11747 = n25 ^ n10724;
assign n1977 = n12049 | n7935;
assign n5271 = ~n11634;
assign n5940 = n12456 | n7180;
assign n11653 = n11356 | n177;
assign n11764 = ~(n4502 ^ n9458);
assign n7514 = ~(n7841 ^ n5149);
assign n5814 = n11653 | n13042;
assign n9730 = ~n2555;
assign n3865 = ~(n12042 ^ n4256);
assign n79 = ~n9531;
assign n9974 = ~(n1299 ^ n8312);
assign n7206 = ~(n2371 ^ n3269);
assign n2999 = n5563 | n11032;
assign n3958 = n3761 | n1014;
assign n11074 = ~(n11780 ^ n11758);
assign n2201 = ~(n9363 | n1566);
assign n12908 = ~n6987;
assign n8098 = ~n1683;
assign n2491 = n477 | n5024;
assign n5717 = n9240 | n7002;
assign n9460 = ~n9115;
assign n4805 = n10113 & n7113;
assign n7721 = ~(n3659 | n8260);
assign n12073 = ~(n12740 ^ n1748);
assign n8615 = ~n8233;
assign n6270 = ~(n9534 | n3192);
assign n9904 = n10966 | n2958;
assign n433 = n5248 | n10299;
assign n11150 = n7868 | n8348;
assign n11750 = ~n4889;
assign n12495 = ~(n551 ^ n2142);
assign n206 = n2557;
assign n10008 = ~n836;
assign n10196 = n11547 | n3689;
assign n10318 = ~n5972;
assign n10272 = ~n10630;
assign n11638 = n12919 & n10533;
assign n340 = ~(n1888 ^ n3464);
assign n489 = n7501 | n11359;
assign n2749 = ~(n1200 | n7645);
assign n1956 = n10837 & n1015;
assign n9493 = n7563 & n7794;
assign n12654 = n9873 & n7856;
assign n12398 = ~(n4262 ^ n8124);
assign n5122 = n2500 | n1371;
assign n5888 = n4473 | n8490;
assign n12929 = ~(n2980 ^ n794);
assign n9432 = ~(n2978 | n10443);
assign n3520 = ~(n11671 | n9062);
assign n1998 = ~n3887;
assign n7821 = n9540 ^ n9510;
assign n7616 = n7914 & n12949;
assign n8558 = n4964 & n1916;
assign n6061 = ~(n7117 ^ n7170);
assign n12662 = ~(n1775 ^ n6316);
assign n2986 = ~(n5272 ^ n5856);
assign n5295 = n11127 & n2355;
assign n11023 = ~(n4379 | n2897);
assign n11985 = n4997 | n3237;
assign n5284 = n1511 | n7935;
assign n3989 = ~(n6071 ^ n10829);
assign n7795 = ~(n12322 | n12374);
assign n9148 = ~n8916;
assign n8934 = ~n11217;
assign n9958 = ~(n7236 ^ n2099);
assign n8462 = n8042 & n2533;
assign n516 = n1319 | n3984;
assign n2552 = n7607 & n3501;
assign n673 = n4220 | n4360;
assign n10006 = n12656 | n10807;
assign n6546 = ~(n5888 ^ n9549);
assign n4742 = ~n10105;
assign n12677 = n7880 | n8348;
assign n3924 = ~n4023;
assign n8601 = n2473 | n11770;
assign n586 = n1449 & n7852;
assign n7510 = n2468 | n12489;
assign n5528 = n5959 | n12889;
assign n13166 = ~(n7686 ^ n12436);
assign n4683 = ~(n3741 | n3551);
assign n10672 = ~(n5680 | n7200);
assign n10427 = n928 | n3287;
assign n10793 = ~n13020;
assign n7058 = ~(n5929 ^ n10215);
assign n5655 = n107 | n5049;
assign n11629 = n4657 | n6404;
assign n11223 = n6008 & n10268;
assign n6196 = n8251 & n12821;
assign n4183 = ~(n6511 ^ n10943);
assign n10023 = n9955 | n10570;
assign n7521 = n12940 & n7496;
assign n5142 = n12982 | n3497;
assign n3018 = n5990 | n4230;
assign n6989 = ~(n6382 | n10175);
assign n13137 = ~(n10113 | n1757);
assign n6928 = n1977 | n9149;
assign n3313 = n8249 | n6635;
assign n5982 = ~(n6618 | n10986);
assign n11969 = ~n12923;
assign n4892 = ~(n8749 ^ n8761);
assign n5134 = n10944 | n6706;
assign n6585 = n2057 & n3076;
assign n8508 = ~n8155;
assign n9479 = n227 | n8268;
assign n6781 = ~(n5794 ^ n11753);
assign n3354 = n11157 | n1463;
assign n5029 = ~(n10485 | n11856);
assign n8149 = ~(n4905 ^ n7757);
assign n6429 = ~(n376 ^ n3921);
assign n4192 = n7084 | n9784;
assign n1512 = ~(n11912 | n9715);
assign n219 = ~(n6065 | n10852);
assign n6925 = n12856 & n6821;
assign n2468 = n1714 & n1475;
assign n12741 = ~n13060;
assign n696 = ~(n2479 ^ n5078);
assign n7880 = ~n5536;
assign n11466 = ~n4006;
assign n11492 = ~(n9869 ^ n7168);
assign n3364 = ~n5758;
assign n3737 = ~(n10967 ^ n13189);
assign n2155 = n5937 | n4165;
assign n971 = ~n389;
assign n4131 = ~(n10339 | n7005);
assign n2619 = ~n4281;
assign n9329 = ~(n91 ^ n9196);
assign n8616 = ~(n6610 ^ n4069);
assign n9988 = ~n824;
assign n140 = ~(n2881 ^ n2751);
assign n9762 = n3231 & n4175;
assign n12763 = n10237 & n6472;
assign n4067 = ~(n5502 | n11452);
assign n998 = ~(n8629 ^ n1852);
assign n824 = n9157 & n11595;
assign n5730 = ~(n7666 ^ n2984);
assign n7813 = n4524 & n9697;
assign n6845 = n13062 | n6176;
assign n9372 = n37 & n5224;
assign n1661 = n1329 | n7723;
assign n1584 = n3166 & n8687;
assign n6627 = n9930 | n3980;
assign n9957 = ~(n1699 ^ n3731);
assign n9566 = ~(n8351 ^ n2213);
assign n865 = n10622 ^ n13157;
assign n12325 = ~(n10056 | n1668);
assign n826 = n2306 & n9247;
assign n6692 = ~(n3510 | n11906);
assign n11927 = ~n12390;
assign n5369 = n2619 | n8012;
assign n3154 = ~(n4764 ^ n7138);
assign n3835 = n8937 & n1141;
assign n8115 = n8795 | n2959;
assign n11728 = n2479 | n8292;
assign n10494 = ~(n6205 ^ n425);
assign n10748 = ~n8954;
assign n561 = ~n3144;
assign n1333 = ~n5984;
assign n5559 = ~n4691;
assign n8697 = ~n10867;
assign n7984 = ~(n3478 ^ n10464);
assign n195 = ~(n5577 ^ n12251);
assign n11757 = ~n22;
assign n1382 = ~(n3988 ^ n2445);
assign n1622 = ~(n32 ^ n4020);
assign n6408 = n4521 & n13099;
assign n11669 = ~(n31 ^ n5051);
assign n4925 = ~(n7435 ^ n7088);
assign n1869 = ~n854;
assign n9052 = ~(n5513 ^ n10251);
assign n2512 = ~(n11233 ^ n7736);
assign n2571 = ~(n4277 | n3046);
assign n12500 = n4298 | n8582;
assign n3478 = n5461 | n6769;
assign n471 = ~(n9401 ^ n3930);
assign n5191 = ~(n1493 | n8624);
assign n7114 = n644 | n7152;
assign n9021 = ~(n9835 ^ n804);
assign n9546 = n11633 & n5829;
assign n6089 = n12336 & n1267;
assign n181 = n588 | n7585;
assign n9224 = n7110 | n9052;
assign n1104 = n3381 | n4819;
assign n1889 = ~n11049;
assign n2962 = n8666 & n6204;
assign n10256 = ~n4470;
assign n10367 = n10717 & n12874;
assign n13061 = ~(n2771 ^ n6168);
assign n6090 = ~(n8785 ^ n197);
assign n6008 = ~n13006;
assign n8419 = ~n7932;
assign n9170 = ~n8713;
assign n468 = ~(n3744 ^ n9184);
assign n6999 = n5412 & n10340;
assign n2220 = n1058 | n12847;
assign n8247 = ~(n7421 | n981);
assign n3119 = ~(n6794 | n5812);
assign n1510 = ~(n548 ^ n2369);
assign n8867 = ~(n2151 ^ n105);
assign n3897 = ~(n10905 ^ n3626);
assign n12944 = n9396 | n9311;
assign n5588 = ~n10594;
assign n8157 = n11683 | n11144;
assign n8463 = ~n10142;
assign n4229 = n4271 | n9348;
assign n4094 = n11078 | n7837;
assign n10435 = n1145 | n10892;
assign n10266 = ~n12605;
assign n11067 = n5675 & n4559;
assign n7787 = ~n5453;
assign n7128 = n10402 | n10319;
assign n3234 = ~(n10785 ^ n429);
assign n3839 = n11447 & n12765;
assign n11756 = n5069 & n123;
assign n9536 = ~(n4663 ^ n8056);
assign n10855 = ~(n7920 | n11034);
assign n6623 = ~(n12039 ^ n4182);
assign n4844 = ~n10606;
assign n6914 = n7668 & n8074;
assign n13041 = n4785 | n7615;
assign n6359 = n10462 | n4724;
assign n6452 = n552 | n3376;
assign n263 = n971 | n2958;
assign n7644 = ~(n7690 ^ n199);
assign n3382 = n4290 | n6364;
assign n11287 = ~(n8812 | n5287);
assign n12980 = n6155 ^ n10670;
assign n6825 = ~n11112;
assign n3020 = n5194 | n5272;
assign n11033 = n8529 | n6404;
assign n1000 = ~n1600;
assign n7608 = ~n13060;
assign n1286 = n11096 ^ n12424;
assign n8097 = ~n2920;
assign n9677 = ~n3121;
assign n6601 = n7561 & n4970;
assign n2223 = n8379 | n5273;
assign n9540 = n2420 | n2287;
assign n5376 = ~(n1507 | n3519);
assign n11046 = ~(n2184 ^ n5486);
assign n8861 = ~(n6688 ^ n8471);
assign n4042 = n7791 & n6469;
assign n92 = ~(n823 ^ n7928);
assign n11037 = ~n5065;
assign n6660 = ~(n1398 ^ n1946);
assign n5754 = ~(n6359 ^ n4255);
assign n10534 = ~(n7709 | n3165);
assign n7410 = ~n8735;
assign n3110 = n5249 & n3614;
assign n838 = ~(n6021 ^ n8227);
assign n4759 = n391 | n12978;
assign n6555 = ~(n3171 ^ n9665);
assign n7790 = ~(n10904 ^ n10777);
assign n9522 = ~(n8881 ^ n3596);
assign n12764 = n9162 | n8702;
assign n8013 = ~(n6740 ^ n9141);
assign n9878 = n5152 | n4495;
assign n5334 = n5990 | n7221;
assign n6309 = ~n11900;
assign n3077 = n182 | n5295;
assign n885 = ~(n477 ^ n8554);
assign n5859 = ~(n3441 | n6909);
assign n996 = n5670 | n7642;
assign n4232 = n11946 & n11481;
assign n12110 = ~(n2043 ^ n5995);
assign n13043 = ~n9941;
assign n5806 = ~n1724;
assign n6816 = ~(n7546 ^ n3610);
assign n4961 = ~(n8864 | n2422);
assign n539 = n4594 & n7588;
assign n4730 = ~(n2304 | n10961);
assign n1491 = n8455 ^ n2229;
assign n6387 = n7599 & n9037;
assign n4244 = n2883 & n1506;
assign n11918 = n7041 | n8348;
assign n661 = n373 & n12309;
assign n11659 = n3628 & n1173;
assign n7234 = ~n12263;
assign n4993 = ~(n7575 ^ n8145);
assign n9466 = n5870 & n528;
assign n7737 = ~(n577 | n2117);
assign n1405 = ~(n7095 ^ n9117);
assign n4162 = ~(n2792 ^ n12911);
assign n3791 = ~n10811;
assign n12442 = n12384 & n7383;
assign n5775 = n2769 & n9660;
assign n308 = ~n2539;
assign n3107 = ~(n11865 ^ n4895);
assign n12901 = n7890 | n10761;
assign n5077 = n3839 | n11346;
assign n10862 = n4021 | n3434;
assign n12987 = ~(n2940 ^ n5741);
assign n6665 = ~(n1095 ^ n9028);
assign n4635 = n8882 | n1850;
assign n13071 = ~n4349;
assign n13086 = ~n11537;
assign n12120 = n9590 & n6509;
assign n2535 = ~(n10373 ^ n10091);
assign n5195 = ~(n3050 ^ n3170);
assign n4390 = n10462 | n2133;
assign n7254 = ~n11488;
assign n7752 = n11941 | n8348;
assign n7649 = n11159 | n10040;
assign n4070 = ~(n9641 | n4873);
assign n4578 = ~(n11444 ^ n3198);
assign n8014 = ~(n455 ^ n5104);
assign n12857 = ~(n9830 ^ n4283);
assign n9251 = ~(n6505 | n13037);
assign n8786 = ~n862;
assign n7292 = ~(n1807 | n6281);
assign n8245 = n2332 | n177;
assign n10311 = n9933 & n7193;
assign n10906 = n8672 | n9195;
assign n8341 = ~n11079;
assign n10087 = ~(n5181 ^ n9295);
assign n2865 = ~(n5102 ^ n4051);
assign n4072 = n5695 | n7339;
assign n6216 = n4850 & n2499;
assign n8302 = n755 | n12967;
assign n12761 = ~(n10774 ^ n5779);
assign n4681 = ~(n10547 ^ n7323);
assign n5583 = ~n3152;
assign n12233 = n11137 | n10319;
assign n4979 = ~n6168;
assign n7678 = ~n12025;
assign n7875 = ~(n2435 ^ n12554);
assign n11848 = ~(n9750 ^ n504);
assign n11239 = ~n9531;
assign n9439 = n2736 | n2659;
assign n11254 = n13001 & n5155;
assign n3013 = n12786 | n8534;
assign n8061 = n5595 | n7530;
assign n7959 = n3945 & n10495;
assign n9655 = n2482 & n12853;
assign n8949 = n13012 | n12188;
assign n2821 = n8183 & n6085;
assign n9248 = ~(n2813 ^ n4691);
assign n8648 = n935 | n2133;
assign n4100 = ~(n4377 ^ n5439);
assign n1222 = n1801 & n2477;
assign n4490 = ~n9915;
assign n4448 = n9486 & n6738;
assign n3744 = n12469 | n12957;
assign n12131 = ~(n1580 | n9463);
assign n5298 = ~(n8651 ^ n2951);
assign n5343 = n10142 & n5962;
assign n13112 = n11336 & n5318;
assign n10022 = n6016 | n8782;
assign n1832 = ~n6879;
assign n7024 = ~(n5233 ^ n12934);
assign n6956 = n10761 | n4936;
assign n2191 = n1795 | n8543;
assign n3932 = n11196 | n9533;
assign n7394 = n2992 & n11262;
assign n1839 = ~(n3749 ^ n801);
assign n2672 = n11576 & n8839;
assign n12974 = n2902 & n1189;
assign n8424 = n7191 | n5939;
assign n4056 = ~(n1025 | n4482);
assign n1140 = ~(n12229 ^ n4019);
assign n1787 = ~n10002;
assign n1948 = ~(n10538 ^ n5650);
assign n10964 = n667 | n5693;
assign n13014 = n4981 | n9110;
assign n9649 = n8060 | n3229;
assign n9452 = ~(n3458 ^ n2964);
assign n10664 = ~(n12204 | n12235);
assign n12206 = n4039 | n9188;
assign n12312 = n12483 | n4194;
assign n40 = ~(n6013 ^ n5232);
assign n11196 = ~(n159 ^ n6154);
assign n10414 = n5200 & n12979;
assign n12842 = n11624 & n5338;
assign n2517 = ~(n6310 | n4414);
assign n12329 = ~(n6460 ^ n5362);
assign n10796 = ~(n12707 ^ n10699);
assign n9279 = n12092 | n10982;
assign n10716 = n1925 | n4407;
assign n9120 = n2480 & n5877;
assign n6000 = n3354 | n6730;
assign n8423 = ~(n8742 | n4816);
assign n1608 = n5665 & n8454;
assign n5803 = n1589 | n2133;
assign n9344 = n5732 & n5504;
assign n5236 = ~(n7697 ^ n4615);
assign n5067 = n151 & n7078;
assign n5455 = ~n11429;
assign n9301 = ~(n10865 | n1004);
assign n4628 = n7437 & n12124;
assign n8162 = ~(n1469 | n7054);
assign n8006 = ~n5969;
assign n5898 = n2742 | n90;
assign n11059 = n2085 & n2149;
assign n4174 = n5322 | n5222;
assign n10772 = ~n12965;
assign n3753 = n10437 | n11107;
assign n10066 = ~n7945;
assign n7185 = ~(n9508 | n10910);
assign n3369 = ~(n3192 ^ n8515);
assign n2942 = ~n11061;
assign n1252 = n7642 | n479;
assign n2363 = n9305 | n10179;
assign n5468 = ~n11991;
assign n7193 = n2884 | n5797;
assign n546 = ~n6236;
assign n4761 = n9402 | n4333;
assign n3836 = n4179 | n2059;
assign n5500 = n2460 & n4750;
assign n547 = ~(n7161 | n1144);
assign n12818 = n10233 & n6218;
assign n1126 = ~n9097;
assign n8927 = n1222 | n10239;
assign n10739 = ~n2023;
assign n5789 = ~(n11711 | n41);
assign n3833 = n5492 | n13135;
assign n7996 = n6682 ^ n6451;
assign n799 = n11512 & n4869;
assign n7461 = n6401 | n306;
assign n11535 = ~n2595;
assign n8562 = ~n3409;
assign n6057 = n349 | n11283;
assign n6225 = ~n4335;
assign n4994 = ~(n8932 ^ n9204);
assign n9157 = n689 | n4626;
assign n2373 = n823 | n4405;
assign n9258 = n3588 & n5967;
assign n11225 = ~n2174;
assign n3809 = n6222 & n3101;
assign n2638 = ~(n8920 ^ n12678);
assign n10820 = n13141 & n11088;
assign n3348 = n542 | n2675;
assign n6227 = ~(n386 | n6482);
assign n6686 = ~(n8850 ^ n632);
assign n2870 = n7385 | n12794;
assign n1053 = ~(n2975 | n12056);
assign n12948 = ~n834;
assign n771 = n9129 | n6404;
assign n5907 = n10182 & n12532;
assign n6004 = ~n4685;
assign n10434 = n8876 ^ n3180;
assign n6568 = ~n2233;
assign n9392 = n10893 | n1144;
assign n2835 = ~(n12553 | n4350);
assign n5845 = n2462 | n8563;
assign n8077 = ~n11760;
assign n10373 = n4161 | n7221;
assign n8994 = n2129 | n7221;
assign n9040 = n7243 | n11232;
assign n12668 = n12963 | n4812;
assign n12774 = n9620 & n8716;
assign n2105 = n9703 | n9064;
assign n1999 = ~n2445;
assign n11881 = ~(n6467 ^ n11112);
assign n12887 = ~(n5394 ^ n4140);
assign n5423 = ~n8233;
assign n1316 = ~(n11023 | n3462);
assign n12883 = ~(n3976 ^ n1884);
assign n2296 = ~n12289;
assign n6224 = ~(n3623 ^ n8917);
assign n11732 = ~(n9258 ^ n4234);
assign n1769 = ~n12594;
assign n5447 = ~(n1494 ^ n9297);
assign n8318 = n8957 | n581;
assign n8249 = ~n5536;
assign n4660 = ~n11607;
assign n10962 = n2851 & n1072;
assign n5327 = ~(n9150 | n8743);
assign n8974 = n2068 & n11109;
assign n4016 = n7396 | n4230;
assign n5628 = ~(n1408 ^ n2239);
assign n12710 = ~(n2143 | n8527);
assign n6312 = n3827 & n5021;
assign n8563 = n3169;
assign n6087 = ~(n11371 ^ n2336);
assign n3646 = ~n3769;
assign n302 = ~(n11590 ^ n11205);
assign n9188 = ~(n8412 ^ n273);
assign n7633 = ~(n3581 | n6331);
assign n950 = ~n7448;
assign n9480 = ~(n3818 ^ n12040);
assign n8682 = ~(n11436 | n5053);
assign n6347 = ~(n12428 ^ n4435);
assign n13100 = ~(n8738 | n5997);
assign n6483 = ~(n6619 ^ n637);
assign n300 = n4464 | n11107;
assign n2522 = ~(n11223 | n3002);
assign n11101 = ~n6668;
assign n5547 = ~n9906;
assign n12572 = n8839 | n11576;
assign n2604 = ~n9412;
assign n10689 = ~n10027;
assign n11162 = ~(n12121 ^ n10458);
assign n7628 = ~(n9033 ^ n12743);
assign n864 = n761 & n11058;
assign n3720 = n11116 | n7976;
assign n795 = ~n11411;
assign n573 = n1065 ^ n7238;
assign n3340 = ~n7541;
assign n9578 = n1505 & n2482;
assign n2599 = ~n8290;
assign n8568 = ~(n12518 | n3041);
assign n4520 = ~(n7311 ^ n12438);
assign n11088 = ~n5228;
assign n5107 = ~n401;
assign n5685 = ~n9092;
assign n3314 = ~(n5523 ^ n2818);
assign n498 = n7257 & n3450;
assign n11624 = n12802 | n4295;
assign n4276 = n11226 | n10106;
assign n3709 = n8541 & n1264;
assign n534 = n12971 | n7344;
assign n12470 = n6313 & n7321;
assign n5681 = n11847 & n7469;
assign n1099 = n3553 | n2544;
assign n10219 = n1370 | n7075;
assign n12078 = n2416 | n2133;
assign n1057 = n1214 ^ n11861;
assign n4958 = n1394 | n3233;
assign n6176 = n8510 | n177;
assign n1085 = n7167 | n7935;
assign n7081 = n3453 | n5335;
assign n13228 = ~n2898;
assign n2179 = n11674 | n7092;
assign n5837 = ~(n7554 ^ n140);
assign n1836 = n2255 ^ n9652;
assign n2405 = ~(n7448 | n194);
assign n5994 = ~(n5730 ^ n6122);
assign n1610 = n2326 & n2267;
assign n7756 = ~(n8001 | n7352);
assign n1781 = ~n2668;
assign n5752 = n6769 | n6404;
assign n8106 = n11903 & n5765;
assign n2919 = ~n834;
assign n8876 = n12343 & n768;
assign n2420 = ~n2758;
assign n1435 = n7119 | n1570;
assign n8021 = ~(n7245 ^ n7007);
assign n6523 = n1976 & n7586;
assign n12534 = ~(n4215 ^ n3983);
assign n477 = ~(n4016 ^ n843);
assign n10053 = n997 & n970;
assign n7668 = ~(n7279 ^ n4532);
assign n405 = n9569 & n10746;
assign n9745 = ~n287;
assign n5093 = n5801 & n9475;
assign n4514 = ~n3130;
assign n2017 = ~(n1847 | n10090);
assign n12979 = ~(n2918 ^ n7259);
assign n3880 = n5705 ^ n10078;
assign n5080 = ~n635;
assign n10732 = ~(n3219 | n739);
assign n6184 = n2678 | n9195;
assign n2257 = n6503 | n310;
assign n8888 = n8139 & n5920;
assign n7565 = n11437 | n10693;
assign n4278 = n4886 & n7810;
assign n4399 = n8704 & n10529;
assign n7975 = n9305 | n7530;
assign n3323 = ~(n486 ^ n1341);
assign n2269 = n1234 | n1934;
assign n9428 = n10761 | n10433;
assign n6974 = n946 | n1985;
assign n8461 = ~(n8125 ^ n1138);
assign n12180 = ~n3860;
assign n12479 = n12592 & n2882;
assign n595 = ~(n10384 | n384);
assign n10713 = n4132 | n12847;
assign n8918 = n2204 & n1546;
assign n283 = n13062 & n6176;
assign n9406 = ~(n3155 | n8656);
assign n4901 = n1524 | n9778;
assign n1010 = ~(n1862 ^ n1283);
assign n5945 = ~(n10859 ^ n11631);
assign n8327 = n12899 & n7710;
assign n10894 = n9806 | n7224;
assign n6946 = n11195 | n10110;
assign n6718 = ~(n10543 ^ n10955);
assign n3212 = ~(n2160 ^ n6198);
assign n1477 = ~n7359;
assign n2637 = ~n11030;
assign n10033 = ~(n6925 ^ n9394);
assign n6275 = n3669 & n3085;
assign n149 = n12159 | n8374;
assign n3207 = ~(n10198 ^ n2832);
assign n9883 = ~(n4170 ^ n1631);
assign n9908 = ~(n5331 ^ n2518);
assign n4269 = n10113 & n12853;
assign n892 = n5088 & n5814;
assign n2150 = n11899 & n383;
assign n2715 = n12592 & n11058;
assign n8724 = n1866 & n8420;
assign n9264 = n5176 | n7868;
assign n11078 = ~n6168;
assign n12362 = n12741 | n8702;
assign n2365 = ~(n5193 ^ n5643);
assign n12988 = n3829 & n11685;
assign n3355 = n12268 | n12401;
assign n11245 = n2688 | n10179;
assign n1529 = n8102 ^ n7717;
assign n13094 = ~n1983;
assign n7601 = ~(n8284 | n4543);
assign n12062 = ~n2590;
assign n628 = ~n12289;
assign n2785 = n10730 | n479;
assign n9184 = n1188 | n4230;
assign n3342 = n6333 & n10063;
assign n11794 = n7502 & n11722;
assign n1682 = ~(n10255 ^ n12985);
assign n10982 = ~n11027;
assign n12649 = ~(n7472 | n10723);
assign n12680 = ~n1660;
assign n9263 = n11523 | n6230;
assign n1159 = ~(n10786 | n7452);
assign n12177 = ~(n7051 | n12820);
assign n466 = ~(n7904 ^ n6);
assign n1819 = ~(n5453 | n9293);
assign n2722 = ~n9163;
assign n883 = n6671 | n6441;
assign n10415 = ~(n10917 ^ n4163);
assign n6220 = ~n7812;
assign n9315 = ~(n4667 ^ n7423);
assign n3777 = ~(n8595 | n7753);
assign n3954 = ~(n1714 ^ n3788);
assign n8146 = n7408 | n8869;
assign n5986 = ~(n10656 | n9292);
assign n12204 = ~n1253;
assign n6694 = n11696 & n7854;
assign n9155 = n4727 & n13196;
assign n12494 = ~(n6491 ^ n8699);
assign n4500 = ~(n12564 | n295);
assign n4603 = ~(n10533 ^ n12919);
assign n12156 = n10199 & n5579;
assign n1837 = ~(n7673 ^ n55);
assign n4297 = ~(n1679 ^ n7042);
assign n2111 = n4411 ^ n388;
assign n4255 = n2491 & n3529;
assign n2471 = n7674 | n532;
assign n3211 = n11665 & n2737;
assign n12697 = n5478 | n479;
assign n9658 = ~n2987;
assign n4190 = ~(n1279 ^ n5831);
assign n4975 = n10592 | n1404;
assign n11038 = ~(n11182 ^ n2932);
assign n1607 = n7507 | n3320;
assign n3651 = ~n3875;
assign n8628 = n5568 & n7113;
assign n4556 = ~(n12631 | n2421);
assign n8783 = ~(n11561 | n1423);
assign n5017 = ~n12245;
assign n257 = ~(n2429 ^ n7014);
assign n3365 = n5838 | n9587;
assign n12522 = ~n1535;
assign n10090 = ~n9419;
assign n8354 = n11334 & n8627;
assign n5123 = ~(n11699 ^ n4806);
assign n1728 = ~n646;
assign n9309 = ~n5536;
assign n2640 = ~n137;
assign n2214 = n10447 | n5076;
assign n5193 = ~(n7189 ^ n5195);
assign n12163 = n4605 & n4134;
assign n647 = ~(n9425 ^ n1146);
assign n10366 = ~(n5706 ^ n403);
assign n5397 = ~(n9677 ^ n2541);
assign n1420 = ~n10333;
assign n5957 = n9890 | n4343;
assign n1746 = n10306 & n5114;
assign n7316 = n3338 & n1171;
assign n6847 = n9783 & n7391;
assign n5653 = n10839 | n368;
assign n679 = n7522 | n8268;
assign n5098 = n12871 | n6265;
assign n7559 = n8310 & n7187;
assign n10419 = n6756 & n9565;
assign n6926 = n13221 ^ n78;
assign n6886 = n5968 | n8702;
assign n686 = n12881 | n9195;
assign n9683 = n592 & n914;
assign n3115 = ~(n6492 ^ n8217);
assign n4360 = ~n5596;
assign n8274 = n12636 & n7009;
assign n11293 = ~(n2920 ^ n11937);
assign n8567 = n10322 & n4604;
assign n6574 = ~(n1922 ^ n11850);
assign n9502 = n4974 | n12188;
assign n8368 = n6519 | n12273;
assign n8309 = ~(n5857 ^ n6177);
assign n7733 = n4627 & n3279;
assign n4328 = ~(n4533 | n12976);
assign n5068 = ~(n9890 ^ n8117);
assign n10009 = ~(n5956 ^ n6803);
assign n10661 = ~n5404;
assign n1060 = ~(n11773 ^ n5026);
assign n5390 = n3970 | n320;
assign n7638 = n5152 | n10552;
assign n9343 = ~(n1425 ^ n4613);
assign n4343 = n12818 & n7680;
assign n12491 = ~n608;
assign n11220 = ~(n10026 | n4542);
assign n4513 = n5047 | n10364;
assign n10138 = n12872 & n12817;
assign n6829 = n7991 & n3899;
assign n9130 = ~(n246 | n11942);
assign n9496 = n3534 | n5242;
assign n4731 = ~(n7011 ^ n6061);
assign n3632 = n6466 & n5512;
assign n10782 = ~(n5799 ^ n4721);
assign n2877 = ~n12263;
assign n776 = ~n10451;
assign n5646 = ~(n7035 ^ n4906);
assign n1689 = ~(n7110 ^ n7614);
assign n2178 = n3191 | n3423;
assign n10626 = n951 & n10063;
assign n5769 = n5365 & n8749;
assign n5208 = n12813 & n2361;
assign n9626 = ~(n10236 | n12438);
assign n3016 = ~(n7550 ^ n3948);
assign n2598 = n5611 | n9159;
assign n12796 = ~(n5669 ^ n5568);
assign n6110 = ~n649;
assign n12621 = ~n3769;
assign n2547 = n6333 & n3085;
assign n5041 = ~n10168;
assign n3618 = ~n12898;
assign n9930 = n11808 | n6770;
assign n10274 = n11272 & n5181;
assign n8572 = ~(n8467 ^ n1263);
assign n12149 = ~(n4374 ^ n7160);
assign n5871 = n12203 | n9075;
assign n11616 = n9120 & n1099;
assign n4625 = n3225 | n12388;
assign n2440 = ~n5143;
assign n1485 = ~(n6171 | n5532);
assign n12066 = ~n11267;
assign n10514 = ~(n3293 | n10866);
assign n1174 = ~(n4715 ^ n913);
assign n12144 = ~(n11335 ^ n1280);
assign n423 = ~n691;
assign n7778 = n5879 ^ n13176;
assign n7629 = n2545 | n9495;
assign n9327 = ~(n11460 ^ n4962);
assign n3457 = ~(n8165 ^ n12191);
assign n9862 = ~(n1855 ^ n11315);
assign n9563 = ~(n191 ^ n3378);
assign n1368 = ~(n11963 | n1924);
assign n7007 = ~(n4346 | n1643);
assign n3407 = ~n11396;
assign n3059 = ~(n1983 ^ n4672);
assign n6610 = n7089 & n12624;
assign n4426 = ~n9621;
assign n10104 = n5359 | n6987;
assign n5267 = ~(n8513 | n10750);
assign n6489 = n1089 | n2449;
assign n12823 = n9298 & n8127;
assign n8265 = ~(n6317 ^ n6134);
assign n8715 = n2449 | n12328;
assign n319 = ~(n7065 ^ n2526);
assign n9164 = ~(n10280 | n8649);
assign n9595 = n1260 & n8418;
assign n3853 = ~n11055;
assign n1873 = n8788 ^ n9202;
assign n3199 = n12668 & n6449;
assign n390 = n3248 | n65;
assign n4221 = ~n5470;
assign n4421 = ~(n408 | n5472);
assign n10738 = n11664 | n10715;
assign n12012 = n11003 | n8044;
assign n11091 = n8139 & n854;
assign n7985 = ~(n11836 ^ n5396);
assign n11499 = n5157 | n6769;
assign n12600 = n9146 | n11802;
assign n12743 = ~(n5843 ^ n6621);
assign n4355 = ~(n10890 | n4090);
assign n6697 = n5433 | n8348;
assign n1946 = ~(n1099 ^ n9120);
assign n7852 = n9019 | n12695;
assign n6728 = n13049 & n13115;
assign n857 = ~(n12055 ^ n12900);
assign n2789 = ~n10568;
assign n5765 = ~(n9929 ^ n5501);
assign n5745 = n1324 | n4315;
assign n12507 = ~(n7412 ^ n5164);
assign n4220 = ~n1617;
assign n1524 = ~n3303;
assign n3980 = n6883 | n10319;
assign n2148 = ~n9591;
assign n12050 = n3259 | n4936;
assign n11075 = n1034 & n12777;
assign n7458 = ~(n10262 ^ n11504);
assign n4649 = ~n5920;
assign n11739 = ~(n5127 ^ n10976);
assign n9523 = ~(n9264 ^ n2400);
assign n10321 = ~n13053;
assign n7496 = ~(n4770 ^ n5777);
assign n7763 = ~(n12192 ^ n5571);
assign n8279 = n4798 & n10519;
assign n1303 = ~(n3214 | n7173);
assign n1905 = n3599 | n773;
assign n12293 = n1052 | n3963;
assign n3125 = ~(n7944 ^ n8726);
assign n12606 = ~(n12085 | n2071);
assign n12350 = ~(n1812 ^ n3567);
assign n8084 = n5801 & n5920;
assign n5571 = n11113 | n2059;
assign n4664 = n9796 | n11794;
assign n1496 = n1696 | n1571;
assign n1290 = ~n8328;
assign n6241 = n8889 | n12068;
assign n9815 = ~(n9529 ^ n5963);
assign n6471 = ~(n878 ^ n6087);
assign n3094 = ~n6292;
assign n12023 = ~n401;
assign n10300 = ~n9446;
assign n4324 = ~(n12960 ^ n611);
assign n13118 = n7295 & n9530;
assign n2578 = n9004 | n9946;
assign n4580 = n7957 | n5495;
assign n689 = n4694 & n4986;
assign n1383 = n6335 & n6221;
assign n3210 = ~n12943;
assign n6441 = n8315 | n8348;
assign n12666 = n6556 & n4635;
assign n907 = n9675 | n12388;
assign n11744 = n8532 | n7723;
assign n1054 = n8710 | n10933;
assign n478 = n4316 & n2924;
assign n12917 = ~(n4241 | n1794);
assign n3553 = ~n12651;
assign n11175 = n11785 | n639;
assign n3050 = ~(n4159 | n11532);
assign n11709 = ~(n6962 ^ n11918);
assign n5450 = ~(n491 | n2990);
assign n579 = ~n12701;
assign n5449 = n586 | n1770;
assign n7913 = n1491 | n8242;
assign n3962 = ~n3832;
assign n6874 = n3700 & n7750;
assign n6708 = ~(n10912 ^ n572);
assign n9101 = n2420 | n9159;
assign n4793 = ~(n6880 ^ n2957);
assign n11805 = ~(n3212 ^ n918);
assign n1503 = n2777 & n9570;
assign n6796 = n12014 | n653;
assign n421 = n2848 | n1463;
assign n12997 = ~n8506;
assign n7311 = ~n10236;
assign n2390 = n5899 | n8578;
assign n10685 = ~(n3711 | n7573);
assign n11563 = ~(n6203 | n2154);
assign n12295 = ~n5065;
assign n11264 = ~(n4682 ^ n5985);
assign n3785 = ~(n10441 | n1355);
assign n3395 = n991 | n8030;
assign n9891 = ~n10643;
assign n7239 = ~n12319;
assign n10154 = n8212 | n9380;
assign n6231 = ~n3112;
assign n6940 = n10938 | n1841;
assign n4454 = ~n510;
assign n12113 = n2952 & n7444;
assign n7865 = ~n4862;
assign n7986 = ~n4711;
assign n4339 = ~n386;
assign n11752 = ~(n3011 ^ n4935);
assign n12877 = n4802 | n8493;
assign n7368 = ~(n5090 | n7638);
assign n4212 = n5766 | n6080;
assign n12804 = n11928 | n2059;
assign n3701 = n8285 & n10933;
assign n7129 = n12736 & n1286;
assign n4630 = n6707 ^ n3760;
assign n8236 = n4561 | n8607;
assign n3479 = ~(n7830 ^ n3875);
assign n8222 = ~(n12333 ^ n9194);
assign n386 = ~(n7464 ^ n4933);
assign n6048 = ~(n8134 ^ n2537);
assign n1492 = ~(n5428 | n11421);
assign n1235 = ~(n12913 ^ n10675);
assign n7372 = ~n10657;
assign n3845 = ~(n10184 ^ n3391);
assign n6711 = n1345 | n8632;
assign n12474 = ~(n10328 ^ n9715);
assign n3564 = ~n4748;
assign n101 = n2951 | n8651;
assign n3623 = n10761 | n7530;
assign n11609 = ~n10408;
assign n6152 = n7001 | n8520;
assign n11163 = n2674 | n10482;
assign n9341 = ~(n2386 ^ n12193);
assign n12915 = n10908 & n5962;
assign n11611 = ~n885;
assign n10410 = n1722 & n4393;
assign n3149 = ~n11324;
assign n9137 = n2771 & n9093;
assign n10255 = ~(n7910 ^ n13092);
assign n9089 = n6861 & n5465;
assign n11850 = ~(n1235 ^ n10494);
assign n9598 = ~(n4489 | n6462);
assign n3404 = n9867 | n10029;
assign n1522 = n12367 | n3673;
assign n12458 = ~n4331;
assign n1642 = ~(n8354 | n6319);
assign n5005 = n5713 | n9195;
assign n299 = n3392 & n7979;
assign n12685 = ~(n1150 ^ n6005);
assign n9573 = n7266 | n7060;
assign n1181 = ~(n11852 ^ n2876);
assign n9624 = n2229 & n2207;
assign n2010 = n10015 & n6608;
assign n12181 = n2641 | n12657;
assign n12822 = n8993 & n8250;
assign n6045 = n1521 | n10272;
assign n11578 = ~(n1449 ^ n6702);
assign n4688 = n7226 & n6912;
assign n13157 = n2404 & n10325;
assign n2799 = ~(n1506 ^ n2883);
assign n4679 = n1434 | n12657;
assign n9211 = n808 | n1720;
assign n9513 = n12490 | n8563;
assign n3066 = ~(n1212 ^ n4546);
assign n2703 = n5050 & n5820;
assign n9376 = ~(n1460 ^ n6050);
assign n9333 = ~(n11610 ^ n12543);
assign n4218 = n3753 | n6819;
assign n9637 = n3854 | n4936;
assign n327 = ~n9578;
assign n9099 = n9620 & n3815;
assign n5543 = n2378 & n8346;
assign n4551 = n30 & n1419;
assign n7937 = n9367 & n1357;
assign n555 = ~(n1312 ^ n12939);
assign n8831 = ~(n10613 ^ n10357);
assign n6882 = ~(n3264 | n1762);
assign n10467 = n4393 | n1722;
assign n4783 = ~n9125;
assign n2085 = n10560 & n1724;
assign n4385 = ~n5758;
assign n3972 = ~n8506;
assign n11737 = ~(n9613 ^ n12534);
assign n3525 = n7416 & n6722;
assign n5484 = n11566 & n453;
assign n4155 = ~(n3766 ^ n12890);
assign n4117 = n10916 & n11402;
assign n10088 = ~(n8911 ^ n7357);
assign n3188 = ~(n17 ^ n9327);
assign n1028 = n392 | n177;
assign n8385 = ~(n939 ^ n1971);
assign n1891 = ~(n11786 ^ n2070);
assign n10388 = n6247 | n11753;
assign n8629 = ~(n585 ^ n12835);
assign n6215 = ~n5189;
assign n9912 = ~(n3917 ^ n7631);
assign n12033 = n9563 & n12216;
assign n12158 = ~(n10365 ^ n10556);
assign n3529 = n3204 | n4729;
assign n5241 = ~(n10284 | n6959);
assign n11551 = ~(n1267 ^ n9779);
assign n9100 = ~(n5747 ^ n3006);
assign n11527 = ~(n2231 | n9295);
assign n11369 = ~n1472;
assign n711 = ~(n6647 ^ n6908);
assign n3518 = ~(n1496 | n5844);
assign n982 = ~(n2898 ^ n4688);
assign n7266 = n7905 & n359;
assign n2686 = ~(n10567 | n2131);
assign n12368 = ~n5352;
assign n10439 = ~n3832;
assign n2313 = ~(n4336 ^ n12222);
assign n7560 = ~n5197;
assign n2263 = ~n6496;
assign n2069 = ~(n12053 | n8910);
assign n12922 = n7543 | n931;
assign n12555 = n6880 | n5072;
assign n1471 = ~(n7650 | n3657);
assign n11195 = n1820 | n12273;
assign n1251 = ~n1956;
assign n1513 = ~(n1757 | n10416);
assign n2642 = ~(n7488 ^ n4738);
assign n9664 = n11053 & n4790;
assign n7541 = n6769 | n10179;
assign n6243 = n7300 & n11156;
assign n12861 = n3598 | n9195;
assign n2218 = ~(n10257 ^ n2879);
assign n3084 = n10637 & n9234;
assign n4864 = ~(n481 ^ n923);
assign n11347 = ~n6107;
assign n11479 = ~(n9123 ^ n380);
assign n1886 = n123 | n5069;
assign n11671 = ~(n9826 ^ n6090);
assign n11478 = ~(n12931 ^ n8641);
assign n2147 = ~(n10882 ^ n12906);
assign n2879 = ~(n6121 ^ n8282);
assign n732 = ~(n9597 | n9372);
assign n4295 = n2922 & n281;
assign n9816 = ~(n2523 | n6237);
assign n10759 = n6996 & n6614;
assign n13081 = n1406 | n5797;
assign n11810 = ~n8506;
assign n7046 = n4391 | n6102;
assign n135 = ~(n5903 ^ n11955);
assign n3998 = ~n8345;
assign n8694 = n11370 | n7221;
assign n2529 = ~(n11953 ^ n6048);
assign n1985 = n3058;
assign n318 = ~n9187;
assign n147 = n1587 | n11668;
assign n7204 = n1629 | n13020;
assign n2033 = ~(n5844 ^ n1496);
assign n2576 = n8582 & n4298;
assign n12933 = ~(n9142 ^ n7740);
assign n1093 = ~(n5342 ^ n2609);
assign n9097 = n2781 & n8440;
assign n10875 = ~(n3767 ^ n11257);
assign n729 = ~(n4397 ^ n3457);
assign n12786 = ~n3769;
assign n2788 = n3528 | n10918;
assign n11346 = n4189 & n1799;
assign n280 = n3460 | n10016;
assign n2808 = n8330 | n5073;
assign n9972 = ~n2037;
assign n10777 = ~(n6357 ^ n12602);
assign n7163 = ~n10013;
assign n7494 = n12028 & n120;
assign n2048 = ~n6937;
assign n2292 = n11245 | n9737;
assign n5170 = n8228 & n13058;
assign n10598 = n2993 & n10480;
assign n11543 = n7864 | n3939;
assign n43 = ~(n8571 ^ n925);
assign n5790 = ~(n1234 ^ n1934);
assign n7025 = ~n1143;
assign n117 = n1609 | n11911;
assign n893 = ~(n5007 ^ n6977);
assign n9724 = n10432 | n10403;
assign n850 = n10829 & n6071;
assign n1355 = ~(n4962 | n10810);
assign n9461 = ~n9277;
assign n8607 = n1314 & n8177;
assign n13194 = ~n4862;
assign n3824 = ~(n3706 ^ n1407);
assign n2863 = n11610 | n1456;
assign n12413 = n3404 | n10984;
assign n1156 = n1196 & n2345;
assign n7023 = n12000 | n8912;
assign n6995 = n8623 | n10581;
assign n1772 = n9016 | n1026;
assign n10694 = ~(n4926 | n5710);
assign n748 = ~(n12745 ^ n4092);
assign n5439 = n6810 | n12501;
assign n6609 = ~(n2477 ^ n1801);
assign n916 = ~(n2240 ^ n1023);
assign n398 = ~(n11217 | n9601);
assign n6403 = n12220 | n2100;
assign n12821 = n2215 & n10052;
assign n9685 = n8959 & n7106;
assign n1347 = ~n1085;
assign n5056 = ~(n7634 ^ n9442);
assign n165 = n5874 | n9122;
assign n1717 = n1548 & n4176;
assign n11960 = ~n9906;
assign n11726 = ~(n6509 ^ n9590);
assign n7141 = ~(n6155 ^ n179);
assign n10026 = n785 | n8268;
assign n6147 = ~(n3682 ^ n4259);
assign n6187 = n7028 | n2092;
assign n1295 = ~(n12531 ^ n2241);
assign n3095 = n6231 | n1043;
assign n5696 = n3835 | n10521;
assign n1444 = ~(n4711 ^ n8540);
assign n4949 = ~n11030;
assign n5175 = ~(n10869 ^ n8359);
assign n9284 = ~(n2334 ^ n2316);
assign n10656 = n2432 & n11637;
assign n11941 = ~n510;
assign n2047 = ~(n10090 ^ n3086);
assign n3217 = n6483 & n9448;
assign n10000 = ~(n608 ^ n3451);
assign n6558 = n8082 | n12388;
assign n10337 = ~(n12139 ^ n3306);
assign n3390 = n9803 & n6946;
assign n9603 = n6422 & n11260;
assign n4428 = ~(n366 ^ n301);
assign n6814 = ~n8183;
assign n9867 = ~n7659;
assign n7590 = ~(n11327 ^ n394);
assign n542 = n3185;
assign n11575 = n12434 | n2544;
assign n9850 = ~(n12341 | n7487);
assign n1319 = n11808 | n3999;
assign n2228 = ~n9915;
assign n2586 = ~(n820 ^ n4295);
assign n953 = n2748 | n7353;
assign n12226 = ~(n4117 ^ n8321);
assign n5555 = ~(n12194 ^ n7727);
assign n11469 = ~(n4650 ^ n13102);
assign n3794 = n6945 & n5108;
assign n10338 = n3714 | n8552;
assign n3614 = n6448 | n11806;
assign n10374 = n11150 & n2034;
assign n12871 = ~n10805;
assign n5616 = n1945 | n1927;
assign n5013 = n2701 | n8038;
assign n1102 = n771 | n478;
assign n2949 = n11823 & n4499;
assign n2431 = n3534 | n121;
assign n13083 = ~n9307;
assign n9176 = n4540 | n10029;
assign n1620 = ~(n4570 ^ n3600);
assign n12627 = n64 & n878;
assign n8505 = ~n11030;
assign n1033 = ~(n8550 | n13119);
assign n3131 = n10024 & n9481;
assign n5103 = n2661 | n2575;
assign n6700 = ~(n2753 ^ n10846);
assign n2061 = ~(n1637 ^ n1844);
assign n9939 = ~(n969 | n7762);
assign n5637 = ~(n4886 ^ n7810);
assign n9307 = ~(n7445 ^ n9876);
assign n11600 = n4248 | n3513;
assign n5347 = n9123 & n8240;
assign n1890 = n5625 & n9539;
assign n162 = n6954 | n1556;
assign n532 = n5874 & n9122;
assign n7860 = ~(n1610 ^ n6678);
assign n1027 = ~(n2802 ^ n11817);
assign n12004 = n8204 | n8128;
assign n4036 = n3130 & n1724;
assign n5604 = n12113 & n8008;
assign n6435 = ~(n6113 ^ n11235);
assign n5517 = n8935 | n12858;
assign n11403 = n8298 & n1821;
assign n8213 = ~(n4118 | n8321);
assign n1244 = n616 | n6117;
assign n2807 = n6519 | n8534;
assign n10747 = ~(n7856 ^ n9873);
assign n2231 = ~(n5181 | n11272);
assign n1230 = n10314 | n1043;
assign n9123 = ~(n2384 ^ n2873);
assign n8322 = ~n1252;
assign n3731 = n13182 | n5939;
assign n7765 = ~n9905;
assign n6346 = n3594 | n4632;
assign n12851 = n10756 | n10871;
assign n9417 = ~n4803;
assign n2038 = n317 & n1557;
assign n5958 = ~(n11039 | n521);
assign n2762 = n3634 | n8268;
assign n11292 = n1894 & n6191;
assign n6386 = ~(n12122 ^ n11788);
assign n6894 = n7255 | n5315;
assign n1189 = ~n7706;
assign n11547 = ~(n4740 ^ n11952);
assign n4645 = ~(n11050 ^ n5046);
assign n6260 = ~n7259;
assign n12346 = n13019 | n507;
assign n8454 = n472 | n1271;
assign n11761 = n8836 & n8766;
assign n10340 = n8488 | n8642;
assign n5422 = ~(n1768 ^ n6626);
assign n3400 = n9461 & n6269;
assign n4643 = ~n11158;
assign n2123 = ~n6273;
assign n6592 = n12999 & n4923;
assign n49 = ~(n7039 ^ n2105);
assign n10707 = ~(n1085 ^ n10860);
assign n11702 = n10281 | n1026;
assign n6549 = ~(n8373 ^ n5519);
assign n11321 = n56 & n4392;
assign n12117 = n11926 & n8657;
assign n3215 = n12019 | n6660;
assign n8714 = ~(n1239 ^ n4747);
assign n1815 = ~n4039;
assign n12057 = n8043 | n7270;
assign n9202 = n12348 & n6937;
assign n3685 = ~(n2530 ^ n9545);
assign n3561 = ~(n5052 | n11325);
assign n4524 = ~n9483;
assign n6888 = n9538 & n7942;
assign n12684 = n3467 & n5577;
assign n3135 = ~(n6222 ^ n6931);
assign n12200 = ~(n1478 | n6547);
assign n453 = n4252 | n9554;
assign n6262 = ~(n1611 ^ n8894);
assign n11491 = ~n3967;
assign n13175 = ~(n10993 ^ n8159);
assign n7757 = ~(n10703 ^ n1566);
assign n5363 = n8550 & n13119;
assign n8000 = ~(n2473 ^ n910);
assign n5174 = n11360 & n11330;
assign n1903 = n5645 | n7935;
assign n9722 = ~n3895;
assign n1267 = n4762 | n4375;
assign n2203 = n6506 | n8360;
assign n2809 = ~n2540;
assign n10570 = ~n3562;
assign n5203 = ~(n10424 | n13076);
assign n12216 = ~(n7832 ^ n9230);
assign n8293 = ~n11366;
assign n8455 = n9606 | n2544;
assign n9674 = ~n12468;
assign n582 = n7500 ^ n567;
assign n2745 = ~(n5987 ^ n6447);
assign n6481 = ~n7830;
assign n1270 = n3244 & n8457;
assign n6921 = n9353 & n3815;
assign n6432 = ~(n8237 ^ n3638);
assign n7149 = n3443 | n6795;
assign n1716 = ~(n5737 ^ n9262);
assign n7146 = ~n12651;
assign n5985 = ~(n5062 ^ n6957);
assign n12497 = ~(n3554 ^ n4108);
assign n10453 = ~(n7452 ^ n4151);
assign n7433 = n7311 | n6251;
assign n4429 = ~(n440 ^ n6827);
assign n9080 = ~n10451;
assign n7538 = n2764 | n7504;
assign n3691 = n3720 & n4079;
assign n8503 = ~(n12970 ^ n995);
assign n133 = n6777 | n10205;
assign n10197 = ~(n4928 ^ n3064);
assign n8875 = n1912 & n11634;
assign n7324 = n4236 & n11989;
assign n11107 = n917;
assign n7014 = ~(n12704 | n10267);
assign n11302 = ~(n10438 | n12849);
assign n8051 = n7329 | n12350;
assign n777 = n3910 ^ n9666;
assign n10108 = ~n3310;
assign n7389 = n4903 & n9015;
assign n10095 = ~(n12317 ^ n9902);
assign n9455 = n9087 & n2453;
assign n10762 = n6988 | n7430;
assign n526 = ~n3862;
assign n2645 = ~(n11520 ^ n7370);
assign n4552 = ~(n7494 | n2815);
assign n828 = n4198 | n7221;
assign n6505 = ~(n6884 | n6424);
assign n11367 = ~(n5125 ^ n12077);
assign n3521 = ~(n3351 ^ n1956);
assign n8291 = n3006 & n7411;
assign n4395 = n73 & n2634;
assign n377 = n5168 | n9159;
assign n9110 = ~(n6737 | n4245);
assign n905 = ~n2771;
assign n10116 = n8866 & n8620;
assign n4786 = ~n4020;
assign n3281 = ~n469;
assign n8304 = ~(n4728 | n10414);
assign n7475 = n6349 | n2408;
assign n9545 = n12473 ^ n11149;
assign n576 = ~(n8059 ^ n10722);
assign n4038 = n4144 | n8030;
assign n11356 = ~n1650;
assign n2692 = ~n7729;
assign n8845 = n1648 & n8952;
assign n2095 = ~n12605;
assign n99 = n9793 | n1144;
assign n9121 = ~(n1072 ^ n10473);
assign n4850 = n4830 | n12089;
assign n9945 = n938 ^ n7006;
assign n9507 = n5164 & n7412;
assign n5249 = n4523 | n10528;
assign n1043 = n3858;
assign n566 = n9479 & n8883;
assign n1310 = ~(n12466 ^ n10742);
assign n9470 = n11018 | n10213;
assign n1829 = n6687 & n432;
assign n4342 = ~n11901;
assign n12939 = n2449 | n1026;
assign n5088 = n10755 | n12831;
assign n9412 = ~(n1285 ^ n857);
assign n9167 = ~(n5858 ^ n7206);
assign n1301 = ~n2592;
assign n11426 = n3907 & n10413;
assign n4653 = ~n13160;
assign n10336 = n12663 | n10535;
assign n3034 = ~(n2120 ^ n3808);
assign n4846 = ~n8314;
assign n1634 = ~n5167;
assign n5908 = ~(n3891 ^ n2833);
assign n9175 = ~(n6603 ^ n10079);
assign n7448 = ~(n9441 ^ n8368);
assign n4880 = n7002 & n9240;
assign n7899 = n5025 | n3893;
assign n13162 = n7878 | n2893;
assign n13218 = n4232 | n6692;
assign n859 = ~(n3978 ^ n8270);
assign n10960 = n9487 | n4870;
assign n10859 = ~(n9318 ^ n10970);
assign n5355 = n3167 & n2995;
assign n8033 = ~n10789;
assign n8441 = ~(n7439 ^ n10963);
assign n8622 = n8863 | n10573;
assign n8617 = ~n9708;
assign n6774 = ~n1418;
assign n10783 = n9643 | n2775;
assign n4886 = ~(n4991 ^ n12980);
assign n11507 = ~(n3151 ^ n11033);
assign n13187 = ~(n6389 ^ n2869);
assign n68 = n10460 & n5589;
assign n1651 = ~n9300;
assign n5724 = n6346 & n1745;
assign n4345 = n3315 & n5760;
assign n4564 = ~n4862;
assign n4267 = n4156 | n10907;
assign n6292 = n10481 | n4514;
assign n6463 = ~n6058;
assign n10158 = ~n3145;
assign n9944 = ~(n1656 | n5376);
assign n226 = n1569 & n7883;
assign n5640 = ~(n4800 ^ n9103);
assign n12107 = ~n6456;
assign n3826 = ~n11891;
assign n4745 = n6890 & n6584;
assign n6933 = ~(n6864 | n4977);
assign n450 = ~(n4210 | n6150);
assign n2787 = ~(n1019 ^ n12245);
assign n1533 = n1041 | n3824;
assign n11594 = ~(n9918 ^ n11339);
assign n4095 = n4927 & n11100;
assign n6810 = ~n6149;
assign n10812 = n6223 | n10029;
assign n5674 = n9994 & n7811;
assign n6972 = ~(n8627 | n11334);
assign n1109 = n7486 & n6159;
assign n12411 = n8562 | n10106;
assign n3166 = n12759 | n356;
assign n3486 = n8625 | n9970;
assign n9472 = n6323 & n10510;
assign n4854 = n4089 & n9059;
assign n4284 = ~(n9096 ^ n1110);
assign n3921 = ~(n4630 ^ n4380);
assign n540 = ~(n10019 ^ n3472);
assign n9250 = ~(n11621 ^ n9175);
assign n9673 = n5806 | n2276;
assign n4593 = ~(n6701 | n7844);
assign n1179 = ~(n9612 ^ n12677);
assign n10662 = ~(n8888 ^ n9707);
assign n10264 = ~(n8023 ^ n12363);
assign n6369 = ~n6550;
assign n247 = ~(n4384 | n2210);
assign n9636 = n932 & n4494;
assign n571 = ~(n4709 ^ n7781);
assign n3052 = ~(n8087 ^ n3403);
assign n4015 = ~(n11010 ^ n9046);
assign n3859 = n12861 | n9661;
assign n2194 = n517 | n1229;
assign n9082 = ~(n695 ^ n6411);
assign n8922 = ~n10067;
assign n11765 = ~(n6599 | n1108);
assign n13 = n4077 | n8348;
assign n1356 = ~n2658;
assign n8790 = ~n4353;
assign n4661 = n12995 & n8433;
assign n2284 = n11113 | n4947;
assign n8638 = ~(n12329 ^ n12);
assign n7642 = ~n9093;
assign n11042 = ~(n3479 ^ n11084);
assign n1556 = ~(n7329 ^ n12350);
assign n10488 = n11333 | n3676;
assign n8850 = n2718 | n6769;
assign n402 = ~(n4196 | n2004);
assign n5496 = n6658 | n4373;
assign n2483 = ~(n12409 ^ n743);
assign n706 = ~(n3360 ^ n2234);
assign n12638 = ~(n11571 ^ n12271);
assign n4325 = n1216 & n8452;
assign n6514 = ~(n1177 ^ n9449);
assign n6416 = ~n4862;
assign n5856 = ~(n5194 ^ n5623);
assign n12469 = ~n9591;
assign n5313 = ~n1465;
assign n5930 = ~n9729;
assign n12626 = n9493 | n9114;
assign n9971 = ~(n6820 | n2915);
assign n458 = n3906 | n10250;
assign n666 = ~n2750;
assign n2589 = n5719 & n6057;
assign n5196 = n9102 & n10368;
assign n2721 = n8723 & n2151;
assign n9869 = n6387 | n7071;
assign n9435 = ~(n12178 ^ n5295);
assign n2197 = ~(n11971 | n9068);
assign n2540 = n542 | n206;
assign n9977 = n1419 | n30;
assign n12387 = n4937 & n978;
assign n11678 = ~(n12081 | n12116);
assign n11519 = ~n12284;
assign n9488 = n10792 | n5087;
assign n2982 = n3864 | n7218;
assign n4375 = ~(n7992 | n6554);
assign n4318 = ~(n2188 ^ n6955);
assign n6782 = ~(n4827 ^ n916);
assign n5257 = n10081 | n7282;
assign n2526 = ~(n3860 ^ n7352);
assign n4501 = ~(n7018 ^ n3328);
assign n8220 = n2088 & n5851;
assign n6839 = n2945 & n8559;
assign n10910 = ~n3824;
assign n5575 = n2559 & n4921;
assign n2499 = n1842 | n6697;
assign n1169 = n12868 & n2755;
assign n1315 = n12924 | n492;
assign n11858 = ~n5750;
assign n1793 = ~(n6558 ^ n9782);
assign n5319 = ~(n12184 ^ n2588);
assign n2524 = ~(n9358 | n4645);
assign n5885 = n5351 & n12659;
assign n11505 = n4861 & n5447;
assign n10625 = n10877 | n8702;
assign n6787 = n4834 & n12580;
assign n7375 = n4385 | n6769;
assign n1071 = ~(n4479 ^ n10582);
assign n2954 = ~(n1031 ^ n1412);
assign n8988 = ~(n8398 ^ n1190);
assign n9845 = ~(n11220 | n10953);
assign n5934 = ~(n351 ^ n4833);
assign n1680 = n1199 | n8030;
assign n11758 = ~(n3263 ^ n12045);
assign n5933 = n9181 | n4237;
assign n9207 = n3814 & n12504;
assign n11809 = ~(n7383 ^ n5068);
assign n10376 = n10908 & n469;
assign n8030 = n5654;
assign n7809 = n11340 | n4601;
assign n1470 = ~(n12947 ^ n43);
assign n13199 = ~(n2950 ^ n3143);
assign n2800 = ~n11068;
assign n4403 = n11291 | n12328;
assign n12105 = n7406 | n11860;
assign n1552 = ~(n7892 ^ n9818);
assign n7270 = ~(n13061 ^ n3066);
assign n6783 = ~n9822;
assign n10294 = n6330 & n3387;
assign n4674 = ~(n7096 | n8340);
assign n5861 = n1756 & n4773;
assign n10448 = ~n12289;
assign n5485 = ~n7540;
assign n11155 = n3616 | n12328;
assign n9973 = ~(n5606 ^ n13129);
assign n8722 = n12677 | n9612;
assign n3235 = ~n6302;
assign n8518 = n12112 ^ n11513;
assign n1059 = n11905 | n3782;
assign n10091 = n542 | n4936;
assign n11820 = ~(n11632 | n4683);
assign n7217 = n1038 ^ n8191;
assign n12599 = n7742 | n12188;
assign n11460 = n4722 | n9075;
assign n8194 = ~n6167;
assign n12229 = ~(n11221 ^ n1382);
assign n13211 = ~(n11691 ^ n11072);
assign n13152 = ~(n8298 | n1821);
assign n1284 = ~(n8049 ^ n5214);
assign n8624 = ~(n6027 ^ n4214);
assign n5165 = n6084 | n8061;
assign n114 = ~n10606;
assign n10951 = ~(n3765 ^ n10734);
assign n11693 = ~(n12715 ^ n3465);
assign n10177 = ~(n3319 ^ n3789);
assign n8229 = n11913 & n3642;
assign n8180 = n6375 | n11144;
assign n1534 = ~(n2894 ^ n806);
assign n239 = n2752 | n7010;
assign n2710 = n11779 | n9195;
assign n12281 = ~n424;
assign n11252 = ~(n3355 ^ n12364);
assign n10310 = n1446 & n11652;
assign n2508 = ~(n7940 | n2152);
assign n5202 = n4827 & n2240;
assign n2605 = ~n5237;
assign n4610 = ~n7659;
assign n2297 = n10418 & n3094;
assign n9859 = ~(n6012 | n8797);
assign n7747 = n2771 & n9531;
assign n7832 = n1390 & n12612;
assign n112 = n5976 & n1372;
assign n4746 = ~(n6495 ^ n2374);
assign n6066 = n9658 | n11809;
assign n9362 = n1605 | n6944;
assign n11373 = n12728 | n11209;
assign n2160 = n13036 | n5076;
assign n6203 = n2135 | n12881;
assign n1500 = ~(n11907 | n12327);
assign n5331 = n10021 | n7837;
assign n4226 = n11476 & n7398;
assign n9634 = n3487 & n4313;
assign n1812 = ~(n9946 ^ n12731);
assign n2991 = ~(n1063 ^ n5147);
assign n7057 = ~(n6259 ^ n3461);
assign n6530 = n12159 | n650;
assign n1929 = ~(n6024 ^ n9038);
assign n3874 = ~(n13009 | n7105);
assign n10950 = ~n9570;
assign n622 = ~n11618;
assign n6534 = ~(n3469 | n11958);
assign n4960 = ~n411;
assign n5478 = ~n12306;
assign n10285 = ~n2629;
assign n7495 = n8587 & n9776;
assign n2190 = ~(n3709 ^ n11769);
assign n7523 = n3225 | n8702;
assign n1318 = ~(n6107 ^ n444);
assign n4857 = n2332 | n4936;
assign n4384 = n4557 & n4703;
assign n7130 = ~n12935;
assign n4780 = ~n1902;
assign n11073 = ~(n414 ^ n945);
assign n1288 = n12799 & n5361;
assign n10224 = ~(n276 ^ n10454);
assign n1453 = n7752 | n10360;
assign n4776 = n12993 | n11274;
assign n8757 = ~n9300;
assign n2606 = ~(n12603 | n1910);
assign n12811 = ~(n645 | n3600);
assign n11198 = ~(n13153 | n4674);
assign n7176 = n10135 | n8030;
assign n6991 = ~(n10842 ^ n10347);
assign n1407 = ~(n2822 ^ n9658);
assign n7285 = ~(n8091 ^ n10382);
assign n697 = ~(n6766 ^ n4292);
assign n5664 = n12153 | n7825;
assign n1589 = ~n8290;
assign n5581 = n10516 & n4171;
assign n1611 = n2591 ^ n11202;
assign n1446 = n4964 & n8506;
assign n9108 = n2547 & n7471;
assign n317 = n8469 | n961;
assign n4563 = n2681 & n9344;
assign n1549 = ~n4946;
assign n6893 = n13214;
assign n8666 = ~n12282;
assign n12637 = n1536 | n6265;
assign n5953 = n8761 | n5769;
assign n102 = n12037 & n10467;
assign n8037 = n6452 & n7190;
assign n11028 = n8597 & n1578;
assign n4740 = n10193 | n5631;
assign n11713 = ~n641;
assign n313 = ~(n600 ^ n11224);
assign n10679 = ~(n2113 ^ n9024);
assign n2889 = ~n6085;
assign n11601 = ~(n2019 | n7696);
assign n5204 = n1099 | n9120;
assign n229 = ~(n5208 ^ n180);
assign n695 = n2723 | n12786;
assign n1884 = ~(n5284 ^ n818);
assign n6235 = n10128 | n12501;
assign n6003 = n10070 & n10053;
assign n664 = n3211 & n7814;
assign n4230 = n482;
assign n9864 = n8764 & n10880;
assign n4486 = n1697 & n12932;
assign n1685 = ~(n11636 ^ n5220);
assign n1674 = ~n11296;
assign n7101 = n11757 | n6265;
assign n5903 = ~(n2171 | n10665);
assign n8055 = ~n9136;
assign n3996 = n2283 | n3762;
assign n10633 = n7715 & n7411;
assign n11888 = n2660 | n6317;
assign n382 = ~(n1294 ^ n11480);
assign n10939 = n7133 | n12695;
assign n1548 = n10184 | n3391;
assign n11999 = n8594 | n12804;
assign n8837 = ~n10185;
assign n12839 = ~(n9514 ^ n9688);
assign n4236 = n6143 | n326;
assign n3773 = n12354 | n11414;
assign n6532 = n9909 ^ n3108;
assign n5057 = n437 | n87;
assign n7330 = ~(n2823 ^ n11962);
assign n10306 = ~(n5288 ^ n2274);
assign n9503 = ~(n3532 ^ n10935);
assign n676 = ~(n527 ^ n3992);
assign n3374 = n11050 & n457;
assign n2951 = n10497;
assign n7322 = n195 | n8198;
assign n600 = n6325 & n2006;
assign n10069 = ~(n11439 ^ n9667);
assign n10106 = n8640;
assign n5625 = n5328 | n10871;
assign n7090 = n10870 & n3937;
assign n2971 = n4732 | n7221;
assign n4496 = ~(n2613 ^ n2172);
assign n6001 = ~n6085;
assign n4982 = ~(n4130 ^ n1201);
assign n5299 = n2884 | n10016;
assign n8605 = ~(n9563 | n12216);
assign n7183 = ~(n12361 ^ n4526);
assign n3727 = ~n3061;
assign n8872 = ~(n2505 ^ n6340);
assign n12968 = ~(n3488 ^ n7965);
assign n11679 = n9392 & n8464;
assign n29 = ~(n5878 | n708);
assign n9899 = ~n10577;
assign n1029 = n2551 | n5501;
assign n13203 = n11972 & n11583;
assign n8646 = ~n22;
assign n4622 = ~(n3088 | n6184);
assign n11990 = n3634 | n8348;
assign n11337 = ~(n2066 ^ n12007);
assign n1635 = ~(n9607 | n1837);
assign n1218 = ~n10408;
assign n613 = n11657 | n7579;
assign n13141 = ~n3330;
assign n8810 = ~(n2897 ^ n4379);
assign n11580 = n2974 | n5240;
assign n3341 = n8760 | n540;
assign n959 = n9010 | n4947;
assign n7549 = ~n5266;
assign n12338 = ~(n5572 ^ n9762);
assign n1436 = ~n12289;
assign n1677 = n13079 | n6474;
assign n7341 = ~(n1378 ^ n9021);
assign n1942 = n6184 & n3088;
assign n375 = n4709 | n526;
assign n12527 = ~(n1389 ^ n11942);
assign n4782 = n11371 | n11292;
assign n1784 = n7932 | n12998;
assign n3175 = n11167 | n3485;
assign n4528 = ~(n6036 ^ n1641);
assign n12036 = ~n6522;
assign n6497 = ~(n473 | n1662);
assign n12007 = n11803 & n7886;
assign n9632 = ~n9591;
assign n3187 = n4523 ^ n11031;
assign n7652 = n8848 | n8227;
assign n5939 = ~n8230;
assign n567 = ~(n2246 ^ n3234);
assign n8471 = n3866 | n11668;
assign n2573 = n4224 | n9864;
assign n1246 = ~n5180;
assign n9144 = n10059 | n12388;
assign n1928 = ~(n12828 | n10732);
assign n3725 = n1135 | n12164;
assign n4527 = ~n7341;
assign n12083 = ~n13214;
assign n4222 = ~(n6555 | n8437);
assign n7783 = ~n2882;
assign n7076 = ~n411;
assign n10937 = n5681 & n5445;
assign n536 = n11810 | n12273;
assign n1387 = n6587 | n10179;
assign n6828 = ~(n1136 ^ n7956);
assign n11341 = ~n6790;
assign n4309 = ~(n6356 | n6989);
assign n10098 = ~n11441;
assign n2417 = ~(n1793 ^ n8178);
assign n12583 = ~(n3203 ^ n7054);
assign n4989 = ~(n5808 ^ n13209);
assign n12195 = n2866 & n12825;
assign n2716 = n10541 & n4260;
assign n12688 = ~(n6943 | n3637);
assign n10517 = n9946 & n9004;
assign n1020 = n147 | n10094;
assign n12751 = ~(n7567 ^ n6097);
assign n3631 = ~(n3298 ^ n1140);
assign n10237 = n1501 | n3971;
assign n5762 = ~(n10389 ^ n1964);
assign n6092 = ~(n11192 ^ n9199);
assign n4370 = ~n12408;
assign n9462 = ~(n12299 | n324);
assign n1172 = ~(n8581 ^ n10330);
assign n4298 = n4143 | n12501;
assign n5256 = n7622 | n8815;
assign n10602 = ~(n5290 ^ n5214);
assign n8733 = n12262 | n3227;
assign n1887 = ~n1307;
assign n4785 = n493 | n5169;
assign n725 = n6649 & n9770;
assign n6487 = ~(n4046 ^ n4603);
assign n8478 = ~(n5850 | n638);
assign n5154 = n5151 & n7843;
assign n2861 = ~n2498;
assign n12958 = ~(n1777 ^ n4029);
assign n10107 = ~(n11314 ^ n1037);
assign n10865 = n445 | n3949;
assign n2165 = ~n5678;
assign n4340 = ~(n8241 | n4807);
assign n10201 = n3110 | n1462;
assign n11318 = n6099 | n8268;
assign n6173 = ~n10606;
assign n12343 = n2965 | n12561;
assign n5891 = ~(n10839 ^ n3559);
assign n7735 = n5142 & n4945;
assign n7005 = ~(n1414 | n8960);
assign n7260 = n3893 & n5025;
assign n6734 = n5568 & n3006;
assign n12080 = n10500 | n11063;
assign n11840 = n5568 & n4470;
assign n10048 = ~(n9994 ^ n9963);
assign n7956 = ~(n6870 ^ n9144);
assign n1851 = ~(n12661 ^ n1196);
assign n9801 = n8648 | n6436;
assign n5721 = ~n2010;
assign n980 = ~n4377;
assign n5235 = n2960 & n3240;
assign n981 = n9054 & n11825;
assign n7267 = ~(n9957 ^ n11036);
assign n10808 = n1364 & n9915;
assign n4790 = n6682 | n7324;
assign n8998 = n5460 | n6306;
assign n2904 = ~(n2668 ^ n5429);
assign n8166 = ~n9611;
assign n10972 = n11345 | n5250;
assign n11741 = n9216 & n5962;
assign n9464 = ~n2279;
assign n1693 = n4185 | n13181;
assign n11646 = n12151 | n1814;
assign n4900 = ~(n2536 ^ n4821);
assign n7168 = ~(n7286 ^ n12377);
assign n10715 = ~n4877;
assign n1931 = n1159 | n6429;
assign n2908 = n8720 | n11300;
assign n5230 = ~(n770 ^ n7115);
assign n10907 = ~(n8273 | n12986);
assign n57 = n12042 | n1836;
assign n680 = ~(n11739 ^ n4324);
assign n7965 = n5835 ^ n11492;
assign n8438 = ~n6669;
assign n6858 = n686 | n11679;
assign n11862 = n2771 & n12289;
assign n6072 = ~(n6744 | n347);
assign n6962 = n12882 | n4373;
assign n11103 = ~(n1626 ^ n11694);
assign n5820 = n9835 | n1378;
assign n6074 = n9061 | n8364;
assign n2064 = ~(n6510 | n5160);
assign n3743 = n4102 | n5002;
assign n1598 = n8139 & n9475;
assign n1106 = ~(n1545 ^ n10438);
assign n6892 = ~(n9494 ^ n11976);
assign n7436 = ~n11565;
assign n12711 = n10775 & n9956;
assign n10068 = ~n1242;
assign n4463 = n2712 & n5640;
assign n2912 = n2669 | n8268;
assign n1365 = n899 | n12501;
assign n2360 = ~(n5958 | n5426);
assign n9642 = n3537 | n12388;
assign n5981 = n3892 | n6404;
assign n8199 = ~n8571;
assign n3339 = n5749 | n2133;
assign n1799 = n4659 | n3151;
assign n7083 = ~(n7552 ^ n13020);
assign n1116 = n6160 & n10010;
assign n10963 = n208 & n9716;
assign n11441 = n5077 & n12702;
assign n4084 = n7772 & n12289;
assign n9581 = ~n9591;
assign n13116 = ~n11971;
assign n12866 = n4799 & n9074;
assign n10461 = n8973 & n2132;
assign n4512 = ~(n7932 ^ n6677);
assign n11857 = n3191 & n3423;
assign n3373 = ~n2464;
assign n6448 = ~n5421;
assign n4710 = n7890 | n2919;
assign n9721 = n7379 | n9116;
assign n5338 = n820 | n4832;
assign n8380 = n4686 | n4796;
assign n3660 = n3784 | n3981;
assign n6898 = n2655 & n12479;
assign n13106 = n117 & n1749;
assign n12266 = n5875 | n12721;
assign n11139 = n8903 | n5432;
assign n7201 = ~(n4184 ^ n11855);
assign n5999 = ~n11061;
assign n6967 = ~n5969;
assign n12462 = n11864 | n12328;
assign n10438 = n4258 | n12501;
assign n4904 = n5070 & n5438;
assign n7430 = ~n10408;
assign n4652 = n10610 & n12525;
assign n0 = ~n7720;
assign n1906 = n12913 | n11351;
assign n8242 = ~(n7821 ^ n4767);
assign n5924 = n5291 & n3288;
assign n2291 = n11605 | n7288;
assign n11093 = ~(n2314 | n1042);
assign n9709 = ~n11236;
assign n1722 = n5352 ^ n7044;
assign n11181 = ~(n856 ^ n2560);
assign n3895 = ~n11974;
assign n5566 = n12354 & n11414;
assign n9046 = ~(n9146 ^ n11802);
assign n1927 = n5709 ^ n10343;
assign n12298 = n8334 & n11717;
assign n8957 = n5226 | n177;
assign n10405 = ~(n10655 ^ n224);
assign n3517 = n4462 | n6265;
assign n8160 = ~n12592;
assign n6332 = ~n2882;
assign n1913 = ~(n11273 ^ n3957);
assign n1574 = n3683 | n9832;
assign n10965 = n3826 | n4194;
assign n2032 = n179 & n9740;
assign n4768 = ~(n4545 | n1834);
assign n10924 = ~n11546;
assign n7059 = ~(n7604 ^ n531);
assign n744 = n7059 ^ n8997;
assign n4071 = ~(n12599 ^ n10350);
assign n7133 = ~n2666;
assign n9770 = n4874 | n9419;
assign n5916 = n9765 | n7491;
assign n9066 = n7872 | n9075;
assign n6998 = n8556 | n1144;
assign n8411 = ~(n12405 ^ n4951);
assign n12052 = ~n8860;
assign n2192 = n12677 & n9612;
assign n10014 = ~n3100;
assign n6341 = n11075 | n13210;
assign n7325 = n3430 | n7557;
assign n9037 = ~(n10980 ^ n3181);
assign n847 = ~(n4145 ^ n12150);
assign n7702 = n1571 | n5841;
assign n8500 = ~n7065;
assign n8705 = ~(n6334 ^ n9719);
assign n12551 = n8407 & n12321;
assign n6132 = n3160 & n10435;
assign n753 = ~(n11138 ^ n10801);
assign n6751 = ~n9531;
assign n5260 = ~(n4265 ^ n2715);
assign n12630 = n4290 | n9195;
assign n10550 = ~(n3384 | n4670);
assign n9544 = ~(n6904 ^ n1875);
assign n1398 = ~(n12669 ^ n8230);
assign n11984 = ~(n10518 ^ n7943);
assign n5569 = ~n3112;
assign n1761 = n3243 | n8702;
assign n4654 = n2452 | n12501;
assign n12021 = ~(n6327 ^ n10499);
assign n4211 = ~(n11666 ^ n2626);
assign n7645 = n9632 | n11354;
assign n10659 = n8073 & n5247;
assign n1083 = ~(n9713 ^ n12136);
assign n7582 = n9455 | n8253;
assign n10153 = ~(n2661 ^ n8195);
assign n6993 = ~(n5114 | n10306);
assign n10860 = n245 & n9099;
assign n3575 = ~(n7516 ^ n10779);
assign n5841 = ~n1364;
assign n12755 = ~(n7822 | n9603);
assign n10841 = n614 & n133;
assign n10719 = n6344 | n2234;
assign n8159 = n3217 | n10246;
assign n7456 = n8264 | n10834;
assign n5552 = ~(n12639 ^ n7698);
assign n11899 = ~(n10638 ^ n606);
assign n7833 = ~n3091;
assign n537 = ~(n8319 ^ n711);
assign n3757 = ~(n11276 ^ n4801);
assign n1655 = n9020 & n5771;
assign n10870 = n11021 | n6999;
assign n7623 = n11519 | n9282;
assign n3209 = ~(n5397 ^ n10933);
assign n5059 = n2373 & n782;
assign n12634 = ~(n2143 ^ n8527);
assign n2869 = ~(n4338 ^ n5618);
assign n7116 = ~(n10825 ^ n2052);
assign n7884 = n11397 & n12558;
assign n13005 = ~n2068;
assign n6924 = ~n4002;
assign n8237 = n10926 | n6564;
assign n10327 = n6220 | n4144;
assign n8978 = n3491 | n4672;
assign n7640 = n1817 & n5904;
assign n8382 = ~(n10269 ^ n5570);
assign n6807 = n2219 | n7052;
assign n8219 = ~(n7572 ^ n6450);
assign n5703 = n10713 | n2994;
assign n9323 = ~n5709;
assign n6588 = n6562 | n2201;
assign n6077 = ~(n12332 ^ n4771);
assign n8707 = n51 & n671;
assign n872 = n621 ^ n9836;
assign n6367 = ~n1724;
assign n9998 = n11821 & n8132;
assign n5813 = ~(n9186 ^ n4081);
assign n553 = ~(n10034 | n5089);
assign n3766 = ~n6660;
assign n9345 = ~n6174;
assign n12982 = n12074 & n1873;
assign n8254 = ~n9669;
assign n4604 = ~n10225;
assign n11973 = ~n8967;
assign n6745 = n12321 | n8407;
assign n5733 = ~n5065;
assign n12164 = ~n854;
assign n11008 = ~n3134;
assign n3359 = n5316 | n9290;
assign n12835 = ~(n6441 ^ n6671);
assign n3780 = n3962 | n8490;
assign n11312 = n9739 | n11101;
assign n8784 = n7690 | n199;
assign n7829 = n8166 & n5434;
assign n2378 = n6463 | n2976;
assign n10588 = n5816 & n136;
assign n1855 = n1111 | n4207;
assign n6190 = n9166 & n4284;
assign n11138 = ~(n6088 ^ n5610);
assign n10312 = ~(n6801 ^ n4476);
assign n3322 = ~(n1527 | n6961);
assign n2628 = n2778 & n12433;
assign n10280 = ~(n9296 | n11838);
assign n6687 = n8658 | n6891;
assign n7619 = n8998 & n12132;
assign n4026 = n1623 & n5001;
assign n7472 = n12106 & n7929;
assign n6128 = n199 & n7690;
assign n1702 = ~(n12936 | n12538);
assign n7248 = ~(n3152 ^ n6017);
assign n10811 = ~(n7220 ^ n12373);
assign n13006 = n11320 | n5076;
assign n4310 = ~(n9656 ^ n1948);
assign n4055 = ~n5332;
assign n9171 = ~(n1611 | n8834);
assign n10573 = ~n11030;
assign n9678 = ~(n1227 ^ n4647);
assign n4723 = ~n4064;
assign n5812 = ~n2977;
assign n10643 = ~(n3398 ^ n9480);
assign n3047 = ~n510;
assign n1101 = ~n2758;
assign n8189 = n1597 & n10618;
assign n3577 = n5070 | n5438;
assign n6744 = n10974 | n8268;
assign n8451 = ~(n3140 ^ n5398);
assign n275 = ~n10963;
assign n11934 = ~(n12580 ^ n4669);
assign n12114 = ~n92;
assign n12973 = ~(n8890 ^ n5955);
assign n12919 = n7297 & n303;
assign n7143 = n8329 | n12847;
assign n11767 = ~(n1873 ^ n3497);
assign n7742 = ~n2252;
assign n1025 = n1945 & n8601;
assign n7064 = n9238 | n2059;
assign n12437 = ~(n12815 | n2874);
assign n12503 = ~(n8218 ^ n3059);
assign n9629 = n12680 & n6636;
assign n839 = n8245 | n12039;
assign n820 = n6381 | n10886;
assign n11768 = n5863 & n5436;
assign n4289 = n10177 | n8075;
assign n6054 = ~(n5214 | n2771);
assign n3350 = n3313 | n14;
assign n2566 = n13177 & n3705;
assign n5860 = n7839 & n3552;
assign n6654 = n11352 | n2544;
assign n6418 = n9974 & n9323;
assign n1831 = n5462 & n11716;
assign n2774 = n5970 & n1687;
assign n5627 = ~(n8856 | n4340);
assign n9942 = ~n7209;
assign n6551 = ~(n6018 ^ n280);
assign n2153 = n359 | n7905;
assign n11774 = n8466 & n11222;
assign n20 = ~(n37 | n5224);
assign n12807 = n9646 | n12984;
assign n3885 = ~n8043;
assign n12607 = ~(n2233 | n1421);
assign n4307 = ~(n2368 ^ n10107);
assign n12090 = n121 | n11609;
assign n138 = ~n1912;
assign n11308 = ~n7517;
assign n4651 = n3340 & n1953;
assign n11063 = n12841 | n9075;
assign n8198 = ~(n9336 | n4152);
assign n4447 = n1251 & n3351;
assign n1922 = n1039 & n10655;
assign n6009 = ~(n5726 ^ n1552);
assign n10781 = ~n497;
assign n3905 = ~(n12901 ^ n8047);
assign n1991 = ~(n9443 ^ n4261);
assign n10473 = n2999 & n10235;
assign n2730 = ~(n11805 ^ n1969);
assign n9190 = ~(n7 ^ n10231);
assign n11640 = n4808 | n12847;
assign n6244 = ~n4646;
assign n9382 = ~n6034;
assign n1578 = n6383 | n10179;
assign n7750 = n4863 | n243;
assign n11296 = ~(n8557 ^ n3704);
assign n8939 = ~(n13156 ^ n11186);
assign n4434 = ~(n4408 ^ n5910);
assign n2881 = ~(n12760 ^ n5012);
assign n8298 = n8681 | n4373;
assign n6033 = ~n3815;
assign n3317 = ~(n4216 ^ n6668);
assign n6417 = n10049 | n9223;
assign n6528 = ~n11394;
assign n1331 = ~n3409;
assign n6040 = ~n3085;
assign n2974 = ~(n9317 ^ n2458);
assign n7732 = n4352 | n9682;
assign n10510 = n7731 | n4596;
assign n7713 = ~(n3512 ^ n6781);
assign n7990 = n4046 | n11638;
assign n3902 = ~(n6357 | n2325);
assign n6679 = ~(n10832 | n13007);
assign n5751 = ~(n5847 ^ n2915);
assign n5779 = n435 & n4776;
assign n442 = ~n6453;
assign n8246 = ~(n2640 | n1858);
assign n1197 = ~n854;
assign n10848 = n7908 | n5302;
assign n10619 = n9649 & n2096;
assign n5317 = n10157 & n400;
assign n1588 = n6368 | n1154;
assign n12517 = n2574 | n11228;
assign n4407 = n11945 & n3773;
assign n6544 = n12196 & n2269;
assign n12461 = ~(n10548 ^ n6281);
assign n1934 = n11119 & n9900;
assign n7868 = ~n4335;
assign n5224 = n8006 | n12242;
assign n5008 = n8379 & n5273;
assign n3096 = ~n4419;
assign n9391 = ~(n10308 | n12917);
assign n3950 = ~(n4439 ^ n10177);
assign n3573 = ~(n2924 ^ n771);
assign n9648 = n11868 | n8030;
assign n3292 = ~(n1911 ^ n9862);
assign n3189 = ~(n5833 | n3095);
assign n13124 = ~(n5648 ^ n7420);
assign n7036 = ~(n10895 ^ n4183);
assign n8386 = n5990 | n7723;
assign n6211 = n8176 | n2221;
assign n1257 = n12533 | n283;
assign n10125 = ~(n6727 ^ n5083);
assign n12681 = n2221 | n7723;
assign n2492 = n3068 | n7530;
assign n12363 = ~(n8488 ^ n8642);
assign n9849 = n11376 ^ n10200;
assign n3852 = n10686 | n1895;
assign n3223 = ~(n12588 ^ n9302);
assign n1279 = ~(n574 | n9405);
assign n2702 = n10936 | n10028;
assign n3158 = ~n12482;
assign n1925 = n8811 & n7284;
assign n5743 = n2444 & n11461;
assign n1708 = ~(n3707 ^ n1371);
assign n8470 = ~n5535;
assign n9907 = n2046 & n12637;
assign n11314 = ~(n2801 ^ n7993);
assign n7180 = n4616 & n8255;
assign n9706 = ~n11076;
assign n5755 = ~(n12477 ^ n9404);
assign n10290 = ~n1650;
assign n3270 = n7062 | n7221;
assign n9820 = ~(n11120 ^ n12459);
assign n7597 = ~n3815;
assign n13129 = ~(n4887 ^ n10523);
assign n4821 = n3509 | n7723;
assign n7690 = n5265 | n4640;
assign n5412 = n8023 | n11569;
assign n3649 = n6916 & n1664;
assign n5580 = ~(n3597 ^ n12050);
assign n6406 = ~(n9133 ^ n5113);
assign n11438 = n4301 & n344;
assign n1872 = ~(n8291 | n783);
assign n11538 = n5367 & n8496;
assign n11518 = n1308 & n4498;
assign n6650 = ~(n1501 ^ n6256);
assign n9813 = n7284 | n8811;
assign n8793 = n7176 & n8366;
assign n5509 = ~(n5637 ^ n8193);
assign n7214 = n2670 ^ n12665;
assign n3151 = n1571 | n1570;
assign n10398 = n10770 & n510;
assign n9064 = ~(n2141 | n10841);
assign n3807 = n9810 | n3805;
assign n6383 = ~n12263;
assign n12355 = n12093 | n12273;
assign n6596 = ~n10522;
assign n12675 = n1130 & n12088;
assign n10774 = n2880 & n11154;
assign n8210 = ~n12414;
assign n5430 = ~n13058;
assign n7799 = ~(n11134 ^ n10687);
assign n3128 = ~n4982;
assign n3533 = n3407 | n177;
assign n4424 = ~(n395 ^ n9659);
assign n2474 = n12441 | n9223;
assign n4913 = ~(n9938 | n3146);
assign n11336 = n3385 | n2005;
assign n11952 = ~(n8137 ^ n10954);
assign n7952 = ~(n7160 | n4374);
assign n8550 = n5688 | n5076;
assign n2012 = ~(n11117 ^ n3093);
assign n8489 = ~(n7048 | n11265);
assign n860 = n11069 & n4158;
assign n10499 = n7281;
assign n597 = n11555 & n9728;
assign n1788 = ~(n8448 ^ n12496);
assign n10726 = ~n5871;
assign n2222 = ~n11030;
assign n7177 = ~(n4041 ^ n7392);
assign n2557 = ~n9353;
assign n5530 = ~(n2460 ^ n10987);
assign n10181 = ~(n5980 ^ n4238);
assign n8132 = n12172 | n10472;
assign n9401 = n6906 & n6186;
assign n3569 = ~(n12582 ^ n1204);
assign n12104 = n2790 | n4546;
assign n12645 = ~(n12276 ^ n1094);
assign n10188 = ~n8468;
assign n3092 = ~n3087;
assign n877 = n6590 | n5076;
assign n8712 = n4406 & n5165;
assign n7211 = n6629 | n11107;
assign n3263 = n2321 | n7998;
assign n2543 = ~(n6111 ^ n8211);
assign n9471 = n9154 | n4640;
assign n12906 = ~n11551;
assign n10834 = n8849 | n6635;
assign n5610 = n6367 | n11521;
assign n3356 = ~(n2343 | n3861);
assign n4794 = ~(n4321 ^ n11749);
assign n8989 = ~n5553;
assign n491 = n410 & n8662;
assign n1923 = n110 & n5946;
assign n7707 = ~n6826;
assign n12819 = n4114 & n2339;
assign n169 = n5007 | n6977;
assign n7352 = n623 & n2863;
assign n5720 = n12563 | n4640;
assign n5215 = ~n4146;
assign n12404 = n8277 & n2337;
assign n9506 = n6318 & n12057;
assign n7635 = ~(n10053 | n10070);
assign n3568 = ~(n1560 ^ n1654);
assign n8846 = n4114 & n1916;
assign n6188 = n8380 | n11981;
assign n5246 = n12697 | n7640;
assign n3205 = ~(n13206 | n5473);
assign n6100 = ~n1964;
assign n1629 = ~n7552;
assign n6237 = n10327 & n6711;
assign n271 = n2352 | n4352;
assign n10896 = n7917 | n2049;
assign n8570 = n5939 | n9159;
assign n4422 = n10710 & n7665;
assign n10283 = ~(n6373 ^ n3663);
assign n7840 = ~(n10139 ^ n1093);
assign n3914 = n11277 | n71;
assign n2189 = n6365 | n8560;
assign n7632 = n5826 | n2831;
assign n5240 = n10526 & n9892;
assign n7067 = ~(n675 ^ n12345);
assign n10905 = ~(n5978 | n8126);
assign n5087 = ~n3085;
assign n6081 = ~(n7010 ^ n9663);
assign n12671 = ~n6937;
assign n2275 = ~(n8880 ^ n7789);
assign n12542 = n8700 & n8382;
assign n936 = n12330 | n2731;
assign n4879 = ~n3121;
assign n6837 = n5182 | n3981;
assign n2902 = ~n679;
assign n12095 = ~n12101;
assign n3371 = n5752 | n2177;
assign n3741 = ~(n307 ^ n2033);
assign n5089 = n4369 & n2951;
assign n364 = ~n6730;
assign n11436 = ~(n11248 | n8200);
assign n11231 = ~n8788;
assign n794 = n5683 | n3949;
assign n2279 = n6236 & n11565;
assign n2840 = ~(n3348 ^ n1167);
assign n3 = n8154 & n8975;
assign n12642 = n1358 & n1766;
assign n4760 = n4875 | n7935;
assign n7145 = ~(n5479 ^ n2648);
assign n8896 = n6768 | n4442;
assign n2423 = ~(n7395 ^ n2131);
assign n3258 = ~(n7267 ^ n11413);
assign n10549 = n5692 & n5834;
assign n9422 = n8242 & n1491;
assign n7220 = n7636 & n4562;
assign n1069 = ~(n307 | n3422);
assign n12251 = ~(n7465 ^ n12357);
assign n8164 = n2066 | n12007;
assign n6672 = ~n772;
assign n417 = n7394 | n5379;
assign n2063 = ~(n1740 | n9881);
assign n3121 = ~n4426;
assign n9936 = ~(n6302 ^ n9032);
assign n5749 = ~n5536;
assign n9672 = n9513 | n1400;
assign n11688 = n13183 | n1570;
assign n4616 = n4537 & n10408;
assign n9510 = n6668 & n4470;
assign n1421 = n13178 & n6576;
assign n829 = ~n6818;
assign n8571 = n3962 | n7935;
assign n9519 = n4741 | n12328;
assign n11627 = ~(n7746 ^ n3856);
assign n13135 = n3280 & n3844;
assign n8555 = ~(n143 ^ n7237);
assign n12795 = ~n10805;
assign n2211 = ~n6362;
assign n8145 = n7568 & n6376;
assign n9760 = n8187 & n3620;
assign n3011 = ~(n1960 ^ n8939);
assign n7524 = n4664 & n2728;
assign n4090 = ~(n3250 ^ n12226);
assign n1712 = ~n1752;
assign n6857 = ~(n7660 ^ n8709);
assign n2685 = n8421 & n5150;
assign n1988 = ~(n7137 ^ n8096);
assign n9776 = ~(n7809 ^ n13232);
assign n9966 = n3433 | n3649;
assign n10692 = ~n472;
assign n9521 = ~(n11448 | n3082);
assign n1233 = ~(n2600 ^ n5000);
assign n12610 = n10792 | n2449;
assign n1394 = n7223 | n9223;
assign n9112 = ~n5065;
assign n4767 = ~(n5039 ^ n1678);
assign n19 = ~n11151;
assign n598 = n896 & n11620;
assign n10807 = n12814 | n5242;
assign n6952 = n2199 & n2385;
assign n6319 = ~(n6972 | n12694);
assign n2945 = ~n1623;
assign n10126 = ~(n9134 ^ n2035);
assign n5042 = ~(n7489 ^ n10836);
assign n9925 = ~(n220 ^ n2548);
assign n10736 = ~(n7885 ^ n1010);
assign n201 = ~(n8304 ^ n7347);
assign n9917 = ~n4743;
assign n5780 = ~(n11318 ^ n2275);
assign n10596 = ~(n3590 ^ n9256);
assign n898 = n12126 | n1144;
assign n8526 = n11994 | n331;
assign n989 = ~(n2521 | n6792);
assign n12242 = ~n1364;
assign n7333 = n6677 | n12714;
assign n11458 = ~(n4428 ^ n3446);
assign n552 = n11500 & n710;
assign n6986 = ~n4862;
assign n98 = ~n11634;
assign n11525 = ~n9540;
assign n10378 = ~(n6805 ^ n5386);
assign n12049 = ~n834;
assign n4877 = ~n12083;
assign n4285 = n10914 ^ n5960;
assign n4944 = ~(n11546 | n7199);
assign n10788 = ~(n7382 | n10461);
assign n8679 = ~n1915;
assign n412 = n10291 & n11439;
assign n6957 = n7069 ^ n5124;
assign n10320 = n2452 | n11522;
assign n3421 = ~(n348 | n4219);
assign n7002 = ~(n3090 ^ n13095);
assign n5838 = ~n1935;
assign n2422 = ~(n1510 ^ n11298);
assign n655 = n3736 & n929;
assign n10233 = n7789 | n4492;
assign n1103 = n12353 & n8316;
assign n9791 = n8648 & n6436;
assign n609 = n3067 | n10985;
assign n4970 = n7242 | n12886;
assign n12549 = ~(n3030 ^ n9878);
assign n10262 = n10112 | n5521;
assign n7916 = n9675 | n1570;
assign n10649 = ~(n2784 ^ n1838);
assign n8190 = ~(n4244 ^ n6547);
assign n5092 = n10277 & n3297;
assign n6249 = ~(n7732 ^ n6035);
assign n7926 = ~(n11447 ^ n12277);
assign n8053 = ~n353;
assign n10714 = ~n8468;
assign n6815 = n5502 ^ n11319;
assign n5772 = n7260 | n523;
assign n8964 = ~(n8654 | n8951);
assign n7716 = ~n11016;
assign n9633 = ~(n6598 ^ n12439);
assign n4547 = n565 | n8593;
assign n2801 = n3364 | n6033;
assign n8011 = ~n8135;
assign n2270 = n3880 | n8953;
assign n13074 = n13021 & n6232;
assign n9410 = ~(n10487 ^ n3904);
assign n6626 = n8415 | n11959;
assign n6049 = n399 & n2596;
assign n643 = ~(n12806 ^ n2589);
assign n5961 = ~(n7043 ^ n8136);
assign n3926 = n2302 & n844;
assign n13167 = ~n13217;
assign n9308 = ~n2466;
assign n2301 = n11683 | n3981;
assign n4085 = n1659 | n10574;
assign n7385 = ~(n12315 | n6495);
assign n12481 = ~(n4592 ^ n5889);
assign n2896 = ~(n11455 ^ n11839);
assign n9178 = n3833 & n2946;
assign n1834 = ~(n10020 | n12884);
assign n7396 = ~n3769;
assign n4968 = ~(n7155 ^ n9825);
assign n3881 = ~(n9670 ^ n7902);
assign n6357 = ~(n12358 ^ n9412);
assign n5593 = n3006 & n12289;
assign n11539 = n2485 | n6032;
assign n8060 = n7291 | n8030;
assign n7444 = n9161 | n6372;
assign n11118 = ~(n6569 | n7169);
assign n10826 = ~(n4298 ^ n8262);
assign n4451 = n2825 | n12388;
assign n754 = n3606 ^ n12632;
assign n232 = ~(n10284 ^ n12513);
assign n11217 = n1731 ^ n4443;
assign n1325 = ~n11061;
assign n11461 = n10017 | n8490;
assign n1037 = ~(n4351 ^ n3482);
assign n2858 = ~n11937;
assign n5876 = ~(n6765 ^ n2572);
assign n10259 = ~(n5637 | n8193);
assign n9534 = ~(n8762 ^ n1397);
assign n8299 = ~(n11211 ^ n5422);
assign n383 = n7074 | n9223;
assign n5919 = ~(n11953 | n578);
assign n3961 = n207 & n12290;
assign n3535 = ~(n12996 ^ n6514);
assign n7904 = ~(n8643 | n7954);
assign n7218 = ~(n2112 | n5614);
assign n75 = ~n13060;
assign n7705 = ~(n4397 | n8165);
assign n12072 = n10500 & n11063;
assign n1664 = n1578 | n8597;
assign n5239 = ~(n12191 | n12700);
assign n12523 = ~(n8714 ^ n7677);
assign n2254 = ~n8860;
assign n7786 = ~(n5120 | n8474);
assign n11455 = n10037 | n8534;
assign n7428 = ~(n4931 ^ n9577);
assign n6869 = ~(n7362 | n12609);
assign n460 = ~(n4273 ^ n7985);
assign n1261 = ~n2882;
assign n12803 = ~(n4275 ^ n76);
assign n8202 = n3101 | n1789;
assign n10047 = ~(n9108 ^ n7036);
assign n10856 = ~n4586;
assign n9751 = n3911 | n4947;
assign n3297 = n3517 | n3571;
assign n10169 = ~(n4314 ^ n5004);
assign n6639 = n6275 & n9993;
assign n10863 = ~(n12137 ^ n3213);
assign n4136 = ~n7307;
assign n7725 = ~(n10025 ^ n12079);
assign n13238 = ~n10770;
assign n6255 = ~n8218;
assign n7122 = n5261 | n3981;
assign n9430 = ~n5815;
assign n12565 = n7435 & n12294;
assign n4909 = ~(n10864 ^ n1757);
assign n9298 = n4352 | n4947;
assign n12722 = n2150 | n3177;
assign n5658 = ~n6791;
assign n6175 = ~n6780;
assign n12450 = n3469 & n11958;
assign n7662 = n9920 | n8423;
assign n12136 = n543 | n6982;
assign n5415 = n8549 & n8919;
assign n12123 = ~(n6832 ^ n13124);
assign n4599 = n2080 | n2463;
assign n1122 = ~(n8518 ^ n6081);
assign n10102 = n7980 & n3846;
assign n3386 = ~(n5403 | n11387);
assign n5513 = n13089 | n6207;
assign n3742 = ~(n884 ^ n11251);
assign n10234 = ~n10409;
assign n6727 = n3830 & n4098;
assign n6472 = n3018 | n6951;
assign n3253 = ~n6222;
assign n1202 = n7358 | n6769;
assign n10936 = n87 & n437;
assign n3755 = ~n6643;
assign n7789 = n6028 | n7221;
assign n7882 = ~(n11501 ^ n8611);
assign n8366 = n11466 | n4640;
assign n12683 = n11511 & n9621;
assign n12451 = ~(n2333 ^ n11830);
assign n12643 = n2382 | n3546;
assign n2639 = ~n5189;
assign n11686 = ~(n3931 | n5119);
assign n11166 = n1735 & n10674;
assign n1300 = ~n1075;
assign n7391 = n5452 | n12681;
assign n10818 = n34 & n701;
assign n6733 = ~n5189;
assign n6271 = ~n9591;
assign n1456 = ~(n6454 ^ n2895);
assign n5127 = ~(n4027 ^ n10952);
assign n1047 = ~n3605;
assign n7225 = n6433 & n6276;
assign n1184 = ~n7387;
assign n1040 = n8838 | n6078;
assign n1565 = ~(n12801 | n9604);
assign n113 = ~(n5734 ^ n6886);
assign n7255 = n1653 & n6479;
assign n4182 = ~(n8245 ^ n3632);
assign n3228 = ~(n11268 ^ n298);
assign n2184 = ~(n4599 ^ n9361);
assign n4531 = n7188 | n8534;
assign n9415 = n1105 & n3136;
assign n4293 = ~n12391;
assign n11358 = ~(n10261 ^ n8820);
assign n6675 = n6725 & n10862;
assign n9767 = ~n9093;
assign n9051 = n8200 | n2216;
assign n3361 = n13077 | n3454;
assign n2632 = ~(n7731 ^ n4596);
assign n5783 = n882 | n8655;
assign n3335 = n11061 & n3769;
assign n11344 = ~n3398;
assign n288 = ~(n4941 | n12229);
assign n736 = ~(n274 ^ n7318);
assign n4873 = n3060 & n7046;
assign n1501 = n3047 | n11354;
assign n12521 = n1933 | n9407;
assign n1540 = ~n5897;
assign n642 = ~(n11904 ^ n6788);
assign n2193 = n1725 | n6769;
assign n6495 = ~(n10036 ^ n3072);
assign n4715 = ~n11837;
assign n2786 = n6178 | n5048;
assign n11099 = ~n8476;
assign n2860 = n11618 | n4136;
assign n4493 = n6336 | n8752;
assign n4611 = n10287 | n12695;
assign n974 = n1786 & n254;
assign n4373 = n12537;
assign n10081 = n10229 | n6288;
assign n9377 = ~(n3227 ^ n12262);
assign n4129 = n6168 & n5729;
assign n8749 = n2768 | n8268;
assign n6303 = n8301 | n6166;
assign n7088 = ~(n12294 ^ n5067);
assign n9557 = ~n1724;
assign n10037 = ~n8233;
assign n10136 = n12841 | n121;
assign n874 = ~(n8703 ^ n4965);
assign n7278 = n7775 | n11483;
assign n6632 = n203 & n4218;
assign n3595 = n1326 | n5476;
assign n1768 = ~(n4555 | n2450);
assign n11798 = n5533 & n5621;
assign n2253 = n475 | n12942;
assign n6492 = n6439 | n6306;
assign n7479 = n12445 & n1681;
assign n8824 = n3852 & n10363;
assign n9454 = n3360 | n10511;
assign n11522 = ~n8230;
assign n4992 = ~(n8211 | n6111);
assign n5342 = n5947 | n7723;
assign n12509 = ~(n6540 ^ n10603);
assign n2765 = ~(n5937 ^ n643);
assign n2429 = ~(n5283 | n2554);
assign n8303 = ~(n13027 ^ n3653);
assign n5444 = ~(n9886 ^ n2218);
assign n7165 = ~(n6718 ^ n2847);
assign n10083 = n4753 & n8570;
assign n4811 = n2516 | n9155;
assign n554 = n11142 | n3792;
assign n223 = ~(n9743 ^ n7946);
assign n2367 = n6776 & n12708;
assign n7387 = ~(n592 ^ n4845);
assign n4813 = n5909 & n12792;
assign n11475 = n12300 & n10972;
assign n11797 = n1256 | n6285;
assign n2810 = n8485 & n12078;
assign n9571 = n7333 & n1784;
assign n8070 = n9215 & n10927;
assign n13222 = ~(n2524 | n3691);
assign n6896 = ~(n9594 ^ n3621);
assign n620 = n11580 & n9937;
assign n843 = ~(n11100 ^ n4927);
assign n10123 = n12545 | n5924;
assign n5827 = ~n8200;
assign n10049 = ~n5962;
assign n10773 = ~(n5322 ^ n7172);
assign n8593 = n10172 ^ n9137;
assign n7337 = n1389 | n3014;
assign n9832 = n3851 & n12382;
assign n8404 = ~(n7402 ^ n2331);
assign n11523 = ~(n10739 | n5824);
assign n5318 = n7828 | n3888;
assign n7490 = ~(n3855 | n1046);
assign n419 = ~(n5678 | n8684);
assign n9379 = n9656 & n10848;
assign n4406 = n4663 | n1127;
assign n9911 = n12732 | n10319;
assign n4550 = ~(n664 | n5759);
assign n4732 = ~n2737;
assign n2819 = ~(n7989 ^ n977);
assign n917 = ~n3006;
assign n5442 = ~(n972 ^ n11071);
assign n6014 = ~(n345 ^ n8054);
assign n10352 = ~n2758;
assign n12318 = n920 | n9079;
assign n5835 = ~(n1645 ^ n6169);
assign n13031 = ~(n4832 ^ n2586);
assign n12447 = ~(n6338 | n5739);
assign n10869 = ~(n2931 ^ n1980);
assign n4207 = ~(n12735 | n11432);
assign n4597 = ~(n4793 ^ n11622);
assign n5557 = ~(n9920 ^ n9991);
assign n7417 = ~(n10824 ^ n8147);
assign n4287 = ~(n288 | n2628);
assign n3840 = n12222 & n4336;
assign n5182 = ~n12965;
assign n2133 = n1301;
assign n5259 = ~(n5906 ^ n1100);
assign n1042 = ~(n5731 | n11108);
assign n635 = n6069 | n11067;
assign n4972 = ~(n13131 ^ n7108);
assign n2714 = n9690 & n10741;
assign n4911 = ~(n11269 ^ n8196);
assign n5426 = ~(n2935 | n31);
assign n1849 = n12107 & n8907;
assign n5161 = ~(n6396 ^ n7425);
assign n11607 = ~(n9079 ^ n10934);
assign n10247 = ~(n11090 ^ n468);
assign n4046 = ~(n1747 ^ n11145);
assign n1219 = n9115 & n6538;
assign n10684 = ~(n2785 ^ n1895);
assign n12186 = n5707 & n1432;
assign n2967 = ~n3954;
assign n5788 = ~(n5216 | n3751);
assign n78 = n951 & n3085;
assign n4444 = ~(n3740 ^ n9599);
assign n9478 = ~n9747;
assign n116 = ~n13221;
assign n12844 = n8351 | n6532;
assign n9143 = ~(n11901 ^ n10809);
assign n12271 = n8020 | n206;
assign n10424 = ~(n1098 ^ n9766);
assign n3174 = n5040 | n11144;
assign n1023 = n8472 | n3981;
assign n3247 = n12837 | n1325;
assign n5166 = n3770 | n3084;
assign n8272 = n2135 | n894;
assign n2653 = ~(n9994 | n7811);
assign n4842 = ~(n12971 ^ n3470);
assign n12989 = n8176 | n11122;
assign n6136 = n1077 | n3960;
assign n5145 = n10031 | n4226;
assign n4332 = n9228 | n3817;
assign n8751 = n3105 | n6746;
assign n9783 = n6685 | n1458;
assign n11047 = n2299 & n12190;
assign n762 = ~(n12943 ^ n2839);
assign n8414 = n3175 & n8731;
assign n862 = ~(n1951 ^ n12739);
assign n2752 = ~n1055;
assign n709 = ~n4036;
assign n5506 = n12451 | n2402;
assign n5294 = ~n1502;
assign n9797 = n406 | n11950;
assign n7788 = ~(n10585 ^ n2696);
assign n6410 = ~(n1559 ^ n6919);
assign n1825 = n6051 & n11998;
assign n11637 = ~n3521;
assign n10677 = n12056 & n2975;
assign n8512 = n10085 | n7530;
assign n12970 = ~(n471 ^ n9472);
assign n2110 = ~(n10064 | n760);
assign n5011 = n8712 & n11092;
assign n2262 = ~(n11183 ^ n10791);
assign n9476 = n7445 & n216;
assign n3200 = ~(n9505 ^ n10596);
assign n2037 = ~n3244;
assign n8284 = ~(n8812 ^ n9532);
assign n8261 = n197 & n8785;
assign n7749 = ~n9347;
assign n3825 = ~n510;
assign n4073 = n6348 & n6936;
assign n10466 = ~n10390;
assign n2376 = ~(n7556 ^ n12291);
assign n7099 = n6279 & n4634;
assign n12801 = ~(n2925 | n4583);
assign n1396 = n5888 | n6572;
assign n2419 = n9216 & n411;
assign n11513 = n5568 & n12853;
assign n8670 = n3969 & n10945;
assign n10758 = ~(n9234 ^ n10637);
assign n11422 = n12635 & n9922;
assign n9789 = n8598 | n1985;
assign n10276 = n9265 & n9286;
assign n4425 = ~(n10498 ^ n5515);
assign n10176 = ~(n2027 ^ n6728);
assign n6637 = n449 | n10302;
assign n7768 = n3478 & n5537;
assign n4491 = n11037 | n9223;
assign n2438 = ~(n10709 ^ n4413);
assign n12994 = ~n5642;
assign n5761 = ~(n7881 ^ n11477);
assign n4176 = n6778 | n12110;
assign n12249 = ~n11180;
assign n10003 = ~(n12216 ^ n9563);
assign n8365 = ~(n1359 ^ n2438);
assign n12640 = n11707 & n6358;
assign n11108 = n12396 | n6978;
assign n207 = n1345 | n10029;
assign n11190 = ~(n6417 ^ n8399);
assign n12022 = n3127 | n8563;
assign n9991 = ~(n235 ^ n4816);
assign n9808 = ~n11537;
assign n8812 = n5688 | n8030;
assign n6907 = n7918 & n1470;
assign n7205 = ~(n4139 ^ n6698);
assign n910 = n12683 | n10617;
assign n6073 = ~(n1774 ^ n83);
assign n9231 = n8167 & n3341;
assign n12931 = ~(n13200 | n6779);
assign n1648 = n1023 | n5202;
assign n264 = ~(n8593 ^ n8921);
assign n1498 = ~(n7000 ^ n4394);
assign n12264 = n2768 | n4230;
assign n179 = ~(n2010 ^ n7685);
assign n9030 = ~(n5612 | n5413);
assign n10481 = ~n1636;
assign n1675 = n10509 | n4844;
assign n3640 = ~n5536;
assign n10229 = ~n9948;
assign n2555 = n7171 & n11684;
assign n12736 = ~(n3244 ^ n7107);
assign n4462 = ~n9915;
assign n4014 = ~(n8473 ^ n3410);
assign n590 = ~(n3115 ^ n6185);
assign n10204 = ~n1327;
assign n3978 = n13025 | n3981;
assign n7543 = n4621 | n121;
assign n4304 = ~(n10183 ^ n11931);
assign n2575 = n5922 & n7874;
assign n2946 = n1957 | n5408;
assign n11610 = n12417 ^ n10376;
assign n8389 = n5086 | n4515;
assign n3684 = n8106 | n5317;
assign n4865 = n10619 & n300;
assign n10062 = ~(n85 ^ n2857);
assign n551 = n6571 & n11124;
assign n6051 = n3225 | n7935;
assign n5026 = ~(n8620 ^ n8866);
assign n1483 = n8325 | n1043;
assign n10919 = n2614 | n1463;
assign n5630 = ~n8394;
assign n11328 = ~n7040;
assign n12016 = n11754 & n8426;
assign n12738 = ~n9367;
assign n7845 = n12174 | n1043;
assign n3180 = ~(n4797 ^ n9311);
assign n9169 = n2128 | n12910;
assign n3062 = ~n12352;
assign n10544 = n8941 | n10016;
assign n9843 = ~(n1232 ^ n10946);
assign n10665 = ~(n1984 | n8963);
assign n1328 = n5190 | n12787;
assign n13220 = ~(n8579 ^ n4008);
assign n6055 = ~n3286;
assign n995 = ~(n4302 ^ n2539);
assign n4280 = ~(n5417 ^ n4541);
assign n10704 = n2217 | n479;
assign n10064 = n12153 | n776;
assign n4379 = n7672 | n4373;
assign n3203 = n2145 & n7006;
assign n7997 = ~(n622 | n7307);
assign n2779 = ~(n1316 ^ n8395);
assign n2200 = ~(n6298 ^ n12529);
assign n904 = ~(n9539 ^ n5625);
assign n4766 = n10664 | n8519;
assign n7688 = n9281 | n6623;
assign n965 = n8498 | n8268;
assign n3758 = ~(n7896 | n851);
assign n1408 = ~(n12131 ^ n12223);
assign n6538 = ~n12452;
assign n4532 = n3311 & n10408;
assign n7893 = ~(n7542 | n4534);
assign n12097 = n1191 | n1463;
assign n11618 = ~(n2021 ^ n12937);
assign n2011 = n9282 | n7158;
assign n7126 = n6250 | n9159;
assign n12493 = ~n11574;
assign n5394 = ~(n6211 ^ n8388);
assign n6932 = ~(n7284 ^ n4407);
assign n4472 = n250 & n2492;
assign n12576 = ~n5600;
assign n6234 = n10092 & n3368;
assign n4726 = ~(n2344 ^ n4956);
assign n4912 = n2254 | n237;
assign n2530 = n6074 & n11191;
assign n7962 = ~n9514;
assign n10543 = ~(n348 ^ n4177);
assign n11533 = n1634 | n12621;
assign n5948 = n2786 | n8972;
assign n69 = ~n772;
assign n2024 = n3854 | n6404;
assign n5822 = n7319 | n12764;
assign n10734 = n5840 & n101;
assign n5932 = n6439 | n12273;
assign n3779 = n11650 & n1121;
assign n6315 = n5927 | n10292;
assign n7964 = ~(n6777 ^ n10205);
assign n7692 = n9995 & n7598;
assign n10590 = ~n6782;
assign n7427 = n6182 | n9223;
assign n3420 = n2726 | n3949;
assign n5598 = ~(n2706 ^ n687);
assign n3898 = ~n11180;
assign n2411 = ~n12156;
assign n9514 = n11197 & n1078;
assign n9796 = ~(n9930 ^ n2565);
assign n10141 = n2563 | n1509;
assign n10751 = ~(n4948 ^ n268);
assign n7506 = n12778 | n11922;
assign n4590 = ~(n7709 ^ n10000);
assign n3971 = n3018 & n6951;
assign n10754 = n12402 & n10456;
assign n5670 = ~n7812;
assign n3071 = n2381 & n5778;
assign n6777 = n10334 | n10179;
assign n11010 = n4642 | n2626;
assign n2325 = ~n10904;
assign n9769 = n4289 & n8878;
assign n1431 = n2558 | n4056;
assign n1640 = ~(n10782 | n12379);
assign n6343 = n11207 & n3033;
assign n5878 = n10988 & n4831;
assign n5002 = ~n7697;
assign n12235 = ~(n3687 ^ n10803);
assign n12846 = ~n892;
assign n1332 = n5205 | n2907;
assign n3504 = ~(n95 | n146);
assign n9838 = ~n12020;
assign n3892 = ~n2498;
assign n2527 = n5942 & n5892;
assign n8528 = ~(n7845 ^ n13098);
assign n6102 = ~(n7713 ^ n5311);
assign n6618 = n11341 & n1954;
assign n10575 = ~(n1667 ^ n11372);
assign n6635 = n4696;
assign n2742 = ~n1611;
assign n12789 = ~n11030;
assign n11651 = n4185 | n8268;
assign n9450 = ~n10805;
assign n2021 = n3092 & n11740;
assign n7624 = ~(n5938 | n2410);
assign n3941 = ~(n3189 | n682);
assign n4762 = n4759 & n2665;
assign n5409 = ~n8684;
assign n5542 = n4995 | n9792;
assign n10930 = ~(n3880 ^ n11670);
assign n1558 = n2994 & n10713;
assign n2473 = ~n10343;
assign n10042 = ~(n7369 ^ n7808);
assign n2688 = ~n817;
assign n608 = n10580 | n815;
assign n105 = ~(n4038 ^ n4424);
assign n6980 = n6479 | n1653;
assign n12664 = n2175 | n7873;
assign n4729 = n10682 & n10896;
assign n3362 = ~(n3633 ^ n12863);
assign n9181 = ~n1636;
assign n4186 = n139 & n3853;
assign n1079 = ~(n3919 | n12108);
assign n3909 = n5671 & n8290;
assign n10997 = n4087 | n8686;
assign n11359 = ~(n1815 | n3555);
assign n12140 = n4104 & n8186;
assign n1281 = ~(n4589 ^ n11503);
assign n6598 = ~(n11378 ^ n1661);
assign n5309 = ~(n2186 ^ n92);
assign n3781 = n5500 | n11475;
assign n7039 = ~(n1809 | n4287);
assign n1240 = n6721 | n1144;
assign n6617 = ~(n10584 ^ n9911);
assign n821 = ~n6357;
assign n5563 = ~(n3333 ^ n7478);
assign n889 = n5999 | n2599;
assign n3236 = ~(n9042 | n10612);
assign n4283 = n6486 | n4640;
assign n9283 = ~n12373;
assign n4613 = ~(n12697 ^ n7640);
assign n5291 = n12253 & n3486;
assign n5896 = n9113 | n8490;
assign n12273 = n5550;
assign n12867 = ~(n4400 ^ n3994);
assign n10904 = n934 & n6674;
assign n6582 = n8085 & n4679;
assign n6657 = n13168 | n12188;
assign n7119 = ~n3076;
assign n10902 = ~(n8986 | n11601);
assign n2708 = ~(n12355 ^ n12264);
assign n9492 = ~n411;
assign n11387 = n9718 & n5933;
assign n4224 = n8672 | n12188;
assign n7643 = n12130 & n12181;
assign n1280 = n6644 ^ n2547;
assign n11531 = n10491 & n13180;
assign n11365 = ~n1717;
assign n5306 = n1671 | n7323;
assign n7584 = ~(n2219 ^ n7509);
assign n10353 = n207 | n12290;
assign n12993 = n2762 ^ n11154;
assign n1862 = ~(n8690 ^ n6995);
assign n5537 = n2228 | n1570;
assign n519 = n8050 | n663;
assign n8767 = n12667 & n1787;
assign n11442 = n3071 | n341;
assign n3122 = n6769 | n6265;
assign n11972 = ~n11939;
assign n13214 = n10681 | n12596;
assign n5498 = ~(n1603 ^ n3455);
assign n5839 = ~n8311;
assign n7181 = n3908 | n1144;
assign n1731 = ~(n10911 ^ n8201);
assign n3540 = ~(n4147 ^ n1981);
assign n11354 = ~n10642;
assign n10585 = n10586 | n12126;
assign n6449 = n6753 | n8573;
assign n11272 = ~(n7398 ^ n8287);
assign n11766 = ~(n9341 ^ n2161);
assign n30 = n554 & n3975;
assign n3611 = ~(n7767 ^ n10372);
assign n11009 = n7780 | n10106;
assign n12815 = n1070 & n12169;
assign n7015 = n5972 | n4987;
assign n7709 = ~n9515;
assign n10460 = n106 | n1266;
assign n5446 = ~n6707;
assign n12116 = n1973 & n6302;
assign n4632 = ~(n12670 ^ n10971);
assign n6707 = n1402 | n9223;
assign n8534 = n6596;
assign n11540 = ~n8745;
assign n8334 = n10924 | n2787;
assign n8713 = ~(n3796 ^ n5325);
assign n11698 = ~(n11733 ^ n9815);
assign n3612 = ~(n8814 ^ n9560);
assign n4080 = ~n497;
assign n8069 = ~(n3810 ^ n4918);
assign n6648 = ~(n9331 ^ n4625);
assign n822 = n7926 & n1334;
assign n4196 = n1391 & n10967;
assign n12695 = n2278;
assign n6533 = ~n4188;
assign n6605 = ~(n2312 ^ n12685);
assign n11235 = n1402 | n2059;
assign n2917 = n8751 & n8344;
assign n4577 = ~(n8366 ^ n7176);
assign n9402 = ~n7896;
assign n5797 = n2278;
assign n9586 = ~n12248;
assign n2144 = n2538 | n3949;
assign n13066 = n6908 | n5819;
assign n3843 = n5900 & n9781;
assign n5596 = n1332 & n11463;
assign n9443 = n7068 | n9159;
assign n12171 = ~n4651;
assign n4571 = ~(n12981 | n6272);
assign n5244 = ~(n7869 ^ n754);
assign n9106 = n12322 & n12374;
assign n6213 = ~(n7926 ^ n236);
assign n8835 = ~n2577;
assign n6951 = n12469 | n12273;
assign n164 = n4761 & n6013;
assign n12310 = n10775 | n9956;
assign n8373 = ~(n12073 ^ n8003);
assign n3761 = ~n10288;
assign n4279 = n7966 | n6404;
assign n1803 = ~(n5399 | n7405);
assign n9134 = n1652 & n10419;
assign n10035 = ~n2212;
assign n8559 = n6595 | n7935;
assign n10192 = ~(n12518 ^ n12024);
assign n9580 = n3365 ^ n11819;
assign n3733 = ~(n3868 | n11143);
assign n12311 = n5803 | n3193;
assign n158 = ~(n13050 ^ n5106);
assign n3786 = n4451 | n5725;
assign n8843 = ~n1302;
assign n5867 = n11455 | n10374;
assign n825 = ~(n11562 ^ n12497);
assign n10443 = ~(n12437 | n3799);
assign n267 = n10314 | n12959;
assign n2500 = n5207 & n3707;
assign n10564 = n11014 & n4770;
assign n4938 = n7283 | n12273;
assign n4388 = ~(n4500 | n1);
assign n2345 = n3619 | n13053;
assign n10263 = ~n10162;
assign n2370 = n1218 | n5242;
assign n2387 = ~n6168;
assign n5199 = n13063 | n5493;
assign n10519 = ~n12078;
assign n11194 = n7091 | n3438;
assign n1417 = n11420 & n2363;
assign n11817 = n3750 & n11399;
assign n2019 = ~(n10496 | n5159);
assign n5248 = n3325 & n4942;
assign n1068 = n10979 ^ n8875;
assign n8642 = n11703 & n8853;
assign n976 = n2717 & n6920;
assign n3484 = ~(n10967 | n1391);
assign n9351 = ~(n11602 ^ n8100);
assign n11437 = ~(n5621 | n5533);
assign n7203 = ~(n6656 | n10036);
assign n13070 = ~(n914 | n592);
assign n2939 = n9253 & n7972;
assign n3304 = n696 | n9352;
assign n8111 = ~n1792;
assign n408 = n5968 | n10179;
assign n7457 = n1554 | n6133;
assign n6565 = n9757 & n6131;
assign n120 = ~(n12035 ^ n2939);
assign n10638 = ~(n8487 ^ n10394);
assign n8056 = ~(n8061 ^ n6084);
assign n9007 = ~(n1282 ^ n11529);
assign n10790 = ~(n2650 ^ n3569);
assign n2796 = ~(n6536 | n4866);
assign n10666 = ~n594;
assign n5143 = ~(n8942 ^ n6632);
assign n1414 = ~(n5850 ^ n187);
assign n2667 = n4205 & n1351;
assign n9631 = ~(n9708 ^ n684);
assign n11210 = n13194 | n10319;
assign n13183 = ~n2295;
assign n1245 = n1018 & n764;
assign n88 = ~(n7583 ^ n6168);
assign n10610 = n5944 | n7305;
assign n8561 = ~n9093;
assign n4894 = ~(n7657 ^ n6795);
assign n565 = n5588 | n10029;
assign n10646 = n1434 | n3459;
assign n156 = ~n6489;
assign n10954 = ~(n12622 ^ n6470);
assign n12246 = ~n2765;
assign n9985 = ~(n4368 | n7716);
assign n10504 = ~(n3122 ^ n6477);
assign n5503 = n7532 | n6635;
assign n11261 = ~(n6668 | n7812);
assign n3222 = ~n4457;
assign n2617 = n4929 & n12060;
assign n1591 = ~(n676 ^ n6432);
assign n9252 = n3224 & n1888;
assign n11471 = ~n5747;
assign n1164 = ~(n4313 ^ n12029);
assign n9756 = ~(n11160 ^ n8069);
assign n10156 = ~(n1380 ^ n5254);
assign n10351 = n10587 | n9159;
assign n11822 = n10136 & n3174;
assign n5337 = n5558 | n13043;
assign n10558 = ~n12579;
assign n3186 = n2931 & n7313;
assign n12991 = ~(n331 ^ n11994);
assign n3075 = ~(n12381 | n4589);
assign n9033 = ~n5498;
assign n10383 = ~n2174;
assign n2938 = n10631 & n10329;
assign n535 = ~(n10327 ^ n10074);
assign n2139 = ~(n9945 ^ n3513);
assign n12907 = ~(n6273 | n12145);
assign n12034 = ~(n9039 ^ n2775);
assign n1970 = n513 | n9027;
assign n11305 = ~(n3834 ^ n9411);
assign n8015 = ~(n9870 ^ n1104);
assign n7669 = n11781 | n902;
assign n8644 = ~n9474;
assign n7321 = n1126 & n13083;
assign n493 = ~n12853;
assign n4812 = n12569 & n7508;
assign n10806 = n9619 & n5382;
assign n2250 = n2753 & n7593;
assign n5494 = ~n6043;
assign n2023 = n2725 & n13228;
assign n12776 = ~(n7316 ^ n4510);
assign n11303 = ~(n2656 ^ n323);
assign n1263 = ~n4789;
assign n7420 = n1485 | n5931;
assign n8813 = ~(n11278 ^ n8482);
assign n7013 = ~n4259;
assign n4 = n11242 | n2133;
assign n8825 = n2504 | n8563;
assign n12812 = ~n10654;
assign n2909 = ~(n2069 ^ n9030);
assign n7637 = ~(n8358 ^ n3087);
assign n10525 = ~n1988;
assign n7764 = ~(n10812 ^ n5074);
assign n1121 = ~(n6555 ^ n12338);
assign n8654 = ~n9580;
assign n5998 = n5659 ^ n11988;
assign n4145 = n8510 | n8702;
assign n13009 = n10558 | n7723;
assign n9553 = ~(n7555 ^ n2864);
assign n4389 = n11249 & n13207;
assign n11115 = n5574 | n5604;
assign n1583 = ~(n6305 ^ n984);
assign n2751 = n1905 & n2608;
assign n8026 = ~n1498;
assign n10988 = ~n13034;
assign n3678 = ~(n2431 ^ n11169);
assign n2580 = ~n11671;
assign n4626 = ~(n7585 ^ n9947);
assign n2888 = ~(n4035 ^ n8902);
assign n7771 = ~n12340;
assign n1794 = n12230 & n4204;
assign n8668 = n7000 | n10937;
assign n8459 = ~(n11899 ^ n2926);
assign n2015 = n2031 | n10130;
assign n3326 = n950 | n3257;
assign n2613 = n10474 | n5782;
assign n7700 = ~n13060;
assign n7353 = n5883 & n7653;
assign n3179 = ~(n10259 | n12454);
assign n5441 = n5973 | n8563;
assign n3995 = n103 & n10408;
assign n5233 = n9606 | n12188;
assign n3559 = n6135 & n4859;
assign n3334 = ~n11386;
assign n10074 = ~(n6711 ^ n2523);
assign n10096 = n6726 | n7530;
assign n9126 = ~(n6431 | n8826);
assign n4060 = ~(n5098 ^ n3647);
assign n1200 = n13181 | n1589;
assign n7105 = n6658 | n7221;
assign n3716 = n8471 & n6688;
assign n9657 = n11313 & n883;
assign n3717 = ~(n4710 | n3840);
assign n9118 = ~n5962;
assign n5139 = n6595 | n7903;
assign n5722 = n10144 & n8545;
assign n6739 = n3465 | n10222;
assign n9765 = ~n4968;
assign n10576 = ~(n12994 | n4422);
assign n3748 = ~(n9151 ^ n2664);
assign n4240 = ~(n1116 ^ n3670);
assign n1868 = n8392 | n9159;
assign n11361 = n1360 | n3531;
assign n8834 = ~n90;
assign n7212 = ~(n7427 ^ n9203);
assign n9697 = ~n2011;
assign n12930 = ~n4470;
assign n6413 = ~(n2739 ^ n975);
assign n1993 = ~(n5025 ^ n523);
assign n12650 = ~(n9974 ^ n11747);
assign n11242 = ~n12408;
assign n3702 = n13163 & n2440;
assign n8504 = ~n429;
assign n2442 = n813 | n10029;
assign n10271 = ~(n6539 ^ n12257);
assign n8039 = ~n5513;
assign n4623 = ~(n9168 ^ n9639);
assign n2630 = n11366 ^ n4269;
assign n9265 = ~n10231;
assign n11781 = ~n4470;
assign n5713 = ~n12651;
assign n7657 = n6733 | n1570;
assign n10957 = ~(n8417 | n10011);
assign n9025 = n7184 | n6635;
assign n13242 = ~n11537;
assign n4680 = ~n3447;
assign n7577 = n5544 ^ n10149;
assign n11462 = n10429 | n252;
assign n9817 = ~(n12797 ^ n4726);
assign n11882 = ~(n8520 ^ n4329);
assign n5384 = ~(n8811 ^ n6932);
assign n10851 = n2985 | n9704;
assign n12040 = ~(n8794 ^ n11814);
assign n8001 = n7065 & n12180;
assign n6768 = ~n4006;
assign n2531 = ~(n12710 | n4193);
assign n7346 = ~n5933;
assign n6281 = n3363 & n2680;
assign n6197 = n10796 ^ n12058;
assign n1136 = n10900 | n2449;
assign n6421 = ~n7670;
assign n585 = ~n1432;
assign n6294 = ~(n6130 ^ n8780);
assign n9295 = n7269 & n9342;
assign n7850 = n5595 | n2875;
assign n5927 = ~n10004;
assign n11604 = ~(n11655 ^ n738);
assign n3856 = n7941 | n4868;
assign n5711 = n3697 | n7655;
assign n4246 = ~(n11987 ^ n3019);
assign n1088 = ~(n11998 ^ n6051);
assign n617 = ~n8233;
assign n12644 = ~(n15 ^ n3056);
assign n5411 = n2013 | n6484;
assign n8566 = n11258 & n11967;
assign n4753 = n7124 | n11550;
assign n4965 = n13084 | n12501;
assign n2943 = ~n13058;
assign n4954 = n3128 & n3203;
assign n6476 = ~(n3627 ^ n13212);
assign n8269 = ~(n10999 ^ n10342);
assign n8618 = n4584 | n4373;
assign n415 = ~(n9261 ^ n11977);
assign n12335 = ~n12003;
assign n11208 = ~(n1205 | n2649);
assign n3952 = ~(n12362 ^ n3987);
assign n7983 = ~(n1395 | n8781);
assign n3482 = ~(n10371 ^ n13015);
assign n2700 = n579 & n7977;
assign n9884 = n7018 | n3016;
assign n1656 = ~(n2107 | n8548);
assign n452 = n216 | n7445;
assign n241 = ~n9534;
assign n13169 = n2711 | n9268;
assign n8004 = ~(n12186 | n6163);
assign n12422 = n7919 ^ n11056;
assign n4818 = ~n1612;
assign n4927 = n5666 | n12273;
assign n12923 = ~(n8889 ^ n6022);
assign n2792 = n5923 | n1026;
assign n6835 = n3347 | n5036;
assign n11142 = n4514 | n11244;
assign n1888 = n1621 | n2133;
assign n1152 = ~n10451;
assign n10316 = n3587 | n9223;
assign n7000 = ~(n8028 ^ n4162);
assign n3850 = ~(n3628 ^ n9218);
assign n2941 = ~n5066;
assign n6012 = n11886 & n4025;
assign n8839 = ~(n4876 ^ n769);
assign n8445 = n3732 & n7438;
assign n7429 = n9332 & n5818;
assign n6712 = n5890 | n8534;
assign n11315 = n12514 | n514;
assign n3955 = ~(n11306 | n8432);
assign n11605 = ~n7326;
assign n1536 = ~n8332;
assign n1455 = ~(n9236 ^ n5023);
assign n10526 = n12517 & n7303;
assign n11319 = ~(n8800 ^ n7628);
assign n12018 = n13061 | n1212;
assign n7142 = ~n1198;
assign n5923 = ~n5189;
assign n7798 = ~n2339;
assign n2900 = n8556 | n11772;
assign n12014 = n1268 ^ n3865;
assign n9686 = n11943 & n2305;
assign n581 = n4737 & n1785;
assign n11192 = n2689 | n8702;
assign n432 = n8141 | n11510;
assign n8125 = n8183 & n5920;
assign n6562 = n4905 & n10703;
assign n2400 = n1406 | n5999;
assign n5890 = ~n2737;
assign n1782 = n3266 & n2224;
assign n2096 = n5004 | n4314;
assign n10554 = ~(n10921 ^ n11675);
assign n8836 = ~n3116;
assign n3550 = n1669 & n1185;
assign n2921 = ~(n2439 ^ n1049);
assign n12406 = ~(n1655 ^ n10082);
assign n12505 = ~(n12867 | n11079);
assign n7717 = ~(n6009 ^ n9055);
assign n8664 = ~n7090;
assign n4538 = n7142 | n2675;
assign n6602 = n8697 | n10648;
assign n4097 = n6988 | n11591;
assign n9644 = ~(n3848 ^ n7484);
assign n7425 = ~(n11189 ^ n6512);
assign n11069 = n10954 | n4504;
assign n6484 = n6132 ^ n6094;
assign n9183 = ~(n4224 ^ n9864);
assign n2561 = ~(n6690 ^ n7141);
assign n3908 = ~n6655;
assign n10024 = n10800 & n8019;
assign n7422 = ~(n744 | n12484);
assign n8020 = ~n1709;
assign n2723 = ~n8768;
assign n11706 = n1387 | n4565;
assign n12552 = ~n11891;
assign n4319 = ~(n9213 ^ n7651);
assign n9828 = ~n1573;
assign n6831 = ~(n4146 ^ n4623);
assign n10720 = ~(n9519 ^ n6541);
assign n7063 = ~(n4012 | n8189);
assign n6192 = ~(n978 ^ n11009);
assign n5459 = n11718 | n5081;
assign n10330 = ~(n7763 ^ n5578);
assign n10210 = ~n7637;
assign n948 = ~(n10795 ^ n12667);
assign n4826 = n12441 | n4063;
assign n1232 = n1420 & n8387;
assign n137 = ~(n3069 ^ n8365);
assign n8807 = ~(n12472 ^ n1926);
assign n3041 = ~n9381;
assign n5147 = ~(n2814 ^ n12123);
assign n5511 = n9422 | n1109;
assign n11390 = ~(n7002 ^ n7308);
assign n10157 = n11903 | n5765;
assign n3814 = n555 | n5677;
assign n6645 = ~n3645;
assign n1324 = ~n4233;
assign n5243 = ~n741;
assign n1406 = ~n9887;
assign n400 = n2566 | n7624;
assign n8689 = n1495 ^ n4518;
assign n3057 = ~(n3394 ^ n12392);
assign n12053 = ~(n672 | n2912);
assign n1779 = n9767 | n8030;
assign n12456 = ~(n8470 | n5469);
assign n1361 = n10232 & n9520;
assign n12099 = ~n9849;
assign n3545 = n3369 | n6227;
assign n70 = ~(n7240 ^ n735);
assign n5649 = n12834 | n2449;
assign n5677 = n8663 & n6476;
assign n12133 = n8466 & n7720;
assign n1100 = ~(n6842 ^ n86);
assign n3439 = n7377 | n9075;
assign n3481 = n12418 & n11713;
assign n10492 = ~n12389;
assign n12726 = n10772 | n11144;
assign n1249 = ~(n9056 ^ n7612);
assign n1208 = ~(n12824 ^ n6897);
assign n3509 = ~n3112;
assign n11156 = n7891 | n8048;
assign n5178 = ~(n3354 ^ n10367);
assign n4700 = n12838 & n4479;
assign n6159 = n6738 | n9486;
assign n80 = ~n951;
assign n4128 = n10281 | n206;
assign n7568 = n8035 | n6565;
assign n6310 = ~(n4277 ^ n9908);
assign n6453 = n7033 | n5521;
assign n6219 = ~n841;
assign n2826 = n79 | n4442;
assign n6953 = n12000 | n4253;
assign n6748 = n3892 | n12069;
assign n11001 = ~(n10918 ^ n3528);
assign n7663 = ~(n4772 ^ n12495);
assign n8958 = ~(n11064 ^ n5237);
assign n1344 = n3602 & n6807;
assign n2070 = n8950 | n6635;
assign n13134 = n5520 | n10761;
assign n10359 = n1706 | n4643;
assign n356 = n8221 & n7261;
assign n276 = ~(n9456 | n1754);
assign n8089 = ~(n10690 ^ n10095);
assign n8285 = ~n6142;
assign n8971 = ~n253;
assign n6706 = ~n1486;
assign n2195 = n13056 & n385;
assign n2935 = n521 & n11039;
assign n876 = n5125 | n12077;
assign n12369 = ~(n7889 ^ n2685);
assign n11106 = ~n12784;
assign n11894 = ~(n2851 ^ n9121);
assign n6890 = n11009 | n12387;
assign n374 = n7017 & n1970;
assign n11762 = ~(n921 ^ n10650);
assign n7712 = ~(n9448 | n6483);
assign n6622 = ~(n6208 ^ n352);
assign n8620 = n6846 | n3703;
assign n9854 = n12084 | n13054;
assign n2719 = ~(n13223 ^ n12822);
assign n47 = ~n5551;
assign n9716 = n1903 | n10931;
assign n1460 = n7047 | n12783;
assign n2928 = ~(n6527 ^ n7278);
assign n12848 = ~n13120;
assign n325 = n5031 & n8506;
assign n8683 = n2232 | n2958;
assign n8344 = n1559 | n6919;
assign n1683 = n1571 | n7530;
assign n9069 = ~n6392;
assign n38 = n6672 | n13238;
assign n6723 = n5943 | n8730;
assign n3876 = ~(n3536 ^ n6857);
assign n4553 = ~(n10790 ^ n4083);
assign n2202 = ~(n12394 ^ n11863);
assign n7861 = n7620 | n9195;
assign n4320 = n7529 & n7772;
assign n12694 = n231 & n8906;
assign n8592 = ~n4008;
assign n2320 = ~(n12260 | n11433);
assign n5009 = n4184 | n12725;
assign n12742 = n8839 ^ n1281;
assign n6806 = n11599 | n7892;
assign n8409 = ~(n3642 ^ n5196);
assign n5176 = ~n8768;
assign n2415 = ~n4740;
assign n4788 = n4803 ^ n256;
assign n523 = n12918 & n5246;
assign n7487 = ~(n10913 | n3746);
assign n3498 = ~n4470;
assign n12005 = n10851 & n3275;
assign n5781 = n9509 & n357;
assign n8991 = ~(n9448 ^ n7389);
assign n8403 = ~(n4654 ^ n1958);
assign n3891 = ~(n7474 | n4068);
assign n4417 = ~(n9554 ^ n3849);
assign n440 = n12871 | n12388;
assign n3087 = n6769 | n1026;
assign n10079 = n7331 & n5204;
assign n8436 = ~n12603;
assign n4835 = n13215 & n150;
assign n11725 = ~(n9523 ^ n11656);
assign n7706 = n6724 | n7723;
assign n3370 = ~(n4251 ^ n3079);
assign n10986 = ~n11445;
assign n4614 = ~(n4101 ^ n9357);
assign n2207 = ~n8455;
assign n5296 = n4667 & n10546;
assign n3901 = n7884 | n12426;
assign n9933 = n10228 & n3915;
assign n9821 = ~n8036;
assign n10399 = ~(n10499 ^ n6893);
assign n1763 = n3299 | n8301;
assign n3324 = ~(n6294 ^ n3034);
assign n13045 = ~(n5505 | n13171);
assign n8672 = ~n9669;
assign n4361 = ~n1228;
assign n1770 = n5314 & n188;
assign n4687 = n9153 & n12001;
assign n2266 = n8528 | n13237;
assign n5105 = ~n4006;
assign n11746 = n9928 & n9445;
assign n7159 = ~n3064;
assign n12628 = ~(n786 | n4428);
assign n632 = ~(n12637 ^ n2046);
assign n3025 = ~n7316;
assign n46 = n2826 & n10965;
assign n1743 = ~(n8689 ^ n6516);
assign n1618 = ~n7720;
assign n10319 = n13005;
assign n833 = ~(n2088 | n5851);
assign n6594 = ~(n12707 | n5333);
assign n3783 = ~n7360;
assign n12771 = n11171 | n12273;
assign n2152 = n3345 & n8112;
assign n8818 = ~(n10920 ^ n5975);
assign n3132 = ~n3711;
assign n1856 = ~(n10033 | n8669);
assign n5071 = n2652 & n11369;
assign n1226 = ~n1312;
assign n7528 = n8146 & n169;
assign n485 = n2535 ^ n11741;
assign n12956 = ~(n11567 ^ n4999);
assign n4093 = n10760 & n5330;
assign n1750 = ~n8228;
assign n504 = n3445 & n6581;
assign n7213 = n7249 | n2836;
assign n11989 = n10525 | n2212;
assign n4143 = ~n7113;
assign n323 = n508 & n6393;
assign n7043 = ~(n10743 ^ n6529);
assign n7588 = n2858 | n8097;
assign n3070 = n1571 | n12388;
assign n10516 = ~(n11893 ^ n6350);
assign n11276 = ~(n1547 ^ n466);
assign n10940 = n1930 | n8348;
assign n9542 = ~(n4204 ^ n4241);
assign n5311 = n4096 & n9072;
assign n2302 = n4692 | n2351;
assign n11846 = n9216 & n13058;
assign n4433 = n6713 | n2989;
assign n3227 = n9723 | n8030;
assign n7112 = n4430 | n68;
assign n6283 = ~(n36 ^ n5219);
assign n6794 = ~(n1935 ^ n9587);
assign n8627 = n1021 & n8628;
assign n7740 = ~(n2233 ^ n1421);
assign n3681 = ~n8543;
assign n3683 = n10481 | n9075;
assign n637 = ~(n382 ^ n3967);
assign n6897 = ~(n5188 ^ n13022);
assign n7630 = n8396 & n11383;
assign n1322 = ~(n8539 | n3525);
assign n12672 = n7894 & n6300;
assign n12457 = ~(n3345 ^ n580);
assign n7658 = n1571 | n8702;
assign n5367 = n5810 | n3133;
assign n10291 = ~n9667;
assign n5144 = n3516 | n5547;
assign n11796 = n4870 & n9487;
assign n3963 = ~n3130;
assign n2283 = n7223 | n3981;
assign n10442 = n5644 & n7179;
assign n6079 = ~(n7669 ^ n10767);
assign n1321 = ~n2630;
assign n10877 = ~n4357;
assign n12225 = n1797 & n9722;
assign n12511 = n7771 & n3524;
assign n11014 = ~n5777;
assign n3823 = ~(n12675 | n3629);
assign n7824 = ~n4543;
assign n10436 = n993 & n6353;
assign n750 = ~(n1442 ^ n9967);
assign n2966 = ~(n877 ^ n12991);
assign n2735 = ~(n13172 ^ n2567);
assign n7167 = ~n11634;
assign n4560 = n4779 & n7832;
assign n9743 = n9822 | n634;
assign n10329 = n2914 | n655;
assign n11297 = ~n10633;
assign n9868 = ~n9570;
assign n11433 = n6915 | n1710;
assign n11267 = n4532 & n7279;
assign n4262 = ~(n6321 ^ n5780);
assign n6095 = n3420 | n6123;
assign n12459 = ~(n12659 ^ n5351);
assign n12794 = ~(n4112 | n4389);
assign n8841 = ~(n6384 ^ n13142);
assign n2251 = ~(n11775 | n12139);
assign n2319 = n8802 & n6235;
assign n9431 = ~n3012;
assign n2582 = ~n9887;
assign n4926 = ~(n9624 | n4914);
assign n8955 = ~(n7264 ^ n1208);
assign n7859 = n1680 & n451;
assign n8435 = n2694 & n12528;
assign n2934 = ~(n8495 ^ n11048);
assign n50 = ~(n10695 ^ n12331);
assign n3163 = n6774 | n10875;
assign n12946 = ~(n3345 | n8112);
assign n6121 = ~(n9548 | n1124);
assign n1543 = n11174 & n13052;
assign n8581 = ~(n8652 ^ n658);
assign n11016 = n3442 & n2191;
assign n9268 = ~n9732;
assign n13131 = ~(n833 | n12706);
assign n9515 = n841 ^ n6734;
assign n11329 = n4022 | n206;
assign n5947 = ~n8860;
assign n3387 = ~n7436;
assign n8750 = ~(n12979 ^ n12589);
assign n7097 = ~(n8548 ^ n2107);
assign n1801 = ~(n3436 ^ n1157);
assign n4050 = ~(n9629 | n6253);
assign n2020 = n9158 & n6902;
assign n129 = n7987 & n12556;
assign n10698 = n12009 | n4947;
assign n11545 = ~n3361;
assign n6603 = ~(n6654 ^ n5180);
assign n9826 = n4620 | n6265;
assign n183 = n11473 ^ n2047;
assign n6065 = n6332 | n2675;
assign n8394 = ~(n7822 ^ n9603);
assign n8350 = n1816 | n10367;
assign n6308 = ~n9394;
assign n11630 = n11134 | n816;
assign n5106 = ~(n9859 ^ n5830);
assign n12134 = n2330 & n7320;
assign n6867 = ~(n3289 ^ n8765);
assign n329 = n10877 | n2675;
assign n5819 = ~(n6647 | n6052);
assign n7851 = ~(n5273 ^ n8379);
assign n8286 = n12264 | n12355;
assign n13130 = ~(n11002 | n3930);
assign n6473 = n4914 & n9624;
assign n2689 = ~n2498;
assign n4172 = n5597 & n5846;
assign n12094 = ~(n4554 ^ n8927);
assign n9547 = ~(n3404 ^ n7704);
assign n4935 = ~(n8737 ^ n1244);
assign n11230 = ~n8616;
assign n12159 = ~n12605;
assign n990 = n6493 & n6517;
assign n9779 = ~(n2081 ^ n9681);
assign n10531 = n3393 & n6812;
assign n7365 = ~(n1821 ^ n8298);
assign n636 = n7900 | n4640;
assign n13226 = ~n10733;
assign n3596 = n7133 | n1043;
assign n3607 = ~(n6413 ^ n12562);
assign n360 = ~(n10204 | n3876);
assign n7179 = n11801 | n1901;
assign n6736 = ~(n5071 ^ n1133);
assign n1742 = n6950 & n10002;
assign n8150 = n9617 & n10359;
assign n6516 = ~(n9833 ^ n9544);
assign n221 = ~(n10745 ^ n5457);
assign n11007 = ~n834;
assign n11246 = ~(n3308 ^ n2349);
assign n2746 = n12911 & n2792;
assign n11729 = ~n2737;
assign n5928 = ~(n4451 ^ n2308);
assign n12963 = n8573 & n6753;
assign n8785 = n11933 | n206;
assign n9739 = ~n11734;
assign n10614 = ~(n5319 ^ n12005);
assign n12379 = n9848 & n7807;
assign n6236 = n691 | n2941;
assign n11113 = ~n12065;
assign n3086 = ~(n4874 ^ n7692);
assign n770 = n8905 & n12625;
assign n11964 = ~(n12083 | n2478);
assign n11585 = ~(n3668 ^ n6560);
assign n8087 = ~(n8170 ^ n662);
assign n3287 = n6187 & n4072;
assign n3308 = ~(n8025 | n9865);
assign n2519 = ~(n7558 ^ n5682);
assign n12625 = ~n9903;
assign n11751 = ~n8768;
assign n10952 = ~(n12440 ^ n1541);
assign n12708 = n9728 | n11555;
assign n10307 = ~(n6479 ^ n5315);
assign n6570 = ~(n5660 ^ n10562);
assign n9047 = ~(n8914 | n7296);
assign n6912 = n11168 | n590;
assign n9314 = ~(n2294 | n12228);
assign n7460 = ~n8031;
assign n6469 = ~n4217;
assign n7760 = n3492 & n8286;
assign n5858 = ~(n1534 ^ n3292);
assign n10888 = n5086 | n12814;
assign n9934 = ~n11634;
assign n2488 = ~(n9571 ^ n12149);
assign n2947 = n10166 | n6497;
assign n2404 = ~n1929;
assign n10993 = n154 | n776;
assign n3507 = n4880 | n10659;
assign n10015 = n9353 & n834;
assign n5893 = n8660 | n2938;
assign n3144 = n10392 & n9655;
assign n6317 = n1931 & n4666;
assign n343 = ~n504;
assign n718 = ~(n2307 | n9258);
assign n10130 = ~(n3973 | n11185);
assign n3565 = ~n7288;
assign n1177 = ~(n9050 ^ n10080);
assign n7869 = n4944 | n12298;
assign n3193 = n9632 | n8268;
assign n4963 = n618 | n9858;
assign n8706 = ~(n6072 | n10840);
assign n10076 = ~(n12699 ^ n11363);
assign n4896 = n6578 & n6712;
assign n7982 = n4527 & n9067;
assign n448 = ~n13003;
assign n5188 = ~(n5574 ^ n5764);
assign n12978 = n12283 & n11543;
assign n9423 = ~(n10568 | n12520);
assign n2467 = ~(n3367 ^ n3938);
assign n1756 = n4129 & n11862;
assign n4149 = ~n397;
assign n7841 = ~(n498 ^ n9459);
assign n11214 = ~(n1942 | n2115);
assign n11050 = ~(n7214 ^ n1237);
assign n778 = n13036 | n4640;
assign n3674 = ~n3411;
assign n6510 = n7798 | n8268;
assign n11167 = ~(n865 | n8055);
assign n7780 = ~n10594;
assign n8961 = n3660 | n8958;
assign n4591 = n9313 ^ n764;
assign n8073 = n2913 | n12654;
assign n6010 = ~(n12809 | n12066);
assign n6640 = n4625 | n9331;
assign n3620 = n8471 | n6688;
assign n342 = n3163 & n286;
assign n86 = ~(n11831 ^ n10647);
assign n426 = ~(n4986 ^ n4626);
assign n3246 = ~(n624 | n12752);
assign n3074 = ~(n9614 ^ n1581);
assign n12145 = ~n11335;
assign n12480 = ~(n4309 ^ n8999);
assign n997 = n4382 & n1724;
assign n11412 = ~(n1096 ^ n5575);
assign n1304 = ~(n11917 ^ n1339);
assign n6344 = n10511 & n3360;
assign n12243 = ~n9315;
assign n3040 = n6056 | n9492;
assign n1454 = ~(n1921 | n933);
assign n2188 = ~(n1340 ^ n9840);
assign n6468 = n9228 | n12273;
assign n12089 = n1842 & n6697;
assign n9984 = n9659 & n395;
assign n10640 = n10021 | n2222;
assign n4058 = ~n8467;
assign n204 = ~n9762;
assign n8085 = n1089 | n8143;
assign n5326 = ~(n3571 ^ n3517);
assign n8802 = n63 | n2544;
assign n13107 = ~(n13008 | n4637);
assign n12879 = n185 | n4431;
assign n8795 = n7162 & n7769;
assign n6415 = ~(n7157 ^ n9742);
assign n3433 = n5188 & n9637;
assign n6171 = ~n7829;
assign n7098 = n3643 | n6544;
assign n4173 = n868 | n8269;
assign n4641 = ~(n10762 | n1675);
assign n12658 = n2606 | n11422;
assign n11965 = ~n5320;
assign n9444 = ~n6392;
assign n7934 = n3460 | n6635;
assign n12124 = n7074 | n5242;
assign n11054 = ~n4006;
assign n1050 = n13090 | n12415;
assign n3415 = n3142 | n2320;
assign n6503 = n7825 | n10029;
assign n2992 = ~(n13056 ^ n3021);
assign n10246 = ~(n7712 | n7389);
assign n13151 = ~(n2602 ^ n13147);
assign n4804 = n2854 | n2853;
assign n3726 = ~n9887;
assign n3831 = n9216 & n5920;
assign n4634 = n8671 | n5796;
assign n12663 = ~n8923;
assign n4209 = ~n287;
assign n624 = ~(n12267 ^ n9495);
assign n12602 = n9061 ^ n5876;
assign n8252 = n6958 | n12360;
assign n5223 = n6634 & n7547;
assign n194 = n1413 & n9398;
assign n6576 = n4814 | n8584;
assign n12937 = ~(n5752 ^ n12827);
assign n4392 = n168 & n1245;
assign n12396 = ~(n4788 | n8122);
assign n10604 = ~(n656 | n9514);
assign n486 = n9653 & n1979;
assign n1370 = ~n11734;
assign n12921 = n354 | n12934;
assign n4636 = n809 & n7404;
assign n1939 = ~(n10351 ^ n1788);
assign n5687 = n9010 | n121;
assign n7563 = ~(n12774 ^ n6228);
assign n5579 = n12124 | n7437;
assign n5116 = ~(n2665 ^ n7992);
assign n4615 = ~(n4102 ^ n8528);
assign n8104 = n12419 & n790;
assign n6198 = n1191 | n2544;
assign n2426 = ~(n4279 ^ n7348);
assign n12558 = n3428 | n4230;
assign n10254 = n5310 & n5630;
assign n2353 = n186 | n7551;
assign n316 = n7529 & n5729;
assign n9133 = n2692 | n5242;
assign n3330 = n13013 | n4454;
assign n4474 = n7973 & n4963;
assign n8578 = ~n1423;
assign n3704 = ~(n12756 ^ n9408);
assign n12015 = ~(n9927 ^ n10493);
assign n8908 = ~(n4025 ^ n11886);
assign n5104 = ~(n11445 ^ n3055);
assign n6770 = ~n10408;
assign n11855 = ~(n2831 ^ n5826);
assign n10571 = n11680 | n9195;
assign n3688 = n2630 | n561;
assign n11860 = n289 & n7934;
assign n2634 = n2950 | n5945;
assign n12086 = ~n5659;
assign n6327 = ~n10105;
assign n6186 = ~n9058;
assign n887 = n5731 ^ n2314;
assign n3202 = n7253 & n8531;
assign n9468 = n8575 | n12423;
assign n9424 = n4778 | n11491;
assign n5118 = n10202 | n8226;
assign n3703 = ~n10642;
assign n9885 = ~n2350;
assign n2926 = ~(n383 ^ n3177);
assign n1600 = ~(n2812 ^ n3207);
assign n4291 = ~(n5365 ^ n4892);
assign n6390 = n636 & n9365;
assign n1575 = n11114 | n1012;
assign n4686 = ~n8139;
assign n5486 = ~(n1079 ^ n1616);
assign n2950 = n10188 | n2958;
assign n912 = n5430 | n9075;
assign n3526 = n7130 & n5489;
assign n2235 = ~(n1543 ^ n426);
assign n11152 = ~n2590;
assign n10579 = ~(n7635 | n12087);
assign n12445 = n10588 | n9744;
assign n10668 = n10253 | n6703;
assign n5254 = ~(n6588 ^ n1115);
assign n8773 = ~(n10069 | n5419);
assign n10238 = ~(n4837 ^ n8013);
assign n9952 = n9552 & n5608;
assign n7100 = n4377 & n10633;
assign n9393 = ~(n4952 | n1133);
assign n7189 = ~(n8300 ^ n148);
assign n1479 = ~(n891 ^ n2082);
assign n9278 = ~(n5879 | n13176);
assign n3597 = n1571 | n1026;
assign n9357 = ~(n4306 ^ n4362);
assign n2931 = ~(n10984 ^ n9547);
assign n3882 = ~(n4035 | n3912);
assign n12646 = n1230 | n9699;
assign n12575 = n5272 & n5194;
assign n7412 = n8472 | n8563;
assign n10297 = ~(n11603 ^ n12776);
assign n10535 = ~n7479;
assign n8123 = n1912 & n12263;
assign n10667 = n7410 & n8070;
assign n12278 = ~(n4233 ^ n8966);
assign n177 = n6210;
assign n6363 = n4221 | n6769;
assign n7135 = ~n10594;
assign n12056 = ~(n3444 ^ n838);
assign n9162 = ~n8332;
assign n4411 = n11701 & n11194;
assign n9456 = ~(n382 | n3967);
assign n8808 = n7680 | n12818;
assign n993 = n3195 | n10470;
assign n12669 = ~(n11550 ^ n2458);
assign n10080 = ~(n1765 ^ n8393);
assign n1381 = ~(n10148 | n8232);
assign n3661 = n11080 | n10155;
assign n2340 = ~(n10609 ^ n13126);
assign n9403 = n5853 | n5658;
assign n2238 = n7672 | n7221;
assign n6256 = ~(n6951 ^ n3018);
assign n9964 = n9700 | n4652;
assign n4573 = n2504 | n2276;
assign n6726 = ~n8859;
assign n11937 = n3516 | n559;
assign n8024 = ~n1364;
assign n3471 = ~(n778 | n10704);
assign n5039 = n11018 | n9159;
assign n9425 = ~(n13171 ^ n5555);
assign n205 = ~n6484;
assign n1652 = ~n2000;
assign n11697 = ~n3352;
assign n2225 = n8729 | n9159;
assign n2336 = ~(n6191 ^ n1894);
assign n2412 = ~n9924;
assign n3194 = ~n11709;
assign n11323 = ~n13172;
assign n599 = n9676 | n5817;
assign n10184 = n10616 | n11578;
assign n5984 = n4756 & n2901;
assign n4728 = n6260 & n2918;
assign n3088 = ~(n11030 ^ n11488);
assign n7437 = ~(n6283 ^ n12779);
assign n2053 = n5348 & n6523;
assign n334 = ~n401;
assign n2476 = ~(n5649 ^ n1685);
assign n11520 = ~(n7197 | n4447);
assign n1465 = n10975 & n6352;
assign n5432 = n5988 & n6992;
assign n9809 = ~n12276;
assign n12837 = ~n12482;
assign n6286 = n10719 & n9454;
assign n2724 = ~(n7360 ^ n10818);
assign n8942 = ~(n7823 ^ n9875);
assign n481 = n13066 & n4468;
assign n11885 = n6772 & n8574;
assign n6691 = ~(n9391 ^ n9057);
assign n10889 = ~(n5816 ^ n6642);
assign n6799 = ~(n12008 | n1863);
assign n7650 = n10334 | n11668;
assign n8429 = ~(n5599 | n6613);
assign n3953 = ~(n6114 ^ n4839);
assign n3940 = ~n12651;
assign n8328 = ~(n12627 ^ n7079);
assign n10387 = ~(n259 | n12138);
assign n7949 = n2140 | n620;
assign n1764 = ~(n11684 ^ n2309);
assign n1528 = n5214 & n3409;
assign n5935 = ~(n3013 ^ n11410);
assign n281 = n9969 | n7732;
assign n5396 = ~(n3475 ^ n11932);
assign n9549 = n11646 & n9976;
assign n8034 = n9288 & n10006;
assign n2310 = n2669 | n6635;
assign n9017 = ~n11222;
assign n4619 = n12926 | n8341;
assign n6116 = ~(n11059 ^ n13091);
assign n3782 = n10241 & n10959;
assign n5605 = ~(n6518 ^ n557);
assign n6589 = n5531 & n5602;
assign n5329 = ~(n3159 ^ n12507);
assign n3241 = n9465 | n9772;
assign n7252 = n8560 & n6365;
assign n9712 = ~n3850;
assign n1544 = ~n6570;
assign n11157 = ~n7411;
assign n8531 = n5095 | n2205;
assign n9836 = ~(n2485 ^ n12752);
assign n11821 = n7446 | n5223;
assign n7636 = ~n1384;
assign n3316 = n481 | n10899;
assign n708 = n6238 & n2137;
assign n12424 = n4964 & n2339;
assign n10853 = ~(n9965 ^ n10831);
assign n3598 = ~n12853;
assign n4369 = ~(n11401 ^ n6899);
assign n11241 = n3496 | n6966;
assign n10837 = n7809 | n13232;
assign n5245 = ~n11064;
assign n7265 = ~(n9530 ^ n13057);
assign n6903 = n4901 & n6403;
assign n7229 = n7608 | n6404;
assign n1581 = ~(n9315 ^ n4399);
assign n11171 = ~n1916;
assign n8112 = n2942 | n1618;
assign n3036 = ~n6075;
assign n7625 = n1490 | n4904;
assign n4658 = n3461 & n6259;
assign n1878 = n7193 | n9933;
assign n7810 = n12476 | n5184;
assign n9270 = n4488 & n3036;
assign n7673 = ~(n3368 ^ n7576);
assign n8479 = n8108 | n8702;
assign n5349 = ~(n7326 | n3565);
assign n6500 = ~(n10423 ^ n3276);
assign n9555 = n8849 | n5414;
assign n6043 = ~(n2482 ^ n10113);
assign n7758 = n7133 | n12847;
assign n10733 = n10751 ^ n1032;
assign n6649 = n2017 | n7692;
assign n8725 = ~(n11417 ^ n11019);
assign n961 = ~(n10811 | n836);
assign n1705 = n2144 | n12421;
assign n11199 = n6308 & n6925;
assign n4747 = ~(n2516 ^ n5728);
assign n6430 = n4355 | n8933;
assign n74 = n2724 & n6455;
assign n12283 = ~(n10697 ^ n2366);
assign n8898 = ~n1812;
assign n8092 = n7450 & n7867;
assign n7315 = n7409 | n2714;
assign n11244 = ~n13058;
assign n7030 = ~(n3637 ^ n12047);
assign n7224 = n6566 & n155;
assign n3752 = ~n2392;
assign n3502 = n4033 & n1503;
assign n5292 = n3250 & n4117;
assign n9477 = n4946 | n4139;
assign n8633 = ~(n11970 ^ n2502);
assign n7648 = n9049 & n2827;
assign n5572 = n12563 | n10029;
assign n10205 = ~(n28 ^ n253);
assign n2955 = n6624 & n7575;
assign n1413 = n6787 | n4669;
assign n3656 = n3270 | n13143;
assign n10057 = ~n5962;
assign n10552 = ~n6668;
assign n5704 = n1887 | n1043;
assign n2050 = ~(n5798 | n9276);
assign n5643 = ~(n4781 ^ n8633);
assign n9421 = ~n11574;
assign n11363 = n161 | n10179;
assign n4620 = ~n2295;
assign n4705 = ~(n5759 ^ n12038);
assign n2584 = ~(n2125 ^ n10118);
assign n7169 = ~(n11530 | n4472);
assign n9048 = n3545 & n13140;
assign n4219 = n7055 & n6292;
assign n4363 = n994 | n1433;
assign n7808 = ~(n6199 ^ n3147);
assign n1758 = ~(n4531 ^ n6077);
assign n3686 = ~(n12468 | n2202);
assign n9414 = n308 & n4302;
assign n310 = n8392 | n8030;
assign n8919 = n8887 ^ n5270;
assign n6698 = ~(n1549 ^ n12611);
assign n12563 = ~n12306;
assign n2337 = n8335 | n6265;
assign n1377 = ~n10424;
assign n8903 = n12776 & n11603;
assign n13119 = n318 | n10106;
assign n9723 = ~n7659;
assign n10225 = n9112 | n4947;
assign n4045 = n1995 | n1081;
assign n2073 = ~(n9389 ^ n9551);
assign n7950 = ~n9915;
assign n8121 = ~(n9436 ^ n3674);
assign n11970 = ~(n494 ^ n11329);
assign n7838 = ~(n7294 ^ n10111);
assign n2828 = ~(n10424 ^ n13076);
assign n11800 = ~n3838;
assign n5061 = n7523 & n7975;
assign n1186 = ~n8227;
assign n1725 = ~n6409;
assign n12137 = n7372 | n11628;
assign n6908 = ~(n1313 ^ n3667);
assign n5732 = n7529 & n10451;
assign n5160 = n7283 | n7723;
assign n10040 = n3987 & n12362;
assign n3871 = n6975 | n7871;
assign n160 = n9934 | n2675;
assign n9247 = n2715 & n4265;
assign n5024 = n4729 & n3204;
assign n1255 = ~n2202;
assign n7781 = ~(n4337 ^ n10478);
assign n7958 = ~(n12716 ^ n9322);
assign n4302 = ~(n1849 ^ n5594);
assign n10506 = ~(n3741 ^ n9143);
assign n3589 = ~n589;
assign n6094 = ~(n11561 ^ n8578);
assign n1519 = ~(n4356 ^ n10499);
assign n6855 = n8400 | n13148;
assign n930 = ~n12577;
assign n2610 = n9945 | n2418;
assign n9937 = n9892 | n10526;
assign n12030 = n3259 | n80;
assign n9465 = ~n4507;
assign n1045 = ~n12443;
assign n5756 = ~(n10341 ^ n3636);
assign n3516 = ~n3311;
assign n11916 = ~(n3728 | n8537);
assign n8250 = n12055 | n1285;
assign n8763 = n12737 & n5956;
assign n8658 = ~n13184;
assign n2406 = ~n2458;
assign n6543 = ~n12641;
assign n4561 = n7924 & n2528;
assign n4941 = n2412 & n5668;
assign n5303 = n6690 & n12772;
assign n7613 = ~(n2514 ^ n13160);
assign n4738 = n74 | n9278;
assign n12916 = n424 ^ n1698;
assign n2509 = n8008 | n12113;
assign n396 = ~(n9292 ^ n11921);
assign n3055 = ~(n6446 ^ n4178);
assign n52 = n6849 | n12526;
assign n456 = ~(n1546 ^ n2204);
assign n11808 = ~n11324;
assign n8826 = n2648 & n9829;
assign n7192 = n5040 | n6370;
assign n3884 = ~(n1676 | n10083);
assign n7855 = n4595 & n11343;
assign n1515 = n12139 & n11775;
assign n2937 = ~(n4175 ^ n3231);
assign n197 = n10290 | n11668;
assign n5815 = n8093 & n7019;
assign n10600 = ~(n145 | n853);
assign n11265 = ~(n12642 | n3291);
assign n8287 = ~(n4713 ^ n11441);
assign n13178 = n11626 | n2891;
assign n3219 = ~(n11488 | n1982);
assign n3997 = n724 & n11163;
assign n8195 = ~(n7874 ^ n5922);
assign n8484 = ~(n12610 ^ n13067);
assign n367 = ~(n5556 | n13198);
assign n9918 = n1320 | n2671;
assign n5365 = n5423 | n2133;
assign n12058 = n4622 | n11214;
assign n6595 = ~n13060;
assign n2177 = n1883 | n6732;
assign n8560 = n1522 & n3483;
assign n2922 = n6035 | n11146;
assign n747 = n626 | n7887;
assign n2813 = ~(n1256 ^ n1619);
assign n3973 = n2198 & n193;
assign n11712 = n11690 & n12743;
assign n2439 = ~(n1803 ^ n7587);
assign n8901 = n11320 | n6293;
assign n2335 = n2747 & n8762;
assign n3863 = ~(n9371 ^ n8323);
assign n3251 = n9828 & n10804;
assign n5221 = ~(n4968 | n11700);
assign n11603 = ~(n2513 ^ n11578);
assign n13020 = ~(n3878 ^ n7248);
assign n10217 = ~(n5407 ^ n2708);
assign n1144 = n8569;
assign n449 = ~(n3764 | n2888);
assign n12587 = ~(n232 | n3580);
assign n6240 = n683 | n4144;
assign n7148 = ~(n13193 ^ n2642);
assign n12530 = n154 | n9962;
assign n7121 = ~(n6184 ^ n2115);
assign n11986 = ~n12417;
assign n9242 = n1582 & n5706;
assign n9535 = n660 | n1530;
assign n1141 = ~(n880 ^ n2856);
assign n6809 = ~(n11518 ^ n10337);
assign n441 = ~(n12737 ^ n10009);
assign n8699 = n6726 | n206;
assign n7174 = n9094 | n6605;
assign n8921 = ~(n565 ^ n10445);
assign n10362 = n1539 & n12633;
assign n13062 = n1296 | n8702;
assign n3904 = ~(n1461 ^ n2303);
assign n5834 = n2482 & n12289;
assign n1337 = ~n11254;
assign n3080 = ~(n6805 | n7691);
assign n10270 = ~(n1744 | n315);
assign n6984 = ~(n10134 ^ n183);
assign n2329 = ~n7974;
assign n3767 = n11291 | n7530;
assign n1326 = n3473 & n8337;
assign n1287 = ~(n5402 | n5149);
assign n11877 = n10263 | n12695;
assign n12712 = n5365 | n8749;
assign n1538 = ~n12418;
assign n8127 = n5667 | n5242;
assign n2118 = ~n12408;
assign n13143 = ~(n10409 ^ n741);
assign n8047 = n9450 | n6968;
assign n9092 = n2458 & n9669;
assign n9208 = ~(n5702 | n7866);
assign n5697 = ~n13098;
assign n3870 = ~n825;
assign n1741 = ~n10606;
assign n2204 = n7158 | n2059;
assign n8863 = ~n3409;
assign n10004 = n4964 & n11222;
assign n10971 = ~(n12812 ^ n2983);
assign n10191 = n545 & n1849;
assign n5237 = n5118 & n6806;
assign n2120 = ~(n2807 ^ n10355);
assign n11843 = ~(n11673 | n42);
assign n1987 = n7869 & n3606;
assign n3310 = n10871 | n1463;
assign n6178 = ~n11537;
assign n4427 = n4708 & n12550;
assign n394 = n12902 & n1684;
assign n4001 = n433 & n9224;
assign n2665 = ~(n10483 ^ n6782);
assign n7680 = n10143 | n12847;
assign n336 = n93 & n7772;
assign n11439 = n6164 & n413;
assign n12760 = n1030 & n4243;
assign n5366 = n5926 | n10884;
assign n12341 = n11985 & n5435;
assign n13111 = ~(n6179 | n5674);
assign n8292 = n11548 | n9159;
assign n11795 = n6010 | n11746;
assign n5262 = n9646 & n12984;
assign n10663 = ~(n10053 ^ n12087);
assign n8678 = ~(n5114 ^ n3506);
assign n9995 = n6498 | n258;
assign n4648 = n10290 | n6265;
assign n5951 = ~(n5935 ^ n8181);
assign n54 = ~(n5438 ^ n5070);
assign n4903 = n12397 | n5235;
assign n703 = n10990 | n13032;
assign n12215 = ~(n3296 ^ n5458);
assign n13150 = ~(n10163 | n4344);
assign n13121 = n855 & n2047;
assign n11652 = n8940 & n5536;
assign n10384 = ~n9895;
assign n9282 = ~n8139;
assign n5650 = ~n5302;
assign n10515 = ~(n149 | n8152);
assign n10703 = n5270 & n5383;
assign n7144 = n4848 & n4984;
assign n3450 = ~n6700;
assign n4799 = n4114 & n8506;
assign n8907 = ~n9610;
assign n2583 = n12592 & n3085;
assign n9090 = ~(n2630 ^ n2561);
assign n13019 = ~(n10048 | n12842);
assign n7761 = n8183 & n9475;
assign n1917 = n3998 & n4486;
assign n7561 = n4411 | n11135;
assign n969 = ~(n3263 | n12045);
assign n529 = ~(n4264 ^ n6287);
assign n132 = n9567 | n7429;
assign n7074 = ~n469;
assign n4929 = n9553 | n6278;
assign n444 = ~(n11433 ^ n12214);
assign n12490 = ~n9475;
assign n7520 = ~(n6800 | n13236);
assign n2614 = ~n1302;
assign n4976 = n9181 | n5740;
assign n7012 = n5890 | n2133;
assign n3491 = ~(n13094 | n8218);
assign n13040 = n4618 & n1232;
assign n6080 = n6421 & n13088;
assign n4412 = ~n1753;
assign n12788 = n12855 | n9088;
assign n4321 = n2877 | n7903;
assign n4047 = n3342 & n8606;
assign n6488 = ~n3076;
assign n10990 = ~(n2431 | n10178);
assign n972 = n12043 & n1005;
assign n8244 = n189 | n11929;
assign n5210 = n1331 | n4455;
assign n5211 = ~(n4021 ^ n6863);
assign n3172 = n11582 | n3801;
assign n10651 = n233 & n11539;
assign n4011 = ~(n7277 ^ n5378);
assign n4942 = n5377 | n12491;
assign n6288 = ~(n1092 ^ n1479);
assign n4601 = ~(n10802 ^ n10684);
assign n1933 = n8532 | n12273;
assign n185 = ~(n6264 | n11458);
assign n12111 = ~(n2063 | n12586);
assign n4784 = n2130 | n8465;
assign n2802 = n6768 | n9195;
assign n3444 = n7228 | n1383;
assign n8364 = ~(n6765 | n10744);
assign n378 = ~(n12374 ^ n12322);
assign n7399 = ~(n11763 ^ n8021);
assign n7388 = ~n6417;
assign n10417 = n10708 & n9588;
assign n9606 = ~n4748;
assign n8513 = ~(n6902 | n9158);
assign n7817 = ~n720;
assign n6335 = n5897 | n159;
assign n1082 = ~n12564;
assign n5392 = ~(n2334 | n3468);
assign n4139 = ~n5753;
assign n6785 = ~(n3951 ^ n5896);
assign n12319 = ~(n4369 ^ n9805);
assign n9992 = ~n1521;
assign n6846 = ~n12482;
assign n3284 = n10761 | n12388;
assign n3890 = ~n9620;
assign n10308 = ~(n12230 | n4204);
assign n6146 = n1359 | n2438;
assign n9792 = ~(n2011 ^ n9483);
assign n4386 = ~(n6097 | n11416);
assign n11454 = ~(n10500 ^ n6542);
assign n505 = n5107 | n1571;
assign n2631 = n7011 & n7117;
assign n10916 = ~n3395;
assign n12478 = ~n4318;
assign n7240 = n10948 & n9137;
assign n9081 = ~(n6242 ^ n10276);
assign n7075 = ~n6168;
assign n5212 = n3159 | n9507;
assign n9892 = n12748 | n12188;
assign n3750 = n6172 | n7610;
assign n11122 = ~n7720;
assign n10073 = ~(n5299 ^ n13072);
assign n9115 = n3435 & n11697;
assign n13139 = n8835 & n8521;
assign n978 = n652 | n5076;
assign n8936 = ~n28;
assign n363 = ~(n1675 ^ n4573);
assign n13011 = n6590 | n1985;
assign n7547 = n6509 | n9590;
assign n9199 = n4736 & n5256;
assign n9240 = n9489 | n5242;
assign n4057 = ~(n4840 | n5887);
assign n10172 = n4495 | n8499;
assign n11583 = n8026 & n9623;
assign n9818 = ~(n11599 ^ n8226);
assign n13052 = ~n5965;
assign n2098 = n7418 | n11744;
assign n6630 = ~n497;
assign n8983 = n4164 & n5441;
assign n5974 = ~n9212;
assign n10155 = n12552 | n8030;
assign n4883 = n5370 | n5983;
assign n5993 = n8646 | n177;
assign n9910 = ~n7671;
assign n7452 = n6533 & n427;
assign n5522 = ~n7919;
assign n5358 = ~(n6254 ^ n4367);
assign n3693 = ~(n3770 ^ n10758);
assign n11895 = ~(n9578 ^ n213);
assign n10146 = n10388 & n10700;
assign n3063 = ~n5576;
assign n3987 = n11596 & n11721;
assign n5346 = n6943 & n3637;
assign n8660 = n5776 & n924;
assign n1614 = ~(n2379 | n690);
assign n7516 = ~(n3138 ^ n7058);
assign n7872 = ~n11109;
assign n10882 = ~n4528;
assign n3579 = n3564 | n10871;
assign n10288 = n6194 & n2721;
assign n3984 = n2889 | n10319;
assign n2663 = n9695 | n8305;
assign n12859 = ~n12670;
assign n7885 = n11878 & n7390;
assign n3295 = ~(n5742 | n12170);
assign n3357 = ~(n7751 ^ n750);
assign n10446 = n9017 | n8534;
assign n1072 = n8131 | n1985;
assign n4189 = n11033 | n2126;
assign n4714 = ~n2856;
assign n6036 = n8248 & n7155;
assign n2374 = ~(n7496 ^ n9981);
assign n844 = n1715 | n8313;
assign n9272 = ~n10063;
assign n1138 = n10142 & n13058;
assign n1051 = ~n7113;
assign n4358 = n5592 & n4607;
assign n12037 = n10410 | n4073;
assign n6251 = ~(n3145 ^ n1583);
assign n9014 = n10943 & n6511;
assign n8396 = n6129 | n4947;
assign n2873 = ~(n5926 ^ n10884);
assign n3257 = ~n194;
assign n4808 = ~n4335;
assign n812 = ~n3431;
assign n9585 = n7772 & n7411;
assign n12709 = n6605 & n9094;
assign n12775 = n10421 | n12388;
assign n87 = ~(n2658 ^ n10396);
assign n2674 = ~n5998;
assign n6577 = n9691 & n217;
assign n1003 = n5097 & n8002;
assign n4876 = n3301 | n1415;
assign n12313 = ~(n11560 ^ n10646);
assign n3849 = ~(n4252 ^ n12666);
assign n10794 = ~n13087;
assign n8444 = n5720 | n8502;
assign n10189 = n6148 | n11494;
assign n3184 = n2528 | n7924;
assign n8760 = n11123;
assign n5654 = ~n8308;
assign n5032 = ~(n589 ^ n7217);
assign n6480 = n5266 | n3380;
assign n8728 = ~n1495;
assign n7655 = n6480 & n6835;
assign n12990 = n3225 | n7530;
assign n1409 = ~(n4760 ^ n12516);
assign n9285 = n8389 & n7192;
assign n3198 = ~(n4042 ^ n2271);
assign n7124 = ~(n2458 | n8230);
assign n7473 = ~n8357;
assign n8184 = ~(n6961 ^ n1527);
assign n11410 = ~(n5353 ^ n4456);
assign n5514 = n7234 | n12718;
assign n9312 = ~(n9883 ^ n8404);
assign n13154 = ~n287;
assign n11298 = ~(n12816 ^ n8037);
assign n2149 = n10908 & n6937;
assign n11963 = n3503 & n11070;
assign n11529 = ~(n3593 ^ n1455);
assign n4881 = n11235 & n6113;
assign n8154 = n10158 | n1583;
assign n8509 = n6119 & n4432;
assign n9932 = ~(n9407 ^ n1933);
assign n12806 = n7532 | n4724;
assign n9853 = n6215 | n4453;
assign n5150 = n8030 | n4640;
assign n842 = n1163 | n3920;
assign n2525 = ~(n8996 ^ n6592);
assign n8997 = n10014 & n8235;
assign n8766 = n12469 | n8534;
assign n8610 = n3730 | n12302;
assign n11082 = ~(n10850 | n1486);
assign n3820 = n3956 & n13123;
assign n1521 = ~n2690;
assign n12232 = ~(n8074 ^ n9615);
assign n12909 = n4771 & n12332;
assign n11026 = n3719 & n9958;
assign n7534 = ~(n4842 ^ n858);
assign n2595 = n2220 ^ n2198;
assign n11204 = n4187 & n10512;
assign n289 = n7927 & n7456;
assign n11176 = n12227 & n11286;
assign n7518 = n8583 | n11524;
assign n11924 = n6112 | n12623;
assign n3137 = ~(n3283 ^ n4281);
assign n9132 = ~n7115;
assign n8018 = ~(n8297 | n13055);
assign n5516 = n1939 | n8116;
assign n1628 = n7516 & n1236;
assign n615 = n6875 | n12847;
assign n8388 = n3344 | n8609;
assign n12865 = ~(n6424 ^ n6884);
assign n5135 = n6175 | n1192;
assign n9857 = ~(n3255 ^ n12672);
assign n1959 = n1215 | n8511;
assign n3243 = ~n11396;
assign n11399 = n3636 | n10341;
assign n11567 = n12990 ^ n1024;
assign n3796 = ~(n4334 ^ n12958);
assign n521 = ~n11873;
assign n963 = ~n6611;
assign n3827 = n12512 | n10249;
assign n10450 = ~(n2282 ^ n5940);
assign n1213 = n12604 | n2449;
assign n8608 = ~(n7199 ^ n10924);
assign n6944 = ~n834;
assign n5431 = ~(n9993 ^ n6275);
assign n413 = ~n3623;
assign n6524 = ~n7417;
assign n1339 = ~(n810 ^ n8138);
assign n61 = ~n11091;
assign n1537 = ~(n12530 ^ n797);
assign n9990 = ~(n6614 ^ n6996);
assign n5200 = ~n12589;
assign n3634 = ~n8860;
assign n7200 = ~(n82 | n2481);
assign n12236 = n7234 | n206;
assign n8426 = n11729 | n5797;
assign n9532 = ~(n10704 ^ n778);
assign n11034 = ~(n9826 | n8261);
assign n9055 = ~n11089;
assign n5648 = ~(n6534 | n3474);
assign n4193 = n7322 & n730;
assign n2872 = ~n9531;
assign n4198 = ~n3769;
assign n3624 = ~(n8311 ^ n6836);
assign n4749 = n8665 | n12655;
assign n12333 = n11157 | n8030;
assign n2797 = ~(n973 ^ n2281);
assign n59 = n3531 | n4230;
assign n9719 = ~(n8429 ^ n11443);
assign n11316 = n10215 & n5929;
assign n2899 = ~n817;
assign n5709 = ~n11974;
assign n9567 = n2129 | n4373;
assign n4371 = ~n7128;
assign n3422 = n1496 & n5844;
assign n10301 = n12166 | n1197;
assign n11980 = n10931 & n1903;
assign n3557 = n8362 | n6181;
assign n2494 = ~(n8004 ^ n2981);
assign n4906 = n3507 & n5717;
assign n53 = ~n761;
assign n2299 = n7129 | n2617;
assign n3303 = n10770 & n287;
assign n10190 = n333 | n12967;
assign n8529 = ~n5969;
assign n4130 = ~(n5934 ^ n12002);
assign n11188 = n10849 & n7784;
assign n9059 = n5947 | n12695;
assign n1410 = n10642 & n7720;
assign n8268 = n765;
assign n6354 = n7608 | n206;
assign n2230 = ~(n12141 ^ n12407);
assign n6362 = n4349 ^ n2419;
assign n3250 = ~(n1121 ^ n12125);
assign n1767 = ~n12950;
assign n9235 = ~(n12237 | n2512);
assign n6264 = ~n2754;
assign n4836 = n7719 | n275;
assign n6325 = n13201 & n3085;
assign n6842 = ~(n4684 | n12927);
assign n8653 = n11103 | n5388;
assign n6207 = ~(n8773 | n4345);
assign n745 = n5569 | n7221;
assign n6729 = n3517 & n3571;
assign n7703 = n12416 | n9159;
assign n13115 = n11450 | n4757;
assign n5865 = ~n11835;
assign n4951 = ~(n5793 ^ n1990);
assign n9772 = ~n1342;
assign n2324 = n10565 & n5585;
assign n810 = n12671 | n10430;
assign n7488 = ~(n11883 | n9598);
assign n2056 = ~n5451;
assign n11055 = n379 | n2816;
assign n928 = n4052 & n109;
assign n1563 = ~(n4509 ^ n875);
assign n7546 = n6680 | n2890;
assign n1593 = n8011 | n2772;
assign n7034 = ~(n94 ^ n6935);
assign n10518 = ~(n10671 ^ n1317);
assign n8866 = n13013 | n0;
assign n7874 = n3826 | n10106;
assign n1073 = ~n7749;
assign n11219 = n5113 & n9133;
assign n5757 = ~(n1077 ^ n11598);
assign n8979 = n2484 | n10552;
assign n9053 = n2391 | n2531;
assign n6971 = n1107 & n10571;
assign n12539 = n8153 & n11275;
assign n11668 = n9280;
assign n238 = n1206 | n11490;
assign n1879 = n8665 | n1720;
assign n6945 = n3796 | n12724;
assign n2812 = n9098 | n6002;
assign n7724 = ~(n1338 ^ n4471);
assign n173 = ~n10906;
assign n10039 = ~n7144;
assign n4078 = n12348 & n5065;
assign n4533 = n10078 & n11040;
assign n2350 = ~n10301;
assign n4829 = n12951 | n7988;
assign n4885 = n9882 | n11300;
assign n12183 = ~n6242;
assign n4354 = n3982 & n752;
assign n7072 = ~n4399;
assign n148 = ~(n10377 ^ n3608);
assign n10350 = n5516 & n6976;
assign n5097 = ~n7605;
assign n2827 = n767 & n3832;
assign n1806 = ~(n10455 ^ n1147);
assign n5487 = ~(n4558 ^ n1811);
assign n5656 = n5530 & n1068;
assign n10612 = ~(n5391 | n9231);
assign n1018 = ~n9313;
assign n5003 = ~(n953 ^ n8746);
assign n12692 = ~(n3607 ^ n2525);
assign n1749 = n6913 | n9650;
assign n208 = n11980 | n8375;
assign n490 = ~n2869;
assign n7106 = n8766 | n2647;
assign n9105 = ~(n1141 ^ n10521);
assign n7515 = n3613 ^ n12527;
assign n6112 = ~n8332;
assign n873 = n4173 & n7275;
assign n4817 = ~(n3502 | n3857);
assign n4467 = n3208 | n7221;
assign n2126 = n4659 & n3151;
assign n12792 = n3818 | n12040;
assign n9611 = n2008 & n12318;
assign n11284 = ~n11222;
assign n3899 = ~(n4568 ^ n2693);
assign n2887 = n1416 | n4967;
assign n7519 = n4478 | n1599;
assign n2424 = n6769 | n7935;
assign n3619 = ~n12661;
assign n10277 = n2424 | n6729;
assign n9558 = ~n12750;
assign n9173 = ~(n9200 | n5471);
assign n6719 = n12607 | n8041;
assign n11161 = ~(n7375 | n10819);
assign n9946 = ~(n1871 ^ n10868);
assign n2644 = n6488 | n6265;
assign n1022 = n10318 ^ n11196;
assign n1679 = n10966 | n9075;
assign n9042 = n9575 | n1500;
assign n657 = ~n2841;
assign n1 = n8430 & n10255;
assign n4177 = ~(n6292 ^ n10418);
assign n8635 = ~(n12815 ^ n3799);
assign n2375 = n1759 & n11382;
assign n4798 = n9239 & n487;
assign n11112 = ~(n2144 ^ n11001);
assign n12210 = n6129 | n11144;
assign n7016 = n3444 & n7652;
assign n3058 = ~n2482;
assign n9662 = n8992 | n541;
assign n6154 = ~(n1540 ^ n6221);
assign n5133 = n5842 | n6033;
assign n3869 = n12465 | n13086;
assign n11090 = ~(n12791 ^ n6666);
assign n3872 = ~(n570 | n3366);
assign n6950 = n103 & n854;
assign n5186 = n7622 & n8815;
assign n10674 = n4844 | n9075;
assign n5136 = ~n7214;
assign n12504 = n6476 | n8663;
assign n11681 = n9417 & n256;
assign n11036 = ~(n8109 ^ n3515);
assign n6261 = ~(n2203 ^ n7623);
assign n3306 = ~(n11775 ^ n665);
assign n10938 = n227 | n6635;
assign n12824 = n8175 & n7616;
assign n2829 = n5786 ^ n1687;
assign n10778 = n5217 & n12011;
assign n11790 = ~n12134;
assign n5599 = ~(n889 | n7897);
assign n7230 = n4890 | n4936;
assign n11825 = n7210 | n12499;
assign n10825 = ~(n6650 ^ n3390);
assign n9814 = n11187 | n8517;
assign n7550 = ~(n4260 ^ n2093);
assign n6881 = ~n12539;
assign n607 = ~(n4708 ^ n10644);
assign n11443 = n6267 & n3400;
assign n11119 = n8105 | n13204;
assign n5763 = ~(n5015 ^ n11380);
assign n8719 = ~n3828;
assign n2394 = ~n9536;
assign n1777 = n2622 | n8268;
assign n2452 = ~n3409;
assign n11968 = n4791 & n11517;
assign n11997 = ~(n13134 ^ n3935);
assign n10603 = n3225 | n2675;
assign n3728 = n11114 | n11522;
assign n9652 = ~(n2294 ^ n13017);
assign n12211 = ~n3756;
assign n5463 = ~(n7192 ^ n8389);
assign n277 = ~(n10323 ^ n1955);
assign n7773 = n10462 | n4230;
assign n3648 = n12264 & n12355;
assign n8913 = ~n2354;
assign n2490 = n12266 & n11625;
assign n4027 = ~(n369 ^ n5339);
assign n4387 = n12987 ^ n3141;
assign n7925 = ~n443;
assign n7533 = ~n9062;
assign n4624 = n9132 & n770;
assign n95 = n2416 | n8534;
assign n3626 = ~(n11098 ^ n4280);
assign n1112 = ~(n13211 ^ n8725);
assign n1117 = ~n2591;
assign n8054 = ~(n5370 ^ n5983);
assign n11445 = ~(n8836 ^ n6953);
assign n2567 = ~(n9654 ^ n2866);
assign n7511 = ~(n3807 ^ n5624);
assign n6735 = n6028 | n7723;
assign n1615 = ~(n2699 ^ n8946);
assign n5680 = ~(n4400 | n12285);
assign n11221 = ~(n2237 ^ n9081);
assign n8511 = ~n3845;
assign n7336 = n879 & n12413;
assign n9976 = n6354 | n8707;
assign n3141 = n8259 & n12511;
assign n12611 = ~(n400 ^ n8596);
assign n10216 = ~(n5133 ^ n10020);
assign n2416 = ~n9570;
assign n5734 = ~(n20 | n732);
assign n3065 = ~(n10191 | n9414);
assign n12324 = ~n7720;
assign n9543 = n684 & n8617;
assign n8884 = n2640 ^ n9983;
assign n8851 = ~(n10600 ^ n3897);
assign n1847 = ~n4874;
assign n4150 = ~(n5140 ^ n6791);
assign n12744 = n971 | n3981;
assign n12748 = ~n12651;
assign n12188 = n9257;
assign n7739 = n3127 | n3949;
assign n2633 = n349 & n11283;
assign n6384 = ~(n10602 ^ n2771);
assign n11149 = n3544 ^ n10553;
assign n3616 = ~n2341;
assign n4043 = ~(n10592 ^ n12502);
assign n11962 = ~(n8883 ^ n9479);
assign n5274 = n4305 & n407;
assign n4294 = ~n12990;
assign n868 = ~n11663;
assign n5456 = n6048 | n5919;
assign n12316 = ~n10142;
assign n10089 = ~(n12339 | n8342);
assign n12425 = ~n1700;
assign n119 = ~n3815;
assign n5121 = n10908 & n5065;
assign n1269 = ~n2388;
assign n7803 = ~(n7613 | n12303);
assign n7759 = ~(n4858 ^ n6896);
assign n10817 = ~(n6694 ^ n11017);
assign n4423 = ~(n5424 ^ n3838);
assign n7187 = n7263 | n12492;
assign n7439 = ~(n1048 ^ n378);
assign n2330 = ~n8267;
assign n1569 = n13147 & n2602;
assign n11931 = ~(n3533 ^ n4754);
assign n8043 = ~(n11386 ^ n1497);
assign n12443 = n2273 & n1598;
assign n8130 = ~(n1471 | n13033);
assign n6518 = n5626 | n12291;
assign n3581 = n9897 & n897;
assign n12208 = ~(n6521 ^ n7565);
assign n7134 = ~(n4689 | n4705);
assign n1820 = ~n8290;
assign n11613 = n1965 & n11784;
assign n10120 = ~n12477;
assign n7607 = n10761 | n2675;
assign n2848 = ~n11111;
assign n12024 = ~(n8432 ^ n8045);
assign n1967 = ~n9481;
assign n2027 = n9868 | n1043;
assign n12139 = ~(n12011 ^ n4897);
assign n9794 = ~(n8387 ^ n10333);
assign n10508 = ~n7384;
assign n7831 = n6880 & n5072;
assign n11663 = n12478 & n13139;
assign n8816 = n36 | n1703;
assign n6248 = n372 & n12572;
assign n7049 = ~n10606;
assign n6923 = n7787 | n6878;
assign n10269 = n12380 & n5082;
assign n1751 = n6735 | n9791;
assign n4383 = ~(n897 ^ n4126);
assign n3328 = n10771 & n1878;
assign n5469 = ~n9847;
assign n9436 = ~n11012;
assign n4132 = ~n2339;
assign n11938 = ~(n8996 | n3607);
assign n12224 = ~n7659;
assign n12254 = ~n2339;
assign n2956 = ~n1344;
assign n3966 = n1354 | n7723;
assign n7822 = ~(n13145 ^ n319);
assign n5631 = n5236 & n9954;
assign n10742 = n8598 | n4640;
assign n3992 = n9113 | n10179;
assign n2959 = n6241 & n1846;
assign n5368 = n4379 & n2897;
assign n10127 = ~n10876;
assign n8492 = ~n6209;
assign n5560 = ~(n2766 ^ n7566);
assign n11886 = ~(n5161 ^ n6116);
assign n3162 = ~(n6780 | n8855);
assign n7544 = ~n11372;
assign n11530 = n4620 | n2675;
assign n10520 = n11392 | n9760;
assign n12733 = ~(n8057 | n4415);
assign n8399 = n8954 ^ n11294;
assign n9113 = ~n10874;
assign n10100 = n2563 & n1509;
assign n7508 = n7438 | n3732;
assign n11288 = n7191 | n1144;
assign n12727 = ~(n12333 | n12640);
assign n10462 = ~n1916;
assign n1673 = n8426 | n11754;
assign n7614 = ~n9052;
assign n8007 = ~(n2804 ^ n10678);
assign n1143 = n10425 & n10380;
assign n9943 = ~(n2618 ^ n11179);
assign n2695 = n10493 & n9927;
assign n5980 = n11864 | n7961;
assign n12000 = ~n9591;
assign n9748 = n2759 | n3653;
assign n12999 = n5296 | n2277;
assign n7674 = n6854 | n8268;
assign n11398 = ~n13212;
assign n1838 = n10784 | n10576;
assign n7853 = ~(n8682 ^ n9351);
assign n1721 = ~(n9579 ^ n7024);
assign n11829 = n8091 | n10932;
assign n793 = ~(n6965 | n1626);
assign n4859 = n1150 | n6005;
assign n11418 = ~n10416;
assign n9753 = ~(n8981 ^ n598);
assign n4257 = ~n2012;
assign n9689 = ~(n4233 | n5229);
assign n5844 = n1335 | n3890;
assign n3436 = ~(n7321 ^ n11993);
assign n10214 = n11074 & n8753;
assign n5413 = n9403 & n4578;
assign n1881 = ~n3910;
assign n8264 = n1618 | n12273;
assign n8877 = ~n1291;
assign n245 = n761 & n5548;
assign n10899 = ~(n5952 | n205);
assign n9646 = n10501 | n4373;
assign n517 = n5384 & n6118;
assign n2990 = ~(n12928 | n2247);
assign n2013 = ~n5952;
assign n10536 = n10637 | n9234;
assign n6724 = ~n12408;
assign n6202 = n8904 | n10029;
assign n1817 = n4038 | n9984;
assign n835 = ~(n344 ^ n6639);
assign n8933 = ~(n2910 | n1430);
assign n2839 = ~(n12020 ^ n964);
assign n7253 = n2097 | n2917;
assign n7915 = ~(n8805 ^ n11623);
assign n12532 = n6369 & n13167;
assign n764 = n8228 & n5920;
assign n12950 = ~(n1125 ^ n12488);
assign n7730 = ~n5167;
assign n3864 = ~(n5294 | n8289);
assign n4167 = n9113 | n177;
assign n3398 = n8877 & n11133;
assign n7268 = ~(n8923 ^ n7479);
assign n973 = n13026 | n177;
assign n7464 = n9303 & n11029;
assign n944 = n9371 | n12016;
assign n6550 = n1586 & n2253;
assign n10437 = ~n1302;
assign n4485 = n1529 | n604;
assign n5418 = ~(n9221 ^ n12344);
assign n11716 = ~(n6952 ^ n8149);
assign n12541 = ~(n7349 | n12447);
assign n6017 = ~(n12821 ^ n9452);
assign n12531 = ~(n10088 ^ n12494);
assign n1183 = n6168 & n12853;
assign n9744 = n13041 & n3661;
assign n7953 = n1261 | n177;
assign n13142 = ~(n9588 ^ n10708);
assign n190 = n9983 | n8246;
assign n1690 = ~(n11837 | n913);
assign n5112 = n6100 & n10389;
assign n13036 = ~n9187;
assign n4449 = ~(n3923 ^ n261);
assign n2082 = n7990 & n3609;
assign n6696 = ~(n4988 ^ n9686);
assign n12198 = n1947 | n8018;
assign n9342 = n1334 | n7926;
assign n128 = ~n13011;
assign n881 = ~n10951;
assign n8401 = n1727 | n8083;
assign n717 = ~(n475 ^ n10012);
assign n9324 = n8948 & n8786;
assign n11234 = ~(n10186 | n10206);
assign n888 = n8295 & n6694;
assign n1353 = ~n4748;
assign n5901 = ~(n3973 ^ n11389);
assign n4570 = ~(n1426 ^ n3751);
assign n11352 = ~n7411;
assign n12446 = n1068 | n5530;
assign n9008 = ~n7164;
assign n1835 = ~(n175 ^ n9377);
assign n5253 = ~(n625 | n9390);
assign n3461 = n10676 & n1091;
assign n6704 = ~(n633 ^ n1000);
assign n5744 = n9739 | n10106;
assign n7219 = n11256 | n9657;
assign n12394 = n1315 & n10174;
assign n5023 = ~(n3179 ^ n11465);
assign n2647 = ~(n8428 ^ n11341);
assign n6730 = ~(n6498 ^ n4246);
assign n1507 = n734 | n10956;
assign n8731 = ~(n962 ^ n11405);
assign n9389 = n11007 | n2675;
assign n11556 = ~(n9823 ^ n2704);
assign n5420 = ~n3181;
assign n11338 = n21 & n2740;
assign n7777 = n2217 | n10871;
assign n9039 = n6068 ^ n5834;
assign n10432 = n3161 & n3249;
assign n7627 = ~(n9678 | n5171);
assign n10731 = n992 | n7239;
assign n8012 = ~n3283;
assign n3816 = ~n5062;
assign n8481 = ~n3939;
assign n5702 = ~(n7096 ^ n7458);
assign n2963 = n9226 | n9521;
assign n7972 = n10919 | n4765;
assign n1449 = ~(n12894 ^ n6459);
assign n10968 = ~(n11710 ^ n11702);
assign n8703 = n7900 | n10106;
assign n2430 = ~n10458;
assign n11056 = n5400 & n4047;
assign n3959 = ~(n7542 ^ n3710);
assign n9205 = n11965 | n4844;
assign n9619 = n4382 & n11109;
assign n2106 = n3327 | n926;
assign n7672 = ~n12579;
assign n10985 = n9135 & n12548;
assign n5770 = n3311 & n6085;
assign n9524 = ~(n4851 | n2998);
assign n9153 = n4213 | n4255;
assign n10119 = ~(n6268 ^ n4358);
assign n8400 = ~n11109;
assign n8 = n8645 | n8563;
assign n5378 = n11430 & n7519;
assign n2364 = ~(n8638 ^ n10679);
assign n5978 = n818 & n6563;
assign n10621 = ~(n12851 ^ n13112);
assign n2062 = n4198 | n4373;
assign n8723 = ~n105;
assign n6638 = ~n7374;
assign n8433 = n325 & n3739;
assign n2385 = ~n7802;
assign n13231 = ~(n4785 ^ n4120);
assign n9318 = n6841 | n8129;
assign n3372 = n4485 & n5936;
assign n7604 = ~(n3032 ^ n847);
assign n11169 = n9707 & n8888;
assign n8540 = ~n10787;
assign n6148 = ~(n11742 ^ n3098);
assign n8833 = n3724 | n7959;
assign n6526 = n3395 ^ n11402;
assign n2944 = n11592 & n4491;
assign n3694 = ~(n6176 ^ n13062);
assign n9617 = n7069 | n1694;
assign n2897 = n12758 | n5797;
assign n5842 = ~n951;
assign n4545 = ~(n12897 | n5133);
assign n9388 = ~(n5323 | n4094);
assign n9124 = n8082 | n1026;
assign n10556 = ~(n29 ^ n7029);
assign n7345 = ~(n10762 ^ n363);
assign n6462 = n11702 & n11710;
assign n10744 = ~(n4232 ^ n5137);
assign n4983 = ~(n2951 | n4369);
assign n11785 = n2465 & n1868;
assign n5875 = ~n5920;
assign n5171 = n10727 & n1967;
assign n2883 = n2068 & n12284;
assign n8984 = n11102 | n2280;
assign n1055 = ~n2791;
assign n3238 = ~(n6892 | n9952);
assign n13219 = ~(n2370 ^ n13161);
assign n6832 = ~(n5627 ^ n9009);
assign n4398 = ~n7059;
assign n4797 = ~(n6352 ^ n9616);
assign n9508 = ~(n12988 ^ n2012);
assign n4482 = n3209 & n8760;
assign n1412 = ~(n3666 ^ n10218);
assign n11976 = ~(n12097 ^ n1375);
assign n7073 = ~n3199;
assign n9467 = ~(n4602 ^ n11487);
assign n8119 = ~(n402 ^ n12679);
assign n813 = ~n9528;
assign n8326 = n7319 & n12764;
assign n5474 = n5993 | n1298;
assign n6535 = ~(n2088 ^ n11731);
assign n6929 = n7730 | n3825;
assign n8675 = n6522 ^ n11840;
assign n4640 = n12128;
assign n9061 = n525 & n10753;
assign n1092 = ~(n7363 ^ n11216);
assign n9326 = n2046 | n12637;
assign n12784 = n5823 & n5381;
assign n11666 = n5522 & n11056;
assign n733 = ~(n8424 ^ n2225);
assign n2597 = ~(n12590 ^ n4410);
assign n6378 = n4983 | n553;
assign n1821 = n8950 | n12695;
assign n1366 = ~n10869;
assign n7569 = n6749 | n7076;
assign n5187 = n12458 | n4303;
assign n9941 = ~(n10312 ^ n4353);
assign n1711 = n1158 | n1713;
assign n5090 = n9913 | n11868;
assign n12826 = ~(n7442 | n12464);
assign n12061 = ~(n7694 ^ n9438);
assign n4827 = n2462 | n10319;
assign n5460 = ~n3769;
assign n2607 = n294 | n11164;
assign n11084 = n3527;
assign n1134 = ~n2619;
assign n8878 = n10332 | n1344;
assign n671 = n3957 | n11273;
assign n3213 = n9383 | n3981;
assign n13233 = ~(n11973 | n12163);
assign n3345 = n2723 | n4209;
assign n7275 = n10999 | n10342;
assign n9500 = ~(n4403 | n1828);
assign n8259 = ~n2966;
assign n4565 = n10920 & n5497;
assign n7172 = ~(n8606 ^ n3342);
assign n6795 = n6136 & n8022;
assign n10829 = ~(n2995 ^ n2840);
assign n8800 = ~n5722;
assign n3116 = ~n2647;
assign n7532 = ~n497;
assign n5849 = ~(n13070 | n6840);
assign n1997 = n7770 | n8066;
assign n9020 = n10149 | n9413;
assign n5242 = n1750;
assign n7468 = n719 | n290;
assign n9773 = n1912 & n13060;
assign n2704 = ~(n10766 ^ n7287);
assign n5364 = ~(n10390 ^ n12034);
assign n7784 = ~n13223;
assign n6963 = ~(n5800 | n1624);
assign n3571 = n9162 | n12328;
assign n5533 = ~n3043;
assign n2135 = ~n1982;
assign n2380 = n5465 | n6861;
assign n7191 = ~n12651;
assign n11626 = n8584 & n4814;
assign n10769 = n8731 ^ n9437;
assign n7107 = ~(n8457 ^ n6903);
assign n13085 = n2789 | n8029;
assign n3615 = n12933 & n3526;
assign n3118 = ~n12217;
assign n10170 = n12202 | n2042;
assign n6457 = n6614 | n6996;
assign n2849 = ~n10395;
assign n10721 = ~(n4266 ^ n483);
assign n7927 = n11407 | n4787;
assign n5943 = n121 | n9118;
assign n9371 = ~(n454 ^ n1179);
assign n12112 = n63 | n479;
assign n4849 = ~(n1508 ^ n4955);
assign n4400 = n12295 | n10319;
assign n7943 = ~(n9498 ^ n6217);
assign n4987 = n8680 & n222;
assign n2822 = ~n11809;
assign n12559 = ~(n8497 ^ n10634);
assign n5280 = n4042 & n1646;
assign n2886 = n10550 | n6258;
assign n12817 = n9174 & n9250;
assign n10944 = ~n10850;
assign n10530 = n10357 | n409;
assign n11942 = ~n3014;
assign n2579 = ~n12429;
assign n3079 = n8378 & n12080;
assign n7355 = n1320 | n9223;
assign n4692 = n4465 | n8534;
assign n5520 = ~n5758;
assign n418 = ~n12622;
assign n4845 = ~(n914 ^ n6840);
assign n5938 = n1602 ^ n1612;
assign n10929 = ~n9846;
assign n3893 = ~(n12199 ^ n13004);
assign n293 = n2743 & n1620;
assign n5967 = n3006 & n5729;
assign n8458 = ~n12614;
assign n3261 = ~(n6016 ^ n8782);
assign n4391 = n10877 | n4936;
assign n1893 = ~n2882;
assign n2413 = n4171 | n10516;
assign n12827 = ~(n2177 ^ n7571);
assign n12428 = n5420 & n10980;
assign n11743 = n2409 & n12026;
assign n3429 = ~n13188;
assign n4924 = ~(n10745 | n5457);
assign n6222 = ~(n5016 ^ n1238);
assign n12852 = ~(n4978 ^ n5236);
assign n9707 = n3311 & n13058;
assign n3621 = n6629 | n12188;
assign n3150 = ~(n4934 ^ n23);
assign n3857 = ~(n1060 | n5860);
assign n4256 = ~n1836;
assign n1850 = n5009 & n7632;
assign n10696 = ~n411;
assign n8311 = ~(n6744 ^ n5263);
assign n2045 = ~n10751;
assign n3627 = n11449 | n12847;
assign n7481 = ~n4708;
assign n9474 = n7068 | n2544;
assign n5083 = ~(n7418 ^ n3015);
assign n12603 = ~(n3695 ^ n4774);
assign n6805 = n10045 | n2675;
assign n9378 = ~n12850;
assign n3934 = ~(n7368 | n11916);
assign n6883 = ~n10606;
assign n1191 = ~n1231;
assign n5794 = ~(n12479 ^ n2655);
assign n7876 = n9112 | n2671;
assign n5407 = n4366 | n2970;
assign n11991 = ~(n5207 ^ n1708);
assign n5040 = ~n6826;
assign n5521 = ~n11030;
assign n1791 = n2940 | n11756;
assign n4489 = n10798 | n6404;
assign n7209 = ~(n8517 ^ n6324);
assign n6717 = n10137 | n8268;
assign n1678 = n4701 & n10507;
assign n7825 = ~n9093;
assign n10660 = n10266 | n1695;
assign n13205 = ~(n11716 ^ n873);
assign n9851 = ~(n6001 | n10866);
assign n3156 = n5163 | n3981;
assign n7060 = n8659 & n2153;
assign n11165 = ~n5311;
assign n2107 = n2296 | n2387;
assign n1780 = ~(n4417 ^ n12156);
assign n9347 = n11509 & n1254;
assign n7653 = ~(n1169 ^ n10401);
assign n12161 = n12109 | n206;
assign n7567 = ~n11416;
assign n9759 = ~(n13104 | n8566);
assign n12546 = ~(n8914 ^ n12231);
assign n7245 = ~(n9347 | n13030);
assign n11715 = ~(n649 ^ n5691);
assign n11002 = ~n9401;
assign n9257 = ~n7772;
assign n9390 = n11365 & n6531;
assign n1627 = n4583 & n2925;
assign n225 = ~(n11026 | n661);
assign n13204 = n2613 & n12233;
assign n5567 = ~(n5872 | n1170);
assign n12336 = n9794 | n9681;
assign n8331 = n8875 & n8491;
assign n12975 = n5206 & n9789;
assign n6166 = ~n11030;
assign n9236 = n4278 ^ n1879;
assign n12415 = n2479 & n8292;
assign n10429 = n2487 | n9075;
assign n12270 = n6220 | n8225;
assign n4841 = ~n9824;
assign n8200 = n6231 | n5797;
assign n3424 = n109 | n4052;
assign n475 = n1893 | n206;
assign n9670 = n98 | n10286;
assign n9601 = ~n4423;
assign n1800 = n8837 | n5100;
assign n167 = n9330 & n11357;
assign n720 = n785 | n4373;
assign n3022 = n10412 | n5262;
assign n6053 = ~(n13024 | n6887);
assign n7423 = ~(n10546 ^ n2277);
assign n9019 = ~n1916;
assign n6172 = n11781 | n8505;
assign n10792 = ~n6409;
assign n2125 = ~(n819 | n2324);
assign n11212 = ~n7974;
assign n12829 = n10830 | n7530;
assign n82 = n8645 | n3981;
assign n2611 = n8576 & n8825;
assign n2444 = n1571 | n11668;
assign n11558 = n11400 | n111;
assign n7896 = ~(n6382 ^ n5183);
assign n1171 = n11132 & n1854;
assign n6349 = n7805 | n11144;
assign n12203 = ~n8468;
assign n6277 = ~(n5563 ^ n1118);
assign n3091 = ~n2376;
assign n925 = n4846 & n7678;
assign n7449 = ~(n5091 ^ n907);
assign n8192 = ~(n4445 ^ n6970);
assign n8407 = ~(n8385 ^ n3406);
assign n7509 = ~(n13053 ^ n1851);
assign n2562 = n7557 & n3430;
assign n6279 = n13106 | n6963;
assign n4907 = n2118 | n4230;
assign n11874 = n1323 | n13238;
assign n2916 = n3026 | n13209;
assign n2572 = ~n10744;
assign n10830 = ~n8163;
assign n12544 = ~n7428;
assign n5968 = ~n11574;
assign n7585 = n10041 & n11741;
assign n1078 = n821 | n10904;
assign n8926 = n7930 | n7935;
assign n2979 = ~(n2091 ^ n5580);
assign n6834 = n3313 & n14;
assign n8886 = ~(n5250 ^ n11345);
assign n11955 = ~(n9254 ^ n5635);
assign n12393 = n8325 | n12695;
assign n12863 = n9891 ^ n4997;
assign n13103 = n1688 | n10871;
assign n3090 = ~(n3563 ^ n12460);
assign n2711 = ~n11109;
assign n11933 = ~n2341;
assign n3821 = n319 & n13145;
assign n5590 = n4132 | n7723;
assign n3759 = ~(n3042 | n12403);
assign n13189 = n9724 & n11956;
assign n12620 = ~n11181;
assign n4503 = n12017 & n2474;
assign n1723 = ~(n6948 ^ n4395);
assign n2198 = n3178 & n834;
assign n10942 = ~(n9624 ^ n5710);
assign n8384 = ~n4713;
assign n3136 = n9345 & n4003;
assign n2003 = n5321 | n1013;
assign n11584 = ~(n59 ^ n12209);
assign n2563 = n8143 | n12328;
assign n6580 = ~n6632;
assign n11557 = n11237 | n8494;
assign n4468 = n713 | n8319;
assign n7274 = ~(n10653 ^ n7397);
assign n5525 = ~(n4896 | n7910);
assign n93 = ~n7161;
assign n3668 = ~(n9960 | n9393);
assign n4153 = n2148 | n2133;
assign n13091 = n5122 & n35;
assign n3035 = n5586 & n2498;
assign n9614 = n7966 | n177;
assign n13243 = n5347 | n5373;
assign n96 = ~n9039;
assign n10876 = n2691 & n8363;
assign n8266 = n1783 | n2757;
assign n7207 = ~(n2987 | n2822);
assign n13010 = n5704 | n10194;
assign n6374 = n12212 | n3379;
assign n1617 = ~(n7064 ^ n11317);
assign n5776 = ~(n1722 ^ n12103);
assign n7139 = n575 | n12870;
assign n8917 = n5048 | n8702;
assign n3003 = n11893 & n11705;
assign n5914 = n7518 & n7112;
assign n2687 = n12178 | n7840;
assign n6135 = n2312 | n7820;
assign n8657 = n5055 & n5593;
assign n4932 = ~(n6757 | n11000);
assign n10824 = n3595 & n9109;
assign n634 = n1237 & n3216;
assign n11996 = n9527 | n4469;
assign n2137 = ~(n4831 ^ n13034);
assign n10325 = n10989 & n1226;
assign n6676 = n6347 | n12377;
assign n10828 = ~(n8584 ^ n4119);
assign n12238 = ~(n310 ^ n6503);
assign n1852 = ~(n9695 ^ n8305);
assign n7378 = n4516 & n5121;
assign n11917 = n12834 | n7950;
assign n2901 = n4566 | n8719;
assign n6157 = n7564 | n11415;
assign n5634 = ~n1084;
assign n10867 = n3239 & n3037;
assign n11146 = n9969 & n7732;
assign n1604 = ~(n12076 ^ n13162);
assign n7466 = ~(n7250 | n1822);
assign n9787 = n4619 & n5288;
assign n6020 = ~(n9094 ^ n431);
assign n8521 = n3870 & n5584;
assign n3576 = n7418 & n11744;
assign n3101 = n1621 | n8534;
assign n7734 = n4288 & n10503;
assign n6612 = n1868 | n2465;
assign n3485 = n940 & n568;
assign n1539 = n5857 | n6177;
assign n1026 = n8160;
assign n13148 = ~n8183;
assign n7697 = n9639 & n9168;
assign n10333 = ~(n1163 ^ n5022);
assign n4215 = n3940 | n8038;
assign n10934 = ~(n920 ^ n11282);
assign n2817 = ~(n2350 | n1073);
assign n6915 = ~(n1393 | n7708);
assign n6958 = n11719 & n8158;
assign n6291 = n12806 | n2589;
assign n6071 = ~(n2285 ^ n5304);
assign n13225 = n5032 & n6426;
assign n1391 = ~(n387 ^ n10887);
assign n10221 = ~n6794;
assign n12230 = n12023 | n3698;
assign n8258 = ~(n7503 ^ n3794);
assign n10800 = n937 & n3769;
assign n880 = n7661 | n11668;
assign n7280 = ~(n10048 ^ n12842);
assign n12739 = ~(n6526 ^ n8066);
assign n5829 = n7607 | n3501;
assign n12617 = ~n3832;
assign n2173 = n7167 | n12657;
assign n9556 = ~(n5335 ^ n3453);
assign n278 = ~n8714;
assign n9445 = n8243 | n11267;
assign n8649 = n351 & n9764;
assign n3265 = n9711 | n1463;
assign n12143 = n6515 & n2393;
assign n12595 = ~n9666;
assign n5307 = n3995 & n9899;
assign n12896 = ~(n1617 | n5596);
assign n8557 = ~(n12883 ^ n8441);
assign n4505 = n6492 & n11464;
assign n4668 = n114 | n121;
assign n3262 = ~(n1361 ^ n4849);
assign n5716 = n8926 & n5736;
assign n7190 = n710 | n11500;
assign n580 = ~(n8112 ^ n7940);
assign n10121 = ~(n8127 ^ n9298);
assign n8173 = ~n12284;
assign n1447 = ~n3076;
assign n12028 = ~(n4389 ^ n4746);
assign n2973 = n829 | n5242;
assign n9332 = n3013 | n2398;
assign n13237 = ~(n7697 | n11172);
assign n884 = n3096 | n12383;
assign n10093 = n3584 | n376;
assign n12778 = ~n7882;
assign n7898 = n4653 & n2514;
assign n6713 = ~(n3385 ^ n6485);
assign n10345 = ~n1148;
assign n11129 = ~(n2754 ^ n11458);
assign n11481 = n740 | n4847;
assign n524 = n5788 | n12811;
assign n11954 = n445 | n121;
assign n584 = ~n2771;
assign n6669 = n1571 | n13086;
assign n2740 = n3005 | n13017;
assign n6498 = ~(n8604 ^ n11030);
assign n4494 = n6371 | n10071;
assign n6856 = n12431 | n8385;
assign n3385 = n1152 | n9195;
assign n5635 = ~(n2532 ^ n8140);
assign n12082 = ~n32;
assign n11333 = ~n772;
assign n6445 = ~(n8009 ^ n6628);
assign n6293 = ~n2771;
assign n1064 = n937 & n8233;
assign n5007 = n10641 | n6635;
assign n11914 = ~n5012;
assign n11701 = n2546 | n8076;
assign n7930 = ~n3085;
assign n4270 = ~(n12047 | n5346);
assign n1932 = n11910 | n4490;
assign n9005 = ~n7087;
assign n5261 = ~n12912;
assign n8514 = ~n2071;
assign n12952 = ~n10544;
assign n3046 = n2518 & n5331;
assign n6106 = ~(n11637 | n2432);
assign n12426 = n11373 & n8829;
assign n9740 = n10066 | n6690;
assign n10617 = ~(n1233 | n13213);
assign n1289 = ~n2656;
assign n2925 = ~(n12167 ^ n11586);
assign n8072 = ~(n505 ^ n3377);
assign n5899 = ~n11561;
assign n4260 = ~n6920;
assign n12142 = ~(n8745 ^ n919);
assign n7154 = ~n3567;
assign n10304 = n2868 | n10350;
assign n2091 = n542 | n6404;
assign n4337 = n2122 & n7388;
assign n6424 = ~(n3775 ^ n3756);
assign n12533 = n2449 | n2675;
assign n5251 = ~n3226;
assign n4823 = n12795 | n4453;
assign n6214 = n2456 | n13233;
assign n1379 = n10920 | n5497;
assign n6440 = ~(n4154 ^ n898);
assign n3514 = ~n1038;
assign n234 = n6299 & n8064;
assign n7615 = n11080 & n10155;
assign n4945 = n1873 | n12074;
assign n2857 = ~(n4436 ^ n642);
assign n1947 = ~(n10211 | n3734);
assign n6155 = ~(n4742 ^ n11084);
assign n8029 = ~n12520;
assign n12740 = ~(n12720 ^ n12175);
assign n1206 = n5595 | n12388;
assign n5965 = n956 | n12188;
assign n11117 = ~(n1319 ^ n957);
assign n6684 = n4364 & n12165;
assign n2657 = ~n5920;
assign n6133 = ~n4335;
assign n9967 = n10929 | n6635;
assign n10881 = ~(n3753 ^ n6819);
assign n5942 = ~(n7984 ^ n12261);
assign n8821 = ~(n8474 ^ n1827);
assign n6517 = n44 | n4947;
assign n9594 = ~(n6473 | n10694);
assign n9667 = ~(n7931 ^ n915);
assign n2381 = ~(n3631 ^ n10841);
assign n12356 = n2605 & n5245;
assign n10992 = ~(n1658 ^ n7233);
assign n2311 = n1740 & n9881;
assign n10017 = ~n5969;
assign n10814 = ~n13060;
assign n4605 = n9625 | n1767;
assign n970 = n11236 & n6937;
assign n12596 = ~n854;
assign n7500 = ~(n9996 ^ n1721);
assign n454 = n3972 | n8534;
assign n13170 = ~n3085;
assign n7923 = n4885 & n585;
assign n1217 = ~(n8771 ^ n3842);
assign n12241 = ~n6009;
assign n8306 = ~n9906;
assign n4777 = ~(n4449 ^ n9077);
assign n6911 = n4387 | n726;
assign n9710 = ~n7208;
assign n6296 = ~(n12386 ^ n6261);
assign n9348 = ~(n3684 ^ n9189);
assign n3171 = n795 | n12930;
assign n5768 = n10770 & n6392;
assign n8103 = ~(n4617 | n5162);
assign n11140 = n1344 ^ n3950;
assign n6345 = n5176 | n3640;
assign n6401 = n5841 | n542;
assign n11930 = ~(n2555 ^ n11479);
assign n7235 = n11723 | n2893;
assign n8794 = ~(n10472 ^ n12148);
assign n10474 = ~n11324;
assign n3177 = n13068 & n7361;
assign n4725 = n10023 | n11042;
assign n9299 = n1989 | n7805;
assign n4549 = ~(n3592 ^ n11811);
assign n9784 = ~n1364;
assign n8923 = ~(n3441 ^ n3277);
assign n8372 = n9421 | n6732;
assign n11866 = n5801 & n10408;
assign n7350 = n2733 | n1272;
assign n9909 = n24 & n1593;
assign n13098 = n3646 | n6635;
assign n10495 = n8518 | n11750;
assign n4311 = ~(n729 ^ n1071);
assign n12227 = n7363 | n10;
assign n5786 = n10814 | n2675;
assign n9446 = ~(n6483 ^ n8991);
assign n8815 = n8529 | n8702;
assign n8686 = ~(n2283 ^ n3762);
assign n6391 = n8390 | n2076;
assign n6104 = ~(n9320 ^ n10449);
assign n7617 = ~(n67 ^ n5587);
assign n2317 = ~(n6468 ^ n8599);
assign n1874 = n2279 | n9126;
assign n5558 = n2346 | n12695;
assign n5992 = ~n10738;
assign n11834 = ~(n1642 ^ n12280);
assign n9316 = n2720 ^ n12645;
assign n9311 = ~n1405;
assign n5000 = ~(n8710 ^ n10933);
assign n13024 = n737 | n8702;
assign n8735 = ~(n5321 ^ n6351);
assign n6465 = n3516 | n3126;
assign n4923 = n10546 | n4667;
assign n11718 = n3222 | n4925;
assign n786 = n4758 & n6420;
assign n9453 = ~n12842;
assign n11655 = n12969 & n12686;
assign n2660 = ~n8867;
assign n13168 = ~n4330;
assign n270 = n3241 & n601;
assign n4115 = ~(n1343 | n11047);
assign n2706 = ~(n3879 | n4115);
assign n13021 = ~n4074;
assign n10838 = n10762 & n1675;
assign n1853 = ~(n13162 | n3883);
assign n9154 = ~n8522;
assign n738 = n9029 & n7679;
assign n2588 = ~(n12161 ^ n12455);
assign n4396 = ~n4698;
assign n10749 = n12448 | n7838;
assign n4127 = ~(n5499 | n5363);
assign n8708 = n6268 | n4358;
assign n186 = n9792 & n4995;
assign n13053 = n8508 & n13235;
assign n9680 = ~(n12928 ^ n2247);
assign n3111 = ~n2431;
assign n8234 = ~n10763;
assign n1097 = ~(n7716 ^ n7103);
assign n4092 = ~(n1968 ^ n9572);
assign n3331 = ~(n7286 | n8798);
assign n286 = n3767 | n11257;
assign n11534 = ~(n5199 ^ n2039);
assign n10670 = n6289 | n1614;
assign n611 = ~(n610 ^ n1275);
assign n7056 = n3268 | n6270;
assign n8968 = ~(n120 | n12028);
assign n7573 = n9627 | n12195;
assign n7356 = ~n9750;
assign n11121 = ~n691;
assign n8395 = ~(n1385 ^ n10554);
assign n11802 = ~(n13217 ^ n6550);
assign n8510 = ~n817;
assign n446 = ~(n5075 ^ n1430);
assign n5518 = n4473 | n7935;
assign n1914 = n3273 | n1780;
assign n658 = ~(n2259 ^ n949);
assign n12302 = n1933 & n9407;
assign n6205 = n1783 | n2958;
assign n6183 = ~n4591;
assign n512 = ~(n10645 | n7583);
assign n3285 = n12598 & n1003;
assign n4515 = ~n9475;
assign n11656 = ~(n1805 ^ n8694);
assign n10455 = n3729 & n11006;
assign n7498 = n596 | n1825;
assign n2984 = ~(n3009 ^ n10488);
assign n8412 = n11858 | n5873;
assign n6334 = ~(n10335 ^ n3966);
assign n6548 = ~(n3188 ^ n4002);
assign n13207 = n5360 | n6601;
assign n10903 = ~n4623;
assign n7826 = ~(n5255 | n10436);
assign n9416 = n9374 & n3389;
assign n12147 = ~(n1003 | n12598);
assign n11127 = n4793 | n10165;
assign n4187 = ~n5827;
assign n4592 = ~(n12532 ^ n1330);
assign n6513 = n11975 & n8408;
assign n8356 = n6689 | n10049;
assign n11661 = n13 | n2127;
assign n8830 = ~(n329 ^ n8479);
assign n9663 = n2791 ^ n4138;
assign n2097 = n2205 & n5095;
assign n3358 = n6808 & n1289;
assign n1268 = n10768 & n10154;
assign n2154 = n5872 & n1170;
assign n13215 = n10895 | n9014;
assign n12077 = n11060 & n5633;
assign n8596 = ~(n11903 ^ n5765);
assign n6798 = ~(n12805 ^ n4);
assign n3942 = ~(n3230 | n10486);
assign n6395 = ~(n277 ^ n7050);
assign n8316 = n9668 | n5242;
assign n10797 = n13011 ^ n13219;
assign n2099 = n7037 & n5337;
assign n7348 = n12109 | n6732;
assign n12374 = n3243 | n206;
assign n9395 = n8576 | n8825;
assign n10546 = ~(n3722 ^ n3903);
assign n7581 = ~(n13152 | n5950);
assign n7164 = n12722 & n2134;
assign n1699 = n11680 | n2542;
assign n3399 = n8892 & n4522;
assign n2455 = ~n1774;
assign n11289 = ~(n4853 ^ n12337);
assign n6877 = n4584 | n7723;
assign n5632 = ~(n1865 ^ n7922);
assign n1340 = ~(n12855 ^ n1670);
assign n9863 = ~(n3471 | n11287);
assign n3397 = n10830 | n6265;
assign n8105 = n8759 | n9075;
assign n243 = n9581 | n8348;
assign n3922 = n1284 | n10885;
assign n9714 = n9477 & n12611;
assign n6137 = n7505 | n8278;
assign n2514 = n4780 & n10623;
assign n8218 = n2211 & n7772;
assign n12098 = n7251 | n9229;
assign n1411 = ~(n11297 ^ n4100);
assign n11057 = ~(n2377 ^ n2147);
assign n4179 = ~n411;
assign n3610 = ~(n11625 ^ n12266);
assign n8993 = n12785 | n12900;
assign n3473 = n6280 | n742;
assign n12290 = n1113 | n8030;
assign n9387 = n13181 | n9444;
assign n1472 = n1035 | n8702;
assign n4848 = n10223 | n2082;
assign n10403 = n12105 & n10129;
assign n11853 = ~n11968;
assign n12941 = n11611 & n3985;
assign n5602 = n5342 | n2609;
assign n8564 = ~(n390 ^ n6328);
assign n1653 = ~(n5757 ^ n10119);
assign n1715 = n0 | n8348;
assign n4333 = ~n851;
assign n10647 = ~(n2780 ^ n7314);
assign n9260 = ~(n5469 ^ n8470);
assign n3739 = n8466 & n5536;
assign n2205 = ~(n10662 ^ n8303);
assign n1739 = n12619 | n5344;
assign n6272 = ~(n6363 | n6582);
assign n10131 = ~n12845;
assign n4584 = ~n11350;
assign n7849 = ~(n11188 ^ n7387);
assign n6129 = ~n443;
assign n2545 = ~n12267;
assign n7051 = ~(n11275 ^ n8459);
assign n7687 = ~(n3327 ^ n10729);
assign n2729 = n9842 & n4275;
assign n4331 = ~(n2721 ^ n9343);
assign n11187 = n4166 | n7530;
assign n12889 = ~n11290;
assign n10394 = ~(n3174 ^ n10136);
assign n10117 = ~n12005;
assign n12330 = ~n11715;
assign n11815 = ~n3378;
assign n1089 = ~n3669;
assign n3411 = n6174 ^ n4003;
assign n7694 = n6557 | n13108;
assign n7405 = ~(n11938 | n6592);
assign n6250 = ~n12651;
assign n8858 = ~n5981;
assign n2233 = ~(n5160 ^ n6510);
assign n583 = ~n962;
assign n12201 = ~(n13138 ^ n564);
assign n5419 = ~(n12866 ^ n9214);
assign n7870 = ~(n5113 | n9133);
assign n12127 = ~(n3642 | n11913);
assign n8172 = ~(n8543 ^ n582);
assign n9608 = n2786 & n8972;
assign n2654 = ~(n5095 ^ n2917);
assign n10933 = n10301;
assign n9073 = ~(n8507 ^ n9852);
assign n4617 = n8006 | n6178;
assign n8152 = n1200 & n7645;
assign n3276 = n9451 & n5366;
assign n5120 = n6755 | n2556;
assign n7381 = ~(n12147 | n4733);
assign n7555 = ~n3303;
assign n9244 = n12777 | n1034;
assign n8583 = ~(n11027 ^ n11693);
assign n5912 = ~(n739 ^ n11488);
assign n2408 = n10208 & n8683;
assign n1167 = ~(n8512 ^ n7658);
assign n1937 = ~(n491 ^ n9680);
assign n6120 = ~n9893;
assign n8791 = ~(n3785 ^ n12185);
assign n3185 = ~n11058;
assign n6238 = ~n342;
assign n12499 = ~(n10572 ^ n2703);
assign n12843 = n1194 | n206;
assign n5601 = n12102 | n2197;
assign n1894 = n4811 & n8787;
assign n10028 = n8355 & n2663;
assign n13033 = ~(n2644 | n2803);
assign n1585 = n45 | n9075;
assign n268 = ~(n7564 ^ n11415);
assign n11836 = ~(n5293 ^ n4409);
assign n2504 = ~n12965;
assign n7844 = n11175 & n6612;
assign n9700 = n8562 | n1985;
assign n7908 = ~n10538;
assign n1180 = n8391 & n5762;
assign n12855 = n12483 | n10573;
assign n7323 = n4293 ^ n7877;
assign n253 = n9434 & n3466;
assign n11266 = n3225 | n4936;
assign n9989 = n7072 & n12243;
assign n3907 = n8275 | n11712;
assign n2268 = n2944 | n7733;
assign n5710 = n5511 & n7913;
assign n5922 = n6751 | n5076;
assign n4663 = n6769 | n2675;
assign n10173 = n9699 & n1230;
assign n11745 = ~n4086;
assign n6086 = ~n9747;
assign n3097 = n5214 & n9669;
assign n12810 = ~(n568 ^ n7246);
assign n9485 = n4750 | n2460;
assign n12169 = ~n1494;
assign n2241 = ~(n5908 ^ n11469);
assign n7138 = ~(n3291 ^ n9198);
assign n10324 = n11680 | n11078;
assign n7836 = n2861 | n1026;
assign n12501 = n9257;
assign n9780 = n6447 | n5987;
assign n12830 = n8446 & n6413;
assign n12758 = ~n6023;
assign n508 = n4531 | n12909;
assign n4943 = n10911 | n2181;
assign n9078 = n1892 & n1679;
assign n5362 = ~(n1859 ^ n7816);
assign n8337 = n9436 | n3411;
assign n13232 = ~(n1427 ^ n5591);
assign n12403 = ~n10207;
assign n7080 = n11015 & n7955;
assign n7745 = ~(n6170 ^ n11181);
assign n514 = ~(n1625 | n1829);
assign n2379 = n4396 & n6893;
assign n8759 = ~n6826;
assign n2249 = n8685 & n3780;
assign n7250 = n504 & n7356;
assign n2354 = n11457 ^ n5991;
assign n2627 = n4497 & n8619;
assign n3928 = ~n11734;
assign n8640 = ~n7529;
assign n13089 = n10069 & n5419;
assign n3531 = ~n510;
assign n8914 = n8985 & n6585;
assign n11674 = n10898 | n12695;
assign n9919 = ~n4335;
assign n12115 = ~n10497;
assign n4281 = ~(n4457 ^ n4925);
assign n7104 = n1893 | n1570;
assign n3280 = n7745 | n418;
assign n12106 = ~(n6812 ^ n6548);
assign n13026 = ~n12263;
assign n1775 = n8646 | n6404;
assign n3159 = n121 | n2890;
assign n11849 = n1835 | n8509;
assign n5760 = n1700 | n11045;
assign n4754 = n6743 | n8702;
assign n4809 = n12039 & n8245;
assign n9156 = ~(n1760 ^ n8451);
assign n7299 = n1601 | n10508;
assign n10295 = ~(n5846 ^ n5597);
assign n10420 = ~(n6342 | n4093);
assign n3700 = n8428 | n8530;
assign n8765 = ~(n9845 ^ n7800);
assign n6167 = n12629 | n6732;
assign n7536 = ~(n95 ^ n4579);
assign n9086 = n11570 & n4239;
assign n10199 = n4628 | n12205;
assign n12932 = n9216 & n10606;
assign n6069 = ~(n9837 | n7290);
assign n2141 = ~n3631;
assign n5990 = ~n8290;
assign n372 = n1281 | n2672;
assign n9565 = n1857 & n9096;
assign n12914 = ~n4113;
assign n1646 = n2592 & n497;
assign n12728 = n11920 | n237;
assign n8630 = ~n4325;
assign n1958 = n10894 & n2503;
assign n12869 = ~(n8157 | n9086);
assign n1188 = ~n11222;
assign n7941 = ~(n7045 | n4069);
assign n8507 = ~(n7654 ^ n8555);
assign n5712 = n390 & n9439;
assign n13234 = n5013 | n84;
assign n2629 = ~(n3136 ^ n587);
assign n5340 = n5528 & n11377;
assign n1950 = ~(n2603 ^ n10224);
assign n2953 = ~(n5192 ^ n722);
assign n4049 = ~(n7609 | n11924);
assign n10471 = ~n12965;
assign n7416 = n189 | n5875;
assign n8392 = ~n10594;
assign n6545 = ~(n12880 | n8478);
assign n10815 = ~(n247 ^ n7995);
assign n8969 = n4837 & n6740;
assign n4402 = n11567 | n7526;
assign n10406 = ~(n335 ^ n10349);
assign n1424 = n3965 | n8941;
assign n10839 = ~(n3579 ^ n6998);
assign n3008 = n11236 & n10408;
assign n6307 = ~(n10415 ^ n6415);
assign n3437 = ~n10928;
assign n12706 = ~(n7413 | n8220);
assign n13018 = ~(n5625 | n9539);
assign n3249 = ~(n12819 ^ n7960);
assign n11780 = n2018 & n411;
assign n5148 = ~n10162;
assign n9331 = n2639 | n2675;
assign n6531 = ~(n6888 ^ n4671);
assign n2739 = ~(n6363 ^ n2328);
assign n5881 = n4660 & n6633;
assign n1173 = n12578 & n7163;
assign n964 = ~(n3939 ^ n9006);
assign n4984 = n891 | n1092;
assign n12381 = ~(n10867 ^ n10648);
assign n2121 = ~(n8750 ^ n12481);
assign n2659 = ~(n12091 ^ n9752);
assign n6646 = ~(n5030 ^ n11547);
assign n5192 = ~(n4699 ^ n13101);
assign n3183 = n6790 & n10398;
assign n2698 = n7534 & n7427;
assign n9811 = ~(n4609 | n2461);
assign n1015 = n1427 | n5591;
assign n1467 = n2636 & n7815;
assign n8684 = n3781 & n9485;
assign n7978 = ~(n3735 ^ n8484);
assign n10175 = n9025 & n11374;
assign n5344 = n252 & n10429;
assign n246 = ~(n4562 ^ n1384);
assign n2446 = ~n7012;
assign n5624 = n4657 | n1605;
assign n12025 = n2228 | n12604;
assign n1599 = n1438 | n479;
assign n1738 = n10724 & n9880;
assign n572 = n9723 | n12501;
assign n12384 = ~n5068;
assign n4838 = ~(n4920 | n6049);
assign n5502 = ~n5477;
assign n4160 = ~(n12276 | n5244);
assign n8869 = n6977 & n5007;
assign n9755 = ~(n359 ^ n7905);
assign n3800 = ~n5570;
assign n906 = ~n7569;
assign n10059 = ~n3815;
assign n4138 = ~(n7728 ^ n12956);
assign n32 = ~(n6212 ^ n6406);
assign n3537 = ~n1198;
assign n2977 = n5248 ^ n1689;
assign n10687 = ~(n6080 ^ n3463);
assign n3173 = ~n10482;
assign n2051 = n1029 & n10252;
assign n5163 = ~n1392;
assign n1883 = ~n9915;
assign n11514 = ~n4452;
assign n6823 = n10599 ^ n5117;
assign n11983 = n11514 | n7430;
assign n10082 = ~(n47 ^ n1728);
assign n9418 = n11020 & n2727;
assign n5546 = ~(n11719 ^ n5629);
assign n8081 = ~n4395;
assign n1389 = ~n246;
assign n785 = ~n12408;
assign n6942 = ~n7285;
assign n503 = n3008 & n9005;
assign n9888 = ~n2062;
assign n10132 = n5588 | n4640;
assign n11282 = n613 & n4137;
assign n11949 = ~(n1762 ^ n11003);
assign n8717 = n4453 | n3225;
assign n724 = ~(n10873 ^ n4512);
assign n6520 = n8020 | n10179;
assign n4779 = ~n9230;
assign n4063 = ~n9732;
assign n2618 = n8033 & n2949;
assign n5620 = n6524 & n5380;
assign n10344 = ~(n10064 ^ n12549);
assign n5785 = n7683 & n4592;
assign n7386 = n8966 | n9689;
assign n11389 = ~(n1278 ^ n2031);
assign n3718 = ~(n7794 ^ n9114);
assign n12444 = n5146 | n2958;
assign n693 = n5199 | n2039;
assign n8613 = ~n12936;
assign n11092 = n10439 | n7530;
assign n7492 = ~(n11776 ^ n3290);
assign n6720 = ~(n5907 | n5785);
assign n11710 = n3616 | n10179;
assign n10182 = ~n1330;
assign n5996 = n8609 | n9919;
assign n10163 = n11777 & n10774;
assign n4736 = n371 | n5186;
assign n5282 = ~(n535 | n8274);
assign n12349 = n12199 | n9582;
assign n8207 = n1051 | n5076;
assign n1296 = ~n3815;
assign n1926 = n11212 | n8702;
assign n5445 = n75 | n4936;
assign n10 = n11768 & n7836;
assign n12441 = ~n1636;
assign n12079 = ~(n11777 ^ n12761);
assign n2601 = n2434 | n2036;
assign n9360 = ~(n4681 | n1313);
assign n11998 = n6699 | n6265;
assign n6554 = ~(n2665 | n4759);
assign n5173 = n6981 & n1020;
assign n3312 = n673 & n366;
assign n170 = n7350 & n4180;
assign n13055 = n7213 & n8961;
assign n6096 = n11557 & n3375;
assign n9288 = n12122 | n6091;
assign n9837 = ~n336;
assign n5748 = n8778 | n1999;
assign n1935 = n6219 & n6734;
assign n12911 = n3225 | n6404;
assign n8676 = n6810 | n10871;
assign n4594 = n2018 & n13058;
assign n10331 = ~n13064;
assign n8066 = n12349 & n8444;
assign n11173 = n1850 & n8882;
assign n1647 = n4999 | n5652;
assign n1166 = ~(n6712 | n6578);
assign n1911 = ~(n11024 ^ n3156);
assign n5913 = ~(n5228 ^ n3330);
assign n10019 = n1431 & n10856;
assign n11005 = n11929 | n9268;
assign n10999 = n6063 | n1463;
assign n7551 = n1305 & n747;
assign n8726 = n7134 | n8247;
assign n6647 = ~(n5584 ^ n825);
assign n11216 = ~(n7836 ^ n11768);
assign n9448 = n909 & n4805;
assign n6619 = ~(n5702 ^ n12201);
assign n7802 = ~(n8549 ^ n5804);
assign n7779 = n11559 ^ n8542;
assign n5225 = ~(n9037 | n7599);
assign n9286 = ~n7;
assign n1919 = ~n8290;
assign n2661 = n7741 | n9159;
assign n11213 = n718 | n12862;
assign n12168 = n5565 | n1144;
assign n7359 = ~(n13031 ^ n3073);
assign n6747 = ~(n8 ^ n4401);
assign n9277 = n1325 | n3825;
assign n5740 = ~n8139;
assign n11571 = n7819 | n2449;
assign n9560 = ~(n10431 ^ n9299);
assign n6761 = ~(n2518 | n5331);
assign n8544 = ~(n5185 ^ n9650);
assign n2957 = ~(n5072 ^ n9289);
assign n6446 = n10411 | n11239;
assign n2074 = n6447 & n5987;
assign n6988 = ~n10657;
assign n11864 = ~n3832;
assign n1187 = n6180 & n1862;
assign n8217 = ~(n11464 ^ n11651);
assign n4034 = n11094 | n4936;
assign n2929 = ~(n10630 ^ n2690);
assign n5153 = n11648 | n8805;
assign n7517 = n6749 | n2943;
assign n11736 = ~(n12312 ^ n12239);
assign n10722 = ~(n223 ^ n1590);
assign n7873 = n8915 & n12012;
assign n4897 = ~(n9138 ^ n11254);
assign n8565 = n12254 | n4230;
assign n9530 = ~(n13171 ^ n7536);
assign n1870 = ~(n2388 ^ n4186);
assign n4499 = ~n5603;
assign n5728 = ~(n13196 ^ n4727);
assign n3506 = n1328 & n6741;
assign n12354 = n6173 | n4116;
assign n8650 = ~n7725;
assign n3594 = ~(n5324 ^ n3074);
assign n12773 = n9580 | n486;
assign n5995 = n5449 & n5855;
assign n593 = n10351 | n8448;
assign n8124 = ~(n9247 ^ n2979);
assign n11719 = ~(n6926 ^ n746);
assign n5964 = n6901 | n11670;
assign n10252 = n745 | n982;
assign n4843 = ~(n1932 ^ n7850);
assign n10827 = ~(n3708 ^ n5496);
assign n12986 = ~n8520;
assign n7545 = n6086 | n5076;
assign n7921 = n7862 | n9861;
assign n11096 = n2416 | n8348;
assign n12864 = ~(n9878 | n3030);
assign n5096 = n10147 & n2564;
assign n7445 = ~(n5431 ^ n4429);
assign n1254 = n8183 & n854;
assign n6901 = n8953 & n3880;
assign n9384 = n10509 | n11928;
assign n9600 = n5233 | n9579;
assign n7726 = ~(n3161 ^ n251);
assign n8177 = n6492 | n11464;
assign n3344 = ~n10162;
assign n12670 = n12615 & n7667;
assign n2119 = ~(n4187 ^ n2216);
assign n3152 = ~(n6607 ^ n7116);
assign n12087 = n2194 & n5109;
assign n11548 = ~n9093;
assign n6479 = n10798 | n10179;
assign n4787 = n8264 & n10834;
assign n8443 = n12894 | n2969;
assign n3988 = ~(n12652 ^ n10076);
assign n6351 = ~(n615 ^ n8386);
assign n11228 = n3928 | n12501;
assign n4882 = ~(n3886 ^ n8899);
assign n1630 = n2823 | n566;
assign n8959 = n11761 | n6874;
assign n12223 = ~(n5615 | n805);
assign n11134 = ~(n3006 ^ n5568);
assign n12468 = ~(n5616 ^ n5332);
assign n6059 = ~(n11203 ^ n3926);
assign n2265 = n11084 | n3479;
assign n10489 = n5923 | n8188;
assign n8082 = ~n2295;
assign n8283 = ~(n2437 ^ n691);
assign n6553 = ~(n1450 ^ n703);
assign n8996 = n3903 & n3722;
assign n2736 = ~(n2137 ^ n342);
assign n5738 = n9019 | n8348;
assign n7854 = n5671 & n4335;
assign n5333 = n11745 & n1920;
assign n1133 = n13127 & n452;
assign n11614 = ~n6857;
assign n13159 = ~n6818;
assign n10055 = ~(n9384 ^ n2401);
assign n7945 = ~n12391;
assign n5771 = n5544 | n3372;
assign n10150 = n2062 ^ n6394;
assign n1400 = n11928 | n2958;
assign n14 = n6672 | n1043;
assign n8321 = n1997 & n4054;
assign n11434 = n11324 & n12284;
assign n5501 = ~(n2536 ^ n982);
assign n9675 = ~n353;
assign n3286 = n629 & n5153;
assign n901 = ~(n7545 ^ n4276);
assign n5549 = ~(n2569 ^ n4590);
assign n5137 = ~(n3974 ^ n11906);
assign n13032 = n1009 & n8296;
assign n6478 = n9032 & n3235;
assign n6624 = ~(n9190 ^ n9503);
assign n8185 = n9776 | n8587;
assign n8238 = ~(n6513 | n2475);
assign n6771 = ~(n6310 ^ n9950);
assign n296 = ~(n12649 ^ n11983);
assign n7942 = ~n2043;
assign n1124 = ~(n5649 | n8695);
assign n2655 = n10168 & n3832;
assign n4286 = n3413 & n9708;
assign n2833 = n3062 | n542;
assign n4169 = n4133 & n11915;
assign n5250 = n2688 | n6265;
assign n5458 = ~(n3683 ^ n9832);
assign n5817 = n12077 & n5125;
assign n12321 = n9474 ^ n11854;
assign n8383 = ~n2771;
assign n1345 = ~n2758;
assign n4365 = n304 | n10079;
assign n5044 = n13075 & n2390;
assign n11696 = ~n12560;
assign n5848 = n6543 & n13187;
assign n12121 = ~(n8242 ^ n10209);
assign n991 = ~n12306;
assign n9865 = ~(n8238 | n725);
assign n6273 = n4888 & n6579;
assign n3221 = ~(n8989 | n3);
assign n6084 = n4462 | n8702;
assign n3049 = ~n9732;
assign n1559 = n10481 | n8563;
assign n3799 = n3795 & n1736;
assign n2448 = n11105 & n9355;
assign n7791 = ~n3029;
assign n9969 = n4536 | n10057;
assign n2677 = n7291 | n5076;
assign n6600 = ~(n11587 ^ n2684);
assign n10605 = n12235 & n12204;
assign n11784 = ~n4703;
assign n12935 = n10950 | n8268;
assign n564 = n3867 & n442;
assign n12420 = ~(n11501 | n7630);
assign n1011 = n536 | n6834;
assign n8206 = ~n5962;
assign n1137 = n1428 & n9191;
assign n1736 = n5447 | n4861;
assign n1036 = ~(n9958 ^ n12461);
assign n11951 = n4716 | n6055;
assign n1131 = n2449 | n7935;
assign n5006 = ~(n11774 | n3828);
assign n2166 = ~n4709;
assign n10343 = n7342;
assign n7282 = ~(n434 ^ n3787);
assign n2131 = ~n8535;
assign n12888 = n3265 | n2188;
assign n2443 = ~n11553;
assign n9304 = n1484 | n3432;
assign n4077 = ~n3769;
assign n12222 = n3459 | n3225;
assign n4367 = ~(n12764 ^ n7319);
assign n853 = ~(n1523 | n9002);
assign n4364 = n6803 | n8763;
assign n983 = n1876 ^ n9303;
assign n683 = ~n7061;
assign n1021 = n8308 & n3409;
assign n5493 = ~(n11184 ^ n8258);
assign n12754 = n6769 | n1570;
assign n4544 = n13080 | n4337;
assign n12731 = ~(n9004 ^ n11735);
assign n6118 = ~(n970 ^ n997);
assign n12380 = ~n11814;
assign n12955 = ~n103;
assign n10635 = ~(n6929 ^ n12664);
assign n2776 = ~(n163 ^ n3065);
assign n4870 = n5238 & n5350;
assign n4159 = n10270 | n9595;
assign n10070 = ~(n3603 ^ n1622);
assign n2418 = ~(n9792 ^ n11428);
assign n7042 = n5547 | n3981;
assign n7583 = n1480 | n905;
assign n9065 = ~(n3477 ^ n7861);
assign n9550 = ~(n10834 ^ n8264);
assign n1308 = ~n13044;
assign n9901 = ~(n4830 ^ n10541);
assign n715 = ~n11396;
assign n10822 = n3288 | n5291;
assign n962 = n8840 & n13157;
assign n10299 = ~(n6574 | n7614);
assign n4088 = n6960 | n4723;
assign n743 = ~(n11585 ^ n12094);
assign n8305 = n9060 & n8722;
assign n10041 = ~n2535;
assign n9000 = ~(n12411 ^ n4745);
assign n11179 = ~(n2896 ^ n1061);
assign n1234 = n5973 | n9075;
assign n7955 = n12481 | n8750;
assign n5054 = n3296 | n3114;
assign n9562 = ~(n1827 | n13059);
assign n716 = n9144 & n6870;
assign n1638 = ~n5729;
assign n2463 = ~n12289;
assign n10537 = n2045 & n1032;
assign n9983 = ~(n4152 ^ n2159);
assign n10959 = n511 | n12162;
assign n6613 = ~(n2495 | n2026);
assign n1526 = ~n2813;
assign n12 = ~(n6593 ^ n2511);
assign n4719 = n3040 ^ n7761;
assign n12276 = ~(n7898 ^ n11285);
assign n12174 = ~n6392;
assign n1974 = ~(n12736 ^ n1994);
assign n9583 = ~(n1304 ^ n4718);
assign n1506 = n12348 & n469;
assign n2484 = ~n10594;
assign n5515 = n5138 & n8784;
assign n3469 = n8324 | n8702;
assign n10523 = ~(n9914 ^ n697);
assign n8148 = n3070 | n4930;
assign n8943 = n6156 | n10207;
assign n9699 = n1011 & n3350;
assign n4675 = ~(n2010 | n10661);
assign n12452 = n7608 | n12388;
assign n1017 = ~n5881;
assign n7527 = ~(n3846 ^ n6277);
assign n10392 = n6209 ^ n11084;
assign n5286 = ~n7573;
assign n5 = ~n11511;
assign n9335 = ~(n3988 | n2445);
assign n6615 = n12390 & n1075;
assign n6502 = n10150 | n9512;
assign n10167 = ~(n10746 ^ n4712);
assign n6634 = n2230 | n12120;
assign n7574 = ~(n4391 ^ n6102);
assign n11351 = n3420 & n6123;
assign n2495 = n6755 | n8374;
assign n5621 = ~(n5391 ^ n9231);
assign n4819 = n7947 & n12601;
assign n2862 = n9484 | n2842;
assign n11598 = ~(n7227 ^ n5231);
assign n3201 = ~n7713;
assign n3740 = ~(n11688 ^ n5374);
assign n2157 = ~n11692;
assign n3855 = ~(n8331 | n798);
assign n1311 = n2933 | n13225;
assign n3770 = n2041 | n1144;
assign n1740 = n787 | n4947;
assign n10705 = ~(n1321 | n3144);
assign n3383 = ~(n6107 | n9988);
assign n12008 = ~(n4754 | n3533);
assign n8743 = n11291 | n1026;
assign n12365 = n4227 | n3418;
assign n1790 = n8469 ^ n9473;
assign n1274 = n4308 | n3820;
assign n5904 = n9659 | n395;
assign n702 = n8234 & n10820;
assign n2743 = ~(n6153 ^ n2392);
assign n9830 = n5079 | n8030;
assign n9149 = n1158 & n1713;
assign n633 = ~n5309;
assign n11022 = n361 | n3039;
assign n265 = n3847 & n10065;
assign n11048 = ~(n12458 ^ n1151);
assign n4771 = n1919 | n8348;
assign n2843 = ~(n11720 ^ n4045);
assign n10565 = ~n8092;
assign n7485 = ~n8518;
assign n2757 = ~n9732;
assign n4655 = ~n3188;
assign n10485 = n7040 ^ n3763;
assign n106 = ~(n9592 | n2668);
assign n3347 = ~(n9209 | n6528);
assign n6792 = ~(n3749 | n46);
assign n538 = n1141 | n8937;
assign n773 = ~(n172 ^ n4973);
assign n5818 = n4456 | n5353;
assign n8651 = ~(n3558 ^ n11766);
assign n12719 = ~(n9138 | n11254);
assign n3546 = ~(n8867 | n9827);
assign n520 = ~(n3236 ^ n9197);
assign n10935 = n1102 & n11908;
assign n531 = ~(n12135 ^ n6714);
assign n2852 = ~(n11881 ^ n6991);
assign n5505 = n146 & n95;
assign n1776 = ~(n12056 ^ n446);
assign n9735 = n9152 & n6457;
assign n7160 = ~(n12949 ^ n8818);
assign n9561 = ~(n9220 | n8333);
assign n1149 = ~(n9496 ^ n8034);
assign n3580 = n2838 & n2388;
assign n1482 = n646 & n47;
assign n6965 = ~(n11279 ^ n11454);
assign n601 = ~(n8241 ^ n7462);
assign n5535 = n3311 & n10606;
assign n10381 = ~n8284;
assign n8248 = ~n9825;
assign n4039 = ~(n5655 ^ n2206);
assign n10629 = ~(n4199 | n6938);
assign n12275 = ~(n2173 ^ n3490);
assign n5465 = n5433 | n4230;
assign n10212 = n12832 | n1690;
assign n9970 = n9723 | n10871;
assign n3608 = ~(n4026 | n1243);
assign n1168 = ~n10162;
assign n8144 = ~(n7578 ^ n6775);
assign n12845 = ~(n264 ^ n6500);
assign n10682 = n856 | n8602;
assign n11487 = n5226 | n8024;
assign n11077 = ~(n5073 ^ n12962);
assign n9098 = n2932 & n11182;
assign n3708 = n2346 | n8348;
assign n6490 = n9066 | n7681;
assign n10566 = n9444 | n4373;
assign n13047 = ~(n11338 ^ n6609);
assign n3650 = n9864 & n4224;
assign n8702 = n4013;
assign n12291 = ~(n6583 ^ n1142);
assign n9855 = n7673 & n1223;
assign n5335 = n11404 | n12273;
assign n9325 = ~n8827;
assign n6223 = ~n4006;
assign n5750 = n11969 & n4560;
assign n6076 = n10220 | n12215;
assign n1004 = n570 & n3366;
assign n8295 = ~n11017;
assign n2005 = n7828 & n3888;
assign n12067 = ~(n7734 ^ n1374);
assign n2040 = ~(n11722 ^ n7502);
assign n12615 = ~n12961;
assign n487 = n2590 & n7720;
assign n1120 = ~(n10160 ^ n10625);
assign n4734 = ~(n4094 ^ n5323);
assign n4869 = n3095 | n2983;
assign n9653 = n3480 | n3119;
assign n8023 = ~(n8801 ^ n12509);
assign n5110 = ~(n11456 ^ n7589);
assign n7070 = ~(n2065 ^ n1565);
assign n9458 = ~(n8547 ^ n416);
assign n10500 = n5782 | n10319;
assign n3883 = n12270 & n12076;
assign n1726 = ~(n6372 ^ n10624);
assign n806 = ~(n271 ^ n12647);
assign n1170 = n5105 | n8505;
assign n1691 = n385 | n13056;
assign n6964 = ~(n2564 ^ n10147);
assign n4393 = n7748 | n2133;
assign n12589 = n12705 & n9051;
assign n9825 = ~(n2677 ^ n6708);
assign n687 = ~(n2886 ^ n8854);
assign n3275 = n9559 | n4690;
assign n9045 = ~(n5439 | n10315);
assign n6477 = ~(n1509 ^ n2563);
assign n1606 = n10498 | n10889;
assign n5534 = ~(n8825 ^ n8576);
assign n5857 = ~(n9625 ^ n12950);
assign n602 = ~n2824;
assign n2093 = ~(n6697 ^ n1842);
assign n5603 = n8941 | n5797;
assign n13078 = n840 & n6667;
assign n427 = n3006 & n4470;
assign n12813 = ~n11897;
assign n4789 = n8940 & n11222;
assign n8028 = n9761 | n1570;
assign n4305 = ~n10111;
assign n8346 = n9502 | n2719;
assign n3760 = n10908 & n10408;
assign n11102 = ~(n6426 ^ n5032);
assign n6616 = ~(n109 ^ n3287);
assign n3232 = ~n62;
assign n126 = n2488 | n793;
assign n7227 = n2825 | n6404;
assign n4068 = ~(n9630 | n12359);
assign n12253 = n3333 | n6715;
assign n4102 = n1978 ^ n3168;
assign n10977 = ~n2174;
assign n11673 = n11236 & n854;
assign n9923 = ~(n12389 | n7539);
assign n3930 = ~(n11913 ^ n8409);
assign n3896 = ~(n10969 ^ n2843);
assign n9628 = n2625 | n4386;
assign n9754 = ~(n7833 | n791);
assign n2209 = n12141 & n10513;
assign n3630 = ~n22;
assign n3655 = ~n3123;
assign n5705 = n8817 | n10106;
assign n10391 = n898 | n4154;
assign n4959 = n2860 & n10125;
assign n1062 = n6038 | n1468;
assign n1707 = ~(n9248 ^ n6872);
assign n1384 = ~(n7201 ^ n11337);
assign n2226 = ~n12605;
assign n7283 = ~n1307;
assign n8370 = n2444 | n11461;
assign n2114 = n11094 | n7530;
assign n6442 = n1452 & n5503;
assign n13030 = ~(n4097 | n12876);
assign n12279 = ~(n6573 ^ n9671);
assign n9420 = n3974 | n9018;
assign n5353 = n8498 | n4373;
assign n8609 = ~n11061;
assign n9737 = n6024 & n4915;
assign n9340 = ~n13161;
assign n8439 = ~(n11444 | n12430);
assign n5850 = n9679 | n9118;
assign n5894 = ~(n11332 ^ n4240);
assign n11586 = ~(n10316 ^ n12022);
assign n12772 = ~n4293;
assign n11126 = ~(n7796 ^ n4829);
assign n3391 = ~(n6778 ^ n12110);
assign n187 = ~(n11005 ^ n1896);
assign n8849 = ~n12482;
assign n6969 = ~(n155 ^ n9806);
assign n9440 = ~(n8536 ^ n3896);
assign n9346 = n3425 | n1028;
assign n11645 = n2888 & n3764;
assign n10697 = n5483 & n6889;
assign n1553 = n583 | n11405;
assign n2927 = n12022 & n10316;
assign n2594 = ~(n691 | n1874);
assign n8196 = n1751 & n9801;
assign n1924 = ~(n10054 | n10651);
assign n1386 = ~(n9944 ^ n1898);
assign n8696 = n8124 & n4262;
assign n10743 = ~(n6943 ^ n7030);
assign n9823 = ~(n12021 ^ n11695);
assign n4915 = n7597 | n6732;
assign n596 = n10286 | n6944;
assign n6305 = n10898 | n12847;
assign n11095 = n9400 | n8030;
assign n18 = ~n4357;
assign n3566 = n13096 & n6146;
assign n11566 = n8431 | n12666;
assign n2116 = n7891 & n8048;
assign n9574 = ~(n6513 ^ n725);
assign n9734 = ~(n3964 | n6879);
assign n3453 = n0 | n4230;
assign n1430 = n6444 & n11489;
assign n12178 = n11171 | n12847;
assign n8280 = ~n4368;
assign n10241 = n12312 | n12781;
assign n3925 = ~(n4953 ^ n8119);
assign n556 = ~(n8313 ^ n1715);
assign n13051 = ~n9669;
assign n10232 = n7677 | n12048;
assign n1044 = n11951 & n11936;
assign n2985 = n4690 & n9559;
assign n7397 = ~(n11875 ^ n11755);
assign n6575 = ~n4695;
assign n5371 = n1183 & n7747;
assign n6134 = ~(n8867 ^ n2382);
assign n10813 = n8208 & n12375;
assign n4548 = ~(n2208 ^ n3402);
assign n9512 = ~n2334;
assign n3393 = n4655 | n6924;
assign n8049 = ~(n10878 ^ n8308);
assign n361 = n1510 & n12816;
assign n2008 = n8090 | n11282;
assign n8225 = ~n5729;
assign n8924 = n4967 | n3981;
assign n3567 = n1499 & n1210;
assign n11427 = ~n12937;
assign n4348 = n12003 & n11109;
assign n9201 = ~(n6131 ^ n9757);
assign n4684 = n4977 & n6864;
assign n3644 = n12920 & n9727;
assign n7695 = n12477 | n8231;
assign n3586 = ~n3263;
assign n9429 = ~n9528;
assign n36 = n3049 | n5264;
assign n473 = ~n4459;
assign n7125 = n11588 | n8748;
assign n12247 = ~(n7671 | n8078);
assign n430 = n10138 | n9386;
assign n3289 = ~(n8944 ^ n6567);
assign n2803 = n7650 & n3657;
assign n6329 = n345 | n1961;
assign n1590 = ~(n10294 ^ n13222);
assign n4051 = ~(n10992 ^ n8015);
assign n7600 = n3564 | n10029;
assign n8554 = ~(n3204 ^ n4729);
assign n4699 = ~(n7161 | n8030);
assign n11704 = n2262 | n4865;
assign n290 = ~n5457;
assign n6366 = ~n3625;
assign n10699 = ~(n4086 ^ n1920);
assign n2026 = n889 & n7897;
assign n1329 = ~n11429;
assign n1451 = ~n9906;
assign n3318 = ~n6604;
assign n763 = ~(n1170 ^ n5872);
assign n2196 = ~(n5128 ^ n6200);
assign n2783 = n987 | n10319;
assign n2039 = ~(n4467 ^ n12142);
assign n482 = ~n2777;
assign n6865 = ~(n346 ^ n5755);
assign n2528 = n3726 | n2133;
assign n3494 = ~(n8476 ^ n10689);
assign n788 = ~(n9892 ^ n10526);
assign n3756 = ~(n13 ^ n11687);
assign n4579 = n5832 & n3303;
assign n12436 = ~(n4508 ^ n11432);
assign n11947 = n4715 | n6561;
assign n11926 = ~n9127;
assign n7033 = ~n9093;
assign n6985 = ~(n11393 ^ n2997);
assign n1551 = ~(n12247 | n10754);
assign n12571 = ~(n4525 ^ n7684);
assign n979 = n4931 & n11084;
assign n7846 = ~n2590;
assign n3190 = ~(n8747 ^ n10737);
assign n11807 = ~n8359;
assign n328 = ~(n6525 ^ n8232);
assign n12401 = n6995 & n8690;
assign n2306 = ~n2979;
assign n6062 = n11263 & n13081;
assign n13192 = n6830 & n3786;
assign n1297 = n8197 & n10245;
assign n10413 = n13146 | n8564;
assign n1811 = ~(n6700 ^ n5277);
assign n7162 = ~(n9553 ^ n6059);
assign n5679 = ~n6655;
assign n11205 = ~(n3699 ^ n4976);
assign n4831 = n8111 & n2967;
assign n370 = ~(n12453 ^ n7766);
assign n5228 = n1737 | n9638;
assign n3155 = n925 & n8199;
assign n3103 = ~n11332;
assign n10681 = ~n3130;
assign n12438 = ~n6251;
assign n1766 = n12568 | n8534;
assign n7811 = n829 | n9075;
assign n4988 = n6986 | n10430;
assign n123 = n991 | n12501;
assign n4350 = n9662 & n10386;
assign n4359 = n1536 | n2675;
assign n5205 = n2044 & n12293;
assign n12639 = ~(n3542 ^ n5418);
assign n9292 = n7434 & n8185;
assign n7040 = n2163 & n2618;
assign n9775 = ~(n5689 ^ n2467);
assign n12655 = ~n10408;
assign n13174 = n2698 | n9203;
assign n1621 = ~n10162;
assign n11087 = ~n5470;
assign n9790 = ~n9965;
assign n2436 = n2407 & n2578;
assign n8277 = n1571 | n7935;
assign n3396 = n10884 & n5926;
assign n9841 = ~(n12074 ^ n11767);
assign n7409 = n11490 & n1206;
assign n6259 = n13182 | n1985;
assign n2327 = n794 | n2980;
assign n7182 = n3336 & n5685;
assign n11177 = ~(n752 ^ n3982);
assign n13097 = ~n9049;
assign n3887 = ~(n3836 ^ n11892);
assign n2676 = n7722 & n11485;
assign n5843 = n1987 | n285;
assign n13092 = ~(n6712 ^ n12186);
assign n10958 = n7010 & n2752;
assign n8758 = ~(n9609 ^ n3134);
assign n2626 = ~(n12942 ^ n717);
assign n12182 = ~(n10109 ^ n3232);
assign n7231 = n560 | n8490;
assign n3927 = n7231 | n6583;
assign n1352 = ~(n12816 | n1510);
assign n9684 = n3102 & n10385;
assign n2083 = ~n791;
assign n1342 = n6137 & n6379;
assign n1944 = ~(n3357 ^ n3012);
assign n9281 = ~n11508;
assign n886 = ~(n8122 ^ n8995);
assign n7303 = n5076 | n10106;
assign n5532 = ~(n1391 ^ n3737);
assign n11958 = n12493 | n177;
assign n6644 = n10761 | n206;
assign n6298 = ~(n7161 | n5076);
assign n3392 = n9353 & n10063;
assign n1700 = ~(n9074 ^ n4799);
assign n414 = ~(n9939 ^ n2356);
assign n3366 = n8174 | n2958;
assign n12732 = ~n12965;
assign n9870 = ~(n6053 | n3080);
assign n4765 = ~(n6661 ^ n6675);
assign n4581 = ~(n14 ^ n3313);
assign n7284 = n3505 | n6689;
assign n6180 = ~n1283;
assign n2453 = ~n11890;
assign n380 = ~(n8240 ^ n5373);
assign n6433 = n1912 & n2498;
assign n11060 = n12660 | n4881;
assign n11873 = n5768 & n10563;
assign n5682 = ~(n8823 ^ n4434);
assign n2782 = n1250 | n3113;
assign n7011 = n12395 | n4960;
assign n6701 = ~(n8207 ^ n1106);
assign n8963 = n8847 & n3007;
assign n5979 = ~(n12279 ^ n9210);
assign n10140 = n848 & n10620;
assign n7379 = n10196 & n10104;
assign n8700 = ~n4813;
assign n9764 = n5770 | n4312;
assign n11541 = ~(n4639 ^ n1457);
assign n4919 = n7468 & n8442;
assign n12347 = ~(n7910 ^ n11358);
assign n7115 = ~(n5126 ^ n1363);
assign n5870 = n4964 & n510;
assign n13088 = ~n6537;
assign n4413 = n5661 & n7174;
assign n6786 = n5092 & n12462;
assign n7738 = n2829 | n228;
assign n10627 = ~(n4661 ^ n8713);
assign n4874 = n11288 ^ n8408;
assign n5084 = n2643 & n4629;
assign n7455 = n4828 ^ n8197;
assign n11683 = ~n6937;
assign n6070 = n10792 | n542;
assign n8530 = n4863 & n243;
assign n667 = n11239 | n8030;
assign n7003 = n8240 | n9123;
assign n141 = ~(n7289 ^ n5463);
assign n10484 = ~(n1756 ^ n6380);
assign n8456 = ~(n9871 ^ n9350);
assign n2036 = ~(n5810 ^ n10720);
assign n9407 = n2582 | n6635;
assign n4053 = n4201 | n11144;
assign n5433 = ~n9887;
assign n8129 = ~n5962;
assign n11238 = n1053 | n9491;
assign n11004 = ~(n9433 ^ n5628);
assign n7222 = n6651 | n2658;
assign n9659 = n8585 | n4640;
assign n4116 = ~n3130;
assign n13096 = n3069 | n8365;
assign n7909 = ~(n9602 ^ n2870);
assign n3723 = n8900 & n5284;
assign n85 = ~(n8256 ^ n5582);
assign n6405 = ~n124;
assign n9245 = ~n9214;
assign n2515 = ~n8924;
assign n10725 = n12007 & n2066;
assign n677 = n1558 | n1692;
assign n13028 = ~n9732;
assign n12687 = ~(n4458 | n9091);
assign n4701 = n2214 | n10589;
assign n395 = n11466 | n479;
assign n5258 = ~(n6009 | n11089);
assign n5372 = ~n6998;
assign n10430 = ~n3130;
assign n3970 = ~n11306;
assign n2994 = ~(n13144 ^ n4911);
assign n12619 = ~(n2767 ^ n6617);
assign n8135 = ~(n10623 ^ n1902);
assign n1547 = ~(n986 ^ n9471);
assign n1882 = ~(n8064 ^ n3843);
assign n1573 = ~(n7476 ^ n11948);
assign n13241 = n11915 | n4133;
assign n7586 = ~n8398;
assign n6011 = n590 & n11168;
assign n6539 = ~(n7100 | n9045);
assign n6145 = ~(n10785 | n429);
assign n12361 = ~(n9901 ^ n1350);
assign n6107 = ~(n9344 ^ n5735);
assign n11006 = ~n1065;
assign n10809 = n864 & n8458;
assign n1350 = ~(n11801 ^ n6216);
assign n11680 = ~n11891;
assign n2763 = n1280 | n12907;
assign n8718 = n1346 & n5839;
assign n13015 = ~(n1537 ^ n5464);
assign n8623 = ~(n2323 | n183);
assign n8046 = n937 & n287;
assign n212 = n5257 & n8425;
assign n11158 = ~(n11108 ^ n887);
assign n153 = ~n1721;
assign n8022 = n5231 | n7227;
assign n1445 = n3780 | n8685;
assign n2186 = n3639 & n503;
assign n9213 = ~(n10540 ^ n8343);
assign n3459 = ~n3669;
assign n3906 = ~n11881;
assign n6466 = n7604 | n4585;
assign n6927 = ~(n659 ^ n1591);
assign n1802 = ~(n5465 ^ n7760);
assign n2755 = n7986 | n8540;
assign n6859 = n8776 | n10761;
assign n1979 = n10221 | n2977;
assign n8158 = n12953 ^ n6140;
assign n2462 = ~n13058;
assign n7194 = n6971 | n3798;
assign n11274 = ~(n3224 ^ n340);
assign n8606 = n9353 & n9915;
assign n13146 = ~n3868;
assign n5014 = ~(n9858 ^ n618);
assign n6295 = ~n2758;
assign n5124 = ~(n10167 ^ n4643);
assign n5213 = ~(n11572 | n1584);
assign n10970 = ~(n7887 ^ n626);
assign n3964 = ~(n9938 ^ n8184);
assign n8577 = n9797 & n12584;
assign n9527 = ~(n2541 | n11280);
assign n12417 = n48 | n11144;
assign n4206 = n3755 | n2845;
assign n7933 = n13168 | n1985;
assign n2466 = n2861 | n12388;
assign n4414 = n12734 & n2441;
assign n10761 = n6405;
assign n6379 = n5700 | n9975;
assign n3527 = n12596 | n5242;
assign n7900 = ~n9747;
assign n1778 = n12745 & n1968;
assign n11511 = n10343 | n6983;
assign n11676 = ~(n6296 ^ n11073);
assign n7089 = ~n6286;
assign n8621 = ~n9415;
assign n7123 = ~(n11004 ^ n5994);
assign n12423 = ~(n90 ^ n6262);
assign n8377 = ~(n5447 ^ n2367);
assign n7226 = n6011 | n13105;
assign n5035 = ~n13040;
assign n474 = ~(n11930 ^ n9316);
assign n12766 = n595 | n3221;
assign n7660 = ~(n1490 ^ n54);
assign n1854 = n3017 & n6921;
assign n12969 = ~n7229;
assign n7731 = n6638 | n1043;
assign n2156 = n10000 | n10534;
assign n1505 = ~n7779;
assign n7238 = n4957 ^ n8452;
assign n10441 = ~(n17 | n11460);
assign n12486 = ~(n10502 ^ n7617);
assign n8140 = ~(n11765 ^ n8851);
assign n12959 = ~n10770;
assign n249 = n1680 | n451;
assign n1415 = ~(n3434 ^ n5211);
assign n4936 = n2623;
assign n10923 = n1378 & n9835;
assign n7689 = n12757 | n225;
assign n6557 = ~n8332;
assign n4908 = n6668 & n10451;
assign n12433 = n7575 | n6624;
assign n796 = ~(n12506 ^ n4631);
assign n10821 = n7857 & n1396;
assign n4763 = ~(n9555 | n1830);
assign n1224 = ~(n2166 | n3862);
assign n899 = ~n9187;
assign n467 = ~n10572;
assign n7269 = n822 | n11176;
assign n1278 = n5334 ^ n9215;
assign n4980 = ~n11634;
assign n2615 = n11051 & n7953;
assign n13132 = n1682 & n1306;
assign n10360 = n3302 & n8133;
assign n2920 = n12814 | n5740;
assign n8930 = ~(n484 | n7618);
assign n9599 = ~(n9853 ^ n12044);
assign n2933 = ~(n3589 | n7217);
assign n4253 = ~n10770;
assign n335 = ~(n688 | n9816);
assign n769 = ~(n10919 ^ n4765);
assign n9409 = n5441 | n4164;
assign n11041 = n7769 | n7162;
assign n4032 = ~(n6530 | n4950);
assign n12476 = ~(n10499 | n12269);
assign n1963 = ~n9204;
assign n9334 = n11381 | n1848;
assign n11081 = ~(n4800 | n2089);
assign n578 = ~n7959;
assign n4111 = n7772 & n12853;
assign n10249 = n944 & n1673;
assign n3588 = ~n6831;
assign n1272 = ~(n4325 ^ n1743);
assign n2754 = n2411 & n757;
assign n10112 = ~n10594;
assign n3104 = n11108 & n5731;
assign n9227 = ~(n9166 | n4284);
assign n6143 = n1609 ^ n8544;
assign n9009 = ~(n8215 | n270);
assign n9665 = ~(n7843 ^ n5151);
assign n12647 = n12316 | n11960;
assign n7342 = ~n9249;
assign n2104 = ~n1202;
assign n10901 = ~(n6559 | n8071);
assign n8142 = ~n1731;
assign n12564 = ~(n6338 ^ n9644);
assign n11141 = n759 & n12035;
assign n1367 = ~n3558;
assign n2100 = n9931 | n8348;
assign n3672 = ~(n7769 ^ n2959);
assign n8938 = n7201 | n10725;
assign n6323 = n9378 | n2632;
assign n8427 = ~(n7514 ^ n10305);
assign n10317 = ~(n1148 ^ n13003);
assign n8227 = ~(n7973 ^ n5014);
assign n7862 = n10256 | n9159;
assign n11123 = n1869 | n3981;
assign n11950 = ~n13058;
assign n12690 = ~(n12449 ^ n7104);
assign n11631 = ~(n3109 ^ n5275);
assign n6300 = n2767 | n10584;
assign n2171 = ~(n8847 | n3007);
assign n6404 = n5041;
assign n9616 = ~(n1669 ^ n4820);
assign n8369 = ~(n12771 ^ n5813);
assign n4916 = n12411 | n4745;
assign n8937 = ~(n4690 ^ n11435);
assign n13117 = ~n9531;
assign n3994 = ~(n12285 ^ n82);
assign n8486 = ~n12987;
assign n7340 = n10929 | n12273;
assign n5453 = ~(n1245 ^ n6386);
assign n8485 = ~n4798;
assign n91 = n6796 & n8984;
assign n6210 = ~n13201;
assign n12267 = n5554 & n11321;
assign n10105 = ~n9125;
assign n9062 = n12626 & n1562;
assign n12212 = ~n3448;
assign n6 = ~(n5791 | n2517);
assign n1341 = ~(n8654 ^ n2457);
assign n13072 = n10977 | n4230;
assign n12608 = ~(n4649 | n10866);
assign n5345 = ~(n5206 | n9789);
assign n6872 = ~(n3828 ^ n4566);
assign n358 = ~(n530 ^ n1022);
assign n3279 = n2474 | n12017;
assign n12762 = n785 | n8534;
assign n8359 = n6341 & n9244;
assign n4477 = ~(n9824 ^ n13078);
assign n11343 = n11929 | n2958;
assign n1830 = n6873 & n7555;
assign n6682 = ~(n3599 ^ n773);
assign n3508 = ~n7702;
assign n5594 = ~(n7296 ^ n12546);
assign n958 = ~n13065;
assign n698 = n4114 & n510;
assign n7383 = n1672 & n6321;
assign n6611 = n12324 | n4724;
assign n2841 = n11771 & n128;
assign n7246 = ~(n8055 ^ n712);
assign n5667 = ~n9906;
assign n1623 = n6228 & n12774;
assign n8170 = n6630 | n8005;
assign n5612 = ~(n5140 | n6791);
assign n10447 = ~n4006;
assign n5276 = ~(n11301 ^ n5444);
assign n4898 = n12465 | n644;
assign n12562 = ~(n5052 ^ n11325);
assign n4156 = n5044 ^ n1444;
assign n12409 = ~(n3905 ^ n9111);
assign n6274 = ~n10560;
assign n11684 = n9148 & n282;
assign n464 = ~n11448;
assign n9645 = n18 | n6732;
assign n12898 = ~(n5558 ^ n9941);
assign n3133 = n6541 & n9519;
assign n6643 = n153 & n9996;
assign n8590 = n2057 & n1198;
assign n4259 = n5559 & n1526;
assign n1305 = n9318 | n10532;
assign n10671 = n8925 & n2930;
assign n9104 = n11170 | n5575;
assign n2080 = ~n7812;
assign n3208 = ~n9846;
assign n2780 = ~(n8338 | n4200);
assign n2441 = ~n3097;
assign n9812 = n13009 & n7105;
assign n6002 = ~(n10133 | n8052);
assign n639 = n1050 & n11728;
assign n3560 = n9868 | n7846;
assign n5647 = n11807 & n1366;
assign n3938 = n8720 | n1554;
assign n947 = ~n11324;
assign n10563 = n10770 & n3769;
assign n5639 = n495 | n6853;
assign n2090 = n947 | n11950;
assign n11622 = ~(n8994 ^ n6847);
assign n1694 = ~(n10167 | n11158);
assign n5855 = n7852 | n1449;
assign n5238 = n3032 | n12244;
assign n1550 = n9867 | n5076;
assign n4476 = ~(n3358 ^ n5927);
assign n1429 = ~(n8180 | n2667);
assign n11658 = ~(n2248 ^ n462);
assign n619 = n8919 | n8549;
assign n10258 = ~n9875;
assign n9189 = ~(n10945 ^ n3969);
assign n3245 = n4491 | n11592;
assign n8965 = n2773 & n6380;
assign n9529 = n11864 | n8079;
assign n12130 = n6968 | n10761;
assign n12836 = ~(n13037 ^ n12865);
assign n6779 = ~(n1839 | n7182);
assign n8755 = ~n2393;
assign n5956 = n8249 | n7723;
assign n8430 = n1082 | n12258;
assign n12580 = n12837 | n4230;
assign n6731 = ~n10809;
assign n457 = n2941 | n9822;
assign n2138 = ~(n1068 ^ n11538);
assign n3548 = ~(n9775 ^ n4282);
assign n4250 = n2284 & n8770;
assign n848 = ~n1569;
assign n9726 = ~(n2359 ^ n4871);
assign n7319 = n3805 | n2675;
assign n4109 = ~(n9838 | n12943);
assign n12591 = ~(n10310 ^ n12414);
assign n2733 = ~(n12272 | n10455);
assign n11280 = ~(n8285 ^ n5481);
assign n7096 = n3572 | n9080;
assign n9955 = n5306 | n12544;
assign n7631 = ~(n7648 | n11208);
assign n8941 = ~n4335;
assign n11240 = n9035 | n3794;
assign n1745 = n3104 | n11093;
assign n8956 = n8277 | n2337;
assign n9232 = n2136 & n13069;
assign n1201 = ~(n2925 ^ n4583);
assign n2016 = ~(n10152 ^ n8810);
assign n7834 = n4530 & n7256;
assign n957 = ~(n3984 ^ n12964);
assign n9367 = n1064 & n12952;
assign n7897 = n6271 | n8754;
assign n12488 = ~(n1535 ^ n5775);
assign n1747 = n542 | n1570;
assign n8406 = n2705 | n5387;
assign n13212 = n7396 | n7723;
assign n1659 = ~n11327;
assign n5747 = ~(n6537 ^ n7670);
assign n2536 = ~n6917;
assign n10611 = n10795 | n5992;
assign n2707 = n3684 & n11672;
assign n7562 = n5696 & n538;
assign n11425 = n6512 & n11189;
assign n919 = n11240 & n2322;
assign n6547 = n7098 & n9349;
assign n9538 = ~n5995;
assign n6439 = ~n8233;
assign n10030 = n12455 & n12161;
assign n10582 = n5343 & n2821;
assign n1960 = ~(n7340 ^ n9287);
assign n3617 = n3255 | n6823;
assign n9011 = n368 & n10839;
assign n5504 = n7772 & n9093;
assign n5231 = n3225 | n1570;
assign n7152 = ~n3815;
assign n2669 = ~n2174;
assign n10688 = ~(n3191 ^ n8588);
assign n3343 = n4961 | n7292;
assign n10253 = n126 & n5783;
assign n6606 = ~n10785;
assign n8457 = n6846 | n8534;
assign n7108 = n12711 | n11259;
assign n8452 = n8228 & n5962;
assign n3647 = n10761 | n7935;
assign n8754 = ~n2590;
assign n606 = ~(n5441 ^ n4164);
assign n915 = ~(n1028 ^ n3425);
assign n12326 = n12558 | n11397;
assign n2513 = n12304 & n12574;
assign n4526 = ~(n10317 ^ n3023);
assign n3176 = n2402 & n12451;
assign n11597 = n1634 | n12997;
assign n1458 = n5452 & n12681;
assign n2906 = ~(n13110 ^ n5005);
assign n6075 = ~(n11500 ^ n4769);
assign n7237 = ~(n3776 ^ n1551);
assign n146 = ~n4579;
assign n8631 = ~n12091;
assign n10491 = n5839 | n1346;
assign n352 = n7621 | n2077;
assign n11400 = ~n12260;
assign n8774 = ~(n6436 ^ n6735);
assign n4947 = n9709;
assign n11770 = ~(n9621 | n7888);
assign n7300 = n11210 | n2116;
assign n1426 = n12371 & n12297;
assign n10084 = ~(n10358 ^ n3574);
assign n4481 = ~n3579;
assign n3252 = ~(n8369 ^ n3286);
assign n9979 = ~(n6233 ^ n5598);
assign n1266 = ~(n1797 ^ n4676);
assign n627 = n5134 & n6311;
assign n2245 = ~(n9763 | n11812);
assign n5615 = n6639 & n12031;
assign n10601 = n9484 & n2842;
assign n8241 = ~(n9597 ^ n7531);
assign n8881 = n2095 | n2599;
assign n10368 = n5395 | n7915;
assign n10779 = ~(n7378 ^ n3202);
assign n863 = n7263 & n12492;
assign n10802 = ~(n13231 ^ n7644);
assign n6326 = n1456 & n11610;
assign n11827 = n12090 | n2611;
assign n10857 = n6590 | n10029;
assign n768 = n633 | n1600;
assign n8320 = ~(n7355 ^ n9259);
assign n1892 = n8129 | n10319;
assign n4228 = ~(n4015 | n7465);
assign n12268 = ~(n2403 | n11348);
assign n1645 = n6110 | n5691;
assign n7173 = ~(n6165 ^ n2448);
assign n5305 = n863 | n7559;
assign n4815 = ~n6017;
assign n2778 = n2955 | n8145;
assign n674 = n8325 | n7221;
assign n6063 = ~n6655;
assign n1969 = ~(n10406 ^ n11126);
assign n13236 = ~(n88 ^ n11411);
assign n8602 = n7917 & n2049;
assign n5302 = ~(n661 ^ n1036);
assign n13235 = ~n2948;
assign n2775 = ~(n3977 ^ n7175);
assign n10974 = ~n1916;
assign n7819 = ~n12352;
assign n12508 = ~n9151;
assign n7477 = ~(n7091 ^ n10440);
assign n9368 = ~(n10876 ^ n6645);
assign n7384 = ~(n4586 ^ n1431);
assign n4647 = ~(n9997 ^ n9387);
assign n8367 = ~(n3511 | n11738);
assign n10034 = n10230 & n8525;
assign n5064 = ~(n930 ^ n2055);
assign n321 = ~n6826;
assign n568 = n6190 | n1861;
assign n7646 = ~(n7399 ^ n11984);
assign n6614 = n4980 | n10179;
assign n11890 = n7772 & n4470;
assign n13063 = ~n3499;
assign n9749 = n5752 & n2177;
assign n6170 = n5697 & n10636;
assign n9129 = ~n817;
assign n4037 = ~(n12889 ^ n171);
assign n9713 = ~(n5112 | n1180);
assign n3542 = ~(n8901 ^ n11552);
assign n4830 = ~n6920;
assign n3259 = ~n5969;
assign n7801 = n10571 | n1107;
assign n12781 = n511 & n12162;
assign n248 = n8349 | n12823;
assign n11178 = n2590 & n6392;
assign n8362 = ~(n495 ^ n461);
assign n8600 = n8263 & n2988;
assign n9621 = n12348 & n854;
assign n9882 = ~n5536;
assign n12213 = n766 | n129;
assign n4600 = n787 | n9223;
assign n12802 = n4832 & n820;
assign n11920 = ~n8506;
assign n12698 = ~n2389;
assign n3505 = ~n12965;
assign n9016 = ~n8332;
assign n8182 = n2449 | n6265;
assign n4509 = n5671 & n510;
assign n8223 = n6245 | n2449;
assign n7236 = ~(n8418 ^ n1260);
assign n6620 = ~(n1752 ^ n12367);
assign n5778 = ~(n7725 ^ n13023);
assign n9876 = ~(n216 ^ n3772);
assign n2286 = ~(n1409 ^ n5657);
assign n338 = ~n12853;
assign n4041 = n8079 | n542;
assign n11828 = n2478 & n10715;
assign n4306 = n8254 | n12789;
assign n6499 = ~n7270;
assign n5798 = ~(n3183 ^ n11445);
assign n12519 = n12689 & n4103;
assign n12299 = ~(n11189 | n6512);
assign n2845 = ~(n1365 ^ n11162);
assign n4126 = ~(n10366 ^ n12474);
assign n3918 = n8168 & n12944;
assign n3877 = ~(n8689 | n8630);
assign n8680 = n6957 | n9370;
assign n1354 = ~n6023;
assign n4939 = n8796 | n10214;
assign n7335 = n4108 & n3554;
assign n2506 = n10908 & n411;
assign n9913 = ~n7812;
assign n4035 = ~(n11812 ^ n1066);
assign n10599 = n8463 | n12655;
assign n7995 = ~(n5622 | n10531);
assign n2347 = ~(n2653 | n13111);
assign n10559 = ~(n12993 ^ n6589);
assign n1909 = ~(n4245 ^ n5866);
assign n2258 = ~(n8953 ^ n10930);
assign n8598 = ~n499;
assign n7367 = ~(n3612 ^ n9312);
assign n1397 = ~(n8349 ^ n10121);
assign n678 = ~(n5056 ^ n2819);
assign n8720 = ~n10162;
assign n11667 = ~(n11826 ^ n8353);
assign n5410 = ~(n6108 | n4091);
assign n11486 = ~(n4049 | n11161);
assign n2836 = ~(n3660 ^ n8958);
assign n6130 = n10143 | n13238;
assign n10730 = ~n9528;
assign n7147 = n6825 & n6467;
assign n9139 = ~(n5774 ^ n2236);
assign n11335 = ~(n11652 ^ n1446);
assign n2646 = ~(n3310 ^ n4909);
assign n6738 = n202 | n10106;
assign n307 = n5520 | n542;
assign n2328 = ~(n4679 ^ n8085);
assign n3788 = ~(n1475 ^ n12489);
assign n9322 = ~(n4810 ^ n3936);
assign n1687 = n2057 & n2295;
assign n7151 = n1136 | n716;
assign n10553 = ~(n12936 ^ n7312);
assign n3423 = n119 | n6404;
assign n7866 = n6764 & n13138;
assign n4420 = ~n10642;
assign n10061 = ~(n11820 ^ n9979);
assign n751 = ~(n5868 ^ n5805);
assign n10909 = n12775 & n4359;
assign n10580 = ~(n9856 | n6101);
assign n5181 = n8858 & n8194;
assign n12250 = n8557 & n12756;
assign n6458 = ~(n1087 ^ n9546);
assign n4263 = ~(n10853 ^ n1311);
assign n4791 = n5028 | n2735;
assign n8153 = ~n8459;
assign n12366 = ~(n9833 | n5746);
assign n9805 = n10034 ^ n2951;
assign n11191 = n11677 | n2572;
assign n4031 = ~(n12984 ^ n9646);
assign n10470 = ~n11885;
assign n7277 = n1331 | n11107;
assign n2464 = n3854 | n11668;
assign n4511 = ~(n4552 ^ n3324);
assign n3968 = n9940 & n8397;
assign n4028 = ~n7792;
assign n9365 = n13084 | n479;
assign n10700 = n5794 | n3512;
assign n4161 = ~n287;
assign n5669 = n5168 | n11107;
assign n73 = n3129 | n3143;
assign n5954 = ~n1978;
assign n6221 = ~(n1745 ^ n3349);
assign n10709 = ~(n368 ^ n5891);
assign n506 = ~(n3314 ^ n9583);
assign n2142 = ~(n5621 ^ n3043);
assign n1907 = n10835 | n10843;
assign n9359 = ~(n8627 ^ n12694);
assign n6597 = ~(n8573 ^ n12096);
assign n9076 = n7506 & n10543;
assign n9049 = n10626 & n8271;
assign n5688 = ~n4748;
assign n12360 = n11115 & n2509;
assign n11331 = ~n2751;
assign n789 = ~n9216;
assign n11277 = ~(n12577 | n2055);
assign n7805 = ~n13058;
assign n12214 = ~(n12260 ^ n3142);
assign n1096 = n9668 | n10886;
assign n1256 = n1058 | n3817;
assign n13080 = ~n5556;
assign n8151 = ~(n6964 ^ n4539);
assign n6685 = n10263 | n7221;
assign n4347 = ~(n1306 ^ n7753);
assign n4376 = n6040 | n10179;
assign n8805 = n8410 ^ n10800;
assign n6758 = n8308 & n4330;
assign n2670 = ~n10103;
assign n6759 = ~(n2638 ^ n415);
assign n4096 = n2527 | n2030;
assign n12473 = ~(n7299 ^ n4082);
assign n12682 = n3225 | n6041;
assign n626 = n2889 | n121;
assign n8240 = n6419 | n11107;
assign n1639 = n3982 | n752;
assign n7310 = n9383 | n2958;
assign n7271 = n10400 | n8348;
assign n13068 = n1235 | n8673;
assign n11552 = n12416 | n10029;
assign n9087 = ~(n2948 ^ n8155);
assign n12150 = n3866 | n2675;
assign n10160 = n6438 | n7530;
assign n7431 = ~(n4304 ^ n11885);
assign n11842 = ~n10615;
assign n6027 = ~(n11896 ^ n7120);
assign n8216 = n3302 | n8133;
assign n13181 = ~n937;
assign n244 = ~(n13093 | n4338);
assign n349 = n9919 | n6635;
assign n4523 = n2520 & n255;
assign n934 = n5914 | n3356;
assign n10208 = n11628 | n8563;
assign n5316 = ~(n5943 ^ n12929);
assign n5019 = ~(n12422 | n10198);
assign n7390 = n1214 | n9418;
assign n6968 = ~n3669;
assign n5971 = ~n11766;
assign n3282 = n11319 | n4067;
assign n9195 = n11418;
assign n8131 = ~n2252;
assign n84 = n6503 & n310;
assign n136 = n9339 | n10029;
assign n7261 = n10136 | n3174;
assign n2267 = n5835 | n3488;
assign n3903 = n5586 & n3832;
assign n8371 = ~(n229 | n651);
assign n11975 = ~n11288;
assign n5735 = ~(n6566 ^ n6969);
assign n6451 = n13106 ^ n7447;
assign n9219 = ~(n3711 ^ n8294);
assign n11268 = ~(n10254 | n4730);
assign n1034 = ~(n1835 ^ n11349);
assign n10953 = ~(n12259 | n3048);
assign n10228 = n122 | n6062;
assign n11893 = n12614 ^ n864;
assign n3991 = ~(n404 ^ n6759);
assign n8418 = n8790 & n10312;
assign n8235 = n5954 & n3168;
assign n11375 = n2677 & n10912;
assign n2878 = ~(n9387 | n9997);
assign n6721 = ~n11891;
assign n6853 = n1779 & n10132;
assign n1087 = n7234 | n8702;
assign n530 = ~n4987;
assign n12793 = n6191 | n1894;
assign n8339 = ~n11559;
assign n2864 = ~(n2100 ^ n12220);
assign n670 = n1220 & n3878;
assign n12038 = ~(n664 ^ n3968);
assign n6955 = ~(n3265 ^ n1433);
assign n7818 = ~(n9065 ^ n3332);
assign n1239 = n12281 & n1698;
assign n5959 = ~n7806;
assign n10002 = n9732 & n854;
assign n3732 = n6414 & n12770;
assign n7946 = n8327 | n3374;
assign n13023 = n7022 & n3656;
assign n9746 = ~(n10395 ^ n102);
assign n8357 = ~(n10294 ^ n8283);
assign n10613 = ~(n10549 ^ n3693);
assign n10949 = n406 | n7998;
assign n7281 = n11218 | n2059;
assign n2697 = ~(n10475 ^ n7021);
assign n6340 = ~(n10718 ^ n10124);
assign n9223 = n12954;
assign n10723 = ~(n12152 | n7735);
assign n2224 = n12754 | n11714;
assign n10849 = ~n12822;
assign n10767 = ~(n9101 ^ n2214);
assign n125 = n9039 | n10466;
assign n2465 = n3361 ^ n4908;
assign n1146 = ~(n5727 ^ n13175);
assign n3983 = n11352 | n10029;
assign n1466 = n12613 & n375;
assign n13158 = ~(n12296 ^ n10096);
assign n4438 = n12493 | n11668;
assign n10027 = ~(n6992 ^ n10297);
assign n7308 = ~(n9240 ^ n10659);
assign n3911 = ~n11180;
assign n12913 = n121 | n4960;
assign n8498 = ~n10162;
assign n3244 = ~(n1524 ^ n6873);
assign n6509 = n13168 | n2544;
assign n12981 = ~(n8085 | n4679);
assign n3028 = n75 | n8024;
assign n11249 = n7970 | n3075;
assign n4329 = ~(n8273 ^ n4156);
assign n11606 = n9199 & n11192;
assign n12938 = n3489 | n3715;
assign n10364 = n9987 & n7901;
assign n10917 = ~(n6240 ^ n7211);
assign n11024 = n11514 | n8777;
assign n984 = ~(n3123 ^ n9212);
assign n2182 = n1515 | n7004;
assign n4233 = ~(n11133 ^ n1291);
assign n707 = ~(n2811 ^ n11250);
assign n13210 = n11704 & n2348;
assign n7610 = n3636 & n10341;
assign n8342 = ~(n2476 | n2510);
assign n6182 = ~n6937;
assign n1450 = ~(n2616 | n5285);
assign n1058 = ~n510;
assign n1030 = ~n4017;
assign n9160 = ~n12892;
assign n2460 = ~(n9099 ^ n245);
assign n11202 = n11236 & n411;
assign n1936 = ~n3566;
assign n7634 = n5733 | n10474;
assign n2960 = n7038 | n1833;
assign n13090 = n10112 | n5076;
assign n8282 = ~(n11804 ^ n4548);
assign n6328 = ~(n2659 ^ n2736);
assign n11086 = n1747 & n11423;
assign n12118 = ~(n7637 ^ n5038);
assign n11493 = n10857 | n8793;
assign n9002 = ~(n10796 | n12058);
assign n5078 = ~(n8292 ^ n13090);
assign n9238 = ~n469;
assign n2684 = ~(n12974 ^ n10038);
assign n3862 = n5490 & n10740;
assign n5075 = ~(n9324 ^ n4090);
assign n1840 = ~(n12873 | n8756);
assign n6844 = n1323 | n12062;
assign n258 = n3019 & n11987;
assign n1990 = n2899 | n11910;
assign n4631 = ~(n1276 ^ n184);
assign n507 = n2243 & n4311;
assign n2546 = n7056 & n7432;
assign n6688 = n12032 | n8490;
assign n7223 = ~n3677;
assign n8352 = n2530 & n12473;
assign n6422 = n6881 | n10702;
assign n9146 = n13190 | n206;
assign n1875 = n4135 ^ n12612;
assign n11330 = n9698 | n4023;
assign n10989 = ~n12939;
assign n10013 = n9429 | n4640;
assign n1371 = n6934 & n3871;
assign n2875 = ~n11537;
assign n12525 = n7566 | n2766;
assign n1885 = ~n3977;
assign n11172 = ~n4102;
assign n5970 = ~n5786;
assign n10823 = n3957 & n11273;
assign n11372 = n2449 | n8490;
assign n7158 = ~n6085;
assign n4508 = n8974 & n10726;
assign n2981 = ~(n1373 ^ n10721);
assign n7153 = n7073 & n1477;
assign n5132 = n10527 | n11107;
assign n12624 = ~n10238;
assign n2976 = ~(n9502 ^ n2719);
assign n8374 = ~n510;
assign n5686 = ~(n4171 ^ n5173);
assign n7077 = ~(n8279 | n802);
assign n145 = n12058 & n10796;
assign n9575 = n11996 & n12650;
assign n7670 = ~(n2006 ^ n6325);
assign n10741 = n12775 | n4359;
assign n12715 = ~(n10671 ^ n1927);
assign n12934 = n1791 & n1886;
assign n9067 = n11614 & n3536;
assign n7247 = ~n5470;
assign n373 = n10824 | n9923;
assign n7137 = n4361 & n4563;
assign n11021 = n3458 & n4475;
assign n8643 = ~(n8923 | n7479);
assign n9804 = ~n11567;
assign n1438 = ~n10594;
assign n2162 = n1513 | n2298;
assign n5489 = ~n5590;
assign n7886 = n12353 | n8316;
assign n10370 = n6231 | n12273;
assign n4120 = ~(n10155 ^ n11080);
assign n2459 = ~(n2854 ^ n2853);
assign n8541 = n10897 | n1856;
assign n10502 = n8664 & n10161;
assign n3474 = ~(n4538 | n12450);
assign n1145 = ~n4681;
assign n10555 = n2614 | n5076;
assign n4044 = n6823 & n3255;
assign n5753 = n11515 & n1542;
assign n3574 = ~(n3131 | n7627);
assign n1734 = ~(n4706 ^ n7851);
assign n10305 = ~n7778;
assign n7037 = n10608 | n3618;
assign n11935 = ~(n10282 | n5859);
assign n6160 = ~n3774;
assign n11476 = n8384 | n10098;
assign n11912 = ~(n10328 | n10366);
assign n5889 = n5773 & n12600;
assign n5524 = n8120 & n9334;
assign n12102 = n3110 ^ n7083;
assign n6607 = n6046 & n2333;
assign n4637 = ~(n6844 | n11085);
assign n7612 = n845 | n9075;
assign n3699 = n6506 | n7865;
assign n10463 = ~(n12850 ^ n2632);
assign n9179 = ~(n3387 | n12115);
assign n2501 = n10997 & n3996;
assign n9982 = ~(n6075 ^ n10821);
assign n11379 = ~n8291;
assign n10948 = ~n10172;
assign n12660 = n11982 | n10764;
assign n1753 = ~(n4489 ^ n10968);
assign n8932 = n2757 | n6001;
assign n6254 = n6769 | n12388;
assign n12713 = ~n10378;
assign n9950 = ~(n5371 ^ n2441);
assign n5836 = ~(n7527 | n8913);
assign n11910 = ~n951;
assign n6105 = ~(n544 ^ n6025);
assign n5975 = ~(n5497 ^ n1387);
assign n10404 = ~(n5998 | n3173);
assign n7656 = n7415 & n3436;
assign n337 = n3647 | n5098;
assign n8031 = ~(n2798 ^ n4670);
assign n1842 = n4808 | n8534;
assign n2280 = n10422 & n12773;
assign n12659 = n10471 | n5242;
assign n3056 = n3900 | n5443;
assign n4712 = ~(n7534 ^ n7212);
assign n7086 = ~n8824;
assign n2891 = n2471 & n165;
assign n11348 = ~(n2475 ^ n9574);
assign n5963 = n1261 | n7935;
assign n1735 = n6770 | n10319;
assign n5853 = ~n5140;
assign n7948 = ~(n1368 ^ n10042);
assign n12588 = ~(n215 | n10629);
assign n2577 = ~(n11845 ^ n7057);
assign n7858 = ~(n3480 ^ n2859);
assign n1046 = n3539 & n12446;
assign n2565 = ~(n3980 ^ n3714);
assign n297 = n6517 | n6493;
assign n12720 = n4166 | n1570;
assign n215 = ~(n2024 | n6508);
assign n10994 = n1989 | n6770;
assign n1986 = n10889 & n10498;
assign n4720 = n9637 | n5188;
assign n12184 = n7783 | n6265;
assign n7393 = ~(n4345 ^ n12570);
assign n11237 = ~n6701;
assign n2287 = ~n8230;
assign n5232 = ~(n7896 ^ n851);
assign n4498 = ~n5546;
assign n9151 = n4638 & n7453;
assign n1434 = ~n8332;
assign n9704 = n867 & n9326;
assign n1876 = n11548 | n1985;
assign n3817 = ~n2590;
assign n3455 = ~(n4600 ^ n1723);
assign n12631 = ~(n7439 | n10963);
assign n6819 = ~(n12845 ^ n13087);
assign n6880 = n13039 | n2133;
assign n5976 = n1875 | n12366;
assign n2403 = ~n13121;
assign n12400 = ~(n1774 | n8413);
assign n13155 = ~(n10547 ^ n7689);
assign n9897 = ~n4126;
assign n12832 = n3662 & n6664;
assign n12427 = n3091 | n2083;
assign n1579 = ~n10075;
assign n12838 = ~n10582;
assign n7377 = ~n5962;
assign n3692 = n13025 | n2059;
assign n10872 = ~n4906;
assign n12179 = n11779 | n7254;
assign n11306 = ~(n5357 ^ n3887);
assign n713 = ~n6647;
assign n5577 = n9564 | n5029;
assign n6007 = ~(n6388 ^ n6243);
assign n236 = ~(n1334 ^ n11176);
assign n1309 = ~(n9066 ^ n7681);
assign n9172 = ~n2073;
assign n5072 = n9069 | n8268;
assign n4349 = n4376 ^ n11813;
assign n1844 = ~(n7754 ^ n775);
assign n12598 = ~(n9922 ^ n6031);
assign n12439 = ~(n9083 ^ n4390);
assign n5554 = ~n748;
assign n5001 = ~n8559;
assign n5693 = n12573 | n4640;
assign n9579 = ~(n6079 ^ n1293);
assign n11353 = ~(n7067 ^ n5979);
assign n6976 = n6657 | n265;
assign n8897 = ~(n5693 ^ n667);
assign n12535 = ~n4042;
assign n384 = ~(n12933 ^ n6158);
assign n1452 = n8610 & n12521;
assign n7004 = ~(n2251 | n665);
assign n932 = n5655 | n2206;
assign n5666 = ~n6392;
assign n1035 = ~n353;
assign n1603 = n3570 & n7898;
assign n10281 = ~n1650;
assign n4535 = ~(n300 ^ n10619);
assign n6677 = n6956 ^ n2583;
assign n451 = n11779 | n4640;
assign n11031 = ~(n5421 ^ n11806);
assign n11405 = ~(n3747 ^ n999);
assign n8093 = n3550 | n5059;
assign n13133 = ~n7465;
assign n4353 = n1867 & n1448;
assign n11459 = n161 | n12328;
assign n557 = ~(n12448 ^ n7838);
assign n6652 = ~n4645;
assign n3861 = ~n3913;
assign n10551 = n10094 & n147;
assign n5645 = ~n10805;
assign n2087 = ~(n9797 | n12584);
assign n3296 = ~(n7891 ^ n6693);
assign n315 = n12585 & n6315;
assign n6678 = ~(n12235 ^ n1253);
assign n9800 = ~(n5933 ^ n6670);
assign n12953 = n1035 | n6732;
assign n4261 = n4974 | n5076;
assign n1654 = n3587 | n4947;
assign n7279 = n8139 & n10606;
assign n8520 = n3316 & n5411;
assign n11273 = n2639 | n8490;
assign n5206 = n9131 | n10871;
assign n8165 = n2109 | n488;
assign n6716 = ~n68;
assign n4180 = n983 | n9177;
assign n7914 = ~n8818;
assign n4930 = n8335 | n2675;
assign n1282 = ~(n11556 ^ n3745);
assign n6664 = n12241 | n9055;
assign n9136 = ~(n9565 ^ n4597);
assign n735 = ~n1528;
assign n4314 = n4610 | n479;
assign n12166 = ~n11324;
assign n6443 = ~(n12167 | n2927);
assign n7290 = n72 ^ n9250;
assign n3113 = n7780 | n1144;
assign n8099 = ~(n5327 | n4421);
assign n11959 = n1311 & n10853;
assign n67 = ~(n3899 ^ n4195);
assign n7935 = n9558;
assign n1373 = n8727 | n6824;
assign n8829 = n2236 | n5774;
assign n10577 = n13028 | n6173;
assign n1695 = ~n7720;
assign n10151 = ~(n13188 ^ n1288);
assign n2042 = ~(n2486 | n979);
assign n7480 = ~n11129;
assign n10021 = ~n11891;
assign n5564 = n11099 | n10689;
assign n9152 = n10688 | n10759;
assign n2890 = ~n13058;
assign n11366 = n6751 | n1463;
assign n6078 = ~(n8476 | n10027);
assign n3999 = ~n5962;
assign n5690 = ~(n7457 | n3117);
assign n10586 = ~n11411;
assign n11971 = ~(n11199 ^ n4601);
assign n7244 = n5166 & n10536;
assign n1601 = n5616 | n4055;
assign n3810 = ~(n5763 ^ n459);
assign n4670 = ~(n7265 ^ n12100);
assign n12054 = n8715 ^ n6921;
assign n8873 = n3802 | n12189;
assign n1493 = ~n2169;
assign n5556 = n9904 ^ n12915;
assign n8090 = n9079 & n920;
assign n8537 = n5090 & n7638;
assign n7744 = ~(n1262 ^ n5235);
assign n10941 = ~n8422;
assign n12573 = ~n11891;
assign n12377 = ~n8798;
assign n10478 = ~(n5556 ^ n6073);
assign n272 = n9399 | n13031;
assign n3060 = n11790 | n7574;
assign n9681 = ~n12810;
assign n1369 = ~(n2289 ^ n4569);
assign n10145 = n8457 | n9972;
assign n9287 = n6922 | n6635;
assign n8171 = n10287 | n12847;
assign n12652 = n1447 | n6404;
assign n4586 = ~(n1233 ^ n10632);
assign n1291 = ~(n941 ^ n4071);
assign n6302 = n6383 | n1570;
assign n4203 = ~n9841;
assign n1334 = ~(n6167 ^ n5981);
assign n11695 = ~(n1742 | n8475);
assign n11813 = n8466 & n8506;
assign n13120 = ~(n7752 ^ n9274);
assign n4795 = n5561 | n2315;
assign n3687 = n3331 | n952;
assign n5266 = ~(n13040 ^ n859);
assign n12309 = n10492 | n6138;
assign n8769 = n9298 | n8127;
assign n4542 = n10929 | n7723;
assign n8437 = n204 & n5572;
assign n8752 = ~(n5546 ^ n13044);
assign n8780 = n8329 | n5797;
assign n10315 = n980 & n11297;
assign n2717 = ~n10541;
assign n5387 = n842 & n4274;
assign n3515 = n946 | n12501;
assign n6282 = ~(n1206 ^ n2714);
assign n612 = ~(n2743 | n1620);
assign n7320 = n8142 & n4443;
assign n12047 = n8759 | n13148;
assign n4112 = n6495 & n12315;
assign n6174 = ~(n12151 ^ n12540);
assign n9924 = n5271 | n6404;
assign n3001 = n10411 | n4208;
assign n1194 = ~n8163;
assign n5464 = ~(n12638 ^ n736);
assign n7578 = ~(n8538 | n12200);
assign n7188 = ~n510;
assign n11472 = ~(n5913 ^ n10379);
assign n13173 = n761 & n3085;
assign n8693 = ~n5307;
assign n5793 = n5107 | n119;
assign n12756 = n8123 & n3373;
assign n8945 = ~(n3578 ^ n4766);
assign n4633 = ~(n12127 | n5196);
assign n6732 = n8160;
assign n8483 = ~(n3397 ^ n11459);
assign n7361 = n6205 | n425;
assign n891 = n12629 | n4936;
assign n1306 = n12576 & n7817;
assign n7084 = ~n817;
assign n8573 = ~(n12485 ^ n1309);
assign n9690 = n11499 | n10909;
assign n9584 = n9499 | n1381;
assign n1437 = ~n11376;
assign n2331 = n5809 | n9759;
assign n7883 = ~n10620;
assign n3256 = n3295 | n4751;
assign n1463 = n3058;
assign n1403 = ~(n10324 ^ n7202);
assign n13050 = ~(n9863 ^ n11128);
assign n11628 = ~n5920;
assign n134 = ~(n68 ^ n6246);
assign n669 = ~(n8972 ^ n6125);
assign n7698 = ~(n2340 ^ n1386);
assign n6496 = n7629 & n3197;
assign n5361 = n11705 | n11893;
assign n9994 = n10714 | n10319;
assign n6427 = ~(n2372 ^ n9785);
assign n823 = ~(n12660 ^ n6435);
assign n8317 = ~n3379;
assign n11992 = ~(n9037 ^ n7599);
assign n12998 = ~n10873;
assign n757 = ~n4417;
assign n10475 = ~(n11676 ^ n2483);
assign n11143 = ~n8564;
assign n9140 = n6384 | n10417;
assign n5452 = n12786 | n8268;
assign n8387 = n10590 & n10483;
assign n956 = ~n10451;
assign n8762 = n8728 & n4518;
assign n10630 = ~(n9466 ^ n13120);
assign n10728 = ~(n12356 ^ n3734);
assign n9986 = n3172 & n1773;
assign n4135 = n4465 | n4373;
assign n6119 = n7215 & n249;
assign n2115 = n692 & n12676;
assign n2129 = ~n8860;
assign n11641 = n7772 & n9531;
assign n11572 = ~(n8180 ^ n4872);
assign n9872 = ~(n259 ^ n10227);
assign n5736 = n2581 | n12328;
assign n12448 = n11757 | n8490;
assign n8585 = ~n2758;
assign n3142 = ~(n1608 ^ n12398);
assign n331 = n11054 | n12188;
assign n4326 = n8599 & n6468;
assign n9559 = n6112 | n7935;
assign n2502 = ~(n11022 ^ n3343);
assign n1473 = ~(n12390 ^ n1300);
assign n7676 = n4991 & n10066;
assign n774 = ~(n10949 ^ n7122);
assign n3947 = ~(n9956 ^ n10775);
assign n5523 = n4080 | n11300;
assign n11861 = ~(n4866 ^ n908);
assign n3268 = ~(n112 ^ n10003);
assign n6352 = n12114 & n2186;
assign n7296 = ~(n12601 ^ n9036);
assign n766 = ~(n9992 | n10630);
assign n5714 = ~n7183;
assign n4504 = ~(n8137 | n4740);
assign n11650 = n10381 | n7824;
assign n730 = n7272 | n3918;
assign n11555 = n5953 & n12712;
assign n10840 = ~(n6797 | n3294);
assign n7501 = n9304 & n6475;
assign n12176 = n1440 & n8741;
assign n7863 = ~(n888 ^ n2765);
assign n10512 = ~n3412;
assign n3447 = n1520 & n10145;
assign n6052 = ~n8319;
assign n8811 = n10577 ^ n3995;
assign n10898 = ~n1307;
assign n1798 = n11030 & n9531;
assign n5585 = ~(n5234 ^ n11201);
assign n7842 = ~(n10973 ^ n2761);
assign n8310 = n9626 | n130;
assign n13084 = ~n5884;
assign n5273 = ~(n12442 ^ n9839);
assign n3662 = n8102 | n5258;
assign n6670 = n1138 & n8125;
assign n9102 = n10545 | n11639;
assign n12074 = ~(n6823 ^ n9857);
assign n8999 = n3758 | n164;
assign n1113 = ~n4006;
assign n4554 = ~(n1877 | n1429);
assign n8975 = n6305 | n984;
assign n5472 = n9150 & n8743;
assign n7305 = n7566 & n2766;
assign n630 = n5307 & n4036;
assign n4618 = ~n10946;
assign n8916 = ~(n9648 ^ n955);
assign n8853 = n7523 | n7975;
assign n2651 = n9605 & n1054;
assign n2377 = n10260 & n5916;
assign n6714 = n1257 & n6845;
assign n7969 = n4875 | n12328;
assign n2874 = ~(n4578 ^ n4150);
assign n4708 = n906 & n2056;
assign n4178 = n12552 | n10213;
assign n5380 = ~(n10023 ^ n11042);
assign n1204 = ~(n5918 ^ n811);
assign n11700 = ~n7491;
assign n7797 = n11751 | n617;
assign n4247 = ~(n12321 ^ n5781);
assign n6659 = n8009 | n6628;
assign n3528 = n7049 | n8563;
assign n11945 = n3307 | n5566;
assign n11064 = ~(n2451 ^ n9034);
assign n8118 = n3822 & n3339;
assign n9819 = n8817 | n9159;
assign n13082 = ~n2174;
assign n1362 = ~(n4968 ^ n756);
assign n4475 = n13183 | n177;
assign n3666 = ~(n9269 ^ n515);
assign n4887 = ~(n12606 | n7020);
assign n5508 = n10452 | n6243;
assign n8491 = ~n10979;
assign n2489 = ~(n3959 | n4286);
assign n9077 = ~(n6852 ^ n6307);
assign n11494 = n9546 & n1087;
assign n3990 = ~(n3606 | n7869);
assign n6093 = n10351 & n8448;
assign n803 = ~n11990;
assign n9442 = n4855 | n10319;
assign n3418 = ~n3319;
assign n9847 = n8139 & n12965;
assign n10584 = n1741 | n9537;
assign n9668 = ~n6826;
assign n9114 = n7498 & n4225;
assign n6290 = ~n1421;
assign n12808 = ~n6607;
assign n927 = ~(n12784 ^ n6620);
assign n4158 = n1663 | n2415;
assign n6153 = ~(n5274 ^ n11296);
assign n10798 = ~n2295;
assign n8900 = ~n818;
assign n11326 = ~(n11414 ^ n12354);
assign n7847 = ~n10575;
assign n10587 = ~n5729;
assign n9777 = ~(n9796 ^ n2040);
assign n1399 = ~(n11125 ^ n10249);
assign n3746 = ~(n5711 ^ n6895);
assign n12193 = ~(n1137 ^ n6899);
assign n3148 = ~(n2053 | n7834);
assign n10538 = ~(n5509 ^ n12875);
assign n12257 = n8732 | n3882;
assign n11062 = ~(n10640 ^ n3382);
assign n12679 = n1634 | n9745;
assign n4792 = ~n10451;
assign n5764 = ~(n8008 ^ n12113);
assign n9215 = n5031 & n510;
assign n1624 = ~n5796;
assign n5055 = n5568 & n5729;
assign n3117 = n2582 | n2816;
assign n9411 = n6416 | n9075;
assign n8739 = ~n4978;
assign n9612 = n7748 | n4373;
assign n11561 = ~(n5306 ^ n7428);
assign n9196 = ~(n4263 ^ n11816);
assign n7156 = n8776 | n6769;
assign n2560 = ~(n2049 ^ n7917);
assign n4103 = n12236 | n4835;
assign n4629 = n6215 | n10433;
assign n4013 = ~n2057;
assign n2255 = n10248 & n5369;
assign n12725 = n5826 & n2831;
assign n7719 = ~n7439;
assign n5060 = ~(n9048 ^ n6105);
assign n3204 = n3634 | n1043;
assign n12569 = n11117 | n8445;
assign n3878 = n3176 | n10652;
assign n3696 = ~n1432;
assign n3937 = n4475 | n3458;
assign n5252 = n10153 | n3650;
assign n4711 = ~(n9955 ^ n3562);
assign n4303 = n1719 ^ n2423;
assign n2006 = n5671 & n8506;
assign n11995 = n3922 & n2428;
assign n1086 = ~(n31 ^ n8872);
assign n12964 = n11960 | n9075;
assign n2044 = ~(n5451 ^ n7569);
assign n9874 = ~(n6151 | n5033);
assign n6904 = ~(n11692 ^ n7309);
assign n7743 = n1087 | n9546;
assign n1002 = n1909 | n3955;
assign n7987 = n4739 | n4675;
assign n3923 = ~(n7875 ^ n4856);
assign n9131 = ~n1302;
assign n1865 = ~(n9423 | n3206);
assign n11786 = n7062 | n12273;
assign n12977 = ~(n11168 ^ n13105);
assign n6414 = n7042 | n9078;
assign n6525 = n803 & n8558;
assign n3889 = ~(n5678 ^ n8684);
assign n7009 = ~n10457;
assign n1697 = ~n1938;
assign n8428 = ~n10398;
assign n2574 = ~(n7529 | n7715);
assign n931 = n4564 | n3949;
assign n10071 = ~(n9903 ^ n3644);
assign n7309 = n542 | n11668;
assign n10995 = ~(n4057 ^ n10994);
assign n4450 = n6029 & n2179;
assign n10465 = ~n7659;
assign n11474 = ~(n7330 ^ n11760);
assign n5428 = n7142 | n6265;
assign n7556 = n812 & n9717;
assign n16 = ~n12348;
assign n7540 = ~(n8827 ^ n6378);
assign n3123 = ~(n10828 ^ n5651);
assign n807 = ~(n3274 ^ n49);
assign n6515 = n4908 & n11545;
assign n2544 = n8640;
assign n6034 = n1453 & n8216;
assign n10218 = ~(n2054 ^ n4575);
assign n10038 = n5893 & n3124;
assign n6407 = ~n834;
assign n4048 = ~(n8483 ^ n3881);
assign n10482 = n13071 & n2419;
assign n1864 = n6967 | n12328;
assign n8008 = n1511 | n1026;
assign n2146 = n1544 & n7611;
assign n8450 = ~(n5568 | n8308);
assign n13067 = n8020 | n7530;
assign n6891 = ~(n8141 ^ n11510);
assign n6695 = ~(n8559 ^ n1623);
assign n7618 = n80 | n1571;
assign n9433 = ~(n8224 ^ n7449);
assign n2234 = n2155 & n6291;
assign n6813 = n6587 | n2675;
assign n994 = n2188 & n3265;
assign n3434 = ~(n7038 ^ n10621);
assign n7398 = ~(n4210 ^ n1473);
assign n1497 = n7146 | n8030;
assign n6475 = n6244 | n9043;
assign n12747 = ~n11518;
assign n12103 = ~(n4393 ^ n4073);
assign n3402 = ~(n2360 ^ n9128);
assign n8575 = ~(n5494 | n9578);
assign n11672 = n3969 | n10945;
assign n2503 = n6566 | n155;
assign n11961 = ~(n2887 ^ n8244);
assign n5359 = ~n5030;
assign n11012 = ~(n3549 ^ n11151);
assign n9385 = ~(n3152 | n4815);
assign n397 = ~(n3401 ^ n1555);
assign n7415 = ~n1157;
assign n9306 = ~(n5292 | n8213);
assign n9180 = n6740 | n4837;
assign n5540 = ~n9777;
assign n3242 = ~(n1277 ^ n11627);
assign n3032 = n2449 | n12388;
assign n2511 = ~(n3223 ^ n1518);
assign n10109 = ~n13220;
assign n4588 = n5466 | n11025;
assign n5109 = n6118 | n5384;
assign n9660 = n13128 | n10858;
assign n11720 = ~(n3414 | n5708);
assign n9981 = n6602 & n9255;
assign n6233 = ~(n4579 | n4763);
assign n12825 = n5854 | n13172;
assign n11300 = ~n10770;
assign n5473 = ~(n7289 | n9285);
assign n9987 = n1208 | n7264;
assign n9717 = n5341 & n9108;
assign n3706 = n8696 | n12351;
assign n3401 = ~(n12090 ^ n5534);
assign n4435 = ~(n10469 ^ n4404);
assign n8870 = ~(n1753 ^ n1915);
assign n5480 = n11582 ^ n751;
assign n3609 = n10533 | n12919;
assign n10655 = n2506 & n5093;
assign n740 = ~n3511;
assign n11859 = n3208 | n8268;
assign n1972 = n7188 | n5797;
assign n4437 = ~(n1003 ^ n4733);
assign n2541 = ~n10343;
assign n6540 = n6733 | n8702;
assign n10012 = n2168 & n1445;
assign n12051 = n10604 | n1516;
assign n1209 = n10670 & n5172;
assign n7118 = ~(n13136 ^ n702);
assign n7979 = n8940 & n8233;
assign n10152 = n1188 | n8348;
assign n7294 = ~(n4052 ^ n6616);
assign n3639 = ~n9820;
assign n10727 = ~n10024;
assign n1730 = ~(n12946 | n2508);
assign n3464 = n2272 & n4704;
assign n2366 = ~(n6476 ^ n555);
assign n890 = n3456 & n5355;
assign n6641 = ~(n7094 ^ n1086);
assign n4755 = n9557 | n2958;
assign n10766 = ~(n948 ^ n9211);
assign n6683 = ~(n2697 ^ n12160);
assign n10631 = n10001 | n5209;
assign n11076 = ~(n9193 ^ n2797);
assign n700 = ~(n13188 | n1288);
assign n2169 = n11165 & n3201;
assign n3067 = n13151 & n2598;
assign n11872 = n80 | n542;
assign n7830 = n10170 & n12221;
assign n366 = ~(n141 ^ n607);
assign n7753 = n2702 & n5057;
assign n8057 = ~(n2774 | n67);
assign n629 = n6126 | n2627;
assign n11011 = ~(n9664 | n6047);
assign n3803 = ~(n1048 | n9106);
assign n10750 = n7510 & n3812;
assign n10983 = ~(n3267 ^ n33);
assign n1349 = ~n3682;
assign n1984 = n4385 | n7930;
assign n7570 = n7355 | n9259;
assign n11401 = ~(n9829 ^ n423);
assign n7078 = n973 | n2281;
assign n6436 = n11122 | n8268;
assign n2696 = n946 | n479;
assign n11414 = n1422 | n2059;
assign n214 = ~(n32 | n4020);
assign n12574 = n12211 & n3775;
assign n1957 = ~n744;
assign n11907 = ~(n12650 ^ n11996);
assign n3910 = n1638 | n12188;
assign n1495 = n10057 | n4947;
assign n2892 = ~(n8310 ^ n3081);
assign n5300 = ~(n11597 ^ n1483);
assign n3346 = ~(n5590 ^ n12935);
assign n1275 = ~(n8144 ^ n1666);
assign n12167 = n12203 | n3949;
assign n2995 = n5177 & n8098;
assign n7903 = ~n9620;
assign n8929 = ~(n4331 | n1151);
assign n5348 = ~n9241;
assign n2172 = ~(n12233 ^ n8105);
assign n9953 = n8580 & n6242;
assign n10835 = n11446 | n3949;
assign n7579 = n6728 & n2027;
assign n130 = n7433 & n9107;
assign n4123 = ~(n3113 ^ n1250);
assign n3445 = ~n9362;
assign n3680 = ~(n4388 ^ n11246);
assign n13079 = n8517 & n11187;
assign n1518 = ~(n9524 ^ n2947);
assign n2520 = n6865 | n5792;
assign n6591 = n6686 | n6786;
assign n13114 = ~(n6679 ^ n9573);
assign n3763 = ~(n3016 ^ n4501);
assign n11517 = n12916 | n657;
assign n3160 = n11979 | n9360;
assign n4861 = ~(n7924 ^ n7994);
assign n5324 = n958 & n11681;
assign n8036 = n10903 & n5215;
assign n10273 = n10276 & n12183;
assign n479 = n917;
assign n4536 = ~n8183;
assign n8656 = ~(n12947 | n9568);
assign n1070 = ~n9297;
assign n11144 = n6274;
assign n10418 = n11308 & n9321;
assign n6124 = ~(n1892 ^ n4297);
assign n8603 = ~(n989 ^ n11575);
assign n9886 = ~(n11844 | n9076);
assign n12942 = ~(n6686 ^ n2760);
assign n7867 = n8890 | n5955;
assign n10686 = n10802 & n2785;
assign n6772 = n11310 | n6827;
assign n3129 = n5945 & n2950;
assign n3977 = n7847 & n5170;
assign n2213 = ~n6532;
assign n8742 = ~(n4563 ^ n1228);
assign n11349 = ~(n4432 ^ n6119);
assign n12962 = ~(n9095 ^ n11103);
assign n10118 = ~(n7633 ^ n77);
assign n1203 = ~(n2495 ^ n9246);
assign n7940 = n6854 | n8754;
assign n152 = n12882 | n8268;
assign n1899 = n2912 & n672;
assign n5944 = n8499 | n1144;
assign n5477 = ~(n6337 ^ n10881);
assign n11451 = n10293 | n2038;
assign n2181 = n3622 & n7230;
assign n3664 = n2176 & n881;
assign n10186 = n1437 & n10200;
assign n11133 = n9145 & n6036;
assign n12891 = ~(n1227 | n4024);
assign n3403 = ~(n4821 ^ n4268);
assign n4237 = ~n11324;
assign n6841 = ~n8139;
assign n3495 = ~(n4735 ^ n2972);
assign n6285 = n5803 & n3193;
assign n2058 = n10117 & n10005;
assign n2043 = ~(n3135 ^ n4989);
assign n7991 = n3727 | n118;
assign n8745 = ~(n5776 ^ n9457);
assign n3419 = ~n9134;
assign n7018 = n10977 | n5797;
assign n9960 = n10861 & n5071;
assign n2818 = n13082 | n8534;
assign n4566 = ~n11774;
assign n5385 = n9917 | n2943;
assign n2243 = n436 | n9453;
assign n9671 = n9335 | n8524;
assign n3912 = ~(n1411 | n476);
assign n2784 = ~(n954 | n1996);
assign n5906 = ~(n630 | n12753);
assign n2124 = n7230 | n3622;
assign n8885 = n4143 | n9195;
assign n9043 = ~n2820;
assign n1783 = ~n12284;
assign n7140 = ~(n2094 | n738);
assign n11325 = n7315 & n238;
assign n4099 = n3401 | n9233;
assign n2690 = ~(n2676 ^ n6868);
assign n3488 = n8405 & n936;
assign n12453 = ~(n2365 ^ n9007);
assign n34 = n7842 | n176;
assign n2988 = n1327 | n9375;
assign n2880 = ~n2762;
assign n5283 = ~(n3382 | n10640);
assign n9012 = n5901 & n12119;
assign n8467 = n9382 & n10361;
assign n4985 = n5565 | n9195;
assign n10185 = ~(n13104 ^ n8566);
assign n9194 = ~(n2409 ^ n6358);
assign n5997 = n2158 & n11271;
assign n9750 = n7700 | n1570;
assign n12940 = ~n9981;
assign n2333 = n6942 & n13240;
assign n11432 = n6501 & n272;
assign n6742 = n7277 | n5378;
assign n5661 = n12709 | n431;
assign n2989 = n4652 & n9700;
assign n8709 = ~(n1230 ^ n9699);
assign n2140 = ~(n9585 | n3766);
assign n2247 = ~(n6850 ^ n8553);
assign n5866 = ~(n12591 ^ n10047);
assign n8588 = ~(n3423 ^ n2357);
assign n6642 = ~(n136 ^ n9744);
assign n339 = n7699 & n8703;
assign n11787 = n10077 | n4994;
assign n10928 = n6575 | n9504;
assign n4899 = n2091 & n3597;
assign n9261 = ~(n4752 ^ n10561);
assign n8904 = ~n12853;
assign n6425 = n5161 & n9119;
assign n13153 = ~(n11504 | n10262);
assign n640 = ~n405;
assign n5229 = ~n4315;
assign n6571 = n11149 | n8352;
assign n6522 = n10352 | n11107;
assign n2285 = n1047 & n963;
assign n9738 = n11829 & n6940;
assign n5434 = ~n7726;
assign n3051 = n45 | n8563;
assign n2958 = n12954;
assign n6722 = n4564 | n6370;
assign n1160 = n7044 & n12368;
assign n6983 = ~n9885;
assign n10380 = ~n465;
assign n11776 = ~(n9205 ^ n5425);
assign n12092 = ~n12715;
assign n5440 = n899 | n11107;
assign n665 = n8252 & n3120;
assign n11691 = ~(n6927 ^ n3107);
assign n5689 = ~(n4912 ^ n7773);
assign n8538 = n5961 & n4244;
assign n9795 = ~n12269;
assign n8838 = n8460 & n2291;
assign n10480 = n5351 | n12659;
assign n9489 = ~n8468;
assign n4418 = n9450 | n1570;
assign n3412 = ~n11248;
assign n11200 = n695 & n7483;
assign n9898 = n1246 & n10597;
assign n3501 = n12795 | n8702;
assign n7992 = ~(n9207 ^ n12207);
assign n2277 = n500 & n13241;
assign n6209 = n1972 ^ n10015;
assign n1262 = ~(n4805 ^ n909);
assign n4487 = ~n9904;
assign n12961 = ~(n10511 ^ n706);
assign n779 = ~(n8731 | n3175);
assign n7198 = ~(n6717 | n9812);
assign n10036 = n489 & n12206;
assign n3440 = ~(n3309 | n4513);
assign n6996 = n2292 & n2362;
assign n5085 = n7774 | n11355;
assign n4495 = ~n6168;
assign n5831 = ~(n4924 | n4919);
assign n7665 = n3978 | n8270;
assign n5611 = ~n7659;
assign n4518 = n8228 & n6085;
assign n1065 = n1152 | n1463;
assign n8814 = ~(n12608 ^ n7310);
assign n8986 = n5159 & n10496;
assign n8549 = ~(n1107 ^ n9541);
assign n12044 = n12741 | n13086;
assign n7701 = n12754 & n11714;
assign n5652 = ~(n7728 | n9804);
assign n189 = ~n103;
assign n3583 = n1017 | n8281;
assign n543 = n9348 & n4271;
assign n3894 = ~n7436;
assign n2709 = ~(n6987 ^ n6646);
assign n7440 = n2090 & n3834;
assign n7620 = ~n4748;
assign n4569 = ~(n3417 ^ n12432);
assign n4264 = ~(n7023 ^ n11497);
assign n9147 = n4358 & n6268;
assign n12633 = n9385 | n670;
assign n6960 = ~n6535;
assign n12132 = n5666 | n2133;
assign n8982 = n10208 | n8683;
assign n8296 = n3111 | n11169;
assign n3851 = n9411 | n7440;
assign n5592 = n8028 | n2746;
assign n8133 = n2183 | n12695;
assign n560 = ~n353;
assign n1681 = n136 | n5816;
assign n3305 = ~(n6203 ^ n763);
assign n11104 = n4948 | n11362;
assign n5691 = ~(n1034 ^ n12925);
assign n12382 = n2090 | n3834;
assign n12623 = ~n9620;
assign n7453 = n1508 | n5454;
assign n6111 = n115 | n479;
assign n3787 = ~(n6213 ^ n7144);
assign n2066 = n11519 | n5242;
assign n6947 = n700 | n6284;
assign n5622 = ~(n3188 | n4002);
assign n11573 = ~(n9500 | n1492);
assign n4018 = ~(n11715 | n5289);
assign n1961 = n5983 & n5370;
assign n6864 = n4714 & n3690;
assign n5792 = ~(n8357 | n8134);
assign n10202 = n7892 & n11599;
assign n5272 = ~(n6453 ^ n11647);
assign n7513 = ~(n3868 ^ n8564);
assign n4868 = ~(n11230 | n799);
assign n122 = n5423 | n8348;
assign n2059 = n11148;
assign n5101 = ~(n547 ^ n8676);
assign n8167 = n7299 | n4082;
assign n10407 = n6374 & n3933;
assign n1992 = ~(n6014 ^ n5754);
assign n6889 = ~n828;
assign n3106 = n10113 & n2252;
assign n2705 = n12215 & n10220;
assign n12035 = ~(n5027 ^ n9446);
assign n11327 = ~(n8550 ^ n1114);
assign n1013 = n8386 & n615;
assign n7400 = n1538 & n641;
assign n2518 = n13117 | n2387;
assign n8278 = n7461 & n8148;
assign n9596 = ~n13138;
assign n13037 = n13216 & n6502;
assign n7491 = n9978 & n4322;
assign n10393 = ~(n3845 ^ n1215);
assign n10799 = ~(n549 ^ n4441);
assign n2798 = n4744 & n10244;
assign n2304 = n13047 & n8394;
assign n2679 = n1319 & n3984;
assign n3642 = n4440 & n8846;
assign n6590 = ~n4470;
assign n1504 = n871 | n8514;
assign n7066 = ~(n11725 ^ n3052);
assign n11915 = n12617 | n8702;
assign n2965 = n6918 & n4061;
assign n8002 = ~n2310;
assign n3873 = ~(n9601 ^ n8934);
assign n7414 = n10402 | n3981;
assign n8952 = n4827 | n2240;
assign n5808 = n11990 ^ n8558;
assign n9197 = ~(n9084 ^ n12744);
assign n10010 = ~n11266;
assign n3771 = ~(n4867 ^ n10995);
assign n11730 = ~(n12022 | n10316);
assign n1976 = ~n1190;
assign n3416 = n618 & n9858;
assign n8946 = n9696 | n11011;
assign n4657 = ~n8332;
assign n8447 = n13137 | n5130;
assign n11125 = n11242 | n5797;
assign n4315 = n6320 & n127;
assign n8488 = n75 | n7530;
assign n10458 = n12921 & n9600;
assign n9243 = ~(n7126 | n2227);
assign n2903 = ~(n8461 ^ n6007);
assign n2055 = ~n10463;
assign n11612 = ~n817;
assign n12472 = n1194 | n2675;
assign n12258 = ~n295;
assign n320 = ~n8432;
assign n941 = ~(n2230 ^ n11726);
assign n4000 = ~(n8931 ^ n10416);
assign n10892 = ~n1313;
assign n11232 = ~n10442;
assign n12897 = n12023 | n2449;
assign n12237 = n7963 & n3334;
assign n13209 = n8443 & n132;
assign n10209 = ~(n1491 ^ n1109);
assign n3593 = ~(n257 ^ n4190);
assign n4469 = n910 & n178;
assign n3657 = n11212 | n206;
assign n4642 = ~n11666;
assign n251 = ~(n3249 ^ n10403);
assign n10257 = ~(n13018 | n355);
assign n4893 = n11514 | n11244;
assign n12460 = ~(n2076 ^ n8390);
assign n1442 = n6922 | n4724;
assign n6226 = n12997 | n5797;
assign n13145 = n9008 & n3118;
assign n4488 = ~n10821;
assign n7839 = ~n4033;
assign n4416 = ~(n8605 | n112);
assign n11722 = n5806 | n3981;
assign n203 = n6337 | n10881;
assign n2369 = ~(n11671 ^ n9062);
assign n1804 = ~(n1134 | n3283);
assign n7800 = ~(n11304 | n4463);
assign n4200 = ~(n9494 | n2996);
assign n1846 = n3530 | n5676;
assign n755 = ~n8820;
assign n2773 = ~n1756;
assign n9056 = ~(n4641 | n6817);
assign n4986 = ~(n5504 ^ n5732);
assign n1192 = n12027 & n11502;
assign n10287 = ~n4075;
assign n12613 = n1224 | n7781;
assign n5921 = ~n925;
assign n7626 = ~(n7806 | n11290);
assign n10357 = ~(n9293 ^ n6400);
assign n13048 = ~(n12293 ^ n2907);
assign n9517 = n12599 | n941;
assign n12566 = n6073 & n4544;
assign n31 = ~(n1789 ^ n2908);
assign n8536 = ~(n8205 ^ n11834);
assign n10486 = ~(n4328 | n12320);
assign n1205 = ~(n7156 ^ n4843);
assign n4300 = n3820 & n4308;
assign n7837 = ~n2771;
assign n4750 = n11612 | n7935;
assign n6827 = n5301 & n422;
assign n11258 = n11431 | n4435;
assign n2134 = n383 | n11899;
assign n1075 = n767 & n2498;
assign n3042 = ~(n1917 ^ n9777);
assign n12358 = n2722 & n2146;
assign n1277 = ~(n8799 ^ n1665);
assign n13126 = n11226 | n4640;
assign n11549 = n11450 & n4757;
assign n7993 = ~(n7876 ^ n3692);
assign n12378 = ~n5161;
assign n7312 = ~n12538;
assign n4516 = n10560 & n1636;
assign n9024 = ~(n6867 ^ n2454);
assign n2391 = n8527 & n2143;
assign n3458 = ~(n11159 ^ n3952);
assign n11883 = ~(n11702 | n11710);
assign n9761 = ~n834;
assign n12873 = n10876 & n3645;
assign n495 = n2701 | n10029;
assign n5275 = n6723 & n2327;
assign n4981 = n10047 & n12591;
assign n3168 = n13201 & n3815;
assign n2854 = n10814 | n11668;
assign n12277 = ~(n12765 ^ n11346);
assign n7373 = ~(n437 ^ n10028);
assign n952 = n6676 & n9869;
assign n10693 = ~(n11798 | n551);
assign n11013 = ~(n1531 ^ n2001);
assign n1582 = n9490 | n9618;
assign n10390 = n12095 & n6464;
assign n10016 = ~n10642;
assign n5683 = ~n6085;
assign n1216 = ~n4957;
assign n5034 = n9762 & n3038;
assign n12590 = n8414 | n4124;
assign n11854 = n7715 & n9669;
assign n5382 = ~n7419;
assign n4338 = ~(n12559 ^ n6026);
assign n8161 = ~n1356;
assign n10784 = ~(n7025 | n6994);
assign n13012 = ~n5715;
assign n4199 = n715 | n4936;
assign n8442 = ~(n6754 ^ n4009);
assign n10789 = ~(n122 ^ n10303);
assign n4464 = ~n4330;
assign n488 = ~n6085;
assign n7054 = n11600 & n2610;
assign n9902 = ~(n12541 ^ n3680);
assign n6032 = ~(n11139 ^ n10393);
assign n10452 = n8461 & n6388;
assign n2847 = ~(n8567 ^ n12176);
assign n8911 = n6967 | n11871;
assign n5467 = ~n3627;
assign n12872 = ~(n2888 ^ n11066);
assign n11788 = ~(n10807 ^ n12656);
assign n11447 = ~(n6669 ^ n11872);
assign n9896 = ~(n11270 ^ n6899);
assign n72 = n7949 & n3215;
assign n7526 = ~n7728;
assign n4163 = ~(n9306 ^ n6430);
assign n12653 = ~(n6930 | n377);
assign n6342 = ~(n1753 | n1915);
assign n749 = n8500 & n3860;
assign n9192 = n7681 & n9066;
assign n9218 = ~(n1173 ^ n8347);
assign n10058 = ~(n4308 ^ n3820);
assign n3721 = n2048 | n121;
assign n8067 = ~(n5096 ^ n9536);
assign n9938 = n10730 | n5076;
assign n4241 = n392 | n6041;
assign n9729 = n8131 | n4640;
assign n975 = ~(n13069 ^ n1130);
assign n9498 = ~(n2102 | n4838);
assign n11052 = n4588 & n1914;
assign n8035 = ~(n4316 ^ n3573);
assign n11182 = ~(n2949 ^ n10789);
assign n3811 = ~(n3664 | n6408);
assign n8887 = n813 | n10871;
assign n10139 = ~(n8998 ^ n4076);
assign n10313 = n10439 | n1026;
assign n2065 = ~(n11730 | n6443);
assign n5565 = ~n2252;
assign n10268 = n7529 & n2252;
assign n3543 = n6630 | n4230;
assign n6885 = ~(n10925 | n4256);
assign n13213 = n563 & n9677;
assign n1828 = n9421 | n8490;
assign n7989 = ~(n2087 | n10557);
assign n4751 = n5934 & n4461;
assign n1142 = ~(n7231 ^ n12519);
assign n3153 = ~(n5139 ^ n5518);
assign n5028 = ~(n8626 | n2841);
assign n2072 = n912 ^ n3831;
assign n11724 = ~(n1172 ^ n6681);
assign n1077 = n12069 | n9761;
assign n10925 = ~(n12539 ^ n10702);
assign n9711 = ~n9528;
assign n5869 = n3586 | n1771;
assign n11647 = n1012 | n956;
assign n923 = ~(n2013 ^ n205);
assign n11903 = ~(n12134 ^ n7574);
assign n10991 = ~n772;
assign n9921 = ~n7572;
assign n7782 = ~(n11499 ^ n6784);
assign n2187 = ~(n8717 | n3869);
assign n6411 = ~(n7483 ^ n4332);
assign n3367 = n2226 | n9622;
assign n2273 = n3311 & n411;
assign n2130 = ~n12567;
assign n1238 = ~n5768;
assign n5049 = ~(n9842 ^ n12803);
assign n8527 = ~(n11015 ^ n2121);
assign n1698 = n2482 & n2758;
assign n2671 = ~n3130;
assign n7654 = ~(n901 ^ n4775);
assign n9481 = n2777 & n8860;
assign n726 = n12475 ^ n5488;
assign n6866 = n10733 | n10331;
assign n7085 = n11553 ^ n11641;
assign n1215 = ~n6445;
assign n3837 = n1579 & n11307;
assign n5851 = n3784 | n9075;
assign n11045 = ~n600;
assign n4953 = ~(n10660 ^ n7351);
assign n9094 = n7620 | n1985;
assign n1968 = n5733 | n5242;
assign n8589 = ~(n11541 ^ n3742);
assign n1114 = ~(n13119 ^ n5499);
assign n8548 = n4610 | n5169;
assign n6361 = ~(n12857 ^ n7804);
assign n8335 = ~n5969;
assign n6507 = n490 & n6389;
assign n6382 = n11284 | n12273;
assign n11510 = ~(n7359 ^ n3199);
assign n4800 = ~(n5120 ^ n8821);
assign n3790 = ~(n10897 ^ n4996);
assign n13125 = n3284 & n6813;
assign n3021 = ~(n385 ^ n3523);
assign n10768 = n4001 | n12177;
assign n9929 = n4818 & n1602;
assign n12992 = n10638 | n8983;
assign n10349 = ~(n10578 | n5282);
assign n2163 = ~n11179;
assign n8179 = n870 & n11655;
assign n3868 = ~(n7382 ^ n10461);
assign n359 = ~(n8967 ^ n12163);
assign n1259 = n3090 | n990;
assign n2351 = n1715 & n8313;
assign n6165 = ~(n4645 ^ n2447);
assign n5629 = ~(n8158 ^ n12360);
assign n869 = n5902 | n11606;
assign n9592 = ~n7085;
assign n9233 = n10289 & n4755;
assign n8690 = ~(n13121 ^ n11348);
assign n987 = ~n12065;
assign n11229 = n11751 | n1820;
assign n1499 = n10962 | n10473;
assign n513 = ~n229;
assign n4727 = n1101 | n10871;
assign n8612 = ~(n690 ^ n6893);
assign n4952 = ~(n5071 | n10861);
assign n2718 = ~n9620;
assign n7971 = n9515 | n2569;
assign n10654 = ~n3095;
assign n3157 = ~n103;
assign n5673 = ~n7153;
assign n4824 = n5965 ^ n485;
assign n570 = n7925 | n8563;
assign n1395 = n10479 & n11434;
assign n7815 = ~(n9989 ^ n12692);
assign n2450 = ~(n9235 | n9506);
assign n4713 = ~(n9150 ^ n2397);
assign n9482 = n11845 | n4658;
assign n13193 = ~(n11361 ^ n13016);
assign n12765 = n10085 | n1570;
assign n10595 = n8717 & n3869;
assign n2893 = ~n8230;
assign n6789 = n6066 & n3706;
assign n1385 = ~(n10446 ^ n10939);
assign n3145 = n7443 & n12442;
assign n9028 = ~(n10046 ^ n5259);
assign n2079 = n7872 | n8744;
assign n4737 = n3348 | n11748;
assign n1995 = ~(n2440 | n13163);
assign n3842 = n3733 | n11426;
assign n8005 = ~n2590;
assign n7166 = ~(n9861 ^ n1207);
assign n5846 = n1168 | n8348;
assign n7276 = n1757 & n4330;
assign n11211 = ~(n2261 ^ n7061);
assign n7901 = n1633 | n5524;
assign n10911 = ~(n12754 ^ n7451);
assign n10454 = ~(n705 | n9208);
assign n11072 = ~(n2730 ^ n11440);
assign n12471 = ~n767;
assign n9679 = ~n5320;
assign n10411 = ~n1982;
assign n6164 = ~n8917;
assign n1346 = ~n6836;
assign n2795 = n6054 | n5290;
assign n12185 = n8670 | n2707;
assign n388 = ~(n6195 ^ n12886);
assign n11270 = ~n691;
assign n11569 = n8642 & n8488;
assign n7664 = ~(n7671 ^ n8078);
assign n9916 = ~(n8718 | n11531);
assign n10846 = ~(n7593 ^ n10701);
assign n8543 = n104 & n6911;
assign n11833 = ~(n7500 | n3681);
assign n9150 = n4166 | n6404;
assign n9225 = n12361 & n10317;
assign n2923 = ~(n12217 ^ n7164);
assign n6850 = n4966 | n9714;
assign n10987 = ~(n4750 ^ n11475);
assign n9267 = ~(n3309 ^ n11534);
assign n4440 = n11665 & n8860;
assign n4669 = n8736 & n7081;
assign n8852 = ~n5214;
assign n2293 = ~(n6722 ^ n7416);
assign n8909 = n9634 | n12029;
assign n10816 = ~(n10331 ^ n13226);
assign n7068 = ~n9528;
assign n2089 = n5268 & n7012;
assign n9275 = ~(n7715 | n2458);
assign n1710 = n5442 & n181;
assign n10785 = ~(n10804 ^ n1573);
assign n3288 = n11320 | n10871;
assign n1920 = ~n6064;
assign n2781 = n12565 | n5067;
assign n13029 = ~(n6780 ^ n2111);
assign n11602 = ~(n2058 | n6907);
assign n4059 = ~(n2731 ^ n5880);
assign n3191 = n2449 | n1570;
assign n4461 = n4348 | n7813;
assign n8009 = n3025 | n4510;
assign n4733 = n5129 & n9180;
assign n9206 = ~(n7118 ^ n12480);
assign n6861 = n10544 ^ n1064;
assign n12667 = ~n6950;
assign n4832 = ~(n2821 ^ n5343);
assign n7980 = ~n6277;
assign n1877 = ~(n4205 | n1351);
assign n6871 = n12522 | n5775;
assign n3981 = n789;
assign n2824 = ~n5833;
assign n9451 = n2384 | n3396;
assign n11085 = n7797 & n5996;
assign n3818 = n6086 | n12188;
assign n800 = ~(n8587 ^ n4707);
assign n2768 = ~n4335;
assign n4739 = n5784 ^ n7722;
assign n8137 = ~(n2361 ^ n11897);
assign n4890 = ~n3832;
assign n12949 = n2583 & n10673;
assign n1762 = n2472 & n11593;
assign n7960 = n11665 & n9570;
assign n7932 = ~(n3739 ^ n325);
assign n8778 = ~n3988;
assign n9736 = ~n11474;
assign n10469 = n4855 | n2958;
assign n11355 = ~(n52 ^ n11923);
assign n2014 = ~(n8411 ^ n807);
assign n6981 = n7177 | n10551;
assign n4587 = n6884 & n6424;
assign n6737 = ~(n10047 | n12591);
assign n4724 = n3858;
assign n2678 = ~n11734;
assign n8239 = n2576 | n8262;
assign n12833 = n13190 | n6265;
assign n1480 = ~n11734;
assign n10711 = ~n3715;
assign n10771 = n2896 | n10311;
assign n9361 = n7878 | n10552;
assign n10650 = n4649 | n2059;
assign n12716 = n11965 | n10764;
assign n10624 = n5645 | n6732;
assign n11867 = n12648 | n8561;
assign n12231 = n417 & n7109;
assign n13099 = n881 | n2176;
assign n11083 = ~(n11572 ^ n1584);
assign n4322 = n12020 | n3210;
assign n10658 = n12010 & n11451;
assign n12315 = ~n2374;
assign n12187 = ~(n3862 ^ n571);
assign n6434 = ~(n824 ^ n1318);
assign n13144 = ~(n5874 ^ n10468);
assign n4752 = ~(n3615 | n5507);
assign n4721 = ~(n9645 ^ n10056);
assign n4778 = ~n382;
assign n7924 = ~(n4217 ^ n3029);
assign n10561 = n1360 | n9511;
assign n11340 = ~n11199;
assign n2396 = n9593 | n8806;
assign n1554 = ~n937;
assign n5222 = ~n299;
assign n11105 = n9341 | n2594;
assign n6572 = ~(n3802 ^ n2459);
assign n12431 = n9339 | n9159;
assign n710 = ~(n4576 ^ n9773);
assign n8323 = ~(n8426 ^ n11754);
assign n8515 = ~(n9534 ^ n3268);
assign n10459 = ~n9901;
assign n8107 = n13205 | n4310;
assign n3967 = n7470 & n3020;
assign n4290 = ~n9531;
assign n2548 = ~(n6067 ^ n1076);
assign n8756 = ~(n3305 | n5662);
assign n845 = ~n7729;
assign n723 = n3429 | n4030;
assign n7785 = n3936 & n4810;
assign n2382 = ~(n9535 ^ n2852);
assign n5796 = ~(n9107 ^ n4520);
assign n11408 = n10593 | n3063;
assign n12561 = ~(n5309 | n1000);
assign n1228 = ~(n2128 ^ n8403);
assign n2832 = ~n12422;
assign n6039 = n9252 | n3464;
assign n8027 = ~(n10913 ^ n3746);
assign n1789 = ~n3253;
assign n8314 = n53 | n6769;
assign n2825 = ~n5189;
assign n11919 = n6043 | n327;
assign n9951 = ~(n10514 ^ n7293);
assign n11413 = ~(n1991 ^ n8603);
assign n7362 = ~n13128;
assign n12543 = n12992 & n9409;
assign n9539 = n4665 | n1985;
assign n5695 = n1511 | n11668;
assign n10879 = ~n5031;
assign n10092 = n7258 | n12234;
assign n5617 = ~(n9874 ^ n6397);
assign n5491 = n10354 | n12763;
assign n8584 = ~(n487 ^ n9239);
assign n6218 = n11318 | n8880;
assign n9752 = n3583 & n13010;
assign n2348 = n300 | n10619;
assign n4744 = ~n1595;
assign n5036 = n10346 & n2534;
assign n11362 = n11415 & n7564;
assign n5966 = n7984 | n11470;
assign n2067 = ~n7137;
assign n4802 = ~(n11142 ^ n11762);
assign n7419 = n10188 | n4947;
assign n7887 = n5667 | n11144;
assign n5676 = n3022 & n12807;
assign n12344 = n12224 | n4979;
assign n12011 = ~(n12081 ^ n9936);
assign n11633 = n1265 | n2552;
assign n2673 = ~n1552;
assign n9877 = n5079 | n1144;
assign n9661 = n898 & n4154;
assign n11649 = ~(n244 | n2436);
assign n9313 = n4796 | n4947;
assign n7751 = n2118 | n12273;
assign n12735 = ~(n4508 | n7686);
assign n10339 = n11339 & n1080;
assign n9198 = ~(n12061 ^ n753);
assign n12375 = n8934 | n4423;
assign n1351 = n3898 | n9223;
assign n10690 = ~(n3254 | n3979);
assign n1292 = n581 & n8957;
assign n11742 = n12242 | n5087;
assign n5285 = ~(n3138 | n11316);
assign n3643 = n2451 & n2799;
assign n11771 = ~n13219;
assign n12928 = ~(n10197 ^ n10615);
assign n9520 = n278 | n11968;
assign n11987 = n12748 | n10871;
assign n6287 = ~(n11229 ^ n7758);
assign n13221 = n10761 | n13242;
assign n9269 = ~(n9683 | n5849);
assign n2034 = n97 | n4373;
assign n12831 = ~(n11653 ^ n13042);
assign n5379 = n12129 & n10960;
assign n6494 = ~(n3518 | n1069);
assign n3860 = n11986 & n10376;
assign n4567 = ~(n4568 | n3353);
assign n4837 = ~(n6861 ^ n1802);
assign n6269 = n2590 & n8290;
assign n9827 = ~n6317;
assign n11898 = n11994 & n331;
assign n1532 = ~(n12584 ^ n3045);
assign n4409 = ~(n7788 ^ n8007);
assign n6426 = n11819 & n8775;
assign n6775 = n6710 | n5782;
assign n11402 = n5568 & n4748;
assign n10426 = n4235 | n3576;
assign n5177 = ~n12557;
assign n10891 = n9011 | n3559;
assign n841 = ~(n12796 ^ n8308);
assign n8523 = n3944 & n3541;
assign n10402 = ~n1636;
assign n4772 = ~(n7849 ^ n5543);
assign n7558 = ~(n8830 ^ n10181);
assign n171 = ~(n7806 ^ n11377);
assign n9317 = ~(n5744 ^ n7715);
assign n12172 = n13006 ^ n10268;
assign n6569 = ~(n250 | n2492);
assign n7233 = ~(n9543 | n2489);
assign n5544 = ~(n4559 ^ n5675);
assign n6817 = ~(n4573 | n10838);
assign n714 = n8324 | n2675;
assign n4471 = n2405 | n8614;
assign n4459 = ~(n5197 ^ n6600);
assign n5030 = ~(n8657 ^ n9127);
assign n10166 = ~(n7560 | n6600);
assign n6239 = n1607 & n9780;
assign n12345 = ~(n4768 ^ n3943);
assign n11660 = n6183 | n3977;
assign n8804 = ~(n3501 ^ n7607);
assign n9214 = ~(n536 ^ n4581);
assign n6438 = ~n1165;
assign n5381 = n6314 | n2354;
assign n1125 = n10558 | n4724;
assign n9117 = n4211 ^ n10485;
assign n5151 = n1101 | n2387;
assign n11449 = ~n6392;
assign n10652 = n1460 & n5506;
assign n12328 = n9280;
assign n2368 = ~(n11035 ^ n1439);
assign n9920 = n100 & n9725;
assign n3417 = n10128 | n11107;
assign n11407 = n935 | n4230;
assign n6314 = ~n7527;
assign n8995 = ~n4788;
assign n11707 = ~n2409;
assign n9505 = ~(n12769 ^ n2909);
assign n8474 = n8912 | n2622;
assign n10623 = n12915 & n4487;
assign n4231 = n1024 & n4294;
assign n6854 = ~n12482;
assign n5787 = ~n7240;
assign n12745 = ~(n6816 ^ n7332);
assign n10669 = ~(n8317 ^ n12212);
assign n10861 = ~(n6353 ^ n7431);
assign n4351 = ~(n2830 ^ n10833);
assign n10086 = ~(n7416 | n6722);
assign n2472 = ~n3390;
assign n1098 = n9489 | n2059;
assign n6725 = n2662 | n6863;
assign n8582 = ~(n696 ^ n9000);
assign n9999 = ~(n10024 ^ n1967);
assign n6812 = ~(n7345 ^ n8895);
assign n3353 = n9460 & n12452;
assign n1132 = n715 | n11668;
assign n10286 = ~n9620;
assign n3949 = n6274;
assign n11467 = ~(n9843 ^ n6528);
assign n7347 = ~(n6720 ^ n2584);
assign n4507 = ~(n4538 ^ n8667);
assign n11473 = n8350 & n6000;
assign n660 = ~(n4630 | n5312);
assign n428 = ~n10599;
assign n6169 = ~(n9926 ^ n5175);
assign n6949 = n7476 & n2301;
assign n2811 = n9478 | n1144;
assign n1714 = ~(n9975 ^ n7482);
assign n4693 = ~(n3885 | n6499);
assign n10468 = ~(n9122 ^ n7674);
assign n12416 = ~n2252;
assign n4069 = ~(n12598 ^ n4437);
assign n11711 = ~(n4081 | n9186);
assign n5360 = ~n12381;
assign n11579 = ~(n4065 ^ n3226);
assign n6587 = ~n10805;
assign n5830 = n13202 | n7016;
assign n11263 = n6133 | n4373;
assign n10883 = ~n5920;
assign n9191 = n11121 | n6899;
assign n8771 = ~(n4992 | n2399);
assign n322 = n2546 ^ n7477;
assign n13104 = ~(n2700 ^ n3575);
assign n7497 = n6670 & n7346;
assign n2656 = ~(n1954 ^ n1488);
assign n9107 = n5008 | n4110;
assign n4871 = n9383 | n5242;
assign n4213 = n6014 & n6359;
assign n5312 = ~n376;
assign n3441 = n9711 | n8030;
assign n2322 = n7503 | n11184;
assign n11332 = ~(n8070 ^ n8735);
assign n9873 = n248 & n8769;
assign n9962 = ~n5729;
assign n1809 = n12229 & n4941;
assign n10836 = ~(n8130 ^ n3190);
assign n330 = ~(n8866 | n8620);
assign n4676 = ~(n25 ^ n5901);
assign n6201 = ~(n4922 ^ n365);
assign n12903 = ~(n12558 ^ n12426);
assign n9940 = n8104 | n7528;
assign n9320 = n4519 | n7080;
assign n8340 = n11504 & n10262;
assign n1703 = n8594 & n12804;
assign n7770 = n1951 & n6526;
assign n4691 = n1630 & n5807;
assign n8324 = ~n9300;
assign n12749 = ~(n12301 ^ n2180);
assign n10372 = ~(n7676 | n1209);
assign n7232 = n175 | n9369;
assign n2315 = n10712 & n1864;
assign n11832 = ~(n9855 | n7063);
assign n10382 = ~(n1841 ^ n10938);
assign n4595 = n4967 | n8563;
assign n4366 = ~n8233;
assign n2559 = n7170 | n2631;
assign n8420 = n10225 ^ n10322;
assign n4238 = n7783 | n12388;
assign n9350 = ~n1826;
assign n2480 = n9275 | n5744;
assign n2581 = ~n10805;
assign n3307 = n4063 | n1218;
assign n10680 = n1563 ^ n2951;
assign n8525 = n423 | n9179;
assign n2691 = ~n10190;
assign n6358 = ~n12026;
assign n10400 = ~n9846;
assign n3804 = ~n1992;
assign n8761 = n3726 | n7723;
assign n11253 = n3911 | n9075;
assign n1785 = n7658 | n8512;
assign n11430 = n9648 | n8677;
assign n3414 = n10258 & n7823;
assign n12782 = ~(n11773 | n10116);
assign n11257 = ~(n3954 ^ n1792);
assign n8431 = n9554 & n4252;
assign n2952 = n10624 | n11708;
assign n3192 = n3877 | n8874;
assign n8740 = n12316 | n1422;
assign n3534 = ~n1636;
assign n347 = n8681 | n7723;
assign n12002 = ~(n7813 ^ n5742);
assign n1555 = ~(n4755 ^ n10289);
assign n10831 = ~(n2512 ^ n131);
assign n8856 = n11068 & n9308;
assign n3105 = ~(n8380 ^ n7596);
assign n8652 = ~(n11295 ^ n1982);
assign n11826 = ~(n10983 ^ n12154);
assign n11648 = n5148 | n4230;
assign n9903 = ~(n10516 ^ n5686);
assign n8262 = n9169 & n1796;
assign n8517 = ~(n5902 ^ n6092);
assign n3975 = n10650 | n921;
assign n920 = n12254 | n1043;
assign n12129 = n6828 | n11796;
assign n12244 = n12150 & n4145;
assign n1965 = ~n4557;
assign n4346 = n1073 & n6983;
assign n6560 = ~(n12470 | n7656);
assign n180 = ~(n5329 ^ n5701);
assign n12850 = n3804 & n12941;
assign n11490 = n1202 ^ n10808;
assign n2451 = ~(n4719 ^ n11412);
assign n7938 = n10977 | n8348;
assign n5391 = ~(n11907 ^ n12327);
assign n11320 = ~n4330;
assign n21 = n2255 | n9314;
assign n7603 = ~(n8331 ^ n1046);
assign n1904 = n755 | n3598;
assign n6900 = n12630 | n1240;
assign n8906 = n10423 | n264;
assign n10724 = n10854 | n837;
assign n12632 = n6633 ^ n11607;
assign n8361 = n6630 | n4373;
assign n5043 = ~(n6212 | n11219);
assign n314 = ~(n12688 | n4270);
assign n2505 = ~(n12840 ^ n4611);
assign n7973 = n305 | n5724;
assign n37 = n7358 | n1571;
assign n3254 = ~(n2284 | n8770);
assign n805 = ~(n1716 | n11438);
assign n10231 = n11910 | n2449;
assign n8868 = ~n13058;
assign n66 = n2595 ^ n8760;
assign n58 = ~(n8766 ^ n6874);
assign n11868 = ~n10451;
assign n10133 = ~(n2932 | n11182);
assign n12996 = ~(n2417 ^ n4319);
assign n12108 = ~(n2522 | n9998);
assign n8954 = n6099 | n1043;
assign n9355 = n11121 | n5802;
assign n11731 = ~(n5851 ^ n7413);
assign n1154 = n8307 & n4940;
assign n5510 = n8447 & n12292;
assign n12790 = n3676 | n3640;
assign n11773 = n10266 | n9745;
assign n12537 = ~n4964;
assign n3572 = ~n1982;
assign n5499 = n6486 | n12501;
assign n13002 = ~(n11190 ^ n10740);
assign n11863 = ~(n740 ^ n11738);
assign n2693 = ~(n12452 ^ n9115);
assign n7593 = ~(n9124 ^ n7229);
assign n10868 = ~(n2710 ^ n541);
assign n6875 = ~n9591;
assign n8168 = n8876 | n12487;
assign n8701 = ~(n2280 ^ n2185);
assign n4140 = ~(n7999 ^ n8171);
assign n690 = n10611 & n11307;
assign n2312 = ~(n6172 ^ n5756);
assign n11259 = n1062 & n12310;
assign n11639 = n6329 & n4883;
assign n3844 = ~(n8235 ^ n3100);
assign n11160 = ~(n5123 ^ n2029);
assign n756 = ~(n4759 ^ n5116);
assign n5481 = ~(n2651 ^ n10933);
assign n312 = ~n12112;
assign n12367 = n8838 ^ n3494;
assign n13161 = ~(n7979 ^ n3392);
assign n2978 = n2874 & n12815;
assign n3126 = ~n12965;
assign n3014 = ~(n13014 ^ n12751);
assign n11203 = n10143 | n4373;
assign n8432 = n9171 | n6257;
assign n10574 = ~n394;
assign n12376 = ~(n7485 | n4889);
assign n294 = n5157 | n12049;
assign n5052 = ~(n6065 ^ n1120);
assign n7010 = n9497 & n6330;
assign n6397 = ~(n12879 ^ n2494);
assign n8446 = n2022 | n1193;
assign n8114 = ~(n10915 ^ n10226);
assign n9419 = ~(n3088 ^ n7121);
assign n8260 = n12738 & n3543;
assign n10529 = n7953 | n11051;
assign n9413 = n3372 & n5544;
assign n1713 = n12465 | n11668;
assign n6878 = ~n9293;
assign n9607 = ~n5647;
assign n76 = n11104 & n6157;
assign n8614 = n3326 & n387;
assign n2756 = ~(n9522 ^ n10635);
assign n8552 = n9930 & n3980;
assign n11371 = ~(n686 ^ n2885);
assign n3599 = n2067 | n8096;
assign n4558 = n8977 | n10179;
assign n840 = n1778 | n9572;
assign n4690 = ~(n12025 ^ n8314);
assign n5949 = ~n6392;
assign n662 = n11225 | n2133;
assign n6931 = ~(n3101 ^ n2290);
assign n12096 = ~(n6753 ^ n4812);
assign n6455 = n1333 & n8842;
assign n5882 = ~(n7379 ^ n9165);
assign n11690 = n5498 | n8800;
assign n12984 = n11404 | n5797;
assign n2859 = ~(n10221 ^ n5812);
assign n6656 = ~(n9374 | n3389);
assign n6820 = ~(n1242 ^ n12173);
assign n9956 = ~(n4459 ^ n1662);
assign n6030 = ~(n8813 ^ n2470);
assign n10740 = n3006 & n10451;
assign n10641 = ~n2737;
assign n3570 = ~n11285;
assign n9875 = ~(n11334 ^ n9359);
assign n5550 = ~n11665;
assign n6067 = n795 | n10135;
assign n2316 = ~(n10150 ^ n12054);
assign n6564 = ~(n9526 | n10146);
assign n7682 = n11345 & n5250;
assign n3277 = ~(n7776 ^ n518);
assign n12878 = n10991 | n8268;
assign n10220 = n12295 | n3981;
assign n1665 = n11370 | n4724;
assign n13177 = n398 | n10813;
assign n3460 = ~n9570;
assign n11497 = n10137 | n2133;
assign n7332 = ~(n1419 ^ n30);
assign n391 = ~(n2072 | n8481);
assign n8044 = ~n1762;
assign n858 = ~(n6975 ^ n7871);
assign n10159 = ~(n4033 ^ n3552);
assign n496 = n9328 & n5948;
assign n9185 = ~(n10844 ^ n5042);
assign n2358 = n12648 | n9962;
assign n3408 = n3259 | n6732;
assign n1358 = ~n976;
assign n6636 = n10039 & n11110;
assign n11763 = ~(n1299 ^ n5397);
assign n7988 = n4085 & n10348;
assign n11953 = ~(n6821 ^ n1369);
assign n5774 = n69 | n12273;
assign n7462 = ~(n2466 ^ n11068);
assign n12570 = ~(n5419 ^ n10069);
assign n9088 = n12630 & n1240;
assign n3600 = n11818 & n10022;
assign n12207 = ~(n4284 ^ n9166);
assign n1061 = ~(n7193 ^ n9933);
assign n3776 = ~(n242 | n6941);
assign n11783 = ~n10025;
assign n2357 = n9129 | n1026;
assign n12567 = n12370 & n12824;
assign n13163 = ~(n3907 ^ n7513);
assign n4534 = n7114 & n4192;
assign n12146 = ~(n9049 ^ n1577);
assign n8208 = n7997 | n4959;
assign n11803 = n3836 | n1103;
assign n10328 = n5372 & n4481;
assign n1848 = ~(n7952 | n9571);
assign n13206 = ~(n8389 | n7192);
assign n11692 = n1571 | n8490;
assign n7435 = ~(n6148 ^ n6458);
assign n11642 = n10499 | n11843;
assign n3368 = ~(n10477 ^ n10484);
assign n6396 = ~(n9928 ^ n12314);
assign n8094 = n7765 & n10906;
assign n10242 = ~(n7156 | n1932);
assign n11281 = n1489 & n10806;
assign n2334 = n7544 & n198;
assign n7053 = ~(n3543 ^ n9367);
assign n11988 = n9216 & n9475;
assign n4967 = ~n6085;
assign n11956 = n3249 | n3161;
assign n12017 = n7475 & n8982;
assign n8788 = n6367 | n10319;
assign n1108 = ~(n7885 | n1187);
assign n8947 = ~(n8567 | n6718);
assign n8691 = ~(n7136 ^ n10698);
assign n12947 = ~(n7375 ^ n12618);
assign n6743 = ~n22;
assign n6990 = ~n5475;
assign n13160 = ~(n5316 ^ n8320);
assign n10527 = ~n10122;
assign n12153 = ~n11411;
assign n10589 = n7669 & n9101;
assign n1119 = ~(n8299 ^ n11752);
assign n1052 = ~n6826;
assign n6504 = ~n498;
assign n7418 = n8615 | n8268;
assign n12151 = ~(n1977 ^ n849);
assign n9339 = ~n11891;
assign n4860 = ~(n3148 ^ n4902);
assign n4722 = ~n3677;
assign n2071 = n5811 & n8202;
assign n913 = ~n6561;
assign n6566 = n11868 | n5076;
assign n7928 = ~(n4480 ^ n10598);
assign n3442 = n567 | n11833;
assign n437 = ~(n720 ^ n5600);
assign n12217 = ~(n1456 ^ n9333);
assign n3214 = n1367 | n5971;
assign n13039 = ~n3769;
assign n8493 = n8034 & n9496;
assign n2308 = n2607 & n6640;
assign n8016 = n9418 & n1214;
assign n4922 = ~(n3872 | n9301);
assign n12876 = n4441 & n2600;
assign n4033 = n8046 & n1410;
assign n12967 = ~n4470;
assign n801 = ~(n10965 ^ n2826);
assign n5657 = ~(n6494 ^ n4438);
assign n5587 = ~(n2774 ^ n4415);
assign n5051 = ~(n11039 ^ n11873);
assign n1105 = ~n587;
assign n792 = n4138 & n239;
assign n3431 = ~(n6206 ^ n2170);
assign n11871 = ~n761;
assign n8553 = ~(n4271 ^ n9348);
assign n12221 = ~n8156;
assign n8042 = n2296 | n7254;
assign n5209 = n655 & n2914;
assign n8075 = ~(n4439 | n2956);
assign n12388 = n7424;
assign n1684 = n5039 | n7821;
assign n12516 = n1651 | n6265;
assign n9068 = ~n3709;
assign n12498 = n12013 & n1632;
assign n908 = n10293 ^ n5480;
assign n10222 = ~(n12715 | n11027);
assign n3100 = ~(n12533 ^ n3694);
assign n4962 = n2692 | n3981;
assign n4277 = n734 | n493;
assign n7092 = ~(n1974 ^ n1595);
assign n12874 = n5795 | n5510;
assign n2352 = ~n10657;
assign n1196 = ~(n4651 ^ n12118);
assign n8710 = ~n10343;
assign n8892 = ~n10479;
assign n6753 = n10018 | n3981;
assign n8120 = n9350 | n10627;
assign n3957 = n3225 | n11668;
assign n12301 = ~(n9516 ^ n11789);
assign n8746 = ~(n13205 ^ n4310);
assign n11313 = n3696 | n447;
assign n9635 = ~n1603;
assign n9276 = ~n9685;
assign n7289 = n1416 | n10696;
assign n8360 = ~n6826;
assign n10379 = ~(n6412 ^ n12763);
assign n6671 = n5749 | n8534;
assign n8574 = n440 | n5431;
assign n12160 = ~(n7123 ^ n1119);
assign n11079 = n5508 & n861;
assign n7804 = ~(n8276 ^ n2905);
assign n7489 = ~(n11873 | n4529);
assign n7947 = n12713 | n7082;
assign n12305 = ~(n10077 ^ n9229);
assign n4583 = n2353 & n5542;
assign n12101 = n10575 ^ n5170;
assign n3462 = ~(n10152 | n5368);
assign n1612 = ~(n590 ^ n12977);
assign n6773 = ~(n7645 ^ n1200);
assign n11132 = ~n1273;
assign n8212 = ~n7051;
assign n11392 = n5271 | n8490;
assign n9881 = n5634 | n5242;
assign n10289 = n1705 & n2788;
assign n9457 = ~(n924 ^ n2938);
assign n4796 = ~n13058;
assign n12780 = n5581 | n5173;
assign n6324 = ~(n11187 ^ n6474);
assign n10775 = ~(n6809 ^ n11000);
assign n8393 = n4022 | n177;
assign n12703 = ~(n733 ^ n2200);
assign n3792 = n10650 & n921;
assign n1535 = ~(n11472 ^ n11949);
assign n2918 = n3318 & n5714;
assign n1564 = n11411 & n6168;
assign n2109 = ~n10142;
assign n7019 = n1185 | n1669;
assign n11279 = n12086 & n11988;
assign n11896 = ~(n1205 ^ n12146);
assign n4937 = n9080 | n9159;
assign n827 = ~(n9726 ^ n8962);
assign n9927 = n13051 | n2544;
assign n6973 = n7386 & n5745;
assign n2278 = ~n8940;
assign n5918 = ~(n11961 ^ n12571);
assign n13105 = n2713 & n7325;
assign n2332 = ~n3076;
assign n6994 = ~(n10306 ^ n8678);
assign n11168 = n13082 | n7221;
assign n4834 = ~(n1410 ^ n8046);
assign n4627 = n5329 | n4503;
assign n10260 = n756 | n5221;
assign n11186 = ~(n6838 | n12587);
assign n11043 = ~(n1730 ^ n7077);
assign n11290 = n10201 & n7204;
assign n2001 = ~(n4556 ^ n135);
assign n12322 = n3630 | n12328;
assign n4608 = n3986 | n5716;
assign n3489 = ~n10613;
assign n8874 = n6516 & n9085;
assign n5659 = n10696 | n9075;
assign n142 = ~n2370;
assign n5207 = ~(n7668 ^ n12232);
assign n8864 = ~n9270;
assign n10147 = n2057 & n10063;
assign n9728 = n4080 | n7723;
assign n5352 = n9309 | n8005;
assign n5113 = n5694 | n4947;
assign n6437 = ~(n2358 | n8462);
assign n11482 = n10928 ^ n4155;
assign n1895 = n7301 & n1274;
assign n4807 = n2800 & n2466;
assign n1032 = n11815 & n191;
assign n8737 = ~(n9173 ^ n13100);
assign n8064 = n6557 | n1570;
assign n10847 = ~(n11384 | n11141);
assign n2469 = n8639 | n10935;
assign n3206 = n13085 & n12696;
assign n9949 = n5358 | n5011;
assign n10423 = ~(n8628 ^ n1021);
assign n11065 = n5757 | n9147;
assign n4757 = n3158 | n4724;
assign n9708 = n9934 | n12388;
assign n5660 = n338 | n5076;
assign n7530 = n6210;
assign n108 = ~(n3841 ^ n1829);
assign n8215 = ~(n4507 | n1342);
assign n12526 = n8416 & n12590;
assign n650 = ~n8233;
assign n6388 = n7865 | n3149;
assign n6793 = n1353 | n9159;
assign n1357 = ~n3543;
assign n12068 = n5676 & n3530;
assign n7922 = ~(n2621 | n3220);
assign n4996 = ~(n11799 ^ n8669);
assign n866 = n1248 | n10878;
assign n5541 = ~(n966 | n7336);
assign n7257 = ~n5277;
assign n11608 = ~(n12682 ^ n9362);
assign n5301 = n11742 | n13125;
assign n12510 = n5415 | n167;
assign n5168 = ~n11734;
assign n6338 = n4370 | n8348;
assign n1502 = ~(n4383 ^ n3566);
assign n11723 = ~n4330;
assign n7531 = ~(n5224 ^ n37);
assign n9427 = ~(n9879 | n12983);
assign n10803 = ~(n5100 ^ n10185);
assign n7807 = n8064 | n6299;
assign n11635 = ~n7161;
assign n1376 = n2301 | n7476;
assign n11841 = n6139 & n6490;
assign n2553 = n1067 | n1195;
assign n12528 = n5265 | n10871;
assign n9613 = ~(n10219 ^ n11411);
assign n8738 = ~(n3357 | n3012);
assign n3377 = n6726 | n10179;
assign n2180 = ~(n2395 ^ n1615);
assign n10032 = ~n11734;
assign n1359 = n318 | n1985;
assign n4004 = n6572 & n5888;
assign n10717 = n4000 | n4223;
assign n4098 = ~n11640;
assign n13149 = n4161 | n2970;
assign n11250 = n4665 | n10871;
assign n4142 = ~(n1575 ^ n8622);
assign n3493 = ~n10860;
assign n6025 = ~n322;
assign n1320 = ~n11109;
assign n231 = n4969 | n3276;
assign n10180 = n6518 | n557;
assign n7069 = n654 & n230;
assign n2747 = ~n1397;
assign n13122 = ~n4376;
assign n10735 = ~(n2297 | n3421);
assign n2585 = ~(n3941 ^ n12658);
assign n13007 = n12846 & n12486;
assign n10278 = n11232 & n7243;
assign n6393 = n4771 | n12332;
assign n2356 = n12249 | n8563;
assign n5773 = n11010 | n9046;
assign n1774 = n11294 & n10748;
assign n1443 = ~(n4825 ^ n7165);
assign n2170 = ~(n12236 ^ n4835);
assign n882 = ~n6965;
assign n10248 = n8600 | n1804;
assign n10864 = ~(n5130 ^ n10113);
assign n9159 = n2406;
assign n3933 = n4587 | n9251;
assign n13102 = n9416 | n7203;
assign n5265 = ~n9669;
assign n6242 = n9934 | n1570;
assign n10358 = ~(n2878 | n12891);
assign n12556 = n5404 | n5721;
assign n2726 = ~n9475;
assign n11286 = n7836 | n11768;
assign n12197 = ~(n314 ^ n11253);
assign n1461 = ~(n5567 | n11563);
assign n1609 = n8449 & n1533;
assign n9071 = n12843 | n8988;
assign n4066 = ~n7745;
assign n175 = n2041 | n584;
assign n3793 = ~(n10765 | n852);
assign n1898 = ~(n5861 | n7548);
assign n4934 = n3364 | n11007;
assign n6402 = ~n11339;
assign n1091 = n4108 | n3554;
assign n3986 = n10761 | n6265;
assign n2002 = n5725 & n4451;
assign n2392 = n10180 & n10749;
assign n2485 = ~n624;
assign n3730 = n8615 | n4230;
assign n10616 = ~n2513;
assign n12064 = n12342 & n9977;
assign n4007 = ~(n976 | n260);
assign n11457 = n2570 & n6923;
assign n12314 = ~(n12809 ^ n11267);
assign n1509 = n9016 | n206;
assign n11512 = n12859 | n10971;
assign n4977 = ~(n1470 ^ n10614);
assign n4405 = n10598 & n4480;
assign n12957 = ~n937;
assign n1264 = n11799 | n3187;
assign n6177 = ~(n6196 ^ n12831);
assign n8408 = n10113 & n7411;
assign n4955 = ~n5454;
assign n8889 = ~(n4692 ^ n556);
assign n11502 = n544 | n322;
assign n7131 = n3522 | n8086;
assign n3009 = n2226 | n9309;
assign n10926 = n6027 & n6898;
assign n625 = n5638 & n6888;
assign n1214 = ~(n1297 ^ n6984);
assign n11944 = ~(n903 ^ n12197);
assign n8178 = ~(n2936 ^ n9356);
assign n6060 = n1238 & n3819;
assign n2609 = n5613 & n12555;
assign n967 = ~n5322;
assign n12218 = ~(n2101 ^ n4794);
assign n11769 = ~(n11971 ^ n12102);
assign n3602 = n8980 | n7509;
assign n8378 = n8862 | n12072;
assign n11993 = ~(n10861 ^ n6736);
assign n4853 = n1725 | n12948;
assign n2117 = n3837 & n6327;
assign n406 = ~n10657;
assign n12152 = ~(n7929 | n12106);
assign n11819 = ~(n783 ^ n8893);
assign n10776 = ~(n8135 ^ n11536);
assign n8645 = ~n11835;
assign n9486 = n7951 & n7921;
assign n5022 = ~(n7414 ^ n8845);
assign n237 = ~n10642;
assign n2240 = n10883 | n9075;
assign n9437 = n10419 ^ n2000;
assign n1669 = ~(n9676 ^ n11367);
assign n6191 = n202 | n1985;
assign n3690 = ~n880;
assign n8880 = n10591 | n7723;
assign n1658 = ~(n11496 | n7893);
assign n3866 = ~n3815;
assign n11536 = ~(n12140 ^ n3989);
assign n434 = n1651 | n4936;
assign n10101 = n10392 ^ n9655;
assign n6961 = n9154 | n12501;
assign n13022 = ~(n9637 ^ n3649);
assign n4074 = n3335 & n11178;
assign n2432 = ~(n4521 ^ n2497);
assign n7553 = ~(n2841 ^ n11528);
assign n3181 = ~(n11592 ^ n4656);
assign n1462 = ~(n7552 | n10793);
assign n2088 = n6375 | n10319;
assign n11484 = ~(n12581 ^ n12905);
assign n5037 = ~n4413;
assign n17 = n11683 | n10319;
assign n4888 = n9353 & n3085;
assign n5219 = ~(n12804 ^ n8594);
assign n11151 = ~(n1758 ^ n6034);
assign n7967 = ~(n1810 ^ n1755);
assign n11664 = ~n5375;
assign n9034 = ~(n2799 ^ n6544);
assign n2183 = ~n9591;
assign n4164 = n1906 & n6095;
assign n10683 = n9917 | n11446;
assign n9835 = n4370 | n4724;
assign n3039 = ~(n1352 | n8037);
assign n5782 = ~n411;
assign n12357 = ~n4015;
assign n250 = n11356 | n8702;
assign n10897 = n5456 & n8833;
assign n4695 = n1889 & n4320;
assign n4607 = n12911 | n2792;
assign n10511 = ~(n10217 ^ n2837);
assign n1824 = ~(n8067 | n10817);
assign n9954 = n8739 | n8036;
assign n8201 = ~(n7230 ^ n3622);
assign n11374 = n12758 | n4724;
assign n6765 = ~(n1601 ^ n7384);
assign n9161 = n12768 | n1570;
assign n3266 = n1772 | n7701;
assign n6702 = ~(n7852 ^ n1770);
assign n1546 = n6381 | n4947;
assign n12609 = n4891 & n6360;
assign n11183 = n1638 | n10029;
assign n5095 = ~(n5121 ^ n4516);
assign n7354 = n542 | n6265;
assign n7912 = ~(n11709 | n3447);
assign n6400 = ~(n5453 ^ n12836);
assign n3492 = n5407 | n3648;
assign n8417 = ~(n6535 | n4064);
assign n9254 = ~(n12467 | n9561);
assign n5277 = n6894 & n6980;
assign n4810 = n5182 | n11521;
assign n4249 = n5526 & n1691;
assign n12449 = n12617 | n9808;
assign n10342 = ~(n7802 ^ n5336);
assign n2101 = ~(n267 ^ n12762);
assign n8727 = ~(n5251 | n4065);
assign n3606 = ~(n890 ^ n7209);
assign n968 = n11113 | n9223;
assign n3784 = ~n12065;
assign n176 = ~(n1349 | n4259);
assign n2206 = ~(n6371 ^ n10071);
assign n3530 = n3460 | n12695;
assign n6047 = n7554 & n591;
assign n719 = ~n10745;
assign n10900 = ~n1364;
assign n2102 = n7514 & n7778;
assign n12467 = ~(n5005 | n13110);
assign n8348 = n3671;
assign n9310 = ~n5470;
assign n6447 = ~(n7256 ^ n832);
assign n651 = ~n9027;
assign n3633 = ~n6973;
assign n3854 = ~n353;
assign n5784 = n3225 | n8490;
assign n8275 = ~(n9033 | n5722);
assign n5847 = ~n6820;
assign n4756 = n9248 | n5006;
assign n1613 = ~(n3339 ^ n12878);
assign n3336 = ~n6189;
assign n4378 = n5911 & n3603;
assign n9839 = ~(n2994 ^ n8110);
assign n5531 = n10139 | n8101;
assign n4430 = ~n1225;
assign n11913 = ~(n11936 ^ n3252);
assign n10706 = ~(n1640 | n1704);
assign n10075 = n10738 & n11673;
assign n11416 = ~(n10385 ^ n3863);
assign n1258 = ~n6597;
assign n2806 = n872 | n7252;
assign n11943 = n7546 | n2490;
assign n9166 = ~(n10325 ^ n1929);
assign n445 = ~n5065;
assign n4716 = ~n8369;
assign n6150 = n11927 & n1300;
assign n3915 = n11263 | n13081;
assign n6752 = ~(n3171 | n5154);
assign n5694 = ~n3677;
assign n3143 = n3359 & n7570;
assign n784 = n930 | n10463;
assign n5255 = ~(n4304 | n11885);
assign n7155 = n316 & n4084;
assign n12414 = ~(n11793 ^ n11177);
assign n1468 = ~(n11534 | n3440);
assign n1402 = ~n10606;
assign n7736 = ~(n12013 ^ n8222);
assign n9807 = n6672 | n4420;
assign n875 = n13201 & n834;
assign n3225 = n6193;
assign n8950 = ~n11429;
assign n3563 = n13028 | n8777;
assign n3438 = ~(n11900 ^ n10816);
assign n3808 = ~(n2286 ^ n647);
assign n8068 = n7637 | n12171;
assign n6082 = n3800 & n10269;
assign n13176 = n11408 & n7911;
assign n9293 = n8865 | n8819;
assign n5719 = n5932 | n2633;
assign n351 = n4537 & n5962;
assign n4251 = n48 | n3981;
assign n4689 = ~n3797;
assign n12337 = n332 | n12733;
assign n1560 = n787 | n2059;
assign n3273 = n987 | n5242;
assign n10054 = ~(n11070 | n3503);
assign n9858 = ~(n8616 ^ n799);
assign n4484 = ~n919;
assign n11779 = ~n7659;
assign n8473 = ~(n2347 ^ n12346);
assign n5184 = n4356 & n4010;
assign n12069 = ~n11537;
assign n2748 = ~(n6750 | n7572);
assign n6141 = n11247 & n2812;
assign n1587 = ~n2498;
assign n9497 = ~n1563;
assign n12340 = n3498 | n10106;
assign n9405 = ~(n11215 | n2375);
assign n10955 = ~(n7882 ^ n1923);
assign n3551 = n6731 & n11901;
assign n6821 = n11513 & n312;
assign n9487 = n98 | n8702;
assign n1786 = n1645 | n6169;
assign n6467 = n3760 & n5446;
assign n4024 = n9387 & n9997;
assign n8080 = ~(n12270 ^ n1604);
assign n7127 = ~n7452;
assign n2022 = ~n5052;
assign n5529 = n7176 | n8366;
assign n12256 = n8891 | n3961;
assign n4208 = ~n12289;
assign n2159 = n7272 ^ n195;
assign n1845 = ~(n6322 ^ n10649);
assign n3388 = ~(n10829 | n6071);
assign n4662 = n11 & n8956;
assign n12905 = ~(n6314 ^ n8913);
assign n7696 = n10212 & n11947;
assign n7710 = ~n7906;
assign n4546 = n2795 & n11654;
assign n2421 = n4836 & n12883;
assign n3255 = n3505 | n9537;
assign n500 = n7782 | n4169;
assign n528 = n8940 & n8290;
assign n605 = n11914 & n12760;
assign n4121 = n3006 & n12853;
assign n3605 = n13154 | n6635;
assign n3679 = n5478 | n6293;
assign n1439 = n10974 | n8534;
assign n242 = ~(n7699 | n8703);
assign n8480 = n12942 & n475;
assign n12286 = ~(n9642 ^ n714);
assign n2264 = ~n10606;
assign n7754 = ~(n27 ^ n11353);
assign n1765 = n4221 | n3225;
assign n4696 = ~n4114;
assign n12524 = ~(n12829 ^ n6461);
assign n2910 = ~n5075;
assign n10097 = n12024 | n8568;
assign n3231 = n6168 & n4470;
assign n10497 = n11218 | n2958;
assign n5102 = ~(n8807 ^ n12275);
assign n1427 = n5679 | n11107;
assign n2009 = ~(n2533 ^ n8042);
assign n1151 = ~n4303;
assign n5218 = n6926 & n4418;
assign n5872 = n10893 | n6364;
assign n385 = n12032 | n12388;
assign n12039 = ~(n6828 ^ n4917);
assign n12390 = n7371 & n8438;
assign n6941 = ~(n4965 | n339);
assign n2850 = n877 | n11898;
assign n7094 = ~(n707 ^ n4307);
assign n8848 = ~n6021;
assign n11830 = ~(n11584 ^ n9738);
assign n11532 = ~(n7236 | n2099);
assign n960 = ~(n7618 ^ n4617);
assign n638 = n1896 & n11005;
assign n3124 = n924 | n5776;
assign n775 = ~(n11046 ^ n6030);
assign n8661 = ~n7161;
assign n3847 = n572 | n11375;
assign n6348 = n12878 | n8118;
assign n5911 = n12082 | n4786;
assign n6778 = n8681 | n5797;
assign n13196 = n11054 | n1463;
assign n12383 = ~n834;
assign n10753 = n9674 | n1255;
assign n4480 = n2487 | n5242;
assign n3332 = ~(n3139 ^ n9470);
assign n9463 = ~(n5737 | n7643);
assign n9290 = n9259 & n7355;
assign n10895 = n12768 | n6265;
assign n3044 = ~n10102;
assign n1795 = ~n7500;
assign n256 = n2394 & n5096;
assign n12440 = ~(n7403 ^ n4034);
assign n35 = n3707 | n5207;
assign n9605 = n549 | n5;
assign n1155 = ~n1910;
assign n6368 = n10828 & n3346;
assign n11875 = ~(n8302 ^ n7366);
assign n8502 = n11493 & n5529;
assign n1090 = ~(n371 ^ n439);
assign n7671 = ~(n7699 ^ n874);
assign n11397 = n11055 ^ n139;
assign n11870 = n8390 & n2076;
assign n4181 = ~(n1166 | n5525);
assign n9625 = n12808 | n8857;
assign n12674 = n10217 | n6442;
assign n11851 = n12084 & n13054;
assign n6353 = ~(n1716 ^ n835);
assign n13054 = ~(n12941 ^ n1992);
assign n1626 = n10404 | n3997;
assign n6339 = ~(n3388 | n12140);
assign n9400 = ~n2252;
assign n9396 = ~n4797;
assign n9833 = n2809 & n9013;
assign n2487 = ~n1724;
assign n11260 = n968 | n2923;
assign n3037 = n9160 & n2335;
assign n9618 = ~n9952;
assign n7450 = n5313 | n12973;
assign n8905 = ~n3644;
assign n6710 = ~n4452;
assign n2132 = n4600 | n1723;
assign n12918 = n1425 | n11689;
assign n8347 = n9003 & n1606;
assign n11966 = ~(n3427 | n3949);
assign n8935 = ~n12553;
assign n12421 = n3528 & n10918;
assign n9852 = ~(n11206 ^ n1845);
assign n11120 = n2538 | n2059;
assign n11404 = ~n12482;
assign n11015 = n4228 | n12684;
assign n8224 = ~(n9860 ^ n1761);
assign n4195 = ~(n3061 ^ n13192);
assign n6031 = ~(n12603 ^ n1910);
assign n3719 = ~n12461;
assign n10005 = ~n5319;
assign n3452 = ~(n11964 | n10766);
assign n1285 = ~(n11736 ^ n12015);
assign n10421 = ~n9915;
assign n6936 = n3822 | n3339;
assign n369 = ~(n5514 ^ n7916);
assign n659 = ~(n12690 ^ n7511);
assign n4086 = n93 & n10113;
assign n11581 = n3016 & n7018;
assign n1989 = ~n9041;
assign n7823 = n10794 & n10131;
assign n4194 = ~n8230;
assign n2834 = n10731 | n5485;
assign n1253 = ~(n5475 ^ n974);
assign n5263 = ~(n347 ^ n6797);
assign n12435 = n6970 | n4445;
assign n2437 = ~n1055;
assign n6370 = ~n9732;
assign n1530 = n4380 & n10093;
assign n8639 = n9190 & n3532;
assign n9398 = n12580 | n4834;
assign n12020 = ~(n4084 ^ n316);
assign n12192 = n3281 | n4116;
assign n1918 = n8926 | n5736;
assign n5114 = n4371 & n4078;
assign n924 = ~(n7706 ^ n679);
assign n6131 = n5271 | n1026;
assign n11811 = n10274 | n11527;
assign n3109 = n7872 | n8563;
assign n3522 = n5482 | n1303;
assign n7370 = n6106 | n5986;
assign n11299 = ~(n11832 ^ n4040);
assign n2407 = n10517 | n11735;
assign n10428 = n10029 | n8030;
assign n8687 = n1975 | n6454;
assign n6852 = ~(n2519 ^ n8591);
assign n10457 = n2458 & n12306;
assign n9177 = ~n10455;
assign n8973 = n9635 | n3455;
assign n4107 = ~n5962;
assign n9593 = ~(n11783 | n12079);
assign n4023 = n4580 & n12844;
assign n7301 = n9364 | n4300;
assign n7966 = ~n4357;
assign n11376 = n6769 | n177;
assign n8634 = n5679 | n8030;
assign n787 = ~n6818;
assign n12976 = ~(n3375 ^ n480);
assign n362 = ~(n6930 ^ n9031);
assign n6083 = ~(n13227 ^ n2770);
assign n7891 = n2276 | n5430;
assign n12767 = n8593 & n565;
assign n4005 = n6438 | n11668;
assign n11339 = n1963 & n1008;
assign n2805 = ~(n6831 ^ n5967);
assign n2410 = ~(n3705 | n13177);
assign n2793 = ~n102;
assign n9914 = n7647 | n10387;
assign n12513 = ~(n9807 ^ n12790);
assign n2343 = ~(n2146 ^ n9163);
assign n1871 = n7792 ^ n6851;
assign n11619 = ~(n1169 | n5620);
assign n2658 = ~(n3696 ^ n4885);
assign n782 = n4480 | n10598;
assign n2086 = n4772 | n12495;
assign n10618 = n7313 | n2931;
assign n8156 = ~(n577 ^ n780);
assign n2914 = n11729 | n7723;
assign n9074 = n5671 & n5536;
assign n143 = ~(n562 ^ n6398);
assign n10493 = n5103 & n3768;
assign n9961 = ~(n12989 ^ n7143);
assign n410 = n7205 | n9985;
assign n12515 = ~(n8647 ^ n4168);
assign n1625 = ~n3841;
assign n8313 = n9931 | n4373;
assign n1759 = n5679 | n10871;
assign n4312 = n8139 & n9906;
assign n7293 = n5261 | n9223;
assign n832 = n6659 & n9071;
assign n1541 = ~(n2182 ^ n5278);
assign n235 = ~n8742;
assign n5091 = n13026 | n7961;
assign n5156 = ~(n2598 ^ n10985);
assign n10346 = n9843 | n11394;
assign n41 = ~(n12771 | n5538);
assign n9036 = ~(n10378 ^ n4249);
assign n3024 = n11328 | n3763;
assign n4856 = ~(n10639 ^ n2921);
assign n3027 = ~(n12222 | n4336);
assign n7263 = ~(n9294 ^ n212);
assign n10193 = ~(n4978 | n9821);
assign n1484 = n10060 & n6866;
assign n10978 = ~n9609;
assign n2049 = n5148 | n4724;
assign n6997 = ~(n3934 ^ n2414);
assign n527 = n6245 | n6769;
assign n13239 = ~n6487;
assign n12292 = n1144 | n10871;
assign n6126 = n8805 & n11648;
assign n4243 = ~n2258;
assign n9459 = ~(n870 ^ n11604);
assign n12797 = ~(n8546 ^ n1585);
assign n955 = ~(n1599 ^ n4478);
assign n6371 = n8757 | n8490;
assign n10282 = ~(n518 | n7776);
assign n139 = n937 & n8506;
assign n11824 = n4065 & n5251;
assign n5010 = n12475 | n3759;
assign n831 = ~(n3953 ^ n796);
assign n262 = ~(n6993 | n3506);
assign n3108 = ~(n1067 ^ n12303);
assign n7044 = n11061 & n8506;
assign n6232 = ~n12255;
assign n9217 = n10705 | n2561;
assign n11283 = n97 | n1043;
assign n12043 = ~n10091;
assign n12729 = ~(n5158 ^ n3861);
assign n11226 = ~n5884;
assign n6905 = n8196 & n11269;
assign n1577 = ~n2827;
assign n9370 = ~(n5062 | n7262);
assign n11939 = ~(n1653 ^ n10307);
assign n109 = n2464 ^ n8123;
assign n10533 = n2689 | n10179;
assign n3858 = ~n5671;
assign n5675 = ~(n336 ^ n7290);
assign n12085 = ~(n5738 ^ n7365);
assign n8281 = ~(n5704 ^ n10194);
assign n591 = ~n140;
assign n4559 = n4155 & n3437;
assign n12714 = ~(n10873 | n8419);
assign n1110 = ~(n5452 ^ n12307);
assign n12657 = ~n1364;
assign n7295 = n3194 | n4680;
assign n1983 = ~(n7772 ^ n7529);
assign n5321 = n4454 | n8268;
assign n12297 = ~n11589;
assign n654 = n1719 | n2686;
assign n691 = n11966;
assign n819 = n10203 & n5234;
assign n10240 = ~n5548;
assign n1147 = ~(n983 ^ n1272);
assign n3073 = ~(n9399 ^ n11841);
assign n10645 = ~(n6168 | n11411);
assign n2175 = ~n40;
assign n12847 = n11940;
assign n341 = n52 & n144;
assign n10708 = n866 & n10428;
assign n2804 = ~(n11659 | n12945);
assign n6163 = ~(n38 | n7923);
assign n2876 = ~(n2991 ^ n9440);
assign n791 = ~(n9684 ^ n12691);
assign n3578 = ~(n5789 ^ n5437);
assign n11506 = ~(n2982 ^ n11764);
assign n12816 = n9773 & n4576;
assign n6115 = ~(n10429 ^ n252);
assign n5561 = n542 | n7935;
assign n12884 = n12897 & n5133;
assign n9638 = ~n10642;
assign n11792 = ~(n4188 ^ n427);
assign n5357 = n11202 & n1117;
assign n9495 = ~(n5018 ^ n4477);
assign n10608 = n10978 | n11008;
assign n154 = ~n8820;
assign n3134 = ~(n11303 ^ n8572);
assign n2846 = ~(n5440 ^ n2244);
assign n8931 = ~(n2298 ^ n1757);
assign n3427 = ~n854;
assign n7755 = ~(n9769 ^ n11388);
assign n3102 = ~n3863;
assign n7828 = n7825 | n1144;
assign n11019 = ~(n7759 ^ n3200);
assign n11304 = ~(n10395 | n102);
assign n1860 = ~(n3144 ^ n9090);
assign n6803 = n8315 | n12847;
assign n5304 = ~(n4317 ^ n5405);
assign n3638 = n5191 | n4070;
assign n10852 = n10625 & n10160;
assign n10745 = ~(n11215 ^ n8214);
assign n6365 = ~(n6954 ^ n1556);
assign n5462 = ~n873;
assign n8122 = ~n7863;
assign n6887 = n2329 | n177;
assign n10675 = ~(n6123 ^ n3420);
assign n11247 = n2832 | n9943;
assign n3082 = ~n1466;
assign n3762 = ~(n9841 ^ n12219);
assign n3224 = ~(n11178 ^ n3335);
assign n6674 = n5158 | n3913;
assign n11687 = ~(n11877 ^ n10566);
assign n5977 = n8909 & n3004;
assign n8109 = n2080 | n13117;
assign n3745 = ~(n3611 ^ n13155);
assign n8817 = ~n7113;
assign n731 = ~(n1424 ^ n1693);
assign n13027 = n6416 | n121;
assign n12419 = ~(n11397 ^ n12903);
assign n2767 = n4536 | n7430;
assign n5220 = n8188 | n2738;
assign n10223 = n1092 & n891;
assign n2753 = ~(n11608 ^ n4894);
assign n8475 = ~(n9211 | n8767);
assign n4671 = ~(n12730 ^ n328);
assign n7580 = n11723 | n2222;
assign n12702 = n12765 | n11447;
assign n6757 = ~n6809;
assign n675 = ~(n8779 ^ n5828);
assign n3670 = ~(n6229 ^ n6263);
assign n10932 = n10938 & n1841;
assign n3226 = ~(n11129 ^ n11052);
assign n7026 = n6202 | n721;
assign n10375 = n5016 | n4172;
assign n12862 = ~(n8036 ^ n12852);
assign n4774 = n602 ^ n10654;
assign n8074 = n12732 | n121;
assign n12359 = n12780 & n2413;
assign n3449 = ~(n12078 ^ n4798);
assign n10509 = ~n10142;
assign n494 = n7819 | n12383;
assign n7317 = n10195 | n12691;
assign n6044 = ~(n6811 | n11364);
assign n2602 = n8230 & n12289;
assign n4828 = n10068 | n12173;
assign n11625 = n6986 | n2059;
assign n9866 = ~(n12341 ^ n8027);
assign n12506 = ~(n2865 ^ n3548);
assign n8155 = n7541 ^ n1953;
assign n2856 = n4890 | n6265;
assign n10760 = n4412 | n8679;
assign n10880 = n8802 | n6235;
assign n5437 = n9501 | n1044;
assign n11812 = ~(n3317 ^ n7812);
assign n7401 = n4107 | n11144;
assign n8519 = ~(n1610 | n10605);
assign n7407 = ~n12746;
assign n7606 = n10941 | n12746;
assign n11110 = ~n6213;
assign n12890 = ~(n12019 ^ n620);
assign n4895 = ~(n10815 ^ n8791);
assign n11755 = ~(n6785 ^ n8691);
assign n11852 = ~(n7711 ^ n9756);
assign n7329 = n5328 | n1463;
assign n8276 = ~(n3405 | n6752);
assign n8143 = ~n9915;
assign n6265 = n138;
assign n9504 = ~(n2974 ^ n788);
assign n13200 = n6189 & n9092;
assign n12429 = ~(n5384 ^ n4296);
assign n1260 = ~(n8203 ^ n315);
assign n7504 = n1250 & n3113;
assign n10334 = ~n8163;
assign n11685 = n8533 & n2515;
assign n3216 = n11091 | n12665;
assign n4466 = n5808 | n3135;
assign n3463 = ~(n9856 ^ n313);
assign n5436 = n1747 | n11423;
assign n11345 = n2738 | n7935;
assign n6584 = n4937 | n978;
assign n1081 = ~(n8647 | n3702);
assign n11215 = n813 | n1144;
assign n7343 = ~(n8043 ^ n814);
assign n5833 = n3509 | n6635;
assign n5471 = ~(n7751 | n7093);
assign n5512 = n12135 | n6714;
assign n2300 = ~(n6747 ^ n6553);
assign n198 = ~n1667;
assign n6456 = n6428 & n839;
assign n305 = n3594 & n4632;
assign n7395 = ~n10567;
assign n10921 = ~(n5982 ^ n10827);
assign n11689 = n7640 & n12697;
assign n9072 = n5892 | n5942;
assign n2760 = ~(n12462 ^ n5092);
assign n5883 = n2734 | n9921;
assign n11322 = n6837 | n11166;
assign n6916 = n13227 | n11028;
assign n13190 = ~n4357;
assign n10326 = ~(n3725 ^ n263);
assign n8050 = ~n10782;
assign n4621 = ~n5920;
assign n4374 = ~(n8433 ^ n441);
assign n28 = ~(n6624 ^ n4993);
assign n10444 = n5100 & n8837;
assign n11749 = n8053 | n7935;
assign n420 = n11488 & n12853;
assign n11705 = n8529 | n7935;
assign n11623 = ~(n11648 ^ n2627);
assign n656 = ~n3713;
assign n3554 = n12573 | n1463;
assign n7685 = ~(n5404 ^ n4739);
assign n8497 = ~(n2358 ^ n2009);
assign n6018 = n3158 | n12957;
assign n11957 = n640 | n1808;
assign n12331 = ~(n13208 ^ n7070);
assign n1063 = ~(n9271 ^ n3925);
assign n7404 = n1290 | n9151;
assign n2769 = n10825 | n6869;
assign n9111 = ~(n9488 ^ n2114);
assign n8925 = ~n209;
assign n8251 = ~n9452;
assign n11218 = ~n854;
assign n5955 = ~(n12429 ^ n5815);
assign n2318 = n4191 | n5074;
assign n7471 = ~n6644;
assign n1938 = n5562 | n9075;
assign n1038 = n3164 & n8928;
assign n4568 = ~(n4710 ^ n2313);
assign n3195 = ~n4304;
assign n9280 = ~n6333;
assign n3675 = ~(n11082 | n627);
assign n10791 = ~(n451 ^ n1680);
assign n8806 = ~(n8650 | n13023);
assign n4323 = ~(n5203 | n309);
assign n4217 = n6225 | n12717;
assign n2635 = ~(n11363 | n10539);
assign n371 = n542 | n12388;
assign n10178 = ~n11169;
assign n7087 = n2264 | n5242;
assign n12088 = ~n13069;
assign n5325 = ~(n2971 ^ n6684);
assign n8405 = n2968 | n4018;
assign n3919 = n3002 & n11223;
assign n13049 = n4317 | n11549;
assign n4408 = ~(n7364 | n219);
assign n3487 = ~(n4994 ^ n12305);
assign n6689 = ~n3130;
assign n1900 = n1484 ^ n9771;
assign n6493 = n12597 & n9834;
assign n13057 = ~(n11709 ^ n3447);
assign n5457 = n7194 & n7801;
assign n8692 = ~(n11577 | n9408);
assign n9640 = ~(n9467 ^ n13158);
assign n4356 = n10075 | n7737;
assign n7679 = n7593 | n2753;
assign n7954 = n10336 & n6771;
assign n11417 = ~(n7066 ^ n9156);
assign n9926 = n9478 | n479;
assign n7718 = ~n9475;
assign n1221 = ~(n6864 ^ n7562);
assign n13076 = n12098 & n11787;
assign n9246 = ~(n7897 ^ n889);
assign n4265 = n3178 & n1007;
assign n7641 = n1649 & n4263;
assign n2622 = ~n5536;
assign n42 = ~n3527;
assign n8797 = ~(n8908 | n8376);
assign n7443 = ~n9839;
assign n7766 = ~(n7380 ^ n10156);
assign n5862 = n1888 | n3224;
assign n8243 = ~n12809;
assign n1314 = n11651 | n4505;
assign n9922 = ~(n3659 ^ n7053);
assign n6423 = n12496 | n6093;
assign n2305 = n12266 | n11625;
assign n151 = n9193 | n12287;
assign n2447 = n9358 ^ n3720;
assign n5421 = ~(n992 ^ n12319);
assign n10539 = n12652 & n12699;
assign n10787 = ~(n1326 ^ n11406);
assign n11000 = n4784 & n4493;
assign n5288 = ~(n5403 ^ n9800);
assign n9889 = ~n13078;
assign n465 = ~(n2903 ^ n10922);
assign n254 = n9926 | n5175;
assign n8422 = ~(n12117 ^ n12594);
assign n5892 = n7661 | n4936;
assign n8464 = n6223 | n10871;
assign n13179 = ~(n5881 ^ n8281);
assign n483 = ~(n12826 ^ n5761);
assign n3351 = ~(n1592 ^ n3850);
assign n6930 = ~(n8230 ^ n6668);
assign n1631 = n5541 | n6234;
assign n1686 = n7871 & n6975;
assign n5025 = n3564 | n11107;
assign n4009 = ~(n10906 ^ n9905);
assign n8307 = n13144 | n6905;
assign n3375 = ~(n10765 ^ n6662);
assign n10501 = ~n7720;
assign n344 = n2877 | n12388;
assign n4030 = ~n1288;
assign n5638 = ~n4671;
assign n261 = ~(n9222 ^ n1348);
assign n9015 = n1262 | n2986;
assign n7376 = ~(n6611 ^ n3605);
assign n2838 = ~n4186;
assign n3164 = n1872 | n11995;
assign n4216 = n1480 | n902;
assign n13017 = ~n12228;
assign n13136 = ~(n2749 | n10515);
assign n11378 = n1930 | n8268;
assign n13188 = ~(n5428 ^ n9774);
assign n33 = ~(n6395 ^ n7148);
assign n6330 = ~n11544;
assign n1080 = ~n9918;
assign n12063 = n137 | n4636;
assign n3711 = ~(n503 ^ n9820);
assign n2623 = ~n3178;
assign n7796 = ~(n1033 | n4127);
assign n7136 = ~(n3993 | n2007);
assign n5164 = n2657 | n3949;
assign n5197 = n4484 & n11540;
assign n211 = n10680 ^ n4121;
assign n1135 = ~n9041;
assign n2217 = ~n1231;
assign n11456 = ~(n4954 | n8162);
assign n3170 = ~(n10855 ^ n3547);
assign n10568 = ~(n668 ^ n2543);
assign n518 = n3908 | n4640;
assign n7062 = ~n7374;
assign n8764 = n5660 | n2319;
assign n5279 = ~n7514;
assign n9127 = ~(n8060 ^ n10169);
assign n11386 = n8729 | n4640;
assign n2823 = n11941 | n2133;
assign n3360 = n10383 | n4724;
assign n291 = ~(n7105 ^ n13009);
assign n12353 = n7718 | n4947;
assign n9449 = ~(n11289 ^ n13114);
assign n12288 = n9496 | n8034;
assign n11694 = ~(n6965 ^ n2488);
assign n9774 = ~(n1828 ^ n4403);
assign n10115 = ~(n2643 | n4629);
assign n6902 = n3035 & n8590;
assign n10490 = n9131 | n1144;
assign n4188 = n9849 ^ n11866;
assign n9844 = ~(n7594 ^ n7512);
assign n6245 = ~n4419;
assign n3838 = ~(n4291 ^ n2256);
assign n333 = ~n11488;
assign n6862 = ~(n12051 ^ n7663);
assign n11463 = n12293 | n2044;
assign n13140 = n4339 | n170;
assign n4273 = ~(n3535 ^ n393);
assign n11905 = n8385 & n12431;
assign n184 = ~(n13197 ^ n8945);
assign n7288 = ~(n3933 ^ n10669);
assign n8048 = n2657 | n3149;
assign n6041 = ~n11537;
assign n7675 = ~n7411;
assign n12717 = ~n2590;
assign n3015 = ~(n11744 ^ n4235);
assign n4822 = n8113 | n7032;
assign n12392 = n12441 | n6814;
assign n8741 = n8420 | n1866;
assign n12084 = ~(n11508 ^ n6623);
assign n12091 = ~(n7829 ^ n5532);
assign n3735 = ~(n781 ^ n4582);
assign n8569 = ~n1757;
assign n6208 = ~(n9243 | n2245);
assign n3754 = ~(n12484 ^ n1957);
assign n4867 = ~(n5539 ^ n12444);
assign n3072 = ~(n3389 ^ n9374);
assign n11097 = n4835 & n12236;
assign n12269 = ~(n4396 ^ n8612);
assign n1949 = n4754 & n3533;
assign n7566 = n8561 | n10871;
assign n8899 = n13130 | n8828;
assign n3120 = n8158 | n11719;
assign n4517 = ~n10113;
assign n10702 = ~(n968 ^ n2923);
assign n3900 = n2892 & n108;
assign n8985 = ~n160;
assign n10890 = ~n9324;
assign n10873 = n13122 & n11813;
assign n6501 = n7327 | n11841;
assign n8669 = ~n3187;
assign n8257 = n10313 | n1782;
assign n5591 = ~(n2750 ^ n8824);
assign n5576 = ~(n2238 ^ n12248);
assign n3712 = ~n3973;
assign n10483 = n5527 & n3831;
assign n8102 = n10668 & n5141;
assign n1596 = n7427 | n7534;
assign n11925 = n7159 & n4928;
assign n8744 = ~n8139;
assign n8966 = ~(n2534 ^ n11467);
assign n9715 = n10891 & n5653;
assign n10967 = n7960 & n12819;
assign n3920 = n8845 & n7414;
assign n9200 = ~(n9967 | n1442);
assign n10226 = ~(n7937 | n7721);
assign n5527 = ~n912;
assign n8175 = ~n6083;
assign n5323 = n5713 | n10029;
assign n5310 = ~n13047;
assign n7178 = ~(n9701 ^ n7009);
assign n12868 = n5044 | n12860;
assign n2510 = n3493 & n1085;
assign n2294 = ~n3005;
assign n12858 = ~n4350;
endmodule
