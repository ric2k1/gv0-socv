module top( 2_n11 , 2_n21 , 2_n22 , 2_n23 , 2_n27 , 2_n29 , 2_n30 , 2_n40 , 2_n45 , 2_n50 , 2_n52 , 2_n54 , 2_n56 , 2_n58 , 2_n71 , 2_n77 , 2_n82 , 2_n85 , 2_n86 , 2_n87 , 2_n94 , 2_n107 , 2_n112 , 2_n117 , 2_n126 , 2_n130 , 2_n138 , 2_n143 , 2_n153 , 2_n155 , 2_n156 , 2_n159 , 2_n161 , 2_n164 , 2_n173 , 2_n181 , 2_n184 , 2_n200 , 2_n216 , 2_n219 , 2_n220 , 2_n222 , 2_n223 , 2_n230 , 2_n233 , 2_n243 , 2_n244 , 2_n246 , 2_n247 , 2_n251 , 2_n254 , 2_n262 , 2_n268 , 2_n273 , 2_n275 , 2_n284 , 2_n288 , 2_n292 , 2_n293 , 2_n299 , 2_n300 , 2_n301 , 2_n304 , 2_n307 , 2_n310 , 2_n312 , 2_n314 , 2_n315 , 2_n318 , 2_n337 , 2_n341 , 2_n344 , 2_n346 , 2_n352 , 2_n362 , 2_n364 , 2_n370 , 2_n374 , 2_n376 , 2_n378 , 2_n380 , 2_n391 , 2_n392 , 2_n396 , 2_n399 , 2_n408 , 2_n409 , 2_n416 , 2_n417 , 2_n420 , 2_n428 , 2_n430 , 2_n453 , 2_n457 , 2_n460 , 2_n477 , 2_n478 , 2_n487 , 2_n489 , 2_n497 , 2_n498 , 2_n501 , 2_n502 , 2_n506 , 2_n507 , 2_n509 , 2_n510 , 2_n516 , 2_n517 , 2_n534 , 2_n545 , 2_n553 , 2_n559 , 2_n560 , 2_n561 , 2_n567 , 2_n574 , 2_n581 , 2_n582 , 2_n585 , 2_n589 , 2_n593 , 2_n595 , 2_n597 , 2_n598 , 2_n600 , 2_n607 , 2_n608 , 2_n609 , 2_n625 , 2_n626 , 2_n638 , 2_n640 , 2_n641 , 2_n645 , 2_n663 , 2_n669 , 2_n671 , 2_n676 , 2_n690 , 2_n693 , 2_n695 , 2_n701 , 2_n710 , 2_n714 , 2_n719 , 2_n726 , 2_n727 , 2_n729 , 2_n734 , 2_n742 , 2_n743 , 2_n755 , 2_n769 , 2_n773 , 2_n775 , 2_n778 , 2_n779 , 2_n782 , 2_n787 , 2_n790 , 2_n794 , 2_n821 , 2_n823 , 2_n831 , 2_n832 , 2_n839 , 2_n842 , 2_n849 , 2_n879 , 2_n882 , 2_n885 , 2_n894 , 2_n905 , 2_n916 , 2_n918 , 2_n920 , 2_n936 , 2_n947 , 2_n952 , 2_n953 , 2_n961 , 2_n969 , 2_n980 , 2_n984 , 2_n986 , 2_n990 , 2_n992 , 2_n997 , 2_n1006 , 2_n1017 , 2_n1023 , 2_n1040 , 2_n1042 , 2_n1044 , 2_n1050 , 2_n1051 , 2_n1054 , 2_n1058 , 2_n1060 , 2_n1061 , 2_n1063 , 2_n1065 , 2_n1071 , 2_n1095 , 2_n1103 , 2_n1114 , 2_n1121 , 2_n1138 , 2_n1152 , 2_n1154 , 2_n1156 , 2_n1164 , 2_n1172 , 2_n1175 , 2_n1177 , 2_n1186 , 2_n1187 , 2_n1191 , 2_n1193 , 2_n1195 , 2_n1205 , 2_n1209 , 2_n1211 , 2_n1225 , 2_n1227 , 2_n1231 , 2_n1234 , 2_n1239 , 2_n1246 , 2_n1250 , 2_n1253 , 2_n1263 , 2_n1278 , 2_n1281 , 2_n1283 , 2_n1285 , 2_n1286 , 2_n1288 , 2_n1289 , 2_n1292 , 2_n1296 , 2_n1299 , 2_n1301 , 2_n1302 , 2_n1305 , 2_n1306 , 2_n1320 , 2_n1322 , 2_n1337 , 2_n1345 , 2_n1346 , 2_n1350 , 2_n1359 , 2_n1361 , 2_n1368 , 2_n1375 , 2_n1386 , 2_n1387 , 2_n1389 , 2_n1391 , 2_n1393 , 2_n1401 , 2_n1411 , 2_n1415 , 2_n1418 , 2_n1420 , 2_n1421 , 2_n1427 , 2_n1428 , 2_n1435 , 2_n1438 , 2_n1443 , 2_n1446 , 2_n1448 , 2_n1463 , 2_n1470 , 2_n1474 , 2_n1476 , 2_n1500 , 2_n1502 , 2_n1506 , 2_n1516 , 2_n1520 , 2_n1521 , 2_n1523 , 2_n1527 , 2_n1534 , 2_n1536 , 2_n1547 , 2_n1548 , 2_n1566 , 2_n1569 , 2_n1576 , 2_n1586 , 2_n1588 , 2_n1592 , 2_n1594 , 2_n1609 , 2_n1613 , 2_n1616 , 2_n1626 , 2_n1627 , 2_n1632 , 2_n1639 , 2_n1644 , 2_n1645 , 2_n1647 , 2_n1656 , 2_n1687 , 2_n1729 , 2_n1738 , 2_n1750 , 2_n1752 , 2_n1753 );
    input 2_n11 , 2_n21 , 2_n29 , 2_n40 , 2_n45 , 2_n50 , 2_n52 , 2_n54 , 2_n56 , 2_n58 , 2_n71 , 2_n77 , 2_n82 , 2_n86 , 2_n87 , 2_n94 , 2_n107 , 2_n117 , 2_n138 , 2_n143 , 2_n153 , 2_n155 , 2_n156 , 2_n159 , 2_n200 , 2_n219 , 2_n220 , 2_n222 , 2_n223 , 2_n243 , 2_n244 , 2_n246 , 2_n251 , 2_n254 , 2_n262 , 2_n268 , 2_n273 , 2_n284 , 2_n288 , 2_n293 , 2_n299 , 2_n300 , 2_n307 , 2_n310 , 2_n312 , 2_n314 , 2_n315 , 2_n318 , 2_n341 , 2_n344 , 2_n346 , 2_n374 , 2_n376 , 2_n380 , 2_n391 , 2_n392 , 2_n399 , 2_n408 , 2_n409 , 2_n416 , 2_n420 , 2_n430 , 2_n477 , 2_n478 , 2_n487 , 2_n489 , 2_n502 , 2_n506 , 2_n507 , 2_n510 , 2_n545 , 2_n559 , 2_n560 , 2_n561 , 2_n567 , 2_n574 , 2_n581 , 2_n582 , 2_n589 , 2_n593 , 2_n598 , 2_n600 , 2_n607 , 2_n608 , 2_n609 , 2_n626 , 2_n641 , 2_n645 , 2_n663 , 2_n671 , 2_n676 , 2_n690 , 2_n695 , 2_n701 , 2_n710 , 2_n727 , 2_n729 , 2_n734 , 2_n742 , 2_n743 , 2_n755 , 2_n769 , 2_n775 , 2_n778 , 2_n779 , 2_n787 , 2_n790 , 2_n823 , 2_n831 , 2_n832 , 2_n839 , 2_n849 , 2_n879 , 2_n882 , 2_n885 , 2_n905 , 2_n920 , 2_n936 , 2_n947 , 2_n953 , 2_n961 , 2_n969 , 2_n980 , 2_n984 , 2_n986 , 2_n992 , 2_n997 , 2_n1023 , 2_n1040 , 2_n1044 , 2_n1054 , 2_n1061 , 2_n1071 , 2_n1095 , 2_n1103 , 2_n1114 , 2_n1121 , 2_n1138 , 2_n1152 , 2_n1154 , 2_n1156 , 2_n1164 , 2_n1172 , 2_n1175 , 2_n1187 , 2_n1191 , 2_n1193 , 2_n1205 , 2_n1225 , 2_n1227 , 2_n1239 , 2_n1246 , 2_n1250 , 2_n1263 , 2_n1278 , 2_n1281 , 2_n1283 , 2_n1286 , 2_n1289 , 2_n1299 , 2_n1301 , 2_n1305 , 2_n1345 , 2_n1346 , 2_n1350 , 2_n1361 , 2_n1386 , 2_n1387 , 2_n1389 , 2_n1393 , 2_n1401 , 2_n1411 , 2_n1415 , 2_n1418 , 2_n1428 , 2_n1435 , 2_n1438 , 2_n1443 , 2_n1446 , 2_n1448 , 2_n1463 , 2_n1470 , 2_n1474 , 2_n1476 , 2_n1500 , 2_n1502 , 2_n1506 , 2_n1516 , 2_n1520 , 2_n1521 , 2_n1523 , 2_n1536 , 2_n1566 , 2_n1569 , 2_n1576 , 2_n1586 , 2_n1592 , 2_n1609 , 2_n1613 , 2_n1616 , 2_n1626 , 2_n1627 , 2_n1644 , 2_n1647 , 2_n1656 , 2_n1750 , 2_n1753 ;
    output 2_n22 , 2_n23 , 2_n27 , 2_n30 , 2_n85 , 2_n112 , 2_n126 , 2_n130 , 2_n161 , 2_n164 , 2_n173 , 2_n181 , 2_n184 , 2_n216 , 2_n230 , 2_n233 , 2_n247 , 2_n275 , 2_n292 , 2_n301 , 2_n304 , 2_n337 , 2_n352 , 2_n362 , 2_n364 , 2_n370 , 2_n378 , 2_n396 , 2_n417 , 2_n428 , 2_n453 , 2_n457 , 2_n460 , 2_n497 , 2_n498 , 2_n501 , 2_n509 , 2_n516 , 2_n517 , 2_n534 , 2_n553 , 2_n585 , 2_n595 , 2_n597 , 2_n625 , 2_n638 , 2_n640 , 2_n669 , 2_n693 , 2_n714 , 2_n719 , 2_n726 , 2_n773 , 2_n782 , 2_n794 , 2_n821 , 2_n842 , 2_n894 , 2_n916 , 2_n918 , 2_n952 , 2_n990 , 2_n1006 , 2_n1017 , 2_n1042 , 2_n1050 , 2_n1051 , 2_n1058 , 2_n1060 , 2_n1063 , 2_n1065 , 2_n1177 , 2_n1186 , 2_n1195 , 2_n1209 , 2_n1211 , 2_n1231 , 2_n1234 , 2_n1253 , 2_n1285 , 2_n1288 , 2_n1292 , 2_n1296 , 2_n1302 , 2_n1306 , 2_n1320 , 2_n1322 , 2_n1337 , 2_n1359 , 2_n1368 , 2_n1375 , 2_n1391 , 2_n1420 , 2_n1421 , 2_n1427 , 2_n1527 , 2_n1534 , 2_n1547 , 2_n1548 , 2_n1588 , 2_n1594 , 2_n1632 , 2_n1639 , 2_n1645 , 2_n1687 , 2_n1729 , 2_n1738 , 2_n1752 ;
    wire 2_n0 , 2_n1 , 2_n2 , 2_n3 , 2_n4 , 2_n5 , 2_n6 , 2_n7 , 2_n8 , 2_n9 , 2_n10 , 2_n12 , 2_n13 , 2_n14 , 2_n15 , 2_n16 , 2_n17 , 2_n18 , 2_n19 , 2_n20 , 2_n24 , 2_n25 , 2_n26 , 2_n28 , 2_n31 , 2_n32 , 2_n33 , 2_n34 , 2_n35 , 2_n36 , 2_n37 , 2_n38 , 2_n39 , 2_n41 , 2_n42 , 2_n43 , 2_n44 , 2_n46 , 2_n47 , 2_n48 , 2_n49 , 2_n51 , 2_n53 , 2_n55 , 2_n57 , 2_n59 , 2_n60 , 2_n61 , 2_n62 , 2_n63 , 2_n64 , 2_n65 , 2_n66 , 2_n67 , 2_n68 , 2_n69 , 2_n70 , 2_n72 , 2_n73 , 2_n74 , 2_n75 , 2_n76 , 2_n78 , 2_n79 , 2_n80 , 2_n81 , 2_n83 , 2_n84 , 2_n88 , 2_n89 , 2_n90 , 2_n91 , 2_n92 , 2_n93 , 2_n95 , 2_n96 , 2_n97 , 2_n98 , 2_n99 , 2_n100 , 2_n101 , 2_n102 , 2_n103 , 2_n104 , 2_n105 , 2_n106 , 2_n108 , 2_n109 , 2_n110 , 2_n111 , 2_n113 , 2_n114 , 2_n115 , 2_n116 , 2_n118 , 2_n119 , 2_n120 , 2_n121 , 2_n122 , 2_n123 , 2_n124 , 2_n125 , 2_n127 , 2_n128 , 2_n129 , 2_n131 , 2_n132 , 2_n133 , 2_n134 , 2_n135 , 2_n136 , 2_n137 , 2_n139 , 2_n140 , 2_n141 , 2_n142 , 2_n144 , 2_n145 , 2_n146 , 2_n147 , 2_n148 , 2_n149 , 2_n150 , 2_n151 , 2_n152 , 2_n154 , 2_n157 , 2_n158 , 2_n160 , 2_n162 , 2_n163 , 2_n165 , 2_n166 , 2_n167 , 2_n168 , 2_n169 , 2_n170 , 2_n171 , 2_n172 , 2_n174 , 2_n175 , 2_n176 , 2_n177 , 2_n178 , 2_n179 , 2_n180 , 2_n182 , 2_n183 , 2_n185 , 2_n186 , 2_n187 , 2_n188 , 2_n189 , 2_n190 , 2_n191 , 2_n192 , 2_n193 , 2_n194 , 2_n195 , 2_n196 , 2_n197 , 2_n198 , 2_n199 , 2_n201 , 2_n202 , 2_n203 , 2_n204 , 2_n205 , 2_n206 , 2_n207 , 2_n208 , 2_n209 , 2_n210 , 2_n211 , 2_n212 , 2_n213 , 2_n214 , 2_n215 , 2_n217 , 2_n218 , 2_n221 , 2_n224 , 2_n225 , 2_n226 , 2_n227 , 2_n228 , 2_n229 , 2_n231 , 2_n232 , 2_n234 , 2_n235 , 2_n236 , 2_n237 , 2_n238 , 2_n239 , 2_n240 , 2_n241 , 2_n242 , 2_n245 , 2_n248 , 2_n249 , 2_n250 , 2_n252 , 2_n253 , 2_n255 , 2_n256 , 2_n257 , 2_n258 , 2_n259 , 2_n260 , 2_n261 , 2_n263 , 2_n264 , 2_n265 , 2_n266 , 2_n267 , 2_n269 , 2_n270 , 2_n271 , 2_n272 , 2_n274 , 2_n276 , 2_n277 , 2_n278 , 2_n279 , 2_n280 , 2_n281 , 2_n282 , 2_n283 , 2_n285 , 2_n286 , 2_n287 , 2_n289 , 2_n290 , 2_n291 , 2_n294 , 2_n295 , 2_n296 , 2_n297 , 2_n298 , 2_n302 , 2_n303 , 2_n305 , 2_n306 , 2_n308 , 2_n309 , 2_n311 , 2_n313 , 2_n316 , 2_n317 , 2_n319 , 2_n320 , 2_n321 , 2_n322 , 2_n323 , 2_n324 , 2_n325 , 2_n326 , 2_n327 , 2_n328 , 2_n329 , 2_n330 , 2_n331 , 2_n332 , 2_n333 , 2_n334 , 2_n335 , 2_n336 , 2_n338 , 2_n339 , 2_n340 , 2_n342 , 2_n343 , 2_n345 , 2_n347 , 2_n348 , 2_n349 , 2_n350 , 2_n351 , 2_n353 , 2_n354 , 2_n355 , 2_n356 , 2_n357 , 2_n358 , 2_n359 , 2_n360 , 2_n361 , 2_n363 , 2_n365 , 2_n366 , 2_n367 , 2_n368 , 2_n369 , 2_n371 , 2_n372 , 2_n373 , 2_n375 , 2_n377 , 2_n379 , 2_n381 , 2_n382 , 2_n383 , 2_n384 , 2_n385 , 2_n386 , 2_n387 , 2_n388 , 2_n389 , 2_n390 , 2_n393 , 2_n394 , 2_n395 , 2_n397 , 2_n398 , 2_n400 , 2_n401 , 2_n402 , 2_n403 , 2_n404 , 2_n405 , 2_n406 , 2_n407 , 2_n410 , 2_n411 , 2_n412 , 2_n413 , 2_n414 , 2_n415 , 2_n418 , 2_n419 , 2_n421 , 2_n422 , 2_n423 , 2_n424 , 2_n425 , 2_n426 , 2_n427 , 2_n429 , 2_n431 , 2_n432 , 2_n433 , 2_n434 , 2_n435 , 2_n436 , 2_n437 , 2_n438 , 2_n439 , 2_n440 , 2_n441 , 2_n442 , 2_n443 , 2_n444 , 2_n445 , 2_n446 , 2_n447 , 2_n448 , 2_n449 , 2_n450 , 2_n451 , 2_n452 , 2_n454 , 2_n455 , 2_n456 , 2_n458 , 2_n459 , 2_n461 , 2_n462 , 2_n463 , 2_n464 , 2_n465 , 2_n466 , 2_n467 , 2_n468 , 2_n469 , 2_n470 , 2_n471 , 2_n472 , 2_n473 , 2_n474 , 2_n475 , 2_n476 , 2_n479 , 2_n480 , 2_n481 , 2_n482 , 2_n483 , 2_n484 , 2_n485 , 2_n486 , 2_n488 , 2_n490 , 2_n491 , 2_n492 , 2_n493 , 2_n494 , 2_n495 , 2_n496 , 2_n499 , 2_n500 , 2_n503 , 2_n504 , 2_n505 , 2_n508 , 2_n511 , 2_n512 , 2_n513 , 2_n514 , 2_n515 , 2_n518 , 2_n519 , 2_n520 , 2_n521 , 2_n522 , 2_n523 , 2_n524 , 2_n525 , 2_n526 , 2_n527 , 2_n528 , 2_n529 , 2_n530 , 2_n531 , 2_n532 , 2_n533 , 2_n535 , 2_n536 , 2_n537 , 2_n538 , 2_n539 , 2_n540 , 2_n541 , 2_n542 , 2_n543 , 2_n544 , 2_n546 , 2_n547 , 2_n548 , 2_n549 , 2_n550 , 2_n551 , 2_n552 , 2_n554 , 2_n555 , 2_n556 , 2_n557 , 2_n558 , 2_n562 , 2_n563 , 2_n564 , 2_n565 , 2_n566 , 2_n568 , 2_n569 , 2_n570 , 2_n571 , 2_n572 , 2_n573 , 2_n575 , 2_n576 , 2_n577 , 2_n578 , 2_n579 , 2_n580 , 2_n583 , 2_n584 , 2_n586 , 2_n587 , 2_n588 , 2_n590 , 2_n591 , 2_n592 , 2_n594 , 2_n596 , 2_n599 , 2_n601 , 2_n602 , 2_n603 , 2_n604 , 2_n605 , 2_n606 , 2_n610 , 2_n611 , 2_n612 , 2_n613 , 2_n614 , 2_n615 , 2_n616 , 2_n617 , 2_n618 , 2_n619 , 2_n620 , 2_n621 , 2_n622 , 2_n623 , 2_n624 , 2_n627 , 2_n628 , 2_n629 , 2_n630 , 2_n631 , 2_n632 , 2_n633 , 2_n634 , 2_n635 , 2_n636 , 2_n637 , 2_n639 , 2_n642 , 2_n643 , 2_n644 , 2_n646 , 2_n647 , 2_n648 , 2_n649 , 2_n650 , 2_n651 , 2_n652 , 2_n653 , 2_n654 , 2_n655 , 2_n656 , 2_n657 , 2_n658 , 2_n659 , 2_n660 , 2_n661 , 2_n662 , 2_n664 , 2_n665 , 2_n666 , 2_n667 , 2_n668 , 2_n670 , 2_n672 , 2_n673 , 2_n674 , 2_n675 , 2_n677 , 2_n678 , 2_n679 , 2_n680 , 2_n681 , 2_n682 , 2_n683 , 2_n684 , 2_n685 , 2_n686 , 2_n687 , 2_n688 , 2_n689 , 2_n691 , 2_n692 , 2_n694 , 2_n696 , 2_n697 , 2_n698 , 2_n699 , 2_n700 , 2_n702 , 2_n703 , 2_n704 , 2_n705 , 2_n706 , 2_n707 , 2_n708 , 2_n709 , 2_n711 , 2_n712 , 2_n713 , 2_n715 , 2_n716 , 2_n717 , 2_n718 , 2_n720 , 2_n721 , 2_n722 , 2_n723 , 2_n724 , 2_n725 , 2_n728 , 2_n730 , 2_n731 , 2_n732 , 2_n733 , 2_n735 , 2_n736 , 2_n737 , 2_n738 , 2_n739 , 2_n740 , 2_n741 , 2_n744 , 2_n745 , 2_n746 , 2_n747 , 2_n748 , 2_n749 , 2_n750 , 2_n751 , 2_n752 , 2_n753 , 2_n754 , 2_n756 , 2_n757 , 2_n758 , 2_n759 , 2_n760 , 2_n761 , 2_n762 , 2_n763 , 2_n764 , 2_n765 , 2_n766 , 2_n767 , 2_n768 , 2_n770 , 2_n771 , 2_n772 , 2_n774 , 2_n776 , 2_n777 , 2_n780 , 2_n781 , 2_n783 , 2_n784 , 2_n785 , 2_n786 , 2_n788 , 2_n789 , 2_n791 , 2_n792 , 2_n793 , 2_n795 , 2_n796 , 2_n797 , 2_n798 , 2_n799 , 2_n800 , 2_n801 , 2_n802 , 2_n803 , 2_n804 , 2_n805 , 2_n806 , 2_n807 , 2_n808 , 2_n809 , 2_n810 , 2_n811 , 2_n812 , 2_n813 , 2_n814 , 2_n815 , 2_n816 , 2_n817 , 2_n818 , 2_n819 , 2_n820 , 2_n822 , 2_n824 , 2_n825 , 2_n826 , 2_n827 , 2_n828 , 2_n829 , 2_n830 , 2_n833 , 2_n834 , 2_n835 , 2_n836 , 2_n837 , 2_n838 , 2_n840 , 2_n841 , 2_n843 , 2_n844 , 2_n845 , 2_n846 , 2_n847 , 2_n848 , 2_n850 , 2_n851 , 2_n852 , 2_n853 , 2_n854 , 2_n855 , 2_n856 , 2_n857 , 2_n858 , 2_n859 , 2_n860 , 2_n861 , 2_n862 , 2_n863 , 2_n864 , 2_n865 , 2_n866 , 2_n867 , 2_n868 , 2_n869 , 2_n870 , 2_n871 , 2_n872 , 2_n873 , 2_n874 , 2_n875 , 2_n876 , 2_n877 , 2_n878 , 2_n880 , 2_n881 , 2_n883 , 2_n884 , 2_n886 , 2_n887 , 2_n888 , 2_n889 , 2_n890 , 2_n891 , 2_n892 , 2_n893 , 2_n895 , 2_n896 , 2_n897 , 2_n898 , 2_n899 , 2_n900 , 2_n901 , 2_n902 , 2_n903 , 2_n904 , 2_n906 , 2_n907 , 2_n908 , 2_n909 , 2_n910 , 2_n911 , 2_n912 , 2_n913 , 2_n914 , 2_n915 , 2_n917 , 2_n919 , 2_n921 , 2_n922 , 2_n923 , 2_n924 , 2_n925 , 2_n926 , 2_n927 , 2_n928 , 2_n929 , 2_n930 , 2_n931 , 2_n932 , 2_n933 , 2_n934 , 2_n935 , 2_n937 , 2_n938 , 2_n939 , 2_n940 , 2_n941 , 2_n942 , 2_n943 , 2_n944 , 2_n945 , 2_n946 , 2_n948 , 2_n949 , 2_n950 , 2_n951 , 2_n954 , 2_n955 , 2_n956 , 2_n957 , 2_n958 , 2_n959 , 2_n960 , 2_n962 , 2_n963 , 2_n964 , 2_n965 , 2_n966 , 2_n967 , 2_n968 , 2_n970 , 2_n971 , 2_n972 , 2_n973 , 2_n974 , 2_n975 , 2_n976 , 2_n977 , 2_n978 , 2_n979 , 2_n981 , 2_n982 , 2_n983 , 2_n985 , 2_n987 , 2_n988 , 2_n989 , 2_n991 , 2_n993 , 2_n994 , 2_n995 , 2_n996 , 2_n998 , 2_n999 , 2_n1000 , 2_n1001 , 2_n1002 , 2_n1003 , 2_n1004 , 2_n1005 , 2_n1007 , 2_n1008 , 2_n1009 , 2_n1010 , 2_n1011 , 2_n1012 , 2_n1013 , 2_n1014 , 2_n1015 , 2_n1016 , 2_n1018 , 2_n1019 , 2_n1020 , 2_n1021 , 2_n1022 , 2_n1024 , 2_n1025 , 2_n1026 , 2_n1027 , 2_n1028 , 2_n1029 , 2_n1030 , 2_n1031 , 2_n1032 , 2_n1033 , 2_n1034 , 2_n1035 , 2_n1036 , 2_n1037 , 2_n1038 , 2_n1039 , 2_n1041 , 2_n1043 , 2_n1045 , 2_n1046 , 2_n1047 , 2_n1048 , 2_n1049 , 2_n1052 , 2_n1053 , 2_n1055 , 2_n1056 , 2_n1057 , 2_n1059 , 2_n1062 , 2_n1064 , 2_n1066 , 2_n1067 , 2_n1068 , 2_n1069 , 2_n1070 , 2_n1072 , 2_n1073 , 2_n1074 , 2_n1075 , 2_n1076 , 2_n1077 , 2_n1078 , 2_n1079 , 2_n1080 , 2_n1081 , 2_n1082 , 2_n1083 , 2_n1084 , 2_n1085 , 2_n1086 , 2_n1087 , 2_n1088 , 2_n1089 , 2_n1090 , 2_n1091 , 2_n1092 , 2_n1093 , 2_n1094 , 2_n1096 , 2_n1097 , 2_n1098 , 2_n1099 , 2_n1100 , 2_n1101 , 2_n1102 , 2_n1104 , 2_n1105 , 2_n1106 , 2_n1107 , 2_n1108 , 2_n1109 , 2_n1110 , 2_n1111 , 2_n1112 , 2_n1113 , 2_n1115 , 2_n1116 , 2_n1117 , 2_n1118 , 2_n1119 , 2_n1120 , 2_n1122 , 2_n1123 , 2_n1124 , 2_n1125 , 2_n1126 , 2_n1127 , 2_n1128 , 2_n1129 , 2_n1130 , 2_n1131 , 2_n1132 , 2_n1133 , 2_n1134 , 2_n1135 , 2_n1136 , 2_n1137 , 2_n1139 , 2_n1140 , 2_n1141 , 2_n1142 , 2_n1143 , 2_n1144 , 2_n1145 , 2_n1146 , 2_n1147 , 2_n1148 , 2_n1149 , 2_n1150 , 2_n1151 , 2_n1153 , 2_n1155 , 2_n1157 , 2_n1158 , 2_n1159 , 2_n1160 , 2_n1161 , 2_n1162 , 2_n1163 , 2_n1165 , 2_n1166 , 2_n1167 , 2_n1168 , 2_n1169 , 2_n1170 , 2_n1171 , 2_n1173 , 2_n1174 , 2_n1176 , 2_n1178 , 2_n1179 , 2_n1180 , 2_n1181 , 2_n1182 , 2_n1183 , 2_n1184 , 2_n1185 , 2_n1188 , 2_n1189 , 2_n1190 , 2_n1192 , 2_n1194 , 2_n1196 , 2_n1197 , 2_n1198 , 2_n1199 , 2_n1200 , 2_n1201 , 2_n1202 , 2_n1203 , 2_n1204 , 2_n1206 , 2_n1207 , 2_n1208 , 2_n1210 , 2_n1212 , 2_n1213 , 2_n1214 , 2_n1215 , 2_n1216 , 2_n1217 , 2_n1218 , 2_n1219 , 2_n1220 , 2_n1221 , 2_n1222 , 2_n1223 , 2_n1224 , 2_n1226 , 2_n1228 , 2_n1229 , 2_n1230 , 2_n1232 , 2_n1233 , 2_n1235 , 2_n1236 , 2_n1237 , 2_n1238 , 2_n1240 , 2_n1241 , 2_n1242 , 2_n1243 , 2_n1244 , 2_n1245 , 2_n1247 , 2_n1248 , 2_n1249 , 2_n1251 , 2_n1252 , 2_n1254 , 2_n1255 , 2_n1256 , 2_n1257 , 2_n1258 , 2_n1259 , 2_n1260 , 2_n1261 , 2_n1262 , 2_n1264 , 2_n1265 , 2_n1266 , 2_n1267 , 2_n1268 , 2_n1269 , 2_n1270 , 2_n1271 , 2_n1272 , 2_n1273 , 2_n1274 , 2_n1275 , 2_n1276 , 2_n1277 , 2_n1279 , 2_n1280 , 2_n1282 , 2_n1284 , 2_n1287 , 2_n1290 , 2_n1291 , 2_n1293 , 2_n1294 , 2_n1295 , 2_n1297 , 2_n1298 , 2_n1300 , 2_n1303 , 2_n1304 , 2_n1307 , 2_n1308 , 2_n1309 , 2_n1310 , 2_n1311 , 2_n1312 , 2_n1313 , 2_n1314 , 2_n1315 , 2_n1316 , 2_n1317 , 2_n1318 , 2_n1319 , 2_n1321 , 2_n1323 , 2_n1324 , 2_n1325 , 2_n1326 , 2_n1327 , 2_n1328 , 2_n1329 , 2_n1330 , 2_n1331 , 2_n1332 , 2_n1333 , 2_n1334 , 2_n1335 , 2_n1336 , 2_n1338 , 2_n1339 , 2_n1340 , 2_n1341 , 2_n1342 , 2_n1343 , 2_n1344 , 2_n1347 , 2_n1348 , 2_n1349 , 2_n1351 , 2_n1352 , 2_n1353 , 2_n1354 , 2_n1355 , 2_n1356 , 2_n1357 , 2_n1358 , 2_n1360 , 2_n1362 , 2_n1363 , 2_n1364 , 2_n1365 , 2_n1366 , 2_n1367 , 2_n1369 , 2_n1370 , 2_n1371 , 2_n1372 , 2_n1373 , 2_n1374 , 2_n1376 , 2_n1377 , 2_n1378 , 2_n1379 , 2_n1380 , 2_n1381 , 2_n1382 , 2_n1383 , 2_n1384 , 2_n1385 , 2_n1388 , 2_n1390 , 2_n1392 , 2_n1394 , 2_n1395 , 2_n1396 , 2_n1397 , 2_n1398 , 2_n1399 , 2_n1400 , 2_n1402 , 2_n1403 , 2_n1404 , 2_n1405 , 2_n1406 , 2_n1407 , 2_n1408 , 2_n1409 , 2_n1410 , 2_n1412 , 2_n1413 , 2_n1414 , 2_n1416 , 2_n1417 , 2_n1419 , 2_n1422 , 2_n1423 , 2_n1424 , 2_n1425 , 2_n1426 , 2_n1429 , 2_n1430 , 2_n1431 , 2_n1432 , 2_n1433 , 2_n1434 , 2_n1436 , 2_n1437 , 2_n1439 , 2_n1440 , 2_n1441 , 2_n1442 , 2_n1444 , 2_n1445 , 2_n1447 , 2_n1449 , 2_n1450 , 2_n1451 , 2_n1452 , 2_n1453 , 2_n1454 , 2_n1455 , 2_n1456 , 2_n1457 , 2_n1458 , 2_n1459 , 2_n1460 , 2_n1461 , 2_n1462 , 2_n1464 , 2_n1465 , 2_n1466 , 2_n1467 , 2_n1468 , 2_n1469 , 2_n1471 , 2_n1472 , 2_n1473 , 2_n1475 , 2_n1477 , 2_n1478 , 2_n1479 , 2_n1480 , 2_n1481 , 2_n1482 , 2_n1483 , 2_n1484 , 2_n1485 , 2_n1486 , 2_n1487 , 2_n1488 , 2_n1489 , 2_n1490 , 2_n1491 , 2_n1492 , 2_n1493 , 2_n1494 , 2_n1495 , 2_n1496 , 2_n1497 , 2_n1498 , 2_n1499 , 2_n1501 , 2_n1503 , 2_n1504 , 2_n1505 , 2_n1507 , 2_n1508 , 2_n1509 , 2_n1510 , 2_n1511 , 2_n1512 , 2_n1513 , 2_n1514 , 2_n1515 , 2_n1517 , 2_n1518 , 2_n1519 , 2_n1522 , 2_n1524 , 2_n1525 , 2_n1526 , 2_n1528 , 2_n1529 , 2_n1530 , 2_n1531 , 2_n1532 , 2_n1533 , 2_n1535 , 2_n1537 , 2_n1538 , 2_n1539 , 2_n1540 , 2_n1541 , 2_n1542 , 2_n1543 , 2_n1544 , 2_n1545 , 2_n1546 , 2_n1549 , 2_n1550 , 2_n1551 , 2_n1552 , 2_n1553 , 2_n1554 , 2_n1555 , 2_n1556 , 2_n1557 , 2_n1558 , 2_n1559 , 2_n1560 , 2_n1561 , 2_n1562 , 2_n1563 , 2_n1564 , 2_n1565 , 2_n1567 , 2_n1568 , 2_n1570 , 2_n1571 , 2_n1572 , 2_n1573 , 2_n1574 , 2_n1575 , 2_n1577 , 2_n1578 , 2_n1579 , 2_n1580 , 2_n1581 , 2_n1582 , 2_n1583 , 2_n1584 , 2_n1585 , 2_n1587 , 2_n1589 , 2_n1590 , 2_n1591 , 2_n1593 , 2_n1595 , 2_n1596 , 2_n1597 , 2_n1598 , 2_n1599 , 2_n1600 , 2_n1601 , 2_n1602 , 2_n1603 , 2_n1604 , 2_n1605 , 2_n1606 , 2_n1607 , 2_n1608 , 2_n1610 , 2_n1611 , 2_n1612 , 2_n1614 , 2_n1615 , 2_n1617 , 2_n1618 , 2_n1619 , 2_n1620 , 2_n1621 , 2_n1622 , 2_n1623 , 2_n1624 , 2_n1625 , 2_n1628 , 2_n1629 , 2_n1630 , 2_n1631 , 2_n1633 , 2_n1634 , 2_n1635 , 2_n1636 , 2_n1637 , 2_n1638 , 2_n1640 , 2_n1641 , 2_n1642 , 2_n1643 , 2_n1646 , 2_n1648 , 2_n1649 , 2_n1650 , 2_n1651 , 2_n1652 , 2_n1653 , 2_n1654 , 2_n1655 , 2_n1657 , 2_n1658 , 2_n1659 , 2_n1660 , 2_n1661 , 2_n1662 , 2_n1663 , 2_n1664 , 2_n1665 , 2_n1666 , 2_n1667 , 2_n1668 , 2_n1669 , 2_n1670 , 2_n1671 , 2_n1672 , 2_n1673 , 2_n1674 , 2_n1675 , 2_n1676 , 2_n1677 , 2_n1678 , 2_n1679 , 2_n1680 , 2_n1681 , 2_n1682 , 2_n1683 , 2_n1684 , 2_n1685 , 2_n1686 , 2_n1688 , 2_n1689 , 2_n1690 , 2_n1691 , 2_n1692 , 2_n1693 , 2_n1694 , 2_n1695 , 2_n1696 , 2_n1697 , 2_n1698 , 2_n1699 , 2_n1700 , 2_n1701 , 2_n1702 , 2_n1703 , 2_n1704 , 2_n1705 , 2_n1706 , 2_n1707 , 2_n1708 , 2_n1709 , 2_n1710 , 2_n1711 , 2_n1712 , 2_n1713 , 2_n1714 , 2_n1715 , 2_n1716 , 2_n1717 , 2_n1718 , 2_n1719 , 2_n1720 , 2_n1721 , 2_n1722 , 2_n1723 , 2_n1724 , 2_n1725 , 2_n1726 , 2_n1727 , 2_n1728 , 2_n1730 , 2_n1731 , 2_n1732 , 2_n1733 , 2_n1734 , 2_n1735 , 2_n1736 , 2_n1737 , 2_n1739 , 2_n1740 , 2_n1741 , 2_n1742 , 2_n1743 , 2_n1744 , 2_n1745 , 2_n1746 , 2_n1747 , 2_n1748 , 2_n1749 , 2_n1751 , 2_n1754 , 2_n1755 , 2_n1756 ;
assign 2_n426 = 2_n422 | 2_n1543;
assign 2_n1664 = 2_n889 | 2_n1101;
assign 2_n1637 = ~(2_n456 ^ 2_n1142);
assign 2_n1067 = ~(2_n1402 ^ 2_n145);
assign 2_n993 = ~(2_n780 ^ 2_n1263);
assign 2_n1517 = 2_n206 ^ 2_n1725;
assign 2_n1735 = 2_n1116 | 2_n1429;
assign 2_n1539 = 2_n1683 & 2_n1276;
assign 2_n154 = ~2_n1002;
assign 2_n1347 = ~(2_n142 | 2_n1105);
assign 2_n1537 = ~2_n1540;
assign 2_n1608 = ~(2_n1573 ^ 2_n866);
assign 2_n960 = ~2_n1377;
assign 2_n476 = 2_n768 & 2_n1126;
assign 2_n805 = 2_n1485 | 2_n192;
assign 2_n752 = ~(2_n88 ^ 2_n540);
assign 2_n1048 = ~2_n654;
assign 2_n1698 = ~(2_n1343 | 2_n109);
assign 2_n1326 = ~(2_n289 | 2_n1230);
assign 2_n721 = ~2_n728;
assign 2_n1555 = ~2_n886;
assign 2_n1578 = 2_n1194 | 2_n25;
assign 2_n1383 = 2_n802 | 2_n218;
assign 2_n821 = 2_n374;
assign 2_n802 = ~2_n837;
assign 2_n103 = 2_n1706 | 2_n1557;
assign 2_n175 = 2_n717 | 2_n943;
assign 2_n468 = ~2_n1419;
assign 2_n38 = ~(2_n1207 ^ 2_n557);
assign 2_n1585 = 2_n1115 | 2_n238;
assign 2_n1105 = 2_n1416 | 2_n467;
assign 2_n1648 = 2_n935 | 2_n266;
assign 2_n165 = ~2_n1664;
assign 2_n212 = 2_n1721 | 2_n500;
assign 2_n624 = 2_n885 & 2_n197;
assign 2_n1218 = 2_n986 & 2_n0;
assign 2_n1002 = 2_n228 | 2_n1551;
assign 2_n256 = 2_n1357 | 2_n1533;
assign 2_n102 = 2_n1531 | 2_n686;
assign 2_n1617 = ~(2_n1373 ^ 2_n1417);
assign 2_n123 = ~(2_n1512 ^ 2_n1355);
assign 2_n272 = 2_n1100 & 2_n177;
assign 2_n305 = 2_n1481 | 2_n272;
assign 2_n104 = ~(2_n721 | 2_n1401);
assign 2_n973 = 2_n1408 | 2_n379;
assign 2_n70 = ~2_n923;
assign 2_n1365 = ~2_n1506;
assign 2_n1316 = ~(2_n632 ^ 2_n1595);
assign 2_n1015 = 2_n376 & 2_n1168;
assign 2_n1302 = ~(2_n837 ^ 2_n933);
assign 2_n1480 = 2_n779 & 2_n721;
assign 2_n1719 = 2_n251 & 2_n1555;
assign 2_n1188 = 2_n1268 | 2_n1458;
assign 2_n148 = ~(2_n721 | 2_n1138);
assign 2_n436 = ~(2_n777 ^ 2_n194);
assign 2_n1247 = ~(2_n1037 ^ 2_n72);
assign 2_n747 = ~2_n1708;
assign 2_n579 = ~2_n1293;
assign 2_n1556 = ~(2_n723 ^ 2_n518);
assign 2_n471 = 2_n1558 & 2_n1312;
assign 2_n327 = ~2_n843;
assign 2_n846 = ~2_n324;
assign 2_n1488 = ~(2_n623 ^ 2_n1382);
assign 2_n1237 = ~(2_n380 & 2_n701);
assign 2_n785 = 2_n63 & 2_n807;
assign 2_n1370 = 2_n559 & 2_n491;
assign 2_n388 = ~2_n1559;
assign 2_n658 = 2_n1696 | 2_n835;
assign 2_n914 = ~2_n1387;
assign 2_n331 = ~(2_n1107 ^ 2_n1707);
assign 2_n1212 = ~(2_n999 ^ 2_n24);
assign 2_n1623 = ~2_n891;
assign 2_n488 = ~(2_n1535 | 2_n1628);
assign 2_n681 = 2_n1172 & 2_n602;
assign 2_n1017 = 2_n1476;
assign 2_n298 = ~2_n1521;
assign 2_n923 = 2_n1692 & 2_n474;
assign 2_n670 = ~2_n626;
assign 2_n554 = 2_n134 & 2_n1400;
assign 2_n1515 = ~2_n1008;
assign 2_n1325 = 2_n1579 | 2_n423;
assign 2_n1201 = 2_n1623 | 2_n1511;
assign 2_n549 = ~(2_n63 | 2_n32);
assign 2_n1158 = 2_n1241 | 2_n1354;
assign 2_n197 = ~2_n1314;
assign 2_n861 = 2_n64 | 2_n1244;
assign 2_n801 = ~(2_n1615 | 2_n1336);
assign 2_n151 = 2_n312 & 2_n1458;
assign 2_n516 = 2_n1187;
assign 2_n1075 = 2_n124 & 2_n1482;
assign 2_n946 = 2_n568 | 2_n999;
assign 2_n1525 = ~(2_n1339 ^ 2_n615);
assign 2_n587 = ~(2_n1734 | 2_n772);
assign 2_n1179 = ~2_n545;
assign 2_n686 = ~(2_n1178 | 2_n175);
assign 2_n1465 = 2_n1254 | 2_n1167;
assign 2_n1477 = 2_n89 & 2_n495;
assign 2_n1687 = 2_n523 | 2_n73;
assign 2_n1538 = 2_n1013 | 2_n444;
assign 2_n1355 = ~2_n188;
assign 2_n1736 = 2_n687 | 2_n979;
assign 2_n1119 = ~(2_n257 | 2_n200);
assign 2_n26 = ~2_n778;
assign 2_n1714 = ~(2_n1445 ^ 2_n1084);
assign 2_n1658 = 2_n1261 | 2_n10;
assign 2_n1596 = 2_n1393 & 2_n530;
assign 2_n1673 = ~2_n993;
assign 2_n1743 = 2_n359 | 2_n434;
assign 2_n1335 = ~(2_n1686 | 2_n1073);
assign 2_n1612 = ~(2_n721 | 2_n56);
assign 2_n1458 = ~2_n808;
assign 2_n182 = 2_n1346 & 2_n602;
assign 2_n1468 = ~(2_n1597 ^ 2_n980);
assign 2_n195 = 2_n1251 & 2_n1598;
assign 2_n1307 = ~(2_n1273 ^ 2_n427);
assign 2_n324 = ~(2_n1721 ^ 2_n732);
assign 2_n828 = 2_n1752 | 2_n493;
assign 2_n958 = 2_n1673 & 2_n798;
assign 2_n301 = 2_n318;
assign 2_n316 = ~2_n1201;
assign 2_n174 = ~(2_n1597 ^ 2_n923);
assign 2_n119 = ~2_n567;
assign 2_n124 = 2_n395 & 2_n1034;
assign 2_n460 = 2_n21;
assign 2_n1496 = ~(2_n1049 ^ 2_n630);
assign 2_n1214 = ~2_n339;
assign 2_n504 = ~(2_n49 ^ 2_n1406);
assign 2_n1107 = ~(2_n83 ^ 2_n724);
assign 2_n811 = ~2_n1475;
assign 2_n1189 = 2_n2 & 2_n323;
assign 2_n17 = ~2_n865;
assign 2_n474 = 2_n803 | 2_n905;
assign 2_n1084 = ~(2_n1648 ^ 2_n1018);
assign 2_n1287 = ~(2_n261 ^ 2_n1727);
assign 2_n252 = ~(2_n522 | 2_n132);
assign 2_n760 = 2_n1230 & 2_n873;
assign 2_n1497 = 2_n721 | 2_n346;
assign 2_n606 = ~(2_n1537 ^ 2_n60);
assign 2_n481 = 2_n1182 | 2_n1238;
assign 2_n306 = 2_n1577 | 2_n1203;
assign 2_n99 = ~(2_n1535 ^ 2_n1442);
assign 2_n35 = 2_n636 | 2_n1620;
assign 2_n1394 = ~2_n1681;
assign 2_n1099 = 2_n1489 | 2_n806;
assign 2_n1306 = 2_n1204 | 2_n1619;
assign 2_n302 = ~(2_n1173 ^ 2_n608);
assign 2_n1600 = ~(2_n32 ^ 2_n1473);
assign 2_n308 = ~2_n1239;
assign 2_n611 = ~(2_n1166 ^ 2_n1699);
assign 2_n1058 = ~(2_n1667 ^ 2_n810);
assign 2_n687 = ~2_n1711;
assign 2_n1430 = ~2_n307;
assign 2_n414 = ~(2_n1470 | 2_n910);
assign 2_n1511 = ~2_n907;
assign 2_n340 = 2_n613 & 2_n698;
assign 2_n1621 = 2_n934 & 2_n1697;
assign 2_n1532 = ~(2_n1667 | 2_n840);
assign 2_n1404 = 2_n133 ^ 2_n375;
assign 2_n921 = 2_n1644 & 2_n1136;
assign 2_n835 = ~2_n413;
assign 2_n1395 = ~2_n738;
assign 2_n1072 = ~(2_n899 ^ 2_n938);
assign 2_n492 = ~(2_n900 | 2_n86);
assign 2_n637 = 2_n1672 & 2_n1475;
assign 2_n213 = 2_n142 ^ 2_n1083;
assign 2_n1269 = ~(2_n999 | 2_n703);
assign 2_n999 = ~2_n1419;
assign 2_n373 = ~(2_n740 ^ 2_n407);
assign 2_n1170 = 2_n903 | 2_n694;
assign 2_n271 = 2_n1750 & 2_n238;
assign 2_n177 = ~(2_n1230 | 2_n1335);
assign 2_n1689 = ~(2_n1200 ^ 2_n707);
assign 2_n1282 = 2_n454 | 2_n639;
assign 2_n1235 = 2_n1722 | 2_n649;
assign 2_n900 = ~2_n413;
assign 2_n1747 = 2_n1102 | 2_n75;
assign 2_n1148 = 2_n798 | 2_n1390;
assign 2_n96 = 2_n687 | 2_n1139;
assign 2_n140 = 2_n651 & 2_n248;
assign 2_n1194 = ~(2_n1099 | 2_n189);
assign 2_n635 = 2_n1668 | 2_n197;
assign 2_n137 = 2_n1415 & 2_n530;
assign 2_n1018 = 2_n479 & 2_n840;
assign 2_n530 = ~2_n808;
assign 2_n1085 = 2_n899 & 2_n1264;
assign 2_n1162 = 2_n803 | 2_n1191;
assign 2_n357 = ~(2_n367 | 2_n158);
assign 2_n91 = 2_n985 | 2_n443;
assign 2_n1083 = 2_n1015 | 2_n804;
assign 2_n1091 = ~(2_n876 ^ 2_n33);
assign 2_n367 = 2_n1360 & 2_n575;
assign 2_n1274 = 2_n1698 | 2_n1075;
assign 2_n379 = 2_n964 | 2_n717;
assign 2_n1229 = ~(2_n922 ^ 2_n1651);
assign 2_n1126 = ~2_n852;
assign 2_n1197 = ~2_n179;
assign 2_n962 = ~(2_n1686 ^ 2_n1498);
assign 2_n47 = 2_n1083 & 2_n1492;
assign 2_n1113 = ~2_n1188;
assign 2_n1457 = ~(2_n206 ^ 2_n1343);
assign 2_n1155 = 2_n1405 | 2_n567;
assign 2_n866 = ~(2_n654 ^ 2_n1629);
assign 2_n1353 = 2_n204 | 2_n577;
assign 2_n537 = 2_n1291 | 2_n1098;
assign 2_n1618 = 2_n761 | 2_n465;
assign 2_n1397 = 2_n219 & 2_n1168;
assign 2_n758 = ~2_n565;
assign 2_n1582 = ~(2_n1641 ^ 2_n1476);
assign 2_n1272 = ~(2_n146 | 2_n481);
assign 2_n592 = 2_n760 | 2_n1327;
assign 2_n1226 = 2_n1585 & 2_n569;
assign 2_n1642 = 2_n1561 | 2_n250;
assign 2_n1380 = ~(2_n1573 ^ 2_n1133);
assign 2_n1132 = ~(2_n324 | 2_n241);
assign 2_n1135 = ~2_n888;
assign 2_n746 = 2_n1493 | 2_n503;
assign 2_n1320 = 2_n1263;
assign 2_n100 = ~(2_n354 | 2_n1137);
assign 2_n1009 = ~(2_n1340 ^ 2_n1636);
assign 2_n259 = ~2_n908;
assign 2_n719 = 2_n1361 | 2_n1225;
assign 2_n245 = ~(2_n803 | 2_n769);
assign 2_n486 = 2_n614 | 2_n1012;
assign 2_n1604 = ~(2_n572 | 2_n1682);
assign 2_n525 = ~(2_n1673 ^ 2_n1148);
assign 2_n1056 = ~(2_n555 ^ 2_n730);
assign 2_n9 = ~2_n1284;
assign 2_n1738 = 2_n45;
assign 2_n718 = 2_n629 | 2_n636;
assign 2_n266 = 2_n1552 | 2_n1222;
assign 2_n120 = 2_n1288 | 2_n1322;
assign 2_n807 = 2_n1136 | 2_n1435;
assign 2_n1565 = ~2_n1747;
assign 2_n812 = 2_n1623 ^ 2_n907;
assign 2_n874 = ~(2_n1535 | 2_n1695);
assign 2_n1190 = 2_n695 | 2_n653;
assign 2_n646 = ~(2_n852 | 2_n1436);
assign 2_n1133 = 2_n883 | 2_n1048;
assign 2_n229 = 2_n793 | 2_n59;
assign 2_n383 = ~(2_n948 ^ 2_n1148);
assign 2_n1709 = 2_n849 & 2_n776;
assign 2_n1358 = 2_n1700 | 2_n212;
assign 2_n1215 = ~(2_n1601 | 2_n998);
assign 2_n348 = ~2_n1307;
assign 2_n731 = ~2_n1694;
assign 2_n1716 = 2_n1304 | 2_n333;
assign 2_n798 = 2_n249 & 2_n1129;
assign 2_n1381 = ~2_n1043;
assign 2_n1493 = ~2_n225;
assign 2_n180 = ~2_n1386;
assign 2_n1399 = 2_n930 & 2_n655;
assign 2_n1740 = 2_n824 | 2_n618;
assign 2_n777 = 2_n137 | 2_n207;
assign 2_n1315 = 2_n1328 | 2_n900;
assign 2_n1513 = ~(2_n1405 | 2_n823);
assign 2_n199 = 2_n915 | 2_n257;
assign 2_n1267 = 2_n416 & 2_n444;
assign 2_n239 = ~2_n50;
assign 2_n48 = ~(2_n613 ^ 2_n405);
assign 2_n800 = ~(2_n318 | 2_n781);
assign 2_n1033 = 2_n514 | 2_n989;
assign 2_n738 = 2_n682 | 2_n668;
assign 2_n536 = 2_n790 & 2_n240;
assign 2_n551 = ~2_n1007;
assign 2_n93 = ~(2_n899 ^ 2_n960);
assign 2_n639 = 2_n1657 | 2_n403;
assign 2_n1037 = ~(2_n469 ^ 2_n1055);
assign 2_n511 = 2_n637 & 2_n1078;
assign 2_n326 = 2_n1333 | 2_n1150;
assign 2_n1297 = ~2_n1077;
assign 2_n1741 = 2_n1141 | 2_n1731;
assign 2_n80 = ~2_n938;
assign 2_n1243 = 2_n47 | 2_n1022;
assign 2_n1624 = 2_n838 | 2_n983;
assign 2_n240 = ~2_n808;
assign 2_n483 = 2_n238 | 2_n839;
assign 2_n1718 = 2_n5 | 2_n1722;
assign 2_n303 = 2_n691 & 2_n639;
assign 2_n134 = ~2_n1261;
assign 2_n1016 = 2_n755 & 2_n721;
assign 2_n1150 = ~2_n668;
assign 2_n422 = ~(2_n675 ^ 2_n1398);
assign 2_n817 = ~(2_n736 | 2_n1422);
assign 2_n88 = 2_n20 | 2_n864;
assign 2_n1482 = 2_n170 | 2_n1545;
assign 2_n1599 = ~2_n887;
assign 2_n963 = 2_n1461 | 2_n444;
assign 2_n1106 = 2_n119 & 2_n1002;
assign 2_n230 = 2_n831;
assign 2_n1526 = ~(2_n630 | 2_n1355);
assign 2_n1570 = 2_n1673 & 2_n1390;
assign 2_n1661 = ~(2_n99 ^ 2_n129);
assign 2_n242 = ~(2_n1637 ^ 2_n606);
assign 2_n1324 = ~2_n1396;
assign 2_n1043 = 2_n1724 | 2_n386;
assign 2_n509 = 2_n769;
assign 2_n1614 = 2_n1298 | 2_n1394;
assign 2_n249 = ~2_n1116;
assign 2_n1437 = 2_n1542 | 2_n875;
assign 2_n378 = ~(2_n224 ^ 2_n211);
assign 2_n1087 = ~(2_n721 | 2_n1502);
assign 2_n1221 = ~(2_n1438 & 2_n1536);
assign 2_n437 = ~(2_n1220 ^ 2_n394);
assign 2_n1427 = 2_n1407 | 2_n1562;
assign 2_n235 = 2_n1377 | 2_n1756;
assign 2_n570 = ~(2_n708 ^ 2_n948);
assign 2_n1375 = 2_n229 | 2_n770;
assign 2_n1455 = 2_n1004 & 2_n1044;
assign 2_n90 = ~(2_n265 ^ 2_n24);
assign 2_n1486 = ~2_n1635;
assign 2_n227 = 2_n150 | 2_n1290;
assign 2_n1094 = 2_n1319 & 2_n205;
assign 2_n1384 = 2_n309 | 2_n444;
assign 2_n749 = ~2_n419;
assign 2_n1417 = ~(2_n1303 ^ 2_n1641);
assign 2_n883 = ~2_n1629;
assign 2_n1045 = ~(2_n43 ^ 2_n33);
assign 2_n387 = 2_n217 | 2_n877;
assign 2_n820 = ~2_n203;
assign 2_n1314 = ~2_n263;
assign 2_n1144 = ~2_n212;
assign 2_n466 = 2_n441 | 2_n636;
assign 2_n950 = 2_n1692 & 2_n483;
assign 2_n655 = 2_n971 | 2_n530;
assign 2_n112 = ~(2_n42 ^ 2_n907);
assign 2_n794 = ~(2_n225 ^ 2_n1208);
assign 2_n167 = 2_n238 | 2_n222;
assign 2_n1251 = 2_n1293 | 2_n708;
assign 2_n1019 = 2_n651 | 2_n527;
assign 2_n1396 = 2_n100 & 2_n1666;
assign 2_n660 = 2_n676 & 2_n197;
assign 2_n1078 = 2_n248 & 2_n527;
assign 2_n135 = ~2_n1073;
assign 2_n1051 = ~(2_n689 ^ 2_n168);
assign 2_n496 = 2_n564 & 2_n473;
assign 2_n1339 = ~(2_n66 ^ 2_n336);
assign 2_n1629 = 2_n2 | 2_n684;
assign 2_n1177 = 2_n487;
assign 2_n1639 = ~(2_n302 ^ 2_n801);
assign 2_n465 = 2_n1152 & 2_n491;
assign 2_n433 = ~(2_n315 & 2_n997);
assign 2_n677 = 2_n1648 | 2_n1232;
assign 2_n1011 = 2_n1513 | 2_n1426;
assign 2_n740 = 2_n1309 | 2_n1742;
assign 2_n1321 = ~2_n691;
assign 2_n534 = ~(2_n248 ^ 2_n472);
assign 2_n515 = 2_n579 | 2_n706;
assign 2_n386 = ~2_n1174;
assign 2_n1459 = ~(2_n321 ^ 2_n1507);
assign 2_n490 = 2_n1029 | 2_n748;
assign 2_n519 = 2_n1682 & 2_n994;
assign 2_n1060 = 2_n762 | 2_n1702;
assign 2_n850 = ~2_n1061;
assign 2_n803 = ~2_n413;
assign 2_n14 = ~2_n1279;
assign 2_n1151 = 2_n868 | 2_n212;
assign 2_n1501 = 2_n1140 | 2_n148;
assign 2_n429 = ~2_n1629;
assign 2_n1700 = ~2_n1582;
assign 2_n231 = 2_n565 & 2_n1150;
assign 2_n463 = 2_n836 | 2_n240;
assign 2_n32 = 2_n884 | 2_n745;
assign 2_n1527 = ~(2_n311 ^ 2_n1706);
assign 2_n768 = 2_n214 & 2_n981;
assign 2_n1219 = ~2_n561;
assign 2_n406 = 2_n845 | 2_n1070;
assign 2_n662 = 2_n282 | 2_n496;
assign 2_n943 = 2_n1491 | 2_n1722;
assign 2_n1035 = 2_n732 & 2_n340;
assign 2_n451 = 2_n979 | 2_n647;
assign 2_n1454 = ~(2_n1742 | 2_n1035);
assign 2_n1349 = 2_n1630 | 2_n1405;
assign 2_n228 = 2_n268 & 2_n1168;
assign 2_n926 = 2_n1413 | 2_n356;
assign 2_n991 = 2_n1059 & 2_n946;
assign 2_n928 = ~(2_n1089 | 2_n787);
assign 2_n1216 = 2_n1057 | 2_n226;
assign 2_n1597 = 2_n1692 & 2_n1509;
assign 2_n1522 = 2_n1103 & 2_n491;
assign 2_n292 = 2_n408;
assign 2_n1462 = ~(2_n1572 ^ 2_n769);
assign 2_n858 = ~(2_n490 | 2_n1229);
assign 2_n359 = 2_n1216 | 2_n932;
assign 2_n419 = 2_n591 | 2_n530;
assign 2_n221 = ~2_n605;
assign 2_n867 = 2_n1555 & 2_n117;
assign 2_n442 = ~(2_n1515 ^ 2_n1487);
assign 2_n765 = 2_n774 | 2_n982;
assign 2_n533 = 2_n1367 | 2_n149;
assign 2_n1142 = ~(2_n371 ^ 2_n1665);
assign 2_n784 = ~2_n1648;
assign 2_n1020 = 2_n906 & 2_n1371;
assign 2_n1607 = 2_n679 | 2_n389;
assign 2_n41 = 2_n721 | 2_n223;
assign 2_n1117 = ~(2_n408 | 2_n704);
assign 2_n1602 = 2_n63 & 2_n1374;
assign 2_n1007 = 2_n1349 & 2_n1077;
assign 2_n717 = ~(2_n1402 ^ 2_n895);
assign 2_n1086 = 2_n1479 | 2_n738;
assign 2_n1228 = 2_n84 & 2_n777;
assign 2_n289 = 2_n811 | 2_n1432;
assign 2_n1708 = 2_n529 | 2_n1555;
assign 2_n1715 = ~2_n1064;
assign 2_n697 = 2_n1493 | 2_n677;
assign 2_n121 = ~(2_n1623 ^ 2_n739);
assign 2_n1694 = ~(2_n841 ^ 2_n1470);
assign 2_n1080 = ~(2_n994 | 2_n242);
assign 2_n1467 = 2_n1655 | 2_n1119;
assign 2_n69 = 2_n1049 | 2_n368;
assign 2_n1655 = 2_n589 & 2_n835;
assign 2_n989 = ~(2_n1399 | 2_n452);
assign 2_n1734 = ~(2_n1232 ^ 2_n225);
assign 2_n809 = ~(2_n1493 | 2_n435);
assign 2_n588 = ~(2_n18 | 2_n1726);
assign 2_n1076 = ~2_n1250;
assign 2_n1169 = ~(2_n321 ^ 2_n1336);
assign 2_n1357 = ~2_n1432;
assign 2_n1434 = ~(2_n1535 | 2_n659);
assign 2_n653 = 2_n1528 & 2_n1703;
assign 2_n25 = ~(2_n144 | 2_n306);
assign 2_n956 = ~(2_n1364 | 2_n901);
assign 2_n930 = 2_n238 | 2_n1071;
assign 2_n1323 = 2_n40 & 2_n257;
assign 2_n364 = 2_n1477 | 2_n1508;
assign 2_n1407 = 2_n1212 & 2_n1650;
assign 2_n1279 = ~(2_n1530 ^ 2_n138);
assign 2_n183 = ~(2_n741 | 2_n891);
assign 2_n1484 = 2_n467 | 2_n363;
assign 2_n1483 = ~(2_n1159 ^ 2_n610);
assign 2_n682 = 2_n545 & 2_n758;
assign 2_n564 = ~2_n479;
assign 2_n139 = ~2_n78;
assign 2_n187 = ~(2_n38 ^ 2_n1009);
assign 2_n142 = 2_n735 & 2_n887;
assign 2_n772 = ~(2_n859 ^ 2_n825);
assign 2_n661 = ~(2_n803 | 2_n94);
assign 2_n1028 = 2_n921 | 2_n1541;
assign 2_n126 = 2_n1449 | 2_n566;
assign 2_n12 = ~(2_n236 ^ 2_n1496);
assign 2_n869 = 2_n1127 | 2_n197;
assign 2_n1543 = ~(2_n1659 ^ 2_n111);
assign 2_n1332 = 2_n1379 | 2_n578;
assign 2_n1340 = ~(2_n874 ^ 2_n1635);
assign 2_n735 = 2_n524 | 2_n257;
assign 2_n1173 = 2_n1553 | 2_n198;
assign 2_n443 = ~(2_n1575 | 2_n402);
assign 2_n913 = 2_n1106 | 2_n1559;
assign 2_n1727 = 2_n949 ^ 2_n857;
assign 2_n896 = ~2_n1734;
assign 2_n269 = ~2_n750;
assign 2_n253 = ~(2_n1537 | 2_n1307);
assign 2_n1240 = 2_n689 & 2_n576;
assign 2_n1545 = 2_n169 | 2_n1728;
assign 2_n1196 = 2_n1021 ^ 2_n1301;
assign 2_n659 = ~(2_n1405 | 2_n1389);
assign 2_n484 = ~2_n1202;
assign 2_n250 = 2_n1193 & 2_n491;
assign 2_n427 = ~(2_n470 ^ 2_n157);
assign 2_n819 = 2_n159 & 2_n835;
assign 2_n390 = ~(2_n1026 | 2_n340);
assign 2_n190 = ~2_n1627;
assign 2_n1253 = 2_n1050;
assign 2_n369 = ~(2_n66 ^ 2_n172);
assign 2_n1293 = 2_n980 | 2_n358;
assign 2_n1166 = ~(2_n1249 ^ 2_n957);
assign 2_n683 = 2_n1126 & 2_n1204;
assign 2_n333 = 2_n1121 & 2_n491;
assign 2_n89 = ~(2_n249 ^ 2_n327);
assign 2_n1184 = 2_n1672 & 2_n1634;
assign 2_n448 = 2_n98 | 2_n1383;
assign 2_n505 = 2_n976 | 2_n1705;
assign 2_n774 = ~(2_n205 | 2_n1390);
assign 2_n542 = ~(2_n654 ^ 2_n1380);
assign 2_n754 = ~(2_n752 ^ 2_n851);
assign 2_n602 = ~2_n413;
assign 2_n1590 = 2_n1483 | 2_n1030;
assign 2_n461 = ~2_n302;
assign 2_n753 = ~(2_n543 ^ 2_n1716);
assign 2_n1414 = 2_n446 & 2_n476;
assign 2_n0 = 2_n627 | 2_n1341;
assign 2_n750 = 2_n1210 | 2_n747;
assign 2_n1273 = ~(2_n1604 ^ 2_n505);
assign 2_n1392 = 2_n1275 | 2_n1046;
assign 2_n1128 = ~(2_n896 | 2_n783);
assign 2_n211 = 2_n1080 | 2_n1621;
assign 2_n815 = 2_n1649 | 2_n1088;
assign 2_n1693 = ~(2_n1217 | 2_n911);
assign 2_n1571 = 2_n879 & 2_n900;
assign 2_n573 = 2_n1007 | 2_n145;
assign 2_n1717 = 2_n1200 & 2_n1664;
assign 2_n1079 = ~2_n538;
assign 2_n906 = ~2_n1733;
assign 2_n181 = ~(2_n1468 ^ 2_n1505);
assign 2_n804 = 2_n262 & 2_n602;
assign 2_n42 = ~2_n1743;
assign 2_n512 = 2_n369 | 2_n1271;
assign 2_n20 = 2_n1419 & 2_n237;
assign 2_n1490 = 2_n1518 | 2_n1053;
assign 2_n1171 = ~(2_n1260 ^ 2_n1725);
assign 2_n1070 = 2_n409 & 2_n1136;
assign 2_n557 = ~(2_n1530 ^ 2_n841);
assign 2_n698 = 2_n1324 | 2_n61;
assign 2_n377 = 2_n1414 | 2_n583;
assign 2_n1507 = ~(2_n302 ^ 2_n473);
assign 2_n1622 = ~2_n941;
assign 2_n1460 = ~(2_n811 | 2_n1079);
assign 2_n23 = 2_n346;
assign 2_n863 = 2_n835 | 2_n1500;
assign 2_n957 = 2_n653 ^ 2_n972;
assign 2_n97 = 2_n1189 | 2_n449;
assign 2_n1534 = 2_n920;
assign 2_n616 = 2_n687 | 2_n979;
assign 2_n418 = ~(2_n471 ^ 2_n332);
assign 2_n893 = ~(2_n1700 ^ 2_n339);
assign 2_n1676 = 2_n1660 | 2_n681;
assign 2_n1568 = ~2_n1476;
assign 2_n1050 = 2_n1361 | 2_n1237;
assign 2_n771 = 2_n1144 | 2_n1579;
assign 2_n651 = 2_n287 & 2_n1382;
assign 2_n1352 = ~2_n972;
assign 2_n129 = ~(2_n1434 ^ 2_n488);
assign 2_n432 = ~(2_n1135 | 2_n265);
assign 2_n618 = 2_n87 & 2_n602;
assign 2_n709 = 2_n110 | 2_n377;
assign 2_n908 = 2_n1739 | 2_n1116;
assign 2_n813 = ~(2_n721 | 2_n775);
assign 2_n578 = ~2_n635;
assign 2_n1236 = 2_n531 | 2_n1701;
assign 2_n736 = 2_n1190 | 2_n1493;
assign 2_n49 = 2_n1180 & 2_n163;
assign 2_n1359 = ~(2_n654 ^ 2_n901);
assign 2_n1270 = 2_n313 | 2_n105;
assign 2_n877 = 2_n1276 & 2_n757;
assign 2_n1160 = ~(2_n570 | 2_n1505);
assign 2_n1318 = 2_n668 & 2_n754;
assign 2_n363 = ~(2_n1416 ^ 2_n142);
assign 2_n1531 = ~(2_n573 | 2_n759);
assign 2_n1681 = 2_n1560 & 2_n1025;
assign 2_n940 = ~(2_n579 ^ 2_n756);
assign 2_n886 = ~2_n728;
assign 2_n1124 = ~(2_n257 | 2_n1616);
assign 2_n85 = 2_n153;
assign 2_n1207 = ~(2_n1317 ^ 2_n1572);
assign 2_n1542 = ~(2_n644 | 2_n1484);
assign 2_n1475 = ~(2_n1392 ^ 2_n1592);
assign 2_n619 = 2_n107 & 2_n1206;
assign 2_n711 = ~(2_n1574 | 2_n1650);
assign 2_n1248 = 2_n1321 | 2_n1217;
assign 2_n295 = 2_n1396 & 2_n326;
assign 2_n766 = ~(2_n1019 ^ 2_n203);
assign 2_n53 = 2_n1591 | 2_n1478;
assign 2_n173 = 2_n823;
assign 2_n384 = ~(2_n471 ^ 2_n68);
assign 2_n36 = 2_n1681 & 2_n1539;
assign 2_n263 = ~2_n308;
assign 2_n907 = ~(2_n750 ^ 2_n293);
assign 2_n297 = 2_n345 | 2_n384;
assign 2_n558 = ~2_n977;
assign 2_n844 = ~2_n1468;
assign 2_n909 = 2_n26 | 2_n238;
assign 2_n873 = 2_n858 | 2_n978;
assign 2_n517 = 2_n398 | 2_n1198;
assign 2_n751 = ~(2_n1021 ^ 2_n725);
assign 2_n453 = 2_n1359;
assign 2_n925 = ~2_n248;
assign 2_n623 = 2_n258 | 2_n1113;
assign 2_n1487 = 2_n271 | 2_n51;
assign 2_n1029 = 2_n1184 | 2_n1153;
assign 2_n208 = ~(2_n478 & 2_n1095);
assign 2_n672 = 2_n468 & 2_n322;
assign 2_n767 = ~(2_n580 ^ 2_n1043);
assign 2_n1518 = 2_n361 | 2_n1272;
assign 2_n1654 = 2_n19 | 2_n1098;
assign 2_n1529 = 2_n199 & 2_n1451;
assign 2_n72 = ~(2_n929 ^ 2_n650);
assign 2_n713 = 2_n36 | 2_n387;
assign 2_n636 = ~(2_n133 ^ 2_n857);
assign 2_n464 = ~(2_n868 | 2_n829);
assign 2_n19 = ~(2_n353 ^ 2_n1291);
assign 2_n237 = ~(2_n722 ^ 2_n222);
assign 2_n1046 = ~2_n1310;
assign 2_n351 = ~2_n613;
assign 2_n825 = ~(2_n8 ^ 2_n1262);
assign 2_n1704 = 2_n902 & 2_n1650;
assign 2_n68 = 2_n909 & 2_n1703;
assign 2_n1595 = 2_n1447 | 2_n819;
assign 2_n1588 = 2_n956 | 2_n1334;
assign 2_n783 = ~2_n772;
assign 2_n1453 = ~2_n441;
assign 2_n786 = ~(2_n7 | 2_n911);
assign 2_n366 = 2_n776 | 2_n608;
assign 2_n878 = 2_n1041 & 2_n899;
assign 2_n1669 = 2_n1713 & 2_n1269;
assign 2_n1294 = ~2_n1251;
assign 2_n1062 = 2_n900 | 2_n727;
assign 2_n1178 = 2_n614 | 2_n649;
assign 2_n1258 = 2_n1378 | 2_n1348;
assign 2_n1678 = 2_n988 | 2_n1743;
assign 2_n945 = 2_n508 | 2_n1460;
assign 2_n1304 = 2_n1222 & 2_n314;
assign 2_n797 = ~2_n33;
assign 2_n270 = 2_n837 & 2_n519;
assign 2_n1697 = ~(2_n911 | 2_n253);
assign 2_n1587 = 2_n1375 | 2_n120;
assign 2_n1112 = ~2_n945;
assign 2_n583 = 2_n446 & 2_n646;
assign 2_n44 = ~(2_n1583 ^ 2_n856);
assign 2_n1649 = ~(2_n721 | 2_n399);
assign 2_n1643 = ~(2_n636 | 2_n1409);
assign 2_n604 = 2_n977 & 2_n1756;
assign 2_n995 = ~(2_n201 | 2_n1395);
assign 2_n8 = 2_n784 | 2_n321;
assign 2_n792 = ~2_n1572;
assign 2_n81 = 2_n1120 | 2_n994;
assign 2_n1322 = 2_n1590 | 2_n426;
assign 2_n446 = ~2_n28;
assign 2_n205 = ~2_n993;
assign 2_n428 = 2_n1588;
assign 2_n1755 = ~(2_n602 | 2_n45);
assign 2_n555 = 2_n1331 | 2_n1601;
assign 2_n74 = ~2_n1226;
assign 2_n1466 = 2_n254 & 2_n491;
assign 2_n1561 = 2_n1289 & 2_n197;
assign 2_n1632 = 2_n1186;
assign 2_n133 = 2_n853 & 2_n959;
assign 2_n1254 = 2_n673 & 2_n1224;
assign 2_n1422 = 2_n461 | 2_n1667;
assign 2_n1611 = 2_n1199 | 2_n325;
assign 2_n1424 = ~(2_n603 | 2_n715);
assign 2_n1111 = ~2_n489;
assign 2_n854 = 2_n1720 | 2_n39;
assign 2_n657 = 2_n669 | 2_n126;
assign 2_n1042 = 2_n1566;
assign 2_n360 = 2_n672 | 2_n1395;
assign 2_n493 = 2_n1594 | 2_n1587;
assign 2_n540 = ~(2_n888 ^ 2_n134);
assign 2_n22 = 2_n1027 | 2_n1549;
assign 2_n255 = ~(2_n1054 & 2_n1040);
assign 2_n322 = 2_n568 & 2_n703;
assign 2_n1514 = 2_n598 & 2_n444;
assign 2_n216 = ~(2_n1462 ^ 2_n1746);
assign 2_n708 = ~2_n706;
assign 2_n757 = 2_n462 | 2_n1;
assign 2_n902 = ~(2_n1311 ^ 2_n991);
assign 2_n725 = 2_n660 | 2_n1599;
assign 2_n1089 = ~2_n1388;
assign 2_n1598 = 2_n515 & 2_n495;
assign 2_n1082 = ~(2_n611 ^ 2_n1109);
assign 2_n935 = ~2_n612;
assign 2_n1729 = 2_n138;
assign 2_n1153 = 2_n140 & 2_n637;
assign 2_n43 = 2_n624 | 2_n250;
assign 2_n576 = 2_n311 & 2_n789;
assign 2_n726 = 2_n1296;
assign 2_n903 = 2_n1652 & 2_n1708;
assign 2_n1410 = ~(2_n613 ^ 2_n968);
assign 2_n1505 = ~2_n982;
assign 2_n92 = ~(2_n513 ^ 2_n90);
assign 2_n1580 = ~(2_n587 | 2_n1554);
assign 2_n723 = 2_n1579 ^ 2_n1026;
assign 2_n1285 = 2_n1401;
assign 2_n440 = ~(2_n846 | 2_n1610);
assign 2_n1102 = ~2_n984;
assign 2_n884 = ~(2_n602 | 2_n1656);
assign 2_n1653 = ~(2_n1135 | 2_n1125);
assign 2_n585 = 2_n553;
assign 2_n281 = ~2_n295;
assign 2_n319 = ~(2_n593 & 2_n1286);
assign 2_n445 = 2_n1523 & 2_n900;
assign 2_n501 = 2_n200;
assign 2_n1257 = 2_n1656 | 2_n1486;
assign 2_n450 = 2_n1047 | 2_n528;
assign 2_n1665 = ~(2_n1694 ^ 2_n1279);
assign 2_n1141 = ~(2_n1196 | 2_n342);
assign 2_n356 = ~(2_n49 | 2_n1718);
assign 2_n528 = ~(2_n1248 | 2_n320);
assign 2_n186 = 2_n19 | 2_n1199;
assign 2_n834 = 2_n302 & 2_n496;
assign 2_n818 = 2_n172 ^ 2_n1456;
assign 2_n330 = ~(2_n14 | 2_n1284);
assign 2_n122 = ~(2_n1640 | 2_n718);
assign 2_n791 = ~2_n998;
assign 2_n28 = 2_n1235 | 2_n486;
assign 2_n1450 = ~2_n742;
assign 2_n597 = ~(2_n1179 ^ 2_n321);
assign 2_n1337 = 2_n1138;
assign 2_n402 = 2_n1499 | 2_n466;
assign 2_n1031 = 2_n34 | 2_n1168;
assign 2_n875 = ~(2_n974 | 2_n1170);
assign 2_n1010 = 2_n303 | 2_n160;
assign 2_n656 = 2_n190 | 2_n1168;
assign 2_n1110 = ~2_n323;
assign 2_n495 = ~2_n982;
assign 2_n1130 = ~(2_n79 ^ 2_n535);
assign 2_n1385 = 2_n1596 | 2_n1466;
assign 2_n146 = 2_n632 | 2_n763;
assign 2_n1198 = ~(2_n1072 | 2_n42);
assign 2_n1261 = ~(2_n154 ^ 2_n567);
assign 2_n1104 = ~2_n138;
assign 2_n1485 = 2_n1163 | 2_n826;
assign 2_n210 = 2_n926 | 2_n252;
assign 2_n888 = ~(2_n1740 ^ 2_n374);
assign 2_n1619 = ~(2_n28 | 2_n1754);
assign 2_n898 = 2_n68 ^ 2_n406;
assign 2_n796 = ~2_n243;
assign 2_n1165 = ~2_n950;
assign 2_n780 = ~2_n880;
assign 2_n24 = ~2_n568;
assign 2_n1147 = 2_n1550 | 2_n629;
assign 2_n704 = ~2_n1303;
assign 2_n1489 = 2_n1535 | 2_n928;
assign 2_n1367 = ~(2_n769 | 2_n792);
assign 2_n497 = 2_n1656;
assign 2_n1351 = 2_n1694 & 2_n39;
assign 2_n841 = 2_n63 & 2_n382;
assign 2_n1402 = 2_n1680 & 2_n656;
assign 2_n1711 = ~(2_n74 ^ 2_n1344);
assign 2_n904 = 2_n558 & 2_n960;
assign 2_n584 = 2_n471 | 2_n647;
assign 2_n1579 = 2_n870 | 2_n601;
assign 2_n890 = ~2_n671;
assign 2_n793 = ~(2_n1287 ^ 2_n1661);
assign 2_n168 = ~(2_n1228 | 2_n576);
assign 2_n538 = 2_n140 | 2_n1078;
assign 2_n1266 = ~2_n1616;
assign 2_n62 = ~2_n506;
assign 2_n795 = ~(2_n385 ^ 2_n92);
assign 2_n688 = ~(2_n545 | 2_n264);
assign 2_n531 = 2_n562 & 2_n1356;
assign 2_n277 = ~(2_n1577 ^ 2_n815);
assign 2_n629 = ~(2_n949 ^ 2_n375);
assign 2_n1328 = ~2_n1114;
assign 2_n1115 = ~2_n392;
assign 2_n1341 = ~2_n487;
assign 2_n1720 = 2_n1104 & 2_n1530;
assign 2_n304 = 2_n420 & 2_n832;
assign 2_n543 = ~2_n1529;
assign 2_n1131 = ~2_n1717;
assign 2_n1309 = ~2_n500;
assign 2_n164 = ~(2_n1672 ^ 2_n482);
assign 2_n739 = 2_n37 & 2_n1511;
assign 2_n1161 = 2_n1136 | 2_n980;
assign 2_n876 = 2_n1093 & 2_n1384;
assign 2_n527 = 2_n1228 & 2_n689;
assign 2_n264 = ~(2_n1714 ^ 2_n954);
assign 2_n1074 = ~2_n1283;
assign 2_n901 = 2_n639 | 2_n1693;
assign 2_n513 = 2_n237 ^ 2_n468;
assign 2_n548 = 2_n847 | 2_n1222;
assign 2_n983 = ~(2_n335 | 2_n1663);
assign 2_n523 = ~(2_n276 | 2_n1134);
assign 2_n762 = ~(2_n183 | 2_n1678);
assign 2_n467 = ~(2_n1083 ^ 2_n1492);
assign 2_n1635 = 2_n1692 & 2_n1372;
assign 2_n565 = 2_n1422 | 2_n746;
assign 2_n1343 = 2_n658 & 2_n869;
assign 2_n1090 = ~(2_n1291 ^ 2_n1165);
assign 2_n191 = ~2_n604;
assign 2_n703 = ~2_n237;
assign 2_n149 = 2_n586 & 2_n1462;
assign 2_n569 = 2_n193 | 2_n1222;
assign 2_n613 = ~(2_n543 ^ 2_n1401);
assign 2_n401 = ~2_n589;
assign 2_n675 = ~(2_n1546 ^ 2_n1091);
assign 2_n413 = ~2_n308;
assign 2_n978 = 2_n490 & 2_n158;
assign 2_n1097 = 2_n1377 | 2_n1201;
assign 2_n345 = ~2_n101;
assign 2_n415 = 2_n958 & 2_n490;
assign 2_n1680 = 2_n1089 | 2_n153;
assign 2_n1737 = ~(2_n785 ^ 2_n1392);
assign 2_n1030 = ~(2_n285 ^ 2_n215);
assign 2_n1731 = 2_n899 & 2_n499;
assign 2_n1260 = 2_n1605 | 2_n618;
assign 2_n918 = 2_n657 | 2_n828;
assign 2_n700 = 2_n1223 | 2_n279;
assign 2_n1159 = ~(2_n1404 ^ 2_n1233);
assign 2_n127 = ~(2_n1733 | 2_n1000);
assign 2_n518 = ~(2_n1742 ^ 2_n893);
assign 2_n939 = ~2_n1018;
assign 2_n2 = ~2_n986;
assign 2_n837 = ~(2_n1317 ^ 2_n626);
assign 2_n673 = ~2_n698;
assign 2_n1388 = ~2_n1314;
assign 2_n911 = ~2_n994;
assign 2_n625 = ~(2_n1236 ^ 2_n1465);
assign 2_n1176 = 2_n1260 & 2_n1725;
assign 2_n870 = 2_n1631 & 2_n580;
assign 2_n16 = ~(2_n322 ^ 2_n1270);
assign 2_n508 = 2_n296 | 2_n1634;
assign 2_n720 = ~(2_n996 | 2_n1284);
assign 2_n836 = ~2_n1156;
assign 2_n605 = 2_n291 | 2_n530;
assign 2_n1671 = ~(2_n1385 ^ 2_n722);
assign 2_n761 = ~(2_n257 | 2_n408);
assign 2_n521 = ~2_n1451;
assign 2_n1329 = 2_n979 | 2_n647;
assign 2_n816 = ~(2_n688 | 2_n1580);
assign 2_n354 = ~(2_n374 | 2_n1646);
assign 2_n1638 = 2_n627 | 2_n559;
assign 2_n1705 = 2_n533 | 2_n9;
assign 2_n196 = 2_n835 | 2_n1566;
assign 2_n724 = 2_n425 | 2_n333;
assign 2_n1503 = ~2_n347;
assign 2_n1426 = 2_n882 & 2_n1405;
assign 2_n472 = ~(2_n1019 | 2_n1240);
assign 2_n1232 = ~(2_n653 ^ 2_n695);
assign 2_n325 = 2_n1118 | 2_n404;
assign 2_n381 = 2_n267 | 2_n705;
assign 2_n1510 = ~2_n321;
assign 2_n1577 = 2_n1161 & 2_n1538;
assign 2_n1391 = ~(2_n14 ^ 2_n833);
assign 2_n696 = ~(2_n899 | 2_n1264);
assign 2_n398 = ~(2_n1085 | 2_n830);
assign 2_n1650 = ~2_n738;
assign 2_n1100 = 2_n1039 | 2_n135;
assign 2_n404 = ~2_n1593;
assign 2_n1262 = 2_n1677 | 2_n939;
assign 2_n666 = 2_n607 & 2_n1004;
assign 2_n1723 = ~2_n502;
assign 2_n782 = 2_n222;
assign 2_n630 = ~2_n1295;
assign 2_n347 = 2_n1614 | 2_n295;
assign 2_n830 = 2_n696 | 2_n1743;
assign 2_n1003 = ~2_n227;
assign 2_n1724 = 2_n1576 & 2_n1458;
assign 2_n462 = 2_n594 | 2_n1741;
assign 2_n1284 = 2_n98 | 2_n1064;
assign 2_n294 = ~(2_n1263 | 2_n780);
assign 2_n648 = ~(2_n311 ^ 2_n820);
assign 2_n938 = 2_n1584 | 2_n1264;
assign 2_n336 = ~2_n631;
assign 2_n57 = 2_n116 | 2_n1405;
assign 2_n1200 = 2_n666 | 2_n207;
assign 2_n1362 = 2_n1020 & 2_n583;
assign 2_n1421 = 2_n695;
assign 2_n892 = ~2_n507;
assign 2_n1049 = 2_n1535 | 2_n661;
assign 2_n1564 = ~2_n1385;
assign 2_n612 = 2_n1369 | 2_n530;
assign 2_n1 = ~(2_n1245 | 2_n1444);
assign 2_n759 = 2_n1722 | 2_n614;
assign 2_n27 = 2_n947;
assign 2_n1001 = ~2_n622;
assign 2_n1116 = ~(2_n278 ^ 2_n346);
assign 2_n83 = 2_n1259 | 2_n521;
assign 2_n1423 = ~(2_n1145 | 2_n1318);
assign 2_n840 = 2_n736 & 2_n697;
assign 2_n912 = 2_n187 | 2_n1130;
assign 2_n1211 = 2_n1241 | 2_n897;
assign 2_n342 = ~2_n904;
assign 2_n61 = ~(2_n1333 | 2_n1395);
assign 2_n1535 = ~2_n1747;
assign 2_n1651 = ~(2_n1123 ^ 2_n940);
assign 2_n1185 = ~(2_n721 | 2_n1301);
assign 2_n238 = ~2_n413;
assign 2_n715 = ~(2_n680 | 2_n622);
assign 2_n1127 = ~2_n600;
assign 2_n339 = ~(2_n1303 ^ 2_n408);
assign 2_n1601 = ~2_n266;
assign 2_n37 = 2_n293 | 2_n269;
assign 2_n827 = 2_n127 | 2_n1158;
assign 2_n1575 = 2_n629 | 2_n1620;
assign 2_n1280 = 2_n1020 & 2_n1414;
assign 2_n1431 = 2_n248 & 2_n1240;
assign 2_n355 = ~(2_n721 | 2_n374);
assign 2_n343 = 2_n1453 | 2_n1499;
assign 2_n1620 = ~(2_n1494 ^ 2_n664);
assign 2_n5 = 2_n57 & 2_n605;
assign 2_n634 = ~(2_n1581 | 2_n1606);
assign 2_n31 = 2_n721 | 2_n1592;
assign 2_n714 = 2_n1036 | 2_n995;
assign 2_n1055 = 2_n1412 ^ 2_n74;
assign 2_n296 = 2_n1342 & 2_n1392;
assign 2_n7 = 2_n14 | 2_n448;
assign 2_n108 = ~2_n722;
assign 2_n891 = ~(2_n1642 ^ 2_n920);
assign 2_n226 = ~(2_n1149 | 2_n868);
assign 2_n1412 = 2_n1732 & 2_n635;
assign 2_n1390 = ~2_n756;
assign 2_n352 = 2_n1463;
assign 2_n1630 = ~2_n77;
assign 2_n1192 = ~(2_n547 | 2_n942);
assign 2_n417 = 2_n399;
assign 2_n1732 = 2_n890 | 2_n257;
assign 2_n1242 = ~2_n601;
assign 2_n1319 = 2_n125 & 2_n1602;
assign 2_n942 = ~(2_n1181 | 2_n599);
assign 2_n494 = 2_n1607 | 2_n122;
assign 2_n328 = ~(2_n900 | 2_n831);
assign 2_n603 = 2_n680 & 2_n274;
assign 2_n915 = ~2_n82;
assign 2_n1032 = 2_n1376 | 2_n238;
assign 2_n965 = 2_n1755 | 2_n1709;
assign 2_n321 = ~(2_n266 ^ 2_n612);
assign 2_n130 = 2_n1592;
assign 2_n553 = 2_n450 | 2_n1010;
assign 2_n1498 = ~(2_n311 ^ 2_n945);
assign 2_n1068 = 2_n1722 | 2_n614;
assign 2_n1296 = ~2_n992;
assign 2_n1615 = 2_n545 & 2_n283;
assign 2_n1583 = 2_n1129 | 2_n843;
assign 2_n1667 = ~2_n473;
assign 2_n1581 = 2_n494 | 2_n91;
assign 2_n1252 = ~2_n1569;
assign 2_n1540 = ~(2_n98 ^ 2_n837);
assign 2_n562 = ~(2_n698 | 2_n1108);
assign 2_n55 = ~(2_n628 | 2_n1469);
assign 2_n1186 = 2_n1047 | 2_n872;
assign 2_n716 = 2_n231 & 2_n795;
assign 2_n1101 = 2_n969 & 2_n1206;
assign 2_n457 = 2_n827 | 2_n1452;
assign 2_n1063 = ~(2_n613 ^ 2_n136);
assign 2_n1356 = 2_n1444 | 2_n1001;
assign 2_n1331 = 2_n1222 & 2_n1411;
assign 2_n1238 = 2_n1171 | 2_n1457;
assign 2_n405 = 2_n1353 | 2_n290;
assign 2_n756 = 2_n141 & 2_n1688;
assign 2_n1069 = 2_n257 | 2_n220;
assign 2_n1683 = 2_n1669 & 2_n682;
assign 2_n1093 = 2_n257 | 2_n293;
assign 2_n1004 = ~2_n1314;
assign 2_n642 = 2_n1450 | 2_n530;
assign 2_n217 = 2_n550 | 2_n415;
assign 2_n160 = 2_n485 | 2_n563;
assign 2_n1136 = ~2_n413;
assign 2_n1373 = ~(2_n753 ^ 2_n767);
assign 2_n403 = 2_n1351 | 2_n720;
assign 2_n763 = ~(2_n179 ^ 2_n1595);
assign 2_n1077 = 2_n298 | 2_n1458;
assign 2_n730 = 2_n1455 | 2_n1348;
assign 2_n1065 = ~(2_n592 ^ 2_n305);
assign 2_n1419 = ~(2_n1385 ^ 2_n1463);
assign 2_n678 = ~2_n1595;
assign 2_n491 = ~2_n413;
assign 2_n1000 = ~2_n1581;
assign 2_n954 = ~(2_n896 ^ 2_n1169);
assign 2_n833 = 2_n1705 | 2_n480;
assign 2_n198 = ~2_n569;
assign 2_n776 = ~2_n1388;
assign 2_n1657 = 2_n414 | 2_n329;
assign 2_n162 = ~2_n1428;
assign 2_n1471 = 2_n316 | 2_n191;
assign 2_n951 = 2_n19 | 2_n1098;
assign 2_n475 = ~2_n1149;
assign 2_n1554 = 2_n1179 | 2_n1128;
assign 2_n193 = ~2_n54;
assign 2_n1330 = ~(2_n1165 | 2_n970);
assign 2_n110 = 2_n1567 | 2_n683;
assign 2_n948 = 2_n1293 & 2_n844;
assign 2_n1744 = ~(2_n55 | 2_n911);
assign 2_n1547 = 2_n420;
assign 2_n897 = ~(2_n1733 | 2_n634);
assign 2_n1405 = ~2_n728;
assign 2_n1726 = ~(2_n1206 | 2_n1205);
assign 2_n712 = ~(2_n1041 | 2_n904);
assign 2_n1491 = ~2_n964;
assign 2_n1377 = 2_n725 ^ 2_n1566;
assign 2_n498 = 2_n293;
assign 2_n1672 = ~(2_n785 ^ 2_n318);
assign 2_n1433 = 2_n95 | 2_n332;
assign 2_n1157 = 2_n712 & 2_n235;
assign 2_n1591 = ~(2_n1512 | 2_n69);
assign 2_n1605 = 2_n1753 & 2_n1222;
assign 2_n194 = 2_n867 | 2_n1522;
assign 2_n1552 = ~2_n510;
assign 2_n224 = 2_n699 | 2_n1744;
assign 2_n407 = 2_n1358 & 2_n178;
assign 2_n1473 = 2_n182 | 2_n328;
assign 2_n649 = ~(2_n551 ^ 2_n1011);
assign 2_n1139 = 2_n101 | 2_n384;
assign 2_n141 = ~(2_n1319 | 2_n259);
assign 2_n421 = ~(2_n652 ^ 2_n1467);
assign 2_n826 = 2_n282 & 2_n302;
assign 2_n1464 = 2_n784 | 2_n1544;
assign 2_n1574 = ~(2_n134 | 2_n88);
assign 2_n1610 = ~(2_n431 ^ 2_n411);
assign 2_n591 = ~2_n1647;
assign 2_n1546 = ~(2_n1416 ^ 2_n115);
assign 2_n1551 = ~2_n869;
assign 2_n1013 = ~2_n71;
assign 2_n456 = 2_n1705 ^ 2_n572;
assign 2_n1038 = ~(2_n283 | 2_n1336);
assign 2_n1181 = 2_n1179 | 2_n716;
assign 2_n1682 = ~(2_n1635 ^ 2_n1656);
assign 2_n1066 = ~2_n1059;
assign 2_n566 = ~(2_n1520 & 2_n1613);
assign 2_n1012 = 2_n973 | 2_n17;
assign 2_n1557 = 2_n367 & 2_n1229;
assign 2_n919 = 2_n1658 & 2_n711;
assign 2_n852 = 2_n1654 | 2_n1611;
assign 2_n1436 = ~2_n1490;
assign 2_n974 = 2_n876 | 2_n1045;
assign 2_n972 = 2_n1397 | 2_n1070;
assign 2_n722 = 2_n151 | 2_n484;
assign 2_n1369 = ~2_n1205;
assign 2_n131 = 2_n1117 | 2_n106;
assign 2_n934 = 2_n1540 | 2_n348;
assign 2_n1451 = 2_n850 | 2_n1555;
assign 2_n275 = 2_n1296;
assign 2_n917 = ~(2_n846 ^ 2_n48);
assign 2_n1118 = 2_n232 | 2_n67;
assign 2_n444 = ~2_n808;
assign 2_n1203 = 2_n368 | 2_n1014;
assign 2_n479 = 2_n45 | 2_n1352;
assign 2_n60 = ~(2_n1682 ^ 2_n941);
assign 2_n218 = ~2_n1682;
assign 2_n459 = 2_n300 & 2_n835;
assign 2_n1206 = ~2_n413;
assign 2_n1298 = ~2_n1276;
assign 2_n1005 = ~(2_n467 | 2_n363);
assign 2_n1544 = ~2_n571;
assign 2_n1666 = ~(2_n338 | 2_n1653);
assign 2_n439 = ~(2_n814 ^ 2_n256);
assign 2_n215 = ~(2_n1439 ^ 2_n1525);
assign 2_n1008 = 2_n104 | 2_n15;
assign 2_n1652 = 2_n239 | 2_n1405;
assign 2_n1452 = 2_n1280 | 2_n1362;
assign 2_n225 = ~(2_n972 ^ 2_n45);
assign 2_n449 = ~(2_n1638 ^ 2_n986);
assign 2_n1195 = 2_n1704 | 2_n919;
assign 2_n764 = 2_n1674 | 2_n1143;
assign 2_n368 = ~(2_n1295 ^ 2_n188);
assign 2_n499 = ~2_n235;
assign 2_n526 = 2_n294 | 2_n1094;
assign 2_n1685 = ~(2_n876 ^ 2_n903);
assign 2_n1413 = 2_n1676 & 2_n1618;
assign 2_n982 = 2_n490 | 2_n937;
assign 2_n1690 = 2_n975 | 2_n139;
assign 2_n532 = ~2_n1573;
assign 2_n1686 = ~2_n1039;
assign 2_n1492 = 2_n1185 | 2_n1480;
assign 2_n334 = ~(2_n405 | 2_n855);
assign 2_n6 = ~(2_n1489 ^ 2_n806);
assign 2_n106 = 2_n204 & 2_n339;
assign 2_n931 = ~(2_n1123 ^ 2_n383);
assign 2_n105 = 2_n913 | 2_n554;
assign 2_n773 = 2_n980;
assign 2_n1174 = 2_n1074 | 2_n1555;
assign 2_n628 = ~(2_n1608 | 2_n1282);
assign 2_n1702 = ~(2_n121 | 2_n42);
assign 2_n814 = ~(2_n1228 | 2_n311);
assign 2_n1241 = 2_n986 & 2_n737;
assign 2_n1567 = 2_n1578 | 2_n286;
assign 2_n397 = ~2_n664;
assign 2_n679 = 2_n949 & 2_n375;
assign 2_n111 = ~(2_n438 ^ 2_n410);
assign 2_n353 = 2_n31 & 2_n1031;
assign 2_n1308 = 2_n1111 | 2_n1555;
assign 2_n1312 = 2_n1723 | 2_n444;
assign 2_n1679 = ~(2_n962 ^ 2_n860);
assign 2_n317 = 2_n834 | 2_n817;
assign 2_n247 = ~(2_n1700 ^ 2_n1325);
assign 2_n640 = 2_n1345;
assign 2_n1376 = ~2_n953;
assign 2_n855 = ~(2_n1358 | 2_n673);
assign 2_n1027 = ~(2_n1570 | 2_n765);
assign 2_n1223 = ~(2_n993 | 2_n908);
assign 2_n349 = 2_n1624 | 2_n861;
assign 2_n309 = ~2_n1448;
assign 2_n985 = ~(2_n1147 | 2_n1096);
assign 2_n868 = 2_n1214 | 2_n1700;
assign 2_n1026 = ~2_n267;
assign 2_n617 = 2_n685 | 2_n336;
assign 2_n535 = ~(2_n174 ^ 2_n674);
assign 2_n853 = 2_n1206 | 2_n138;
assign 2_n971 = ~2_n341;
assign 2_n1631 = ~2_n823;
assign 2_n1208 = 2_n78 & 2_n435;
assign 2_n370 = ~(2_n339 ^ 2_n334);
assign 2_n59 = ~(2_n546 ^ 2_n12);
assign 2_n851 = ~(2_n513 ^ 2_n16);
assign 2_n541 = 2_n162 | 2_n238;
assign 2_n889 = ~(2_n257 | 2_n1345);
assign 2_n203 = ~(2_n811 ^ 2_n1672);
assign 2_n158 = ~(2_n44 ^ 2_n931);
assign 2_n748 = 2_n1684 | 2_n511;
assign 2_n95 = ~2_n406;
assign 2_n395 = ~(2_n1171 | 2_n1457);
assign 2_n201 = ~(2_n888 ^ 2_n1270);
assign 2_n937 = ~(2_n1360 | 2_n1230);
assign 2_n18 = 2_n729 & 2_n900;
assign 2_n575 = ~2_n490;
assign 2_n842 = 2_n1205;
assign 2_n1628 = ~(2_n257 | 2_n246);
assign 2_n144 = 2_n1751 | 2_n6;
assign 2_n998 = 2_n197 | 2_n18;
assign 2_n994 = 2_n1503 | 2_n713;
assign 2_n529 = ~2_n641;
assign 2_n1721 = ~2_n539;
assign 2_n1562 = ~(2_n1748 | 2_n360);
assign 2_n741 = ~2_n37;
assign 2_n1549 = ~(2_n525 | 2_n495);
assign 2_n3 = ~(2_n1206 | 2_n487);
assign 2_n684 = ~2_n1092;
assign 2_n234 = ~(2_n93 ^ 2_n1471);
assign 2_n789 = 2_n757 | 2_n944;
assign 2_n1429 = ~2_n1583;
assign 2_n685 = 2_n692 & 2_n1188;
assign 2_n371 = 2_n586 | 2_n1715;
assign 2_n996 = 2_n731 | 2_n14;
assign 2_n280 = 2_n1418 & 2_n257;
assign 2_n241 = ~2_n1610;
assign 2_n881 = ~(2_n166 ^ 2_n520);
assign 2_n1006 = ~(2_n237 ^ 2_n1395);
assign 2_n361 = ~(2_n702 | 2_n147);
assign 2_n1081 = 2_n865 & 2_n621;
assign 2_n615 = ~(2_n165 ^ 2_n1028);
assign 2_n65 = ~(2_n368 | 2_n1014);
assign 2_n988 = ~2_n1756;
assign 2_n622 = ~(2_n1441 ^ 2_n234);
assign 2_n860 = ~(2_n1256 ^ 2_n766);
assign 2_n1024 = ~(2_n812 ^ 2_n1662);
assign 2_n594 = 2_n1603 | 2_n878;
assign 2_n632 = 2_n167 & 2_n1730;
assign 2_n848 = 2_n1516 & 2_n1222;
assign 2_n1096 = 2_n924 | 2_n35;
assign 2_n455 = ~(2_n648 ^ 2_n881);
assign 2_n1508 = 2_n1735 & 2_n1710;
assign 2_n101 = 2_n266 | 2_n791;
assign 2_n922 = ~(2_n843 ^ 2_n856);
assign 2_n283 = 2_n473 & 2_n1677;
assign 2_n236 = ~(2_n1489 ^ 2_n1751);
assign 2_n737 = 2_n1638 | 2_n1110;
assign 2_n1379 = 2_n310 & 2_n240;
assign 2_n172 = 2_n541 & 2_n419;
assign 2_n1699 = ~(2_n1173 ^ 2_n1332);
assign 2_n707 = 2_n400 | 2_n1522;
assign 2_n880 = 2_n63 & 2_n1069;
assign 2_n1728 = ~(2_n451 | 2_n96);
assign 2_n1288 = 2_n912 | 2_n128;
assign 2_n1047 = 2_n1218 | 2_n429;
assign 2_n1703 = 2_n1076 | 2_n1004;
assign 2_n788 = ~2_n1282;
assign 2_n520 = 2_n289 & 2_n1112;
assign 2_n1137 = 2_n1106 & 2_n888;
assign 2_n976 = ~2_n448;
assign 2_n1039 = ~(2_n689 ^ 2_n925);
assign 2_n1233 = ~(2_n924 ^ 2_n1494);
assign 2_n214 = 2_n690 & 2_n1711;
assign 2_n1122 = 2_n542 & 2_n639;
assign 2_n1593 = 2_n65 & 2_n365;
assign 2_n643 = 2_n637 & 2_n1357;
assign 2_n1408 = ~(2_n83 | 2_n1008);
assign 2_n1363 = ~(2_n1045 | 2_n1685);
assign 2_n1752 = 2_n118 | 2_n208;
assign 2_n358 = ~2_n1597;
assign 2_n1742 = 2_n1472 | 2_n1633;
assign 2_n1371 = 2_n590 & 2_n1643;
assign 2_n932 = 2_n131 | 2_n464;
assign 2_n480 = 2_n1462 & 2_n270;
assign 2_n680 = 2_n1151 & 2_n1444;
assign 2_n424 = ~2_n1071;
assign 2_n176 = ~(2_n1683 | 2_n281);
assign 2_n114 = 2_n1533 | 2_n1431;
assign 2_n1053 = 2_n1176 | 2_n1274;
assign 2_n1559 = 2_n1066 & 2_n1311;
assign 2_n1589 = 2_n154 ^ 2_n1740;
assign 2_n1528 = 2_n1252 | 2_n1136;
assign 2_n702 = 2_n1197 | 2_n678;
assign 2_n15 = 2_n1227 & 2_n602;
assign 2_n169 = ~(2_n1433 | 2_n616);
assign 2_n1707 = 2_n895 ^ 2_n551;
assign 2_n862 = ~2_n36;
assign 2_n84 = ~2_n1345;
assign 2_n1249 = ~(2_n871 ^ 2_n1258);
assign 2_n150 = ~2_n689;
assign 2_n705 = ~2_n732;
assign 2_n1603 = ~(2_n1301 | 2_n1675);
assign 2_n1670 = ~(2_n93 ^ 2_n604);
assign 2_n1245 = 2_n1196 | 2_n1097;
assign 2_n610 = ~(2_n1600 ^ 2_n421);
assign 2_n1378 = 2_n240 & 2_n1281;
assign 2_n857 = 2_n1535 | 2_n492;
assign 2_n1368 = 2_n420;
assign 2_n1021 = 2_n733 | 2_n804;
assign 2_n434 = ~(2_n1151 | 2_n673);
assign 2_n1445 = ~(2_n78 ^ 2_n1507);
assign 2_n1469 = ~(2_n542 | 2_n788);
assign 2_n454 = ~2_n1217;
assign 2_n692 = 2_n1749 | 2_n835;
assign 2_n824 = 2_n645 & 2_n1555;
assign 2_n400 = 2_n240 & 2_n1023;
assign 2_n1641 = 2_n848 | 2_n221;
assign 2_n571 = 2_n1179 | 2_n1510;
assign 2_n964 = 2_n83 & 2_n1008;
assign 2_n1398 = ~(2_n504 ^ 2_n1265);
assign 2_n941 = 2_n330 | 2_n854;
assign 2_n1572 = 2_n63 & 2_n393;
assign 2_n952 = ~(2_n539 ^ 2_n1454);
assign 2_n1584 = ~2_n1097;
assign 2_n1684 = 2_n800 | 2_n1425;
assign 2_n627 = ~2_n156;
assign 2_n1606 = 2_n1371 & 2_n709;
assign 2_n1754 = ~(2_n768 | 2_n1490);
assign 2_n1333 = ~2_n1669;
assign 2_n1696 = ~2_n288;
assign 2_n291 = ~2_n710;
assign 2_n39 = 2_n1279 & 2_n533;
assign 2_n706 = ~(2_n923 ^ 2_n399);
assign 2_n1277 = ~(2_n1038 ^ 2_n1690);
assign 2_n968 = ~2_n893;
assign 2_n157 = ~(2_n1519 ^ 2_n1300);
assign 2_n1550 = 2_n1535 | 2_n1087;
assign 2_n411 = ~(2_n1410 ^ 2_n373);
assign 2_n147 = 2_n1171 | 2_n1457;
assign 2_n621 = 2_n210 | 2_n102;
assign 2_n1633 = ~2_n381;
assign 2_n1725 = 2_n355 | 2_n1016;
assign 2_n118 = ~(2_n581 & 2_n743);
assign 2_n1677 = ~2_n746;
assign 2_n1220 = ~(2_n331 ^ 2_n556);
assign 2_n1271 = 2_n1131 | 2_n1098;
assign 2_n1478 = 2_n1593 & 2_n349;
assign 2_n1264 = ~2_n1157;
assign 2_n1213 = ~(2_n249 | 2_n1583);
assign 2_n547 = ~(2_n545 | 2_n1423);
assign 2_n669 = 2_n1221 | 2_n433;
assign 2_n1014 = ~(2_n1512 ^ 2_n1049);
assign 2_n1311 = ~2_n1261;
assign 2_n375 = 2_n1146 | 2_n459;
assign 2_n1553 = 2_n1609 & 2_n1555;
assign 2_n966 = ~(2_n721 | 2_n1263);
assign 2_n577 = 2_n870 & 2_n1582;
assign 2_n1634 = 2_n987 & 2_n1475;
assign 2_n1640 = 2_n397 | 2_n260;
assign 2_n620 = 2_n153 | 2_n1381;
assign 2_n320 = ~2_n387;
assign 2_n76 = 2_n1136 | 2_n626;
assign 2_n1733 = 2_n97;
assign 2_n1134 = 2_n1712 | 2_n1743;
assign 2_n163 = 2_n180 | 2_n1168;
assign 2_n1342 = ~2_n1592;
assign 2_n500 = 2_n705 | 2_n351;
assign 2_n596 = ~(2_n667 ^ 2_n751);
assign 2_n595 = 2_n1301;
assign 2_n1303 = 2_n1719 | 2_n681;
assign 2_n1143 = ~2_n124;
assign 2_n665 = ~2_n829;
assign 2_n1209 = 2_n1071;
assign 2_n394 = ~(2_n458 ^ 2_n213);
assign 2_n887 = 2_n1625 | 2_n1458;
assign 2_n1057 = 2_n339 & 2_n577;
assign 2_n125 = ~2_n346;
assign 2_n66 = 2_n1440 & 2_n463;
assign 2_n1509 = 2_n835 | 2_n1278;
assign 2_n654 = ~(2_n1092 ^ 2_n986);
assign 2_n638 = 2_n420;
assign 2_n278 = ~2_n1602;
assign 2_n539 = ~(2_n580 ^ 2_n823);
assign 2_n552 = ~2_n1739;
assign 2_n674 = ~(2_n1602 ^ 2_n880);
assign 2_n843 = 2_n552 | 2_n1294;
assign 2_n438 = ~(2_n1399 ^ 2_n1344);
assign 2_n745 = 2_n663 & 2_n1136;
assign 2_n799 = ~(2_n436 ^ 2_n1488);
assign 2_n1123 = 2_n708 ^ 2_n1468;
assign 2_n1125 = ~2_n554;
assign 2_n644 = 2_n1052 | 2_n797;
assign 2_n145 = ~2_n1011;
assign 2_n1439 = ~(2_n353 ^ 2_n970);
assign 2_n1691 = ~2_n1173;
assign 2_n599 = ~(2_n231 | 2_n754);
assign 2_n650 = 2_n1343 ^ 2_n1260;
assign 2_n1292 = 2_n1616;
assign 2_n544 = 2_n673 | 2_n440;
assign 2_n116 = ~2_n1586;
assign 2_n550 = 2_n526 | 2_n700;
assign 2_n1224 = ~(2_n917 ^ 2_n1556);
assign 2_n1230 = ~2_n789;
assign 2_n1073 = ~(2_n439 ^ 2_n455);
assign 2_n1530 = 2_n1692 & 2_n863;
assign 2_n894 = ~(2_n811 ^ 2_n114);
assign 2_n1745 = ~(2_n1617 ^ 2_n596);
assign 2_n1374 = 2_n900 | 2_n391;
assign 2_n977 = 2_n920 | 2_n1504;
assign 2_n1668 = ~2_n1175;
assign 2_n452 = 2_n1412 | 2_n687;
assign 2_n1425 = 2_n296 & 2_n1672;
assign 2_n1268 = ~2_n1443;
assign 2_n838 = ~(2_n617 | 2_n1313);
assign 2_n335 = 2_n66 | 2_n1199;
assign 2_n1548 = 2_n567;
assign 2_n441 = 2_n1535 | 2_n209;
assign 2_n847 = ~2_n936;
assign 2_n51 = ~(2_n721 | 2_n947);
assign 2_n206 = 2_n1155 & 2_n548;
assign 2_n189 = 2_n368 | 2_n1014;
assign 2_n435 = 2_n571 | 2_n1232;
assign 2_n232 = ~(2_n1200 | 2_n1664);
assign 2_n161 = 2_n457;
assign 2_n568 = 2_n222 | 2_n108;
assign 2_n1265 = ~(2_n1067 ^ 2_n442);
assign 2_n425 = 2_n1222 & 2_n560;
assign 2_n1499 = ~(2_n924 ^ 2_n1550);
assign 2_n469 = ~(2_n1056 ^ 2_n898);
assign 2_n1291 = 2_n1032 & 2_n1310;
assign 2_n412 = ~(2_n941 | 2_n786);
assign 2_n276 = 2_n960 & 2_n191;
assign 2_n1025 = ~2_n1151;
assign 2_n113 = 2_n892 | 2_n1458;
assign 2_n856 = ~(2_n205 ^ 2_n249);
assign 2_n808 = ~2_n263;
assign 2_n1256 = 2_n1228 ^ 2_n1533;
assign 2_n1701 = ~(2_n136 | 2_n1424);
assign 2_n1646 = ~2_n1740;
assign 2_n689 = ~(2_n1382 ^ 2_n1446);
assign 2_n46 = ~2_n1566;
assign 2_n152 = ~(2_n960 ^ 2_n1471);
assign 2_n1558 = 2_n803 | 2_n695;
assign 2_n372 = ~(2_n353 | 2_n537);
assign 2_n1730 = 2_n796 | 2_n1168;
assign 2_n1259 = 2_n344 & 2_n197;
assign 2_n546 = ~(2_n1366 ^ 2_n1090);
assign 2_n1441 = ~(2_n812 ^ 2_n13);
assign 2_n1713 = ~(2_n1135 | 2_n1261);
assign 2_n128 = 2_n1745 | 2_n1082;
assign 2_n1674 = 2_n1215 | 2_n297;
assign 2_n423 = 2_n539 & 2_n1035;
assign 2_n694 = 2_n467 | 2_n363;
assign 2_n1533 = 2_n987 | 2_n538;
assign 2_n1751 = 2_n1535 | 2_n350;
assign 2_n1746 = ~(2_n371 | 2_n270);
assign 2_n179 = 2_n1267 | 2_n1466;
assign 2_n927 = ~(2_n257 | 2_n920);
assign 2_n1041 = 2_n46 & 2_n725;
assign 2_n652 = ~(2_n1370 | 2_n3);
assign 2_n899 = ~2_n1196;
assign 2_n580 = 2_n536 | 2_n1297;
assign 2_n389 = ~(2_n133 | 2_n1495);
assign 2_n1059 = 2_n1463 | 2_n1564;
assign 2_n1659 = ~(2_n1517 ^ 2_n1316);
assign 2_n115 = ~2_n1492;
assign 2_n949 = 2_n63 & 2_n41;
assign 2_n458 = 2_n903 ^ 2_n43;
assign 2_n274 = ~(2_n1670 ^ 2_n1024);
assign 2_n987 = 2_n1266 & 2_n623;
assign 2_n967 = ~(2_n1577 ^ 2_n1751);
assign 2_n1145 = ~(2_n668 | 2_n795);
assign 2_n258 = 2_n58 & 2_n240;
assign 2_n1354 = 2_n1020 & 2_n110;
assign 2_n313 = 2_n134 & 2_n20;
assign 2_n601 = 2_n475 | 2_n665;
assign 2_n845 = 2_n29 & 2_n1004;
assign 2_n1449 = ~(2_n284 & 2_n574);
assign 2_n1519 = 2_n1403 | 2_n371;
assign 2_n1442 = ~(2_n1535 | 2_n1612);
assign 2_n1494 = 2_n245 | 2_n1571;
assign 2_n1749 = ~2_n52;
assign 2_n1199 = ~(2_n1456 ^ 2_n631);
assign 2_n279 = 2_n205 & 2_n1183;
assign 2_n1406 = ~2_n1618;
assign 2_n207 = 2_n1246 & 2_n491;
assign 2_n1366 = ~(2_n1689 ^ 2_n818);
assign 2_n924 = 2_n76 & 2_n963;
assign 2_n482 = ~(2_n945 | 2_n1326);
assign 2_n1400 = ~2_n946;
assign 2_n13 = ~(2_n739 ^ 2_n80);
assign 2_n10 = ~2_n88;
assign 2_n1036 = ~(2_n432 | 2_n1086);
assign 2_n1108 = ~(2_n359 | 2_n274);
assign 2_n1204 = 2_n1437 | 2_n1243;
assign 2_n188 = 2_n966 | 2_n1323;
assign 2_n1594 = 2_n255 | 2_n319;
assign 2_n73 = ~(2_n152 | 2_n42);
assign 2_n1146 = ~(2_n1405 | 2_n1470);
assign 2_n1180 = 2_n1405 | 2_n1476;
assign 2_n1710 = ~(2_n1213 | 2_n495);
assign 2_n1098 = ~(2_n950 ^ 2_n633);
assign 2_n1120 = 2_n1608 & 2_n744;
assign 2_n1663 = 2_n172 | 2_n951;
assign 2_n202 = ~(2_n1026 | 2_n613);
assign 2_n1688 = ~2_n1183;
assign 2_n209 = ~2_n32;
assign 2_n171 = 2_n1458 & 2_n961;
assign 2_n136 = ~2_n698;
assign 2_n975 = ~2_n503;
assign 2_n396 = 2_n195 | 2_n1160;
assign 2_n34 = ~2_n1305;
assign 2_n1472 = ~2_n620;
assign 2_n1244 = ~(2_n186 | 2_n512);
assign 2_n1625 = ~2_n1154;
assign 2_n257 = ~2_n728;
assign 2_n1348 = 2_n299 & 2_n491;
assign 2_n781 = ~2_n785;
assign 2_n944 = ~(2_n1394 | 2_n176);
assign 2_n4 = 2_n1136 | 2_n1299;
assign 2_n1722 = ~(2_n1676 ^ 2_n1618);
assign 2_n1034 = ~(2_n763 | 2_n185);
assign 2_n1313 = 2_n19 | 2_n1098;
assign 2_n1560 = ~2_n1245;
assign 2_n1675 = ~2_n1021;
assign 2_n431 = ~(2_n202 ^ 2_n771);
assign 2_n1310 = 2_n1365 | 2_n1458;
assign 2_n871 = 2_n171 | 2_n1601;
assign 2_n633 = 2_n447 | 2_n445;
assign 2_n338 = ~(2_n1135 | 2_n388);
assign 2_n1222 = ~2_n886;
assign 2_n285 = ~(2_n123 ^ 2_n277);
assign 2_n1129 = 2_n706 & 2_n1468;
assign 2_n1255 = 2_n62 | 2_n1206;
assign 2_n910 = ~2_n841;
assign 2_n260 = ~2_n1494;
assign 2_n1275 = 2_n1474 & 2_n1168;
assign 2_n1512 = 2_n1497 & 2_n1308;
assign 2_n1364 = ~(2_n1573 ^ 2_n1629);
assign 2_n1088 = 2_n1164 & 2_n257;
assign 2_n859 = ~(2_n1459 ^ 2_n1277);
assign 2_n332 = ~2_n965;
assign 2_n1416 = 2_n196 & 2_n113;
assign 2_n572 = ~2_n1257;
assign 2_n647 = ~(2_n406 ^ 2_n965);
assign 2_n916 = ~(2_n1682 ^ 2_n911);
assign 2_n1660 = 2_n734 & 2_n240;
assign 2_n1563 = ~2_n200;
assign 2_n524 = ~2_n273;
assign 2_n556 = 2_n5 ^ 2_n1676;
assign 2_n1756 = 2_n37 | 2_n1623;
assign 2_n1327 = ~(2_n357 | 2_n103);
assign 2_n166 = 2_n1003 | 2_n1019;
assign 2_n1168 = ~2_n1314;
assign 2_n732 = ~(2_n1043 ^ 2_n153);
assign 2_n362 = 2_n914 | 2_n1361;
assign 2_n1461 = ~2_n143;
assign 2_n265 = ~2_n105;
assign 2_n1432 = 2_n925 | 2_n227;
assign 2_n282 = 2_n424 & 2_n1332;
assign 2_n204 = 2_n1568 & 2_n1641;
assign 2_n810 = 2_n809 | 2_n939;
assign 2_n1440 = 2_n1206 | 2_n1446;
assign 2_n1573 = ~(2_n0 ^ 2_n986);
assign 2_n970 = ~2_n633;
assign 2_n929 = 2_n1182 ^ 2_n179;
assign 2_n822 = ~(2_n584 | 2_n1524);
assign 2_n1456 = ~2_n685;
assign 2_n1276 = 2_n958 & 2_n643;
assign 2_n1092 = 2_n627 | 2_n1563;
assign 2_n1479 = 2_n1135 & 2_n265;
assign 2_n192 = ~(2_n1422 | 2_n697);
assign 2_n981 = ~(2_n1329 | 2_n764);
assign 2_n1210 = 2_n244 & 2_n197;
assign 2_n614 = ~(2_n49 ^ 2_n5);
assign 2_n1217 = 2_n996 | 2_n448;
assign 2_n329 = 2_n1720 & 2_n1694;
assign 2_n959 = 2_n1219 | 2_n444;
assign 2_n1334 = 2_n1380 & 2_n901;
assign 2_n955 = ~(2_n588 ^ 2_n1501);
assign 2_n586 = 2_n670 & 2_n1317;
assign 2_n770 = 2_n437 | 2_n1247;
assign 2_n1662 = ~(2_n741 ^ 2_n1157);
assign 2_n79 = ~(2_n799 ^ 2_n1737);
assign 2_n1234 = 2_n608;
assign 2_n1692 = ~2_n1565;
assign 2_n473 = ~(2_n1332 ^ 2_n1071);
assign 2_n1739 = 2_n399 | 2_n70;
assign 2_n1338 = ~(2_n1535 | 2_n813);
assign 2_n590 = ~(2_n629 | 2_n1620);
assign 2_n184 = 2_n420;
assign 2_n1420 = ~(2_n1232 ^ 2_n1464);
assign 2_n1712 = ~(2_n960 | 2_n191);
assign 2_n1300 = 2_n7 & 2_n1622;
assign 2_n311 = ~(2_n777 ^ 2_n1345);
assign 2_n979 = ~(2_n1399 ^ 2_n1412);
assign 2_n631 = 2_n1124 | 2_n280;
assign 2_n1444 = ~2_n359;
assign 2_n1706 = ~2_n789;
assign 2_n1202 = 2_n1430 | 2_n240;
assign 2_n1290 = ~2_n311;
assign 2_n664 = 2_n63 & 2_n4;
assign 2_n30 = 2_n362;
assign 2_n78 = 2_n1190 & 2_n677;
assign 2_n287 = ~2_n1446;
assign 2_n337 = 2_n626;
assign 2_n733 = 2_n1350 & 2_n530;
assign 2_n323 = 2_n156 & 2_n401;
assign 2_n1447 = ~(2_n1405 | 2_n1463);
assign 2_n1372 = 2_n803 | 2_n430;
assign 2_n667 = ~(2_n1642 ^ 2_n750);
assign 2_n1524 = 2_n68 | 2_n1736;
assign 2_n1064 = 2_n1257 | 2_n802;
assign 2_n990 = ~(2_n1694 ^ 2_n412);
assign 2_n563 = ~(2_n1248 | 2_n347);
assign 2_n1403 = ~2_n1383;
assign 2_n1295 = 2_n1692 & 2_n1062;
assign 2_n267 = 2_n1401 | 2_n1529;
assign 2_n1382 = 2_n1514 | 2_n749;
assign 2_n895 = 2_n1315 & 2_n1174;
assign 2_n1149 = 2_n620 | 2_n1721;
assign 2_n261 = ~(2_n1550 ^ 2_n397);
assign 2_n1183 = 2_n249 & 2_n1294;
assign 2_n1495 = 2_n857 | 2_n629;
assign 2_n248 = ~(2_n623 ^ 2_n1616);
assign 2_n185 = ~(2_n632 ^ 2_n1182);
assign 2_n806 = ~2_n815;
assign 2_n393 = 2_n602 | 2_n477;
assign 2_n382 = 2_n1206 | 2_n582;
assign 2_n447 = ~(2_n803 | 2_n318);
assign 2_n1636 = ~(2_n1535 ^ 2_n1338);
assign 2_n64 = 2_n1330 | 2_n372;
assign 2_n1317 = 2_n1692 & 2_n1162;
assign 2_n233 = ~(2_n1192 ^ 2_n816);
assign 2_n691 = 2_n532 & 2_n1048;
assign 2_n1163 = ~(2_n608 | 2_n1691);
assign 2_n33 = 2_n927 | 2_n619;
assign 2_n365 = ~(2_n6 | 2_n967);
assign 2_n744 = ~2_n639;
assign 2_n286 = 2_n1526 | 2_n53;
assign 2_n410 = ~(2_n418 ^ 2_n955);
assign 2_n1409 = 2_n549 | 2_n343;
assign 2_n1748 = ~(2_n999 | 2_n322);
assign 2_n865 = 2_n1005 & 2_n1363;
assign 2_n1344 = 2_n366 & 2_n642;
assign 2_n1052 = ~2_n43;
assign 2_n1481 = 2_n1706 & 2_n1679;
assign 2_n470 = ~(2_n1682 ^ 2_n1665);
assign 2_n1182 = 2_n1255 & 2_n1202;
assign 2_n290 = ~(2_n1700 | 2_n1242);
assign 2_n1504 = ~2_n1642;
assign 2_n132 = 2_n895 | 2_n1068;
assign 2_n350 = ~(2_n257 | 2_n609);
assign 2_n178 = ~2_n405;
assign 2_n109 = 2_n206 | 2_n1171;
assign 2_n1336 = 2_n662 | 2_n1532;
assign 2_n98 = ~2_n1462;
assign 2_n699 = ~(2_n1122 | 2_n81);
assign 2_n668 = 2_n317 | 2_n805;
assign 2_n1109 = ~(2_n1671 ^ 2_n1589);
assign 2_n693 = ~(2_n732 ^ 2_n390);
assign 2_n385 = ~(2_n864 ^ 2_n540);
assign 2_n1645 = 2_n1446;
assign 2_n829 = 2_n1721 | 2_n381;
assign 2_n75 = ~2_n11;
assign 2_n170 = 2_n1033 | 2_n822;
assign 2_n503 = 2_n1510 | 2_n1232;
assign 2_n1140 = 2_n155 & 2_n803;
assign 2_n1360 = ~2_n643;
assign 2_n1231 = 2_n1470;
assign 2_n63 = ~2_n1565;
assign 2_n728 = ~2_n308;
assign 2_n864 = ~2_n991;
assign 2_n1695 = ~(2_n257 | 2_n1626);
assign 2_n1167 = ~(2_n1132 | 2_n544);
assign 2_n522 = 2_n1402 | 2_n649;
assign 2_n1022 = 2_n1347 | 2_n1081;
assign 2_n485 = ~(2_n1248 | 2_n862);
assign 2_n67 = 2_n1717 | 2_n369;
assign 2_n872 = 2_n691 & 2_n901;
assign 2_n514 = ~(2_n1226 | 2_n1344);
assign 2_n933 = ~(2_n572 | 2_n519);
assign 2_n1541 = ~(2_n721 | 2_n21);
endmodule
