module top(in1, in2, in3, out1);
  input [3:0] in1, in2, in3;
  output [3:0] out1;
  wire [3:0] in1, in2, in3;
  wire [3:0] out1;
  wire csa_tree_ADD_TC_OP_groupi_n_0, csa_tree_ADD_TC_OP_groupi_n_1, csa_tree_ADD_TC_OP_groupi_n_2, csa_tree_ADD_TC_OP_groupi_n_3, csa_tree_ADD_TC_OP_groupi_n_4, csa_tree_ADD_TC_OP_groupi_n_5, csa_tree_ADD_TC_OP_groupi_n_6, csa_tree_ADD_TC_OP_groupi_n_7;
  wire csa_tree_ADD_TC_OP_groupi_n_8, csa_tree_ADD_TC_OP_groupi_n_9, csa_tree_ADD_TC_OP_groupi_n_10, csa_tree_ADD_TC_OP_groupi_n_11, csa_tree_ADD_TC_OP_groupi_n_12, csa_tree_ADD_TC_OP_groupi_n_13, csa_tree_ADD_TC_OP_groupi_n_14, csa_tree_ADD_TC_OP_groupi_n_15;
  wire csa_tree_ADD_TC_OP_groupi_n_16, csa_tree_ADD_TC_OP_groupi_n_17, csa_tree_ADD_TC_OP_groupi_n_18, csa_tree_ADD_TC_OP_groupi_n_19, csa_tree_ADD_TC_OP_groupi_n_20, csa_tree_ADD_TC_OP_groupi_n_21, csa_tree_ADD_TC_OP_groupi_n_22, csa_tree_ADD_TC_OP_groupi_n_23;
  wire csa_tree_ADD_TC_OP_groupi_n_24, csa_tree_ADD_TC_OP_groupi_n_25, csa_tree_ADD_TC_OP_groupi_n_26, csa_tree_ADD_TC_OP_groupi_n_27, csa_tree_ADD_TC_OP_groupi_n_28, csa_tree_ADD_TC_OP_groupi_n_29, csa_tree_ADD_TC_OP_groupi_n_30, csa_tree_ADD_TC_OP_groupi_n_31;
  wire csa_tree_ADD_TC_OP_groupi_n_32, csa_tree_ADD_TC_OP_groupi_n_33, csa_tree_ADD_TC_OP_groupi_n_34, csa_tree_ADD_TC_OP_groupi_n_35, csa_tree_ADD_TC_OP_groupi_n_36, csa_tree_ADD_TC_OP_groupi_n_37, csa_tree_ADD_TC_OP_groupi_n_39, csa_tree_ADD_TC_OP_groupi_n_40;
  wire csa_tree_ADD_TC_OP_groupi_n_41, csa_tree_ADD_TC_OP_groupi_n_42, csa_tree_ADD_TC_OP_groupi_n_43, csa_tree_ADD_TC_OP_groupi_n_44, csa_tree_ADD_TC_OP_groupi_n_45, csa_tree_ADD_TC_OP_groupi_n_46, csa_tree_ADD_TC_OP_groupi_n_47, csa_tree_ADD_TC_OP_groupi_n_48;
  wire csa_tree_ADD_TC_OP_groupi_n_49, csa_tree_ADD_TC_OP_groupi_n_50, csa_tree_ADD_TC_OP_groupi_n_51, csa_tree_ADD_TC_OP_groupi_n_53, csa_tree_ADD_TC_OP_groupi_n_54, csa_tree_ADD_TC_OP_groupi_n_55;
  xnor csa_tree_ADD_TC_OP_groupi_g168__2398(out1[3] ,csa_tree_ADD_TC_OP_groupi_n_54 ,csa_tree_ADD_TC_OP_groupi_n_55);
  xnor csa_tree_ADD_TC_OP_groupi_g169__5107(out1[2] ,csa_tree_ADD_TC_OP_groupi_n_48 ,csa_tree_ADD_TC_OP_groupi_n_0);
  xnor csa_tree_ADD_TC_OP_groupi_g170__6260(csa_tree_ADD_TC_OP_groupi_n_55 ,csa_tree_ADD_TC_OP_groupi_n_46 ,csa_tree_ADD_TC_OP_groupi_n_51);
  nor csa_tree_ADD_TC_OP_groupi_g171__4319(csa_tree_ADD_TC_OP_groupi_n_54 ,csa_tree_ADD_TC_OP_groupi_n_50 ,csa_tree_ADD_TC_OP_groupi_n_53);
  nor csa_tree_ADD_TC_OP_groupi_g172__8428(csa_tree_ADD_TC_OP_groupi_n_53 ,csa_tree_ADD_TC_OP_groupi_n_48 ,csa_tree_ADD_TC_OP_groupi_n_49);
  xnor csa_tree_ADD_TC_OP_groupi_g174__5526(out1[1] ,csa_tree_ADD_TC_OP_groupi_n_31 ,csa_tree_ADD_TC_OP_groupi_n_45);
  xnor csa_tree_ADD_TC_OP_groupi_g175__6783(csa_tree_ADD_TC_OP_groupi_n_51 ,csa_tree_ADD_TC_OP_groupi_n_42 ,csa_tree_ADD_TC_OP_groupi_n_43);
  and csa_tree_ADD_TC_OP_groupi_g176__3680(csa_tree_ADD_TC_OP_groupi_n_50 ,csa_tree_ADD_TC_OP_groupi_n_30 ,csa_tree_ADD_TC_OP_groupi_n_44);
  nor csa_tree_ADD_TC_OP_groupi_g177__1617(csa_tree_ADD_TC_OP_groupi_n_49 ,csa_tree_ADD_TC_OP_groupi_n_30 ,csa_tree_ADD_TC_OP_groupi_n_44);
  and csa_tree_ADD_TC_OP_groupi_g178__2802(csa_tree_ADD_TC_OP_groupi_n_48 ,csa_tree_ADD_TC_OP_groupi_n_39 ,csa_tree_ADD_TC_OP_groupi_n_47);
  or csa_tree_ADD_TC_OP_groupi_g179__1705(csa_tree_ADD_TC_OP_groupi_n_47 ,csa_tree_ADD_TC_OP_groupi_n_31 ,csa_tree_ADD_TC_OP_groupi_n_41);
  nor csa_tree_ADD_TC_OP_groupi_g180__5122(csa_tree_ADD_TC_OP_groupi_n_46 ,csa_tree_ADD_TC_OP_groupi_n_28 ,csa_tree_ADD_TC_OP_groupi_n_40);
  xnor csa_tree_ADD_TC_OP_groupi_g181__8246(csa_tree_ADD_TC_OP_groupi_n_45 ,csa_tree_ADD_TC_OP_groupi_n_21 ,csa_tree_ADD_TC_OP_groupi_n_36);
  xnor csa_tree_ADD_TC_OP_groupi_g182__7098(csa_tree_ADD_TC_OP_groupi_n_44 ,csa_tree_ADD_TC_OP_groupi_n_37 ,csa_tree_ADD_TC_OP_groupi_n_33);
  xnor csa_tree_ADD_TC_OP_groupi_g183__6131(csa_tree_ADD_TC_OP_groupi_n_43 ,csa_tree_ADD_TC_OP_groupi_n_22 ,csa_tree_ADD_TC_OP_groupi_n_34);
  xnor csa_tree_ADD_TC_OP_groupi_g184__1881(csa_tree_ADD_TC_OP_groupi_n_42 ,csa_tree_ADD_TC_OP_groupi_n_29 ,csa_tree_ADD_TC_OP_groupi_n_32);
  nor csa_tree_ADD_TC_OP_groupi_g185__5115(csa_tree_ADD_TC_OP_groupi_n_41 ,csa_tree_ADD_TC_OP_groupi_n_20 ,csa_tree_ADD_TC_OP_groupi_n_36);
  and csa_tree_ADD_TC_OP_groupi_g186__7482(csa_tree_ADD_TC_OP_groupi_n_40 ,csa_tree_ADD_TC_OP_groupi_n_27 ,csa_tree_ADD_TC_OP_groupi_n_37);
  or csa_tree_ADD_TC_OP_groupi_g187__4733(csa_tree_ADD_TC_OP_groupi_n_39 ,csa_tree_ADD_TC_OP_groupi_n_21 ,csa_tree_ADD_TC_OP_groupi_n_35);
  xnor csa_tree_ADD_TC_OP_groupi_g188__6161(out1[0] ,csa_tree_ADD_TC_OP_groupi_n_16 ,in3[0]);
  xnor csa_tree_ADD_TC_OP_groupi_g189__9315(csa_tree_ADD_TC_OP_groupi_n_37 ,csa_tree_ADD_TC_OP_groupi_n_23 ,in3[2]);
  not csa_tree_ADD_TC_OP_groupi_g190(csa_tree_ADD_TC_OP_groupi_n_35 ,csa_tree_ADD_TC_OP_groupi_n_36);
  xnor csa_tree_ADD_TC_OP_groupi_g191__9945(csa_tree_ADD_TC_OP_groupi_n_36 ,csa_tree_ADD_TC_OP_groupi_n_25 ,in3[1]);
  xnor csa_tree_ADD_TC_OP_groupi_g192__2883(csa_tree_ADD_TC_OP_groupi_n_34 ,csa_tree_ADD_TC_OP_groupi_n_17 ,csa_tree_ADD_TC_OP_groupi_n_24);
  xnor csa_tree_ADD_TC_OP_groupi_g193__2346(csa_tree_ADD_TC_OP_groupi_n_33 ,csa_tree_ADD_TC_OP_groupi_n_15 ,csa_tree_ADD_TC_OP_groupi_n_19);
  xnor csa_tree_ADD_TC_OP_groupi_g194__1666(csa_tree_ADD_TC_OP_groupi_n_32 ,csa_tree_ADD_TC_OP_groupi_n_13 ,in3[3]);
  or csa_tree_ADD_TC_OP_groupi_g195__7410(csa_tree_ADD_TC_OP_groupi_n_31 ,csa_tree_ADD_TC_OP_groupi_n_10 ,csa_tree_ADD_TC_OP_groupi_n_16);
  and csa_tree_ADD_TC_OP_groupi_g197__6417(csa_tree_ADD_TC_OP_groupi_n_30 ,in3[1] ,csa_tree_ADD_TC_OP_groupi_n_26);
  or csa_tree_ADD_TC_OP_groupi_g198__5477(csa_tree_ADD_TC_OP_groupi_n_29 ,csa_tree_ADD_TC_OP_groupi_n_6 ,csa_tree_ADD_TC_OP_groupi_n_23);
  nor csa_tree_ADD_TC_OP_groupi_g199__2398(csa_tree_ADD_TC_OP_groupi_n_28 ,csa_tree_ADD_TC_OP_groupi_n_15 ,csa_tree_ADD_TC_OP_groupi_n_19);
  or csa_tree_ADD_TC_OP_groupi_g200__5107(csa_tree_ADD_TC_OP_groupi_n_27 ,csa_tree_ADD_TC_OP_groupi_n_14 ,csa_tree_ADD_TC_OP_groupi_n_18);
  not csa_tree_ADD_TC_OP_groupi_g201(csa_tree_ADD_TC_OP_groupi_n_26 ,csa_tree_ADD_TC_OP_groupi_n_25);
  or csa_tree_ADD_TC_OP_groupi_g202__6260(csa_tree_ADD_TC_OP_groupi_n_25 ,csa_tree_ADD_TC_OP_groupi_n_9 ,csa_tree_ADD_TC_OP_groupi_n_3);
  or csa_tree_ADD_TC_OP_groupi_g203__4319(csa_tree_ADD_TC_OP_groupi_n_24 ,csa_tree_ADD_TC_OP_groupi_n_8 ,csa_tree_ADD_TC_OP_groupi_n_5);
  or csa_tree_ADD_TC_OP_groupi_g204__8428(csa_tree_ADD_TC_OP_groupi_n_23 ,csa_tree_ADD_TC_OP_groupi_n_8 ,csa_tree_ADD_TC_OP_groupi_n_3);
  or csa_tree_ADD_TC_OP_groupi_g205__5526(csa_tree_ADD_TC_OP_groupi_n_22 ,csa_tree_ADD_TC_OP_groupi_n_9 ,csa_tree_ADD_TC_OP_groupi_n_7);
  not csa_tree_ADD_TC_OP_groupi_g206(csa_tree_ADD_TC_OP_groupi_n_20 ,csa_tree_ADD_TC_OP_groupi_n_21);
  or csa_tree_ADD_TC_OP_groupi_g207__6783(csa_tree_ADD_TC_OP_groupi_n_21 ,csa_tree_ADD_TC_OP_groupi_n_4 ,csa_tree_ADD_TC_OP_groupi_n_5);
  not csa_tree_ADD_TC_OP_groupi_g208(csa_tree_ADD_TC_OP_groupi_n_19 ,csa_tree_ADD_TC_OP_groupi_n_18);
  and csa_tree_ADD_TC_OP_groupi_g209__3680(csa_tree_ADD_TC_OP_groupi_n_18 ,in1[1] ,in2[1]);
  or csa_tree_ADD_TC_OP_groupi_g210__1617(csa_tree_ADD_TC_OP_groupi_n_17 ,csa_tree_ADD_TC_OP_groupi_n_4 ,csa_tree_ADD_TC_OP_groupi_n_12);
  or csa_tree_ADD_TC_OP_groupi_g211__2802(csa_tree_ADD_TC_OP_groupi_n_16 ,csa_tree_ADD_TC_OP_groupi_n_4 ,csa_tree_ADD_TC_OP_groupi_n_2);
  not csa_tree_ADD_TC_OP_groupi_g212(csa_tree_ADD_TC_OP_groupi_n_15 ,csa_tree_ADD_TC_OP_groupi_n_14);
  and csa_tree_ADD_TC_OP_groupi_g213__1705(csa_tree_ADD_TC_OP_groupi_n_14 ,in1[0] ,in2[2]);
  or csa_tree_ADD_TC_OP_groupi_g214__5122(csa_tree_ADD_TC_OP_groupi_n_13 ,csa_tree_ADD_TC_OP_groupi_n_11 ,csa_tree_ADD_TC_OP_groupi_n_2);
  not csa_tree_ADD_TC_OP_groupi_g215(csa_tree_ADD_TC_OP_groupi_n_12 ,in2[3]);
  not csa_tree_ADD_TC_OP_groupi_g216(csa_tree_ADD_TC_OP_groupi_n_11 ,in1[3]);
  not csa_tree_ADD_TC_OP_groupi_g217(csa_tree_ADD_TC_OP_groupi_n_10 ,in3[0]);
  not csa_tree_ADD_TC_OP_groupi_g218(csa_tree_ADD_TC_OP_groupi_n_9 ,in1[1]);
  not csa_tree_ADD_TC_OP_groupi_g219(csa_tree_ADD_TC_OP_groupi_n_8 ,in1[2]);
  not csa_tree_ADD_TC_OP_groupi_g220(csa_tree_ADD_TC_OP_groupi_n_7 ,in2[2]);
  not csa_tree_ADD_TC_OP_groupi_g221(csa_tree_ADD_TC_OP_groupi_n_6 ,in3[2]);
  not csa_tree_ADD_TC_OP_groupi_g222(csa_tree_ADD_TC_OP_groupi_n_5 ,in2[1]);
  not csa_tree_ADD_TC_OP_groupi_g223(csa_tree_ADD_TC_OP_groupi_n_4 ,in1[0]);
  not csa_tree_ADD_TC_OP_groupi_g224(csa_tree_ADD_TC_OP_groupi_n_3 ,in2[0]);
  not csa_tree_ADD_TC_OP_groupi_drc_bufs225(csa_tree_ADD_TC_OP_groupi_n_2 ,csa_tree_ADD_TC_OP_groupi_n_1);
  not csa_tree_ADD_TC_OP_groupi_drc_bufs226(csa_tree_ADD_TC_OP_groupi_n_1 ,csa_tree_ADD_TC_OP_groupi_n_3);
  xor csa_tree_ADD_TC_OP_groupi_g2__8246(csa_tree_ADD_TC_OP_groupi_n_0 ,csa_tree_ADD_TC_OP_groupi_n_30 ,csa_tree_ADD_TC_OP_groupi_n_44);
endmodule
