module top( 1_n5 , 1_n16 , 1_n23 , 1_n24 , 1_n31 , 1_n38 , 1_n41 , 1_n44 , 1_n46 , 1_n53 , 1_n55 , 1_n57 , 1_n62 , 1_n63 , 1_n68 , 1_n71 , 1_n72 , 1_n78 , 1_n79 , 1_n84 , 1_n92 , 1_n96 , 1_n98 , 1_n101 , 1_n106 , 1_n107 , 1_n120 , 1_n123 , 1_n126 , 1_n136 , 1_n142 , 1_n144 , 1_n145 , 1_n153 , 1_n165 , 1_n177 , 1_n182 , 1_n216 , 1_n220 );
    input 1_n16 , 1_n23 , 1_n24 , 1_n31 , 1_n38 , 1_n41 , 1_n44 , 1_n46 , 1_n53 , 1_n55 , 1_n57 , 1_n62 , 1_n68 , 1_n71 , 1_n72 , 1_n79 , 1_n84 , 1_n92 , 1_n96 , 1_n98 , 1_n101 , 1_n106 , 1_n107 , 1_n120 , 1_n123 , 1_n136 , 1_n145 , 1_n165 , 1_n177 , 1_n182 , 1_n216 , 1_n220 ;
    output 1_n5 , 1_n63 , 1_n78 , 1_n126 , 1_n142 , 1_n144 , 1_n153 ;
    wire 1_n0 , 1_n1 , 1_n2 , 1_n3 , 1_n4 , 1_n6 , 1_n7 , 1_n8 , 1_n9 , 1_n10 , 1_n11 , 1_n12 , 1_n13 , 1_n14 , 1_n15 , 1_n17 , 1_n18 , 1_n19 , 1_n20 , 1_n21 , 1_n22 , 1_n25 , 1_n26 , 1_n27 , 1_n28 , 1_n29 , 1_n30 , 1_n32 , 1_n33 , 1_n34 , 1_n35 , 1_n36 , 1_n37 , 1_n39 , 1_n40 , 1_n42 , 1_n43 , 1_n45 , 1_n47 , 1_n48 , 1_n49 , 1_n50 , 1_n51 , 1_n52 , 1_n54 , 1_n56 , 1_n58 , 1_n59 , 1_n60 , 1_n61 , 1_n64 , 1_n65 , 1_n66 , 1_n67 , 1_n69 , 1_n70 , 1_n73 , 1_n74 , 1_n75 , 1_n76 , 1_n77 , 1_n80 , 1_n81 , 1_n82 , 1_n83 , 1_n85 , 1_n86 , 1_n87 , 1_n88 , 1_n89 , 1_n90 , 1_n91 , 1_n93 , 1_n94 , 1_n95 , 1_n97 , 1_n99 , 1_n100 , 1_n102 , 1_n103 , 1_n104 , 1_n105 , 1_n108 , 1_n109 , 1_n110 , 1_n111 , 1_n112 , 1_n113 , 1_n114 , 1_n115 , 1_n116 , 1_n117 , 1_n118 , 1_n119 , 1_n121 , 1_n122 , 1_n124 , 1_n125 , 1_n127 , 1_n128 , 1_n129 , 1_n130 , 1_n131 , 1_n132 , 1_n133 , 1_n134 , 1_n135 , 1_n137 , 1_n138 , 1_n139 , 1_n140 , 1_n141 , 1_n143 , 1_n146 , 1_n147 , 1_n148 , 1_n149 , 1_n150 , 1_n151 , 1_n152 , 1_n154 , 1_n155 , 1_n156 , 1_n157 , 1_n158 , 1_n159 , 1_n160 , 1_n161 , 1_n162 , 1_n163 , 1_n164 , 1_n166 , 1_n167 , 1_n168 , 1_n169 , 1_n170 , 1_n171 , 1_n172 , 1_n173 , 1_n174 , 1_n175 , 1_n176 , 1_n178 , 1_n179 , 1_n180 , 1_n181 , 1_n183 , 1_n184 , 1_n185 , 1_n186 , 1_n187 , 1_n188 , 1_n189 , 1_n190 , 1_n191 , 1_n192 , 1_n193 , 1_n194 , 1_n195 , 1_n196 , 1_n197 , 1_n198 , 1_n199 , 1_n200 , 1_n201 , 1_n202 , 1_n203 , 1_n204 , 1_n205 , 1_n206 , 1_n207 , 1_n208 , 1_n209 , 1_n210 , 1_n211 , 1_n212 , 1_n213 , 1_n214 , 1_n215 , 1_n217 , 1_n218 , 1_n219 , 1_n221 , 1_n222 , 1_n223 , 1_n224 , 1_n225 , 1_n226 , 1_n227 , 1_n228 , 1_n229 , 1_n230 ;
assign 1_n17 = ~1_n38;
assign 1_n211 = 1_n18 & 1_n116;
assign 1_n193 = ~1_n195;
assign 1_n81 = 1_n118 & 1_n84;
assign 1_n75 = 1_n173 | 1_n113;
assign 1_n180 = 1_n132 & 1_n55;
assign 1_n89 = 1_n125 & 1_n136;
assign 1_n103 = 1_n164 | 1_n131;
assign 1_n127 = 1_n226 & 1_n176;
assign 1_n155 = ~(1_n198 | 1_n179);
assign 1_n18 = ~1_n195;
assign 1_n21 = 1_n180 & 1_n59;
assign 1_n42 = 1_n121 & 1_n170;
assign 1_n209 = 1_n159 & 1_n98;
assign 1_n28 = ~(1_n107 | 1_n70);
assign 1_n135 = 1_n139 & 1_n96;
assign 1_n100 = 1_n209 | 1_n1;
assign 1_n172 = 1_n8 | 1_n230;
assign 1_n78 = 1_n97 | 1_n115;
assign 1_n186 = 1_n229 | 1_n86;
assign 1_n111 = 1_n28 & 1_n68;
assign 1_n88 = ~1_n37;
assign 1_n95 = ~1_n129;
assign 1_n199 = 1_n193 & 1_n71;
assign 1_n2 = ~(1_n190 | 1_n118);
assign 1_n47 = ~1_n61;
assign 1_n179 = 1_n199 | 1_n81;
assign 1_n200 = ~(1_n58 | 1_n194);
assign 1_n205 = 1_n155 & 1_n38;
assign 1_n26 = ~(1_n75 | 1_n115);
assign 1_n105 = ~1_n170;
assign 1_n152 = 1_n153 & 1_n120;
assign 1_n131 = 1_n88 & 1_n31;
assign 1_n201 = ~1_n212;
assign 1_n80 = 1_n227 & 1_n53;
assign 1_n217 = ~1_n67;
assign 1_n51 = 1_n41 | 1_n7;
assign 1_n109 = 1_n218 & 1_n10;
assign 1_n11 = ~(1_n33 | 1_n64);
assign 1_n215 = 1_n80 & 1_n50;
assign 1_n52 = ~1_n106;
assign 1_n159 = ~1_n47;
assign 1_n114 = ~(1_n157 | 1_n125);
assign 1_n110 = ~(1_n79 | 1_n82);
assign 1_n83 = 1_n95 & 1_n79;
assign 1_n133 = 1_n171 | 1_n2;
assign 1_n162 = 1_n66 & 1_n9;
assign 1_n112 = ~1_n182;
assign 1_n138 = ~(1_n89 | 1_n102);
assign 1_n174 = ~1_n217;
assign 1_n39 = 1_n50 | 1_n204;
assign 1_n99 = 1_n0 & 1_n35;
assign 1_n116 = 1_n71 | 1_n17;
assign 1_n50 = 1_n25 & 1_n53;
assign 1_n70 = 1_n5 & 1_n206;
assign 1_n194 = 1_n138 & 1_n53;
assign 1_n160 = 1_n6 & 1_n11;
assign 1_n82 = 1_n159 & 1_n163;
assign 1_n212 = 1_n223 & 1_n51;
assign 1_n161 = 1_n193 & 1_n165;
assign 1_n183 = 1_n171 & 1_n162;
assign 1_n6 = ~(1_n181 | 1_n196);
assign 1_n158 = 1_n80 | 1_n137;
assign 1_n91 = 1_n29 & 1_n48;
assign 1_n29 = 1_n210 & 1_n38;
assign 1_n204 = 1_n29 | 1_n221;
assign 1_n102 = 1_n166 | 1_n60;
assign 1_n35 = 1_n169 | 1_n180;
assign 1_n169 = 1_n168 & 1_n182;
assign 1_n32 = 1_n147 | 1_n191;
assign 1_n25 = ~(1_n136 | 1_n54);
assign 1_n33 = 1_n119 | 1_n85;
assign 1_n154 = 1_n141 & 1_n51;
assign 1_n73 = 1_n46 | 1_n112;
assign 1_n139 = ~(1_n62 | 1_n186);
assign 1_n227 = ~(1_n177 | 1_n54);
assign 1_n143 = 1_n172 | 1_n78;
assign 1_n184 = ~(1_n31 | 1_n128);
assign 1_n141 = 1_n44 | 1_n77;
assign 1_n59 = 1_n110 & 1_n55;
assign 1_n27 = 1_n213 & 1_n230;
assign 1_n178 = 1_n137 & 1_n111;
assign 1_n124 = ~1_n145;
assign 1_n22 = 1_n111 | 1_n108;
assign 1_n148 = 1_n52 | 1_n76;
assign 1_n86 = 1_n153 & 1_n32;
assign 1_n45 = ~1_n195;
assign 1_n153 = ~1_n49;
assign 1_n214 = ~1_n75;
assign 1_n173 = ~1_n68;
assign 1_n66 = ~1_n190;
assign 1_n74 = 1_n169 & 1_n189;
assign 1_n9 = ~1_n92;
assign 1_n134 = 1_n83 | 1_n222;
assign 1_n208 = 1_n34 & 1_n36;
assign 1_n7 = ~1_n84;
assign 1_n163 = 1_n165 | 1_n56;
assign 1_n170 = 1_n147 | 1_n104;
assign 1_n30 = ~(1_n182 | 1_n143);
assign 1_n54 = 1_n45 & 1_n141;
assign 1_n128 = 1_n90 & 1_n10;
assign 1_n130 = ~1_n103;
assign 1_n157 = ~(1_n48 | 1_n34);
assign 1_n225 = ~1_n13;
assign 1_n5 = ~1_n192;
assign 1_n15 = ~(1_n185 | 1_n140);
assign 1_n34 = 1_n184 & 1_n84;
assign 1_n12 = ~1_n101;
assign 1_n48 = 1_n228 & 1_n7;
assign 1_n10 = ~1_n185;
assign 1_n140 = 1_n195 & 1_n84;
assign 1_n171 = 1_n66 & 1_n24;
assign 1_n206 = 1_n57 | 1_n173;
assign 1_n226 = 1_n20 & 1_n116;
assign 1_n4 = 1_n87 & 1_n73;
assign 1_n122 = ~1_n211;
assign 1_n63 = 1_n149 & 1_n103;
assign 1_n13 = ~1_n40;
assign 1_n20 = 1_n154 & 1_n73;
assign 1_n207 = 1_n91 | 1_n208;
assign 1_n164 = 1_n15 | 1_n152;
assign 1_n166 = 1_n45 & 1_n44;
assign 1_n228 = 1_n122 & 1_n38;
assign 1_n67 = ~1_n203;
assign 1_n121 = ~(1_n200 | 1_n26);
assign 1_n0 = 1_n203;
assign 1_n65 = ~(1_n189 | 1_n39);
assign 1_n40 = ~1_n76;
assign 1_n189 = 1_n175 & 1_n182;
assign 1_n132 = ~(1_n16 | 1_n82);
assign 1_n168 = ~(1_n220 | 1_n4);
assign 1_n175 = ~(1_n123 | 1_n4);
assign 1_n156 = ~(1_n216 | 1_n70);
assign 1_n119 = 1_n215 | 1_n178;
assign 1_n94 = 1_n127 & 1_n163;
assign 1_n56 = ~1_n55;
assign 1_n60 = 1_n225 & 1_n177;
assign 1_n187 = 1_n201 & 1_n52;
assign 1_n149 = 1_n3 | 1_n42;
assign 1_n76 = 1_n160 & 1_n219;
assign 1_n142 = ~1_n13;
assign 1_n198 = 1_n146 & 1_n23;
assign 1_n19 = 1_n146 & 1_n72;
assign 1_n3 = 1_n148 & 1_n201;
assign 1_n185 = 1_n12 & 1_n84;
assign 1_n144 = ~(1_n205 | 1_n30);
assign 1_n167 = 1_n74 | 1_n21;
assign 1_n117 = 1_n18 & 1_n57;
assign 1_n181 = 1_n167 | 1_n99;
assign 1_n190 = 1_n124 | 1_n87;
assign 1_n230 = 1_n194 | 1_n214;
assign 1_n210 = ~(1_n23 | 1_n211);
assign 1_n191 = 1_n72 | 1_n229;
assign 1_n150 = 1_n88 & 1_n216;
assign 1_n8 = ~1_n58;
assign 1_n113 = 1_n224 | 1_n93;
assign 1_n126 = ~(1_n97 | 1_n27);
assign 1_n36 = 1_n43 & 1_n84;
assign 1_n64 = 1_n207 | 1_n114;
assign 1_n176 = 1_n98 | 1_n147;
assign 1_n196 = 1_n183 | 1_n135;
assign 1_n129 = ~1_n67;
assign 1_n43 = ~(1_n120 | 1_n128);
assign 1_n218 = 1_n94 & 1_n206;
assign 1_n213 = ~1_n115;
assign 1_n137 = 1_n156 & 1_n68;
assign 1_n104 = 1_n19 | 1_n100;
assign 1_n146 = ~1_n129;
assign 1_n61 = ~1_n109;
assign 1_n49 = ~1_n174;
assign 1_n97 = 1_n130 | 1_n3;
assign 1_n188 = ~1_n32;
assign 1_n203 = 1_n65 & 1_n212;
assign 1_n197 = 1_n59 | 1_n22;
assign 1_n223 = ~1_n140;
assign 1_n202 = 1_n133 & 1_n151;
assign 1_n221 = 1_n36 | 1_n197;
assign 1_n90 = ~1_n47;
assign 1_n195 = 1_n109;
assign 1_n229 = 1_n90 & 1_n176;
assign 1_n85 = 1_n0 & 1_n158;
assign 1_n147 = ~1_n96;
assign 1_n69 = 1_n225 & 1_n16;
assign 1_n87 = ~1_n192;
assign 1_n224 = 1_n95 & 1_n107;
assign 1_n151 = 1_n9 | 1_n0;
assign 1_n125 = ~1_n217;
assign 1_n108 = 1_n188 | 1_n162;
assign 1_n93 = 1_n117 | 1_n150;
assign 1_n115 = 1_n202 | 1_n105;
assign 1_n77 = ~1_n53;
assign 1_n1 = 1_n142 & 1_n62;
assign 1_n58 = 1_n56 | 1_n134;
assign 1_n192 = ~1_n61;
assign 1_n37 = ~1_n40;
assign 1_n222 = 1_n161 | 1_n69;
assign 1_n219 = ~(1_n187 | 1_n14);
assign 1_n118 = ~1_n37;
assign 1_n14 = 1_n0 & 1_n171;
endmodule
