module top( 2_n0 , 2_n2 , 2_n17 , 2_n18 , 2_n23 , 2_n24 , 2_n26 , 2_n27 , 2_n29 , 2_n37 , 2_n43 , 2_n58 , 2_n59 , 2_n61 , 2_n66 , 2_n70 , 2_n73 , 2_n75 , 2_n80 , 2_n81 , 2_n84 , 2_n86 , 2_n88 , 2_n89 , 2_n90 , 2_n91 , 2_n94 , 2_n98 , 2_n104 , 2_n107 , 2_n123 , 2_n129 , 2_n130 , 2_n133 , 2_n137 , 2_n145 , 2_n151 , 2_n160 , 2_n164 , 2_n168 , 2_n169 , 2_n174 , 2_n179 , 2_n187 , 2_n194 , 2_n196 , 2_n199 , 2_n210 , 2_n211 , 2_n212 , 2_n213 , 2_n214 , 2_n217 , 2_n221 , 2_n226 , 2_n234 , 2_n237 , 2_n238 , 2_n246 , 2_n249 , 2_n253 , 2_n256 , 2_n260 , 2_n261 , 2_n265 , 2_n272 , 2_n278 , 2_n281 , 2_n286 , 2_n289 , 2_n292 , 2_n304 , 2_n310 );
    input 2_n0 , 2_n2 , 2_n17 , 2_n18 , 2_n23 , 2_n27 , 2_n29 , 2_n37 , 2_n43 , 2_n58 , 2_n59 , 2_n70 , 2_n75 , 2_n84 , 2_n90 , 2_n91 , 2_n107 , 2_n130 , 2_n133 , 2_n137 , 2_n169 , 2_n174 , 2_n179 , 2_n187 , 2_n194 , 2_n196 , 2_n210 , 2_n211 , 2_n214 , 2_n226 , 2_n234 , 2_n237 , 2_n238 , 2_n249 , 2_n256 , 2_n260 , 2_n272 , 2_n278 , 2_n281 , 2_n289 , 2_n292 ;
    output 2_n24 , 2_n26 , 2_n61 , 2_n66 , 2_n73 , 2_n80 , 2_n81 , 2_n86 , 2_n88 , 2_n89 , 2_n94 , 2_n98 , 2_n104 , 2_n123 , 2_n129 , 2_n145 , 2_n151 , 2_n160 , 2_n164 , 2_n168 , 2_n199 , 2_n212 , 2_n213 , 2_n217 , 2_n221 , 2_n246 , 2_n253 , 2_n261 , 2_n265 , 2_n286 , 2_n304 , 2_n310 ;
    wire 2_n1 , 2_n3 , 2_n4 , 2_n5 , 2_n6 , 2_n7 , 2_n8 , 2_n9 , 2_n10 , 2_n11 , 2_n12 , 2_n13 , 2_n14 , 2_n15 , 2_n16 , 2_n19 , 2_n20 , 2_n21 , 2_n22 , 2_n25 , 2_n28 , 2_n30 , 2_n31 , 2_n32 , 2_n33 , 2_n34 , 2_n35 , 2_n36 , 2_n38 , 2_n39 , 2_n40 , 2_n41 , 2_n42 , 2_n44 , 2_n45 , 2_n46 , 2_n47 , 2_n48 , 2_n49 , 2_n50 , 2_n51 , 2_n52 , 2_n53 , 2_n54 , 2_n55 , 2_n56 , 2_n57 , 2_n60 , 2_n62 , 2_n63 , 2_n64 , 2_n65 , 2_n67 , 2_n68 , 2_n69 , 2_n71 , 2_n72 , 2_n74 , 2_n76 , 2_n77 , 2_n78 , 2_n79 , 2_n82 , 2_n83 , 2_n85 , 2_n87 , 2_n92 , 2_n93 , 2_n95 , 2_n96 , 2_n97 , 2_n99 , 2_n100 , 2_n101 , 2_n102 , 2_n103 , 2_n105 , 2_n106 , 2_n108 , 2_n109 , 2_n110 , 2_n111 , 2_n112 , 2_n113 , 2_n114 , 2_n115 , 2_n116 , 2_n117 , 2_n118 , 2_n119 , 2_n120 , 2_n121 , 2_n122 , 2_n124 , 2_n125 , 2_n126 , 2_n127 , 2_n128 , 2_n131 , 2_n132 , 2_n134 , 2_n135 , 2_n136 , 2_n138 , 2_n139 , 2_n140 , 2_n141 , 2_n142 , 2_n143 , 2_n144 , 2_n146 , 2_n147 , 2_n148 , 2_n149 , 2_n150 , 2_n152 , 2_n153 , 2_n154 , 2_n155 , 2_n156 , 2_n157 , 2_n158 , 2_n159 , 2_n161 , 2_n162 , 2_n163 , 2_n165 , 2_n166 , 2_n167 , 2_n170 , 2_n171 , 2_n172 , 2_n173 , 2_n175 , 2_n176 , 2_n177 , 2_n178 , 2_n180 , 2_n181 , 2_n182 , 2_n183 , 2_n184 , 2_n185 , 2_n186 , 2_n188 , 2_n189 , 2_n190 , 2_n191 , 2_n192 , 2_n193 , 2_n195 , 2_n197 , 2_n198 , 2_n200 , 2_n201 , 2_n202 , 2_n203 , 2_n204 , 2_n205 , 2_n206 , 2_n207 , 2_n208 , 2_n209 , 2_n215 , 2_n216 , 2_n218 , 2_n219 , 2_n220 , 2_n222 , 2_n223 , 2_n224 , 2_n225 , 2_n227 , 2_n228 , 2_n229 , 2_n230 , 2_n231 , 2_n232 , 2_n233 , 2_n235 , 2_n236 , 2_n239 , 2_n240 , 2_n241 , 2_n242 , 2_n243 , 2_n244 , 2_n245 , 2_n247 , 2_n248 , 2_n250 , 2_n251 , 2_n252 , 2_n254 , 2_n255 , 2_n257 , 2_n258 , 2_n259 , 2_n262 , 2_n263 , 2_n264 , 2_n266 , 2_n267 , 2_n268 , 2_n269 , 2_n270 , 2_n271 , 2_n273 , 2_n274 , 2_n275 , 2_n276 , 2_n277 , 2_n279 , 2_n280 , 2_n282 , 2_n283 , 2_n284 , 2_n285 , 2_n287 , 2_n288 , 2_n290 , 2_n291 , 2_n293 , 2_n294 , 2_n295 , 2_n296 , 2_n297 , 2_n298 , 2_n299 , 2_n300 , 2_n301 , 2_n302 , 2_n303 , 2_n305 , 2_n306 , 2_n307 , 2_n308 , 2_n309 , 2_n311 ;
assign 2_n163 = ~(2_n174 ^ 2_n169);
assign 2_n129 = ~(2_n153 ^ 2_n210);
assign 2_n53 = 2_n205 | 2_n155;
assign 2_n28 = 2_n279 | 2_n298;
assign 2_n14 = ~(2_n124 ^ 2_n126);
assign 2_n66 = ~(2_n30 ^ 2_n29);
assign 2_n143 = 2_n140 | 2_n216;
assign 2_n38 = 2_n301 | 2_n72;
assign 2_n262 = ~(2_n238 ^ 2_n29);
assign 2_n259 = ~2_n180;
assign 2_n251 = 2_n96 | 2_n51;
assign 2_n45 = ~(2_n43 ^ 2_n214);
assign 2_n60 = ~(2_n8 ^ 2_n114);
assign 2_n19 = 2_n273 | 2_n297;
assign 2_n34 = ~(2_n70 ^ 2_n174);
assign 2_n209 = 2_n140 | 2_n175;
assign 2_n275 = 2_n53 | 2_n276;
assign 2_n239 = ~(2_n14 ^ 2_n288);
assign 2_n308 = ~(2_n70 ^ 2_n2);
assign 2_n255 = 2_n251 | 2_n172;
assign 2_n166 = 2_n305 | 2_n181;
assign 2_n198 = 2_n252 | 2_n173;
assign 2_n86 = ~(2_n200 ^ 2_n196);
assign 2_n223 = 2_n250 | 2_n46;
assign 2_n5 = 2_n62 | 2_n85;
assign 2_n161 = 2_n178 | 2_n64;
assign 2_n204 = ~2_n58;
assign 2_n1 = ~(2_n189 ^ 2_n296);
assign 2_n301 = ~2_n119;
assign 2_n9 = 2_n283 | 2_n291;
assign 2_n304 = ~(2_n224 ^ 2_n214);
assign 2_n208 = ~(2_n225 ^ 2_n83);
assign 2_n21 = 2_n110 | 2_n82;
assign 2_n57 = ~(2_n135 ^ 2_n197);
assign 2_n296 = ~(2_n179 ^ 2_n0);
assign 2_n203 = 2_n171 | 2_n103;
assign 2_n243 = 2_n205 | 2_n155;
assign 2_n303 = ~(2_n237 ^ 2_n210);
assign 2_n191 = ~(2_n278 ^ 2_n272);
assign 2_n171 = ~2_n226;
assign 2_n233 = 2_n149 ^ 2_n309;
assign 2_n140 = ~2_n78;
assign 2_n279 = ~2_n119;
assign 2_n63 = ~(2_n130 ^ 2_n107);
assign 2_n220 = 2_n235 | 2_n274;
assign 2_n65 = 2_n128 | 2_n68;
assign 2_n103 = ~2_n281;
assign 2_n150 = 2_n60;
assign 2_n149 = ~(2_n32 ^ 2_n141);
assign 2_n270 = 2_n112 | 2_n190;
assign 2_n41 = 2_n155 | 2_n230;
assign 2_n248 = ~(2_n17 ^ 2_n75);
assign 2_n267 = 2_n56 | 2_n273;
assign 2_n294 = 2_n204 | 2_n103;
assign 2_n85 = 2_n152 | 2_n276;
assign 2_n62 = 2_n140 | 2_n216;
assign 2_n274 = 2_n95 | 2_n76;
assign 2_n311 = ~(2_n130 ^ 2_n256);
assign 2_n114 = ~(2_n294 ^ 2_n87);
assign 2_n222 = ~(2_n77 ^ 2_n191);
assign 2_n69 = 2_n156 | 2_n76;
assign 2_n263 = 2_n162 | 2_n51;
assign 2_n221 = ~(2_n219 ^ 2_n179);
assign 2_n36 = 2_n258 | 2_n33;
assign 2_n254 = ~(2_n23 ^ 2_n249);
assign 2_n306 = ~(2_n290 ^ 2_n10);
assign 2_n297 = ~2_n279;
assign 2_n286 = ~(2_n49 ^ 2_n238);
assign 2_n141 = ~(2_n256 ^ 2_n289);
assign 2_n67 = 2_n167 | 2_n159;
assign 2_n104 = ~(2_n142 ^ 2_n289);
assign 2_n26 = ~(2_n115 ^ 2_n169);
assign 2_n92 = 2_n127 | 2_n113;
assign 2_n244 = 2_n243 | 2_n232;
assign 2_n269 = 2_n56 | 2_n72;
assign 2_n142 = 2_n209 | 2_n9;
assign 2_n10 = ~(2_n234 ^ 2_n196);
assign 2_n215 = 2_n15 | 2_n33;
assign 2_n216 = ~2_n134;
assign 2_n154 = 2_n263 | 2_n198;
assign 2_n113 = 2_n183 | 2_n230;
assign 2_n186 = 2_n184 | 2_n103;
assign 2_n68 = 2_n206 | 2_n255;
assign 2_n93 = ~2_n74;
assign 2_n52 = ~(2_n238 ^ 2_n17);
assign 2_n49 = 2_n28 | 2_n159;
assign 2_n188 = 2_n162 | 2_n106;
assign 2_n250 = 2_n301 | 2_n298;
assign 2_n115 = 2_n105 | 2_n64;
assign 2_n240 = ~(2_n229 ^ 2_n303);
assign 2_n33 = 2_n267 | 2_n173;
assign 2_n197 = ~(2_n285 ^ 2_n42);
assign 2_n87 = ~(2_n278 ^ 2_n234);
assign 2_n88 = ~(2_n299 ^ 2_n107);
assign 2_n117 = ~(2_n194 ^ 2_n27);
assign 2_n227 = ~(2_n242 ^ 2_n240);
assign 2_n89 = ~(2_n271 ^ 2_n43);
assign 2_n290 = ~(2_n260 ^ 2_n27);
assign 2_n202 = 2_n101 | 2_n9;
assign 2_n280 = 2_n177 | 2_n297;
assign 2_n155 = ~2_n60;
assign 2_n46 = 2_n7 | 2_n181;
assign 2_n258 = 2_n301 | 2_n138;
assign 2_n126 = ~(2_n249 ^ 2_n214);
assign 2_n190 = ~2_n100;
assign 2_n158 = 2_n112 | 2_n190;
assign 2_n177 = ~2_n233;
assign 2_n30 = 2_n13 | 2_n274;
assign 2_n175 = ~2_n134;
assign 2_n232 = 2_n301 | 2_n25;
assign 2_n252 = 2_n96 | 2_n93;
assign 2_n156 = 2_n96 | 2_n93;
assign 2_n160 = ~(2_n16 ^ 2_n70);
assign 2_n167 = 2_n177 | 2_n51;
assign 2_n159 = 2_n266 | 2_n92;
assign 2_n152 = 2_n150 | 2_n230;
assign 2_n172 = 2_n298 | 2_n93;
assign 2_n287 = ~(2_n83 ^ 2_n222);
assign 2_n101 = 2_n112 | 2_n231;
assign 2_n235 = 2_n177 | 2_n259;
assign 2_n94 = ~(2_n223 ^ 2_n137);
assign 2_n310 = ~(2_n65 ^ 2_n237);
assign 2_n25 = 2_n138 | 2_n106;
assign 2_n299 = 2_n144 | 2_n244;
assign 2_n31 = 2_n38 | 2_n69;
assign 2_n81 = ~(2_n132 ^ 2_n90);
assign 2_n39 = 2_n301 | 2_n298;
assign 2_n72 = ~2_n50;
assign 2_n134 = ~2_n71;
assign 2_n246 = ~(2_n277 ^ 2_n249);
assign 2_n245 = ~(2_n136 ^ 2_n108);
assign 2_n11 = 2_n39 | 2_n201;
assign 2_n183 = ~2_n110;
assign 2_n298 = ~2_n50;
assign 2_n162 = ~2_n233;
assign 2_n213 = ~(2_n220 ^ 2_n75);
assign 2_n305 = 2_n56 | 2_n273;
assign 2_n82 = ~2_n241;
assign 2_n164 = ~(2_n161 ^ 2_n2);
assign 2_n131 = ~(2_n102 ^ 2_n120);
assign 2_n122 = ~(2_n208 ^ 2_n45);
assign 2_n132 = 2_n158 | 2_n85;
assign 2_n293 = 2_n157 | 2_n103;
assign 2_n95 = 2_n56 | 2_n273;
assign 2_n205 = 2_n57;
assign 2_n257 = ~2_n91;
assign 2_n148 = 2_n112 | 2_n41;
assign 2_n120 = ~(2_n187 ^ 2_n211);
assign 2_n283 = 2_n205 | 2_n155;
assign 2_n99 = 2_n307 | 2_n147;
assign 2_n284 = 2_n55 | 2_n46;
assign 2_n6 = ~(2_n306 ^ 2_n222);
assign 2_n73 = ~(2_n284 ^ 2_n260);
assign 2_n178 = 2_n112 | 2_n231;
assign 2_n78 = 2_n131 ^ 2_n44;
assign 2_n173 = 2_n140 | 2_n3;
assign 2_n125 = ~(2_n287 ^ 2_n63);
assign 2_n136 = ~(2_n163 ^ 2_n195);
assign 2_n195 = ~(2_n210 ^ 2_n59);
assign 2_n105 = 2_n110 | 2_n175;
assign 2_n7 = 2_n96 | 2_n93;
assign 2_n199 = ~(2_n36 ^ 2_n187);
assign 2_n277 = 2_n21 | 2_n147;
assign 2_n118 = ~(2_n293 ^ 2_n34);
assign 2_n145 = ~(2_n11 ^ 2_n278);
assign 2_n218 = ~(2_n97 ^ 2_n268);
assign 2_n291 = 2_n297 | 2_n188;
assign 2_n32 = ~(2_n225 ^ 2_n306);
assign 2_n121 = ~(2_n137 ^ 2_n260);
assign 2_n48 = 2_n279 | 2_n138;
assign 2_n153 = 2_n143 | 2_n68;
assign 2_n80 = ~(2_n116 ^ 2_n174);
assign 2_n229 = 2_n257 | 2_n103;
assign 2_n61 = ~(2_n67 ^ 2_n17);
assign 2_n54 = ~(2_n2 ^ 2_n169);
assign 2_n200 = 2_n236 | 2_n69;
assign 2_n96 = 2_n227;
assign 2_n193 = 2_n150 | 2_n230;
assign 2_n176 = 2_n280 | 2_n166;
assign 2_n185 = 2_n162 | 2_n297;
assign 2_n128 = 2_n112 | 2_n183;
assign 2_n100 = ~2_n78;
assign 2_n24 = ~(2_n5 ^ 2_n59);
assign 2_n77 = ~(2_n137 ^ 2_n194);
assign 2_n207 = ~(2_n29 ^ 2_n75);
assign 2_n276 = 2_n269 | 2_n19;
assign 2_n139 = 2_n96 | 2_n93;
assign 2_n212 = ~(2_n99 ^ 2_n23);
assign 2_n217 = ~(2_n202 ^ 2_n256);
assign 2_n302 = 2_n185 | 2_n201;
assign 2_n146 = ~(2_n179 ^ 2_n187);
assign 2_n268 = ~(2_n90 ^ 2_n59);
assign 2_n206 = 2_n150 | 2_n230;
assign 2_n230 = ~2_n57;
assign 2_n12 = 2_n241 | 2_n183;
assign 2_n3 = 2_n82 | 2_n41;
assign 2_n109 = 2_n47 | 2_n232;
assign 2_n236 = 2_n162 | 2_n259;
assign 2_n135 = ~(2_n239 ^ 2_n207);
assign 2_n47 = 2_n150 | 2_n230;
assign 2_n64 = 2_n193 | 2_n291;
assign 2_n4 = 2_n35 | 2_n198;
assign 2_n56 = 2_n74;
assign 2_n264 = 2_n12 | 2_n244;
assign 2_n74 = ~(2_n122 ^ 2_n218);
assign 2_n168 = ~(2_n264 ^ 2_n130);
assign 2_n112 = ~2_n71;
assign 2_n189 = ~(2_n288 ^ 2_n108);
assign 2_n102 = ~(2_n14 ^ 2_n136);
assign 2_n8 = ~(2_n245 ^ 2_n52);
assign 2_n71 = 2_n1 ^ 2_n182;
assign 2_n300 = 2_n155 | 2_n82;
assign 2_n242 = ~(2_n6 ^ 2_n254);
assign 2_n79 = ~2_n84;
assign 2_n123 = ~(2_n215 ^ 2_n211);
assign 2_n151 = ~(2_n302 ^ 2_n234);
assign 2_n127 = 2_n150 | 2_n175;
assign 2_n266 = 2_n56 | 2_n273;
assign 2_n50 = ~2_n233;
assign 2_n295 = ~(2_n23 ^ 2_n43);
assign 2_n22 = 2_n247 | 2_n103;
assign 2_n16 = 2_n270 | 2_n109;
assign 2_n42 = ~(2_n272 ^ 2_n196);
assign 2_n116 = 2_n20 | 2_n109;
assign 2_n147 = 2_n165 | 2_n255;
assign 2_n181 = 2_n183 | 2_n148;
assign 2_n170 = 2_n241 | 2_n231;
assign 2_n165 = 2_n205 | 2_n155;
assign 2_n225 = ~(2_n111 ^ 2_n248);
assign 2_n241 = ~2_n71;
assign 2_n265 = ~(2_n4 ^ 2_n194);
assign 2_n35 = 2_n301 | 2_n138;
assign 2_n157 = ~2_n37;
assign 2_n192 = ~2_n292;
assign 2_n285 = 2_n79 | 2_n103;
assign 2_n184 = ~2_n18;
assign 2_n55 = 2_n162 | 2_n259;
assign 2_n309 = ~(2_n186 ^ 2_n54);
assign 2_n119 = 2_n125 ^ 2_n118;
assign 2_n97 = 2_n192 | 2_n103;
assign 2_n13 = 2_n279 | 2_n72;
assign 2_n106 = 2_n273 | 2_n93;
assign 2_n273 = ~2_n227;
assign 2_n307 = 2_n241 | 2_n190;
assign 2_n231 = ~2_n100;
assign 2_n51 = ~2_n180;
assign 2_n76 = 2_n282 | 2_n300;
assign 2_n224 = 2_n228 | 2_n275;
assign 2_n247 = ~2_n133;
assign 2_n83 = ~(2_n146 ^ 2_n262);
assign 2_n201 = 2_n139 | 2_n92;
assign 2_n228 = 2_n140 | 2_n82;
assign 2_n182 = ~(2_n203 ^ 2_n121);
assign 2_n124 = ~(2_n107 ^ 2_n289);
assign 2_n15 = 2_n162 | 2_n51;
assign 2_n219 = 2_n48 | 2_n166;
assign 2_n253 = ~(2_n31 ^ 2_n272);
assign 2_n180 = ~2_n119;
assign 2_n138 = ~2_n177;
assign 2_n108 = ~(2_n308 ^ 2_n40);
assign 2_n110 = ~2_n78;
assign 2_n271 = 2_n170 | 2_n275;
assign 2_n20 = 2_n140 | 2_n175;
assign 2_n98 = ~(2_n154 ^ 2_n27);
assign 2_n44 = ~(2_n22 ^ 2_n117);
assign 2_n111 = ~(2_n0 ^ 2_n211);
assign 2_n282 = 2_n205 | 2_n231;
assign 2_n288 = ~(2_n311 ^ 2_n295);
assign 2_n40 = ~(2_n237 ^ 2_n90);
assign 2_n261 = ~(2_n176 ^ 2_n0);
assign 2_n144 = 2_n110 | 2_n216;
endmodule
