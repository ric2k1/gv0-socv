module top( n1 , n4 , n5 , n6 , n11 , n16 , n19 , n24 , n35 , n36 , n39 , n44 , n45 , n46 , n48 , n49 );
    input n1 , n4 , n5 , n11 , n19 , n24 , n35 , n39 , n45 , n46 , n48 , n49 ;
    output n6 , n16 , n36 , n44 ;
    wire n0 , n2 , n3 , n7 , n8 , n9 , n10 , n12 , n13 , n14 , n15 , n17 , n18 , n20 , n21 , n22 , n23 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n37 , n38 , n40 , n41 , n42 , n43 , n47 ;
assign n38 = ~n11;
assign n43 = ~(n47 ^ n49);
assign n10 = ~n30;
assign n6 = ~(n7 ^ n23);
assign n34 = n26 | n8;
assign n15 = ~(n20 | n7);
assign n27 = ~(n35 ^ n48);
assign n41 = ~(n5 ^ n4);
assign n14 = ~(n18 ^ n3);
assign n23 = ~(n14 ^ n19);
assign n31 = ~(n24 ^ n39);
assign n13 = ~(n35 & n48);
assign n25 = ~(n0 ^ n11);
assign n28 = ~(n22 | n18);
assign n36 = ~(n31 ^ n46);
assign n18 = n32 & n13;
assign n8 = ~n39;
assign n30 = n21 & n46;
assign n22 = ~(n45 | n1);
assign n0 = ~(n34 ^ n27);
assign n9 = ~(n35 | n48);
assign n3 = ~(n45 ^ n1);
assign n12 = n38 | n10;
assign n7 = n2 & n12;
assign n20 = n14 & n29;
assign n21 = ~n31;
assign n17 = n40 | n15;
assign n2 = n0 | n37;
assign n32 = n9 | n34;
assign n42 = ~(n41 ^ n17);
assign n16 = ~(n43 ^ n42);
assign n33 = n1 & n45;
assign n37 = ~(n11 | n30);
assign n44 = ~(n10 ^ n25);
assign n26 = ~n24;
assign n29 = ~n19;
assign n40 = ~(n29 | n14);
assign n47 = n33 | n28;
endmodule
