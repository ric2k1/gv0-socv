module top( n9 , n22 , n103 , n124 , n134 , n201 , n211 , n287 , n353 , 
n358 , n370 , n389 , n396 , n401 , n411 , n443 , n460 , n469 , n497 , 
n499 , n510 , n537 , n573 , n603 , n728 , n758 , n761 , n762 , n767 , 
n772 , n777 , n800 , n817 , n831 , n834 , n846 , n854 , n922 , n927 , 
n937 , n951 , n985 , n1007 , n1084 , n1097 , n1112 , n1165 , n1181 , n1198 , 
n1231 , n1302 , n1307 , n1364 , n1392 , n1401 , n1487 , n1561 , n1636 , n1650 , 
n1709 , n1724 , n1757 , n1806 , n1860 , n1912 , n1916 , n1937 , n1982 , n2057 , 
n2061 , n2068 , n2174 , n2190 , n2235 , n2252 , n2295 , n2339 , n2341 , n2458 , 
n2482 , n2498 , n2549 , n2590 , n2592 , n2666 , n2709 , n2737 , n2758 , n2771 , 
n2777 , n2805 , n2882 , n2904 , n2934 , n3006 , n3076 , n3085 , n3112 , n3130 , 
n3178 , n3262 , n3311 , n3323 , n3362 , n3409 , n3591 , n3641 , n3669 , n3677 , 
n3748 , n3769 , n3790 , n3815 , n3832 , n3946 , n4006 , n4059 , n4075 , n4114 , 
n4122 , n4141 , n4202 , n4330 , n4335 , n4357 , n4382 , n4419 , n4452 , n4470 , 
n4553 , n4743 , n4748 , n4777 , n4824 , n4862 , n4864 , n4964 , n4998 , n5003 , 
n5031 , n5060 , n5065 , n5167 , n5189 , n5214 , n5320 , n5356 , n5364 , n5427 , 
n5470 , n5536 , n5548 , n5549 , n5557 , n5568 , n5586 , n5609 , n5671 , n5684 , 
n5715 , n5729 , n5758 , n5801 , n5882 , n5884 , n5920 , n5962 , n5969 , n6019 , 
n6023 , n6085 , n6103 , n6109 , n6149 , n6168 , n6297 , n6301 , n6333 , n6392 , 
n6409 , n6434 , n6586 , n6655 , n6668 , n6683 , n6818 , n6826 , n6843 , n6862 , 
n6937 , n7034 , n7061 , n7111 , n7113 , n7132 , n7161 , n7241 , n7374 , n7411 , 
n7529 , n7553 , n7582 , n7659 , n7687 , n7715 , n7720 , n7729 , n7755 , n7772 , 
n7790 , n7812 , n7858 , n7860 , n7968 , n7974 , n8139 , n8163 , n8172 , n8183 , 
n8219 , n8228 , n8230 , n8233 , n8265 , n8290 , n8308 , n8332 , n8336 , n8466 , 
n8468 , n8506 , n8516 , n8522 , n8701 , n8716 , n8768 , n8820 , n8859 , n8860 , 
n8940 , n9041 , n9093 , n9100 , n9187 , n9216 , n9300 , n9329 , n9353 , n9475 , 
n9528 , n9531 , n9570 , n9591 , n9620 , n9669 , n9732 , n9747 , n9846 , n9866 , 
n9872 , n9887 , n9906 , n9915 , n10063 , n10101 , n10113 , n10122 , n10142 , n10162 , 
n10168 , n10243 , n10408 , n10416 , n10451 , n10453 , n10522 , n10524 , n10560 , n10594 , 
n10606 , n10628 , n10642 , n10657 , n10736 , n10770 , n10797 , n10805 , n10866 , n10874 , 
n10908 , n11030 , n11057 , n11058 , n11061 , n11077 , n11109 , n11111 , n11140 , n11147 , 
n11180 , n11222 , n11236 , n11252 , n11264 , n11324 , n11350 , n11396 , n11411 , n11429 , 
n11484 , n11488 , n11537 , n11574 , n11634 , n11665 , n11667 , n11732 , n11734 , n11778 , 
n11792 , n11835 , n11879 , n11882 , n11891 , n11895 , n12003 , n12059 , n12065 , n12067 , 
n12187 , n12263 , n12284 , n12289 , n12306 , n12334 , n12348 , n12352 , n12372 , n12406 , 
n12408 , n12463 , n12482 , n12503 , n12515 , n12579 , n12592 , n12605 , n12616 , n12651 , 
n12693 , n12750 , n12839 , n12853 , n12912 , n12965 , n12968 , n13002 , n13035 , n13058 , 
n13060 , n13201 );
    input n9 , n22 , n103 , n124 , n287 , n353 , n389 , n401 , n411 , 
n443 , n469 , n497 , n499 , n510 , n603 , n761 , n767 , n772 , n817 , 
n834 , n854 , n937 , n951 , n1007 , n1084 , n1165 , n1198 , n1231 , n1302 , 
n1307 , n1364 , n1392 , n1636 , n1650 , n1709 , n1724 , n1757 , n1912 , n1916 , 
n1982 , n2057 , n2068 , n2174 , n2252 , n2295 , n2339 , n2341 , n2458 , n2482 , 
n2498 , n2590 , n2592 , n2666 , n2737 , n2758 , n2771 , n2777 , n2882 , n3006 , 
n3076 , n3085 , n3112 , n3130 , n3178 , n3311 , n3409 , n3591 , n3641 , n3669 , 
n3677 , n3769 , n3815 , n3832 , n4006 , n4075 , n4114 , n4122 , n4141 , n4330 , 
n4335 , n4357 , n4382 , n4419 , n4452 , n4470 , n4743 , n4748 , n4862 , n4964 , 
n4998 , n5031 , n5065 , n5167 , n5189 , n5214 , n5320 , n5356 , n5427 , n5470 , 
n5536 , n5548 , n5568 , n5586 , n5671 , n5684 , n5715 , n5729 , n5758 , n5801 , 
n5884 , n5920 , n5962 , n5969 , n6023 , n6085 , n6149 , n6168 , n6333 , n6392 , 
n6409 , n6655 , n6668 , n6818 , n6826 , n6843 , n6937 , n7061 , n7113 , n7161 , 
n7374 , n7411 , n7529 , n7659 , n7715 , n7720 , n7729 , n7772 , n7812 , n7974 , 
n8139 , n8163 , n8183 , n8228 , n8230 , n8233 , n8290 , n8308 , n8332 , n8466 , 
n8468 , n8506 , n8522 , n8716 , n8768 , n8820 , n8859 , n8860 , n8940 , n9041 , 
n9093 , n9187 , n9216 , n9300 , n9353 , n9475 , n9528 , n9531 , n9570 , n9591 , 
n9620 , n9669 , n9732 , n9747 , n9846 , n9887 , n9906 , n9915 , n10063 , n10113 , 
n10122 , n10142 , n10162 , n10168 , n10408 , n10416 , n10451 , n10522 , n10560 , n10594 , 
n10606 , n10642 , n10657 , n10770 , n10805 , n10866 , n10874 , n10908 , n11030 , n11058 , 
n11061 , n11109 , n11111 , n11180 , n11222 , n11236 , n11324 , n11350 , n11396 , n11411 , 
n11429 , n11488 , n11537 , n11574 , n11634 , n11665 , n11734 , n11835 , n11891 , n12003 , 
n12065 , n12263 , n12284 , n12289 , n12306 , n12348 , n12352 , n12372 , n12408 , n12482 , 
n12579 , n12592 , n12605 , n12651 , n12693 , n12750 , n12853 , n12912 , n12965 , n13058 , 
n13060 , n13201 ;
    output n134 , n201 , n211 , n358 , n370 , n396 , n460 , n537 , n573 , 
n728 , n758 , n762 , n777 , n800 , n831 , n846 , n922 , n927 , n985 , 
n1097 , n1112 , n1181 , n1401 , n1487 , n1561 , n1806 , n1860 , n1937 , n2061 , 
n2190 , n2235 , n2549 , n2709 , n2805 , n2904 , n2934 , n3262 , n3323 , n3362 , 
n3748 , n3790 , n3946 , n4059 , n4202 , n4553 , n4777 , n4824 , n4864 , n5003 , 
n5060 , n5364 , n5549 , n5557 , n5609 , n5882 , n6019 , n6103 , n6109 , n6297 , 
n6301 , n6434 , n6586 , n6683 , n6862 , n7034 , n7111 , n7132 , n7241 , n7553 , 
n7582 , n7687 , n7755 , n7790 , n7858 , n7860 , n7968 , n8172 , n8219 , n8265 , 
n8336 , n8516 , n8701 , n9100 , n9329 , n9866 , n9872 , n10101 , n10243 , n10453 , 
n10524 , n10628 , n10736 , n10797 , n11057 , n11077 , n11140 , n11147 , n11252 , n11264 , 
n11484 , n11667 , n11732 , n11778 , n11792 , n11879 , n11882 , n11895 , n12059 , n12067 , 
n12187 , n12334 , n12406 , n12463 , n12503 , n12515 , n12616 , n12839 , n12968 , n13002 , 
n13035 ;
    wire n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , 
n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , 
n20 , n21 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , 
n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , 
n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , 
n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , 
n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , 
n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , 
n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , 
n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , 
n101 , n102 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , 
n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , 
n122 , n123 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , 
n133 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , 
n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , 
n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , 
n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , 
n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , 
n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , 
n194 , n195 , n196 , n197 , n198 , n199 , n200 , n202 , n203 , n204 , 
n205 , n206 , n207 , n208 , n209 , n210 , n212 , n213 , n214 , n215 , 
n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , 
n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , 
n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , 
n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , 
n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , 
n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , 
n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , 
n286 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , 
n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , 
n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , 
n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , 
n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , 
n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , 
n347 , n348 , n349 , n350 , n351 , n352 , n354 , n355 , n356 , n357 , 
n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , 
n369 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , 
n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n390 , 
n391 , n392 , n393 , n394 , n395 , n397 , n398 , n399 , n400 , n402 , 
n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n412 , n413 , 
n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , 
n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , 
n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n444 , 
n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , 
n455 , n456 , n457 , n458 , n459 , n461 , n462 , n463 , n464 , n465 , 
n466 , n467 , n468 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , 
n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , 
n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , 
n498 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , 
n509 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , 
n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , 
n530 , n531 , n532 , n533 , n534 , n535 , n536 , n538 , n539 , n540 , 
n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , 
n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , 
n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , 
n571 , n572 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , 
n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , 
n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , 
n602 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , 
n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , 
n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , 
n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , 
n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , 
n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , 
n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , 
n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , 
n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , 
n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , 
n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , 
n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , 
n723 , n724 , n725 , n726 , n727 , n729 , n730 , n731 , n732 , n733 , 
n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , 
n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , 
n754 , n755 , n756 , n757 , n759 , n760 , n763 , n764 , n765 , n766 , 
n768 , n769 , n770 , n771 , n773 , n774 , n775 , n776 , n778 , n779 , 
n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , 
n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , 
n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , 
n811 , n812 , n813 , n814 , n815 , n816 , n818 , n819 , n820 , n821 , 
n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n832 , 
n833 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , 
n844 , n845 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n855 , 
n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , 
n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , 
n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , 
n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , 
n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , 
n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , 
n916 , n917 , n918 , n919 , n920 , n921 , n923 , n924 , n925 , n926 , 
n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n938 , 
n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , 
n949 , n950 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , 
n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , 
n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , 
n980 , n981 , n982 , n983 , n984 , n986 , n987 , n988 , n989 , n990 , 
n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , 
n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1008 , n1009 , n1010 , n1011 , 
n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , 
n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , 
n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , 
n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , 
n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , 
n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , 
n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , 
n1082 , n1083 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , 
n1093 , n1094 , n1095 , n1096 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , 
n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1113 , n1114 , 
n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , 
n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , 
n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , 
n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , 
n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , 
n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , 
n1176 , n1177 , n1178 , n1179 , n1180 , n1182 , n1183 , n1184 , n1185 , n1186 , 
n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , 
n1197 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , 
n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , 
n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , 
n1228 , n1229 , n1230 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , 
n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , 
n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , 
n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , 
n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , 
n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , 
n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , 
n1299 , n1300 , n1301 , n1303 , n1304 , n1305 , n1306 , n1308 , n1309 , n1310 , 
n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , 
n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , 
n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , 
n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , 
n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , 
n1361 , n1362 , n1363 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , 
n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , 
n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , 
n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1402 , n1403 , 
n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , 
n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , 
n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , 
n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , 
n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , 
n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , 
n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , 
n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , 
n1484 , n1485 , n1486 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , 
n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , 
n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , 
n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , 
n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , 
n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , 
n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , 
n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1562 , n1563 , n1564 , n1565 , 
n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , 
n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , 
n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , 
n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , 
n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , 
n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , 
n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , 
n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , 
n1647 , n1648 , n1649 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , 
n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , 
n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , 
n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , 
n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , 
n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , 
n1708 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , 
n1719 , n1720 , n1721 , n1722 , n1723 , n1725 , n1726 , n1727 , n1728 , n1729 , 
n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , 
n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , 
n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1758 , n1759 , n1760 , 
n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , 
n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , 
n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , 
n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , 
n1801 , n1802 , n1803 , n1804 , n1805 , n1807 , n1808 , n1809 , n1810 , n1811 , 
n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , 
n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , 
n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , 
n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , 
n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1861 , n1862 , 
n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , 
n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , 
n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , 
n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , 
n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1913 , 
n1914 , n1915 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , 
n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , 
n1935 , n1936 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , 
n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , 
n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , 
n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , 
n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1983 , n1984 , n1985 , n1986 , 
n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , 
n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , 
n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , 
n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , 
n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , 
n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , 
n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , 
n2058 , n2059 , n2060 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2069 , 
n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , 
n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , 
n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , 
n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , 
n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , 
n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , 
n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , 
n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , 
n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , 
n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , 
n2170 , n2171 , n2172 , n2173 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , 
n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2191 , 
n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , 
n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , 
n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , 
n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , 
n2232 , n2233 , n2234 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , 
n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2253 , 
n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , 
n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , 
n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , 
n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , 
n2294 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , 
n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , 
n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , 
n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , 
n2335 , n2336 , n2337 , n2338 , n2340 , n2342 , n2343 , n2344 , n2345 , n2346 , 
n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , 
n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , 
n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , 
n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , 
n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , 
n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , 
n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , 
n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , 
n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , 
n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , 
n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , 
n2457 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , 
n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , 
n2478 , n2479 , n2480 , n2481 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , 
n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2499 , 
n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , 
n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , 
n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , 
n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , 
n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2550 , 
n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , 
n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , 
n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , 
n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2591 , 
n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , 
n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , 
n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , 
n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , 
n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , 
n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , 
n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , 
n2663 , n2664 , n2665 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , 
n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , 
n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , 
n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , 
n2704 , n2705 , n2706 , n2707 , n2708 , n2710 , n2711 , n2712 , n2713 , n2714 , 
n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , 
n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , 
n2735 , n2736 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , 
n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , 
n2756 , n2757 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , 
n2767 , n2768 , n2769 , n2770 , n2772 , n2773 , n2774 , n2775 , n2776 , n2778 , 
n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , 
n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , 
n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2806 , n2807 , n2808 , n2809 , 
n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , 
n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , 
n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , 
n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , 
n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , 
n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , 
n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , 
n2880 , n2881 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , 
n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , 
n2901 , n2902 , n2903 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , 
n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , 
n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , 
n2932 , n2933 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , 
n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , 
n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , 
n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , 
n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , 
n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , 
n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , 
n3003 , n3004 , n3005 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , 
n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , 
n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , 
n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , 
n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , 
n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , 
n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , 
n3074 , n3075 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , 
n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , 
n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , 
n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3113 , n3114 , n3115 , n3116 , 
n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , 
n3127 , n3128 , n3129 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , 
n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , 
n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , 
n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , 
n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , 
n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , 
n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , 
n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , 
n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , 
n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , 
n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , 
n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , 
n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , 
n3259 , n3260 , n3261 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , 
n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , 
n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , 
n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , 
n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , 
n3310 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , 
n3321 , n3322 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , 
n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , 
n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , 
n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , 
n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , 
n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , 
n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , 
n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , 
n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3410 , n3411 , n3412 , n3413 , 
n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , 
n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , 
n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , 
n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , 
n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , 
n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , 
n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , 
n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , 
n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , 
n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , 
n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , 
n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , 
n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , 
n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , 
n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , 
n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , 
n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , 
n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3592 , n3593 , n3594 , 
n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , 
n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , 
n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , 
n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , 
n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3642 , n3643 , n3644 , n3645 , 
n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , 
n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , 
n3666 , n3667 , n3668 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , 
n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , 
n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , 
n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , 
n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , 
n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , 
n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , 
n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , 
n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , 
n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , 
n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , 
n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , 
n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , 
n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , 
n3811 , n3812 , n3813 , n3814 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , 
n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , 
n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , 
n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , 
n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , 
n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , 
n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , 
n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , 
n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , 
n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , 
n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , 
n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , 
n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , 
n3943 , n3944 , n3945 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , 
n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , 
n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , 
n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , 
n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , 
n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , 
n4004 , n4005 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , 
n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , 
n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , 
n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , 
n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , 
n4055 , n4056 , n4057 , n4058 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , 
n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4076 , 
n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , 
n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , 
n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , 
n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4115 , n4116 , n4117 , 
n4118 , n4119 , n4120 , n4121 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , 
n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , 
n4139 , n4140 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , 
n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , 
n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , 
n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , 
n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , 
n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , 
n4200 , n4201 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , 
n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , 
n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , 
n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , 
n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , 
n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , 
n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , 
n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , 
n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , 
n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , 
n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , 
n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , 
n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4331 , 
n4332 , n4333 , n4334 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , 
n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , 
n4353 , n4354 , n4355 , n4356 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , 
n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , 
n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4383 , n4384 , 
n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , 
n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , 
n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , 
n4415 , n4416 , n4417 , n4418 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , 
n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , 
n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , 
n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4453 , n4454 , n4455 , n4456 , 
n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , 
n4467 , n4468 , n4469 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , 
n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , 
n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , 
n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , 
n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , 
n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , 
n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , 
n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , 
n4548 , n4549 , n4550 , n4551 , n4552 , n4554 , n4555 , n4556 , n4557 , n4558 , 
n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , 
n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , 
n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , 
n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , 
n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , 
n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , 
n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , 
n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , 
n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , 
n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , 
n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , 
n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , 
n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , 
n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , 
n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , 
n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , 
n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , 
n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , 
n4739 , n4740 , n4741 , n4742 , n4744 , n4745 , n4746 , n4747 , n4749 , n4750 , 
n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , 
n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , 
n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4778 , n4779 , n4780 , n4781 , 
n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , 
n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , 
n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , 
n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , 
n4822 , n4823 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , 
n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , 
n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , 
n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4863 , 
n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , 
n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , 
n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , 
n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , 
n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , 
n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , 
n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , 
n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , 
n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , 
n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4965 , 
n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , 
n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , 
n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , 
n4996 , n4997 , n4999 , n5000 , n5001 , n5002 , n5004 , n5005 , n5006 , n5007 , 
n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , 
n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , 
n5028 , n5029 , n5030 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , 
n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , 
n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , 
n5059 , n5061 , n5062 , n5063 , n5064 , n5066 , n5067 , n5068 , n5069 , n5070 , 
n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , 
n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , 
n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , 
n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , 
n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , 
n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , 
n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , 
n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , 
n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , 
n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5168 , n5169 , n5170 , n5171 , 
n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , 
n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5190 , n5191 , n5192 , 
n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , 
n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , 
n5213 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , 
n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , 
n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , 
n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , 
n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , 
n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , 
n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , 
n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , 
n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , 
n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , 
n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5321 , n5322 , n5323 , n5324 , 
n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , 
n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , 
n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , 
n5355 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5365 , n5366 , 
n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , 
n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , 
n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , 
n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , 
n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , 
n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , 
n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , 
n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , 
n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , 
n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , 
n5468 , n5469 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , 
n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , 
n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , 
n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , 
n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , 
n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , 
n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5537 , n5538 , n5539 , 
n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5550 , n5551 , 
n5552 , n5553 , n5554 , n5555 , n5556 , n5558 , n5559 , n5560 , n5561 , n5562 , 
n5563 , n5564 , n5565 , n5566 , n5567 , n5569 , n5570 , n5571 , n5572 , n5573 , 
n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , 
n5584 , n5585 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , 
n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , 
n5605 , n5606 , n5607 , n5608 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , 
n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , 
n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , 
n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , 
n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , 
n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , 
n5666 , n5667 , n5668 , n5669 , n5670 , n5672 , n5673 , n5674 , n5675 , n5676 , 
n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5685 , n5686 , n5687 , 
n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , 
n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , 
n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5716 , n5717 , n5718 , 
n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , 
n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , 
n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , 
n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5759 , n5760 , 
n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , 
n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , 
n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , 
n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , 
n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , 
n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , 
n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , 
n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , 
n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , 
n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , 
n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , 
n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , 
n5883 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , 
n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , 
n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , 
n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5921 , n5922 , n5923 , n5924 , 
n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , 
n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , 
n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , 
n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5963 , n5964 , n5965 , 
n5966 , n5967 , n5968 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , 
n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , 
n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , 
n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , 
n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , 
n6017 , n6018 , n6020 , n6021 , n6022 , n6024 , n6025 , n6026 , n6027 , n6028 , 
n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , 
n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , 
n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , 
n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , 
n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , 
n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6086 , n6087 , n6088 , n6089 , 
n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , 
n6100 , n6101 , n6102 , n6104 , n6105 , n6106 , n6107 , n6108 , n6110 , n6111 , 
n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , 
n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , 
n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , 
n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6150 , n6151 , n6152 , 
n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , 
n6163 , n6164 , n6165 , n6166 , n6167 , n6169 , n6170 , n6171 , n6172 , n6173 , 
n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , 
n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , 
n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , 
n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , 
n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , 
n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , 
n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , 
n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , 
n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , 
n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , 
n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , 
n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , 
n6294 , n6295 , n6296 , n6298 , n6299 , n6300 , n6302 , n6303 , n6304 , n6305 , 
n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , 
n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , 
n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6334 , n6335 , n6336 , 
n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , 
n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , 
n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , 
n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , 
n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , 
n6387 , n6388 , n6389 , n6390 , n6391 , n6393 , n6394 , n6395 , n6396 , n6397 , 
n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , 
n6408 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , 
n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , 
n6429 , n6430 , n6431 , n6432 , n6433 , n6435 , n6436 , n6437 , n6438 , n6439 , 
n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , 
n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , 
n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , 
n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , 
n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , 
n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , 
n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , 
n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , 
n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , 
n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , 
n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , 
n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , 
n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , 
n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , 
n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6587 , n6588 , n6589 , n6590 , 
n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , 
n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , 
n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , 
n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , 
n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , 
n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , 
n6651 , n6652 , n6653 , n6654 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , 
n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6669 , n6670 , n6671 , n6672 , 
n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , 
n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , 
n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , 
n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , 
n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , 
n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , 
n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , 
n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , 
n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , 
n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , 
n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , 
n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , 
n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , 
n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , 
n6814 , n6815 , n6816 , n6817 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , 
n6825 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , 
n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6844 , n6845 , n6846 , 
n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , 
n6857 , n6858 , n6859 , n6860 , n6861 , n6863 , n6864 , n6865 , n6866 , n6867 , 
n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , 
n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , 
n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , 
n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , 
n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , 
n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , 
n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6938 , 
n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , 
n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , 
n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , 
n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , 
n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , 
n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , 
n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , 
n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , 
n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , 
n7029 , n7030 , n7031 , n7032 , n7033 , n7035 , n7036 , n7037 , n7038 , n7039 , 
n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , 
n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , 
n7060 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , 
n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , 
n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , 
n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , 
n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , 
n7112 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , 
n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7133 , 
n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , 
n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , 
n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7162 , n7163 , n7164 , 
n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , 
n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , 
n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , 
n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , 
n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , 
n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , 
n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , 
n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7242 , n7243 , n7244 , n7245 , 
n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , 
n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , 
n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , 
n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , 
n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , 
n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , 
n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , 
n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , 
n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , 
n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , 
n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , 
n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , 
n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7375 , n7376 , 
n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , 
n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , 
n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , 
n7407 , n7408 , n7409 , n7410 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , 
n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , 
n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , 
n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , 
n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , 
n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , 
n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , 
n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , 
n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , 
n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , 
n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , 
n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , 
n7528 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , 
n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , 
n7549 , n7550 , n7551 , n7552 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , 
n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , 
n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , 
n7580 , n7581 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , 
n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , 
n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , 
n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , 
n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , 
n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , 
n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , 
n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7660 , n7661 , 
n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , 
n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , 
n7682 , n7683 , n7684 , n7685 , n7686 , n7688 , n7689 , n7690 , n7691 , n7692 , 
n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , 
n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , 
n7713 , n7714 , n7716 , n7717 , n7718 , n7719 , n7721 , n7722 , n7723 , n7724 , 
n7725 , n7726 , n7727 , n7728 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , 
n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , 
n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7756 , 
n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , 
n7767 , n7768 , n7769 , n7770 , n7771 , n7773 , n7774 , n7775 , n7776 , n7777 , 
n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , 
n7788 , n7789 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , 
n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , 
n7809 , n7810 , n7811 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , 
n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , 
n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , 
n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , 
n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7859 , n7861 , 
n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , 
n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , 
n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , 
n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , 
n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , 
n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , 
n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , 
n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , 
n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , 
n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , 
n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7969 , n7970 , n7971 , n7972 , 
n7973 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , 
n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , 
n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , 
n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , 
n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , 
n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , 
n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , 
n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , 
n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , 
n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , 
n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , 
n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , 
n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , 
n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , 
n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , 
n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , 
n8134 , n8135 , n8136 , n8137 , n8138 , n8140 , n8141 , n8142 , n8143 , n8144 , 
n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , 
n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8164 , n8165 , 
n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8173 , n8174 , n8175 , n8176 , 
n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8184 , n8185 , n8186 , n8187 , 
n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , 
n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , 
n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , 
n8218 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8229 , 
n8231 , n8232 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , 
n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , 
n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , 
n8262 , n8263 , n8264 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , 
n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , 
n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8291 , n8292 , n8293 , 
n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , 
n8304 , n8305 , n8306 , n8307 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , 
n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , 
n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8333 , n8334 , n8335 , 
n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , 
n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , 
n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , 
n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , 
n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , 
n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , 
n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , 
n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , 
n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , 
n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , 
n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , 
n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , 
n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8467 , 
n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , 
n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , 
n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , 
n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8507 , n8508 , n8509 , 
n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8517 , n8518 , n8519 , n8520 , 
n8521 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , 
n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , 
n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , 
n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , 
n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , 
n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , 
n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , 
n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , 
n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , 
n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , 
n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , 
n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , 
n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , 
n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , 
n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , 
n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , 
n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , 
n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8702 , 
n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , 
n8713 , n8714 , n8715 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , 
n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , 
n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , 
n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , 
n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , 
n8764 , n8765 , n8766 , n8767 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , 
n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , 
n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , 
n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , 
n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , 
n8815 , n8816 , n8817 , n8818 , n8819 , n8821 , n8822 , n8823 , n8824 , n8825 , 
n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , 
n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , 
n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , 
n8856 , n8857 , n8858 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , 
n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , 
n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , 
n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , 
n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , 
n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , 
n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , 
n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , 
n8938 , n8939 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , 
n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , 
n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , 
n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , 
n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , 
n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , 
n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , 
n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , 
n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , 
n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , 
n9039 , n9040 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , 
n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , 
n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , 
n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , 
n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , 
n9090 , n9091 , n9092 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9101 , 
n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , 
n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , 
n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , 
n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , 
n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , 
n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , 
n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , 
n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , 
n9182 , n9183 , n9184 , n9185 , n9186 , n9188 , n9189 , n9190 , n9191 , n9192 , 
n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , 
n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , 
n9213 , n9214 , n9215 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , 
n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , 
n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , 
n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , 
n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , 
n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , 
n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , 
n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , 
n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9301 , n9302 , n9303 , n9304 , 
n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , 
n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , 
n9325 , n9326 , n9327 , n9328 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , 
n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , 
n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9354 , n9355 , n9356 , 
n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , 
n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , 
n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , 
n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , 
n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , 
n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , 
n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , 
n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , 
n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , 
n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , 
n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , 
n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9476 , n9477 , 
n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , 
n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , 
n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , 
n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , 
n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , 
n9529 , n9530 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , 
n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , 
n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , 
n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , 
n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , 
n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , 
n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , 
n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , 
n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9621 , n9622 , 
n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , 
n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , 
n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , 
n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , 
n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9670 , n9671 , n9672 , n9673 , 
n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , 
n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , 
n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , 
n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , 
n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , 
n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9733 , n9734 , 
n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , 
n9745 , n9746 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , 
n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , 
n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , 
n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , 
n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , 
n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , 
n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , 
n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , 
n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , 
n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , 
n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , 
n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9867 , 
n9868 , n9869 , n9870 , n9871 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , 
n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9888 , n9889 , 
n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , 
n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9907 , n9908 , n9909 , n9910 , 
n9911 , n9912 , n9913 , n9914 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , 
n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , 
n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , 
n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , 
n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , 
n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , 
n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , 
n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , 
n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , 
n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , 
n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , 
n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , 
n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , 
n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , 
n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , 
n10062 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , 
n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , 
n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , 
n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10102 , n10103 , 
n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10114 , 
n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10123 , n10124 , n10125 , 
n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , 
n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10143 , n10144 , n10145 , n10146 , 
n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , 
n10157 , n10158 , n10159 , n10160 , n10161 , n10163 , n10164 , n10165 , n10166 , n10167 , 
n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , 
n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , 
n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , 
n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , 
n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , 
n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , 
n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , 
n10239 , n10240 , n10241 , n10242 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , 
n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , 
n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , 
n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , 
n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , 
n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , 
n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , 
n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , 
n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , 
n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , 
n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , 
n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , 
n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , 
n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , 
n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , 
n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , 
n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10409 , n10410 , 
n10411 , n10412 , n10413 , n10414 , n10415 , n10417 , n10418 , n10419 , n10420 , n10421 , 
n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , 
n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , 
n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , n10452 , 
n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , 
n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , 
n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , 
n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , 
n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , 
n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , 
n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10523 , n10525 , 
n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , 
n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , 
n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , 
n10556 , n10557 , n10558 , n10559 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , 
n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , 
n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , 
n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10595 , n10596 , n10597 , 
n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10607 , n10608 , 
n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , 
n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10629 , 
n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , 
n10640 , n10641 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , 
n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10658 , n10659 , n10660 , n10661 , 
n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , 
n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , 
n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , 
n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , 
n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , 
n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , 
n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , 
n10732 , n10733 , n10734 , n10735 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , 
n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , 
n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , 
n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10771 , n10772 , n10773 , 
n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , 
n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , 
n10794 , n10795 , n10796 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , 
n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , 
n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , 
n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , 
n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , 
n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , 
n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , 
n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10875 , n10876 , n10877 , 
n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , 
n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , 
n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , 
n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , 
n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , 
n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , 
n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , 
n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , 
n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , 
n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , 
n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , 
n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , 
n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , 
n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , 
n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , 
n11029 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , 
n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , 
n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11059 , n11060 , n11062 , 
n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , 
n11073 , n11074 , n11075 , n11076 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , 
n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , 
n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , 
n11104 , n11105 , n11106 , n11107 , n11108 , n11110 , n11112 , n11113 , n11114 , n11115 , 
n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , 
n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , 
n11136 , n11137 , n11138 , n11139 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , 
n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , 
n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , 
n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , 
n11178 , n11179 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , 
n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , 
n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , 
n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , 
n11219 , n11220 , n11221 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , 
n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11237 , n11238 , n11239 , n11240 , 
n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , 
n11251 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , 
n11262 , n11263 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , 
n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , 
n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , 
n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , 
n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , 
n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , 
n11323 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , 
n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , 
n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11351 , n11352 , n11353 , n11354 , 
n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , 
n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , 
n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , 
n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , 
n11395 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , 
n11406 , n11407 , n11408 , n11409 , n11410 , n11412 , n11413 , n11414 , n11415 , n11416 , 
n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , 
n11427 , n11428 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , 
n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , 
n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , 
n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , 
n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , 
n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11485 , n11486 , n11487 , n11489 , 
n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , 
n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , 
n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , 
n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , 
n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11538 , n11539 , n11540 , 
n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , 
n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , 
n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , 
n11571 , n11572 , n11573 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , 
n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , 
n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , 
n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , 
n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , 
n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , 
n11632 , n11633 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , 
n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , 
n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , 
n11663 , n11664 , n11666 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , 
n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , 
n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , 
n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , 
n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , 
n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , 
n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11733 , n11735 , n11736 , 
n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , 
n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , 
n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , 
n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , 
n11777 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , 
n11788 , n11789 , n11790 , n11791 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , 
n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , 
n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , 
n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , 
n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11836 , n11837 , n11838 , n11839 , 
n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , 
n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , 
n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , 
n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11880 , 
n11881 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11892 , 
n11893 , n11894 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , 
n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , 
n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , 
n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , 
n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , 
n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , 
n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , 
n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , 
n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , 
n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , 
n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12004 , 
n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , 
n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , 
n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , 
n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , 
n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , 
n12055 , n12056 , n12057 , n12058 , n12060 , n12061 , n12062 , n12063 , n12064 , n12066 , 
n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , 
n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , 
n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , 
n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , 
n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , 
n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , 
n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , 
n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , 
n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , 
n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , 
n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , 
n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12188 , 
n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , 
n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , 
n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , 
n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , 
n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , 
n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , 
n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , 
n12259 , n12260 , n12261 , n12262 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , 
n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , 
n12280 , n12281 , n12282 , n12283 , n12285 , n12286 , n12287 , n12288 , n12290 , n12291 , 
n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , 
n12302 , n12303 , n12304 , n12305 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , 
n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , 
n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , 
n12333 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , 
n12344 , n12345 , n12346 , n12347 , n12349 , n12350 , n12351 , n12353 , n12354 , n12355 , 
n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , 
n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12373 , n12374 , n12375 , n12376 , 
n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , 
n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , 
n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12407 , 
n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , 
n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , 
n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , 
n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , 
n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , 
n12459 , n12460 , n12461 , n12462 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , 
n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , 
n12480 , n12481 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , 
n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , 
n12501 , n12502 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , n12511 , 
n12512 , n12513 , n12514 , n12516 , n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , 
n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , 
n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , 
n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , 
n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , 
n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , 
n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12580 , n12581 , n12582 , n12583 , 
n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , n12591 , n12593 , n12594 , 
n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , 
n12606 , n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , 
n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , 
n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , 
n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , 
n12647 , n12648 , n12649 , n12650 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , 
n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , 
n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , 
n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , 
n12688 , n12689 , n12690 , n12691 , n12692 , n12694 , n12695 , n12696 , n12697 , n12698 , 
n12699 , n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , 
n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , 
n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , 
n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , 
n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , 
n12749 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , 
n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , 
n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , 
n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , 
n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , 
n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , 
n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , 
n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , 
n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12840 , 
n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , 
n12851 , n12852 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , n12861 , 
n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , n12871 , 
n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , n12880 , n12881 , 
n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , n12891 , 
n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , n12901 , 
n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , n12911 , 
n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , 
n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , n12929 , n12930 , n12931 , n12932 , 
n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , n12941 , n12942 , 
n12943 , n12944 , n12945 , n12946 , n12947 , n12948 , n12949 , n12950 , n12951 , n12952 , 
n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , n12960 , n12961 , n12962 , 
n12963 , n12964 , n12966 , n12967 , n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , 
n12975 , n12976 , n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , 
n12985 , n12986 , n12987 , n12988 , n12989 , n12990 , n12991 , n12992 , n12993 , n12994 , 
n12995 , n12996 , n12997 , n12998 , n12999 , n13000 , n13001 , n13003 , n13004 , n13005 , 
n13006 , n13007 , n13008 , n13009 , n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , 
n13016 , n13017 , n13018 , n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , 
n13026 , n13027 , n13028 , n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , n13036 , 
n13037 , n13038 , n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , 
n13047 , n13048 , n13049 , n13050 , n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , 
n13057 , n13059 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , 
n13069 , n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , 
n13079 , n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , 
n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , 
n13099 , n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , 
n13109 , n13110 , n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , n13117 , n13118 , 
n13119 , n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , 
n13129 , n13130 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , 
n13139 , n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , 
n13149 , n13150 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , 
n13159 , n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , 
n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , 
n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , 
n13189 , n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , 
n13199 , n13200 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , 
n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , n13219 , 
n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , 
n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , 
n13240 , n13241 , n13242 , n13243 ;
    and g0 ( n3523 , n7151 , n6767 );
    xnor g1 ( n1818 , n11618 , n10125 );
    or g2 ( n6666 , n1354 , n6635 );
    or g3 ( n13003 , n10781 , n8348 );
    or g4 ( n8017 , n995 , n12970 );
    and g5 ( n9879 , n4074 , n12255 );
    xnor g6 ( n849 , n1713 , n1158 );
    nor g7 ( n837 , n3701 , n2651 );
    xnor g8 ( n3470 , n12726 , n4668 );
    xnor g9 ( n6673 , n2914 , n655 );
    xnor g10 ( n8353 , n3258 , n2954 );
    or g11 ( n1644 , n7660 , n10173 );
    xnor g12 ( n4458 , n11074 , n9291 );
    or g13 ( n4154 , n12552 , n10871 );
    not g14 ( n5448 , n13203 );
    or g15 ( n938 , n2711 , n11144 );
    not g16 ( n9174 , n72 );
    or g17 ( n6954 , n3044 , n11894 );
    xnor g18 ( n224 , n10835 , n2683 );
    not g19 ( n7171 , n2309 );
    nor g20 ( n1343 , n8789 , n7265 );
    not g21 ( n3099 , n5324 );
    not g22 ( n12128 , n5568 );
    nor g23 ( n12514 , n5673 , n13166 );
    or g24 ( n5497 , n10761 , n6732 );
    and g25 ( n6006 , n3747 , n4857 );
    xnor g26 ( n8827 , n6431 , n7145 );
    and g27 ( n9763 , n7126 , n2227 );
    or g28 ( n11908 , n4316 , n2924 );
    xnor g29 ( n2161 , n11270 , n1874 );
    xnor g30 ( n618 , n7815 , n4460 );
    not g31 ( n1422 , n12965 );
    xnor g32 ( n9158 , n601 , n9373 );
    or g33 ( n9135 , n1550 , n2209 );
    and g34 ( n12910 , n1958 , n4654 );
    or g35 ( n13069 , n10439 , n12388 );
    xnor g36 ( n13000 , n4381 , n10298 );
    xnor g37 ( n12582 , n1459 , n1950 );
    xnor g38 ( n1273 , n8182 , n8861 );
    not g39 ( n11174 , n485 );
    not g40 ( n5045 , n5586 );
    or g41 ( n7486 , n6079 , n4448 );
    or g42 ( n9434 , n6006 , n9735 );
    or g43 ( n6268 , n7700 , n1026 );
    or g44 ( n11498 , n6991 , n11644 );
    not g45 ( n1005 , n10373 );
    not g46 ( n10206 , n6964 );
    xnor g47 ( n746 , n4418 , n496 );
    or g48 ( n12707 , n7675 , n1144 );
    or g49 ( n11383 , n5865 , n5242 );
    not g50 ( n12636 , n9701 );
    not g51 ( n6506 , n3311 );
    or g52 ( n5217 , n7939 , n1337 );
    not g53 ( n6028 , n12482 );
    xnor g54 ( n7328 , n6204 , n12282 );
    or g55 ( n3430 , n12568 , n12847 );
    xnor g56 ( n13217 , n8937 , n9105 );
    xnor g57 ( n7035 , n3487 , n1164 );
    or g58 ( n11295 , n10032 , n7254 );
    not g59 ( n734 , n11411 );
    xnor g60 ( n11278 , n9811 , n9427 );
    xnor g61 ( n10946 , n12215 , n3738 );
    xnor g62 ( n610 , n10055 , n774 );
    xnor g63 ( n10496 , n10728 , n13055 );
    xnor g64 ( n12601 , n3959 , n9631 );
    or g65 ( n10620 , n6939 , n9159 );
    not g66 ( n5216 , n1426 );
    xnor g67 ( n3802 , n596 , n1088 );
    or g68 ( n12895 , n13027 , n10662 );
    not g69 ( n11521 , n9732 );
    not g70 ( n4884 , n3670 );
    not g71 ( n9741 , n8078 );
    xor g72 ( n1826 , n6083 , n7616 );
    xnor g73 ( n3658 , n12111 , n4323 );
    and g74 ( n6851 , n11030 , n12289 );
    xnor g75 ( n10227 , n10752 , n594 );
    xor g76 ( n11559 , n6226 , n4888 );
    or g77 ( n127 , n10882 , n11551 );
    or g78 ( n8256 , n7819 , n10043 );
    buf g79 ( n10029 , n8852 );
    not g80 ( n4473 , n2295 );
    not g81 ( n10956 , n5729 );
    not g82 ( n3456 , n11682 );
    not g83 ( n9718 , n6670 );
    or g84 ( n7609 , n8188 , n4490 );
    nor g85 ( n10187 , n330 , n12782 );
    and g86 ( n5538 , n4081 , n9186 );
    xnor g87 ( n1464 , n520 , n7499 );
    xnor g88 ( n9928 , n4616 , n9260 );
    buf g89 ( n1570 , n12471 );
    xnor g90 ( n1525 , n8885 , n10490 );
    and g91 ( n3435 , n3669 , n834 );
    or g92 ( n11902 , n2848 , n12501 );
    or g93 ( n2414 , n4258 , n10106 );
    and g94 ( n252 , n10338 , n6627 );
    or g95 ( n9289 , n1168 , n7723 );
    or g96 ( n12010 , n5480 , n2796 );
    xnor g97 ( n13046 , n6622 , n10271 );
    or g98 ( n12280 , n683 , n9080 );
    or g99 ( n7727 , n7912 , n13118 );
    xnor g100 ( n8096 , n8582 , n10826 );
    or g101 ( n9186 , n5455 , n4724 );
    xnor g102 ( n4933 , n5944 , n5560 );
    xnor g103 ( n7994 , n2528 , n8607 );
    not g104 ( n10128 , n11891 );
    or g105 ( n1597 , n3186 , n3500 );
    nor g106 ( n12870 , n1824 , n10842 );
    and g107 ( n11470 , n1782 , n10313 );
    not g108 ( n5626 , n7556 );
    xnor g109 ( n5131 , n7739 , n3051 );
    and g110 ( n425 , n1907 , n9672 );
    xnor g111 ( n7539 , n9415 , n9935 );
    or g112 ( n3425 , n10761 , n8702 );
    xnor g113 ( n8270 , n465 , n727 );
    and g114 ( n12783 , n7695 , n9404 );
    xnor g115 ( n3269 , n6985 , n12644 );
    and g116 ( n12026 , n3006 , n6149 );
    not g117 ( n12042 , n10925 );
    not g118 ( n9682 , n11324 );
    and g119 ( n10094 , n4795 , n8792 );
    not g120 ( n8499 , n10451 );
    or g121 ( n12046 , n10812 , n2937 );
    xnor g122 ( n2932 , n4047 , n10504 );
    and g123 ( n3026 , n3135 , n5808 );
    and g124 ( n12849 , n8207 , n1545 );
    xnor g125 ( n4076 , n12132 , n965 );
    or g126 ( n7769 , n7041 , n12695 );
    xnor g127 ( n11615 , n1868 , n639 );
    xnor g128 ( n12282 , n6713 , n6848 );
    or g129 ( n4146 , n8868 , n2958 );
    not g130 ( n12518 , n2646 );
    and g131 ( n4928 , n2430 , n13186 );
    xnor g132 ( n2372 , n8740 , n9673 );
    xnor g133 ( n1964 , n12106 , n11044 );
    or g134 ( n2158 , n5607 , n9431 );
    or g135 ( n12165 , n12737 , n5956 );
    and g136 ( n9096 , n11398 , n5467 );
    and g137 ( n6181 , n5378 , n7277 );
    xnor g138 ( n10765 , n5090 , n5825 );
    or g139 ( n10235 , n7933 , n7244 );
    or g140 ( n10691 , n4755 , n10289 );
    xnor g141 ( n11500 , n7563 , n3718 );
    xnor g142 ( n2741 , n10187 , n4817 );
    not g143 ( n12881 , n4470 );
    or g144 ( n8882 , n48 , n4947 );
    and g145 ( n12252 , n5759 , n664 );
    xnor g146 ( n11017 , n5932 , n284 );
    or g147 ( n8688 , n2580 , n7533 );
    or g148 ( n6625 , n7931 , n11255 );
    or g149 ( n7215 , n11183 , n7859 );
    not g150 ( n10018 , n8468 );
    and g151 ( n3622 , n8063 , n3371 );
    xnor g152 ( n11049 , n2108 , n7715 );
    nor g153 ( n7369 , n2074 , n6239 );
    xnor g154 ( n7264 , n3499 , n5493 );
    nor g155 ( n15 , n2867 , n11302 );
    and g156 ( n6977 , n7625 , n3577 );
    xnor g157 ( n1657 , n1414 , n11594 );
    and g158 ( n8071 , n11471 , n3006 );
    and g159 ( n8822 , n2106 , n10607 );
    xnor g160 ( n8482 , n8706 , n9916 );
    and g161 ( n6836 , n6039 , n5862 );
    nor g162 ( n8910 , n745 , n1899 );
    not g163 ( n6581 , n12682 );
    and g164 ( n4969 , n264 , n10423 );
    not g165 ( n4875 , n1198 );
    buf g166 ( n7723 , n10879 );
    and g167 ( n4889 , n10680 , n4121 );
    not g168 ( n1511 , n12263 );
    and g169 ( n10200 , n5671 , n8233 );
    and g170 ( n9518 , n6162 , n8361 );
    not g171 ( n3167 , n2840 );
    or g172 ( n12055 , n9429 , n12501 );
    xnor g173 ( n3747 , n8035 , n9201 );
    xnor g174 ( n1459 , n1525 , n4142 );
    xnor g175 ( n7157 , n2593 , n8114 );
    or g176 ( n2025 , n4595 , n11343 );
    not g177 ( n8315 , n772 );
    and g178 ( n5117 , n8183 , n10606 );
    xnor g179 ( n10969 , n2741 , n7724 );
    or g180 ( n9023 , n1365 , n11162 );
    xnor g181 ( n11207 , n4982 , n12583 );
    xnor g182 ( n8844 , n9406 , n3154 );
    xnor g183 ( n5897 , n405 , n1808 );
    or g184 ( n9959 , n5670 , n10135 );
    xnor g185 ( n5651 , n3346 , n1154 );
    or g186 ( n2272 , n965 , n7619 );
    xnor g187 ( n12545 , n6303 , n2855 );
    xnor g188 ( n6019 , n1466 , n5895 );
    not g189 ( n7748 , n772 );
    or g190 ( n1773 , n5605 , n5868 );
    xnor g191 ( n5741 , n123 , n5069 );
    not g192 ( n8776 , n401 );
    or g193 ( n6970 , n7597 , n6265 );
    xnor g194 ( n7467 , n2424 , n5326 );
    and g195 ( n1797 , n11535 , n8925 );
    not g196 ( n663 , n12379 );
    xnor g197 ( n3064 , n4914 , n10942 );
    not g198 ( n3127 , n6818 );
    or g199 ( n5021 , n11125 , n998 );
    xnor g200 ( n7406 , n13149 , n9556 );
    not g201 ( n7055 , n10418 );
    xnor g202 ( n5403 , n9797 , n1532 );
    xnor g203 ( n8895 , n4557 , n11784 );
    nor g204 ( n12945 , n681 , n8347 );
    or g205 ( n6336 , n6743 , n4936 );
    or g206 ( n9803 , n59 , n5406 );
    and g207 ( n8253 , n10998 , n11890 );
    not g208 ( n1039 , n224 );
    and g209 ( n12475 , n7125 , n12365 );
    xnor g210 ( n1123 , n11737 , n2953 );
    or g211 ( n4878 , n3122 , n10100 );
    not g212 ( n12483 , n12853 );
    xnor g213 ( n11066 , n9898 , n2 );
    or g214 ( n9060 , n454 , n2192 );
    xnor g215 ( n6801 , n2647 , n58 );
    or g216 ( n11464 , n4808 , n2133 );
    not g217 ( n56 , n12893 );
    or g218 ( n3394 , n2109 , n2232 );
    xnor g219 ( n8591 , n5698 , n3242 );
    and g220 ( n12397 , n2986 , n1262 );
    or g221 ( n5936 , n11482 , n8822 );
    or g222 ( n12536 , n3346 , n10828 );
    and g223 ( n182 , n7840 , n12178 );
    or g224 ( n5374 , n8977 , n6404 );
    or g225 ( n5665 , n5260 , n7302 );
    or g226 ( n6797 , n1329 , n12847 );
    and g227 ( n11384 , n10300 , n5027 );
    not g228 ( n544 , n7328 );
    and g229 ( n9948 , n13239 , n826 );
    nor g230 ( n7302 , n972 , n10692 );
    xnor g231 ( n12985 , n12564 , n295 );
    or g232 ( n6934 , n4842 , n1686 );
    not g233 ( n10213 , n11488 );
    xnor g234 ( n4065 , n9986 , n9694 );
    nor g235 ( n4118 , n4117 , n3250 );
    xnor g236 ( n548 , n3150 , n6695 );
    or g237 ( n11717 , n850 , n6339 );
    xnor g238 ( n10634 , n641 , n12418 );
    xnor g239 ( n2885 , n8464 , n9392 );
    or g240 ( n7889 , n6250 , n479 );
    and g241 ( n10884 , n5639 , n7441 );
    or g242 ( n4336 , n6699 , n9784 );
    xnor g243 ( n7686 , n4311 , n7280 );
    and g244 ( n4585 , n6714 , n12135 );
    xnor g245 ( n5941 , n7983 , n10957 );
    xnor g246 ( n2699 , n2064 , n6719 );
    or g247 ( n1667 , n12621 , n12695 );
    or g248 ( n1128 , n5597 , n5846 );
    xnor g249 ( n7241 , n1858 , n8884 );
    or g250 ( n4706 , n7207 , n6789 );
    xnor g251 ( n12100 , n8789 , n11047 );
    not g252 ( n1720 , n854 );
    or g253 ( n1727 , n7903 , n12768 );
    and g254 ( n2694 , n3859 , n10391 );
    or g255 ( n11269 , n10950 , n7723 );
    and g256 ( n12665 , n3311 , n854 );
    xnor g257 ( n9038 , n4915 , n11245 );
    xor g258 ( n7103 , n8280 , n7205 );
    xnor g259 ( n11224 , n1700 , n6224 );
    xnor g260 ( n10194 , n7726 , n9611 );
    or g261 ( n8063 , n7571 , n9749 );
    or g262 ( n9003 , n1986 , n5515 );
    xnor g263 ( n2603 , n11198 , n9001 );
    nor g264 ( n12041 , n12652 , n12699 );
    xnor g265 ( n10243 , n9664 , n5837 );
    nor g266 ( n8126 , n3976 , n3723 );
    xnor g267 ( n509 , n11533 , n8434 );
    nor g268 ( n926 , n10067 , n11759 );
    not g269 ( n3428 , n772 );
    and g270 ( n6790 , n10770 , n8290 );
    xnor g271 ( n7120 , n10782 , n12379 );
    and g272 ( n1432 , n10770 , n8506 );
    nor g273 ( n3993 , n3936 , n4810 );
    or g274 ( n8434 , n10287 , n4724 );
    and g275 ( n10369 , n2036 , n2434 );
    xnor g276 ( n2820 , n5750 , n5873 );
    xnor g277 ( n11906 , n11583 , n11939 );
    nor g278 ( n10844 , n6507 , n5848 );
    xnor g279 ( n5991 , n11605 , n3565 );
    xnor g280 ( n3182 , n12290 , n207 );
    and g281 ( n1127 , n6084 , n8061 );
    xnor g282 ( n8535 , n7139 , n886 );
    and g283 ( n6715 , n8625 , n9970 );
    xnor g284 ( n12405 , n9026 , n1435 );
    and g285 ( n12489 , n869 , n11564 );
    or g286 ( n10275 , n12829 , n6461 );
    nor g287 ( n6766 , n10996 , n12420 );
    or g288 ( n895 , n11793 , n4354 );
    xnor g289 ( n6200 , n1966 , n3658 );
    or g290 ( n5125 , n7216 , n4947 );
    and g291 ( n8232 , n2916 , n4466 );
    not g292 ( n3698 , n3085 );
    and g293 ( n9623 , n4884 , n1116 );
    xnor g294 ( n5759 , n11271 , n1944 );
    or g295 ( n7298 , n12955 , n8360 );
    xnor g296 ( n13065 , n11051 , n5718 );
    or g297 ( n4814 , n3158 , n2133 );
    or g298 ( n12076 , n10448 , n11101 );
    and g299 ( n3499 , n9170 , n4661 );
    not g300 ( n7258 , n966 );
    not g301 ( n5466 , n9831 );
    or g302 ( n9354 , n6964 , n1211 );
    and g303 ( n684 , n156 , n2342 );
    xnor g304 ( n13035 , n680 , n2364 );
    or g305 ( n1952 , n10369 , n12854 );
    and g306 ( n7505 , n9975 , n5700 );
    xnor g307 ( n1378 , n7408 , n893 );
    nor g308 ( n3432 , n4910 , n2820 );
    and g309 ( n7681 , n11391 , n516 );
    xnor g310 ( n1009 , n4594 , n11293 );
    xnor g311 ( n11528 , n12916 , n2735 );
    or g312 ( n5451 , n3049 , n11137 );
    xnor g313 ( n870 , n5330 , n8870 );
    or g314 ( n11889 , n11092 , n8712 );
    nor g315 ( n274 , n10086 , n1322 );
    nor g316 ( n1816 , n5099 , n364 );
    and g317 ( n8711 , n3488 , n5835 );
    xnor g318 ( n8045 , n11306 , n1909 );
    not g319 ( n5854 , n9654 );
    and g320 ( n4148 , n6718 , n8567 );
    not g321 ( n6276 , n7969 );
    not g322 ( n2215 , n10264 );
    or g323 ( n10363 , n2785 , n10802 );
    or g324 ( n3736 , n4029 , n12800 );
    not g325 ( n392 , n10805 );
    xnor g326 ( n1523 , n8333 , n2906 );
    or g327 ( n5909 , n11344 , n9480 );
    xnor g328 ( n9058 , n7915 , n4106 );
    not g329 ( n6101 , n6080 );
    or g330 ( n4479 , n1320 , n4237 );
    not g331 ( n1323 , n9887 );
    or g332 ( n2727 , n7455 , n7734 );
    and g333 ( n3146 , n1527 , n6961 );
    nor g334 ( n8865 , n4591 , n1885 );
    not g335 ( n3829 , n6124 );
    xnor g336 ( n3233 , n11991 , n7273 );
    xnor g337 ( n8698 , n11223 , n9998 );
    xnor g338 ( n11480 , n9789 , n5206 );
    or g339 ( n4666 , n8675 , n7127 );
    or g340 ( n6098 , n7657 , n11608 );
    or g341 ( n3812 , n1475 , n1714 );
    xnor g342 ( n10472 , n13151 , n5156 );
    xnor g343 ( n2397 , n8743 , n408 );
    not g344 ( n4537 , n10866 );
    and g345 ( n7474 , n5126 , n7225 );
    xnor g346 ( n7175 , n4591 , n9284 );
    and g347 ( n10810 , n17 , n11460 );
    xnor g348 ( n6935 , n3991 , n12749 );
    nor g349 ( n2867 , n8207 , n1545 );
    or g350 ( n12294 , n560 , n7530 );
    or g351 ( n5141 , n10109 , n62 );
    and g352 ( n5614 , n8289 , n5294 );
    xnor g353 ( n11789 , n996 , n11902 );
    not g354 ( n8977 , n1650 );
    xnor g355 ( n8289 , n4193 , n12634 );
    or g356 ( n230 , n7395 , n8535 );
    xnor g357 ( n3147 , n10089 , n6641 );
    or g358 ( n3582 , n8074 , n7668 );
    and g359 ( n3248 , n8976 , n13179 );
    xnor g360 ( n5393 , n513 , n651 );
    or g361 ( n4574 , n6295 , n12188 );
    not g362 ( n12391 , n6155 );
    nor g363 ( n533 , n6504 , n9459 );
    or g364 ( n51 , n3260 , n10823 );
    or g365 ( n10044 , n6949 , n7524 );
    xnor g366 ( n8003 , n8072 , n4549 );
    xnor g367 ( n2402 , n10052 , n10264 );
    xnor g368 ( n1561 , n11576 , n12742 );
    xor g369 ( n2185 , n11102 , n12014 );
    xnor g370 ( n8205 , n5664 , n3556 );
    or g371 ( n5438 , n694 , n6635 );
    not g372 ( n11137 , n9475 );
    xnor g373 ( n4718 , n7818 , n7274 );
    and g374 ( n2290 , n10375 , n1128 );
    not g375 ( n9296 , n5770 );
    not g376 ( n2386 , n5136 );
    and g377 ( n1843 , n2767 , n10584 );
    not g378 ( n9720 , n7330 );
    not g379 ( n855 , n11473 );
    and g380 ( n332 , n67 , n2774 );
    and g381 ( n10445 , n13234 , n2257 );
    xnor g382 ( n1752 , n10102 , n11894 );
    or g383 ( n12259 , n4272 , n12847 );
    xnor g384 ( n429 , n13177 , n2844 );
    nor g385 ( n9627 , n9654 , n11323 );
    or g386 ( n3695 , n13082 , n12273 );
    or g387 ( n2591 , n7718 , n5242 );
    and g388 ( n90 , n8339 , n8542 );
    not g389 ( n1663 , n8137 );
    nor g390 ( n8095 , n12747 , n10337 );
    nor g391 ( n7881 , n12896 , n3312 );
    xnor g392 ( n10569 , n12468 , n1255 );
    nor g393 ( n7775 , n1632 , n12013 );
    nor g394 ( n1531 , n13132 , n3777 );
    not g395 ( n9569 , n4712 );
    and g396 ( n6228 , n761 , n834 );
    xnor g397 ( n3946 , n11968 , n12523 );
    and g398 ( n9352 , n4745 , n12411 );
    buf g399 ( n2675 , n5045 );
    xor g400 ( n9577 , n2486 , n11084 );
    not g401 ( n6099 , n287 );
    xnor g402 ( n4341 , n4533 , n12320 );
    or g403 ( n1594 , n3613 , n9130 );
    not g404 ( n8671 , n5800 );
    or g405 ( n6873 , n10501 , n12959 );
    or g406 ( n178 , n10343 , n9182 );
    and g407 ( n13113 , n3453 , n5335 );
    xnor g408 ( n11699 , n9176 , n3054 );
    xnor g409 ( n6311 , n3400 , n1203 );
    or g410 ( n11801 , n1406 , n8534 );
    and g411 ( n7251 , n4994 , n10077 );
    and g412 ( n12189 , n2853 , n2854 );
    and g413 ( n5069 , n2850 , n8526 );
    or g414 ( n1955 , n3068 , n6732 );
    not g415 ( n5377 , n10405 );
    not g416 ( n4152 , n3918 );
    buf g417 ( n6769 , n9272 );
    and g418 ( n5399 , n3607 , n8996 );
    nor g419 ( n2997 , n4593 , n6096 );
    and g420 ( n10914 , n3415 , n11558 );
    xnor g421 ( n2496 , n5094 , n7517 );
    and g422 ( n11981 , n7543 , n931 );
    or g423 ( n739 , n9793 , n12789 );
    and g424 ( n3519 , n2107 , n8548 );
    not g425 ( n1193 , n11325 );
    or g426 ( n12300 , n1213 , n7682 );
    xnor g427 ( n5727 , n11867 , n421 );
    or g428 ( n11662 , n1735 , n10674 );
    nor g429 ( n11301 , n6653 , n7490 );
    or g430 ( n7195 , n4016 , n4095 );
    or g431 ( n1514 , n1090 , n1292 );
    xnor g432 ( n2389 , n2023 , n5824 );
    nor g433 ( n2911 , n10278 , n1441 );
    or g434 ( n8704 , n2615 , n2871 );
    not g435 ( n5375 , n7877 );
    xnor g436 ( n2898 , n4861 , n8377 );
    xnor g437 ( n4381 , n3291 , n3601 );
    or g438 ( n7605 , n12568 , n12273 );
    or g439 ( n4105 , n4539 , n11234 );
    nor g440 ( n3697 , n7549 , n2597 );
    xnor g441 ( n463 , n3247 , n3560 );
    or g442 ( n2596 , n8613 , n7312 );
    not g443 ( n2478 , n11468 );
    xor g444 ( n13056 , n6489 , n2342 );
    and g445 ( n2996 , n1375 , n12097 );
    xnor g446 ( n9031 , n377 , n10083 );
    nor g447 ( n3689 , n5030 , n12908 );
    or g448 ( n4506 , n4044 , n12672 );
    or g449 ( n1419 , n3534 , n4947 );
    and g450 ( n8101 , n2609 , n5342 );
    xnor g451 ( n3043 , n6049 , n8427 );
    xnor g452 ( n5126 , n10506 , n10151 );
    xnor g453 ( n3081 , n12492 , n7263 );
    nor g454 ( n11804 , n7304 , n11649 );
    or g455 ( n3982 , n9882 , n4373 );
    xor g456 ( n2457 , n4001 , n9692 );
    xnor g457 ( n3511 , n10667 , n11474 );
    nor g458 ( n4502 , n7870 , n5043 );
    and g459 ( n1971 , n6668 , n12853 );
    or g460 ( n399 , n3544 , n1702 );
    and g461 ( n9564 , n7095 , n4211 );
    nor g462 ( n6266 , n10405 , n608 );
    not g463 ( n12834 , n5758 );
    not g464 ( n9321 , n5094 );
    nor g465 ( n5198 , n2237 , n9953 );
    not g466 ( n12272 , n983 );
    or g467 ( n7857 , n4004 , n9549 );
    xnor g468 ( n7666 , n3916 , n4907 );
    xnor g469 ( n1115 , n5410 , n2779 );
    xnor g470 ( n5408 , n3985 , n885 );
    xor g471 ( n10498 , n10013 , n12578 );
    not g472 ( n6375 , n469 );
    or g473 ( n3083 , n10188 , n3963 );
    xnor g474 ( n10718 , n10888 , n4826 );
    xnor g475 ( n8854 , n11573 , n9844 );
    and g476 ( n210 , n1934 , n1234 );
    or g477 ( n11453 , n4467 , n12142 );
    or g478 ( n11636 , n6355 , n3890 );
    and g479 ( n10322 , n4382 , n1636 );
    and g480 ( n292 , n13229 , n7849 );
    and g481 ( n9220 , n5005 , n13110 );
    not g482 ( n1930 , n7374 );
    xnor g483 ( n9271 , n1880 , n6551 );
    xnor g484 ( n4672 , n10482 , n4254 );
    and g485 ( n2409 , n8661 , n5568 );
    xnor g486 ( n10371 , n10940 , n5821 );
    and g487 ( n9032 , n78 , n116 );
    xnor g488 ( n7027 , n11092 , n8712 );
    xnor g489 ( n7525 , n5996 , n6844 );
    and g490 ( n6474 , n1514 , n8318 );
    or g491 ( n7432 , n241 , n9070 );
    or g492 ( n10678 , n3299 , n7741 );
    xnor g493 ( n2549 , n4889 , n1122 );
    xnor g494 ( n2497 , n2176 , n10951 );
    xnor g495 ( n6026 , n12553 , n4350 );
    not g496 ( n6046 , n11830 );
    not g497 ( n1271 , n972 );
    nor g498 ( n3381 , n10378 , n4249 );
    xnor g499 ( n11526 , n11658 , n5101 );
    xnor g500 ( n5339 , n6859 , n4823 );
    and g501 ( n933 , n2263 , n1443 );
    and g502 ( n10111 , n12972 , n3927 );
    xnor g503 ( n3969 , n988 , n4873 );
    xnor g504 ( n3765 , n3214 , n7173 );
    and g505 ( n2361 , n1175 , n8084 );
    xnor g506 ( n4052 , n10931 , n13164 );
    xnor g507 ( n6662 , n6515 , n8755 );
    not g508 ( n765 , n9 );
    and g509 ( n6541 , n13109 , n12435 );
    and g510 ( n9259 , n5545 , n2025 );
    xnor g511 ( n9554 , n2044 , n13048 );
    and g512 ( n11395 , n11331 , n2881 );
    or g513 ( n11489 , n5440 , n2244 );
    or g514 ( n8091 , n3047 , n12273 );
    xnor g515 ( n8203 , n5798 , n6252 );
    xnor g516 ( n6681 , n3205 , n9751 );
    or g517 ( n8349 , n8206 , n2059 );
    not g518 ( n7052 , n8253 );
    nor g519 ( n7594 , n3504 , n13045 );
    nor g520 ( n12464 , n12628 , n5484 );
    nor g521 ( n5388 , n9095 , n3813 );
    xnor g522 ( n4931 , n12021 , n6893 );
    buf g523 ( n10179 , n2623 );
    xnor g524 ( n2164 , n228 , n6127 );
    or g525 ( n7297 , n12050 , n4899 );
    not g526 ( n2307 , n3496 );
    and g527 ( n1474 , n2247 , n12928 );
    or g528 ( n12274 , n3099 , n3074 );
    xnor g529 ( n4948 , n5561 , n2060 );
    or g530 ( n9880 , n9722 , n9974 );
    not g531 ( n8188 , n761 );
    and g532 ( n1910 , n2425 , n2380 );
    xnor g533 ( n1330 , n4977 , n1221 );
    nor g534 ( n6567 , n2732 , n11081 );
    xnor g535 ( n5706 , n3305 , n9368 );
    not g536 ( n8665 , n4743 );
    and g537 ( n6879 , n1059 , n6856 );
    nor g538 ( n5417 , n4427 , n5663 );
    and g539 ( n2569 , n11617 , n11630 );
    or g540 ( n150 , n10943 , n6511 );
    xnor g541 ( n5642 , n1143 , n6994 );
    and g542 ( n2342 , n1364 , n3815 );
    or g543 ( n10507 , n7669 , n9101 );
    xor g544 ( n5389 , n10253 , n12182 );
    not g545 ( n13198 , n4337 );
    xnor g546 ( n8336 , n7491 , n1362 );
    and g547 ( n11164 , n4625 , n9331 );
    or g548 ( n9237 , n8386 , n615 );
    or g549 ( n6491 , n9702 , n1571 );
    and g550 ( n8204 , n228 , n2829 );
    or g551 ( n1520 , n1270 , n6903 );
    xnor g552 ( n11777 , n13180 , n3624 );
    xnor g553 ( n2242 , n2014 , n13224 );
    xnor g554 ( n11936 , n9678 , n9999 );
    and g555 ( n3480 , n2156 , n7971 );
    and g556 ( n3327 , n8653 , n2808 );
    nor g557 ( n986 , n6761 , n2571 );
    and g558 ( n649 , n1769 , n12117 );
    nor g559 ( n10528 , n5421 , n9376 );
    xnor g560 ( n5825 , n7638 , n3728 );
    and g561 ( n7667 , n12246 , n888 );
    xnor g562 ( n5062 , n10288 , n1014 );
    or g563 ( n809 , n10434 , n12723 );
    or g564 ( n2516 , n12930 , n1144 );
    or g565 ( n12791 , n10558 , n12273 );
    not g566 ( n5917 , n1707 );
    and g567 ( n10134 , n11635 , n2482 );
    not g568 ( n3524 , n4574 );
    or g569 ( n4204 , n5842 , n10761 );
    xnor g570 ( n10913 , n8382 , n4813 );
    or g571 ( n9727 , n4275 , n9842 );
    xnor g572 ( n501 , n11461 , n2444 );
    and g573 ( n3544 , n13218 , n9420 );
    and g574 ( n3000 , n10097 , n12071 );
    not g575 ( n379 , n5536 );
    not g576 ( n12648 , n1982 );
    not g577 ( n107 , n10537 );
    not g578 ( n11887 , n4479 );
    xnor g579 ( n1666 , n10902 , n12198 );
    or g580 ( n9122 , n12324 , n2133 );
    and g581 ( n3828 , n8077 , n9720 );
    not g582 ( n2725 , n4688 );
    xnor g583 ( n3496 , n5593 , n5055 );
    xor g584 ( n10149 , n12832 , n1174 );
    xor g585 ( n5725 , n3352 , n3435 );
    and g586 ( n8495 , n12643 , n11888 );
    xnor g587 ( n10348 , n535 , n7178 );
    not g588 ( n1388 , n9428 );
    or g589 ( n5130 , n3928 , n1985 );
    xnor g590 ( n2031 , n11266 , n3774 );
    not g591 ( n5562 , n10408 );
    and g592 ( n3645 , n10416 , n12306 );
    or g593 ( n12119 , n9323 , n1797 );
    or g594 ( n3302 , n1919 , n4373 );
    xnor g595 ( n10622 , n10688 , n9990 );
    xnor g596 ( n6263 , n2363 , n11420 );
    not g597 ( n39 , n4240 );
    not g598 ( n2081 , n9794 );
    or g599 ( n3477 , n12563 , n4949 );
    and g600 ( n4950 , n7457 , n3117 );
    or g601 ( n1220 , n5583 , n6017 );
    or g602 ( n1176 , n10037 , n4373 );
    xnor g603 ( n502 , n4486 , n8345 );
    and g604 ( n5047 , n1208 , n7264 );
    not g605 ( n45 , n1084 );
    or g606 ( n9656 , n5297 , n11619 );
    and g607 ( n5033 , n3752 , n6153 );
    or g608 ( n2712 , n2849 , n2793 );
    and g609 ( n11275 , n5058 , n1922 );
    xnor g610 ( n13171 , n9972 , n9555 );
    not g611 ( n672 , n192 );
    xnor g612 ( n9274 , n8133 , n3302 );
    xnor g613 ( n11590 , n11954 , n12210 );
    and g614 ( n11495 , n60 , n5230 );
    nor g615 ( n2905 , n5034 , n4222 );
    xnor g616 ( n5159 , n1062 , n3947 );
    not g617 ( n9641 , n988 );
    or g618 ( n7598 , n11987 , n3019 );
    nor g619 ( n2616 , n5929 , n10215 );
    or g620 ( n188 , n9059 , n4089 );
    xnor g621 ( n9469 , n5736 , n3986 );
    and g622 ( n6938 , n2024 , n6508 );
    or g623 ( n1448 , n1263 , n4058 );
    and g624 ( n3772 , n10189 , n7743 );
    xnor g625 ( n11589 , n87 , n7373 );
    and g626 ( n1943 , n6583 , n7231 );
    or g627 ( n12342 , n6816 , n4551 );
    not g628 ( n10636 , n7845 );
    xnor g629 ( n5678 , n2644 , n6709 );
    or g630 ( n4456 , n11449 , n8348 );
    and g631 ( n4644 , n10603 , n6540 );
    xnor g632 ( n7554 , n7099 , n2620 );
    xnor g633 ( n459 , n9851 , n5144 );
    nor g634 ( n7349 , n7484 , n3848 );
    not g635 ( n11018 , n4006 );
    not g636 ( n12926 , n12867 );
    and g637 ( n7704 , n7232 , n8733 );
    not g638 ( n6699 , n5189 );
    or g639 ( n3956 , n2289 , n3538 );
    or g640 ( n10422 , n2457 , n8964 );
    nor g641 ( n4266 , n12250 , n8692 );
    not g642 ( n3169 , n10908 );
    and g643 ( n6909 , n518 , n7776 );
    xnor g644 ( n10542 , n5695 , n7339 );
    not g645 ( n1094 , n5244 );
    nor g646 ( n4697 , n12184 , n10030 );
    or g647 ( n9731 , n1360 , n3972 );
    and g648 ( n12155 , n6177 , n5857 );
    xnor g649 ( n594 , n13187 , n12641 );
    not g650 ( n10143 , n9570 );
    or g651 ( n11515 , n2246 , n6145 );
    xnor g652 ( n3713 , n6058 , n2976 );
    or g653 ( n13109 , n1131 , n1153 );
    nor g654 ( n2260 , n3272 , n12869 );
    or g655 ( n6139 , n12485 , n9192 );
    or g656 ( n8594 , n4515 , n10681 );
    and g657 ( n1229 , n599 , n876 );
    not g658 ( n8019 , n8410 );
    not g659 ( n11928 , n6826 );
    or g660 ( n2766 , n1438 , n1985 );
    xnor g661 ( n6868 , n3260 , n1913 );
    nor g662 ( n8169 , n3448 , n8317 );
    and g663 ( n2393 , n2458 , n3409 );
    or g664 ( n3007 , n9450 , n12623 );
    not g665 ( n5048 , n3085 );
    or g666 ( n9266 , n6254 , n8326 );
    not g667 ( n4453 , n951 );
    and g668 ( n10011 , n4088 , n7043 );
    or g669 ( n10056 , n8108 , n10179 );
    nor g670 ( n6860 , n4528 , n12906 );
    xnor g671 ( n3010 , n3366 , n570 );
    not g672 ( n11130 , n180 );
    nor g673 ( n1338 , n8368 , n9441 );
    xnor g674 ( n2371 , n7879 , n6997 );
    xnor g675 ( n3974 , n4113 , n1707 );
    not g676 ( n10043 , n3085 );
    and g677 ( n6331 , n1936 , n4383 );
    or g678 ( n8636 , n4148 , n900 );
    nor g679 ( n3218 , n8042 , n2533 );
    not g680 ( n6755 , n8768 );
    xnor g681 ( n1336 , n11262 , n5379 );
    and g682 ( n954 , n11355 , n7774 );
    or g683 ( n8211 , n8843 , n4640 );
    not g684 ( n3813 , n5073 );
    xnor g685 ( n5895 , n11448 , n9226 );
    not g686 ( n644 , n3669 );
    xnor g687 ( n10737 , n10735 , n5276 );
    xnor g688 ( n11979 , n129 , n2929 );
    and g689 ( n4557 , n428 , n5117 );
    xnor g690 ( n9241 , n798 , n7603 );
    or g691 ( n1227 , n3965 , n5460 );
    or g692 ( n12060 , n11203 , n3926 );
    or g693 ( n3483 , n1712 , n12784 );
    nor g694 ( n279 , n1801 , n2477 );
    not g695 ( n10673 , n6956 );
    xnor g696 ( n6206 , n8926 , n9469 );
    or g697 ( n9026 , n4980 , n2875 );
    nor g698 ( n6117 , n91 , n7641 );
    or g699 ( n8847 , n53 , n10761 );
    or g700 ( n9255 , n2973 , n5646 );
    xnor g701 ( n27 , n9633 , n12887 );
    and g702 ( n11775 , n6140 , n3031 );
    or g703 ( n3768 , n5922 , n7874 );
    or g704 ( n9249 , n11591 , n10319 );
    and g705 ( n741 , n3077 , n2687 );
    and g706 ( n9369 , n12262 , n3227 );
    or g707 ( n7999 , n5401 , n13039 );
    or g708 ( n3665 , n9392 , n8464 );
    xnor g709 ( n5046 , n12899 , n6899 );
    xnor g710 ( n5929 , n10865 , n3010 );
    xnor g711 ( n11044 , n7929 , n7735 );
    or g712 ( n1542 , n6606 , n8504 );
    or g713 ( n12327 , n12798 , n12240 );
    xnor g714 ( n8181 , n9059 , n4089 );
    not g715 ( n5402 , n7841 );
    xnor g716 ( n1298 , n9307 , n9097 );
    and g717 ( n7463 , n7296 , n8914 );
    xnor g718 ( n8970 , n2205 , n2654 );
    xnor g719 ( n985 , n6362 , n7772 );
    xnor g720 ( n393 , n576 , n3757 );
    not g721 ( n7286 , n6347 );
    or g722 ( n12809 , n5806 , n121 );
    nor g723 ( n8944 , n7786 , n9562 );
    and g724 ( n1592 , n7086 , n666 );
    nor g725 ( n11884 , n9047 , n12231 );
    and g726 ( n11342 , n11842 , n10197 );
    xnor g727 ( n722 , n10007 , n9337 );
    or g728 ( n357 , n9927 , n10493 );
    xnor g729 ( n9798 , n4930 , n3070 );
    xnor g730 ( n6461 , n9610 , n6456 );
    xnor g731 ( n9210 , n13150 , n2396 );
    xnor g732 ( n2113 , n5699 , n3604 );
    not g733 ( n209 , n7888 );
    or g734 ( n7931 , n10043 , n2675 );
    nor g735 ( n616 , n4263 , n1649 );
    and g736 ( n4758 , n4382 , n12284 );
    or g737 ( n7029 , n11311 , n5712 );
    xnor g738 ( n5960 , n1041 , n10910 );
    or g739 ( n3749 , n6220 , n894 );
    nor g740 ( n7186 , n600 , n12425 );
    xor g741 ( n12746 , n860 , n5393 );
    and g742 ( n10843 , n9513 , n1400 );
    xnor g743 ( n8782 , n11589 , n6312 );
    nor g744 ( n6356 , n9025 , n11374 );
    xnor g745 ( n3705 , n7320 , n8267 );
    not g746 ( n569 , n2758 );
    not g747 ( n7199 , n2787 );
    not g748 ( n946 , n5427 );
    not g749 ( n6939 , n4330 );
    xnor g750 ( n10464 , n5537 , n11629 );
    or g751 ( n11596 , n8801 , n4644 );
    and g752 ( n7728 , n875 , n4509 );
    and g753 ( n3797 , n10757 , n467 );
    or g754 ( n623 , n6326 , n12543 );
    or g755 ( n1940 , n2048 , n9682 );
    and g756 ( n5287 , n778 , n10704 );
    and g757 ( n7446 , n10472 , n12172 );
    or g758 ( n7434 , n4037 , n7495 );
    xnor g759 ( n4168 , n13163 , n5143 );
    nor g760 ( n4197 , n12455 , n12161 );
    or g761 ( n12162 , n6721 , n5076 );
    xnor g762 ( n592 , n3541 , n2587 );
    or g763 ( n7031 , n12362 , n3987 );
    or g764 ( n4268 , n10780 , n8268 );
    nor g765 ( n3629 , n2739 , n9232 );
    xor g766 ( n5038 , n11640 , n3830 );
    or g767 ( n11553 , n338 , n2544 );
    or g768 ( n8402 , n9238 , n12166 );
    not g769 ( n12856 , n1369 );
    xnor g770 ( n439 , n8815 , n7622 );
    or g771 ( n3532 , n2899 , n1570 );
    not g772 ( n11799 , n10033 );
    xnor g773 ( n4101 , n7181 , n13103 );
    not g774 ( n5414 , n10770 );
    nor g775 ( n2998 , n9022 , n10038 );
    xnor g776 ( n10067 , n4695 , n9504 );
    or g777 ( n10513 , n1436 , n9159 );
    xnor g778 ( n3707 , n2149 , n2085 );
    xnor g779 ( n2620 , n108 , n2892 );
    xnor g780 ( n6561 , n4513 , n9267 );
    xnor g781 ( n8476 , n11321 , n748 );
    and g782 ( n13184 , n1258 , n4971 );
    xor g783 ( n8721 , n1025 , n8760 );
    xnor g784 ( n455 , n1904 , n6974 );
    xnor g785 ( n6788 , n631 , n11724 );
    xor g786 ( n1487 , n8253 , n7584 );
    or g787 ( n10920 , n13170 , n6404 );
    or g788 ( n10261 , n13012 , n1985 );
    or g789 ( n7017 , n860 , n8371 );
    or g790 ( n921 , n13194 , n4947 );
    and g791 ( n6257 , n8894 , n5898 );
    or g792 ( n12770 , n1892 , n1679 );
    not g793 ( n44 , n11109 );
    xnor g794 ( n2761 , n4153 , n7032 );
    or g795 ( n2359 , n808 , n4621 );
    xnor g796 ( n9541 , n10571 , n3798 );
    or g797 ( n6212 , n6182 , n2059 );
    not g798 ( n7045 , n6610 );
    nor g799 ( n2344 , n7705 , n5239 );
    or g800 ( n11714 , n1883 , n6404 );
    or g801 ( n2076 , n1451 , n2059 );
    or g802 ( n9848 , n234 , n3843 );
    or g803 ( n7843 , n6768 , n4455 );
    not g804 ( n4258 , n499 );
    not g805 ( n1175 , n5845 );
    or g806 ( n7911 , n2238 , n9586 );
    xnor g807 ( n11948 , n2301 , n7524 );
    xnor g808 ( n11444 , n7797 , n7525 );
    xnor g809 ( n12081 , n12230 , n9542 );
    xnor g810 ( n11587 , n5640 , n9746 );
    nor g811 ( n12317 , n550 , n6594 );
    xnor g812 ( n11406 , n8758 , n2629 );
    xnor g813 ( n9771 , n2820 , n4646 );
    and g814 ( n12520 , n7591 , n4547 );
    and g815 ( n431 , n4782 , n12793 );
    not g816 ( n4665 , n5884 );
    nor g817 ( n574 , n1759 , n11382 );
    not g818 ( n3652 , n3203 );
    xnor g819 ( n4946 , n3251 , n8686 );
    or g820 ( n12676 , n6166 , n9195 );
    xnor g821 ( n5868 , n7317 , n3261 );
    and g822 ( n9319 , n3914 , n8017 );
    not g823 ( n1335 , n5969 );
    or g824 ( n9597 , n11087 , n542 );
    and g825 ( n2668 , n66 , n4111 );
    xnor g826 ( n4119 , n4814 , n2891 );
    or g827 ( n12135 , n4741 , n177 );
    xnor g828 ( n3140 , n12399 , n10706 );
    not g829 ( n3867 , n11647 );
    xnor g830 ( n5886 , n296 , n1083 );
    xnor g831 ( n1481 , n11909 , n4125 );
    or g832 ( n3944 , n1897 , n1832 );
    not g833 ( n6015 , n11482 );
    not g834 ( n10292 , n3358 );
    xnor g835 ( n7905 , n12486 , n892 );
    xnor g836 ( n6297 , n3000 , n5751 );
    xnor g837 ( n13095 , n6517 , n6493 );
    and g838 ( n8981 , n448 , n10345 );
    not g839 ( n2636 , n4460 );
    nor g840 ( n9491 , n3271 , n10677 );
    nor g841 ( n4124 , n9437 , n779 );
    not g842 ( n3165 , n2569 );
    or g843 ( n3315 , n6224 , n7186 );
    not g844 ( n4087 , n3251 );
    or g845 ( n3795 , n11505 , n2367 );
    xnor g846 ( n12386 , n5687 , n3300 );
    not g847 ( n1632 , n8222 );
    nor g848 ( n9548 , n5220 , n11636 );
    not g849 ( n12899 , n6783 );
    and g850 ( n12255 , n2592 , n8860 );
    or g851 ( n4863 , n1737 , n8534 );
    not g852 ( n9893 , n42 );
    and g853 ( n65 , n4598 , n5843 );
    xnor g854 ( n7806 , n2834 , n5298 );
    not g855 ( n8065 , n7309 );
    not g856 ( n10998 , n9087 );
    xnor g857 ( n11147 , n4315 , n12278 );
    and g858 ( n6253 , n558 , n9294 );
    or g859 ( n668 , n6419 , n8030 );
    xnor g860 ( n3628 , n6771 , n7268 );
    and g861 ( n6746 , n6919 , n1559 );
    or g862 ( n1805 , n5401 , n617 );
    xnor g863 ( n2052 , n13128 , n12609 );
    not g864 ( n12371 , n6312 );
    and g865 ( n6800 , n5323 , n4094 );
    and g866 ( n1019 , n8058 , n2285 );
    or g867 ( n7622 , n1571 , n2675 );
    nor g868 ( n2461 , n4332 , n11200 );
    and g869 ( n8025 , n2475 , n6513 );
    or g870 ( n4717 , n2352 , n7049 );
    or g871 ( n4362 , n9711 , n9195 );
    not g872 ( n8301 , n5729 );
    and g873 ( n7442 , n4428 , n786 );
    or g874 ( n476 , n12653 , n3884 );
    or g875 ( n2980 , n8306 , n8563 );
    or g876 ( n11793 , n11920 , n8348 );
    not g877 ( n4855 , n443 );
    or g878 ( n4029 , n10991 , n7723 );
    not g879 ( n11544 , n12115 );
    xnor g880 ( n6661 , n2986 , n7744 );
    and g881 ( n12612 , n8940 , n7720 );
    and g882 ( n7327 , n13031 , n9399 );
    or g883 ( n8088 , n11150 , n2034 );
    xnor g884 ( n2256 , n3430 , n7557 );
    xnor g885 ( n5810 , n1213 , n8886 );
    xnor g886 ( n8667 , n11958 , n3469 );
    and g887 ( n10025 , n5243 , n10234 );
    nor g888 ( n6804 , n8930 , n8103 );
    and g889 ( n4576 , n6333 , n2295 );
    not g890 ( n1897 , n3964 );
    or g891 ( n9980 , n5448 , n5487 );
    xnor g892 ( n3410 , n4050 , n5305 );
    or g893 ( n1185 , n12671 , n5242 );
    and g894 ( n914 , n11854 , n8644 );
    xnor g895 ( n12154 , n7646 , n1464 );
    and g896 ( n4175 , n2771 , n2758 );
    not g897 ( n11370 , n3591 );
    or g898 ( n6088 , n3157 , n10471 );
    not g899 ( n7272 , n9336 );
    or g900 ( n2764 , n4792 , n10573 );
    not g901 ( n48 , n12284 );
    not g902 ( n8840 , n10622 );
    xnor g903 ( n4833 , n11838 , n9296 );
    or g904 ( n3951 , n3062 , n6769 );
    or g905 ( n4582 , n9129 , n3459 );
    and g906 ( n5336 , n4363 , n12888 );
    or g907 ( n11391 , n12964 , n2679 );
    or g908 ( n2533 , n10465 , n4949 );
    nor g909 ( n8781 , n10743 , n3399 );
    xnor g910 ( n577 , n1787 , n10399 );
    xnor g911 ( n5081 , n5993 , n1298 );
    or g912 ( n4445 , n11612 , n12328 );
    not g913 ( n9511 , n287 );
    xnor g914 ( n8214 , n11382 , n1759 );
    nor g915 ( n2612 , n11909 , n10595 );
    or g916 ( n12920 , n2729 , n76 );
    xnor g917 ( n811 , n3540 , n7909 );
    and g918 ( n11753 , n5966 , n8257 );
    not g919 ( n11982 , n3130 );
    not g920 ( n6482 , n170 );
    xnor g921 ( n8273 , n13139 , n4318 );
    or g922 ( n5435 , n9891 , n6973 );
    not g923 ( n4698 , n948 );
    and g924 ( n6151 , n1674 , n5274 );
    and g925 ( n6663 , n8211 , n6111 );
    xnor g926 ( n10505 , n302 , n2300 );
    xnor g927 ( n9142 , n12457 , n3449 );
    not g928 ( n2975 , n446 );
    not g929 ( n2493 , n12219 );
    or g930 ( n9441 , n1887 , n6635 );
    or g931 ( n4275 , n3537 , n8490 );
    or g932 ( n11100 , n3344 , n6635 );
    nor g933 ( n5950 , n5738 , n11403 );
    not g934 ( n8580 , n10276 );
    or g935 ( n5823 , n12581 , n5836 );
    not g936 ( n3384 , n2798 );
    and g937 ( n1223 , n6758 , n5930 );
    nor g938 ( n8748 , n502 , n3319 );
    or g939 ( n7202 , n13051 , n8383 );
    nor g940 ( n9337 , n9388 , n7520 );
    or g941 ( n5636 , n7798 , n2133 );
    or g942 ( n12971 , n6841 , n11609 );
    or g943 ( n311 , n4927 , n11100 );
    not g944 ( n5400 , n10504 );
    not g945 ( n11468 , n1742 );
    not g946 ( n5905 , n5083 );
    nor g947 ( n7981 , n2081 , n12810 );
    not g948 ( n12019 , n9585 );
    or g949 ( n5795 , n5713 , n1463 );
    xnor g950 ( n6122 , n5300 , n3125 );
    xnor g951 ( n7079 , n6605 , n6020 );
    and g952 ( n1792 , n1677 , n9814 );
    and g953 ( n9239 , n11061 , n287 );
    not g954 ( n5915 , n9833 );
    xnor g955 ( n7050 , n10420 , n7466 );
    not g956 ( n2600 , n1254 );
    not g957 ( n1857 , n1110 );
    and g958 ( n6280 , n12213 , n6045 );
    not g959 ( n7814 , n7537 );
    or g960 ( n7210 , n10400 , n4724 );
    or g961 ( n7109 , n11262 , n2992 );
    nor g962 ( n3801 , n5805 , n9786 );
    xnor g963 ( n3841 , n7153 , n13166 );
    nor g964 ( n9501 , n8369 , n3286 );
    xnor g965 ( n5429 , n7085 , n1266 );
    xnor g966 ( n11233 , n13236 , n4734 );
    nor g967 ( n5053 , n7938 , n11204 );
    or g968 ( n11035 , n12052 , n4253 );
    xnor g969 ( n2216 , n7183 , n6604 );
    xor g970 ( n4847 , n1498 , n9623 );
    or g971 ( n2972 , n1135 , n5264 );
    not g972 ( n9490 , n6892 );
    xnor g973 ( n11025 , n3273 , n1780 );
    or g974 ( n2507 , n6603 , n362 );
    or g975 ( n6508 , n8646 , n6732 );
    xnor g976 ( n3426 , n7210 , n12499 );
    not g977 ( n12768 , n3085 );
    or g978 ( n1457 , n4022 , n4936 );
    or g979 ( n11 , n4041 , n12404 );
    and g980 ( n12724 , n6684 , n2971 );
    or g981 ( n3916 , n7522 , n3703 );
    not g982 ( n407 , n7294 );
    or g983 ( n1001 , n5503 , n1452 );
    not g984 ( n10966 , n6085 );
    xnor g985 ( n11904 , n7271 , n8618 );
    nor g986 ( n8086 , n3765 , n10734 );
    nor g987 ( n4956 , n3278 , n12385 );
    not g988 ( n12303 , n1195 );
    or g989 ( n8871 , n8995 , n7863 );
    xnor g990 ( n4596 , n9058 , n4687 );
    and g991 ( n6920 , n10770 , n8233 );
    not g992 ( n902 , n8230 );
    not g993 ( n1945 , n10671 );
    or g994 ( n6537 , n7076 , n9223 );
    xnor g995 ( n12553 , n12168 , n904 );
    and g996 ( n4519 , n12481 , n8750 );
    not g997 ( n5607 , n3357 );
    or g998 ( n5900 , n11629 , n7768 );
    or g999 ( n4995 , n1451 , n121 );
    or g1000 ( n8832 , n10714 , n10474 );
    not g1001 ( n8325 , n4122 );
    xnor g1002 ( n9404 , n13240 , n7285 );
    or g1003 ( n12071 , n2646 , n9381 );
    or g1004 ( n12557 , n542 , n8702 );
    xnor g1005 ( n1374 , n3931 , n1790 );
    or g1006 ( n6651 , n69 , n8534 );
    not g1007 ( n9788 , n12692 );
    and g1008 ( n11421 , n4403 , n1828 );
    xnor g1009 ( n7499 , n11478 , n12208 );
    and g1010 ( n12800 , n4334 , n1777 );
    not g1011 ( n9786 , n5868 );
    and g1012 ( n3023 , n10845 , n200 );
    nor g1013 ( n10296 , n6615 , n450 );
    and g1014 ( n10547 , n6120 , n4783 );
    and g1015 ( n376 , n12099 , n11866 );
    xnor g1016 ( n7910 , n8161 , n38 );
    or g1017 ( n3637 , n2109 , n2726 );
    and g1018 ( n3500 , n11849 , n3778 );
    or g1019 ( n12777 , n9400 , n11107 );
    nor g1020 ( n7507 , n6445 , n3845 );
    not g1021 ( n5692 , n6068 );
    or g1022 ( n8255 , n5535 , n9847 );
    xnor g1023 ( n4917 , n9487 , n4870 );
    not g1024 ( n9793 , n11734 );
    or g1025 ( n255 , n7473 , n196 );
    or g1026 ( n10386 , n2710 , n1871 );
    xnor g1027 ( n3734 , n5961 , n8190 );
    and g1028 ( n5739 , n7484 , n3848 );
    xnor g1029 ( n1619 , n3193 , n5803 );
    not g1030 ( n6194 , n9343 );
    not g1031 ( n3380 , n2597 );
    nor g1032 ( n1243 , n3150 , n6839 );
    xnor g1033 ( n1276 , n7592 , n11299 );
    nor g1034 ( n12399 , n2103 , n12325 );
    or g1035 ( n174 , n9588 , n10708 );
    and g1036 ( n4113 , n9736 , n10667 );
    nor g1037 ( n11483 , n11233 , n12498 );
    or g1038 ( n5633 , n11235 , n6113 );
    not g1039 ( n894 , n12853 );
    xnor g1040 ( n3541 , n1839 , n11409 );
    not g1041 ( n2884 , n497 );
    or g1042 ( n3030 , n2484 , n8383 );
    and g1043 ( n9831 , n9283 , n7220 );
    not g1044 ( n4522 , n11434 );
    and g1045 ( n12418 , n4028 , n6851 );
    nor g1046 ( n1517 , n13185 , n10309 );
    nor g1047 ( n9526 , n6898 , n6027 );
    and g1048 ( n3846 , n7827 , n10549 );
    not g1049 ( n2816 , n10642 );
    not g1050 ( n4301 , n6639 );
    xnor g1051 ( n12936 , n10593 , n5576 );
    and g1052 ( n12828 , n1982 , n11488 );
    xnor g1053 ( n11428 , n4995 , n7551 );
    nor g1054 ( n12860 , n4711 , n10787 );
    xnor g1055 ( n6470 , n7745 , n3844 );
    and g1056 ( n705 , n564 , n9596 );
    nor g1057 ( n900 , n8947 , n12176 );
    or g1058 ( n13123 , n12432 , n3417 );
    not g1059 ( n8632 , n6668 );
    or g1060 ( n4575 , n9426 , n3053 );
    and g1061 ( n6653 , n798 , n8331 );
    not g1062 ( n12240 , n3472 );
    xor g1063 ( n216 , n1472 , n2652 );
    not g1064 ( n8809 , n10126 );
    xnor g1065 ( n5902 , n6401 , n9798 );
    or g1066 ( n6376 , n6131 , n9757 );
    or g1067 ( n4317 , n13154 , n12273 );
    or g1068 ( n10110 , n2183 , n6635 );
    nor g1069 ( n2815 , n6248 , n8968 );
    not g1070 ( n10293 , n6536 );
    not g1071 ( n10975 , n9616 );
    xnor g1072 ( n5570 , n3002 , n8698 );
    not g1073 ( n712 , n865 );
    and g1074 ( n9582 , n8502 , n5720 );
    or g1075 ( n2434 , n1447 , n206 );
    and g1076 ( n10165 , n6847 , n8994 );
    or g1077 ( n6992 , n8169 , n10407 );
    xnor g1078 ( n12209 , n10110 , n11195 );
    xnor g1079 ( n2384 , n5013 , n12238 );
    or g1080 ( n8662 , n8280 , n11016 );
    or g1081 ( n2046 , n10421 , n7935 );
    or g1082 ( n11967 , n10469 , n4404 );
    and g1083 ( n1754 , n9424 , n6619 );
    not g1084 ( n11677 , n6765 );
    and g1085 ( n6791 , n8236 , n3184 );
    and g1086 ( n13147 , n6668 , n5729 );
    xnor g1087 ( n11892 , n8316 , n12353 );
    or g1088 ( n100 , n444 , n3383 );
    not g1089 ( n6056 , n10142 );
    or g1090 ( n12635 , n8436 , n1155 );
    and g1091 ( n6038 , n4513 , n3309 );
    xnor g1092 ( n12540 , n6354 , n8707 );
    not g1093 ( n5742 , n4348 );
    xnor g1094 ( n10124 , n4048 , n827 );
    and g1095 ( n11670 , n3304 , n4916 );
    nor g1096 ( n3590 , n11925 , n11342 );
    not g1097 ( n161 , n7974 );
    xnor g1098 ( n4510 , n2036 , n5925 );
    or g1099 ( n6918 , n8294 , n10685 );
    or g1100 ( n2523 , n5105 , n11772 );
    not g1101 ( n1908 , n11454 );
    and g1102 ( n12854 , n4975 , n10520 );
    nor g1103 ( n10854 , n10933 , n10799 );
    xnor g1104 ( n3451 , n10405 , n7393 );
    not g1105 ( n2738 , n3815 );
    not g1106 ( n10795 , n10002 );
    or g1107 ( n12737 , n11810 , n8268 );
    nor g1108 ( n6849 , n10356 , n8809 );
    not g1109 ( n1688 , n8522 );
    nor g1110 ( n2521 , n2826 , n10965 );
    and g1111 ( n1242 , n7907 , n10108 );
    and g1112 ( n9993 , n1364 , n124 );
    nor g1113 ( n3943 , n10273 , n5198 );
    or g1114 ( n8547 , n6399 , n5063 );
    not g1115 ( n12032 , n817 );
    and g1116 ( n6278 , n3926 , n11203 );
    and g1117 ( n1814 , n8707 , n6354 );
    or g1118 ( n8460 , n11457 , n5349 );
    xnor g1119 ( n9766 , n9881 , n1740 );
    xnor g1120 ( n9262 , n12181 , n12130 );
    not g1121 ( n11838 , n4312 );
    and g1122 ( n4245 , n2763 , n9366 );
    xnor g1123 ( n8953 , n2465 , n11615 );
    nor g1124 ( n8796 , n4685 , n1045 );
    not g1125 ( n13073 , n7982 );
    or g1126 ( n12196 , n4731 , n210 );
    xnor g1127 ( n1425 , n10857 , n4577 );
    xnor g1128 ( n5553 , n9895 , n384 );
    or g1129 ( n8421 , n8450 , n5669 );
    not g1130 ( n8329 , n6843 );
    not g1131 ( n2772 , n6822 );
    xnor g1132 ( n11089 , n7901 , n8955 );
    nor g1133 ( n7048 , n1766 , n1358 );
    and g1134 ( n9639 , n13201 , n5548 );
    xnor g1135 ( n9294 , n6636 , n1660 );
    xnor g1136 ( n8842 , n7842 , n6147 );
    or g1137 ( n11847 , n6229 , n1417 );
    not g1138 ( n6267 , n1203 );
    or g1139 ( n3300 , n4612 , n3949 );
    or g1140 ( n12597 , n8356 , n8918 );
    xnor g1141 ( n8136 , n6535 , n4064 );
    and g1142 ( n8226 , n240 , n8734 );
    nor g1143 ( n9057 , n6478 , n11678 );
    xnor g1144 ( n8823 , n4571 , n3823 );
    nor g1145 ( n5910 , n3561 , n12830 );
    not g1146 ( n652 , n9093 );
    not g1147 ( n9375 , n3876 );
    not g1148 ( n8297 , n10728 );
    nor g1149 ( n3272 , n11570 , n4239 );
    xnor g1150 ( n348 , n8539 , n2293 );
    not g1151 ( n64 , n6087 );
    and g1152 ( n9303 , n10113 , n10451 );
    not g1153 ( n2122 , n8399 );
    not g1154 ( n9010 , n469 );
    xnor g1155 ( n4858 , n9959 , n8896 );
    nor g1156 ( n688 , n10327 , n6711 );
    and g1157 ( n10215 , n9748 , n12895 );
    xnor g1158 ( n1182 , n7934 , n289 );
    or g1159 ( n110 , n9273 , n9686 );
    nor g1160 ( n10072 , n11930 , n3924 );
    and g1161 ( n4770 , n10872 , n12308 );
    xor g1162 ( n7208 , n828 , n5483 );
    and g1163 ( n1190 , n1952 , n2601 );
    and g1164 ( n9273 , n2496 , n4988 );
    not g1165 ( n5802 , n1874 );
    not g1166 ( n12370 , n6897 );
    or g1167 ( n4525 , n9917 , n10049 );
    or g1168 ( n1562 , n7794 , n7563 );
    and g1169 ( n10532 , n626 , n7887 );
    not g1170 ( n6306 , n2590 );
    not g1171 ( n9182 , n11280 );
    and g1172 ( n1823 , n10984 , n3404 );
    not g1173 ( n118 , n13192 );
    and g1174 ( n12029 , n1259 , n297 );
    and g1175 ( n6058 , n2604 , n12358 );
    or g1176 ( n5180 , n7146 , n5076 );
    xnor g1177 ( n2454 , n1517 , n430 );
    nor g1178 ( n3237 , n10643 , n3633 );
    and g1179 ( n2794 , n9788 , n9989 );
    xnor g1180 ( n12410 , n3321 , n10190 );
    not g1181 ( n8058 , n5304 );
    and g1182 ( n851 , n5491 , n10171 );
    not g1183 ( n6579 , n6226 );
    and g1184 ( n7339 , n4608 , n1918 );
    not g1185 ( n12170 , n7813 );
    or g1186 ( n5004 , n1436 , n4640 );
    or g1187 ( n11900 , n12033 , n4416 );
    and g1188 ( n1833 , n13112 , n12851 );
    xnor g1189 ( n9840 , n12528 , n2694 );
    and g1190 ( n11760 , n2003 , n9237 );
    nor g1191 ( n12880 , n1896 , n11005 );
    xnor g1192 ( n6754 , n8272 , n11062 );
    or g1193 ( n701 , n3682 , n7013 );
    nor g1194 ( n7402 , n10444 , n8586 );
    xor g1195 ( n4171 , n7969 , n6433 );
    xnor g1196 ( n12463 , n1192 , n13029 );
    xnor g1197 ( n3283 , n9067 , n7341 );
    or g1198 ( n11560 , n7247 , n2228 );
    not g1199 ( n11740 , n8358 );
    not g1200 ( n11431 , n12428 );
    not g1201 ( n10893 , n2758 );
    and g1202 ( n7502 , n11322 , n11662 );
    not g1203 ( n6486 , n1231 );
    or g1204 ( n4225 , n6051 , n11998 );
    and g1205 ( n8980 , n7052 , n2219 );
    xor g1206 ( n4957 , n2540 , n9013 );
    xnor g1207 ( n4999 , n3909 , n698 );
    not g1208 ( n12995 , n441 );
    or g1209 ( n1729 , n12551 , n5781 );
    or g1210 ( n4334 , n12997 , n2133 );
    nor g1211 ( n8641 , n9734 , n8523 );
    or g1212 ( n4446 , n3416 , n4474 );
    nor g1213 ( n2399 , n668 , n6663 );
    or g1214 ( n3539 , n5656 , n11538 );
    not g1215 ( n3671 , n5684 );
    not g1216 ( n11869 , n6515 );
    xnor g1217 ( n699 , n11859 , n6877 );
    not g1218 ( n7421 , n4572 );
    nor g1219 ( n7071 , n374 , n5225 );
    nor g1220 ( n12454 , n5509 , n12875 );
    not g1221 ( n1008 , n8932 );
    xnor g1222 ( n10648 , n2973 , n5646 );
    or g1223 ( n12656 , n559 , n4947 );
    or g1224 ( n11197 , n12602 , n3902 );
    xnor g1225 ( n7111 , n2212 , n9768 );
    not g1226 ( n13182 , n9669 );
    and g1227 ( n10052 , n9172 , n4231 );
    and g1228 ( n3294 , n6744 , n347 );
    xnor g1229 ( n8398 , n5530 , n2138 );
    xnor g1230 ( n1568 , n5636 , n152 );
    xnor g1231 ( n1489 , n1657 , n2828 );
    xnor g1232 ( n9336 , n1465 , n12973 );
    xnor g1233 ( n2237 , n12897 , n10216 );
    and g1234 ( n11565 , n10908 , n854 );
    and g1235 ( n12320 , n5964 , n2270 );
    and g1236 ( n4191 , n2937 , n10812 );
    and g1237 ( n11632 , n10809 , n4342 );
    xnor g1238 ( n5701 , n2474 , n12017 );
    xnor g1239 ( n7465 , n3024 , n2119 );
    xnor g1240 ( n368 , n12410 , n1027 );
    and g1241 ( n259 , n2806 , n2189 );
    or g1242 ( n2479 , n4792 , n3454 );
    xnor g1243 ( n3875 , n12269 , n1519 );
    xnor g1244 ( n12554 , n10450 , n5201 );
    not g1245 ( n2550 , n471 );
    xnor g1246 ( n5281 , n10806 , n5977 );
    xnor g1247 ( n11448 , n282 , n8916 );
    xnor g1248 ( n4125 , n3869 , n8717 );
    or g1249 ( n7537 , n4370 , n6635 );
    and g1250 ( n346 , n1647 , n4402 );
    or g1251 ( n12705 , n3024 , n2119 );
    or g1252 ( n12070 , n9968 , n9850 );
    or g1253 ( n10912 , n628 , n10106 );
    or g1254 ( n4010 , n11664 , n9795 );
    or g1255 ( n4235 , n12093 , n12847 );
    and g1256 ( n5623 , n7538 , n2782 );
    not g1257 ( n6811 , n4387 );
    or g1258 ( n8734 , n4251 , n3079 );
    or g1259 ( n10183 , n8053 , n2675 );
    not g1260 ( n10051 , n3298 );
    nor g1261 ( n8338 , n1375 , n12097 );
    or g1262 ( n1372 , n6904 , n5915 );
    not g1263 ( n3555 , n9188 );
    and g1264 ( n4492 , n11318 , n8880 );
    and g1265 ( n12900 , n5252 , n2573 );
    xnor g1266 ( n7599 , n11193 , n6705 );
    nor g1267 ( n8415 , n9790 , n10831 );
    and g1268 ( n7722 , n6333 , n834 );
    not g1269 ( n9622 , n6392 );
    xnor g1270 ( n728 , n3271 , n1776 );
    or g1271 ( n5129 , n8969 , n9141 );
    xnor g1272 ( n228 , n5725 , n5928 );
    xnor g1273 ( n10763 , n149 , n6773 );
    xnor g1274 ( n6784 , n4359 , n12775 );
    or g1275 ( n4104 , n1567 , n12400 );
    or g1276 ( n1048 , n9675 , n6265 );
    xnor g1277 ( n12199 , n8891 , n3182 );
    or g1278 ( n1158 , n3225 , n6265 );
    not g1279 ( n9537 , n11324 );
    or g1280 ( n2388 , n4732 , n4230 );
    xnor g1281 ( n12173 , n4000 , n8477 );
    or g1282 ( n7542 , n11087 , n2449 );
    not g1283 ( n7184 , n12579 );
    or g1284 ( n5589 , n7085 , n1781 );
    xnor g1285 ( n587 , n6572 , n6546 );
    not g1286 ( n11452 , n5174 );
    or g1287 ( n9366 , n11335 , n2123 );
    and g1288 ( n13087 , n13243 , n7003 );
    and g1289 ( n9572 , n12877 , n12288 );
    nor g1290 ( n7548 , n10477 , n8965 );
    buf g1291 ( n2449 , n10240 );
    xnor g1292 ( n5386 , n6887 , n13024 );
    or g1293 ( n4108 , n13117 , n10871 );
    and g1294 ( n9905 , n420 , n1798 );
    and g1295 ( n575 , n8067 , n10817 );
    or g1296 ( n11909 , n334 , n12948 );
    or g1297 ( n8972 , n10761 , n1570 );
    and g1298 ( n9203 , n4099 , n10691 );
    or g1299 ( n5526 , n2195 , n3523 );
    nor g1300 ( n11135 , n6195 , n1900 );
    xnor g1301 ( n9610 , n2992 , n1336 );
    and g1302 ( n6377 , n8688 , n548 );
    not g1303 ( n8453 , n7165 );
    or g1304 ( n13138 , n10756 , n9195 );
    xnor g1305 ( n10001 , n3822 , n1613 );
    and g1306 ( n2092 , n7339 , n5695 );
    nor g1307 ( n11644 , n11881 , n9535 );
    xor g1308 ( n7968 , n9705 , n12101 );
    or g1309 ( n10341 , n1113 , n1144 );
    xnor g1310 ( n5609 , n5914 , n12729 );
    nor g1311 ( n10239 , n279 , n11338 );
    not g1312 ( n4694 , n1543 );
    and g1313 ( n3653 , n6188 , n12922 );
    and g1314 ( n1996 , n5711 , n5085 );
    xnor g1315 ( n301 , n1617 , n5596 );
    xnor g1316 ( n5404 , n528 , n5870 );
    xnor g1317 ( n10356 , n1553 , n7964 );
    not g1318 ( n4589 , n6601 );
    nor g1319 ( n1095 , n4197 , n4697 );
    and g1320 ( n3443 , n11608 , n7657 );
    xnor g1321 ( n1637 , n2242 , n9073 );
    or g1322 ( n9733 , n1983 , n6255 );
    not g1323 ( n9228 , n10162 );
    not g1324 ( n10757 , n2703 );
    or g1325 ( n8410 , n9622 , n4420 );
    xnor g1326 ( n2288 , n6902 , n10750 );
    or g1327 ( n2534 , n7981 , n6089 );
    or g1328 ( n8801 , n2919 , n12388 );
    and g1329 ( n9590 , n6423 , n593 );
    or g1330 ( n12689 , n6206 , n11097 );
    not g1331 ( n6313 , n11993 );
    or g1332 ( n7917 , n5949 , n6635 );
    not g1333 ( n10198 , n9943 );
    or g1334 ( n929 , n4334 , n1777 );
    or g1335 ( n2355 , n8994 , n6847 );
    or g1336 ( n5155 , n4418 , n6926 );
    not g1337 ( n12841 , n9475 );
    and g1338 ( n3019 , n2162 , n4678 );
    xnor g1339 ( n7936 , n12085 , n2071 );
    or g1340 ( n6428 , n4809 , n3632 );
    xnor g1341 ( n8967 , n3625 , n6871 );
    nor g1342 ( n6527 , n11743 , n12727 );
    and g1343 ( n12622 , n2266 , n3743 );
    or g1344 ( n2993 , n11120 , n5885 );
    not g1345 ( n7708 , n7585 );
    xnor g1346 ( n8345 , n1735 , n10164 );
    or g1347 ( n12548 , n12141 , n10513 );
    xnor g1348 ( n4394 , n5445 , n5681 );
    xnor g1349 ( n4380 , n10186 , n8151 );
    not g1350 ( n3468 , n10150 );
    xor g1351 ( n8803 , n7128 , n4078 );
    xnor g1352 ( n9027 , n3833 , n3754 );
    or g1353 ( n298 , n3821 , n12755 );
    and g1354 ( n4223 , n5510 , n5795 );
    xnor g1355 ( n4271 , n5762 , n2501 );
    not g1356 ( n9209 , n9843 );
    and g1357 ( n5315 , n8668 , n8381 );
    xnor g1358 ( n6536 , n9831 , n11025 );
    or g1359 ( n9900 , n2613 , n12233 );
    nor g1360 ( n10031 , n4713 , n11441 );
    nor g1361 ( n10431 , n2167 , n7535 );
    or g1362 ( n949 , n7675 , n9195 );
    not g1363 ( n10045 , n3076 );
    xnor g1364 ( n2683 , n1400 , n9513 );
    nor g1365 ( n7976 , n11131 , n1137 );
    and g1366 ( n6162 , n5867 , n8088 );
    and g1367 ( n2907 , n8816 , n11999 );
    not g1368 ( n3587 , n1084 );
    xnor g1369 ( n3138 , n1009 , n3678 );
    and g1370 ( n5190 , n2903 , n8803 );
    and g1371 ( n4703 , n11324 , n1724 );
    xnor g1372 ( n11865 , n8551 , n1249 );
    nor g1373 ( n7338 , n11095 , n6390 );
    xnor g1374 ( n2895 , n1975 , n356 );
    or g1375 ( n5989 , n644 , n542 );
    xor g1376 ( n12820 , n8600 , n3137 );
    nor g1377 ( n1643 , n2817 , n1299 );
    or g1378 ( n3004 , n4313 , n3487 );
    nor g1379 ( n4012 , n1223 , n7673 );
    not g1380 ( n63 , n9531 );
    and g1381 ( n13093 , n7276 , n3106 );
    not g1382 ( n4866 , n2038 );
    and g1383 ( n5791 , n5371 , n3097 );
    xnor g1384 ( n3503 , n1607 , n2745 );
    or g1385 ( n5863 , n3408 , n11086 );
    not g1386 ( n12718 , n11537 );
    or g1387 ( n1210 , n1072 , n2851 );
    or g1388 ( n4940 , n11269 , n8196 );
    or g1389 ( n4205 , n4612 , n8563 );
    xnor g1390 ( n10572 , n12419 , n3196 );
    or g1391 ( n5416 , n4668 , n12726 );
    xnor g1392 ( n2968 , n374 , n11992 );
    not g1393 ( n4185 , n9887 );
    or g1394 ( n10712 , n1571 , n6265 );
    nor g1395 ( n3673 , n1752 , n11106 );
    not g1396 ( n7001 , n8273 );
    not g1397 ( n11185 , n1278 );
    xnor g1398 ( n4296 , n6118 , n1229 );
    xnor g1399 ( n9230 , n10412 , n4031 );
    nor g1400 ( n8990 , n3874 , n7198 );
    not g1401 ( n3729 , n7238 );
    xnor g1402 ( n8501 , n8289 , n1502 );
    and g1403 ( n1418 , n9942 , n890 );
    nor g1404 ( n7621 , n8632 , n9913 );
    xnor g1405 ( n7774 , n5642 , n4422 );
    or g1406 ( n6372 , n10761 , n6404 );
    and g1407 ( n8685 , n4878 , n10141 );
    and g1408 ( n1704 , n519 , n11896 );
    xnor g1409 ( n9856 , n5093 , n2506 );
    not g1410 ( n11922 , n1923 );
    xnor g1411 ( n3710 , n4192 , n7114 );
    xnor g1412 ( n6373 , n7101 , n1132 );
    and g1413 ( n11415 , n470 , n8370 );
    not g1414 ( n8174 , n11835 );
    xnor g1415 ( n8604 , n99 , n10416 );
    and g1416 ( n309 , n11876 , n1657 );
    or g1417 ( n9781 , n3478 , n5537 );
    not g1418 ( n9829 , n3894 );
    or g1419 ( n12175 , n8757 , n6404 );
    and g1420 ( n4673 , n1184 , n11188 );
    xor g1421 ( n4252 , n959 , n4758 );
    or g1422 ( n8448 , n10448 , n5076 );
    or g1423 ( n8625 , n4208 , n1144 );
    xnor g1424 ( n10396 , n6651 , n9657 );
    xnor g1425 ( n9128 , n7581 , n9973 );
    or g1426 ( n896 , n9225 , n3023 );
    or g1427 ( n7095 , n5019 , n6141 );
    nor g1428 ( n4966 , n1549 , n5753 );
    xnor g1429 ( n472 , n12133 , n7595 );
    or g1430 ( n3848 , n4272 , n5797 );
    xnor g1431 ( n3806 , n1178 , n10489 );
    or g1432 ( n3592 , n3096 , n542 );
    or g1433 ( n6667 , n1968 , n12745 );
    and g1434 ( n2732 , n1160 , n2446 );
    or g1435 ( n7894 , n9911 , n1843 );
    not g1436 ( n1954 , n10398 );
    xnor g1437 ( n12148 , n12172 , n5223 );
    and g1438 ( n11582 , n12904 , n12427 );
    and g1439 ( n1139 , n9901 , n11801 );
    or g1440 ( n10129 , n7934 , n289 );
    not g1441 ( n11227 , n6868 );
    xnor g1442 ( n6161 , n7978 , n1129 );
    and g1443 ( n3376 , n8873 , n4804 );
    not g1444 ( n10085 , n5969 );
    and g1445 ( n4110 , n2223 , n4706 );
    not g1446 ( n10425 , n727 );
    xor g1447 ( n4707 , n9776 , n4037 );
    or g1448 ( n10637 , n2463 , n10871 );
    not g1449 ( n5016 , n10563 );
    not g1450 ( n5328 , n9747 );
    and g1451 ( n9168 , n5671 , n3769 );
    or g1452 ( n1265 , n13170 , n12388 );
    not g1453 ( n7242 , n6195 );
    xnor g1454 ( n1660 , n11272 , n10087 );
    and g1455 ( n10479 , n12673 , n7761 );
    and g1456 ( n8083 , n3647 , n5098 );
    xnor g1457 ( n8147 , n12389 , n6138 );
    xnor g1458 ( n7426 , n12817 , n12872 );
    or g1459 ( n155 , n652 , n2544 );
    nor g1460 ( n5887 , n6425 , n13091 );
    xnor g1461 ( n12502 , n11392 , n9760 );
    and g1462 ( n2229 , n7715 , n12306 );
    not g1463 ( n10927 , n5334 );
    xnor g1464 ( n10548 , n9270 , n2422 );
    and g1465 ( n6204 , n8040 , n7464 );
    or g1466 ( n12805 , n10641 , n11152 );
    and g1467 ( n8587 , n5601 , n10265 );
    or g1468 ( n4401 , n6304 , n539 );
    and g1469 ( n10819 , n7609 , n11924 );
    and g1470 ( n2648 , n9464 , n9191 );
    xnor g1471 ( n6158 , n3526 , n350 );
    and g1472 ( n6833 , n5517 , n12559 );
    or g1473 ( n303 , n2091 , n3597 );
    xnor g1474 ( n9079 , n7406 , n1182 );
    and g1475 ( n13240 , n698 , n3909 );
    nor g1476 ( n6289 , n6893 , n948 );
    xnor g1477 ( n13230 , n10496 , n5159 );
    or g1478 ( n2425 , n9089 , n7760 );
    not g1479 ( n9305 , n5189 );
    xnor g1480 ( n11592 , n3105 , n6410 );
    xnor g1481 ( n3093 , n7438 , n3732 );
    xnor g1482 ( n10887 , n7448 , n194 );
    and g1483 ( n1024 , n2057 , n834 );
    and g1484 ( n8542 , n8228 , n411 );
    not g1485 ( n8951 , n486 );
    nor g1486 ( n2532 , n293 , n7150 );
    not g1487 ( n11806 , n9376 );
    xnor g1488 ( n11243 , n9365 , n636 );
    xor g1489 ( n9666 , n7208 , n11846 );
    or g1490 ( n4288 , n3000 , n9971 );
    and g1491 ( n12875 , n4725 , n2265 );
    or g1492 ( n10607 , n8922 , n5389 );
    xnor g1493 ( n2054 , n8990 , n3675 );
    not g1494 ( n11509 , n4441 );
    xnor g1495 ( n798 , n217 , n3889 );
    and g1496 ( n4091 , n953 , n8107 );
    nor g1497 ( n10007 , n1564 , n512 );
    not g1498 ( n8729 , n7411 );
    not g1499 ( n6808 , n323 );
    nor g1500 ( n12757 , n9958 , n3719 );
    nor g1501 ( n9022 , n12974 , n11587 );
    nor g1502 ( n2004 , n3484 , n13189 );
    xnor g1503 ( n8611 , n11383 , n8396 );
    or g1504 ( n4316 , n5461 , n2449 );
    xnor g1505 ( n648 , n10568 , n12520 );
    or g1506 ( n9438 , n11370 , n5797 );
    or g1507 ( n4521 , n7626 , n5340 );
    not g1508 ( n7522 , n2737 );
    or g1509 ( n13001 , n5218 , n496 );
    not g1510 ( n12721 , n3130 );
    or g1511 ( n12455 , n18 , n11668 );
    xor g1512 ( n790 , n7537 , n3211 );
    xnor g1513 ( n9394 , n9364 , n10058 );
    xnor g1514 ( n5699 , n11312 , n7812 );
    or g1515 ( n11501 , n11037 , n2059 );
    or g1516 ( n5350 , n12150 , n4145 );
    xnor g1517 ( n13004 , n5720 , n8502 );
    xnor g1518 ( n4806 , n9894 , n5210 );
    xnor g1519 ( n3161 , n4834 , n11934 );
    xnor g1520 ( n2309 , n8362 , n4011 );
    xnor g1521 ( n4019 , n4941 , n2628 );
    or g1522 ( n9044 , n6003 , n10579 );
    not g1523 ( n9651 , n10709 );
    and g1524 ( n5373 , n3557 , n6742 );
    xnor g1525 ( n11923 , n5778 , n2381 );
    and g1526 ( n11508 , n4398 , n8997 );
    xnor g1527 ( n8894 , n6273 , n12144 );
    xnor g1528 ( n1576 , n10620 , n1569 );
    not g1529 ( n4144 , n4470 );
    and g1530 ( n3775 , n9888 , n6394 );
    xnor g1531 ( n9103 , n7012 , n1160 );
    xnor g1532 ( n12059 , n7324 , n7996 );
    not g1533 ( n10755 , n6196 );
    and g1534 ( n12701 , n2268 , n3245 );
    and g1535 ( n8992 , n1871 , n2710 );
    xnor g1536 ( n10729 , n8922 , n11759 );
    and g1537 ( n6919 , n5212 , n6802 );
    xnor g1538 ( n4991 , n10766 , n2078 );
    not g1539 ( n13025 , n443 );
    not g1540 ( n227 , n8290 );
    or g1541 ( n9330 , n1340 , n8435 );
    nor g1542 ( n3220 , n10344 , n266 );
    not g1543 ( n10433 , n9620 );
    nor g1544 ( n2208 , n3218 , n6437 );
    and g1545 ( n6394 , n8940 , n6392 );
    xnor g1546 ( n9358 , n5479 , n2951 );
    or g1547 ( n5094 , n6680 , n7306 );
    or g1548 ( n10335 , n7184 , n8268 );
    xnor g1549 ( n8191 , n6499 , n7343 );
    xnor g1550 ( n4299 , n5941 , n4972 );
    xnor g1551 ( n2143 , n5585 , n8092 );
    xnor g1552 ( n4902 , n1454 , n9185 );
    or g1553 ( n3636 , n569 , n9195 );
    or g1554 ( n12699 , n10830 , n6732 );
    not g1555 ( n10764 , n10408 );
    not g1556 ( n10644 , n12550 );
    xnor g1557 ( n4214 , n6898 , n10146 );
    and g1558 ( n5149 , n9980 , n11424 );
    and g1559 ( n8319 , n9217 , n3688 );
    and g1560 ( n2621 , n7240 , n1528 );
    and g1561 ( n2112 , n190 , n12063 );
    or g1562 ( n9297 , n10781 , n8268 );
    nor g1563 ( n5573 , n4550 , n3968 );
    or g1564 ( n13127 , n9476 , n3772 );
    or g1565 ( n5608 , n2802 , n12410 );
    not g1566 ( n558 , n212 );
    or g1567 ( n11654 , n584 , n10029 );
    xnor g1568 ( n9947 , n1393 , n5442 );
    and g1569 ( n3230 , n12976 , n4533 );
    or g1570 ( n1586 , n8480 , n10012 );
    xnor g1571 ( n4803 , n5358 , n7027 );
    nor g1572 ( n10377 , n10115 , n9799 );
    xnor g1573 ( n12248 , n8842 , n5984 );
    or g1574 ( n7571 , n4657 , n10179 );
    and g1575 ( n760 , n9878 , n3030 );
    nor g1576 ( n5443 , n7454 , n7099 );
    or g1577 ( n2261 , n13012 , n11107 );
    nor g1578 ( n5507 , n12593 , n350 );
    not g1579 ( n10211 , n12356 );
    nor g1580 ( n911 , n8135 , n6822 );
    nor g1581 ( n6258 , n7460 , n4450 );
    xnor g1582 ( n2060 , n1864 , n10712 );
    and g1583 ( n4840 , n12378 , n11059 );
    xnor g1584 ( n12125 , n8284 , n4543 );
    xnor g1585 ( n11932 , n9206 , n2645 );
    xnor g1586 ( n8379 , n9948 , n6288 );
    not g1587 ( n816 , n8071 );
    and g1588 ( n3939 , n9710 , n11846 );
    or g1589 ( n2326 , n11492 , n8711 );
    not g1590 ( n8413 , n7376 );
    xnor g1591 ( n8674 , n2442 , n8634 );
    or g1592 ( n12799 , n3003 , n4662 );
    not g1593 ( n4352 , n6085 );
    xnor g1594 ( n5574 , n2786 , n669 );
    or g1595 ( n1490 , n2556 , n4230 );
    xnor g1596 ( n10592 , n1131 , n8192 );
    nor g1597 ( n324 , n6396 , n11425 );
    and g1598 ( n13044 , n9966 , n4720 );
    or g1599 ( n10503 , n5847 , n7515 );
    and g1600 ( n9568 , n5921 , n8571 );
    not g1601 ( n8655 , n1626 );
    not g1602 ( n5973 , n12284 );
    and g1603 ( n5708 , n6580 , n8942 );
    not g1604 ( n6519 , n2339 );
    xnor g1605 ( n7592 , n1763 , n5132 );
    xnor g1606 ( n9516 , n8979 , n10320 );
    and g1607 ( n9757 , n2427 , n2178 );
    not g1608 ( n4530 , n832 );
    and g1609 ( n11311 , n2736 , n2659 );
    not g1610 ( n2346 , n12579 );
    not g1611 ( n10756 , n3409 );
    or g1612 ( n614 , n1553 , n7964 );
    and g1613 ( n9381 , n9468 , n11919 );
    not g1614 ( n11929 , n9906 );
    or g1615 ( n12122 , n7805 , n2059 );
    nor g1616 ( n11496 , n7114 , n4192 );
    and g1617 ( n8209 , n5275 , n3109 );
    nor g1618 ( n4702 , n7693 , n5977 );
    and g1619 ( n4851 , n11587 , n12974 );
    and g1620 ( n199 , n7026 , n10964 );
    or g1621 ( n943 , n3109 , n5275 );
    and g1622 ( n1719 , n11498 , n458 );
    and g1623 ( n3798 , n12788 , n6900 );
    xnor g1624 ( n3603 , n7958 , n2682 );
    nor g1625 ( n5308 , n10538 , n5650 );
    nor g1626 ( n2210 , n7345 , n11613 );
    xnor g1627 ( n4918 , n5110 , n1217 );
    and g1628 ( n8730 , n794 , n2980 );
    nor g1629 ( n7647 , n10666 , n10752 );
    xnor g1630 ( n7408 , n12728 , n9139 );
    and g1631 ( n1130 , n2104 , n10808 );
    xnor g1632 ( n1966 , n6545 , n4131 );
    xnor g1633 ( n4483 , n3007 , n8847 );
    xnor g1634 ( n12691 , n998 , n1399 );
    xnor g1635 ( n8288 , n7938 , n12966 );
    or g1636 ( n2924 , n7152 , n1570 );
    or g1637 ( n9834 , n2204 , n1546 );
    xnor g1638 ( n11477 , n4181 , n11013 );
    or g1639 ( n867 , n8850 , n9907 );
    xor g1640 ( n1401 , n66 , n4111 );
    and g1641 ( n818 , n13173 , n1388 );
    not g1642 ( n2018 , n10866 );
    and g1643 ( n2759 , n10662 , n13027 );
    or g1644 ( n9256 , n1474 , n5450 );
    not g1645 ( n8038 , n2771 );
    xnor g1646 ( n11816 , n10961 , n6552 );
    or g1647 ( n1527 , n6063 , n2544 );
    and g1648 ( n2652 , n5586 , n12263 );
    xnor g1649 ( n2219 , n4574 , n12340 );
    not g1650 ( n12752 , n6032 );
    xnor g1651 ( n8300 , n4648 , n11155 );
    or g1652 ( n8862 , n321 , n3981 );
    and g1653 ( n7871 , n11827 , n9395 );
    and g1654 ( n7929 , n11231 , n9202 );
    or g1655 ( n6125 , n2641 , n6404 );
    and g1656 ( n2539 , n10099 , n10275 );
    or g1657 ( n12402 , n9910 , n9741 );
    and g1658 ( n10545 , n7915 , n5395 );
    nor g1659 ( n10046 , n3238 , n9242 );
    not g1660 ( n7602 , n8822 );
    or g1661 ( n9253 , n4876 , n769 );
    not g1662 ( n10135 , n2758 );
    xnor g1663 ( n4541 , n1928 , n8089 );
    nor g1664 ( n4344 , n3585 , n5779 );
    or g1665 ( n7196 , n5477 , n5174 );
    xnor g1666 ( n6621 , n8976 , n13179 );
    or g1667 ( n11901 , n3892 , n7935 );
    not g1668 ( n8857 , n7116 );
    xnor g1669 ( n9447 , n791 , n2376 );
    or g1670 ( n3556 , n2848 , n479 );
    buf g1671 ( n5076 , n218 );
    nor g1672 ( n2554 , n8272 , n3337 );
    xnor g1673 ( n8197 , n364 , n5178 );
    or g1674 ( n8496 , n9519 , n6541 );
    not g1675 ( n1199 , n12289 );
    nor g1676 ( n12487 , n4797 , n1405 );
    not g1677 ( n6563 , n5284 );
    or g1678 ( n10676 , n11562 , n7335 );
    and g1679 ( n9778 , n12220 , n2100 );
    xnor g1680 ( n11285 , n5945 , n13199 );
    not g1681 ( n111 , n11433 );
    not g1682 ( n3584 , n4630 );
    not g1683 ( n11114 , n10594 );
    xnor g1684 ( n8117 , n7680 , n12818 );
    and g1685 ( n9408 , n10427 , n3424 );
    nor g1686 ( n5931 , n8631 , n9752 );
    xnor g1687 ( n12894 , n3819 , n10295 );
    not g1688 ( n7262 , n4682 );
    or g1689 ( n6975 , n7216 , n8563 );
    or g1690 ( n4639 , n334 , n3225 );
    xnor g1691 ( n2964 , n4475 , n6999 );
    xnor g1692 ( n166 , n7639 , n4327 );
    and g1693 ( n9229 , n5227 , n6391 );
    and g1694 ( n10578 , n9701 , n10457 );
    xnor g1695 ( n12925 , n12777 , n13210 );
    and g1696 ( n5270 , n1757 , n9669 );
    xnor g1697 ( n94 , n6549 , n9167 );
    and g1698 ( n6321 , n7595 , n12133 );
    or g1699 ( n11465 , n5308 , n9379 );
    nor g1700 ( n6521 , n3322 , n4913 );
    xnor g1701 ( n83 , n7376 , n1567 );
    and g1702 ( n589 , n11635 , n3006 );
    nor g1703 ( n6910 , n6471 , n4955 );
    nor g1704 ( n9602 , n5345 , n11727 );
    not g1705 ( n2271 , n1646 );
    xnor g1706 ( n10401 , n5380 , n7417 );
    nor g1707 ( n7920 , n197 , n8785 );
    or g1708 ( n12560 , n4366 , n6635 );
    xnor g1709 ( n6848 , n9700 , n4652 );
    not g1710 ( n6764 , n564 );
    and g1711 ( n3497 , n1739 , n11462 );
    xnor g1712 ( n3472 , n11280 , n8000 );
    not g1713 ( n1012 , n11488 );
    xnor g1714 ( n4973 , n2258 , n4017 );
    and g1715 ( n1153 , n6970 , n4445 );
    not g1716 ( n1973 , n9032 );
    or g1717 ( n5737 , n9310 , n6040 );
    or g1718 ( n8753 , n6004 , n12443 );
    or g1719 ( n462 , n5261 , n5242 );
    or g1720 ( n8545 , n9809 , n1094 );
    and g1721 ( n1161 , n8305 , n9695 );
    or g1722 ( n4137 , n2027 , n6728 );
    and g1723 ( n7307 , n685 , n8068 );
    or g1724 ( n144 , n2381 , n5778 );
    nor g1725 ( n12593 , n3526 , n12933 );
    xnor g1726 ( n5987 , n6531 , n1717 );
    or g1727 ( n3945 , n12376 , n6081 );
    not g1728 ( n694 , n772 );
    not g1729 ( n2681 , n5735 );
    and g1730 ( n3513 , n11419 , n943 );
    xnor g1731 ( n5332 , n3209 , n8721 );
    not g1732 ( n6608 , n1972 );
    xnor g1733 ( n3406 , n12431 , n3782 );
    or g1734 ( n12584 , n8463 , n7306 );
    xnor g1735 ( n11136 , n11935 , n3811 );
    or g1736 ( n8141 , n13159 , n3981 );
    or g1737 ( n7331 , n1398 , n11616 );
    and g1738 ( n12641 , n162 , n8051 );
    and g1739 ( n1157 , n5459 , n5474 );
    xnor g1740 ( n5952 , n8521 , n2577 );
    not g1741 ( n3676 , n937 );
    xnor g1742 ( n8893 , n11379 , n11995 );
    and g1743 ( n5162 , n484 , n7618 );
    nor g1744 ( n13156 , n10583 , n5241 );
    xnor g1745 ( n6246 , n1225 , n8583 );
    xor g1746 ( n11262 , n160 , n6585 );
    or g1747 ( n5988 , n12776 , n11603 );
    not g1748 ( n5264 , n411 );
    and g1749 ( n11576 , n2624 , n5135 );
    xnor g1750 ( n1283 , n10658 , n11579 );
    and g1751 ( n721 , n667 , n5693 );
    and g1752 ( n4017 , n8239 , n12500 );
    xnor g1753 ( n6552 , n8394 , n5310 );
    xnor g1754 ( n9785 , n4717 , n5115 );
    xnor g1755 ( n11409 , n6189 , n5685 );
    or g1756 ( n6113 , n10772 , n4947 );
    and g1757 ( n12219 , n10044 , n1376 );
    nor g1758 ( n5476 , n12885 , n2629 );
    or g1759 ( n10943 , n10761 , n12328 );
    xnor g1760 ( n8477 , n5795 , n5510 );
    or g1761 ( n12001 , n6359 , n6014 );
    not g1762 ( n7306 , n5920 );
    or g1763 ( n7483 , n8609 , n12174 );
    and g1764 ( n6838 , n4186 , n1269 );
    not g1765 ( n2221 , n6392 );
    and g1766 ( n3613 , n1002 , n5390 );
    xnor g1767 ( n11388 , n6811 , n11364 );
    or g1768 ( n12904 , n10279 , n9754 );
    xnor g1769 ( n4292 , n9584 , n7948 );
    not g1770 ( n11485 , n5784 );
    not g1771 ( n6420 , n959 );
    xnor g1772 ( n12261 , n10313 , n1782 );
    and g1773 ( n5584 , n4269 , n8293 );
    and g1774 ( n9397 , n995 , n12970 );
    xnor g1775 ( n12730 , n11669 , n7936 );
    not g1776 ( n3805 , n9915 );
    or g1777 ( n1896 , n12955 , n488 );
    or g1778 ( n4184 , n3963 , n9492 );
    not g1779 ( n1041 , n9508 );
    xor g1780 ( n10973 , n9277 , n6269 );
    and g1781 ( n5809 , n3575 , n2700 );
    nor g1782 ( n9386 , n7426 , n5080 );
    xnor g1783 ( n6022 , n3530 , n5676 );
    not g1784 ( n4442 , n6668 );
    nor g1785 ( n9363 , n10703 , n4905 );
    and g1786 ( n6189 , n1971 , n939 );
    and g1787 ( n7557 , n10426 , n2098 );
    nor g1788 ( n11727 , n1294 , n12975 );
    xnor g1789 ( n942 , n3721 , n4053 );
    and g1790 ( n12430 , n12535 , n2271 );
    and g1791 ( n5726 , n8592 , n8579 );
    and g1792 ( n8789 , n2744 , n12424 );
    not g1793 ( n12885 , n8758 );
    xnor g1794 ( n5322 , n5603 , n1176 );
    and g1795 ( n12787 , n5054 , n1574 );
    not g1796 ( n1696 , n761 );
    not g1797 ( n12009 , n7729 );
    or g1798 ( n11053 , n6451 , n8032 );
    or g1799 ( n7591 , n12767 , n10445 );
    xnor g1800 ( n2814 , n12286 , n113 );
    or g1801 ( n11818 , n7317 , n3261 );
    not g1802 ( n7358 , n3669 );
    xnor g1803 ( n5488 , n6156 , n12403 );
    xnor g1804 ( n7132 , n8822 , n1162 );
    xnor g1805 ( n1755 , n2928 , n3228 );
    xnor g1806 ( n2108 , n11228 , n7529 );
    not g1807 ( n9698 , n11930 );
    xnor g1808 ( n13208 , n9164 , n3256 );
    or g1809 ( n1545 , n10437 , n2544 );
    nor g1810 ( n7454 , n108 , n2892 );
    and g1811 ( n306 , n3070 , n4930 );
    not g1812 ( n3510 , n3974 );
    xnor g1813 ( n3005 , n11718 , n5081 );
    not g1814 ( n1211 , n10186 );
    xnor g1815 ( n3098 , n6813 , n3284 );
    and g1816 ( n1676 , n377 , n6930 );
    and g1817 ( n6863 , n4433 , n9964 );
    and g1818 ( n6247 , n3512 , n5794 );
    not g1819 ( n10244 , n1974 );
    or g1820 ( n11504 , n7033 , n10213 );
    or g1821 ( n11564 , n11192 , n9199 );
    xnor g1822 ( n12245 , n11657 , n10176 );
    or g1823 ( n5821 , n5455 , n4373 );
    nor g1824 ( n10148 , n6525 , n12730 );
    not g1825 ( n7091 , n6763 );
    xnor g1826 ( n4905 , n8442 , n221 );
    not g1827 ( n6360 , n11584 );
    not g1828 ( n12109 , n1165 );
    xnor g1829 ( n11682 , n1090 , n7835 );
    not g1830 ( n7877 , n7281 );
    not g1831 ( n8494 , n7844 );
    xnor g1832 ( n9050 , n4898 , n3028 );
    xnor g1833 ( n4008 , n4496 , n3370 );
    and g1834 ( n3329 , n7156 , n1932 );
    or g1835 ( n3834 , n10883 , n10319 );
    not g1836 ( n1390 , n4135 );
    or g1837 ( n5644 , n1139 , n6216 );
    or g1838 ( n3321 , n6295 , n2637 );
    not g1839 ( n8533 , n3439 );
    and g1840 ( n354 , n9579 , n5233 );
    not g1841 ( n5119 , n7734 );
    or g1842 ( n6444 , n3958 , n2846 );
    not g1843 ( n1737 , n8290 );
    xnor g1844 ( n1014 , n3893 , n1993 );
    and g1845 ( n6385 , n2673 , n5726 );
    or g1846 ( n2298 , n3928 , n10871 );
    nor g1847 ( n12466 , n12864 , n2110 );
    nor g1848 ( n1248 , n8308 , n5214 );
    or g1849 ( n13101 , n1941 , n4640 );
    and g1850 ( n12578 , n8308 , n9669 );
    xnor g1851 ( n1293 , n6738 , n9486 );
    not g1852 ( n2276 , n8183 );
    xnor g1853 ( n2470 , n3654 , n12070 );
    xnor g1854 ( n7038 , n2764 , n4123 );
    not g1855 ( n1508 , n6471 );
    xnor g1856 ( n2176 , n8659 , n9755 );
    not g1857 ( n6419 , n7113 );
    nor g1858 ( n682 , n3695 , n5723 );
    or g1859 ( n830 , n4153 , n10973 );
    or g1860 ( n3240 , n12851 , n13112 );
    nor g1861 ( n5539 , n114 , n10866 );
    xnor g1862 ( n7259 , n13000 , n9753 );
    xnor g1863 ( n8059 , n10326 , n7793 );
    xnor g1864 ( n4082 , n540 , n8760 );
    and g1865 ( n2212 , n7662 , n1006 );
    nor g1866 ( n1981 , n10564 , n7521 );
    and g1867 ( n2151 , n11840 , n12036 );
    nor g1868 ( n2007 , n12716 , n7785 );
    or g1869 ( n12585 , n6801 , n4062 );
    not g1870 ( n192 , n4821 );
    or g1871 ( n5877 , n9159 , n5076 );
    and g1872 ( n2398 , n4456 , n5353 );
    xnor g1873 ( n6740 , n2310 , n7605 );
    and g1874 ( n6389 , n7154 , n8898 );
    xnor g1875 ( n416 , n6104 , n9053 );
    xnor g1876 ( n846 , n7779 , n2482 );
    not g1877 ( n11591 , n854 );
    nor g1878 ( n6042 , n3061 , n13192 );
    or g1879 ( n1212 , n5168 , n10029 );
    not g1880 ( n10780 , n3112 );
    or g1881 ( n10947 , n6303 , n10601 );
    nor g1882 ( n11577 , n12756 , n8557 );
    xnor g1883 ( n5804 , n8919 , n167 );
    not g1884 ( n4741 , n11634 );
    not g1885 ( n3413 , n684 );
    or g1886 ( n2427 , n2357 , n11857 );
    xnor g1887 ( n7919 , n7467 , n1476 );
    and g1888 ( n2731 , n9721 , n7606 );
    or g1889 ( n1148 , n11225 , n4373 );
    or g1890 ( n12412 , n7172 , n11978 );
    and g1891 ( n5074 , n12256 , n10353 );
    xnor g1892 ( n7065 , n4458 , n11083 );
    and g1893 ( n5406 , n11195 , n10110 );
    not g1894 ( n6381 , n9906 );
    and g1895 ( n4920 , n5279 , n10305 );
    xnor g1896 ( n9373 , n4507 , n1342 );
    xnor g1897 ( n2075 , n8420 , n12064 );
    xnor g1898 ( n9688 , n656 , n3685 );
    or g1899 ( n1975 , n7707 , n121 );
    xnor g1900 ( n6185 , n9728 , n11555 );
    not g1901 ( n8532 , n4335 );
    nor g1902 ( n11524 , n1225 , n6716 );
    or g1903 ( n2428 , n7889 , n2685 );
    or g1904 ( n3547 , n3520 , n6377 );
    or g1905 ( n424 , n10256 , n10871 );
    or g1906 ( n11423 , n1571 , n6404 );
    not g1907 ( n218 , n7715 );
    xnor g1908 ( n4656 , n4491 , n7733 );
    xnor g1909 ( n5201 , n9462 , n11795 );
    and g1910 ( n11209 , n2236 , n5774 );
    and g1911 ( n6108 , n4310 , n13205 );
    or g1912 ( n5807 , n9479 , n8883 );
    or g1913 ( n8792 , n10712 , n1864 );
    xnor g1914 ( n10298 , n8288 , n10442 );
    nor g1915 ( n9338 , n8497 , n7400 );
    nor g1916 ( n1861 , n9227 , n9207 );
    xnor g1917 ( n3196 , n790 , n7528 );
    xnor g1918 ( n10365 , n12157 , n6070 );
    not g1919 ( n1732 , n7617 );
    xnor g1920 ( n5731 , n11681 , n13065 );
    or g1921 ( n4061 , n3132 , n5286 );
    and g1922 ( n4165 , n2589 , n12806 );
    or g1923 ( n7413 , n3898 , n3981 );
    nor g1924 ( n4735 , n749 , n7756 );
    xnor g1925 ( n9291 , n4685 , n12443 );
    xnor g1926 ( n11201 , n10070 , n10663 );
    nor g1927 ( n6703 , n13220 , n3232 );
    or g1928 ( n8736 , n13149 , n13113 );
    and g1929 ( n12287 , n2281 , n973 );
    not g1930 ( n6097 , n1718 );
    xnor g1931 ( n988 , n2169 , n8624 );
    xnor g1932 ( n4781 , n3153 , n3806 );
    xnor g1933 ( n7256 , n6523 , n9241 );
    or g1934 ( n641 , n6939 , n9195 );
    xnor g1935 ( n1163 , n2090 , n11305 );
    and g1936 ( n9212 , n677 , n5703 );
    nor g1937 ( n2094 , n11655 , n870 );
    xnor g1938 ( n6021 , n8908 , n8376 );
    nor g1939 ( n1074 , n1746 , n262 );
    or g1940 ( n3466 , n4857 , n3747 );
    not g1941 ( n6749 , n103 );
    not g1942 ( n737 , n8163 );
    and g1943 ( n9968 , n3746 , n10913 );
    not g1944 ( n5401 , n4998 );
    not g1945 ( n6464 , n9705 );
    or g1946 ( n7564 , n2861 , n206 );
    not g1947 ( n5146 , n603 );
    not g1948 ( n3931 , n7455 );
    xnor g1949 ( n217 , n2476 , n10707 );
    or g1950 ( n10710 , n5035 , n859 );
    not g1951 ( n11446 , n411 );
    xnor g1952 ( n6485 , n3888 , n7828 );
    not g1953 ( n12031 , n344 );
    not g1954 ( n6380 , n4773 );
    xnor g1955 ( n11782 , n9640 , n12158 );
    nor g1956 ( n2456 , n6366 , n6871 );
    or g1957 ( n12529 , n1941 , n10106 );
    or g1958 ( n7351 , n8329 , n4724 );
    and g1959 ( n7895 , n5772 , n7899 );
    xnor g1960 ( n5551 , n7426 , n635 );
    xnor g1961 ( n1902 , n7401 , n5852 );
    or g1962 ( n12323 , n6259 , n3461 );
    or g1963 ( n9860 , n3630 , n2675 );
    not g1964 ( n4227 , n502 );
    xnor g1965 ( n12389 , n10608 , n12898 );
    or g1966 ( n2248 , n9679 , n11137 );
    xnor g1967 ( n3378 , n7354 , n501 );
    or g1968 ( n861 , n6388 , n8461 );
    or g1969 ( n2961 , n6568 , n6290 );
    or g1970 ( n2680 , n4128 , n9982 );
    xnor g1971 ( n12260 , n11685 , n6124 );
    or g1972 ( n222 , n3816 , n4682 );
    not g1973 ( n1706 , n10167 );
    and g1974 ( n3012 , n3901 , n12326 );
    and g1975 ( n4543 , n2318 , n12046 );
    or g1976 ( n104 , n9769 , n6044 );
    nor g1977 ( n12194 , n11918 , n6962 );
    and g1978 ( n10842 , n4105 , n9354 );
    xnor g1979 ( n12407 , n10513 , n1550 );
    or g1980 ( n5946 , n4988 , n2496 );
    xnor g1981 ( n9963 , n7811 , n6179 );
    and g1982 ( n1441 , n9040 , n4381 );
    or g1983 ( n3197 , n5018 , n4477 );
    or g1984 ( n11946 , n12394 , n8367 );
    not g1985 ( n9145 , n1641 );
    or g1986 ( n3888 , n7780 , n10871 );
    or g1987 ( n9484 , n628 , n9195 );
    xnor g1988 ( n461 , n10132 , n1779 );
    not g1989 ( n1813 , n6661 );
    and g1990 ( n5723 , n12812 , n602 );
    xnor g1991 ( n213 , n6043 , n12423 );
    nor g1992 ( n2077 , n11261 , n4216 );
    nor g1993 ( n11844 , n7882 , n1923 );
    and g1994 ( n10521 , n6591 , n11385 );
    nor g1995 ( n6304 , n11937 , n2920 );
    xnor g1996 ( n1118 , n7933 , n7244 );
    not g1997 ( n10161 , n2164 );
    or g1998 ( n4274 , n7414 , n8845 );
    or g1999 ( n8138 , n4201 , n2059 );
    and g2000 ( n6064 , n2482 , n6149 );
    xnor g2001 ( n9138 , n2024 , n12006 );
    or g2002 ( n13016 , n3783 , n10818 );
    or g2003 ( n692 , n8062 , n99 );
    xnor g2004 ( n4410 , n10476 , n8809 );
    and g2005 ( n8647 , n3282 , n7196 );
    xnor g2006 ( n3601 , n1766 , n976 );
    and g2007 ( n4002 , n4506 , n3617 );
    not g2008 ( n10476 , n10356 );
    not g2009 ( n9380 , n12820 );
    or g2010 ( n3069 , n1733 , n7079 );
    not g2011 ( n8079 , n9620 );
    not g2012 ( n168 , n6386 );
    and g2013 ( n4089 , n11661 , n9525 );
    xnor g2014 ( n6693 , n8048 , n11210 );
    not g2015 ( n3038 , n5572 );
    xnor g2016 ( n5925 , n2434 , n12854 );
    xnor g2017 ( n8312 , n9347 , n10933 );
    not g2018 ( n2199 , n5336 );
    xnor g2019 ( n3465 , n492 , n5894 );
    or g2020 ( n3778 , n4432 , n6119 );
    nor g2021 ( n6037 , n13226 , n13064 );
    xnor g2022 ( n8772 , n9877 , n7777 );
    and g2023 ( n191 , n8065 , n2157 );
    and g2024 ( n1469 , n4982 , n3652 );
    not g2025 ( n8855 , n1192 );
    xnor g2026 ( n1348 , n3771 , n158 );
    and g2027 ( n7020 , n1504 , n11669 );
    or g2028 ( n12141 , n7291 , n2287 );
    and g2029 ( n3985 , n12620 , n6170 );
    and g2030 ( n9996 , n8486 , n3141 );
    xnor g2031 ( n9165 , n10941 , n7407 );
    xnor g2032 ( n11588 , n7307 , n1818 );
    and g2033 ( n852 , n11869 , n8755 );
    or g2034 ( n11876 , n1377 , n6760 );
    or g2035 ( n5050 , n10923 , n804 );
    and g2036 ( n2281 , n6625 , n9346 );
    nor g2037 ( n9630 , n7225 , n5126 );
    not g2038 ( n559 , n5920 );
    or g2039 ( n1294 , n1051 , n1144 );
    xnor g2040 ( n2435 , n942 , n2084 );
    xnor g2041 ( n6762 , n12124 , n12205 );
    xnor g2042 ( n9842 , n7177 , n12265 );
    xor g2043 ( n5672 , n6365 , n872 );
    not g2044 ( n2542 , n6668 );
    and g2045 ( n4443 , n11427 , n2021 );
    nor g2046 ( n4170 , n7714 , n7338 );
    not g2047 ( n12304 , n5951 );
    or g2048 ( n525 , n8637 , n3686 );
    or g2049 ( n11880 , n5694 , n10319 );
    not g2050 ( n2791 , n9358 );
    xnor g2051 ( n7382 , n3033 , n11207 );
    xnor g2052 ( n9364 , n6202 , n8897 );
    xnor g2053 ( n10653 , n11248 , n5179 );
    nor g2054 ( n5063 , n4242 , n598 );
    or g2055 ( n6035 , n2338 , n10319 );
    xnor g2056 ( n1476 , n3780 , n8685 );
    xnor g2057 ( n9692 , n7051 , n9380 );
    or g2058 ( n8546 , n13159 , n10319 );
    or g2059 ( n1557 , n3791 , n10008 );
    nor g2060 ( n6398 , n226 , n12075 );
    not g2061 ( n9095 , n8330 );
    and g2062 ( n3320 , n1959 , n11139 );
    or g2063 ( n9861 , n8585 , n5076 );
    not g2064 ( n5169 , n2771 );
    nor g2065 ( n5606 , n419 , n6577 );
    xnor g2066 ( n7711 , n50 , n11782 );
    buf g2067 ( n9075 , n16 );
    xnor g2068 ( n8920 , n6804 , n8372 );
    xnor g2069 ( n6460 , n699 , n6798 );
    xnor g2070 ( n7021 , n1123 , n7967 );
    not g2071 ( n5152 , n9093 );
    nor g2072 ( n13008 , n7797 , n5996 );
    not g2073 ( n12882 , n1307 );
    and g2074 ( n6633 , n5017 , n1019 );
    or g2075 ( n8425 , n434 , n3787 );
    xnor g2076 ( n10449 , n1840 , n8844 );
    or g2077 ( n9525 , n10566 , n11877 );
    nor g2078 ( n6573 , n12041 , n2635 );
    xnor g2079 ( n3290 , n4749 , n9044 );
    xnor g2080 ( n6631 , n3288 , n5291 );
    xnor g2081 ( n11516 , n1568 , n11043 );
    nor g2082 ( n2103 , n5799 , n9645 );
    xnor g2083 ( n2866 , n299 , n10773 );
    and g2084 ( n3830 , n5031 , n8233 );
    or g2085 ( n6179 , n5634 , n3981 );
    or g2086 ( n4598 , n8976 , n13179 );
    and g2087 ( n13185 , n1728 , n5551 );
    xnor g2088 ( n6586 , n9381 , n10192 );
    or g2089 ( n3325 , n7393 , n6266 );
    xnor g2090 ( n4106 , n5395 , n11639 );
    or g2091 ( n5799 , n6332 , n6404 );
    not g2092 ( n2701 , n10451 );
    and g2093 ( n1915 , n7149 , n6098 );
    or g2094 ( n5278 , n8095 , n4932 );
    xnor g2095 ( n1488 , n243 , n4863 );
    xnor g2096 ( n12893 , n4802 , n1149 );
    xnor g2097 ( n7596 , n931 , n7543 );
    xnor g2098 ( n2537 , n8357 , n6865 );
    not g2099 ( n7041 , n2339 );
    and g2100 ( n2486 , n1671 , n11642 );
    xnor g2101 ( n10752 , n10651 , n6876 );
    not g2102 ( n2744 , n11096 );
    or g2103 ( n12027 , n9048 , n3635 );
    xnor g2104 ( n13223 , n8407 , n4247 );
    or g2105 ( n3333 , n9962 , n9195 );
    and g2106 ( n1668 , n5799 , n9645 );
    and g2107 ( n550 , n4086 , n6064 );
    nor g2108 ( n4529 , n2908 , n6060 );
    nor g2109 ( n1478 , n4244 , n5961 );
    xnor g2110 ( n10477 , n1507 , n7097 );
    xnor g2111 ( n11778 , n8560 , n5672 );
    not g2112 ( n7977 , n8970 );
    xnor g2113 ( n13042 , n2164 , n7090 );
    or g2114 ( n4441 , n6056 , n12164 );
    or g2115 ( n1150 , n8556 , n10871 );
    xnor g2116 ( n11435 , n9559 , n9704 );
    xnor g2117 ( n4436 , n11526 , n12347 );
    or g2118 ( n11721 , n10603 , n6540 );
    not g2119 ( n6680 , n9732 );
    xnor g2120 ( n4820 , n1185 , n5059 );
    or g2121 ( n8928 , n11379 , n8841 );
    xnor g2122 ( n11159 , n294 , n6648 );
    not g2123 ( n2538 , n10408 );
    or g2124 ( n4040 , n1635 , n1572 );
    xor g2125 ( n2987 , n6487 , n826 );
    not g2126 ( n7371 , n11872 );
    xnor g2127 ( n11837 , n6385 , n2836 );
    nor g2128 ( n10583 , n12790 , n9807 );
    nor g2129 ( n12927 , n6933 , n7562 );
    not g2130 ( n11823 , n1176 );
    and g2131 ( n1486 , n4822 , n830 );
    xor g2132 ( n5454 , n2965 , n6704 );
    not g2133 ( n3301 , n2962 );
    not g2134 ( n10203 , n11201 );
    or g2135 ( n9349 , n2799 , n2451 );
    xnor g2136 ( n4872 , n1351 , n4205 );
    or g2137 ( n9997 , n8720 , n3703 );
    not g2138 ( n1671 , n10547 );
    or g2139 ( n5600 , n11729 , n8348 );
    and g2140 ( n8116 , n265 , n6657 );
    not g2141 ( n438 , n1007 );
    xnor g2142 ( n5398 , n9432 , n9263 );
    or g2143 ( n13110 , n333 , n2222 );
    and g2144 ( n1516 , n1962 , n3685 );
    xnor g2145 ( n6876 , n11070 , n3503 );
    or g2146 ( n5582 , n11094 , n8490 );
    xnor g2147 ( n6948 , n2418 , n2139 );
    or g2148 ( n7794 , n5923 , n7935 );
    nor g2149 ( n9302 , n12719 , n10778 );
    not g2150 ( n7110 , n6574 );
    not g2151 ( n6750 , n2734 );
    and g2152 ( n4971 , n4257 , n12988 );
    and g2153 ( n1566 , n12510 , n619 );
    buf g2154 ( n10871 , n4517 );
    xnor g2155 ( n5578 , n10683 , n12393 );
    not g2156 ( n9702 , n5758 );
    xnor g2157 ( n3476 , n7549 , n3380 );
    or g2158 ( n1313 , n5303 , n2032 );
    and g2159 ( n7032 , n11797 , n12311 );
    or g2160 ( n5370 , n12052 , n6635 );
    and g2161 ( n4020 , n10716 , n9813 );
    and g2162 ( n2246 , n5010 , n8943 );
    or g2163 ( n9494 , n1353 , n1144 );
    xnor g2164 ( n77 , n4007 , n6665 );
    or g2165 ( n10174 , n39 , n3103 );
    not g2166 ( n2028 , n7273 );
    or g2167 ( n11424 , n4558 , n1811 );
    xnor g2168 ( n8110 , n10713 , n1692 );
    xnor g2169 ( n1748 , n12030 , n6748 );
    not g2170 ( n7102 , n12683 );
    or g2171 ( n4497 , n4157 , n4326 );
    not g2172 ( n3031 , n12953 );
    or g2173 ( n240 , n4496 , n1247 );
    xnor g2174 ( n6195 , n3037 , n11390 );
    xnor g2175 ( n11377 , n12633 , n8309 );
    or g2176 ( n4677 , n2598 , n13151 );
    or g2177 ( n12902 , n4372 , n1678 );
    and g2178 ( n11170 , n4719 , n1096 );
    or g2179 ( n12432 , n79 , n4640 );
    nor g2180 ( n4650 , n4624 , n11495 );
    xnor g2181 ( n9551 , n7975 , n7523 );
    and g2182 ( n4415 , n12004 , n7738 );
    and g2183 ( n3549 , n12848 , n9466 );
    and g2184 ( n1595 , n8115 , n11041 );
    xnor g2185 ( n1363 , n7225 , n12359 );
    or g2186 ( n6822 , n367 , n12566 );
    and g2187 ( n8960 , n6402 , n9918 );
    xnor g2188 ( n10164 , n10674 , n6837 );
    or g2189 ( n13216 , n12054 , n5392 );
    or g2190 ( n1494 , n10383 , n7723 );
    or g2191 ( n7792 , n333 , n10956 );
    not g2192 ( n8987 , n5989 );
    xnor g2193 ( n3267 , n4444 , n8589 );
    and g2194 ( n7273 , n13174 , n1596 );
    and g2195 ( n13165 , n5568 , n10451 );
    or g2196 ( n1207 , n11466 , n10106 );
    not g2197 ( n12308 , n7035 );
    and g2198 ( n3298 , n8971 , n8936 );
    nor g2199 ( n7767 , n11828 , n3452 );
    or g2200 ( n2713 , n4291 , n2562 );
    not g2201 ( n12686 , n9124 );
    or g2202 ( n9029 , n2250 , n10701 );
    xnor g2203 ( n6127 , n2829 , n8128 );
    nor g2204 ( n12586 , n1098 , n2311 );
    not g2205 ( n2323 , n10134 );
    not g2206 ( n8912 , n11061 );
    xor g2207 ( n4313 , n7419 , n9619 );
    nor g2208 ( n515 , n4673 , n292 );
    and g2209 ( n3048 , n10026 , n4542 );
    and g2210 ( n897 , n5037 , n9651 );
    xnor g2211 ( n6299 , n8271 , n10626 );
    or g2212 ( n12296 , n9310 , n1571 );
    or g2213 ( n4478 , n13077 , n4640 );
    not g2214 ( n5058 , n11850 );
    not g2215 ( n2930 , n4426 );
    not g2216 ( n8775 , n3365 );
    or g2217 ( n6318 , n4693 , n814 );
    or g2218 ( n5111 , n9614 , n1581 );
    or g2219 ( n8416 , n10476 , n10126 );
    not g2220 ( n10591 , n7720 );
    or g2221 ( n10355 , n1887 , n8348 );
    not g2222 ( n7827 , n3693 );
    and g2223 ( n10615 , n4206 , n9023 );
    not g2224 ( n7878 , n7659 );
    or g2225 ( n6320 , n2377 , n6860 );
    xnor g2226 ( n6350 , n11705 , n4662 );
    xnor g2227 ( n7576 , n966 , n7336 );
    or g2228 ( n4852 , n1096 , n4719 );
    or g2229 ( n8221 , n8487 , n11822 );
    not g2230 ( n159 , n8150 );
    or g2231 ( n2289 , n8904 , n8030 );
    not g2232 ( n5086 , n103 );
    or g2233 ( n12220 , n10591 , n8534 );
    not g2234 ( n115 , n499 );
    xnor g2235 ( n10567 , n7147 , n397 );
    nor g2236 ( n11911 , n5185 , n1734 );
    or g2237 ( n11080 , n2872 , n10029 );
    not g2238 ( n6156 , n3042 );
    xnor g2239 ( n10303 , n13081 , n11263 );
    xnor g2240 ( n9063 , n9188 , n1815 );
    and g2241 ( n3715 , n10783 , n125 );
    not g2242 ( n4816 , n4285 );
    and g2243 ( n2720 , n7493 , n2553 );
    xnor g2244 ( n903 , n8402 , n2783 );
    xnor g2245 ( n7314 , n11486 , n9410 );
    and g2246 ( n11256 , n8161 , n6651 );
    or g2247 ( n3139 , n3572 , n10352 );
    xnor g2248 ( n2475 , n1523 , n6197 );
    or g2249 ( n11420 , n3225 , n6732 );
    xnor g2250 ( n8902 , n1411 , n476 );
    and g2251 ( n11294 , n13201 , n11058 );
    and g2252 ( n7595 , n5031 , n287 );
    and g2253 ( n7820 , n6005 , n1150 );
    or g2254 ( n8799 , n7730 , n650 );
    xnor g2255 ( n11145 , n11423 , n3408 );
    or g2256 ( n9483 , n2321 , n3999 );
    nor g2257 ( n12753 , n7958 , n5864 );
    and g2258 ( n9701 , n9510 , n11525 );
    not g2259 ( n6917 , n745 );
    or g2260 ( n422 , n3284 , n6813 );
    xnor g2261 ( n10395 , n10026 , n9802 );
    or g2262 ( n8487 , n8744 , n4179 );
    xnor g2263 ( n6109 , n2112 , n8501 );
    and g2264 ( n5662 , n10127 , n6645 );
    not g2265 ( n13013 , n937 );
    or g2266 ( n8879 , n11333 , n2942 );
    xnor g2267 ( n9975 , n7702 , n5989 );
    not g2268 ( n13191 , n6948 );
    and g2269 ( n727 , n8406 , n6076 );
    and g2270 ( n11814 , n10304 , n9517 );
    nor g2271 ( n6199 , n3481 , n9338 );
    or g2272 ( n10284 , n2095 , n11810 );
    xnor g2273 ( n11334 , n12696 , n648 );
    or g2274 ( n10979 , n7119 , n12328 );
    or g2275 ( n9328 , n6125 , n9608 );
    or g2276 ( n10845 , n7550 , n9518 );
    and g2277 ( n653 , n2280 , n11102 );
    or g2278 ( n172 , n8843 , n12501 );
    xnor g2279 ( n2750 , n10889 , n4425 );
    or g2280 ( n4921 , n7011 , n7117 );
    or g2281 ( n12262 , n2296 , n10029 );
    not g2282 ( n11593 , n6650 );
    and g2283 ( n71 , n784 , n2433 );
    or g2284 ( n12840 , n6355 , n1696 );
    nor g2285 ( n7364 , n10625 , n10160 );
    xnor g2286 ( n6103 , n4023 , n474 );
    nor g2287 ( n1380 , n2016 , n2050 );
    not g2288 ( n11148 , n4382 );
    xnor g2289 ( n1107 , n1798 , n420 );
    not g2290 ( n10786 , n8675 );
    and g2291 ( n5483 , n3178 , n5548 );
    not g2292 ( n7961 , n1364 );
    or g2293 ( n7403 , n6245 , n3698 );
    xnor g2294 ( n3562 , n8156 , n10170 );
    or g2295 ( n10060 , n6309 , n6037 );
    xnor g2296 ( n945 , n5269 , n4939 );
    and g2297 ( n563 , n7102 , n1054 );
    not g2298 ( n8556 , n12306 );
    xnor g2299 ( n8267 , n5942 , n7334 );
    or g2300 ( n24 , n11536 , n911 );
    xnor g2301 ( n11657 , n11407 , n9550 );
    xnor g2302 ( n6884 , n1854 , n1273 );
    or g2303 ( n9647 , n9557 , n4686 );
    xnor g2304 ( n2000 , n7840 , n9435 );
    xnor g2305 ( n9374 , n5230 , n9636 );
    and g2306 ( n12512 , n998 , n11125 );
    nor g2307 ( n562 , n3929 , n1853 );
    xnor g2308 ( n11206 , n3057 , n10863 );
    or g2309 ( n10541 , n6225 , n5414 );
    and g2310 ( n2969 , n7429 , n9567 );
    nor g2311 ( n11393 , n12143 , n3793 );
    not g2312 ( n8176 , n8768 );
    xnor g2313 ( n6050 , n12451 , n2402 );
    or g2314 ( n1701 , n1278 , n3712 );
    not g2315 ( n11029 , n1876 );
    not g2316 ( n8663 , n10697 );
    xnor g2317 ( n3789 , n502 , n11588 );
    and g2318 ( n9091 , n1584 , n11572 );
    xnor g2319 ( n11879 , n9418 , n1057 );
    not g2320 ( n12568 , n497 );
    not g2321 ( n9383 , n5356 );
    nor g2322 ( n13202 , n6021 , n1186 );
    xnor g2323 ( n9576 , n4239 , n11570 );
    not g2324 ( n759 , n2939 );
    xnor g2325 ( n7892 , n4731 , n5790 );
    not g2326 ( n4606 , n12488 );
    not g2327 ( n10858 , n12609 );
    or g2328 ( n1841 , n2148 , n1043 );
    or g2329 ( n5700 , n10017 , n12388 );
    xnor g2330 ( n2239 , n6799 , n7826 );
    xnor g2331 ( n2913 , n8356 , n456 );
    or g2332 ( n10065 , n2677 , n10912 );
    nor g2333 ( n604 , n6015 , n7602 );
    or g2334 ( n3352 , n3225 , n10900 );
    xnor g2335 ( n7639 , n11791 , n269 );
    xnor g2336 ( n1810 , n9951 , n3495 );
    xnor g2337 ( n4646 , n10537 , n5049 );
    not g2338 ( n549 , n1254 );
    and g2339 ( n4372 , n7821 , n5039 );
    and g2340 ( n6399 , n13000 , n8981 );
    xnor g2341 ( n5972 , n3958 , n2846 );
    not g2342 ( n11940 , n8466 );
    nor g2343 ( n4062 , n10004 , n3358 );
    xnor g2344 ( n381 , n6657 , n265 );
    or g2345 ( n2168 , n7467 , n2249 );
    and g2346 ( n3538 , n12432 , n3417 );
    or g2347 ( n435 , n5767 , n6589 );
    xnor g2348 ( n1162 , n6015 , n1529 );
    not g2349 ( n1067 , n7613 );
    and g2350 ( n8732 , n476 , n1411 );
    or g2351 ( n3045 , n2232 , n6814 );
    not g2352 ( n11291 , n9300 );
    nor g2353 ( n11831 , n214 , n4378 );
    and g2354 ( n2790 , n1212 , n13061 );
    and g2355 ( n10980 , n11130 , n5208 );
    xnor g2356 ( n6459 , n9567 , n7429 );
    xnor g2357 ( n7392 , n2337 , n8277 );
    xnor g2358 ( n5852 , n11343 , n4595 );
    and g2359 ( n3278 , n10582 , n11887 );
    xnor g2360 ( n2029 , n1310 , n5632 );
    or g2361 ( n3260 , n12948 , n6265 );
    and g2362 ( n8597 , n11706 , n1379 );
    and g2363 ( n5020 , n10366 , n10328 );
    and g2364 ( n2127 , n10566 , n11877 );
    or g2365 ( n4704 , n8998 , n12132 );
    xnor g2366 ( n12538 , n13203 , n5487 );
    xnor g2367 ( n10639 , n12313 , n522 );
    and g2368 ( n1247 , n3079 , n4251 );
    not g2369 ( n9119 , n11059 );
    and g2370 ( n7344 , n4668 , n12726 );
    and g2371 ( n12339 , n10860 , n1347 );
    xnor g2372 ( n12265 , n147 , n10094 );
    nor g2373 ( n3654 , n6082 , n12542 );
    or g2374 ( n6802 , n5164 , n7412 );
    xnor g2375 ( n5185 , n4971 , n6597 );
    xnor g2376 ( n5800 , n13184 , n6891 );
    not g2377 ( n2970 , n10642 );
    and g2378 ( n2167 , n11643 , n7378 );
    xnor g2379 ( n345 , n4157 , n2317 );
    not g2380 ( n2551 , n9929 );
    and g2381 ( n12581 , n10530 , n12938 );
    or g2382 ( n2259 , n3940 , n2637 );
    and g2383 ( n2868 , n941 , n12599 );
    or g2384 ( n9552 , n1241 , n11817 );
    not g2385 ( n7424 , n4141 );
    not g2386 ( n935 , n287 );
    and g2387 ( n8677 , n4478 , n1599 );
    not g2388 ( n6756 , n4597 );
    or g2389 ( n4157 , n4077 , n9638 );
    not g2390 ( n7998 , n9475 );
    and g2391 ( n6959 , n12790 , n9807 );
    xnor g2392 ( n3309 , n12567 , n8465 );
    or g2393 ( n4134 , n1125 , n4606 );
    and g2394 ( n8637 , n6739 , n9279 );
    and g2395 ( n5668 , n12592 , n3076 );
    xnor g2396 ( n3389 , n8031 , n4450 );
    and g2397 ( n8032 , n7324 , n6682 );
    xnor g2398 ( n631 , n7298 , n8266 );
    and g2399 ( n5983 , n7195 , n311 );
    not g2400 ( n5766 , n9856 );
    or g2401 ( n3774 , n6407 , n6732 );
    xnor g2402 ( n10207 , n8208 , n3873 );
    and g2403 ( n2564 , n13201 , n9915 );
    or g2404 ( n9725 , n11347 , n824 );
    xnor g2405 ( n6763 , n2335 , n12892 );
    not g2406 ( n1416 , n5320 );
    not g2407 ( n1672 , n5780 );
    xnor g2408 ( n480 , n6701 , n7844 );
    xnor g2409 ( n11440 , n6427 , n5886 );
    or g2410 ( n781 , n7247 , n10059 );
    or g2411 ( n12614 , n1571 , n2718 );
    nor g2412 ( n9643 , n96 , n10390 );
    or g2413 ( n11020 , n1790 , n11686 );
    xnor g2414 ( n4839 , n5552 , n7367 );
    nor g2415 ( n260 , n11874 , n2716 );
    or g2416 ( n6511 , n12795 , n8490 );
    xnor g2417 ( n8551 , n1940 , n11880 );
    nor g2418 ( n6599 , n1862 , n6180 );
    xnor g2419 ( n11733 , n12833 , n4005 );
    or g2420 ( n11039 , n2254 , n8534 );
    or g2421 ( n7357 , n1587 , n3890 );
    or g2422 ( n7503 , n6724 , n7221 );
    not g2423 ( n5226 , n2498 );
    xnor g2424 ( n2477 , n4572 , n981 );
    or g2425 ( n9588 , n3553 , n4640 );
    not g2426 ( n11738 , n4847 );
    not g2427 ( n12465 , n5189 );
    not g2428 ( n3239 , n11390 );
    and g2429 ( n12013 , n12104 , n12018 );
    or g2430 ( n12191 , n2338 , n13148 );
    not g2431 ( n10195 , n9684 );
    xnor g2432 ( n966 , n11095 , n11243 );
    xnor g2433 ( n11271 , n232 , n1870 );
    xnor g2434 ( n13180 , n9082 , n9687 );
    xnor g2435 ( n4327 , n10672 , n11442 );
    nor g2436 ( n11116 , n6899 , n7214 );
    xnor g2437 ( n3948 , n8361 , n6162 );
    xnor g2438 ( n9768 , n1988 , n6143 );
    nor g2439 ( n4242 , n8981 , n13000 );
    or g2440 ( n4678 , n9195 , n1144 );
    not g2441 ( n202 , n12306 );
    or g2442 ( n8787 , n4727 , n13196 );
    xnor g2443 ( n7028 , n1727 , n4060 );
    or g2444 ( n10878 , n1370 , n4640 );
    or g2445 ( n1616 , n10527 , n12188 );
    xnor g2446 ( n1980 , n7313 , n3500 );
    nor g2447 ( n12157 , n2020 , n5267 );
    xnor g2448 ( n10236 , n10081 , n7282 );
    or g2449 ( n8187 , n8182 , n3716 );
    xnor g2450 ( n11317 , n8770 , n2284 );
    and g2451 ( n12205 , n8938 , n8164 );
    xor g2452 ( n2314 , n7667 , n12961 );
    and g2453 ( n10746 , n4149 , n7147 );
    xnor g2454 ( n3061 , n11530 , n9589 );
    not g2455 ( n4455 , n2771 );
    not g2456 ( n4540 , n7113 );
    nor g2457 ( n1633 , n1826 , n9871 );
    and g2458 ( n7762 , n11780 , n5869 );
    xnor g2459 ( n1859 , n6345 , n8879 );
    and g2460 ( n9499 , n12730 , n6525 );
    nor g2461 ( n7228 , n1540 , n8150 );
    and g2462 ( n1602 , n11800 , n5424 );
    or g2463 ( n7318 , n5865 , n4947 );
    xnor g2464 ( n2770 , n1578 , n8597 );
    nor g2465 ( n4431 , n7480 , n11052 );
    nor g2466 ( n5492 , n4066 , n12622 );
    and g2467 ( n11735 , n10123 , n10822 );
    and g2468 ( n2649 , n13097 , n1577 );
    and g2469 ( n12550 , n3130 , n12284 );
    or g2470 ( n81 , n11581 , n3328 );
    and g2471 ( n541 , n10947 , n2862 );
    or g2472 ( n6556 , n6283 , n11173 );
    not g2473 ( n7683 , n5889 );
    and g2474 ( n282 , n13165 , n8322 );
    xor g2475 ( n4978 , n5845 , n8084 );
    and g2476 ( n3053 , n12051 , n2086 );
    xor g2477 ( n11546 , n11682 , n5355 );
    or g2478 ( n6741 , n8803 , n2903 );
    or g2479 ( n856 , n3646 , n12273 );
    and g2480 ( n8113 , n10973 , n4153 );
    or g2481 ( n1076 , n10447 , n4979 );
    or g2482 ( n2362 , n6024 , n4915 );
    not g2483 ( n9871 , n10627 );
    and g2484 ( n4025 , n2028 , n5468 );
    and g2485 ( n1662 , n693 , n11453 );
    xnor g2486 ( n9890 , n8648 , n8774 );
    and g2487 ( n3114 , n9832 , n3683 );
    xnor g2488 ( n12373 , n7437 , n6762 );
    not g2489 ( n12954 , n5801 );
    nor g2490 ( n6230 , n12698 , n2051 );
    xnor g2491 ( n10976 , n11944 , n4299 );
    xnor g2492 ( n6114 , n10505 , n6161 );
    or g2493 ( n5926 , n8863 , n4640 );
    or g2494 ( n3319 , n11554 , n1156 );
    and g2495 ( n11310 , n5431 , n440 );
    or g2496 ( n4432 , n4464 , n4640 );
    or g2497 ( n1056 , n6914 , n9615 );
    or g2498 ( n3682 , n9017 , n7723 );
    xnor g2499 ( n6013 , n10820 , n10763 );
    nor g2500 ( n12951 , n11327 , n394 );
    xnor g2501 ( n13197 , n1891 , n10084 );
    and g2502 ( n804 , n1644 , n12646 );
    not g2503 ( n97 , n9887 );
    xnor g2504 ( n4439 , n12511 , n2966 );
    xnor g2505 ( n7363 , n4659 , n11507 );
    or g2506 ( n9894 , n7135 , n7075 );
    not g2507 ( n10230 , n10294 );
    xnor g2508 ( n12477 , n4231 , n2073 );
    not g2509 ( n10114 , n39 );
    xnor g2510 ( n1760 , n2426 , n9912 );
    xnor g2511 ( n8333 , n5912 , n1982 );
    or g2512 ( n6870 , n7084 , n2675 );
    xnor g2513 ( n9222 , n9925 , n6361 );
    xnor g2514 ( n1808 , n1394 , n3233 );
    and g2515 ( n8673 , n425 , n6205 );
    xnor g2516 ( n1994 , n1286 , n2617 );
    not g2517 ( n4022 , n12693 );
    and g2518 ( n11154 , n5031 , n1916 );
    not g2519 ( n5157 , n1364 );
    or g2520 ( n8010 , n464 , n1466 );
    xnor g2521 ( n13064 , n4560 , n12923 );
    and g2522 ( n2662 , n3434 , n4021 );
    not g2523 ( n10250 , n9535 );
    xnor g2524 ( n999 , n4857 , n9735 );
    or g2525 ( n9705 , n8225 , n1985 );
    not g2526 ( n2338 , n9906 );
    not g2527 ( n6629 , n3641 );
    nor g2528 ( n3405 , n5151 , n7843 );
    xor g2529 ( n10931 , n9428 , n13173 );
    or g2530 ( n11248 , n5569 , n4373 );
    xnor g2531 ( n404 , n704 , n11516 );
    or g2532 ( n977 , n8174 , n9075 );
    or g2533 ( n6412 , n9581 , n4230 );
    not g2534 ( n8681 , n7374 );
    or g2535 ( n9001 , n115 , n10871 );
    nor g2536 ( n7587 , n2794 , n1467 );
    not g2537 ( n13186 , n12121 );
    xnor g2538 ( n10409 , n11274 , n10559 );
    not g2539 ( n4201 , n3677 );
    xnor g2540 ( n10632 , n4879 , n563 );
    and g2541 ( n6690 , n8492 , n6120 );
    not g2542 ( n7216 , n1724 );
    and g2543 ( n1921 , n8453 , n4825 );
    not g2544 ( n5832 , n6873 );
    or g2545 ( n7493 , n9909 , n7803 );
    nor g2546 ( n11856 , n4211 , n7095 );
    buf g2547 ( n1571 , n438 );
    or g2548 ( n4685 , n8173 , n121 );
    xnor g2549 ( n5475 , n5647 , n1837 );
    nor g2550 ( n12075 , n8080 , n10140 );
    xnor g2551 ( n9004 , n3106 , n7276 );
    and g2552 ( n10885 , n2685 , n7889 );
    and g2553 ( n10581 , n6984 , n1297 );
    not g2554 ( n808 , n5320 );
    not g2555 ( n8472 , n4862 );
    nor g2556 ( n12983 , n9082 , n13074 );
    xnor g2557 ( n3604 , n8949 , n6637 );
    and g2558 ( n8375 , n8401 , n337 );
    nor g2559 ( n8062 , n10416 , n11030 );
    xnor g2560 ( n2593 , n5833 , n10370 );
    xor g2561 ( n12661 , n1938 , n12932 );
    or g2562 ( n5227 , n3563 , n11870 );
    or g2563 ( n1978 , n2449 , n8702 );
    xnor g2564 ( n12616 , n3372 , n7577 );
    and g2565 ( n10389 , n2493 , n4203 );
    not g2566 ( n5479 , n3894 );
    not g2567 ( n12798 , n10019 );
    xnor g2568 ( n3475 , n10247 , n2756 );
    not g2569 ( n11643 , n7516 );
    xnor g2570 ( n10945 , n2389 , n2051 );
    or g2571 ( n2842 , n12224 , n1144 );
    not g2572 ( n10103 , n61 );
    not g2573 ( n3454 , n8230 );
    and g2574 ( n5073 , n8978 , n9733 );
    not g2575 ( n9070 , n3192 );
    xor g2576 ( n9399 , n5871 , n8974 );
    and g2577 ( n492 , n2015 , n1701 );
    or g2578 ( n9054 , n13073 , n3426 );
    xnor g2579 ( n1031 , n529 , n8705 );
    xnor g2580 ( n10251 , n9375 , n10204 );
    xor g2581 ( n12966 , n10512 , n5827 );
    and g2582 ( n4562 , n1998 , n5357 );
    and g2583 ( n4773 , n5214 , n4330 );
    nor g2584 ( n1317 , n6418 , n1738 );
    and g2585 ( n295 , n7219 , n7222 );
    or g2586 ( n2608 , n172 , n4973 );
    and g2587 ( n4003 , n11227 , n2676 );
    and g2588 ( n5354 , n3078 , n6952 );
    not g2589 ( n12395 , n8183 );
    or g2590 ( n484 , n9810 , n542 );
    nor g2591 ( n3089 , n605 , n11395 );
    xnor g2592 ( n4769 , n710 , n3376 );
    xnor g2593 ( n9758 , n3117 , n7457 );
    nor g2594 ( n304 , n6144 , n11621 );
    xnor g2595 ( n4368 , n6643 , n2845 );
    xnor g2596 ( n2084 , n6465 , n9647 );
    or g2597 ( n3363 , n8621 , n9935 );
    nor g2598 ( n6824 , n11824 , n10658 );
    or g2599 ( n2401 , n8173 , n12395 );
    nor g2600 ( n326 , n1988 , n10035 );
    xnor g2601 ( n2128 , n4937 , n6192 );
    and g2602 ( n3960 , n5231 , n7227 );
    xnor g2603 ( n3002 , n10456 , n7664 );
    or g2604 ( n7117 , n3293 , n947 );
    or g2605 ( n470 , n7354 , n5743 );
    or g2606 ( n7459 , n1718 , n7567 );
    or g2607 ( n6316 , n3407 , n1026 );
    not g2608 ( n7888 , n11123 );
    buf g2609 ( n7221 , n11940 );
    xor g2610 ( n7313 , n9729 , n6758 );
    or g2611 ( n7918 , n10005 , n10117 );
    or g2612 ( n9234 , n10465 , n1463 );
    and g2613 ( n6284 , n723 , n10506 );
    or g2614 ( n8390 , n5683 , n12721 );
    or g2615 ( n7906 , n121 , n1869 );
    nor g2616 ( n3635 , n7328 , n6025 );
    or g2617 ( n7469 , n11420 , n2363 );
    and g2618 ( n1404 , n9760 , n11392 );
    xnor g2619 ( n780 , n4742 , n3837 );
    xnor g2620 ( n12696 , n10344 , n70 );
    or g2621 ( n233 , n621 , n3246 );
    and g2622 ( n2481 , n4400 , n12285 );
    not g2623 ( n545 , n5594 );
    xnor g2624 ( n3291 , n1901 , n11874 );
    and g2625 ( n1953 , n8466 , n8233 );
    buf g2626 ( n6899 , n7906 );
    xnor g2627 ( n4801 , n7131 , n11136 );
    and g2628 ( n8524 , n5748 , n11221 );
    or g2629 ( n200 , n8361 , n6162 );
    and g2630 ( n2871 , n9949 , n11889 );
    xnor g2631 ( n12547 , n386 , n3369 );
    or g2632 ( n2570 , n12836 , n1819 );
    nor g2633 ( n409 , n10613 , n10711 );
    or g2634 ( n511 , n2872 , n9159 );
    and g2635 ( n4682 , n10981 , n5187 );
    not g2636 ( n3724 , n11953 );
    xnor g2637 ( n10850 , n6717 , n291 );
    or g2638 ( n5826 , n12490 , n2059 );
    and g2639 ( n1237 , n2018 , n854 );
    or g2640 ( n5828 , n2329 , n1026 );
    xnor g2641 ( n5100 , n3914 , n8503 );
    and g2642 ( n5424 , n5905 , n6727 );
    and g2643 ( n8271 , n11537 , n9915 );
    xnor g2644 ( n6895 , n7774 , n11355 );
    nor g2645 ( n3929 , n12270 , n12076 );
    or g2646 ( n10077 , n8306 , n11982 );
    and g2647 ( n10354 , n5913 , n6412 );
    and g2648 ( n7006 , n10908 , n8468 );
    or g2649 ( n2282 , n845 , n8563 );
    xnor g2650 ( n11568 , n10850 , n1486 );
    xnor g2651 ( n5293 , n8674 , n1403 );
    or g2652 ( n3467 , n12357 , n13133 );
    or g2653 ( n11599 , n3281 , n3981 );
    and g2654 ( n7572 , n4267 , n6152 );
    not g2655 ( n9018 , n11906 );
    not g2656 ( n6355 , n817 );
    or g2657 ( n2643 , n11871 , n3225 );
    or g2658 ( n8193 , n6481 , n3651 );
    not g2659 ( n8777 , n5962 );
    and g2660 ( n3229 , n5004 , n4314 );
    or g2661 ( n6016 , n11542 , n12695 );
    or g2662 ( n940 , n712 , n9136 );
    and g2663 ( n10385 , n8210 , n10310 );
    not g2664 ( n13108 , n761 );
    not g2665 ( n196 , n8134 );
    or g2666 ( n3936 , n5086 , n1741 );
    not g2667 ( n6906 , n4687 );
    or g2668 ( n879 , n1823 , n7704 );
    xnor g2669 ( n758 , n3715 , n8831 );
    xnor g2670 ( n2650 , n2196 , n1295 );
    not g2671 ( n4910 , n6244 );
    not g2672 ( n4272 , n11350 );
    or g2673 ( n11620 , n10317 , n12361 );
    and g2674 ( n12138 , n10752 , n10666 );
    nor g2675 ( n10540 , n1219 , n4567 );
    or g2676 ( n8890 , n5694 , n5242 );
    or g2677 ( n752 , n3428 , n12695 );
    xnor g2678 ( n3625 , n40 , n7873 );
    and g2679 ( n350 , n1588 , n12536 );
    xnor g2680 ( n2664 , n8328 , n10434 );
    or g2681 ( n4602 , n1335 , n1089 );
    xnor g2682 ( n8100 , n2911 , n11506 );
    or g2683 ( n8440 , n12294 , n7435 );
    and g2684 ( n7611 , n2443 , n11641 );
    xnor g2685 ( n403 , n6892 , n9952 );
    or g2686 ( n10981 , n8495 , n8929 );
    and g2687 ( n4064 , n9104 , n4852 );
    xnor g2688 ( n2244 , n862 , n7895 );
    not g2689 ( n2232 , n4862 );
    xnor g2690 ( n10456 , n8080 , n1576 );
    and g2691 ( n909 , n1757 , n3409 );
    nor g2692 ( n3917 , n10242 , n10050 );
    xnor g2693 ( n11309 , n8683 , n10208 );
    nor g2694 ( n10915 , n5690 , n4032 );
    or g2695 ( n10171 , n6412 , n5913 );
    or g2696 ( n5070 , n379 , n12273 );
    xnor g2697 ( n6542 , n11063 , n8862 );
    not g2698 ( n9931 , n12482 );
    xnor g2699 ( n6705 , n13054 , n12084 );
    not g2700 ( n12604 , n9620 );
    and g2701 ( n11381 , n7160 , n4374 );
    or g2702 ( n10099 , n7688 , n12524 );
    or g2703 ( n6776 , n3115 , n597 );
    or g2704 ( n5290 , n10032 , n8030 );
    not g2705 ( n7864 , n2072 );
    xnor g2706 ( n10833 , n3001 , n12179 );
    or g2707 ( n5115 , n5146 , n3981 );
    and g2708 ( n4460 , n12274 , n5111 );
    xnor g2709 ( n918 , n2900 , n6793 );
    nor g2710 ( n10309 , n1655 , n1482 );
    or g2711 ( n7438 , n44 , n3981 );
    xnor g2712 ( n5937 , n3730 , n9932 );
    and g2713 ( n2030 , n4943 , n2124 );
    not g2714 ( n1744 , n8203 );
    and g2715 ( n5027 , n89 , n1813 );
    nor g2716 ( n1822 , n1481 , n7848 );
    xnor g2717 ( n4667 , n11490 , n6282 );
    and g2718 ( n11748 , n7658 , n8512 );
    xor g2719 ( n4539 , n12560 , n7854 );
    xnor g2720 ( n11071 , n472 , n5260 );
    and g2721 ( n7691 , n13024 , n6887 );
    xnor g2722 ( n2734 , n11663 , n8269 );
    not g2723 ( n2556 , n8506 );
    xnor g2724 ( n23 , n4629 , n2643 );
    xnor g2725 ( n5824 , n2874 , n8635 );
    not g2726 ( n8391 , n2501 );
    not g2727 ( n12734 , n5371 );
    not g2728 ( n6760 , n13076 );
    xnor g2729 ( n9226 , n6822 , n10776 );
    nor g2730 ( n1580 , n12130 , n12181 );
    and g2731 ( n9609 , n19 , n3549 );
    xnor g2732 ( n9687 , n4074 , n6232 );
    or g2733 ( n9691 , n2165 , n5409 );
    or g2734 ( n12972 , n1943 , n12519 );
    or g2735 ( n6123 , n1052 , n8563 );
    not g2736 ( n8040 , n4933 );
    and g2737 ( n12759 , n6454 , n1975 );
    not g2738 ( n1901 , n10459 );
    nor g2739 ( n9799 , n4934 , n5084 );
    or g2740 ( n7684 , n5163 , n5242 );
    xnor g2741 ( n1049 , n2260 , n4446 );
    and g2742 ( n447 , n6671 , n6441 );
    nor g2743 ( n5269 , n5213 , n12687 );
    and g2744 ( n8586 , n3687 , n1800 );
    or g2745 ( n9204 , n3157 , n8206 );
    xor g2746 ( n2844 , n3705 , n5938 );
    or g2747 ( n7366 , n6629 , n1985 );
    and g2748 ( n8128 , n7649 , n7031 );
    and g2749 ( n3264 , n4114 , n11222 );
    nor g2750 ( n10323 , n2187 , n2612 );
    or g2751 ( n2948 , n5562 , n3981 );
    or g2752 ( n11153 , n10018 , n121 );
    not g2753 ( n588 , n1393 );
    nor g2754 ( n10487 , n5020 , n1512 );
    not g2755 ( n11772 , n8230 );
    not g2756 ( n1733 , n12627 );
    xnor g2757 ( n522 , n2193 , n4167 );
    not g2758 ( n5268 , n1160 );
    or g2759 ( n1006 , n235 , n4285 );
    not g2760 ( n13229 , n5543 );
    not g2761 ( n12234 , n7336 );
    xnor g2762 ( n13227 , n9161 , n1726 );
    or g2763 ( n4638 , n1361 , n6910 );
    or g2764 ( n9695 , n5890 , n4373 );
    xnor g2765 ( n7552 , n10731 , n7540 );
    or g2766 ( n2728 , n11722 , n7502 );
    or g2767 ( n4054 , n6526 , n1951 );
    xnor g2768 ( n55 , n1223 , n8189 );
    xnor g2769 ( n6529 , n10479 , n4522 );
    not g2770 ( n10597 , n6654 );
    or g2771 ( n5840 , n2834 , n5298 );
    or g2772 ( n1867 , n11303 , n4990 );
    xnor g2773 ( n9802 , n4542 , n12259 );
    xnor g2774 ( n646 , n7696 , n13230 );
    and g2775 ( n4825 , n9889 , n4841 );
    not g2776 ( n6193 , n8716 );
    and g2777 ( n9895 , n5974 , n3655 );
    nor g2778 ( n8595 , n1306 , n1682 );
    not g2779 ( n2041 , n5729 );
    nor g2780 ( n4990 , n4789 , n8467 );
    xnor g2781 ( n13034 , n9158 , n2288 );
    and g2782 ( n7304 , n4338 , n13093 );
    or g2783 ( n7484 , n11542 , n4373 );
    xnor g2784 ( n5777 , n1489 , n5281 );
    and g2785 ( n8819 , n9284 , n11660 );
    or g2786 ( n1178 , n9702 , n3225 );
    or g2787 ( n11124 , n12473 , n2530 );
    or g2788 ( n9109 , n8758 , n10285 );
    xnor g2789 ( n1475 , n8590 , n3035 );
    or g2790 ( n2624 , n2111 , n3162 );
    nor g2791 ( n8343 , n6042 , n6829 );
    xnor g2792 ( n6322 , n1074 , n4893 );
    or g2793 ( n6979 , n1268 , n6885 );
    and g2794 ( n9965 , n3514 , n8191 );
    not g2795 ( n12673 , n3040 );
    and g2796 ( n10961 , n6979 , n57 );
    or g2797 ( n11703 , n9389 , n5061 );
    xnor g2798 ( n8962 , n5385 , n8636 );
    or g2799 ( n2227 , n2542 , n2287 );
    xnor g2800 ( n7512 , n6947 , n4511 );
    not g2801 ( n1360 , n4998 );
    and g2802 ( n9615 , n534 , n5416 );
    xnor g2803 ( n11051 , n7782 , n13038 );
    xnor g2804 ( n11845 , n12861 , n6440 );
    xnor g2805 ( n12678 , n10296 , n5145 );
    xor g2806 ( n4709 , n1252 , n13165 );
    not g2807 ( n7661 , n2882 );
    or g2808 ( n5247 , n7856 , n9873 );
    or g2809 ( n5172 , n12772 , n4991 );
    xnor g2810 ( n6431 , n61 , n9896 );
    xnor g2811 ( n7326 , n4392 , n12893 );
    not g2812 ( n2915 , n7515 );
    nor g2813 ( n9696 , n591 , n7554 );
    xnor g2814 ( n10984 , n11862 , n4129 );
    xnor g2815 ( n10562 , n6235 , n8802 );
    xnor g2816 ( n5873 , n7162 , n3672 );
    xnor g2817 ( n10628 , n8071 , n7799 );
    not g2818 ( n6142 , n10799 );
    xnor g2819 ( n3659 , n6530 , n9758 );
    not g2820 ( n7963 , n1497 );
    or g2821 ( n1440 , n8724 , n12064 );
    xnor g2822 ( n2894 , n6855 , n8832 );
    xnor g2823 ( n11394 , n3175 , n10769 );
    not g2824 ( n5079 , n9187 );
    and g2825 ( n878 , n26 , n1239 );
    xnor g2826 ( n3738 , n10220 , n5387 );
    xnor g2827 ( n11897 , n6349 , n11309 );
    nor g2828 ( n802 , n12457 , n2810 );
    xnor g2829 ( n7677 , n7573 , n9219 );
    or g2830 ( n11595 , n4986 , n4694 );
    xnor g2831 ( n6709 , n3657 , n7650 );
    xor g2832 ( n8330 , n11049 , n4320 );
    or g2833 ( n12190 , n1286 , n12736 );
    not g2834 ( n11040 , n5705 );
    xnor g2835 ( n12485 , n9969 , n6249 );
    not g2836 ( n7907 , n4909 );
    and g2837 ( n939 , n8230 , n9531 );
    nor g2838 ( n10996 , n8396 , n11383 );
    and g2839 ( n6978 , n8871 , n7139 );
    not g2840 ( n5490 , n11190 );
    xnor g2841 ( n12364 , n524 , n5617 );
    and g2842 ( n12785 , n1285 , n12055 );
    or g2843 ( n11550 , n2678 , n5076 );
    xnor g2844 ( n12769 , n13107 , n5619 );
    xor g2845 ( n7970 , n7501 , n9063 );
    xnor g2846 ( n4282 , n509 , n4882 );
    xnor g2847 ( n11977 , n8099 , n12766 );
    xnor g2848 ( n25 , n4879 , n8760 );
    not g2849 ( n4891 , n9738 );
    not g2850 ( n11364 , n726 );
    not g2851 ( n12886 , n1900 );
    xnor g2852 ( n7651 , n11118 , n6214 );
    not g2853 ( n60 , n9636 );
    nor g2854 ( n8747 , n2835 , n6833 );
    not g2855 ( n11621 , n362 );
    xnor g2856 ( n3379 , n12574 , n5951 );
    not g2857 ( n3965 , n12605 );
    and g2858 ( n8579 , n1908 , n11279 );
    or g2859 ( n6767 , n9144 , n6870 );
    xnor g2860 ( n4764 , n8772 , n506 );
    and g2861 ( n814 , n9140 , n174 );
    xnor g2862 ( n387 , n1060 , n10159 );
    xnor g2863 ( n704 , n463 , n9961 );
    not g2864 ( n10245 , n4828 );
    not g2865 ( n5461 , n11537 );
    nor g2866 ( n9703 , n10051 , n1140 );
    xnor g2867 ( n13164 , n1903 , n8375 );
    xnor g2868 ( n7334 , n5892 , n2030 );
    not g2869 ( n3017 , n8715 );
    or g2870 ( n10020 , n8510 , n12718 );
    or g2871 ( n8915 , n11472 , n6882 );
    xor g2872 ( n11503 , n5360 , n7970 );
    and g2873 ( n1433 , n9482 , n12323 );
    or g2874 ( n9978 , n4109 , n964 );
    xnor g2875 ( n11839 , n2034 , n11150 );
    not g2876 ( n9125 , n11673 );
    xnor g2877 ( n12577 , n7688 , n12524 );
    not g2878 ( n8108 , n1165 );
    and g2879 ( n12943 , n12595 , n1881 );
    xnor g2880 ( n5395 , n8846 , n4440 );
    or g2881 ( n10918 , n3126 , n2958 );
    not g2882 ( n783 , n8841 );
    xnor g2883 ( n11921 , n2432 , n3521 );
    xnor g2884 ( n2587 , n3964 , n6879 );
    xnor g2885 ( n5128 , n3568 , n5641 );
    xnor g2886 ( n220 , n3679 , n7600 );
    xnor g2887 ( n11189 , n8157 , n9576 );
    nor g2888 ( n742 , n11012 , n3674 );
    and g2889 ( n12700 , n4397 , n8165 );
    not g2890 ( n12814 , n4862 );
    nor g2891 ( n11098 , n7795 , n3803 );
    nor g2892 ( n12924 , n10114 , n11332 );
    or g2893 ( n11360 , n9316 , n10072 );
    not g2894 ( n7291 , n5729 );
    not g2895 ( n6913 , n5185 );
    nor g2896 ( n11554 , n12661 , n10321 );
    or g2897 ( n6229 , n6407 , n6404 );
    not g2898 ( n11759 , n5389 );
    or g2899 ( n5613 , n9289 , n7831 );
    not g2900 ( n11542 , n9846 );
    or g2901 ( n7170 , n321 , n10319 );
    nor g2902 ( n1863 , n10183 , n1949 );
    xnor g2903 ( n8516 , n7959 , n2529 );
    not g2904 ( n10314 , n2737 );
    nor g2905 ( n10302 , n11645 , n2 );
    not g2906 ( n8351 , n1764 );
    or g2907 ( n8449 , n10914 , n7185 );
    xnor g2908 ( n2940 , n7862 , n7166 );
    xnor g2909 ( n13224 , n678 , n166 );
    nor g2910 ( n7150 , n612 , n9986 );
    not g2911 ( n7890 , n5470 );
    xnor g2912 ( n6780 , n2962 , n1415 );
    not g2913 ( n89 , n6675 );
    or g2914 ( n8381 , n5445 , n5681 );
    xnor g2915 ( n6628 , n12843 , n8988 );
    not g2916 ( n6138 , n7539 );
    nor g2917 ( n5619 , n5280 , n8439 );
    xnor g2918 ( n8976 , n1418 , n10875 );
    not g2919 ( n5383 , n8887 );
    not g2920 ( n7741 , n12853 );
    xnor g2921 ( n5880 , n11715 , n2968 );
    nor g2922 ( n7047 , n10120 , n346 );
    nor g2923 ( n8828 , n2550 , n9472 );
    nor g2924 ( n10267 , n6754 , n8094 );
    or g2925 ( n6024 , n2449 , n6404 );
    or g2926 ( n2383 , n3532 , n9190 );
    and g2927 ( n8376 , n11957 , n4958 );
    xnor g2928 ( n10347 , n10817 , n8067 );
    or g2929 ( n2433 , n11851 , n157 );
    xnor g2930 ( n2851 , n12545 , n6631 );
    nor g2931 ( n2568 , n8124 , n4262 );
    and g2932 ( n11068 , n8987 , n3508 );
    not g2933 ( n3552 , n1503 );
    or g2934 ( n11382 , n1688 , n1463 );
    xnor g2935 ( n1225 , n7611 , n6570 );
    nor g2936 ( n12048 , n8714 , n11853 );
    xnor g2937 ( n8465 , n6336 , n8752 );
    nor g2938 ( n4609 , n695 , n7483 );
    or g2939 ( n8619 , n8599 , n6468 );
    or g2940 ( n12332 , n6875 , n4373 );
    or g2941 ( n10593 , n12914 , n5917 );
    not g2942 ( n7939 , n9138 );
    not g2943 ( n7249 , n6385 );
    or g2944 ( n5194 , n7135 , n9195 );
    nor g2945 ( n3979 , n7064 , n4250 );
    xnor g2946 ( n6454 , n1598 , n2273 );
    not g2947 ( n8363 , n3321 );
    xnor g2948 ( n273 , n11674 , n7092 );
    and g2949 ( n8052 , n12412 , n4174 );
    nor g2950 ( n5495 , n1764 , n2213 );
    and g2951 ( n8469 , n1594 , n7337 );
    or g2952 ( n2236 , n7880 , n4230 );
    or g2953 ( n11027 , n12225 , n9012 );
    xnor g2954 ( n6301 , n11452 , n6815 );
    and g2955 ( n3722 , n2057 , n2882 );
    not g2956 ( n1941 , n6149 );
    or g2957 ( n11307 , n10499 , n6893 );
    not g2958 ( n1649 , n11816 );
    xnor g2959 ( n12779 , n8882 , n1850 );
    xnor g2960 ( n1670 , n1240 , n12630 );
    or g2961 ( n3935 , n2581 , n13108 );
    not g2962 ( n1605 , n951 );
    nor g2963 ( n3886 , n8229 , n4633 );
    not g2964 ( n1807 , n10548 );
    or g2965 ( n3490 , n6488 , n12388 );
    or g2966 ( n11251 , n8179 , n7140 );
    or g2967 ( n7856 , n8400 , n5242 );
    or g2968 ( n3029 , n1325 , n5423 );
    and g2969 ( n2 , n4365 , n2507 );
    and g2970 ( n3271 , n3932 , n7015 );
    or g2971 ( n13075 , n6132 , n8783 );
    and g2972 ( n3558 , n6378 , n9325 );
    and g2973 ( n11131 , n2386 , n6899 );
    and g2974 ( n5767 , n11274 , n12993 );
    and g2975 ( n2853 , n6928 , n1711 );
    xnor g2976 ( n5012 , n12976 , n4341 );
    not g2977 ( n7243 , n8288 );
    not g2978 ( n8626 , n12916 );
    or g2979 ( n8186 , n7376 , n2455 );
    xnor g2980 ( n1880 , n8565 , n4938 );
    xnor g2981 ( n5618 , n13093 , n2436 );
    or g2982 ( n12496 , n5611 , n2544 );
    and g2983 ( n7957 , n2963 , n8010 );
    xnor g2984 ( n4234 , n3496 , n12862 );
    and g2985 ( n157 , n9854 , n11193 );
    xnor g2986 ( n3349 , n3594 , n4632 );
    not g2987 ( n5746 , n6904 );
    or g2988 ( n7902 , n10045 , n7935 );
    and g2989 ( n12704 , n9905 , n173 );
    not g2990 ( n871 , n12085 );
    not g2991 ( n2136 , n1130 );
    or g2992 ( n6337 , n9730 , n11479 );
    not g2993 ( n5066 , n7710 );
    xnor g2994 ( n12239 , n12162 , n511 );
    not g2995 ( n12484 , n5408 );
    xor g2996 ( n836 , n10279 , n9447 );
    not g2997 ( n3819 , n10563 );
    xnor g2998 ( n9587 , n1284 , n12369 );
    xnor g2999 ( n5698 , n10073 , n731 );
    xnor g3000 ( n12892 , n2913 , n10747 );
    xnor g3001 ( n9676 , n3307 , n11326 );
    not g3002 ( n6364 , n11488 );
    xnor g3003 ( n1951 , n2937 , n7764 );
    or g3004 ( n8599 , n5949 , n4230 );
    or g3005 ( n5351 , n6883 , n4947 );
    not g3006 ( n11003 , n3264 );
    not g3007 ( n193 , n2220 );
    and g3008 ( n6604 , n81 , n9884 );
    not g3009 ( n3764 , n9898 );
    and g3010 ( n5234 , n9430 , n2579 );
    xnor g3011 ( n9824 , n1866 , n2075 );
    or g3012 ( n5179 , n10780 , n8348 );
    and g3013 ( n7008 , n7862 , n9861 );
    and g3014 ( n4248 , n2418 , n9945 );
    nor g3015 ( n12385 , n729 , n4700 );
    xnor g3016 ( n1423 , n6280 , n8121 );
    or g3017 ( n11617 , n10901 , n10687 );
    xnor g3018 ( n2303 , n8489 , n7853 );
    or g3019 ( n6068 , n10587 , n10871 );
    xnor g3020 ( n3663 , n11997 , n10062 );
    or g3021 ( n12285 , n6129 , n9075 );
    not g3022 ( n8948 , n7895 );
    xnor g3023 ( n8798 , n2433 , n5064 );
    not g3024 ( n6922 , n11350 );
    not g3025 ( n2145 , n938 );
    xnor g3026 ( n10695 , n5131 , n10397 );
    or g3027 ( n8358 , n7950 , n4936 );
    xnor g3028 ( n7835 , n8957 , n581 );
    or g3029 ( n7951 , n1207 , n7008 );
    and g3030 ( n11708 , n9161 , n6372 );
    or g3031 ( n4397 , n7372 , n4107 );
    xnor g3032 ( n284 , n11283 , n349 );
    or g3033 ( n8770 , n12249 , n5242 );
    nor g3034 ( n2936 , n3027 , n3717 );
    xnor g3035 ( n4210 , n484 , n960 );
    xnor g3036 ( n1129 , n2776 , n6201 );
    xnor g3037 ( n3751 , n1682 , n4347 );
    or g3038 ( n7776 , n12434 , n479 );
    not g3039 ( n5099 , n3354 );
    and g3040 ( n11754 , n895 , n1639 );
    or g3041 ( n1312 , n1296 , n4936 );
    or g3042 ( n4021 , n4540 , n1463 );
    or g3043 ( n992 , n10230 , n8283 );
    or g3044 ( n8576 , n2264 , n11144 );
    and g3045 ( n1771 , n8139 , n6826 );
    and g3046 ( n5864 , n8693 , n709 );
    or g3047 ( n11357 , n12528 , n2694 );
    xnor g3048 ( n13038 , n11915 , n4133 );
    or g3049 ( n8539 , n1416 , n8868 );
    xnor g3050 ( n2837 , n5503 , n1452 );
    xnor g3051 ( n2855 , n2842 , n9484 );
    nor g3052 ( n681 , n1173 , n3628 );
    xnor g3053 ( n6252 , n2016 , n9685 );
    xnor g3054 ( n9473 , n10811 , n10008 );
    nor g3055 ( n10557 , n3045 , n8577 );
    and g3056 ( n6840 , n1729 , n6745 );
    xnor g3057 ( n7447 , n8671 , n1624 );
    xnor g3058 ( n3667 , n4681 , n11979 );
    or g3059 ( n797 , n10527 , n1463 );
    not g3060 ( n8231 , n346 );
    and g3061 ( n7093 , n9967 , n1442 );
    and g3062 ( n815 , n313 , n4212 );
    or g3063 ( n11994 , n569 , n2544 );
    not g3064 ( n3293 , n9475 );
    xnor g3065 ( n9742 , n2585 , n11238 );
    or g3066 ( n7287 , n971 , n5242 );
    xnor g3067 ( n2682 , n5307 , n709 );
    buf g3068 ( n8490 , n2557 );
    or g3069 ( n5597 , n9069 , n8534 );
    nor g3070 ( n5482 , n6165 , n2448 );
    not g3071 ( n9810 , n401 );
    xnor g3072 ( n3274 , n8223 , n6520 );
    xnor g3073 ( n5718 , n7953 , n2871 );
    not g3074 ( n6144 , n6603 );
    not g3075 ( n12045 , n1771 );
    not g3076 ( n3338 , n4043 );
    xnor g3077 ( n12618 , n11924 , n7609 );
    or g3078 ( n5874 , n4209 , n7846 );
    xor g3079 ( n3448 , n4043 , n1171 );
    xnor g3080 ( n9694 , n1620 , n2743 );
    or g3081 ( n11570 , n4722 , n8563 );
    xnor g3082 ( n7816 , n9731 , n674 );
    xnor g3083 ( n4151 , n8675 , n6429 );
    and g3084 ( n9141 , n12674 , n1001 );
    nor g3085 ( n12202 , n11084 , n4931 );
    not g3086 ( n10886 , n11324 );
    xnor g3087 ( n2349 , n12218 , n10283 );
    and g3088 ( n4133 , n9266 , n5822 );
    or g3089 ( n4659 , n9808 , n542 );
    xnor g3090 ( n12228 , n7982 , n3426 );
    or g3091 ( n7 , n6033 , n13242 );
    xnor g3092 ( n1866 , n2496 , n6696 );
    xnor g3093 ( n6593 , n12662 , n6691 );
    not g3094 ( n436 , n10048 );
    or g3095 ( n8134 , n10958 , n792 );
    not g3096 ( n2625 , n13014 );
    xnor g3097 ( n7482 , n5700 , n8278 );
    nor g3098 ( n4147 , n11281 , n4702 );
    or g3099 ( n9083 , n2129 , n12062 );
    xnor g3100 ( n11184 , n10001 , n6673 );
    not g3101 ( n5707 , n4885 );
    xor g3102 ( n7575 , n9924 , n5668 );
    xnor g3103 ( n4572 , n3797 , n4705 );
    not g3104 ( n7082 , n4249 );
    xnor g3105 ( n1393 , n8924 , n3439 );
    or g3106 ( n1250 , n9767 , n9195 );
    xnor g3107 ( n1195 , n11717 , n8608 );
    or g3108 ( n11193 , n7422 , n9178 );
    xnor g3109 ( n10524 , n5253 , n4860 );
    or g3110 ( n4081 , n6638 , n6635 );
    or g3111 ( n10412 , n9511 , n8348 );
    xnor g3112 ( n4202 , n170 , n12547 );
    nor g3113 ( n7380 , n5354 , n1831 );
    xnor g3114 ( n1567 , n1683 , n12557 );
    nor g3115 ( n11978 , n299 , n967 );
    or g3116 ( n13128 , n11284 , n1043 );
    xnor g3117 ( n5816 , n7747 , n1183 );
    nor g3118 ( n12351 , n2568 , n1608 );
    or g3119 ( n9806 , n11114 , n12188 );
    not g3120 ( n5595 , n8332 );
    xnor g3121 ( n4083 , n10847 , n10061 );
    nor g3122 ( n7693 , n10806 , n1489 );
    or g3123 ( n11878 , n11861 , n8016 );
    or g3124 ( n5425 , n5146 , n5242 );
    or g3125 ( n11419 , n10859 , n8209 );
    or g3126 ( n5314 , n5935 , n4854 );
    xnor g3127 ( n12334 , n6248 , n1016 );
    not g3128 ( n12093 , n9887 );
    not g3129 ( n9650 , n1734 );
    or g3130 ( n5108 , n2971 , n6684 );
    nor g3131 ( n10050 , n7850 , n3329 );
    or g3132 ( n11380 , n5163 , n9223 );
    xnor g3133 ( n6583 , n7028 , n10542 );
    not g3134 ( n10332 , n4439 );
    nor g3135 ( n11791 , n7497 , n3386 );
    or g3136 ( n8355 , n8629 , n1161 );
    xnor g3137 ( n6450 , n6750 , n7653 );
    not g3138 ( n10361 , n1758 );
    xnor g3139 ( n12960 , n12703 , n13046 );
    xnor g3140 ( n7451 , n11714 , n1772 );
    or g3141 ( n8659 , n12155 , n10362 );
    and g3142 ( n3337 , n3382 , n10640 );
    or g3143 ( n5545 , n7401 , n7855 );
    not g3144 ( n2321 , n3311 );
    not g3145 ( n11094 , n12372 );
    and g3146 ( n266 , n5787 , n735 );
    xnor g3147 ( n7476 , n12619 , n6115 );
    or g3148 ( n6217 , n533 , n1287 );
    xnor g3149 ( n9163 , n10153 , n9183 );
    nor g3150 ( n163 , n7463 , n11884 );
    or g3151 ( n8397 , n790 , n12419 );
    xnor g3152 ( n1066 , n2227 , n7126 );
    xnor g3153 ( n5405 , n4757 , n11450 );
    not g3154 ( n26 , n4747 );
    xnor g3155 ( n3512 , n6299 , n1882 );
    not g3156 ( n5158 , n2343 );
    nor g3157 ( n5297 , n5380 , n6524 );
    and g3158 ( n6091 , n12656 , n10807 );
    xnor g3159 ( n10801 , n11698 , n7492 );
    and g3160 ( n9426 , n12495 , n4772 );
    not g3161 ( n3078 , n8149 );
    xnor g3162 ( n62 , n9334 , n8456 );
    xnor g3163 ( n11675 , n4614 , n8014 );
    or g3164 ( n5015 , n1989 , n7377 );
    not g3165 ( n9693 , n8689 );
    xnor g3166 ( n1641 , n1939 , n381 );
    and g3167 ( n9822 , n12665 , n11091 );
    not g3168 ( n5289 , n2731 );
    not g3169 ( n4612 , n12065 );
    xnor g3170 ( n922 , n7957 , n9566 );
    and g3171 ( n6005 , n6858 , n3665 );
    xnor g3172 ( n4254 , n5998 , n724 );
    nor g3173 ( n12723 , n8328 , n12508 );
    nor g3174 ( n11368 , n4651 , n10210 );
    and g3175 ( n4377 , n8661 , n7529 );
    or g3176 ( n11385 , n12462 , n5092 );
    xnor g3177 ( n131 , n12237 , n9506 );
    xnor g3178 ( n4914 , n10348 , n7590 );
    or g3179 ( n1375 , n13036 , n10871 );
    xnor g3180 ( n1016 , n120 , n12028 );
    or g3181 ( n6029 , n8412 , n273 );
    or g3182 ( n6830 , n2002 , n2308 );
    xnor g3183 ( n3976 , n1984 , n4483 );
    and g3184 ( n4457 , n9706 , n412 );
    or g3185 ( n685 , n5038 , n11368 );
    xnor g3186 ( n9935 , n4128 , n9982 );
    and g3187 ( n10078 , n7715 , n3409 );
    nor g3188 ( n3585 , n10774 , n11777 );
    xnor g3189 ( n2983 , n10238 , n6286 );
    and g3190 ( n7848 , n343 , n9750 );
    xnor g3191 ( n4997 , n6835 , n3476 );
    not g3192 ( n2641 , n10805 );
    not g3193 ( n3068 , n2341 );
    nor g3194 ( n285 , n12632 , n3990 );
    xnor g3195 ( n7478 , n9970 , n8625 );
    xor g3196 ( n9654 , n7087 , n3008 );
    or g3197 ( n5138 , n13231 , n6128 );
    or g3198 ( n11450 , n1695 , n6635 );
    and g3199 ( n6987 , n11213 , n11241 );
    or g3200 ( n5018 , n7925 , n5242 );
    xnor g3201 ( n5879 , n6455 , n2724 );
    xnor g3202 ( n1299 , n10799 , n4097 );
    not g3203 ( n13077 , n9093 );
    and g3204 ( n9035 , n11184 , n7503 );
    not g3205 ( n12126 , n9531 );
    or g3206 ( n9356 , n11933 , n8702 );
    buf g3207 ( n121 , n12335 );
    or g3208 ( n8891 , n3498 , n905 );
    and g3209 ( n8041 , n2961 , n9142 );
    or g3210 ( n3714 , n12732 , n9075 );
    not g3211 ( n4465 , n287 );
    and g3212 ( n10701 , n11065 , n8708 );
    nor g3213 ( n269 , n12505 , n9787 );
    xnor g3214 ( n9193 , n1265 , n8804 );
    nor g3215 ( n7535 , n1628 , n3202 );
    and g3216 ( n2445 , n2469 , n2383 );
    and g3217 ( n6982 , n6850 , n4229 );
    xnor g3218 ( n4775 , n7235 , n7703 );
    or g3219 ( n1428 , n2670 , n546 );
    xnor g3220 ( n2395 , n3942 , n3089 );
    and g3221 ( n621 , n1040 , n5564 );
    and g3222 ( n8078 , n609 , n4677 );
    and g3223 ( n6140 , n10168 , n12263 );
    nor g3224 ( n7714 , n636 , n9365 );
    not g3225 ( n6559 , n11134 );
    or g3226 ( n11562 , n493 , n1144 );
    not g3227 ( n5341 , n7036 );
    and g3228 ( n13059 , n5120 , n8474 );
    xnor g3229 ( n8294 , n8052 , n11038 );
    nor g3230 ( n9116 , n8422 , n7407 );
    xnor g3231 ( n7360 , n6311 , n11568 );
    or g3232 ( n9084 , n6710 , n1197 );
    not g3233 ( n10440 , n3438 );
    and g3234 ( n1692 , n5957 , n8808 );
    not g3235 ( n6578 , n12186 );
    not g3236 ( n6966 , n9258 );
    xor g3237 ( n3913 , n8637 , n10569 );
    xnor g3238 ( n10397 , n2079 , n11153 );
    xnor g3239 ( n2830 , n7580 , n4985 );
    xnor g3240 ( n3446 , n786 , n5484 );
    and g3241 ( n13172 , n9340 , n142 );
    xnor g3242 ( n2078 , n1742 , n6893 );
    and g3243 ( n1241 , n12410 , n2802 );
    xnor g3244 ( n11070 , n1443 , n6496 );
    not g3245 ( n1858 , n4636 );
    or g3246 ( n7470 , n12575 , n5623 );
    and g3247 ( n13195 , n7481 , n10644 );
    and g3248 ( n1111 , n7686 , n4508 );
    not g3249 ( n4166 , n1198 );
    and g3250 ( n3536 , n9245 , n12866 );
    or g3251 ( n6943 , n406 , n11446 );
    and g3252 ( n10279 , n9628 , n7459 );
    and g3253 ( n4555 , n2512 , n12237 );
    xnor g3254 ( n5330 , n1481 , n11848 );
    not g3255 ( n5805 , n5605 );
    nor g3256 ( n11128 , n7601 , n3779 );
    and g3257 ( n10804 , n5540 , n1917 );
    and g3258 ( n6512 , n1056 , n3582 );
    or g3259 ( n9782 , n10281 , n2675 );
    xnor g3260 ( n9589 , n2492 , n250 );
    nor g3261 ( n8076 , n6763 , n10440 );
    not g3262 ( n1236 , n7378 );
    not g3263 ( n645 , n4570 );
    not g3264 ( n12434 , n8522 );
    xnor g3265 ( n9006 , n2072 , n12283 );
    xnor g3266 ( n4404 , n8970 , n12701 );
    not g3267 ( n3299 , n7061 );
    xnor g3268 ( n5140 , n2912 , n4900 );
    or g3269 ( n2831 , n7707 , n4947 );
    and g3270 ( n7197 , n9712 , n1592 );
    not g3271 ( n5082 , n8794 );
    and g3272 ( n3033 , n8081 , n13191 );
    not g3273 ( n4974 , n6655 );
    xnor g3274 ( n5641 , n13169 , n3083 );
    and g3275 ( n9013 , n8940 , n287 );
    or g3276 ( n8263 , n8039 , n360 );
    or g3277 ( n9221 , n10586 , n1199 );
    or g3278 ( n10144 , n2720 , n4160 );
    xor g3279 ( n1327 , n11076 , n412 );
    not g3280 ( n12629 , n1198 );
    or g3281 ( n9509 , n11736 , n2695 );
    nor g3282 ( n5663 , n141 , n13195 );
    or g3283 ( n10265 , n13116 , n3709 );
    or g3284 ( n1796 , n4654 , n1958 );
    or g3285 ( n3822 , n3972 , n11152 );
    and g3286 ( n8695 , n5220 , n11636 );
    or g3287 ( n4079 , n2437 , n6652 );
    xnor g3288 ( n2035 , n3270 , n13143 );
    xnor g3289 ( n5183 , n11374 , n9025 );
    or g3290 ( n10609 , n7900 , n8030 );
    xnor g3291 ( n12492 , n5553 , n3 );
    or g3292 ( n365 , n9397 , n9319 );
    xnor g3293 ( n10922 , n8803 , n12787 );
    or g3294 ( n7589 , n6343 , n10788 );
    and g3295 ( n10832 , n1732 , n10502 );
    nor g3296 ( n2558 , n8760 , n3209 );
    xnor g3297 ( n12594 , n2262 , n4535 );
    or g3298 ( n8883 , n6271 , n7723 );
    nor g3299 ( n7746 , n3285 , n7381 );
    nor g3300 ( n7944 , n12252 , n5573 );
    nor g3301 ( n9533 , n10318 , n530 );
    xnor g3302 ( n12307 , n12681 , n6685 );
    or g3303 ( n1827 , n694 , n12717 );
    and g3304 ( n11032 , n7244 , n7933 );
    or g3305 ( n8779 , n737 , n6404 );
    or g3306 ( n1962 , n3713 , n7962 );
    not g3307 ( n6658 , n6023 );
    nor g3308 ( n355 , n12168 , n1890 );
    xor g3309 ( n1718 , n3431 , n9717 );
    or g3310 ( n4308 , n8254 , n11107 );
    or g3311 ( n3054 , n9131 , n8030 );
    xnor g3312 ( n12006 , n6508 , n4199 );
    and g3313 ( n3879 , n7265 , n8789 );
    or g3314 ( n7699 , n7742 , n5076 );
    or g3315 ( n5811 , n3809 , n2290 );
    xnor g3316 ( n5519 , n9817 , n4014 );
    nor g3317 ( n9604 , n4130 , n1627 );
    or g3318 ( n7441 , n1779 , n10132 );
    not g3319 ( n10137 , n11222 );
    nor g3320 ( n1572 , n6990 , n974 );
    and g3321 ( n11255 , n3425 , n1028 );
    not g3322 ( n11974 , n25 );
    or g3323 ( n7022 , n3419 , n2035 );
    xnor g3324 ( n2274 , n12867 , n11079 );
    xnor g3325 ( n7879 , n9819 , n10555 );
    or g3326 ( n9085 , n9693 , n4325 );
    or g3327 ( n4239 , n12009 , n9223 );
    xnor g3328 ( n7793 , n11050 , n11401 );
    xor g3329 ( n11747 , n25 , n10724 );
    or g3330 ( n1977 , n12049 , n7935 );
    not g3331 ( n5271 , n11634 );
    or g3332 ( n5940 , n12456 , n7180 );
    or g3333 ( n11653 , n11356 , n177 );
    xnor g3334 ( n11764 , n4502 , n9458 );
    xnor g3335 ( n7514 , n7841 , n5149 );
    or g3336 ( n5814 , n11653 , n13042 );
    not g3337 ( n9730 , n2555 );
    xnor g3338 ( n3865 , n12042 , n4256 );
    not g3339 ( n79 , n9531 );
    xnor g3340 ( n9974 , n1299 , n8312 );
    xnor g3341 ( n7206 , n2371 , n3269 );
    or g3342 ( n2999 , n5563 , n11032 );
    or g3343 ( n3958 , n3761 , n1014 );
    xnor g3344 ( n11074 , n11780 , n11758 );
    nor g3345 ( n2201 , n9363 , n1566 );
    not g3346 ( n12908 , n6987 );
    not g3347 ( n8098 , n1683 );
    or g3348 ( n2491 , n477 , n5024 );
    or g3349 ( n5717 , n9240 , n7002 );
    not g3350 ( n9460 , n9115 );
    and g3351 ( n4805 , n10113 , n7113 );
    nor g3352 ( n7721 , n3659 , n8260 );
    xnor g3353 ( n12073 , n12740 , n1748 );
    not g3354 ( n8615 , n8233 );
    nor g3355 ( n6270 , n9534 , n3192 );
    or g3356 ( n9904 , n10966 , n2958 );
    or g3357 ( n433 , n5248 , n10299 );
    or g3358 ( n11150 , n7868 , n8348 );
    not g3359 ( n11750 , n4889 );
    xnor g3360 ( n12495 , n551 , n2142 );
    buf g3361 ( n206 , n2557 );
    not g3362 ( n10008 , n836 );
    or g3363 ( n10196 , n11547 , n3689 );
    not g3364 ( n10318 , n5972 );
    not g3365 ( n10272 , n10630 );
    and g3366 ( n11638 , n12919 , n10533 );
    xnor g3367 ( n340 , n1888 , n3464 );
    or g3368 ( n489 , n7501 , n11359 );
    nor g3369 ( n2749 , n1200 , n7645 );
    and g3370 ( n1956 , n10837 , n1015 );
    and g3371 ( n9493 , n7563 , n7794 );
    and g3372 ( n12654 , n9873 , n7856 );
    xnor g3373 ( n12398 , n4262 , n8124 );
    or g3374 ( n5122 , n2500 , n1371 );
    or g3375 ( n5888 , n4473 , n8490 );
    xnor g3376 ( n12929 , n2980 , n794 );
    nor g3377 ( n9432 , n2978 , n10443 );
    nor g3378 ( n3520 , n11671 , n9062 );
    not g3379 ( n1998 , n3887 );
    xor g3380 ( n7821 , n9540 , n9510 );
    and g3381 ( n7616 , n7914 , n12949 );
    and g3382 ( n8558 , n4964 , n1916 );
    xnor g3383 ( n6061 , n7117 , n7170 );
    xnor g3384 ( n12662 , n1775 , n6316 );
    xnor g3385 ( n2986 , n5272 , n5856 );
    and g3386 ( n5295 , n11127 , n2355 );
    nor g3387 ( n11023 , n4379 , n2897 );
    or g3388 ( n11985 , n4997 , n3237 );
    or g3389 ( n5284 , n1511 , n7935 );
    xnor g3390 ( n3989 , n6071 , n10829 );
    nor g3391 ( n7795 , n12322 , n12374 );
    not g3392 ( n9148 , n8916 );
    not g3393 ( n8934 , n11217 );
    xnor g3394 ( n9958 , n7236 , n2099 );
    and g3395 ( n8462 , n8042 , n2533 );
    or g3396 ( n516 , n1319 , n3984 );
    and g3397 ( n2552 , n7607 , n3501 );
    or g3398 ( n673 , n4220 , n4360 );
    or g3399 ( n10006 , n12656 , n10807 );
    xnor g3400 ( n6546 , n5888 , n9549 );
    not g3401 ( n4742 , n10105 );
    or g3402 ( n12677 , n7880 , n8348 );
    not g3403 ( n3924 , n4023 );
    or g3404 ( n8601 , n2473 , n11770 );
    and g3405 ( n586 , n1449 , n7852 );
    or g3406 ( n7510 , n2468 , n12489 );
    or g3407 ( n5528 , n5959 , n12889 );
    xnor g3408 ( n13166 , n7686 , n12436 );
    nor g3409 ( n4683 , n3741 , n3551 );
    nor g3410 ( n10672 , n5680 , n7200 );
    or g3411 ( n10427 , n928 , n3287 );
    not g3412 ( n10793 , n13020 );
    xnor g3413 ( n7058 , n5929 , n10215 );
    or g3414 ( n5655 , n107 , n5049 );
    or g3415 ( n11629 , n4657 , n6404 );
    and g3416 ( n11223 , n6008 , n10268 );
    and g3417 ( n6196 , n8251 , n12821 );
    xnor g3418 ( n4183 , n6511 , n10943 );
    or g3419 ( n10023 , n9955 , n10570 );
    and g3420 ( n7521 , n12940 , n7496 );
    or g3421 ( n5142 , n12982 , n3497 );
    or g3422 ( n3018 , n5990 , n4230 );
    nor g3423 ( n6989 , n6382 , n10175 );
    nor g3424 ( n13137 , n10113 , n1757 );
    or g3425 ( n6928 , n1977 , n9149 );
    or g3426 ( n3313 , n8249 , n6635 );
    nor g3427 ( n5982 , n6618 , n10986 );
    not g3428 ( n11969 , n12923 );
    xnor g3429 ( n4892 , n8749 , n8761 );
    or g3430 ( n5134 , n10944 , n6706 );
    and g3431 ( n6585 , n2057 , n3076 );
    not g3432 ( n8508 , n8155 );
    or g3433 ( n9479 , n227 , n8268 );
    xnor g3434 ( n6781 , n5794 , n11753 );
    or g3435 ( n3354 , n11157 , n1463 );
    nor g3436 ( n5029 , n10485 , n11856 );
    xnor g3437 ( n8149 , n4905 , n7757 );
    xnor g3438 ( n6429 , n376 , n3921 );
    or g3439 ( n4192 , n7084 , n9784 );
    nor g3440 ( n1512 , n11912 , n9715 );
    nor g3441 ( n219 , n6065 , n10852 );
    and g3442 ( n6925 , n12856 , n6821 );
    and g3443 ( n2468 , n1714 , n1475 );
    not g3444 ( n12741 , n13060 );
    xnor g3445 ( n696 , n2479 , n5078 );
    not g3446 ( n7880 , n5536 );
    not g3447 ( n11466 , n4006 );
    xnor g3448 ( n11492 , n9869 , n7168 );
    not g3449 ( n3364 , n5758 );
    xnor g3450 ( n3737 , n10967 , n13189 );
    or g3451 ( n2155 , n5937 , n4165 );
    not g3452 ( n971 , n389 );
    nor g3453 ( n4131 , n10339 , n7005 );
    not g3454 ( n2619 , n4281 );
    xnor g3455 ( n9329 , n91 , n9196 );
    xnor g3456 ( n8616 , n6610 , n4069 );
    not g3457 ( n9988 , n824 );
    xnor g3458 ( n140 , n2881 , n2751 );
    and g3459 ( n9762 , n3231 , n4175 );
    and g3460 ( n12763 , n10237 , n6472 );
    nor g3461 ( n4067 , n5502 , n11452 );
    xnor g3462 ( n998 , n8629 , n1852 );
    and g3463 ( n824 , n9157 , n11595 );
    xnor g3464 ( n5730 , n7666 , n2984 );
    and g3465 ( n7813 , n4524 , n9697 );
    or g3466 ( n6845 , n13062 , n6176 );
    and g3467 ( n9372 , n37 , n5224 );
    or g3468 ( n1661 , n1329 , n7723 );
    and g3469 ( n1584 , n3166 , n8687 );
    or g3470 ( n6627 , n9930 , n3980 );
    xnor g3471 ( n9957 , n1699 , n3731 );
    xnor g3472 ( n9566 , n8351 , n2213 );
    xor g3473 ( n865 , n10622 , n13157 );
    nor g3474 ( n12325 , n10056 , n1668 );
    and g3475 ( n826 , n2306 , n9247 );
    nor g3476 ( n6692 , n3510 , n11906 );
    not g3477 ( n11927 , n12390 );
    or g3478 ( n5369 , n2619 , n8012 );
    xnor g3479 ( n3154 , n4764 , n7138 );
    and g3480 ( n3835 , n8937 , n1141 );
    or g3481 ( n8115 , n8795 , n2959 );
    or g3482 ( n11728 , n2479 , n8292 );
    xnor g3483 ( n10494 , n6205 , n425 );
    not g3484 ( n10748 , n8954 );
    not g3485 ( n561 , n3144 );
    not g3486 ( n1333 , n5984 );
    not g3487 ( n5559 , n4691 );
    not g3488 ( n8697 , n10867 );
    xnor g3489 ( n7984 , n3478 , n10464 );
    xnor g3490 ( n195 , n5577 , n12251 );
    not g3491 ( n11757 , n22 );
    xnor g3492 ( n1382 , n3988 , n2445 );
    xnor g3493 ( n1622 , n32 , n4020 );
    and g3494 ( n6408 , n4521 , n13099 );
    xnor g3495 ( n11669 , n31 , n5051 );
    xnor g3496 ( n4925 , n7435 , n7088 );
    not g3497 ( n1869 , n854 );
    xnor g3498 ( n9052 , n5513 , n10251 );
    xnor g3499 ( n2512 , n11233 , n7736 );
    nor g3500 ( n2571 , n4277 , n3046 );
    or g3501 ( n12500 , n4298 , n8582 );
    or g3502 ( n3478 , n5461 , n6769 );
    xnor g3503 ( n471 , n9401 , n3930 );
    nor g3504 ( n5191 , n1493 , n8624 );
    or g3505 ( n7114 , n644 , n7152 );
    xnor g3506 ( n9021 , n9835 , n804 );
    and g3507 ( n9546 , n11633 , n5829 );
    and g3508 ( n6089 , n12336 , n1267 );
    or g3509 ( n181 , n588 , n7585 );
    or g3510 ( n9224 , n7110 , n9052 );
    or g3511 ( n1104 , n3381 , n4819 );
    not g3512 ( n1889 , n11049 );
    and g3513 ( n2962 , n8666 , n6204 );
    not g3514 ( n10256 , n4470 );
    and g3515 ( n10367 , n10717 , n12874 );
    xnor g3516 ( n13061 , n2771 , n6168 );
    xnor g3517 ( n6090 , n8785 , n197 );
    not g3518 ( n6008 , n13006 );
    not g3519 ( n8419 , n7932 );
    not g3520 ( n9170 , n8713 );
    xnor g3521 ( n468 , n3744 , n9184 );
    and g3522 ( n6999 , n5412 , n10340 );
    or g3523 ( n2220 , n1058 , n12847 );
    nor g3524 ( n8247 , n7421 , n981 );
    nor g3525 ( n3119 , n6794 , n5812 );
    xnor g3526 ( n1510 , n548 , n2369 );
    xnor g3527 ( n8867 , n2151 , n105 );
    xnor g3528 ( n3897 , n10905 , n3626 );
    or g3529 ( n12944 , n9396 , n9311 );
    not g3530 ( n5588 , n10594 );
    or g3531 ( n8157 , n11683 , n11144 );
    not g3532 ( n8463 , n10142 );
    or g3533 ( n4229 , n4271 , n9348 );
    or g3534 ( n4094 , n11078 , n7837 );
    or g3535 ( n10435 , n1145 , n10892 );
    not g3536 ( n10266 , n12605 );
    and g3537 ( n11067 , n5675 , n4559 );
    not g3538 ( n7787 , n5453 );
    or g3539 ( n7128 , n10402 , n10319 );
    xnor g3540 ( n3234 , n10785 , n429 );
    and g3541 ( n3839 , n11447 , n12765 );
    and g3542 ( n11756 , n5069 , n123 );
    xnor g3543 ( n9536 , n4663 , n8056 );
    nor g3544 ( n10855 , n7920 , n11034 );
    xnor g3545 ( n6623 , n12039 , n4182 );
    not g3546 ( n4844 , n10606 );
    and g3547 ( n6914 , n7668 , n8074 );
    or g3548 ( n13041 , n4785 , n7615 );
    or g3549 ( n6359 , n10462 , n4724 );
    or g3550 ( n6452 , n552 , n3376 );
    or g3551 ( n263 , n971 , n2958 );
    xnor g3552 ( n7644 , n7690 , n199 );
    or g3553 ( n3382 , n4290 , n6364 );
    nor g3554 ( n11287 , n8812 , n5287 );
    xor g3555 ( n12980 , n6155 , n10670 );
    not g3556 ( n6825 , n11112 );
    or g3557 ( n3020 , n5194 , n5272 );
    or g3558 ( n11033 , n8529 , n6404 );
    not g3559 ( n1000 , n1600 );
    not g3560 ( n7608 , n13060 );
    xor g3561 ( n1286 , n11096 , n12424 );
    not g3562 ( n8097 , n2920 );
    not g3563 ( n9677 , n3121 );
    and g3564 ( n6601 , n7561 , n4970 );
    or g3565 ( n2223 , n8379 , n5273 );
    or g3566 ( n9540 , n2420 , n2287 );
    nor g3567 ( n5376 , n1507 , n3519 );
    xnor g3568 ( n11046 , n2184 , n5486 );
    xnor g3569 ( n8861 , n6688 , n8471 );
    and g3570 ( n4042 , n7791 , n6469 );
    xnor g3571 ( n92 , n823 , n7928 );
    not g3572 ( n11037 , n5065 );
    xnor g3573 ( n6660 , n1398 , n1946 );
    xnor g3574 ( n5754 , n6359 , n4255 );
    nor g3575 ( n10534 , n7709 , n3165 );
    not g3576 ( n7410 , n8735 );
    and g3577 ( n3110 , n5249 , n3614 );
    xnor g3578 ( n838 , n6021 , n8227 );
    or g3579 ( n4759 , n391 , n12978 );
    xnor g3580 ( n6555 , n3171 , n9665 );
    xnor g3581 ( n7790 , n10904 , n10777 );
    xnor g3582 ( n9522 , n8881 , n3596 );
    or g3583 ( n12764 , n9162 , n8702 );
    xnor g3584 ( n8013 , n6740 , n9141 );
    or g3585 ( n9878 , n5152 , n4495 );
    or g3586 ( n5334 , n5990 , n7221 );
    not g3587 ( n6309 , n11900 );
    or g3588 ( n3077 , n182 , n5295 );
    xnor g3589 ( n885 , n477 , n8554 );
    nor g3590 ( n5859 , n3441 , n6909 );
    or g3591 ( n996 , n5670 , n7642 );
    and g3592 ( n4232 , n11946 , n11481 );
    xnor g3593 ( n12110 , n2043 , n5995 );
    not g3594 ( n13043 , n9941 );
    not g3595 ( n5806 , n1724 );
    xnor g3596 ( n6816 , n7546 , n3610 );
    nor g3597 ( n4961 , n8864 , n2422 );
    and g3598 ( n539 , n4594 , n7588 );
    nor g3599 ( n4730 , n2304 , n10961 );
    xor g3600 ( n1491 , n8455 , n2229 );
    and g3601 ( n6387 , n7599 , n9037 );
    and g3602 ( n4244 , n2883 , n1506 );
    or g3603 ( n11918 , n7041 , n8348 );
    and g3604 ( n661 , n373 , n12309 );
    and g3605 ( n11659 , n3628 , n1173 );
    not g3606 ( n7234 , n12263 );
    xnor g3607 ( n4993 , n7575 , n8145 );
    and g3608 ( n9466 , n5870 , n528 );
    nor g3609 ( n7737 , n577 , n2117 );
    xnor g3610 ( n1405 , n7095 , n9117 );
    xnor g3611 ( n4162 , n2792 , n12911 );
    not g3612 ( n3791 , n10811 );
    and g3613 ( n12442 , n12384 , n7383 );
    and g3614 ( n5775 , n2769 , n9660 );
    not g3615 ( n308 , n2539 );
    xnor g3616 ( n3107 , n11865 , n4895 );
    or g3617 ( n12901 , n7890 , n10761 );
    or g3618 ( n5077 , n3839 , n11346 );
    or g3619 ( n10862 , n4021 , n3434 );
    xnor g3620 ( n12987 , n2940 , n5741 );
    xnor g3621 ( n6665 , n1095 , n9028 );
    or g3622 ( n4635 , n8882 , n1850 );
    not g3623 ( n13071 , n4349 );
    not g3624 ( n13086 , n11537 );
    and g3625 ( n12120 , n9590 , n6509 );
    xnor g3626 ( n2535 , n10373 , n10091 );
    xnor g3627 ( n5195 , n3050 , n3170 );
    or g3628 ( n4390 , n10462 , n2133 );
    not g3629 ( n7254 , n11488 );
    or g3630 ( n7752 , n11941 , n8348 );
    or g3631 ( n7649 , n11159 , n10040 );
    nor g3632 ( n4070 , n9641 , n4873 );
    xnor g3633 ( n4578 , n11444 , n3198 );
    xnor g3634 ( n8014 , n455 , n5104 );
    xnor g3635 ( n12857 , n9830 , n4283 );
    nor g3636 ( n9251 , n6505 , n13037 );
    not g3637 ( n8786 , n862 );
    nor g3638 ( n7292 , n1807 , n6281 );
    or g3639 ( n8245 , n2332 , n177 );
    and g3640 ( n10311 , n9933 , n7193 );
    or g3641 ( n10906 , n8672 , n9195 );
    not g3642 ( n8341 , n11079 );
    xnor g3643 ( n10087 , n5181 , n9295 );
    xnor g3644 ( n2865 , n5102 , n4051 );
    or g3645 ( n4072 , n5695 , n7339 );
    and g3646 ( n6216 , n4850 , n2499 );
    or g3647 ( n8302 , n755 , n12967 );
    xnor g3648 ( n12761 , n10774 , n5779 );
    xnor g3649 ( n4681 , n10547 , n7323 );
    not g3650 ( n5583 , n3152 );
    or g3651 ( n12233 , n11137 , n10319 );
    not g3652 ( n4979 , n6168 );
    not g3653 ( n7678 , n12025 );
    xnor g3654 ( n7875 , n2435 , n12554 );
    xnor g3655 ( n11848 , n9750 , n504 );
    not g3656 ( n11239 , n9531 );
    or g3657 ( n9439 , n2736 , n2659 );
    and g3658 ( n11254 , n13001 , n5155 );
    or g3659 ( n3013 , n12786 , n8534 );
    or g3660 ( n8061 , n5595 , n7530 );
    and g3661 ( n7959 , n3945 , n10495 );
    and g3662 ( n9655 , n2482 , n12853 );
    or g3663 ( n8949 , n13012 , n12188 );
    and g3664 ( n2821 , n8183 , n6085 );
    xnor g3665 ( n9248 , n2813 , n4691 );
    or g3666 ( n8648 , n935 , n2133 );
    xnor g3667 ( n4100 , n4377 , n5439 );
    and g3668 ( n1222 , n1801 , n2477 );
    not g3669 ( n4490 , n9915 );
    and g3670 ( n4448 , n9486 , n6738 );
    or g3671 ( n3744 , n12469 , n12957 );
    nor g3672 ( n12131 , n1580 , n9463 );
    xnor g3673 ( n5298 , n8651 , n2951 );
    and g3674 ( n5343 , n10142 , n5962 );
    and g3675 ( n13112 , n11336 , n5318 );
    or g3676 ( n10022 , n6016 , n8782 );
    not g3677 ( n1832 , n6879 );
    xnor g3678 ( n7024 , n5233 , n12934 );
    or g3679 ( n6956 , n10761 , n4936 );
    or g3680 ( n2191 , n1795 , n8543 );
    or g3681 ( n3932 , n11196 , n9533 );
    and g3682 ( n7394 , n2992 , n11262 );
    xnor g3683 ( n1839 , n3749 , n801 );
    and g3684 ( n2672 , n11576 , n8839 );
    and g3685 ( n12974 , n2902 , n1189 );
    or g3686 ( n8424 , n7191 , n5939 );
    nor g3687 ( n4056 , n1025 , n4482 );
    xnor g3688 ( n1140 , n12229 , n4019 );
    not g3689 ( n1787 , n10002 );
    xnor g3690 ( n1948 , n10538 , n5650 );
    or g3691 ( n10964 , n667 , n5693 );
    or g3692 ( n13014 , n4981 , n9110 );
    or g3693 ( n9649 , n8060 , n3229 );
    xnor g3694 ( n9452 , n3458 , n2964 );
    nor g3695 ( n10664 , n12204 , n12235 );
    or g3696 ( n12206 , n4039 , n9188 );
    or g3697 ( n12312 , n12483 , n4194 );
    xnor g3698 ( n40 , n6013 , n5232 );
    xnor g3699 ( n11196 , n159 , n6154 );
    and g3700 ( n10414 , n5200 , n12979 );
    and g3701 ( n12842 , n11624 , n5338 );
    nor g3702 ( n2517 , n6310 , n4414 );
    xnor g3703 ( n12329 , n6460 , n5362 );
    xnor g3704 ( n10796 , n12707 , n10699 );
    or g3705 ( n9279 , n12092 , n10982 );
    or g3706 ( n10716 , n1925 , n4407 );
    and g3707 ( n9120 , n2480 , n5877 );
    or g3708 ( n6000 , n3354 , n6730 );
    nor g3709 ( n8423 , n8742 , n4816 );
    and g3710 ( n1608 , n5665 , n8454 );
    or g3711 ( n5803 , n1589 , n2133 );
    and g3712 ( n9344 , n5732 , n5504 );
    xnor g3713 ( n5236 , n7697 , n4615 );
    and g3714 ( n5067 , n151 , n7078 );
    not g3715 ( n5455 , n11429 );
    nor g3716 ( n9301 , n10865 , n1004 );
    and g3717 ( n4628 , n7437 , n12124 );
    nor g3718 ( n8162 , n1469 , n7054 );
    not g3719 ( n8006 , n5969 );
    or g3720 ( n5898 , n2742 , n90 );
    and g3721 ( n11059 , n2085 , n2149 );
    or g3722 ( n4174 , n5322 , n5222 );
    not g3723 ( n10772 , n12965 );
    or g3724 ( n3753 , n10437 , n11107 );
    not g3725 ( n10066 , n7945 );
    nor g3726 ( n7185 , n9508 , n10910 );
    xnor g3727 ( n3369 , n3192 , n8515 );
    not g3728 ( n2942 , n11061 );
    or g3729 ( n1252 , n7642 , n479 );
    or g3730 ( n2363 , n9305 , n10179 );
    not g3731 ( n5468 , n11991 );
    or g3732 ( n7193 , n2884 , n5797 );
    not g3733 ( n546 , n6236 );
    or g3734 ( n4761 , n9402 , n4333 );
    or g3735 ( n3836 , n4179 , n2059 );
    and g3736 ( n5500 , n2460 , n4750 );
    nor g3737 ( n547 , n7161 , n1144 );
    and g3738 ( n12818 , n10233 , n6218 );
    not g3739 ( n1126 , n9097 );
    or g3740 ( n8927 , n1222 , n10239 );
    not g3741 ( n10739 , n2023 );
    nor g3742 ( n5789 , n11711 , n41 );
    or g3743 ( n3833 , n5492 , n13135 );
    xor g3744 ( n7996 , n6682 , n6451 );
    and g3745 ( n799 , n11512 , n4869 );
    or g3746 ( n7461 , n6401 , n306 );
    not g3747 ( n11535 , n2595 );
    not g3748 ( n8562 , n3409 );
    or g3749 ( n6057 , n349 , n11283 );
    not g3750 ( n6225 , n4335 );
    xnor g3751 ( n4994 , n8932 , n9204 );
    or g3752 ( n9157 , n689 , n4626 );
    or g3753 ( n2373 , n823 , n4405 );
    and g3754 ( n9258 , n3588 , n5967 );
    not g3755 ( n11225 , n2174 );
    and g3756 ( n3809 , n6222 , n3101 );
    xnor g3757 ( n2638 , n8920 , n12678 );
    and g3758 ( n10820 , n13141 , n11088 );
    or g3759 ( n3348 , n542 , n2675 );
    nor g3760 ( n6227 , n386 , n6482 );
    xnor g3761 ( n6686 , n8850 , n632 );
    or g3762 ( n2870 , n7385 , n12794 );
    nor g3763 ( n1053 , n2975 , n12056 );
    not g3764 ( n12948 , n834 );
    or g3765 ( n771 , n9129 , n6404 );
    and g3766 ( n5907 , n10182 , n12532 );
    not g3767 ( n6004 , n4685 );
    xor g3768 ( n10434 , n8876 , n3180 );
    not g3769 ( n6568 , n2233 );
    or g3770 ( n9392 , n10893 , n1144 );
    nor g3771 ( n2835 , n12553 , n4350 );
    or g3772 ( n5845 , n2462 , n8563 );
    not g3773 ( n8077 , n11760 );
    or g3774 ( n10373 , n4161 , n7221 );
    or g3775 ( n8994 , n2129 , n7221 );
    or g3776 ( n9040 , n7243 , n11232 );
    or g3777 ( n12668 , n12963 , n4812 );
    and g3778 ( n12774 , n9620 , n8716 );
    or g3779 ( n2105 , n9703 , n9064 );
    not g3780 ( n1999 , n2445 );
    xnor g3781 ( n11881 , n6467 , n11112 );
    xnor g3782 ( n12887 , n5394 , n4140 );
    not g3783 ( n5423 , n8233 );
    nor g3784 ( n1316 , n11023 , n3462 );
    xnor g3785 ( n12883 , n3976 , n1884 );
    not g3786 ( n2296 , n12289 );
    xnor g3787 ( n6224 , n3623 , n8917 );
    xnor g3788 ( n11732 , n9258 , n4234 );
    not g3789 ( n1769 , n12594 );
    xnor g3790 ( n5447 , n1494 , n9297 );
    or g3791 ( n8318 , n8957 , n581 );
    not g3792 ( n8249 , n5536 );
    not g3793 ( n4660 , n11607 );
    and g3794 ( n10962 , n2851 , n1072 );
    nor g3795 ( n5327 , n9150 , n8743 );
    and g3796 ( n8974 , n2068 , n11109 );
    or g3797 ( n4016 , n7396 , n4230 );
    xnor g3798 ( n5628 , n1408 , n2239 );
    nor g3799 ( n12710 , n2143 , n8527 );
    and g3800 ( n6312 , n3827 , n5021 );
    buf g3801 ( n8563 , n3169 );
    xnor g3802 ( n6087 , n11371 , n2336 );
    not g3803 ( n3646 , n3769 );
    xnor g3804 ( n302 , n11590 , n11205 );
    xnor g3805 ( n9188 , n8412 , n273 );
    nor g3806 ( n7633 , n3581 , n6331 );
    not g3807 ( n950 , n7448 );
    xnor g3808 ( n9480 , n3818 , n12040 );
    nor g3809 ( n8682 , n11436 , n5053 );
    xnor g3810 ( n6347 , n12428 , n4435 );
    nor g3811 ( n13100 , n8738 , n5997 );
    xnor g3812 ( n6483 , n6619 , n637 );
    or g3813 ( n300 , n4464 , n11107 );
    nor g3814 ( n2522 , n11223 , n3002 );
    not g3815 ( n11101 , n6668 );
    not g3816 ( n5547 , n9906 );
    or g3817 ( n12572 , n8839 , n11576 );
    not g3818 ( n2604 , n9412 );
    not g3819 ( n10689 , n10027 );
    xnor g3820 ( n11162 , n12121 , n10458 );
    xnor g3821 ( n7628 , n9033 , n12743 );
    and g3822 ( n864 , n761 , n11058 );
    or g3823 ( n3720 , n11116 , n7976 );
    not g3824 ( n795 , n11411 );
    xor g3825 ( n573 , n1065 , n7238 );
    not g3826 ( n3340 , n7541 );
    and g3827 ( n9578 , n1505 , n2482 );
    not g3828 ( n2599 , n8290 );
    nor g3829 ( n8568 , n12518 , n3041 );
    xnor g3830 ( n4520 , n7311 , n12438 );
    not g3831 ( n11088 , n5228 );
    not g3832 ( n5107 , n401 );
    not g3833 ( n5685 , n9092 );
    xnor g3834 ( n3314 , n5523 , n2818 );
    and g3835 ( n498 , n7257 , n3450 );
    or g3836 ( n11624 , n12802 , n4295 );
    or g3837 ( n4276 , n11226 , n10106 );
    and g3838 ( n3709 , n8541 , n1264 );
    or g3839 ( n534 , n12971 , n7344 );
    and g3840 ( n12470 , n6313 , n7321 );
    and g3841 ( n5681 , n11847 , n7469 );
    or g3842 ( n1099 , n3553 , n2544 );
    or g3843 ( n10219 , n1370 , n7075 );
    or g3844 ( n12078 , n2416 , n2133 );
    xor g3845 ( n1057 , n1214 , n11861 );
    or g3846 ( n4958 , n1394 , n3233 );
    or g3847 ( n6176 , n8510 , n177 );
    or g3848 ( n1085 , n7167 , n7935 );
    or g3849 ( n7081 , n3453 , n5335 );
    not g3850 ( n13228 , n2898 );
    or g3851 ( n2179 , n11674 , n7092 );
    xnor g3852 ( n5837 , n7554 , n140 );
    xor g3853 ( n1836 , n2255 , n9652 );
    nor g3854 ( n2405 , n7448 , n194 );
    xnor g3855 ( n5994 , n5730 , n6122 );
    and g3856 ( n1610 , n2326 , n2267 );
    nor g3857 ( n7756 , n8001 , n7352 );
    not g3858 ( n1781 , n2668 );
    or g3859 ( n5752 , n6769 , n6404 );
    and g3860 ( n8106 , n11903 , n5765 );
    not g3861 ( n2919 , n834 );
    and g3862 ( n8876 , n12343 , n768 );
    not g3863 ( n2420 , n2758 );
    or g3864 ( n1435 , n7119 , n1570 );
    xnor g3865 ( n8021 , n7245 , n7007 );
    and g3866 ( n6523 , n1976 , n7586 );
    xnor g3867 ( n12534 , n4215 , n3983 );
    xnor g3868 ( n477 , n4016 , n843 );
    and g3869 ( n10053 , n997 , n970 );
    xnor g3870 ( n7668 , n7279 , n4532 );
    and g3871 ( n405 , n9569 , n10746 );
    not g3872 ( n9745 , n287 );
    and g3873 ( n5093 , n5801 , n9475 );
    not g3874 ( n4514 , n3130 );
    nor g3875 ( n2017 , n1847 , n10090 );
    xnor g3876 ( n12979 , n2918 , n7259 );
    xor g3877 ( n3880 , n5705 , n10078 );
    not g3878 ( n5080 , n635 );
    nor g3879 ( n10732 , n3219 , n739 );
    or g3880 ( n6184 , n2678 , n9195 );
    or g3881 ( n2257 , n6503 , n310 );
    and g3882 ( n8888 , n8139 , n5920 );
    or g3883 ( n7565 , n11437 , n10693 );
    and g3884 ( n4278 , n4886 , n7810 );
    and g3885 ( n4399 , n8704 , n10529 );
    or g3886 ( n7975 , n9305 , n7530 );
    xnor g3887 ( n3323 , n486 , n1341 );
    or g3888 ( n2269 , n1234 , n1934 );
    or g3889 ( n9428 , n10761 , n10433 );
    or g3890 ( n6974 , n946 , n1985 );
    xnor g3891 ( n8461 , n8125 , n1138 );
    not g3892 ( n12180 , n3860 );
    and g3893 ( n12479 , n12592 , n2882 );
    nor g3894 ( n595 , n10384 , n384 );
    or g3895 ( n10713 , n4132 , n12847 );
    and g3896 ( n8918 , n2204 , n1546 );
    and g3897 ( n283 , n13062 , n6176 );
    nor g3898 ( n9406 , n3155 , n8656 );
    or g3899 ( n4901 , n1524 , n9778 );
    xnor g3900 ( n1010 , n1862 , n1283 );
    xnor g3901 ( n5945 , n10859 , n11631 );
    and g3902 ( n8327 , n12899 , n7710 );
    or g3903 ( n10894 , n9806 , n7224 );
    or g3904 ( n6946 , n11195 , n10110 );
    xnor g3905 ( n6718 , n10543 , n10955 );
    xnor g3906 ( n3212 , n2160 , n6198 );
    not g3907 ( n1477 , n7359 );
    not g3908 ( n2637 , n11030 );
    xnor g3909 ( n10033 , n6925 , n9394 );
    and g3910 ( n6275 , n3669 , n3085 );
    or g3911 ( n149 , n12159 , n8374 );
    xnor g3912 ( n3207 , n10198 , n2832 );
    xnor g3913 ( n9883 , n4170 , n1631 );
    xnor g3914 ( n9908 , n5331 , n2518 );
    and g3915 ( n4269 , n10113 , n12853 );
    and g3916 ( n892 , n5088 , n5814 );
    and g3917 ( n2150 , n11899 , n383 );
    and g3918 ( n2715 , n12592 , n11058 );
    and g3919 ( n8724 , n1866 , n8420 );
    or g3920 ( n9264 , n5176 , n7868 );
    not g3921 ( n11078 , n6168 );
    or g3922 ( n12362 , n12741 , n8702 );
    xnor g3923 ( n2365 , n5193 , n5643 );
    and g3924 ( n12988 , n3829 , n11685 );
    or g3925 ( n3355 , n12268 , n12401 );
    or g3926 ( n11245 , n2688 , n10179 );
    xor g3927 ( n1529 , n8102 , n7717 );
    not g3928 ( n13094 , n1983 );
    nor g3929 ( n7601 , n8284 , n4543 );
    not g3930 ( n12062 , n2590 );
    not g3931 ( n628 , n12289 );
    or g3932 ( n2785 , n10730 , n479 );
    or g3933 ( n9184 , n1188 , n4230 );
    and g3934 ( n3342 , n6333 , n10063 );
    and g3935 ( n11794 , n7502 , n11722 );
    xnor g3936 ( n1682 , n10255 , n12985 );
    not g3937 ( n10982 , n11027 );
    nor g3938 ( n12649 , n7472 , n10723 );
    not g3939 ( n12680 , n1660 );
    or g3940 ( n9263 , n11523 , n6230 );
    nor g3941 ( n1159 , n10786 , n7452 );
    nor g3942 ( n12177 , n7051 , n12820 );
    xnor g3943 ( n466 , n7904 , n6 );
    nor g3944 ( n1819 , n5453 , n9293 );
    not g3945 ( n2722 , n9163 );
    or g3946 ( n883 , n6671 , n6441 );
    xnor g3947 ( n10415 , n10917 , n4163 );
    not g3948 ( n6220 , n7812 );
    xnor g3949 ( n9315 , n4667 , n7423 );
    nor g3950 ( n3777 , n8595 , n7753 );
    xnor g3951 ( n3954 , n1714 , n3788 );
    or g3952 ( n8146 , n7408 , n8869 );
    nor g3953 ( n5986 , n10656 , n9292 );
    not g3954 ( n12204 , n1253 );
    and g3955 ( n6694 , n11696 , n7854 );
    and g3956 ( n9155 , n4727 , n13196 );
    xnor g3957 ( n12494 , n6491 , n8699 );
    nor g3958 ( n4500 , n12564 , n295 );
    xnor g3959 ( n4603 , n10533 , n12919 );
    and g3960 ( n12156 , n10199 , n5579 );
    xnor g3961 ( n1837 , n7673 , n55 );
    xnor g3962 ( n4297 , n1679 , n7042 );
    xor g3963 ( n2111 , n4411 , n388 );
    and g3964 ( n4255 , n2491 , n3529 );
    or g3965 ( n2471 , n7674 , n532 );
    and g3966 ( n3211 , n11665 , n2737 );
    or g3967 ( n12697 , n5478 , n479 );
    not g3968 ( n9658 , n2987 );
    xnor g3969 ( n4190 , n1279 , n5831 );
    or g3970 ( n4975 , n10592 , n1404 );
    xnor g3971 ( n11038 , n11182 , n2932 );
    or g3972 ( n1607 , n7507 , n3320 );
    not g3973 ( n3651 , n3875 );
    and g3974 ( n8628 , n5568 , n7113 );
    nor g3975 ( n4556 , n12631 , n2421 );
    nor g3976 ( n8783 , n11561 , n1423 );
    not g3977 ( n5017 , n12245 );
    xnor g3978 ( n257 , n2429 , n7014 );
    or g3979 ( n3365 , n5838 , n9587 );
    not g3980 ( n12522 , n1535 );
    not g3981 ( n10090 , n9419 );
    and g3982 ( n8354 , n11334 , n8627 );
    xnor g3983 ( n5123 , n11699 , n4806 );
    not g3984 ( n1728 , n646 );
    not g3985 ( n9309 , n5536 );
    not g3986 ( n2640 , n137 );
    or g3987 ( n2214 , n10447 , n5076 );
    xnor g3988 ( n5193 , n7189 , n5195 );
    and g3989 ( n12163 , n4605 , n4134 );
    xnor g3990 ( n647 , n9425 , n1146 );
    xnor g3991 ( n10366 , n5706 , n403 );
    xnor g3992 ( n5397 , n9677 , n2541 );
    not g3993 ( n1420 , n10333 );
    or g3994 ( n5957 , n9890 , n4343 );
    and g3995 ( n1746 , n10306 , n5114 );
    and g3996 ( n7316 , n3338 , n1171 );
    and g3997 ( n6847 , n9783 , n7391 );
    or g3998 ( n5653 , n10839 , n368 );
    or g3999 ( n679 , n7522 , n8268 );
    or g4000 ( n5098 , n12871 , n6265 );
    and g4001 ( n7559 , n8310 , n7187 );
    and g4002 ( n10419 , n6756 , n9565 );
    xor g4003 ( n6926 , n13221 , n78 );
    or g4004 ( n6886 , n5968 , n8702 );
    or g4005 ( n686 , n12881 , n9195 );
    and g4006 ( n9683 , n592 , n914 );
    xnor g4007 ( n3115 , n6492 , n8217 );
    not g4008 ( n4360 , n5596 );
    and g4009 ( n8274 , n12636 , n7009 );
    xnor g4010 ( n11293 , n2920 , n11937 );
    and g4011 ( n8567 , n10322 , n4604 );
    xnor g4012 ( n6574 , n1922 , n11850 );
    or g4013 ( n9502 , n4974 , n12188 );
    or g4014 ( n8368 , n6519 , n12273 );
    xnor g4015 ( n8309 , n5857 , n6177 );
    and g4016 ( n7733 , n4627 , n3279 );
    nor g4017 ( n4328 , n4533 , n12976 );
    xnor g4018 ( n5068 , n9890 , n8117 );
    xnor g4019 ( n10009 , n5956 , n6803 );
    not g4020 ( n10661 , n5404 );
    xnor g4021 ( n1060 , n11773 , n5026 );
    or g4022 ( n5390 , n3970 , n320 );
    or g4023 ( n7638 , n5152 , n10552 );
    xnor g4024 ( n9343 , n1425 , n4613 );
    and g4025 ( n4343 , n12818 , n7680 );
    not g4026 ( n12491 , n608 );
    nor g4027 ( n11220 , n10026 , n4542 );
    or g4028 ( n4513 , n5047 , n10364 );
    and g4029 ( n10138 , n12872 , n12817 );
    and g4030 ( n6829 , n7991 , n3899 );
    nor g4031 ( n9130 , n246 , n11942 );
    or g4032 ( n9496 , n3534 , n5242 );
    xnor g4033 ( n4731 , n7011 , n6061 );
    and g4034 ( n3632 , n6466 , n5512 );
    xnor g4035 ( n10782 , n5799 , n4721 );
    not g4036 ( n2877 , n12263 );
    not g4037 ( n776 , n10451 );
    xnor g4038 ( n5646 , n7035 , n4906 );
    xnor g4039 ( n1689 , n7110 , n7614 );
    or g4040 ( n2178 , n3191 , n3423 );
    and g4041 ( n10626 , n951 , n10063 );
    and g4042 ( n5769 , n5365 , n8749 );
    and g4043 ( n5208 , n12813 , n2361 );
    nor g4044 ( n9626 , n10236 , n12438 );
    xnor g4045 ( n3016 , n7550 , n3948 );
    or g4046 ( n2598 , n5611 , n9159 );
    xnor g4047 ( n12796 , n5669 , n5568 );
    not g4048 ( n6110 , n649 );
    not g4049 ( n12621 , n3769 );
    and g4050 ( n2547 , n6333 , n3085 );
    not g4051 ( n5041 , n10168 );
    not g4052 ( n3618 , n12898 );
    or g4053 ( n9930 , n11808 , n6770 );
    and g4054 ( n10274 , n11272 , n5181 );
    xnor g4055 ( n8572 , n8467 , n1263 );
    xnor g4056 ( n12149 , n4374 , n7160 );
    or g4057 ( n5871 , n12203 , n9075 );
    and g4058 ( n11616 , n9120 , n1099 );
    or g4059 ( n4625 , n3225 , n12388 );
    not g4060 ( n2440 , n5143 );
    nor g4061 ( n1485 , n6171 , n5532 );
    not g4062 ( n12066 , n11267 );
    nor g4063 ( n10514 , n3293 , n10866 );
    xnor g4064 ( n1174 , n4715 , n913 );
    xnor g4065 ( n12144 , n11335 , n1280 );
    not g4066 ( n423 , n691 );
    xor g4067 ( n7778 , n5879 , n13176 );
    or g4068 ( n7629 , n2545 , n9495 );
    xnor g4069 ( n9327 , n11460 , n4962 );
    xnor g4070 ( n3457 , n8165 , n12191 );
    xnor g4071 ( n9862 , n1855 , n11315 );
    xnor g4072 ( n9563 , n191 , n3378 );
    nor g4073 ( n1368 , n11963 , n1924 );
    nor g4074 ( n7007 , n4346 , n1643 );
    not g4075 ( n3407 , n11396 );
    xnor g4076 ( n3059 , n1983 , n4672 );
    and g4077 ( n6610 , n7089 , n12624 );
    not g4078 ( n4426 , n9621 );
    or g4079 ( n10104 , n5359 , n6987 );
    nor g4080 ( n5267 , n8513 , n10750 );
    or g4081 ( n6489 , n1089 , n2449 );
    and g4082 ( n12823 , n9298 , n8127 );
    xnor g4083 ( n8265 , n6317 , n6134 );
    or g4084 ( n8715 , n2449 , n12328 );
    xnor g4085 ( n319 , n7065 , n2526 );
    nor g4086 ( n9164 , n10280 , n8649 );
    and g4087 ( n9595 , n1260 , n8418 );
    not g4088 ( n3853 , n11055 );
    xor g4089 ( n1873 , n8788 , n9202 );
    and g4090 ( n3199 , n12668 , n6449 );
    or g4091 ( n390 , n3248 , n65 );
    not g4092 ( n4221 , n5470 );
    nor g4093 ( n4421 , n408 , n5472 );
    or g4094 ( n10738 , n11664 , n10715 );
    or g4095 ( n12012 , n11003 , n8044 );
    and g4096 ( n11091 , n8139 , n854 );
    xnor g4097 ( n7985 , n11836 , n5396 );
    or g4098 ( n11499 , n5157 , n6769 );
    or g4099 ( n12600 , n9146 , n11802 );
    xnor g4100 ( n12743 , n5843 , n6621 );
    nor g4101 ( n4355 , n10890 , n4090 );
    or g4102 ( n6697 , n5433 , n8348 );
    xnor g4103 ( n1946 , n1099 , n9120 );
    or g4104 ( n7852 , n9019 , n12695 );
    and g4105 ( n6728 , n13049 , n13115 );
    xnor g4106 ( n857 , n12055 , n12900 );
    not g4107 ( n2789 , n10568 );
    xnor g4108 ( n5765 , n9929 , n5501 );
    or g4109 ( n5745 , n1324 , n4315 );
    xnor g4110 ( n12507 , n7412 , n5164 );
    not g4111 ( n4220 , n1617 );
    not g4112 ( n1524 , n3303 );
    or g4113 ( n3980 , n6883 , n10319 );
    not g4114 ( n2148 , n9591 );
    or g4115 ( n12050 , n3259 , n4936 );
    and g4116 ( n11075 , n1034 , n12777 );
    xnor g4117 ( n7458 , n10262 , n11504 );
    not g4118 ( n4649 , n5920 );
    xnor g4119 ( n11739 , n5127 , n10976 );
    xnor g4120 ( n9523 , n9264 , n2400 );
    not g4121 ( n10321 , n13053 );
    xnor g4122 ( n7496 , n4770 , n5777 );
    xnor g4123 ( n7763 , n12192 , n5571 );
    and g4124 ( n8279 , n4798 , n10519 );
    nor g4125 ( n1303 , n3214 , n7173 );
    or g4126 ( n1905 , n3599 , n773 );
    or g4127 ( n12293 , n1052 , n3963 );
    xnor g4128 ( n3125 , n7944 , n8726 );
    nor g4129 ( n12606 , n12085 , n2071 );
    xnor g4130 ( n12350 , n1812 , n3567 );
    and g4131 ( n8084 , n5801 , n5920 );
    or g4132 ( n5571 , n11113 , n2059 );
    or g4133 ( n4664 , n9796 , n11794 );
    or g4134 ( n1496 , n1696 , n1571 );
    not g4135 ( n1290 , n8328 );
    or g4136 ( n6241 , n8889 , n12068 );
    xnor g4137 ( n9815 , n9529 , n5963 );
    xnor g4138 ( n6471 , n878 , n6087 );
    not g4139 ( n3094 , n6292 );
    not g4140 ( n12023 , n401 );
    not g4141 ( n10300 , n9446 );
    xnor g4142 ( n4324 , n12960 , n611 );
    and g4143 ( n13118 , n7295 , n9530 );
    or g4144 ( n2578 , n9004 , n9946 );
    or g4145 ( n4580 , n7957 , n5495 );
    and g4146 ( n689 , n4694 , n4986 );
    and g4147 ( n1383 , n6335 , n6221 );
    not g4148 ( n3210 , n12943 );
    or g4149 ( n6441 , n8315 , n8348 );
    and g4150 ( n12666 , n6556 , n4635 );
    or g4151 ( n907 , n9675 , n12388 );
    or g4152 ( n11744 , n8532 , n7723 );
    or g4153 ( n1054 , n8710 , n10933 );
    and g4154 ( n478 , n4316 , n2924 );
    nor g4155 ( n12917 , n4241 , n1794 );
    not g4156 ( n3553 , n12651 );
    or g4157 ( n11175 , n11785 , n639 );
    nor g4158 ( n3050 , n4159 , n11532 );
    xnor g4159 ( n11709 , n6962 , n11918 );
    nor g4160 ( n5450 , n491 , n2990 );
    not g4161 ( n579 , n12701 );
    or g4162 ( n5449 , n586 , n1770 );
    or g4163 ( n7913 , n1491 , n8242 );
    not g4164 ( n3962 , n3832 );
    and g4165 ( n6874 , n3700 , n7750 );
    xnor g4166 ( n6708 , n10912 , n572 );
    or g4167 ( n9101 , n2420 , n9159 );
    xnor g4168 ( n4793 , n6880 , n2957 );
    xnor g4169 ( n11805 , n3212 , n918 );
    and g4170 ( n1503 , n2777 , n9570 );
    or g4171 ( n6796 , n12014 , n653 );
    or g4172 ( n421 , n2848 , n1463 );
    not g4173 ( n12997 , n8506 );
    not g4174 ( n7311 , n10236 );
    or g4175 ( n2390 , n5899 , n8578 );
    nor g4176 ( n10685 , n3711 , n7573 );
    nor g4177 ( n11563 , n6203 , n2154 );
    not g4178 ( n12295 , n5065 );
    xnor g4179 ( n11264 , n4682 , n5985 );
    nor g4180 ( n3785 , n10441 , n1355 );
    or g4181 ( n3395 , n991 , n8030 );
    not g4182 ( n9891 , n10643 );
    not g4183 ( n7239 , n12319 );
    or g4184 ( n10154 , n8212 , n9380 );
    not g4185 ( n6231 , n3112 );
    or g4186 ( n6940 , n10938 , n1841 );
    not g4187 ( n4454 , n510 );
    and g4188 ( n12113 , n2952 , n7444 );
    not g4189 ( n7865 , n4862 );
    not g4190 ( n7986 , n4711 );
    not g4191 ( n4339 , n386 );
    xnor g4192 ( n11752 , n3011 , n4935 );
    or g4193 ( n12877 , n4802 , n8493 );
    nor g4194 ( n7368 , n5090 , n7638 );
    or g4195 ( n4212 , n5766 , n6080 );
    or g4196 ( n12804 , n11928 , n2059 );
    and g4197 ( n3701 , n8285 , n10933 );
    and g4198 ( n7129 , n12736 , n1286 );
    xor g4199 ( n4630 , n6707 , n3760 );
    or g4200 ( n8236 , n4561 , n8607 );
    xnor g4201 ( n3479 , n7830 , n3875 );
    xnor g4202 ( n8222 , n12333 , n9194 );
    xnor g4203 ( n386 , n7464 , n4933 );
    xnor g4204 ( n6048 , n8134 , n2537 );
    nor g4205 ( n1492 , n5428 , n11421 );
    xnor g4206 ( n1235 , n12913 , n10675 );
    not g4207 ( n7372 , n10657 );
    xnor g4208 ( n3845 , n10184 , n3391 );
    or g4209 ( n6711 , n1345 , n8632 );
    xnor g4210 ( n12474 , n10328 , n9715 );
    not g4211 ( n3564 , n4748 );
    or g4212 ( n101 , n2951 , n8651 );
    or g4213 ( n3623 , n10761 , n7530 );
    not g4214 ( n11609 , n10408 );
    or g4215 ( n6152 , n7001 , n8520 );
    or g4216 ( n11163 , n2674 , n10482 );
    xnor g4217 ( n9341 , n2386 , n12193 );
    and g4218 ( n12915 , n10908 , n5962 );
    not g4219 ( n11611 , n885 );
    and g4220 ( n10410 , n1722 , n4393 );
    not g4221 ( n3149 , n11324 );
    and g4222 ( n9137 , n2771 , n9093 );
    xnor g4223 ( n10255 , n7910 , n13092 );
    and g4224 ( n9089 , n6861 , n5465 );
    xnor g4225 ( n11850 , n1235 , n10494 );
    nor g4226 ( n9598 , n4489 , n6462 );
    or g4227 ( n3404 , n9867 , n10029 );
    or g4228 ( n1522 , n12367 , n3673 );
    not g4229 ( n12458 , n4331 );
    nor g4230 ( n1642 , n8354 , n6319 );
    or g4231 ( n5005 , n5713 , n9195 );
    and g4232 ( n299 , n3392 , n7979 );
    xnor g4233 ( n12685 , n1150 , n6005 );
    or g4234 ( n9573 , n7266 , n7060 );
    xnor g4235 ( n1181 , n11852 , n2876 );
    and g4236 ( n9624 , n2229 , n2207 );
    and g4237 ( n2010 , n10015 , n6608 );
    or g4238 ( n12181 , n2641 , n12657 );
    and g4239 ( n12822 , n8993 , n8250 );
    or g4240 ( n6045 , n1521 , n10272 );
    xnor g4241 ( n11578 , n1449 , n6702 );
    and g4242 ( n4688 , n7226 , n6912 );
    and g4243 ( n13157 , n2404 , n10325 );
    xnor g4244 ( n2799 , n1506 , n2883 );
    or g4245 ( n4679 , n1434 , n12657 );
    or g4246 ( n9211 , n808 , n1720 );
    or g4247 ( n9513 , n12490 , n8563 );
    xnor g4248 ( n3066 , n1212 , n4546 );
    and g4249 ( n2703 , n5050 , n5820 );
    xnor g4250 ( n9376 , n1460 , n6050 );
    xnor g4251 ( n9333 , n11610 , n12543 );
    or g4252 ( n4218 , n3753 , n6819 );
    or g4253 ( n9637 , n3854 , n4936 );
    not g4254 ( n327 , n9578 );
    and g4255 ( n9099 , n9620 , n3815 );
    and g4256 ( n5543 , n2378 , n8346 );
    and g4257 ( n4551 , n30 , n1419 );
    and g4258 ( n7937 , n9367 , n1357 );
    xnor g4259 ( n555 , n1312 , n12939 );
    xnor g4260 ( n8831 , n10613 , n10357 );
    nor g4261 ( n6882 , n3264 , n1762 );
    or g4262 ( n10467 , n4393 , n1722 );
    not g4263 ( n4783 , n9125 );
    and g4264 ( n2085 , n10560 , n1724 );
    not g4265 ( n4385 , n5758 );
    not g4266 ( n3972 , n8506 );
    xnor g4267 ( n11737 , n9613 , n12534 );
    and g4268 ( n3525 , n7416 , n6722 );
    and g4269 ( n5484 , n11566 , n453 );
    xnor g4270 ( n4155 , n3766 , n12890 );
    and g4271 ( n4117 , n10916 , n11402 );
    xnor g4272 ( n10088 , n8911 , n7357 );
    xnor g4273 ( n3188 , n17 , n9327 );
    or g4274 ( n1028 , n392 , n177 );
    xnor g4275 ( n8385 , n939 , n1971 );
    xnor g4276 ( n1891 , n11786 , n2070 );
    or g4277 ( n10388 , n6247 , n11753 );
    xnor g4278 ( n8629 , n585 , n12835 );
    not g4279 ( n6215 , n5189 );
    xnor g4280 ( n9912 , n3917 , n7631 );
    and g4281 ( n12033 , n9563 , n12216 );
    xnor g4282 ( n12158 , n10365 , n10556 );
    or g4283 ( n3529 , n3204 , n4729 );
    nor g4284 ( n5241 , n10284 , n6959 );
    xnor g4285 ( n11551 , n1267 , n9779 );
    xnor g4286 ( n9100 , n5747 , n3006 );
    nor g4287 ( n11527 , n2231 , n9295 );
    not g4288 ( n11369 , n1472 );
    xnor g4289 ( n711 , n6647 , n6908 );
    nor g4290 ( n3518 , n1496 , n5844 );
    xnor g4291 ( n982 , n2898 , n4688 );
    and g4292 ( n7266 , n7905 , n359 );
    nor g4293 ( n2686 , n10567 , n2131 );
    not g4294 ( n12368 , n5352 );
    not g4295 ( n10439 , n3832 );
    xnor g4296 ( n2313 , n4336 , n12222 );
    not g4297 ( n7560 , n5197 );
    not g4298 ( n2263 , n6496 );
    nor g4299 ( n2069 , n12053 , n8910 );
    or g4300 ( n12922 , n7543 , n931 );
    or g4301 ( n12555 , n6880 , n5072 );
    nor g4302 ( n1471 , n7650 , n3657 );
    or g4303 ( n11195 , n1820 , n12273 );
    not g4304 ( n1251 , n1956 );
    nor g4305 ( n1513 , n1757 , n10416 );
    xnor g4306 ( n2642 , n7488 , n4738 );
    and g4307 ( n9664 , n11053 , n4790 );
    or g4308 ( n7541 , n6769 , n10179 );
    and g4309 ( n6243 , n7300 , n11156 );
    or g4310 ( n12861 , n3598 , n9195 );
    xnor g4311 ( n2218 , n10257 , n2879 );
    and g4312 ( n3084 , n10637 , n9234 );
    xnor g4313 ( n4864 , n481 , n923 );
    not g4314 ( n11347 , n6107 );
    xnor g4315 ( n11479 , n9123 , n380 );
    or g4316 ( n1886 , n123 , n5069 );
    xnor g4317 ( n11671 , n9826 , n6090 );
    xnor g4318 ( n11478 , n12931 , n8641 );
    xnor g4319 ( n2147 , n10882 , n12906 );
    xnor g4320 ( n2879 , n6121 , n8282 );
    nor g4321 ( n732 , n9597 , n9372 );
    and g4322 ( n4295 , n2922 , n281 );
    nor g4323 ( n9816 , n2523 , n6237 );
    and g4324 ( n10759 , n6996 , n6614 );
    or g4325 ( n13081 , n1406 , n5797 );
    not g4326 ( n11810 , n8506 );
    or g4327 ( n7046 , n4391 , n6102 );
    xnor g4328 ( n135 , n5903 , n11955 );
    not g4329 ( n3998 , n8345 );
    or g4330 ( n8694 , n11370 , n7221 );
    xnor g4331 ( n2529 , n11953 , n6048 );
    buf g4332 ( n1985 , n3058 );
    not g4333 ( n318 , n9187 );
    or g4334 ( n147 , n1587 , n11668 );
    or g4335 ( n7204 , n1629 , n13020 );
    xnor g4336 ( n2033 , n5844 , n1496 );
    and g4337 ( n2576 , n8582 , n4298 );
    xnor g4338 ( n12933 , n9142 , n7740 );
    xnor g4339 ( n1093 , n5342 , n2609 );
    and g4340 ( n9097 , n2781 , n8440 );
    xnor g4341 ( n10875 , n3767 , n11257 );
    xnor g4342 ( n729 , n4397 , n3457 );
    not g4343 ( n12786 , n3769 );
    or g4344 ( n2788 , n3528 , n10918 );
    and g4345 ( n11346 , n4189 , n1799 );
    or g4346 ( n280 , n3460 , n10016 );
    or g4347 ( n2808 , n8330 , n5073 );
    not g4348 ( n9972 , n2037 );
    xnor g4349 ( n10777 , n6357 , n12602 );
    not g4350 ( n7163 , n10013 );
    and g4351 ( n7494 , n12028 , n120 );
    not g4352 ( n2048 , n6937 );
    or g4353 ( n2292 , n11245 , n9737 );
    and g4354 ( n5170 , n8228 , n13058 );
    and g4355 ( n10598 , n2993 , n10480 );
    or g4356 ( n11543 , n7864 , n3939 );
    xnor g4357 ( n43 , n8571 , n925 );
    xnor g4358 ( n5790 , n1234 , n1934 );
    not g4359 ( n7025 , n1143 );
    or g4360 ( n117 , n1609 , n11911 );
    xnor g4361 ( n893 , n5007 , n6977 );
    or g4362 ( n9724 , n10432 , n10403 );
    and g4363 ( n850 , n10829 , n6071 );
    nor g4364 ( n1355 , n4962 , n10810 );
    not g4365 ( n9461 , n9277 );
    and g4366 ( n8607 , n1314 , n8177 );
    not g4367 ( n13194 , n4862 );
    xnor g4368 ( n3824 , n3706 , n1407 );
    or g4369 ( n2863 , n11610 , n1456 );
    or g4370 ( n12413 , n3404 , n10984 );
    and g4371 ( n1156 , n1196 , n2345 );
    or g4372 ( n7023 , n12000 , n8912 );
    or g4373 ( n6995 , n8623 , n10581 );
    or g4374 ( n1772 , n9016 , n1026 );
    nor g4375 ( n10694 , n4926 , n5710 );
    xnor g4376 ( n748 , n12745 , n4092 );
    or g4377 ( n5439 , n6810 , n12501 );
    xnor g4378 ( n6609 , n2477 , n1801 );
    xnor g4379 ( n916 , n2240 , n1023 );
    nor g4380 ( n398 , n11217 , n9601 );
    or g4381 ( n6403 , n12220 , n2100 );
    and g4382 ( n12821 , n2215 , n10052 );
    and g4383 ( n9685 , n8959 , n7106 );
    not g4384 ( n1347 , n1085 );
    xnor g4385 ( n5056 , n7634 , n9442 );
    or g4386 ( n165 , n5874 , n9122 );
    and g4387 ( n1717 , n1548 , n4176 );
    not g4388 ( n11960 , n9906 );
    xnor g4389 ( n11726 , n6509 , n9590 );
    xnor g4390 ( n7141 , n6155 , n179 );
    or g4391 ( n10026 , n785 , n8268 );
    xnor g4392 ( n6147 , n3682 , n4259 );
    or g4393 ( n6187 , n7028 , n2092 );
    xnor g4394 ( n1295 , n12531 , n2241 );
    or g4395 ( n3095 , n6231 , n1043 );
    or g4396 ( n5696 , n3835 , n10521 );
    xnor g4397 ( n1444 , n4711 , n8540 );
    not g4398 ( n4949 , n11030 );
    xnor g4399 ( n5175 , n10869 , n8359 );
    xnor g4400 ( n9284 , n2334 , n2316 );
    and g4401 ( n10656 , n2432 , n11637 );
    not g4402 ( n11941 , n510 );
    xnor g4403 ( n2047 , n10090 , n3086 );
    and g4404 ( n3217 , n6483 , n9448 );
    xnor g4405 ( n10000 , n608 , n3451 );
    or g4406 ( n6558 , n8082 , n12388 );
    xnor g4407 ( n10337 , n12139 , n3306 );
    and g4408 ( n3390 , n9803 , n6946 );
    and g4409 ( n9603 , n6422 , n11260 );
    xnor g4410 ( n4428 , n366 , n301 );
    not g4411 ( n6814 , n8183 );
    not g4412 ( n9867 , n7659 );
    xnor g4413 ( n7590 , n11327 , n394 );
    buf g4414 ( n542 , n3185 );
    or g4415 ( n11575 , n12434 , n2544 );
    nor g4416 ( n9850 , n12341 , n7487 );
    or g4417 ( n1319 , n11808 , n3999 );
    not g4418 ( n2228 , n9915 );
    xnor g4419 ( n2586 , n820 , n4295 );
    or g4420 ( n953 , n2748 , n7353 );
    xnor g4421 ( n12226 , n4117 , n8321 );
    xnor g4422 ( n5555 , n12194 , n7727 );
    xnor g4423 ( n11469 , n4650 , n13102 );
    and g4424 ( n3794 , n6945 , n5108 );
    or g4425 ( n10338 , n3714 , n8552 );
    or g4426 ( n3614 , n6448 , n11806 );
    and g4427 ( n10374 , n11150 , n2034 );
    not g4428 ( n12871 , n10805 );
    or g4429 ( n5616 , n1945 , n1927 );
    or g4430 ( n5013 , n2701 , n8038 );
    or g4431 ( n1102 , n771 , n478 );
    and g4432 ( n2949 , n11823 , n4499 );
    or g4433 ( n2431 , n3534 , n121 );
    not g4434 ( n13083 , n9307 );
    or g4435 ( n9176 , n4540 , n10029 );
    xnor g4436 ( n1620 , n4570 , n3600 );
    and g4437 ( n12627 , n64 , n878 );
    not g4438 ( n8505 , n11030 );
    nor g4439 ( n1033 , n8550 , n13119 );
    and g4440 ( n3131 , n10024 , n9481 );
    or g4441 ( n5103 , n2661 , n2575 );
    xnor g4442 ( n6700 , n2753 , n10846 );
    xnor g4443 ( n2061 , n1637 , n1844 );
    nor g4444 ( n9939 , n969 , n7762 );
    xnor g4445 ( n5637 , n4886 , n7810 );
    xnor g4446 ( n9307 , n7445 , n9876 );
    or g4447 ( n11600 , n4248 , n3513 );
    and g4448 ( n5347 , n9123 , n8240 );
    and g4449 ( n1890 , n5625 , n9539 );
    or g4450 ( n162 , n6954 , n1556 );
    and g4451 ( n532 , n5874 , n9122 );
    xnor g4452 ( n7860 , n1610 , n6678 );
    xnor g4453 ( n1027 , n2802 , n11817 );
    or g4454 ( n12004 , n8204 , n8128 );
    and g4455 ( n4036 , n3130 , n1724 );
    and g4456 ( n5604 , n12113 , n8008 );
    xnor g4457 ( n6435 , n6113 , n11235 );
    or g4458 ( n5517 , n8935 , n12858 );
    and g4459 ( n11403 , n8298 , n1821 );
    nor g4460 ( n8213 , n4118 , n8321 );
    or g4461 ( n1244 , n616 , n6117 );
    or g4462 ( n2807 , n6519 , n8534 );
    xnor g4463 ( n10747 , n7856 , n9873 );
    nor g4464 ( n2231 , n5181 , n11272 );
    or g4465 ( n1230 , n10314 , n1043 );
    xnor g4466 ( n9123 , n2384 , n2873 );
    not g4467 ( n8322 , n1252 );
    or g4468 ( n3731 , n13182 , n5939 );
    not g4469 ( n7765 , n9905 );
    or g4470 ( n6346 , n3594 , n4632 );
    or g4471 ( n12851 , n10756 , n10871 );
    not g4472 ( n9417 , n4803 );
    and g4473 ( n2038 , n317 , n1557 );
    nor g4474 ( n5958 , n11039 , n521 );
    or g4475 ( n2762 , n3634 , n8268 );
    and g4476 ( n11292 , n1894 , n6191 );
    xnor g4477 ( n6386 , n12122 , n11788 );
    or g4478 ( n6894 , n7255 , n5315 );
    not g4479 ( n1189 , n7706 );
    xnor g4480 ( n11547 , n4740 , n11952 );
    xnor g4481 ( n4645 , n11050 , n5046 );
    not g4482 ( n6260 , n7259 );
    or g4483 ( n12346 , n13019 , n507 );
    or g4484 ( n8454 , n472 , n1271 );
    and g4485 ( n11761 , n8836 , n8766 );
    or g4486 ( n10340 , n8488 , n8642 );
    xnor g4487 ( n5422 , n1768 , n6626 );
    and g4488 ( n3400 , n9461 , n6269 );
    not g4489 ( n4643 , n11158 );
    not g4490 ( n2123 , n6273 );
    and g4491 ( n6592 , n12999 , n4923 );
    xnor g4492 ( n49 , n7039 , n2105 );
    xnor g4493 ( n10707 , n1085 , n10860 );
    or g4494 ( n11702 , n10281 , n1026 );
    xnor g4495 ( n6549 , n8373 , n5519 );
    and g4496 ( n11321 , n56 , n4392 );
    and g4497 ( n12117 , n11926 , n8657 );
    or g4498 ( n3215 , n12019 , n6660 );
    xnor g4499 ( n8714 , n1239 , n4747 );
    not g4500 ( n1815 , n4039 );
    or g4501 ( n12057 , n8043 , n7270 );
    and g4502 ( n9202 , n12348 , n6937 );
    xnor g4503 ( n3685 , n2530 , n9545 );
    nor g4504 ( n3561 , n5052 , n11325 );
    not g4505 ( n4524 , n9483 );
    and g4506 ( n6888 , n9538 , n7942 );
    and g4507 ( n12684 , n3467 , n5577 );
    xnor g4508 ( n3135 , n6222 , n6931 );
    nor g4509 ( n12200 , n1478 , n6547 );
    or g4510 ( n453 , n4252 , n9554 );
    xnor g4511 ( n6262 , n1611 , n8894 );
    not g4512 ( n11491 , n3967 );
    xnor g4513 ( n13175 , n10993 , n8159 );
    xnor g4514 ( n7757 , n10703 , n1566 );
    and g4515 ( n5363 , n8550 , n13119 );
    xnor g4516 ( n8000 , n2473 , n910 );
    and g4517 ( n5174 , n11360 , n11330 );
    or g4518 ( n1903 , n5645 , n7935 );
    not g4519 ( n9722 , n3895 );
    or g4520 ( n1267 , n4762 , n4375 );
    or g4521 ( n2203 , n6506 , n8360 );
    not g4522 ( n2809 , n2540 );
    not g4523 ( n10570 , n3562 );
    nor g4524 ( n5203 , n10424 , n13076 );
    xnor g4525 ( n12216 , n7832 , n9230 );
    not g4526 ( n8293 , n11366 );
    or g4527 ( n8455 , n9606 , n2544 );
    not g4528 ( n9674 , n12468 );
    xor g4529 ( n582 , n7500 , n567 );
    xnor g4530 ( n2745 , n5987 , n6447 );
    not g4531 ( n6481 , n7830 );
    and g4532 ( n1270 , n3244 , n8457 );
    and g4533 ( n6921 , n9353 , n3815 );
    xnor g4534 ( n6432 , n8237 , n3638 );
    or g4535 ( n7149 , n3443 , n6795 );
    xnor g4536 ( n1716 , n5737 , n9262 );
    not g4537 ( n7146 , n12651 );
    xnor g4538 ( n5985 , n5062 , n6957 );
    xnor g4539 ( n12497 , n3554 , n4108 );
    xnor g4540 ( n10453 , n7452 , n4151 );
    or g4541 ( n7433 , n7311 , n6251 );
    xnor g4542 ( n4429 , n440 , n6827 );
    not g4543 ( n9080 , n10451 );
    or g4544 ( n7538 , n2764 , n7504 );
    and g4545 ( n3691 , n3720 , n4079 );
    xnor g4546 ( n8503 , n12970 , n995 );
    or g4547 ( n133 , n6777 , n10205 );
    xnor g4548 ( n10197 , n4928 , n3064 );
    and g4549 ( n8875 , n1912 , n11634 );
    and g4550 ( n7324 , n4236 , n11989 );
    buf g4551 ( n11107 , n917 );
    nor g4552 ( n7014 , n12704 , n10267 );
    nor g4553 ( n11302 , n10438 , n12849 );
    or g4554 ( n8051 , n7329 , n12350 );
    xor g4555 ( n777 , n3910 , n9666 );
    not g4556 ( n10108 , n3310 );
    and g4557 ( n7389 , n4903 , n9015 );
    xnor g4558 ( n10095 , n12317 , n9902 );
    and g4559 ( n9455 , n9087 , n2453 );
    or g4560 ( n10762 , n6988 , n7430 );
    not g4561 ( n526 , n3862 );
    xnor g4562 ( n2645 , n11520 , n7370 );
    nor g4563 ( n4552 , n7494 , n2815 );
    or g4564 ( n828 , n4198 , n7221 );
    nor g4565 ( n6505 , n6884 , n6424 );
    xnor g4566 ( n11367 , n5125 , n12077 );
    xnor g4567 ( n3521 , n3351 , n1956 );
    and g4568 ( n8291 , n3006 , n7411 );
    and g4569 ( n4395 , n73 , n2634 );
    or g4570 ( n377 , n5168 , n9159 );
    nor g4571 ( n9110 , n6737 , n4245 );
    not g4572 ( n905 , n2771 );
    and g4573 ( n10116 , n8866 , n8620 );
    not g4574 ( n4786 , n4020 );
    not g4575 ( n3281 , n469 );
    nor g4576 ( n8304 , n4728 , n10414 );
    or g4577 ( n7475 , n6349 , n2408 );
    xor g4578 ( n9545 , n12473 , n11149 );
    xnor g4579 ( n576 , n8059 , n10722 );
    or g4580 ( n4038 , n4144 , n8030 );
    not g4581 ( n11356 , n1650 );
    not g4582 ( n2692 , n7729 );
    and g4583 ( n8845 , n1648 , n8952 );
    not g4584 ( n2095 , n12605 );
    or g4585 ( n99 , n9793 , n1144 );
    xnor g4586 ( n9121 , n1072 , n10473 );
    or g4587 ( n4850 , n4830 , n12089 );
    xor g4588 ( n9945 , n938 , n7006 );
    and g4589 ( n9507 , n5164 , n7412 );
    or g4590 ( n5249 , n4523 , n10528 );
    buf g4591 ( n1043 , n3858 );
    and g4592 ( n566 , n9479 , n8883 );
    xnor g4593 ( n1310 , n12466 , n10742 );
    or g4594 ( n9470 , n11018 , n10213 );
    and g4595 ( n1829 , n6687 , n432 );
    not g4596 ( n4342 , n11901 );
    or g4597 ( n12939 , n2449 , n1026 );
    or g4598 ( n5088 , n10755 , n12831 );
    xnor g4599 ( n9412 , n1285 , n857 );
    xnor g4600 ( n9167 , n5858 , n7206 );
    not g4601 ( n1301 , n2592 );
    and g4602 ( n11426 , n3907 , n10413 );
    not g4603 ( n4653 , n13160 );
    or g4604 ( n10336 , n12663 , n10535 );
    xnor g4605 ( n3034 , n2120 , n3808 );
    not g4606 ( n4846 , n8314 );
    not g4607 ( n1634 , n5167 );
    xnor g4608 ( n5908 , n3891 , n2833 );
    xnor g4609 ( n9175 , n6603 , n10079 );
    xnor g4610 ( n7448 , n9441 , n8368 );
    and g4611 ( n4880 , n7002 , n9240 );
    or g4612 ( n7899 , n5025 , n3893 );
    or g4613 ( n13162 , n7878 , n2893 );
    or g4614 ( n13218 , n4232 , n6692 );
    xnor g4615 ( n859 , n3978 , n8270 );
    or g4616 ( n10960 , n9487 , n4870 );
    xnor g4617 ( n10859 , n9318 , n10970 );
    and g4618 ( n5355 , n3167 , n2995 );
    not g4619 ( n8033 , n10789 );
    xnor g4620 ( n8441 , n7439 , n10963 );
    or g4621 ( n8622 , n8863 , n10573 );
    not g4622 ( n8617 , n9708 );
    not g4623 ( n6774 , n1418 );
    or g4624 ( n10783 , n9643 , n2775 );
    xnor g4625 ( n4886 , n4991 , n12980 );
    xnor g4626 ( n11507 , n3151 , n11033 );
    xnor g4627 ( n13187 , n6389 , n2869 );
    and g4628 ( n68 , n10460 , n5589 );
    not g4629 ( n1651 , n9300 );
    and g4630 ( n5724 , n6346 , n1745 );
    and g4631 ( n4345 , n3315 , n5760 );
    not g4632 ( n4564 , n4862 );
    or g4633 ( n4267 , n4156 , n10907 );
    or g4634 ( n6292 , n10481 , n4514 );
    not g4635 ( n6463 , n6058 );
    not g4636 ( n10158 , n3145 );
    nor g4637 ( n9944 , n1656 , n5376 );
    and g4638 ( n226 , n1569 , n7883 );
    xnor g4639 ( n5640 , n4800 , n9103 );
    not g4640 ( n12107 , n6456 );
    not g4641 ( n3826 , n11891 );
    and g4642 ( n4745 , n6890 , n6584 );
    nor g4643 ( n6933 , n6864 , n4977 );
    nor g4644 ( n450 , n4210 , n6150 );
    xnor g4645 ( n2787 , n1019 , n12245 );
    or g4646 ( n1533 , n1041 , n3824 );
    xnor g4647 ( n11594 , n9918 , n11339 );
    and g4648 ( n4095 , n4927 , n11100 );
    not g4649 ( n6810 , n6149 );
    or g4650 ( n10812 , n6223 , n10029 );
    and g4651 ( n5674 , n9994 , n7811 );
    nor g4652 ( n6972 , n8627 , n11334 );
    and g4653 ( n1109 , n7486 , n6159 );
    or g4654 ( n12411 , n8562 , n10106 );
    or g4655 ( n3166 , n12759 , n356 );
    or g4656 ( n3486 , n8625 , n9970 );
    and g4657 ( n9472 , n6323 , n10510 );
    and g4658 ( n4854 , n4089 , n9059 );
    xnor g4659 ( n4284 , n9096 , n1110 );
    xnor g4660 ( n3921 , n4630 , n4380 );
    xnor g4661 ( n540 , n10019 , n3472 );
    xnor g4662 ( n9250 , n11621 , n9175 );
    or g4663 ( n9673 , n5806 , n2276 );
    nor g4664 ( n4593 , n6701 , n7844 );
    xnor g4665 ( n1179 , n9612 , n12677 );
    xnor g4666 ( n10662 , n8888 , n9707 );
    xnor g4667 ( n10264 , n8023 , n12363 );
    not g4668 ( n6369 , n6550 );
    nor g4669 ( n247 , n4384 , n2210 );
    and g4670 ( n9636 , n932 , n4494 );
    xnor g4671 ( n571 , n4709 , n7781 );
    xnor g4672 ( n3052 , n8087 , n3403 );
    xnor g4673 ( n4015 , n11010 , n9046 );
    or g4674 ( n3859 , n12861 , n9661 );
    or g4675 ( n2194 , n517 , n1229 );
    xnor g4676 ( n9082 , n695 , n6411 );
    not g4677 ( n8922 , n10067 );
    nor g4678 ( n11765 , n6599 , n1108 );
    or g4679 ( n13 , n4077 , n8348 );
    not g4680 ( n1356 , n2658 );
    not g4681 ( n8790 , n4353 );
    and g4682 ( n4661 , n12995 , n8433 );
    or g4683 ( n2284 , n11113 , n4947 );
    xnor g4684 ( n8638 , n12329 , n12 );
    not g4685 ( n7642 , n9093 );
    xnor g4686 ( n11042 , n3479 , n11084 );
    xnor g4687 ( n1556 , n7329 , n12350 );
    or g4688 ( n10488 , n11333 , n3676 );
    or g4689 ( n8850 , n2718 , n6769 );
    nor g4690 ( n402 , n4196 , n2004 );
    or g4691 ( n5496 , n6658 , n4373 );
    xnor g4692 ( n2483 , n12409 , n743 );
    xnor g4693 ( n706 , n3360 , n2234 );
    xnor g4694 ( n12638 , n11571 , n12271 );
    and g4695 ( n4325 , n1216 , n8452 );
    xnor g4696 ( n6514 , n1177 , n9449 );
    not g4697 ( n6416 , n4862 );
    xnor g4698 ( n5856 , n5194 , n5623 );
    not g4699 ( n12469 , n9591 );
    not g4700 ( n5313 , n1465 );
    not g4701 ( n5930 , n9729 );
    or g4702 ( n12626 , n9493 , n9114 );
    nor g4703 ( n9971 , n6820 , n2915 );
    or g4704 ( n458 , n3906 , n10250 );
    not g4705 ( n666 , n2750 );
    and g4706 ( n2589 , n5719 , n6057 );
    and g4707 ( n5196 , n9102 , n10368 );
    and g4708 ( n2721 , n8723 , n2151 );
    or g4709 ( n9869 , n6387 , n7071 );
    xnor g4710 ( n9435 , n12178 , n5295 );
    nor g4711 ( n2197 , n11971 , n9068 );
    or g4712 ( n2540 , n542 , n206 );
    or g4713 ( n9977 , n1419 , n30 );
    and g4714 ( n12387 , n4937 , n978 );
    nor g4715 ( n11678 , n12081 , n12116 );
    not g4716 ( n11519 , n12284 );
    or g4717 ( n9488 , n10792 , n5087 );
    or g4718 ( n2982 , n3864 , n7218 );
    nor g4719 ( n4375 , n7992 , n6554 );
    xnor g4720 ( n4318 , n2188 , n6955 );
    xnor g4721 ( n6782 , n4827 , n916 );
    or g4722 ( n5257 , n10081 , n7282 );
    xnor g4723 ( n2526 , n3860 , n7352 );
    xnor g4724 ( n4501 , n7018 , n3328 );
    and g4725 ( n8220 , n2088 , n5851 );
    and g4726 ( n6839 , n2945 , n8559 );
    not g4727 ( n10910 , n3824 );
    and g4728 ( n5575 , n2559 , n4921 );
    or g4729 ( n2499 , n1842 , n6697 );
    and g4730 ( n1169 , n12868 , n2755 );
    or g4731 ( n1315 , n12924 , n492 );
    not g4732 ( n11858 , n5750 );
    xnor g4733 ( n1793 , n6558 , n9782 );
    xnor g4734 ( n5319 , n12184 , n2588 );
    nor g4735 ( n2524 , n9358 , n4645 );
    and g4736 ( n5885 , n5351 , n12659 );
    and g4737 ( n11505 , n4861 , n5447 );
    or g4738 ( n10625 , n10877 , n8702 );
    and g4739 ( n6787 , n4834 , n12580 );
    or g4740 ( n7375 , n4385 , n6769 );
    xnor g4741 ( n1071 , n4479 , n10582 );
    xnor g4742 ( n2954 , n1031 , n1412 );
    xnor g4743 ( n8988 , n8398 , n1190 );
    nor g4744 ( n9845 , n11220 , n10953 );
    xnor g4745 ( n5934 , n351 , n4833 );
    or g4746 ( n1680 , n1199 , n8030 );
    xnor g4747 ( n11758 , n3263 , n12045 );
    or g4748 ( n5933 , n9181 , n4237 );
    and g4749 ( n9207 , n3814 , n12504 );
    xnor g4750 ( n11809 , n7383 , n5068 );
    and g4751 ( n10376 , n10908 , n469 );
    buf g4752 ( n8030 , n5654 );
    or g4753 ( n7809 , n11340 , n4601 );
    xnor g4754 ( n1470 , n12947 , n43 );
    xnor g4755 ( n13199 , n2950 , n3143 );
    not g4756 ( n2800 , n11068 );
    or g4757 ( n4403 , n11291 , n12328 );
    or g4758 ( n12105 , n7406 , n11860 );
    xnor g4759 ( n1552 , n7892 , n9818 );
    xnor g4760 ( n7270 , n13061 , n3066 );
    not g4761 ( n6783 , n9822 );
    and g4762 ( n10294 , n6330 , n3387 );
    nor g4763 ( n4674 , n7096 , n8340 );
    and g4764 ( n5861 , n1756 , n4773 );
    not g4765 ( n10448 , n12289 );
    not g4766 ( n5485 , n7540 );
    or g4767 ( n11155 , n3616 , n12328 );
    xnor g4768 ( n9973 , n5606 , n13129 );
    or g4769 ( n8722 , n12677 , n9612 );
    not g4770 ( n3235 , n6302 );
    xor g4771 ( n8518 , n12112 , n11513 );
    or g4772 ( n1059 , n11905 , n3782 );
    or g4773 ( n10091 , n542 , n4936 );
    nor g4774 ( n11820 , n11632 , n4683 );
    xor g4775 ( n7217 , n1038 , n8191 );
    or g4776 ( n12599 , n7742 , n12188 );
    or g4777 ( n11460 , n4722 , n9075 );
    not g4778 ( n8194 , n6167 );
    xnor g4779 ( n12229 , n11221 , n1382 );
    xnor g4780 ( n13211 , n11691 , n11072 );
    nor g4781 ( n13152 , n8298 , n1821 );
    xnor g4782 ( n1284 , n8049 , n5214 );
    xnor g4783 ( n8624 , n6027 , n4214 );
    or g4784 ( n5165 , n6084 , n8061 );
    not g4785 ( n114 , n10606 );
    xnor g4786 ( n10951 , n3765 , n10734 );
    xnor g4787 ( n11693 , n12715 , n3465 );
    xnor g4788 ( n10177 , n3319 , n3789 );
    and g4789 ( n8229 , n11913 , n3642 );
    or g4790 ( n8180 , n6375 , n11144 );
    xnor g4791 ( n1534 , n2894 , n806 );
    or g4792 ( n239 , n2752 , n7010 );
    or g4793 ( n2710 , n11779 , n9195 );
    not g4794 ( n12281 , n424 );
    xnor g4795 ( n11252 , n3355 , n12364 );
    and g4796 ( n10310 , n1446 , n11652 );
    nor g4797 ( n2508 , n7940 , n2152 );
    and g4798 ( n5202 , n4827 , n2240 );
    not g4799 ( n2605 , n5237 );
    not g4800 ( n4610 , n7659 );
    and g4801 ( n2297 , n10418 , n3094 );
    nor g4802 ( n9859 , n6012 , n8797 );
    and g4803 ( n7747 , n2771 , n9531 );
    and g4804 ( n7832 , n1390 , n12612 );
    and g4805 ( n112 , n5976 , n1372 );
    xnor g4806 ( n4746 , n6495 , n2374 );
    or g4807 ( n6066 , n9658 , n11809 );
    or g4808 ( n9362 , n1605 , n6944 );
    or g4809 ( n11373 , n12728 , n11209 );
    or g4810 ( n2160 , n13036 , n5076 );
    or g4811 ( n6203 , n2135 , n12881 );
    nor g4812 ( n1500 , n11907 , n12327 );
    or g4813 ( n5331 , n10021 , n7837 );
    and g4814 ( n4226 , n11476 , n7398 );
    and g4815 ( n9634 , n3487 , n4313 );
    xnor g4816 ( n1812 , n9946 , n12731 );
    xnor g4817 ( n2991 , n1063 , n5147 );
    xnor g4818 ( n7057 , n6259 , n3461 );
    or g4819 ( n6530 , n12159 , n650 );
    xnor g4820 ( n1929 , n6024 , n9038 );
    nor g4821 ( n3874 , n13009 , n7105 );
    not g4822 ( n10950 , n9570 );
    not g4823 ( n622 , n11618 );
    nor g4824 ( n6534 , n3469 , n11958 );
    not g4825 ( n4960 , n411 );
    not g4826 ( n5478 , n12306 );
    not g4827 ( n10285 , n2629 );
    and g4828 ( n7495 , n8587 , n9776 );
    xnor g4829 ( n2190 , n3709 , n11769 );
    or g4830 ( n7523 , n3225 , n8702 );
    xnor g4831 ( n1318 , n6107 , n444 );
    or g4832 ( n4857 , n2332 , n4936 );
    and g4833 ( n4384 , n4557 , n4703 );
    not g4834 ( n7130 , n12935 );
    not g4835 ( n4780 , n1902 );
    xnor g4836 ( n11073 , n414 , n945 );
    and g4837 ( n1288 , n12799 , n5361 );
    xnor g4838 ( n10224 , n276 , n10454 );
    or g4839 ( n1453 , n7752 , n10360 );
    or g4840 ( n4776 , n12993 , n11274 );
    not g4841 ( n8757 , n9300 );
    nor g4842 ( n2606 , n12603 , n1910 );
    nor g4843 ( n12811 , n645 , n3600 );
    nor g4844 ( n11198 , n13153 , n4674 );
    or g4845 ( n7176 , n10135 , n8030 );
    xnor g4846 ( n6991 , n10842 , n10347 );
    xnor g4847 ( n1407 , n2822 , n9658 );
    xnor g4848 ( n7285 , n8091 , n10382 );
    xnor g4849 ( n697 , n6766 , n4292 );
    or g4850 ( n5664 , n12153 , n7825 );
    not g4851 ( n1589 , n8290 );
    and g4852 ( n5581 , n10516 , n4171 );
    xor g4853 ( n1611 , n2591 , n11202 );
    and g4854 ( n1446 , n4964 , n8506 );
    and g4855 ( n9108 , n2547 , n7471 );
    or g4856 ( n317 , n8469 , n961 );
    and g4857 ( n4563 , n2681 , n9344 );
    not g4858 ( n1549 , n4946 );
    buf g4859 ( n6893 , n13214 );
    not g4860 ( n8666 , n12282 );
    or g4861 ( n12637 , n1536 , n6265 );
    or g4862 ( n5953 , n8761 , n5769 );
    and g4863 ( n102 , n12037 , n10467 );
    and g4864 ( n8037 , n6452 , n7190 );
    and g4865 ( n11028 , n8597 , n1578 );
    or g4866 ( n4740 , n10193 , n5631 );
    not g4867 ( n11713 , n641 );
    xnor g4868 ( n313 , n600 , n11224 );
    xnor g4869 ( n10679 , n2113 , n9024 );
    not g4870 ( n2889 , n6085 );
    nor g4871 ( n11601 , n2019 , n7696 );
    or g4872 ( n5204 , n1099 , n9120 );
    xnor g4873 ( n229 , n5208 , n180 );
    or g4874 ( n695 , n2723 , n12786 );
    xnor g4875 ( n1884 , n5284 , n818 );
    or g4876 ( n6235 , n10128 , n12501 );
    and g4877 ( n6003 , n10070 , n10053 );
    and g4878 ( n664 , n3211 , n7814 );
    buf g4879 ( n4230 , n482 );
    and g4880 ( n9864 , n8764 , n10880 );
    and g4881 ( n4486 , n1697 , n12932 );
    xnor g4882 ( n1685 , n11636 , n5220 );
    not g4883 ( n1674 , n11296 );
    or g4884 ( n7101 , n11757 , n6265 );
    nor g4885 ( n5903 , n2171 , n10665 );
    not g4886 ( n8055 , n9136 );
    or g4887 ( n3996 , n2283 , n3762 );
    and g4888 ( n10633 , n7715 , n7411 );
    or g4889 ( n11888 , n2660 , n6317 );
    xnor g4890 ( n382 , n1294 , n11480 );
    or g4891 ( n10939 , n7133 , n12695 );
    or g4892 ( n1548 , n10184 , n3391 );
    or g4893 ( n11999 , n8594 , n12804 );
    not g4894 ( n8837 , n10185 );
    xnor g4895 ( n12839 , n9514 , n9688 );
    or g4896 ( n4236 , n6143 , n326 );
    or g4897 ( n3773 , n12354 , n11414 );
    xor g4898 ( n6532 , n9909 , n3108 );
    or g4899 ( n5057 , n437 , n87 );
    xnor g4900 ( n7330 , n2823 , n11962 );
    xnor g4901 ( n10306 , n5288 , n2274 );
    xnor g4902 ( n9503 , n3532 , n10935 );
    xnor g4903 ( n676 , n527 , n3992 );
    and g4904 ( n3374 , n11050 , n457 );
    buf g4905 ( n2951 , n10497 );
    or g4906 ( n7322 , n195 , n8198 );
    and g4907 ( n600 , n6325 , n2006 );
    xnor g4908 ( n10069 , n11439 , n9667 );
    buf g4909 ( n10106 , n8640 );
    or g4910 ( n5625 , n5328 , n10871 );
    and g4911 ( n7090 , n10870 , n3937 );
    or g4912 ( n2971 , n4732 , n7221 );
    xnor g4913 ( n4496 , n2613 , n2172 );
    not g4914 ( n6001 , n6085 );
    xnor g4915 ( n4982 , n4130 , n1201 );
    or g4916 ( n5299 , n2884 , n10016 );
    nor g4917 ( n8605 , n9563 , n12216 );
    xnor g4918 ( n7183 , n12361 , n4526 );
    not g4919 ( n3727 , n3061 );
    xnor g4920 ( n8872 , n2505 , n6340 );
    xnor g4921 ( n12968 , n3488 , n7965 );
    and g4922 ( n11679 , n9392 , n8464 );
    nor g4923 ( n29 , n5878 , n708 );
    not g4924 ( n9899 , n10577 );
    or g4925 ( n1029 , n2551 , n5501 );
    and g4926 ( n13203 , n11972 , n11583 );
    not g4927 ( n8646 , n22 );
    nor g4928 ( n4622 , n3088 , n6184 );
    or g4929 ( n11990 , n3634 , n8348 );
    xnor g4930 ( n11337 , n2066 , n12007 );
    nor g4931 ( n1635 , n9607 , n1837 );
    not g4932 ( n1218 , n10408 );
    or g4933 ( n613 , n11657 , n7579 );
    not g4934 ( n13141 , n3330 );
    xnor g4935 ( n8810 , n2897 , n4379 );
    or g4936 ( n11580 , n2974 , n5240 );
    or g4937 ( n3341 , n8760 , n540 );
    or g4938 ( n959 , n9010 , n4947 );
    not g4939 ( n7549 , n5266 );
    xnor g4940 ( n12338 , n5572 , n9762 );
    not g4941 ( n1436 , n12289 );
    or g4942 ( n1677 , n13079 , n6474 );
    xnor g4943 ( n7341 , n1378 , n9021 );
    and g4944 ( n1942 , n6184 , n3088 );
    or g4945 ( n375 , n4709 , n526 );
    xnor g4946 ( n12527 , n1389 , n11942 );
    or g4947 ( n4782 , n11371 , n11292 );
    or g4948 ( n1784 , n7932 , n12998 );
    or g4949 ( n3175 , n11167 , n3485 );
    xnor g4950 ( n4528 , n6036 , n1641 );
    not g4951 ( n12036 , n6522 );
    nor g4952 ( n6497 , n473 , n1662 );
    and g4953 ( n12007 , n11803 , n7886 );
    not g4954 ( n9632 , n9591 );
    xor g4955 ( n3187 , n4523 , n11031 );
    or g4956 ( n7652 , n8848 , n8227 );
    not g4957 ( n5939 , n8230 );
    xnor g4958 ( n567 , n2246 , n3234 );
    or g4959 ( n8471 , n3866 , n11668 );
    or g4960 ( n2573 , n4224 , n9864 );
    not g4961 ( n1246 , n5180 );
    or g4962 ( n9144 , n10059 , n12388 );
    nor g4963 ( n1928 , n12828 , n10732 );
    or g4964 ( n3725 , n1135 , n12164 );
    not g4965 ( n4527 , n7341 );
    not g4966 ( n12083 , n13214 );
    nor g4967 ( n4222 , n6555 , n8437 );
    not g4968 ( n7783 , n2882 );
    not g4969 ( n7076 , n411 );
    and g4970 ( n10937 , n5681 , n5445 );
    or g4971 ( n536 , n11810 , n12273 );
    or g4972 ( n1387 , n6587 , n10179 );
    xnor g4973 ( n6828 , n1136 , n7956 );
    not g4974 ( n11341 , n6790 );
    nor g4975 ( n4309 , n6356 , n6989 );
    not g4976 ( n10098 , n11441 );
    xnor g4977 ( n2417 , n1793 , n8178 );
    xnor g4978 ( n12583 , n3203 , n7054 );
    xnor g4979 ( n4989 , n5808 , n13209 );
    and g4980 ( n12195 , n2866 , n12825 );
    and g4981 ( n2716 , n10541 , n4260 );
    nor g4982 ( n12688 , n6943 , n3637 );
    and g4983 ( n10517 , n9946 , n9004 );
    or g4984 ( n1020 , n147 , n10094 );
    xnor g4985 ( n12751 , n7567 , n6097 );
    xnor g4986 ( n3631 , n3298 , n1140 );
    or g4987 ( n10237 , n1501 , n3971 );
    xnor g4988 ( n5762 , n10389 , n1964 );
    xnor g4989 ( n6092 , n11192 , n9199 );
    not g4990 ( n4370 , n12408 );
    nor g4991 ( n9462 , n12299 , n324 );
    xnor g4992 ( n1172 , n8581 , n10330 );
    or g4993 ( n4298 , n4143 , n12501 );
    or g4994 ( n5256 , n7622 , n8815 );
    xnor g4995 ( n10602 , n5290 , n5214 );
    or g4996 ( n8733 , n12262 , n3227 );
    not g4997 ( n1887 , n1307 );
    or g4998 ( n4785 , n493 , n5169 );
    and g4999 ( n725 , n6649 , n9770 );
    xnor g5000 ( n6487 , n4046 , n4603 );
    nor g5001 ( n8478 , n5850 , n638 );
    and g5002 ( n5154 , n5151 , n7843 );
    not g5003 ( n2861 , n2498 );
    xnor g5004 ( n12958 , n1777 , n4029 );
    xnor g5005 ( n10107 , n11314 , n1037 );
    or g5006 ( n10865 , n445 , n3949 );
    not g5007 ( n2165 , n5678 );
    nor g5008 ( n4340 , n8241 , n4807 );
    or g5009 ( n10201 , n3110 , n1462 );
    or g5010 ( n11318 , n6099 , n8268 );
    not g5011 ( n6173 , n10606 );
    or g5012 ( n12343 , n2965 , n12561 );
    xnor g5013 ( n5891 , n10839 , n3559 );
    and g5014 ( n7735 , n5142 , n4945 );
    nor g5015 ( n7005 , n1414 , n8960 );
    and g5016 ( n7260 , n3893 , n5025 );
    and g5017 ( n6734 , n5568 , n3006 );
    or g5018 ( n12080 , n10500 , n11063 );
    and g5019 ( n11840 , n5568 , n4470 );
    xnor g5020 ( n10048 , n9994 , n9963 );
    xnor g5021 ( n7956 , n6870 , n9144 );
    xnor g5022 ( n1851 , n12661 , n1196 );
    or g5023 ( n9801 , n8648 , n6436 );
    not g5024 ( n5721 , n2010 );
    not g5025 ( n980 , n4377 );
    and g5026 ( n5235 , n2960 , n3240 );
    and g5027 ( n981 , n9054 , n11825 );
    xnor g5028 ( n7267 , n9957 , n11036 );
    and g5029 ( n10808 , n1364 , n9915 );
    or g5030 ( n4790 , n6682 , n7324 );
    or g5031 ( n8998 , n5460 , n6306 );
    xnor g5032 ( n2904 , n2668 , n5429 );
    not g5033 ( n8166 , n9611 );
    or g5034 ( n10972 , n11345 , n5250 );
    and g5035 ( n11741 , n9216 , n5962 );
    not g5036 ( n9464 , n2279 );
    or g5037 ( n1693 , n4185 , n13181 );
    or g5038 ( n11646 , n12151 , n1814 );
    xnor g5039 ( n4900 , n2536 , n4821 );
    xnor g5040 ( n7168 , n7286 , n12377 );
    not g5041 ( n10715 , n4877 );
    or g5042 ( n1931 , n1159 , n6429 );
    or g5043 ( n2908 , n8720 , n11300 );
    xnor g5044 ( n5230 , n770 , n7115 );
    nor g5045 ( n10907 , n8273 , n12986 );
    or g5046 ( n57 , n12042 , n1836 );
    xnor g5047 ( n680 , n11739 , n4324 );
    xor g5048 ( n7965 , n5835 , n11492 );
    not g5049 ( n8438 , n6669 );
    or g5050 ( n6858 , n686 , n11679 );
    and g5051 ( n11862 , n2771 , n12289 );
    nor g5052 ( n6072 , n6744 , n347 );
    or g5053 ( n6962 , n12882 , n4373 );
    xnor g5054 ( n11103 , n1626 , n11694 );
    or g5055 ( n5820 , n9835 , n1378 );
    or g5056 ( n6074 , n9061 , n8364 );
    nor g5057 ( n2064 , n6510 , n5160 );
    or g5058 ( n3743 , n4102 , n5002 );
    and g5059 ( n1598 , n8139 , n9475 );
    xnor g5060 ( n1106 , n1545 , n10438 );
    xnor g5061 ( n6892 , n9494 , n11976 );
    not g5062 ( n7436 , n11565 );
    and g5063 ( n12711 , n10775 , n9956 );
    not g5064 ( n10068 , n1242 );
    and g5065 ( n4463 , n2712 , n5640 );
    or g5066 ( n2912 , n2669 , n8268 );
    or g5067 ( n1365 , n899 , n12501 );
    nor g5068 ( n2360 , n5958 , n5426 );
    or g5069 ( n9642 , n3537 , n12388 );
    or g5070 ( n5981 , n3892 , n6404 );
    not g5071 ( n8199 , n8571 );
    or g5072 ( n3339 , n5749 , n2133 );
    or g5073 ( n1799 , n4659 , n3151 );
    xnor g5074 ( n7083 , n7552 , n13020 );
    and g5075 ( n1116 , n6160 , n10010 );
    and g5076 ( n10963 , n208 , n9716 );
    and g5077 ( n11441 , n5077 , n12702 );
    and g5078 ( n4084 , n7772 , n12289 );
    not g5079 ( n9581 , n9591 );
    not g5080 ( n13116 , n11971 );
    and g5081 ( n12866 , n4799 , n9074 );
    and g5082 ( n10461 , n8973 , n2132 );
    xnor g5083 ( n4512 , n7932 , n6677 );
    and g5084 ( n11857 , n3191 , n3423 );
    not g5085 ( n3373 , n2464 );
    not g5086 ( n6448 , n5421 );
    or g5087 ( n4710 , n7890 , n2919 );
    or g5088 ( n9721 , n7379 , n9116 );
    or g5089 ( n5338 , n820 , n4832 );
    or g5090 ( n8380 , n4686 , n4796 );
    or g5091 ( n3660 , n3784 , n3981 );
    and g5092 ( n6898 , n2655 , n12479 );
    and g5093 ( n13106 , n117 , n1749 );
    or g5094 ( n12266 , n5875 , n12721 );
    or g5095 ( n11139 , n8903 , n5432 );
    xnor g5096 ( n7201 , n4184 , n11855 );
    not g5097 ( n5999 , n11061 );
    not g5098 ( n6967 , n5969 );
    or g5099 ( n12462 , n11864 , n12328 );
    or g5100 ( n10438 , n4258 , n12501 );
    and g5101 ( n4904 , n5070 , n5438 );
    not g5102 ( n7430 , n10408 );
    and g5103 ( n4652 , n10610 , n12525 );
    not g5104 ( n0 , n7720 );
    or g5105 ( n1906 , n12913 , n11351 );
    xnor g5106 ( n8242 , n7821 , n4767 );
    and g5107 ( n5924 , n5291 , n3288 );
    or g5108 ( n2291 , n11605 , n7288 );
    nor g5109 ( n11093 , n2314 , n1042 );
    not g5110 ( n9709 , n11236 );
    xor g5111 ( n1722 , n5352 , n7044 );
    xnor g5112 ( n11181 , n856 , n2560 );
    not g5113 ( n3895 , n11974 );
    and g5114 ( n5566 , n12354 , n11414 );
    xnor g5115 ( n9046 , n9146 , n11802 );
    xor g5116 ( n1927 , n5709 , n10343 );
    and g5117 ( n12298 , n8334 , n11717 );
    or g5118 ( n8957 , n5226 , n177 );
    xnor g5119 ( n10405 , n10655 , n224 );
    or g5120 ( n3517 , n4462 , n6265 );
    not g5121 ( n8160 , n12592 );
    not g5122 ( n6332 , n2882 );
    xnor g5123 ( n1913 , n11273 , n3957 );
    or g5124 ( n1574 , n3683 , n9832 );
    or g5125 ( n10965 , n3826 , n4194 );
    and g5126 ( n2032 , n179 , n9740 );
    nor g5127 ( n4768 , n4545 , n1834 );
    not g5128 ( n10924 , n11546 );
    xnor g5129 ( n7059 , n7604 , n531 );
    xor g5130 ( n744 , n7059 , n8997 );
    xnor g5131 ( n4071 , n12599 , n10350 );
    not g5132 ( n7133 , n2666 );
    or g5133 ( n9770 , n4874 , n9419 );
    or g5134 ( n5916 , n9765 , n7491 );
    or g5135 ( n9066 , n7872 , n9075 );
    or g5136 ( n6998 , n8556 , n1144 );
    xnor g5137 ( n8411 , n12405 , n4951 );
    not g5138 ( n12052 , n8860 );
    and g5139 ( n2192 , n12677 , n9612 );
    not g5140 ( n10014 , n3100 );
    or g5141 ( n6341 , n11075 , n13210 );
    or g5142 ( n7325 , n3430 , n7557 );
    xnor g5143 ( n9037 , n10980 , n3181 );
    xnor g5144 ( n847 , n4145 , n12150 );
    or g5145 ( n7702 , n1571 , n5841 );
    not g5146 ( n8500 , n7065 );
    xnor g5147 ( n8705 , n6334 , n9719 );
    and g5148 ( n12551 , n8407 , n12321 );
    and g5149 ( n6132 , n3160 , n10435 );
    xnor g5150 ( n753 , n11138 , n10801 );
    not g5151 ( n6751 , n9531 );
    xnor g5152 ( n5260 , n4265 , n2715 );
    or g5153 ( n12630 , n4290 , n9195 );
    nor g5154 ( n10550 , n3384 , n4670 );
    xnor g5155 ( n9544 , n6904 , n1875 );
    xnor g5156 ( n1398 , n12669 , n8230 );
    xnor g5157 ( n11984 , n10518 , n7943 );
    not g5158 ( n5569 , n3112 );
    or g5159 ( n1761 , n3243 , n8702 );
    or g5160 ( n4654 , n2452 , n12501 );
    xnor g5161 ( n12021 , n6327 , n10499 );
    xnor g5162 ( n4211 , n11666 , n2626 );
    or g5163 ( n7645 , n9632 , n11354 );
    and g5164 ( n10659 , n8073 , n5247 );
    xnor g5165 ( n1083 , n9713 , n12136 );
    or g5166 ( n7582 , n9455 , n8253 );
    xnor g5167 ( n10153 , n2661 , n8195 );
    nor g5168 ( n6993 , n5114 , n10306 );
    and g5169 ( n10860 , n245 , n9099 );
    xnor g5170 ( n3575 , n7516 , n10779 );
    not g5171 ( n5841 , n1364 );
    nor g5172 ( n12755 , n7822 , n9603 );
    and g5173 ( n10841 , n614 , n133 );
    or g5174 ( n10719 , n6344 , n2234 );
    or g5175 ( n8159 , n3217 , n10246 );
    or g5176 ( n7456 , n8264 , n10834 );
    xnor g5177 ( n5552 , n12639 , n7698 );
    xnor g5178 ( n11899 , n10638 , n606 );
    not g5179 ( n7833 , n3091 );
    xnor g5180 ( n537 , n8319 , n711 );
    xnor g5181 ( n3757 , n11276 , n4801 );
    and g5182 ( n1655 , n9020 , n5771 );
    or g5183 ( n10870 , n11021 , n6999 );
    or g5184 ( n7623 , n11519 , n9282 );
    xnor g5185 ( n3209 , n5397 , n10933 );
    and g5186 ( n5059 , n2373 , n782 );
    xnor g5187 ( n12634 , n2143 , n8527 );
    xnor g5188 ( n2869 , n4338 , n5618 );
    xnor g5189 ( n7116 , n10825 , n2052 );
    and g5190 ( n7884 , n11397 , n12558 );
    not g5191 ( n13005 , n2068 );
    not g5192 ( n6924 , n4002 );
    or g5193 ( n8237 , n10926 , n6564 );
    or g5194 ( n10327 , n6220 , n4144 );
    or g5195 ( n8978 , n3491 , n4672 );
    and g5196 ( n7640 , n1817 , n5904 );
    xnor g5197 ( n8382 , n10269 , n5570 );
    or g5198 ( n6807 , n2219 , n7052 );
    xnor g5199 ( n8219 , n7572 , n6450 );
    or g5200 ( n5703 , n10713 , n2994 );
    not g5201 ( n9323 , n5709 );
    or g5202 ( n6588 , n6562 , n2201 );
    xnor g5203 ( n6077 , n12332 , n4771 );
    and g5204 ( n8707 , n51 , n671 );
    xor g5205 ( n872 , n621 , n9836 );
    not g5206 ( n6367 , n1724 );
    and g5207 ( n9998 , n11821 , n8132 );
    xnor g5208 ( n5813 , n9186 , n4081 );
    nor g5209 ( n553 , n10034 , n5089 );
    not g5210 ( n3766 , n6660 );
    not g5211 ( n9345 , n6174 );
    and g5212 ( n12982 , n12074 , n1873 );
    not g5213 ( n8254 , n9669 );
    not g5214 ( n4604 , n10225 );
    not g5215 ( n11973 , n8967 );
    or g5216 ( n6745 , n12321 , n8407 );
    not g5217 ( n5733 , n5065 );
    not g5218 ( n12164 , n854 );
    not g5219 ( n11008 , n3134 );
    or g5220 ( n3359 , n5316 , n9290 );
    xnor g5221 ( n12835 , n6441 , n6671 );
    or g5222 ( n3780 , n3962 , n8490 );
    or g5223 ( n11312 , n9739 , n11101 );
    or g5224 ( n8784 , n7690 , n199 );
    and g5225 ( n7829 , n8166 , n5434 );
    or g5226 ( n2378 , n6463 , n2976 );
    and g5227 ( n10588 , n5816 , n136 );
    or g5228 ( n1855 , n1111 , n4207 );
    and g5229 ( n6190 , n9166 , n4284 );
    xnor g5230 ( n11138 , n6088 , n5610 );
    xnor g5231 ( n10312 , n6801 , n4476 );
    nor g5232 ( n3322 , n1527 , n6961 );
    and g5233 ( n2628 , n2778 , n12433 );
    nor g5234 ( n10280 , n9296 , n11838 );
    or g5235 ( n6687 , n8658 , n6891 );
    and g5236 ( n7619 , n8998 , n12132 );
    and g5237 ( n4026 , n1623 , n5001 );
    and g5238 ( n7472 , n12106 , n7929 );
    and g5239 ( n6128 , n199 , n7690 );
    nor g5240 ( n1702 , n12936 , n12538 );
    xnor g5241 ( n7248 , n3152 , n6017 );
    xnor g5242 ( n10811 , n7220 , n12373 );
    or g5243 ( n13006 , n11320 , n5076 );
    xnor g5244 ( n4310 , n9656 , n1948 );
    not g5245 ( n4055 , n5332 );
    nor g5246 ( n9171 , n1611 , n8834 );
    not g5247 ( n10573 , n11030 );
    xnor g5248 ( n9678 , n1227 , n4647 );
    not g5249 ( n4723 , n4064 );
    not g5250 ( n5812 , n2977 );
    xnor g5251 ( n10643 , n3398 , n9480 );
    not g5252 ( n3047 , n510 );
    not g5253 ( n1101 , n2758 );
    and g5254 ( n8189 , n1597 , n10618 );
    or g5255 ( n3577 , n5070 , n5438 );
    or g5256 ( n6744 , n10974 , n8268 );
    xnor g5257 ( n8451 , n3140 , n5398 );
    not g5258 ( n275 , n10963 );
    xnor g5259 ( n11934 , n12580 , n4669 );
    not g5260 ( n12114 , n92 );
    xnor g5261 ( n12973 , n8890 , n5955 );
    and g5262 ( n12919 , n7297 , n303 );
    or g5263 ( n7143 , n8329 , n12847 );
    xnor g5264 ( n11767 , n1873 , n3497 );
    not g5265 ( n7742 , n2252 );
    and g5266 ( n1025 , n1945 , n8601 );
    or g5267 ( n7064 , n9238 , n2059 );
    nor g5268 ( n12437 , n12815 , n2874 );
    xnor g5269 ( n12503 , n8218 , n3059 );
    and g5270 ( n9629 , n12680 , n6636 );
    or g5271 ( n839 , n8245 , n12039 );
    or g5272 ( n820 , n6381 , n10886 );
    and g5273 ( n11768 , n5863 , n5436 );
    or g5274 ( n4289 , n10177 , n8075 );
    nor g5275 ( n6054 , n5214 , n2771 );
    or g5276 ( n3350 , n3313 , n14 );
    and g5277 ( n2566 , n13177 , n3705 );
    and g5278 ( n5860 , n7839 , n3552 );
    or g5279 ( n6654 , n11352 , n2544 );
    and g5280 ( n6418 , n9974 , n9323 );
    and g5281 ( n1831 , n5462 , n11716 );
    and g5282 ( n2774 , n5970 , n1687 );
    nor g5283 ( n5627 , n8856 , n4340 );
    not g5284 ( n9942 , n7209 );
    xnor g5285 ( n6551 , n6018 , n280 );
    or g5286 ( n2153 , n359 , n7905 );
    and g5287 ( n11774 , n8466 , n11222 );
    nor g5288 ( n20 , n37 , n5224 );
    or g5289 ( n12807 , n9646 , n12984 );
    not g5290 ( n3885 , n8043 );
    nor g5291 ( n12607 , n2233 , n1421 );
    xnor g5292 ( n4307 , n2368 , n10107 );
    or g5293 ( n12090 , n121 , n11609 );
    not g5294 ( n138 , n1912 );
    not g5295 ( n11308 , n7517 );
    and g5296 ( n4651 , n3340 , n1953 );
    or g5297 ( n11063 , n12841 , n9075 );
    nor g5298 ( n8198 , n9336 , n4152 );
    and g5299 ( n4447 , n1251 , n3351 );
    and g5300 ( n1922 , n1039 , n10655 );
    xnor g5301 ( n6009 , n5726 , n1552 );
    not g5302 ( n10781 , n497 );
    xnor g5303 ( n3905 , n12901 , n8047 );
    xnor g5304 ( n1991 , n9443 , n4261 );
    and g5305 ( n10473 , n2999 , n10235 );
    xnor g5306 ( n2730 , n11805 , n1969 );
    xnor g5307 ( n9190 , n7 , n10231 );
    or g5308 ( n11640 , n4808 , n12847 );
    not g5309 ( n6244 , n4646 );
    not g5310 ( n9382 , n6034 );
    or g5311 ( n1578 , n6383 , n10179 );
    or g5312 ( n7750 , n4863 , n243 );
    xnor g5313 ( n11296 , n8557 , n3704 );
    xnor g5314 ( n8939 , n13156 , n11186 );
    xnor g5315 ( n4434 , n4408 , n5910 );
    xnor g5316 ( n2881 , n12760 , n5012 );
    or g5317 ( n8298 , n8681 , n4373 );
    not g5318 ( n6033 , n3815 );
    xnor g5319 ( n3317 , n4216 , n6668 );
    or g5320 ( n6417 , n10049 , n9223 );
    not g5321 ( n6528 , n11394 );
    not g5322 ( n1331 , n3409 );
    not g5323 ( n6040 , n3085 );
    xnor g5324 ( n2974 , n9317 , n2458 );
    or g5325 ( n7732 , n4352 , n9682 );
    or g5326 ( n10510 , n7731 , n4596 );
    xnor g5327 ( n7713 , n3512 , n6781 );
    or g5328 ( n7990 , n4046 , n11638 );
    nor g5329 ( n3902 , n6357 , n2325 );
    nor g5330 ( n6679 , n10832 , n13007 );
    xnor g5331 ( n5751 , n5847 , n2915 );
    and g5332 ( n5779 , n435 , n4776 );
    not g5333 ( n442 , n6453 );
    nor g5334 ( n8246 , n2640 , n1858 );
    not g5335 ( n1197 , n854 );
    or g5336 ( n10848 , n7908 , n5302 );
    and g5337 ( n10619 , n9649 , n2096 );
    and g5338 ( n5317 , n10157 , n400 );
    or g5339 ( n1588 , n6368 , n1154 );
    or g5340 ( n12517 , n2574 , n11228 );
    and g5341 ( n4407 , n11945 , n3773 );
    and g5342 ( n6544 , n12196 , n2269 );
    xnor g5343 ( n12461 , n10548 , n6281 );
    and g5344 ( n1934 , n11119 , n9900 );
    not g5345 ( n7868 , n4335 );
    or g5346 ( n5224 , n8006 , n12242 );
    and g5347 ( n5008 , n8379 , n5273 );
    not g5348 ( n3096 , n4419 );
    nor g5349 ( n9391 , n10308 , n12917 );
    xnor g5350 ( n3950 , n4439 , n10177 );
    xnor g5351 ( n3573 , n2924 , n771 );
    or g5352 ( n9648 , n11868 , n8030 );
    xnor g5353 ( n3292 , n1911 , n9862 );
    nor g5354 ( n3189 , n5833 , n3095 );
    xnor g5355 ( n13124 , n5648 , n7420 );
    xnor g5356 ( n7036 , n10895 , n4183 );
    or g5357 ( n8386 , n5990 , n7723 );
    or g5358 ( n6211 , n8176 , n2221 );
    or g5359 ( n1257 , n12533 , n283 );
    xnor g5360 ( n10125 , n6727 , n5083 );
    or g5361 ( n12681 , n2221 , n7723 );
    or g5362 ( n2492 , n3068 , n7530 );
    xnor g5363 ( n12363 , n8488 , n8642 );
    xor g5364 ( n9849 , n11376 , n10200 );
    or g5365 ( n3852 , n10686 , n1895 );
    xnor g5366 ( n3223 , n12588 , n9302 );
    nor g5367 ( n1279 , n574 , n9405 );
    or g5368 ( n2702 , n10936 , n10028 );
    not g5369 ( n3158 , n12482 );
    and g5370 ( n1925 , n8811 , n7284 );
    and g5371 ( n5743 , n2444 , n11461 );
    xnor g5372 ( n1708 , n3707 , n1371 );
    not g5373 ( n8470 , n5535 );
    and g5374 ( n9907 , n2046 , n12637 );
    xnor g5375 ( n11314 , n2801 , n7993 );
    and g5376 ( n7180 , n4616 , n8255 );
    not g5377 ( n9706 , n11076 );
    xnor g5378 ( n5755 , n12477 , n9404 );
    not g5379 ( n10290 , n1650 );
    or g5380 ( n3270 , n7062 , n7221 );
    xnor g5381 ( n9820 , n11120 , n12459 );
    not g5382 ( n7597 , n3815 );
    xnor g5383 ( n13129 , n4887 , n10523 );
    or g5384 ( n4821 , n3509 , n7723 );
    or g5385 ( n7690 , n5265 , n4640 );
    or g5386 ( n5412 , n8023 , n11569 );
    and g5387 ( n3649 , n6916 , n1664 );
    xnor g5388 ( n5580 , n3597 , n12050 );
    xnor g5389 ( n6406 , n9133 , n5113 );
    and g5390 ( n11438 , n4301 , n344 );
    nor g5391 ( n1872 , n8291 , n783 );
    and g5392 ( n11538 , n5367 , n8496 );
    and g5393 ( n11518 , n1308 , n4498 );
    xnor g5394 ( n6650 , n1501 , n6256 );
    or g5395 ( n9813 , n7284 , n8811 );
    and g5396 ( n8793 , n7176 , n8366 );
    xnor g5397 ( n5509 , n5637 , n8193 );
    xor g5398 ( n7214 , n2670 , n12665 );
    or g5399 ( n3151 , n1571 , n1570 );
    and g5400 ( n10398 , n10770 , n510 );
    nor g5401 ( n9064 , n2141 , n10841 );
    or g5402 ( n3807 , n9810 , n3805 );
    not g5403 ( n6383 , n12263 );
    or g5404 ( n12355 , n12093 , n12273 );
    not g5405 ( n6596 , n10522 );
    and g5406 ( n12675 , n1130 , n12088 );
    and g5407 ( n10774 , n2880 , n11154 );
    not g5408 ( n8210 , n12414 );
    not g5409 ( n5430 , n13058 );
    xnor g5410 ( n7799 , n11134 , n10687 );
    not g5411 ( n3128 , n4982 );
    or g5412 ( n3533 , n3407 , n177 );
    xnor g5413 ( n4424 , n395 , n9659 );
    or g5414 ( n2474 , n12441 , n9223 );
    nor g5415 ( n4913 , n9938 , n3146 );
    or g5416 ( n11336 , n3385 , n2005 );
    xnor g5417 ( n11952 , n8137 , n10954 );
    nor g5418 ( n7952 , n7160 , n4374 );
    or g5419 ( n8550 , n5688 , n5076 );
    xnor g5420 ( n2012 , n11117 , n3093 );
    nor g5421 ( n8489 , n7048 , n11265 );
    and g5422 ( n860 , n11069 , n4158 );
    buf g5423 ( n10499 , n7281 );
    and g5424 ( n597 , n11555 , n9728 );
    xnor g5425 ( n1788 , n8448 , n12496 );
    not g5426 ( n10726 , n5871 );
    not g5427 ( n2222 , n11030 );
    xnor g5428 ( n7177 , n4041 , n7392 );
    not g5429 ( n2557 , n9353 );
    xnor g5430 ( n5530 , n2460 , n10987 );
    xnor g5431 ( n10181 , n5980 , n4238 );
    or g5432 ( n8132 , n12172 , n10472 );
    and g5433 ( n9401 , n6906 , n6186 );
    xnor g5434 ( n3569 , n12582 , n1204 );
    or g5435 ( n12104 , n2790 , n4546 );
    xnor g5436 ( n12645 , n12276 , n1094 );
    not g5437 ( n10188 , n8468 );
    not g5438 ( n3092 , n3087 );
    or g5439 ( n877 , n6590 , n5076 );
    and g5440 ( n8712 , n4406 , n5165 );
    or g5441 ( n7211 , n6629 , n11107 );
    or g5442 ( n3263 , n2321 , n7998 );
    xnor g5443 ( n2543 , n6111 , n8211 );
    or g5444 ( n9471 , n9154 , n4640 );
    not g5445 ( n12906 , n11551 );
    or g5446 ( n10834 , n8849 , n6635 );
    or g5447 ( n5610 , n6367 , n11521 );
    nor g5448 ( n3356 , n2343 , n3861 );
    xnor g5449 ( n4794 , n4321 , n11749 );
    not g5450 ( n8989 , n5553 );
    and g5451 ( n491 , n410 , n8662 );
    and g5452 ( n1923 , n110 , n5946 );
    not g5453 ( n7707 , n6826 );
    and g5454 ( n12819 , n4114 , n2339 );
    or g5455 ( n169 , n5007 , n6977 );
    and g5456 ( n7352 , n623 , n2863 );
    or g5457 ( n5720 , n12563 , n4640 );
    not g5458 ( n5215 , n4146 );
    and g5459 ( n12404 , n8277 , n2337 );
    and g5460 ( n9506 , n6318 , n12057 );
    nor g5461 ( n7635 , n10053 , n10070 );
    xnor g5462 ( n3568 , n1560 , n1654 );
    and g5463 ( n8846 , n4114 , n1916 );
    or g5464 ( n6188 , n8380 , n11981 );
    or g5465 ( n5246 , n12697 , n7640 );
    nor g5466 ( n3205 , n13206 , n5473 );
    not g5467 ( n6100 , n1964 );
    not g5468 ( n1629 , n7552 );
    and g5469 ( n6237 , n10327 , n6711 );
    or g5470 ( n271 , n2352 , n4352 );
    or g5471 ( n10896 , n7917 , n2049 );
    or g5472 ( n8570 , n5939 , n9159 );
    and g5473 ( n4422 , n10710 , n7665 );
    xnor g5474 ( n10283 , n6373 , n3663 );
    xnor g5475 ( n7840 , n10139 , n1093 );
    or g5476 ( n3914 , n11277 , n71 );
    or g5477 ( n2189 , n6365 , n8560 );
    or g5478 ( n7632 , n5826 , n2831 );
    and g5479 ( n5240 , n10526 , n9892 );
    xnor g5480 ( n7067 , n675 , n12345 );
    nor g5481 ( n10905 , n5978 , n8126 );
    not g5482 ( n5087 , n3085 );
    xnor g5483 ( n6081 , n7010 , n9663 );
    not g5484 ( n12671 , n6937 );
    xnor g5485 ( n2275 , n8880 , n7789 );
    and g5486 ( n12542 , n8700 , n8382 );
    or g5487 ( n936 , n12330 , n2731 );
    not g5488 ( n4879 , n3121 );
    or g5489 ( n6837 , n5182 , n3981 );
    not g5490 ( n2902 , n679 );
    not g5491 ( n12095 , n12101 );
    or g5492 ( n3371 , n5752 , n2177 );
    xnor g5493 ( n3741 , n307 , n2033 );
    and g5494 ( n5089 , n4369 , n2951 );
    not g5495 ( n364 , n6730 );
    nor g5496 ( n11436 , n11248 , n8200 );
    not g5497 ( n11231 , n8788 );
    or g5498 ( n794 , n5683 , n3949 );
    and g5499 ( n2279 , n6236 , n11565 );
    xnor g5500 ( n2840 , n3348 , n1167 );
    and g5501 ( n3 , n8154 , n8975 );
    and g5502 ( n12642 , n1358 , n1766 );
    or g5503 ( n4760 , n4875 , n7935 );
    xnor g5504 ( n7145 , n5479 , n2648 );
    or g5505 ( n8896 , n6768 , n4442 );
    xnor g5506 ( n2423 , n7395 , n2131 );
    xnor g5507 ( n3258 , n7267 , n11413 );
    and g5508 ( n10549 , n5692 , n5834 );
    and g5509 ( n9422 , n8242 , n1491 );
    and g5510 ( n7220 , n7636 , n4562 );
    nor g5511 ( n1069 , n307 , n3422 );
    xnor g5512 ( n12251 , n7465 , n12357 );
    or g5513 ( n8164 , n2066 , n12007 );
    not g5514 ( n6672 , n772 );
    or g5515 ( n417 , n7394 , n5379 );
    nor g5516 ( n2063 , n1740 , n9881 );
    not g5517 ( n3121 , n4426 );
    xnor g5518 ( n9936 , n6302 , n9032 );
    not g5519 ( n5749 , n5536 );
    or g5520 ( n9672 , n9513 , n1400 );
    or g5521 ( n11688 , n13183 , n1570 );
    and g5522 ( n4616 , n4537 , n10408 );
    and g5523 ( n9510 , n6668 , n4470 );
    and g5524 ( n1421 , n13178 , n6576 );
    not g5525 ( n829 , n6818 );
    or g5526 ( n8571 , n3962 , n7935 );
    or g5527 ( n9519 , n4741 , n12328 );
    xnor g5528 ( n11627 , n7746 , n3856 );
    and g5529 ( n13135 , n3280 , n3844 );
    xnor g5530 ( n8555 , n143 , n7237 );
    not g5531 ( n12795 , n10805 );
    not g5532 ( n2211 , n6362 );
    and g5533 ( n8145 , n7568 , n6376 );
    and g5534 ( n9760 , n8187 , n3620 );
    xnor g5535 ( n3011 , n1960 , n8939 );
    and g5536 ( n7524 , n4664 , n2728 );
    xnor g5537 ( n4090 , n3250 , n12226 );
    not g5538 ( n1712 , n1752 );
    xnor g5539 ( n6857 , n7660 , n8709 );
    and g5540 ( n2685 , n8421 , n5150 );
    xnor g5541 ( n1988 , n7137 , n8096 );
    xnor g5542 ( n9776 , n7809 , n13232 );
    or g5543 ( n9966 , n3433 , n3649 );
    not g5544 ( n10692 , n472 );
    nor g5545 ( n9521 , n11448 , n3082 );
    xnor g5546 ( n1233 , n2600 , n5000 );
    or g5547 ( n12610 , n10792 , n2449 );
    or g5548 ( n1394 , n7223 , n9223 );
    not g5549 ( n9112 , n5065 );
    xnor g5550 ( n4767 , n5039 , n1678 );
    not g5551 ( n19 , n11151 );
    and g5552 ( n598 , n896 , n11620 );
    or g5553 ( n10807 , n12814 , n5242 );
    and g5554 ( n6952 , n2199 , n2385 );
    nor g5555 ( n6319 , n6972 , n12694 );
    not g5556 ( n2945 , n1623 );
    xnor g5557 ( n10126 , n9134 , n2035 );
    xnor g5558 ( n5042 , n7489 , n10836 );
    xnor g5559 ( n9925 , n220 , n2548 );
    xnor g5560 ( n10736 , n7885 , n1010 );
    xnor g5561 ( n201 , n8304 , n7347 );
    not g5562 ( n9917 , n4743 );
    xnor g5563 ( n5780 , n11318 , n2275 );
    xnor g5564 ( n10596 , n3590 , n9256 );
    or g5565 ( n898 , n12126 , n1144 );
    or g5566 ( n8526 , n11994 , n331 );
    nor g5567 ( n989 , n2521 , n6792 );
    not g5568 ( n12242 , n1364 );
    or g5569 ( n7333 , n6677 , n12714 );
    xnor g5570 ( n11458 , n4428 , n3446 );
    and g5571 ( n552 , n11500 , n710 );
    not g5572 ( n6986 , n4862 );
    not g5573 ( n98 , n11634 );
    not g5574 ( n11525 , n9540 );
    xnor g5575 ( n10378 , n6805 , n5386 );
    not g5576 ( n12049 , n834 );
    not g5577 ( n4877 , n12083 );
    xor g5578 ( n4285 , n10914 , n5960 );
    nor g5579 ( n4944 , n11546 , n7199 );
    nor g5580 ( n10788 , n7382 , n10461 );
    not g5581 ( n8679 , n1915 );
    and g5582 ( n412 , n10291 , n11439 );
    xor g5583 ( n6957 , n7069 , n5124 );
    or g5584 ( n10320 , n2452 , n11522 );
    nor g5585 ( n3421 , n348 , n4219 );
    xnor g5586 ( n7002 , n3090 , n13095 );
    not g5587 ( n5838 , n1935 );
    xnor g5588 ( n2422 , n1510 , n11298 );
    and g5589 ( n655 , n3736 , n929 );
    or g5590 ( n10233 , n7789 , n4492 );
    and g5591 ( n1103 , n12353 , n8316 );
    and g5592 ( n9791 , n8648 , n6436 );
    or g5593 ( n609 , n3067 , n10985 );
    or g5594 ( n4970 , n7242 , n12886 );
    xnor g5595 ( n12549 , n3030 , n9878 );
    or g5596 ( n10262 , n10112 , n5521 );
    or g5597 ( n7916 , n9675 , n1570 );
    xnor g5598 ( n10649 , n2784 , n1838 );
    xnor g5599 ( n8190 , n4244 , n6547 );
    and g5600 ( n5092 , n10277 , n3297 );
    xnor g5601 ( n6249 , n7732 , n6035 );
    xnor g5602 ( n7926 , n11447 , n12277 );
    not g5603 ( n8053 , n353 );
    not g5604 ( n10714 , n8468 );
    xor g5605 ( n6815 , n5502 , n11319 );
    or g5606 ( n5772 , n7260 , n523 );
    nor g5607 ( n8964 , n8654 , n8951 );
    not g5608 ( n7716 , n11016 );
    xnor g5609 ( n9633 , n6598 , n12439 );
    or g5610 ( n4547 , n565 , n8593 );
    or g5611 ( n2801 , n3364 , n6033 );
    not g5612 ( n8011 , n8135 );
    or g5613 ( n2270 , n3880 , n8953 );
    and g5614 ( n13074 , n13021 , n6232 );
    xnor g5615 ( n9410 , n10487 , n3904 );
    or g5616 ( n6626 , n8415 , n11959 );
    and g5617 ( n6049 , n399 , n2596 );
    xnor g5618 ( n643 , n12806 , n2589 );
    xnor g5619 ( n5961 , n7043 , n8136 );
    and g5620 ( n3926 , n2302 , n844 );
    not g5621 ( n13167 , n13217 );
    not g5622 ( n9308 , n2466 );
    or g5623 ( n2301 , n11683 , n3981 );
    or g5624 ( n4085 , n1659 , n10574 );
    nor g5625 ( n7385 , n12315 , n6495 );
    xnor g5626 ( n12481 , n4592 , n5889 );
    xnor g5627 ( n2896 , n11455 , n11839 );
    and g5628 ( n9178 , n3833 , n2946 );
    nor g5629 ( n1834 , n10020 , n12884 );
    not g5630 ( n7396 , n3769 );
    xnor g5631 ( n4968 , n7155 , n9825 );
    xnor g5632 ( n3881 , n9670 , n7902 );
    xnor g5633 ( n6357 , n12358 , n9412 );
    and g5634 ( n5593 , n3006 , n12289 );
    or g5635 ( n11539 , n2485 , n6032 );
    or g5636 ( n8060 , n7291 , n8030 );
    or g5637 ( n7444 , n9161 , n6372 );
    nor g5638 ( n11118 , n6569 , n7169 );
    xnor g5639 ( n10826 , n4298 , n8262 );
    or g5640 ( n4451 , n2825 , n12388 );
    xor g5641 ( n754 , n3606 , n12632 );
    xnor g5642 ( n232 , n10284 , n12513 );
    xor g5643 ( n11217 , n1731 , n4443 );
    not g5644 ( n1325 , n11061 );
    or g5645 ( n11461 , n10017 , n8490 );
    xnor g5646 ( n1037 , n4351 , n3482 );
    not g5647 ( n2858 , n11937 );
    xnor g5648 ( n5876 , n6765 , n2572 );
    nor g5649 ( n10259 , n5637 , n8193 );
    xnor g5650 ( n9534 , n8762 , n1397 );
    xnor g5651 ( n8299 , n11211 , n5422 );
    or g5652 ( n383 , n7074 , n9223 );
    nor g5653 ( n5919 , n11953 , n578 );
    and g5654 ( n3961 , n207 , n12290 );
    xnor g5655 ( n3535 , n12996 , n6514 );
    nor g5656 ( n7904 , n8643 , n7954 );
    nor g5657 ( n7218 , n2112 , n5614 );
    not g5658 ( n75 , n13060 );
    nor g5659 ( n7705 , n4397 , n8165 );
    and g5660 ( n12072 , n10500 , n11063 );
    or g5661 ( n1664 , n1578 , n8597 );
    nor g5662 ( n5239 , n12191 , n12700 );
    xnor g5663 ( n12523 , n8714 , n7677 );
    not g5664 ( n2254 , n8860 );
    nor g5665 ( n7786 , n5120 , n8474 );
    or g5666 ( n11455 , n10037 , n8534 );
    xnor g5667 ( n7428 , n4931 , n9577 );
    nor g5668 ( n6869 , n7362 , n12609 );
    xnor g5669 ( n460 , n4273 , n7985 );
    not g5670 ( n1261 , n2882 );
    xnor g5671 ( n12803 , n4275 , n76 );
    or g5672 ( n8202 , n3101 , n1789 );
    xnor g5673 ( n10047 , n9108 , n7036 );
    not g5674 ( n10856 , n4586 );
    or g5675 ( n9751 , n3911 , n4947 );
    or g5676 ( n3297 , n3517 , n3571 );
    xnor g5677 ( n10169 , n4314 , n5004 );
    and g5678 ( n6639 , n6275 , n9993 );
    xnor g5679 ( n10863 , n12137 , n3213 );
    not g5680 ( n4136 , n7307 );
    xnor g5681 ( n7725 , n10025 , n12079 );
    not g5682 ( n13238 , n10770 );
    not g5683 ( n6255 , n8218 );
    or g5684 ( n7122 , n5261 , n3981 );
    not g5685 ( n9430 , n5815 );
    and g5686 ( n12565 , n7435 , n12294 );
    xnor g5687 ( n4909 , n10864 , n1757 );
    or g5688 ( n9298 , n4352 , n4947 );
    or g5689 ( n12722 , n2150 , n3177 );
    not g5690 ( n5658 , n6791 );
    not g5691 ( n6175 , n6780 );
    and g5692 ( n12450 , n3469 , n11958 );
    or g5693 ( n7662 , n9920 , n8423 );
    or g5694 ( n12136 , n543 , n6982 );
    and g5695 ( n5415 , n8549 , n8919 );
    xnor g5696 ( n12123 , n6832 , n13124 );
    or g5697 ( n4599 , n2080 , n2463 );
    xnor g5698 ( n1122 , n8518 , n6081 );
    and g5699 ( n10102 , n7980 , n3846 );
    nor g5700 ( n3386 , n5403 , n11387 );
    or g5701 ( n5513 , n13089 , n6207 );
    xnor g5702 ( n3742 , n884 , n11251 );
    not g5703 ( n10234 , n10409 );
    and g5704 ( n6727 , n3830 , n4098 );
    or g5705 ( n6472 , n3018 , n6951 );
    not g5706 ( n3253 , n6222 );
    or g5707 ( n1202 , n7358 , n6769 );
    and g5708 ( n10936 , n87 , n437 );
    not g5709 ( n3755 , n6643 );
    or g5710 ( n7789 , n6028 , n7221 );
    xnor g5711 ( n7882 , n11501 , n8611 );
    or g5712 ( n8366 , n11466 , n4640 );
    and g5713 ( n12683 , n11511 , n9621 );
    xnor g5714 ( n12451 , n2333 , n11830 );
    or g5715 ( n12643 , n2382 , n3546 );
    not g5716 ( n2639 , n5189 );
    nor g5717 ( n11686 , n3931 , n5119 );
    and g5718 ( n11166 , n1735 , n10674 );
    not g5719 ( n1300 , n1075 );
    or g5720 ( n7391 , n5452 , n12681 );
    and g5721 ( n10818 , n34 , n701 );
    not g5722 ( n6733 , n5189 );
    not g5723 ( n6271 , n9591 );
    xnor g5724 ( n1456 , n6454 , n2895 );
    xnor g5725 ( n5127 , n4027 , n10952 );
    not g5726 ( n1047 , n3605 );
    and g5727 ( n7225 , n6433 , n6276 );
    not g5728 ( n1184 , n7387 );
    or g5729 ( n1040 , n8838 , n6078 );
    nor g5730 ( n1565 , n12801 , n9604 );
    xnor g5731 ( n113 , n5734 , n6886 );
    and g5732 ( n7255 , n1653 , n6479 );
    xnor g5733 ( n4182 , n8245 , n3632 );
    xnor g5734 ( n3228 , n11268 , n298 );
    xnor g5735 ( n2184 , n4599 , n9361 );
    or g5736 ( n4531 , n7188 , n8534 );
    and g5737 ( n9415 , n1105 , n3136 );
    not g5738 ( n4293 , n12391 );
    xnor g5739 ( n11358 , n10261 , n8820 );
    and g5740 ( n6675 , n6725 , n10862 );
    not g5741 ( n9767 , n9093 );
    or g5742 ( n9051 , n8200 , n2216 );
    or g5743 ( n3361 , n13077 , n3454 );
    xnor g5744 ( n2632 , n7731 , n4596 );
    or g5745 ( n5783 , n882 , n8655 );
    and g5746 ( n3335 , n11061 , n3769 );
    not g5747 ( n11344 , n3398 );
    nor g5748 ( n288 , n4941 , n12229 );
    xnor g5749 ( n736 , n274 , n7318 );
    and g5750 ( n4873 , n3060 , n7046 );
    or g5751 ( n1501 , n3047 , n11354 );
    or g5752 ( n12521 , n1933 , n9407 );
    not g5753 ( n1540 , n5897 );
    xnor g5754 ( n642 , n11904 , n6788 );
    or g5755 ( n2193 , n1725 , n6769 );
    xnor g5756 ( n6495 , n10036 , n3072 );
    not g5757 ( n4715 , n11837 );
    or g5758 ( n2786 , n6178 , n5048 );
    not g5759 ( n11099 , n8476 );
    or g5760 ( n2860 , n11618 , n4136 );
    or g5761 ( n4493 , n6336 , n8752 );
    or g5762 ( n4611 , n10287 , n12695 );
    and g5763 ( n974 , n1786 , n254 );
    buf g5764 ( n4373 , n12537 );
    or g5765 ( n10081 , n10229 , n6288 );
    xnor g5766 ( n9377 , n3227 , n12262 );
    and g5767 ( n4129 , n6168 , n5729 );
    or g5768 ( n8749 , n2768 , n8268 );
    or g5769 ( n6303 , n8301 , n6166 );
    xnor g5770 ( n7088 , n12294 , n5067 );
    not g5771 ( n9557 , n1724 );
    not g5772 ( n10037 , n8233 );
    or g5773 ( n10136 , n12841 , n121 );
    xnor g5774 ( n874 , n8703 , n4965 );
    or g5775 ( n7278 , n7775 , n11483 );
    and g5776 ( n6632 , n203 , n4218 );
    or g5777 ( n3595 , n1326 , n5476 );
    nor g5778 ( n1768 , n4555 , n2450 );
    and g5779 ( n11798 , n5533 , n5621 );
    or g5780 ( n2253 , n475 , n12942 );
    or g5781 ( n6492 , n6439 , n6306 );
    and g5782 ( n7479 , n12445 , n1681 );
    and g5783 ( n8824 , n3852 , n10363 );
    or g5784 ( n9454 , n3360 , n10511 );
    not g5785 ( n11522 , n8230 );
    nor g5786 ( n4992 , n8211 , n6111 );
    or g5787 ( n5342 , n5947 , n7723 );
    xnor g5788 ( n12509 , n6540 , n10603 );
    xnor g5789 ( n2765 , n5937 , n643 );
    nor g5790 ( n2429 , n5283 , n2554 );
    xnor g5791 ( n8303 , n13027 , n3653 );
    xnor g5792 ( n5444 , n9886 , n2218 );
    xnor g5793 ( n7165 , n6718 , n2847 );
    and g5794 ( n10083 , n4753 , n8570 );
    or g5795 ( n4811 , n2516 , n9155 );
    or g5796 ( n554 , n11142 , n3792 );
    xnor g5797 ( n223 , n9743 , n7946 );
    and g5798 ( n2367 , n6776 , n12708 );
    xnor g5799 ( n7387 , n592 , n4845 );
    and g5800 ( n4813 , n5909 , n12792 );
    and g5801 ( n11475 , n12300 , n10972 );
    or g5802 ( n11797 , n1256 , n6285 );
    and g5803 ( n2810 , n8485 , n12078 );
    and g5804 ( n9571 , n7333 , n1784 );
    and g5805 ( n8070 , n9215 , n10927 );
    nor g5806 ( n13222 , n2524 , n3691 );
    xnor g5807 ( n6896 , n9594 , n3621 );
    and g5808 ( n620 , n11580 , n9937 );
    xnor g5809 ( n843 , n11100 , n4927 );
    or g5810 ( n10123 , n12545 , n5924 );
    not g5811 ( n5827 , n8200 );
    not g5812 ( n10049 , n5962 );
    xnor g5813 ( n10773 , n5322 , n7172 );
    xor g5814 ( n8593 , n10172 , n9137 );
    or g5815 ( n7337 , n1389 , n3014 );
    and g5816 ( n9832 , n3851 , n12382 );
    xnor g5817 ( n8404 , n7402 , n2331 );
    nor g5818 ( n11523 , n10739 , n5824 );
    or g5819 ( n5318 , n7828 , n3888 );
    nor g5820 ( n7490 , n3855 , n1046 );
    nor g5821 ( n419 , n5678 , n8684 );
    and g5822 ( n9379 , n9656 , n10848 );
    or g5823 ( n4406 , n4663 , n1127 );
    or g5824 ( n9911 , n12732 , n10319 );
    nor g5825 ( n4550 , n664 , n5759 );
    not g5826 ( n4732 , n2737 );
    xnor g5827 ( n2819 , n7989 , n977 );
    not g5828 ( n917 , n3006 );
    xnor g5829 ( n5442 , n972 , n11071 );
    xnor g5830 ( n6014 , n345 , n8054 );
    not g5831 ( n10352 , n2758 );
    or g5832 ( n12318 , n920 , n9079 );
    xnor g5833 ( n5835 , n1645 , n6169 );
    xnor g5834 ( n13031 , n4832 , n2586 );
    nor g5835 ( n12447 , n6338 , n5739 );
    xnor g5836 ( n10869 , n2931 , n1980 );
    nor g5837 ( n4207 , n12735 , n11432 );
    xnor g5838 ( n4597 , n4793 , n11622 );
    xnor g5839 ( n5557 , n9920 , n9991 );
    xnor g5840 ( n7417 , n10824 , n8147 );
    nor g5841 ( n4287 , n288 , n2628 );
    and g5842 ( n3840 , n12222 , n4336 );
    not g5843 ( n5182 , n12965 );
    buf g5844 ( n2133 , n1301 );
    xnor g5845 ( n5259 , n5906 , n1100 );
    nor g5846 ( n1042 , n5731 , n11108 );
    or g5847 ( n635 , n6069 , n11067 );
    xnor g5848 ( n4972 , n13131 , n7108 );
    and g5849 ( n2714 , n9690 , n10741 );
    xnor g5850 ( n4911 , n11269 , n8196 );
    nor g5851 ( n5426 , n2935 , n31 );
    and g5852 ( n1849 , n12107 , n8907 );
    xnor g5853 ( n5161 , n6396 , n7425 );
    xnor g5854 ( n11607 , n9079 , n10934 );
    xnor g5855 ( n10247 , n11090 , n468 );
    xnor g5856 ( n4046 , n1747 , n11145 );
    and g5857 ( n1219 , n9115 , n6538 );
    xnor g5858 ( n10684 , n2785 , n1895 );
    and g5859 ( n12186 , n5707 , n1432 );
    not g5860 ( n2967 , n3954 );
    nor g5861 ( n5788 , n5216 , n3751 );
    and g5862 ( n78 , n951 , n3085 );
    xnor g5863 ( n4444 , n3740 , n9599 );
    not g5864 ( n9478 , n9747 );
    not g5865 ( n116 , n13221 );
    or g5866 ( n12844 , n8351 , n6532 );
    xnor g5867 ( n9143 , n11901 , n10809 );
    or g5868 ( n12271 , n8020 , n206 );
    xnor g5869 ( n10424 , n1098 , n9766 );
    or g5870 ( n3174 , n5040 , n11144 );
    or g5871 ( n1023 , n8472 , n3981 );
    or g5872 ( n3247 , n12837 , n1325 );
    or g5873 ( n5166 , n3770 , n3084 );
    or g5874 ( n8272 , n2135 , n894 );
    nor g5875 ( n2653 , n9994 , n7811 );
    xnor g5876 ( n4842 , n12971 , n3470 );
    or g5877 ( n12989 , n8176 , n11122 );
    or g5878 ( n6136 , n1077 , n3960 );
    or g5879 ( n5145 , n10031 , n4226 );
    or g5880 ( n4332 , n9228 , n3817 );
    or g5881 ( n8751 , n3105 , n6746 );
    or g5882 ( n9783 , n6685 , n1458 );
    and g5883 ( n11047 , n2299 , n12190 );
    xnor g5884 ( n762 , n12943 , n2839 );
    and g5885 ( n8414 , n3175 , n8731 );
    xnor g5886 ( n862 , n1951 , n12739 );
    not g5887 ( n2752 , n1055 );
    not g5888 ( n709 , n4036 );
    or g5889 ( n5506 , n12451 , n2402 );
    not g5890 ( n5294 , n1502 );
    or g5891 ( n9797 , n406 , n11950 );
    xnor g5892 ( n7788 , n10585 , n2696 );
    xnor g5893 ( n6410 , n1559 , n6919 );
    and g5894 ( n1825 , n6051 , n11998 );
    not g5895 ( n11637 , n3521 );
    and g5896 ( n10677 , n12056 , n2975 );
    or g5897 ( n8512 , n10085 , n7530 );
    xnor g5898 ( n12970 , n471 , n9472 );
    nor g5899 ( n2110 , n10064 , n760 );
    and g5900 ( n5011 , n8712 , n11092 );
    xnor g5901 ( n2262 , n11183 , n10791 );
    and g5902 ( n9476 , n7445 , n216 );
    xnor g5903 ( n3200 , n9505 , n10596 );
    not g5904 ( n2037 , n3244 );
    xnor g5905 ( n8284 , n8812 , n9532 );
    and g5906 ( n8261 , n197 , n8785 );
    not g5907 ( n7749 , n9347 );
    not g5908 ( n3825 , n510 );
    and g5909 ( n4073 , n6348 , n6936 );
    not g5910 ( n10466 , n10390 );
    xnor g5911 ( n2376 , n7556 , n12291 );
    and g5912 ( n7099 , n6279 , n4634 );
    nor g5913 ( n12801 , n2925 , n4583 );
    or g5914 ( n1396 , n5888 , n6572 );
    and g5915 ( n2419 , n9216 , n411 );
    and g5916 ( n11513 , n5568 , n12853 );
    and g5917 ( n8670 , n3969 , n10945 );
    xnor g5918 ( n10758 , n9234 , n10637 );
    and g5919 ( n11422 , n12635 , n9922 );
    or g5920 ( n9789 , n8598 , n1985 );
    and g5921 ( n10276 , n9265 , n9286 );
    xnor g5922 ( n4425 , n10498 , n5515 );
    xnor g5923 ( n10176 , n2027 , n6728 );
    or g5924 ( n6637 , n449 , n10302 );
    and g5925 ( n7768 , n3478 , n5537 );
    or g5926 ( n4491 , n11037 , n9223 );
    xnor g5927 ( n2438 , n10709 , n4413 );
    not g5928 ( n12994 , n5642 );
    xnor g5929 ( n5761 , n7881 , n11477 );
    or g5930 ( n4176 , n6778 , n12110 );
    not g5931 ( n12249 , n11180 );
    xnor g5932 ( n10003 , n12216 , n9563 );
    xnor g5933 ( n8365 , n1359 , n2438 );
    and g5934 ( n12640 , n11707 , n6358 );
    or g5935 ( n11108 , n12396 , n6978 );
    or g5936 ( n207 , n1345 , n10029 );
    xnor g5937 ( n11190 , n6417 , n8399 );
    or g5938 ( n12022 , n3127 , n8563 );
    xnor g5939 ( n9991 , n235 , n4816 );
    not g5940 ( n9808 , n11537 );
    or g5941 ( n8812 , n5688 , n8030 );
    and g5942 ( n6907 , n7918 , n1470 );
    xnor g5943 ( n7205 , n4139 , n6698 );
    or g5944 ( n910 , n12683 , n10617 );
    xnor g5945 ( n6073 , n1774 , n83 );
    and g5946 ( n9231 , n8167 , n3341 );
    nor g5947 ( n12931 , n13200 , n6779 );
    or g5948 ( n1648 , n1023 , n5202 );
    xnor g5949 ( n264 , n8593 , n8921 );
    xnor g5950 ( n1498 , n7000 , n4394 );
    or g5951 ( n12264 , n2768 , n4230 );
    xnor g5952 ( n179 , n2010 , n7685 );
    nor g5953 ( n9030 , n5612 , n5413 );
    not g5954 ( n10481 , n1636 );
    or g5955 ( n1675 , n10509 , n4844 );
    not g5956 ( n3640 , n5536 );
    not g5957 ( n10229 , n9948 );
    and g5958 ( n2555 , n7171 , n11684 );
    xnor g5959 ( n12736 , n3244 , n7107 );
    not g5960 ( n4462 , n9915 );
    xnor g5961 ( n4014 , n8473 , n3410 );
    xnor g5962 ( n590 , n3115 , n6185 );
    not g5963 ( n10204 , n1327 );
    or g5964 ( n3978 , n13025 , n3981 );
    or g5965 ( n7543 , n4621 , n121 );
    xnor g5966 ( n4304 , n10183 , n11931 );
    and g5967 ( n2575 , n5922 , n7874 );
    or g5968 ( n2946 , n1957 , n5408 );
    xor g5969 ( n11610 , n12417 , n10376 );
    or g5970 ( n8389 , n5086 , n4515 );
    or g5971 ( n3684 , n8106 , n5317 );
    and g5972 ( n4865 , n10619 , n300 );
    xnor g5973 ( n10062 , n85 , n2857 );
    and g5974 ( n551 , n6571 , n11124 );
    or g5975 ( n6051 , n3225 , n7935 );
    xnor g5976 ( n5026 , n8620 , n8866 );
    or g5977 ( n1483 , n8325 , n1043 );
    or g5978 ( n10919 , n2614 , n1463 );
    not g5979 ( n5630 , n8394 );
    not g5980 ( n11328 , n7040 );
    and g5981 ( n12016 , n11754 , n8426 );
    not g5982 ( n12738 , n9367 );
    or g5983 ( n7845 , n12174 , n1043 );
    xnor g5984 ( n3180 , n4797 , n9311 );
    or g5985 ( n9169 , n2128 , n12910 );
    not g5986 ( n3062 , n12352 );
    or g5987 ( n10544 , n8941 , n10016 );
    xnor g5988 ( n9843 , n1232 , n10946 );
    nor g5989 ( n10665 , n1984 , n8963 );
    or g5990 ( n1328 , n5190 , n12787 );
    xnor g5991 ( n13220 , n8579 , n4008 );
    not g5992 ( n6055 , n3286 );
    xnor g5993 ( n995 , n4302 , n2539 );
    xnor g5994 ( n4280 , n5417 , n4541 );
    or g5995 ( n10704 , n2217 , n479 );
    or g5996 ( n10064 , n12153 , n776 );
    or g5997 ( n4379 , n7672 , n4373 );
    and g5998 ( n3203 , n2145 , n7006 );
    nor g5999 ( n7997 , n622 , n7307 );
    xnor g6000 ( n2779 , n1316 , n8395 );
    xnor g6001 ( n2200 , n6298 , n12529 );
    xnor g6002 ( n904 , n9539 , n5625 );
    or g6003 ( n4766 , n10664 , n8519 );
    or g6004 ( n7688 , n9281 , n6623 );
    or g6005 ( n965 , n8498 , n8268 );
    nor g6006 ( n3758 , n7896 , n851 );
    xnor g6007 ( n1408 , n12131 , n12223 );
    not g6008 ( n6538 , n12452 );
    and g6009 ( n4532 , n3311 , n10408 );
    nor g6010 ( n7893 , n7542 , n4534 );
    or g6011 ( n12097 , n1191 , n1463 );
    xnor g6012 ( n11618 , n2021 , n12937 );
    or g6013 ( n2011 , n9282 , n7158 );
    or g6014 ( n7126 , n6250 , n9159 );
    not g6015 ( n12493 , n11574 );
    xnor g6016 ( n5394 , n6211 , n8388 );
    xnor g6017 ( n6932 , n7284 , n4407 );
    and g6018 ( n4472 , n250 , n2492 );
    not g6019 ( n12576 , n5600 );
    and g6020 ( n6234 , n10092 , n3368 );
    xnor g6021 ( n4726 , n2344 , n4956 );
    or g6022 ( n4912 , n2254 , n237 );
    and g6023 ( n2530 , n6074 , n11191 );
    not g6024 ( n7962 , n9514 );
    xnor g6025 ( n10543 , n348 , n4177 );
    or g6026 ( n11533 , n1634 , n12621 );
    or g6027 ( n5948 , n2786 , n8972 );
    not g6028 ( n69 , n772 );
    or g6029 ( n2024 , n3854 , n6404 );
    or g6030 ( n5822 , n7319 , n12764 );
    and g6031 ( n10734 , n5840 , n101 );
    or g6032 ( n5932 , n6439 , n12273 );
    and g6033 ( n3779 , n11650 , n1121 );
    or g6034 ( n6315 , n5927 , n10292 );
    xnor g6035 ( n7964 , n6777 , n10205 );
    and g6036 ( n7692 , n9995 , n7598 );
    not g6037 ( n10590 , n6782 );
    or g6038 ( n7427 , n6182 , n9223 );
    or g6039 ( n3420 , n2726 , n3949 );
    xnor g6040 ( n5598 , n2706 , n687 );
    not g6041 ( n3898 , n11180 );
    not g6042 ( n2411 , n12156 );
    and g6043 ( n9514 , n11197 , n1078 );
    xnor g6044 ( n9796 , n9930 , n2565 );
    or g6045 ( n10141 , n2563 , n1509 );
    xnor g6046 ( n10751 , n4948 , n268 );
    or g6047 ( n7506 , n12778 , n11922 );
    xnor g6048 ( n4590 , n7709 , n10000 );
    and g6049 ( n3971 , n3018 , n6951 );
    and g6050 ( n10754 , n12402 , n10456 );
    not g6051 ( n5670 , n7812 );
    and g6052 ( n3071 , n2381 , n5778 );
    or g6053 ( n6777 , n10334 , n10179 );
    or g6054 ( n11010 , n4642 , n2626 );
    not g6055 ( n2325 , n10904 );
    and g6056 ( n9769 , n4289 , n8878 );
    or g6057 ( n1431 , n2558 , n4056 );
    nor g6058 ( n1640 , n10782 , n12379 );
    and g6059 ( n6343 , n11207 , n3033 );
    and g6060 ( n5878 , n10988 , n4831 );
    not g6061 ( n5002 , n7697 );
    xnor g6062 ( n12235 , n3687 , n10803 );
    not g6063 ( n12846 , n892 );
    or g6064 ( n1332 , n5205 , n2907 );
    nor g6065 ( n3504 , n95 , n146 );
    not g6066 ( n9838 , n12020 );
    not g6067 ( n3892 , n2498 );
    and g6068 ( n2527 , n5942 , n5892 );
    xnor g6069 ( n8528 , n7845 , n13098 );
    xnor g6070 ( n6102 , n7713 , n5311 );
    and g6071 ( n6618 , n11341 , n1954 );
    xnor g6072 ( n10575 , n1667 , n11372 );
    buf g6073 ( n6635 , n4696 );
    not g6074 ( n2742 , n1611 );
    not g6075 ( n12789 , n11030 );
    or g6076 ( n11651 , n4185 , n8268 );
    not g6077 ( n9450 , n10805 );
    and g6078 ( n2021 , n3092 , n11740 );
    nor g6079 ( n7624 , n5938 , n2410 );
    nor g6080 ( n3941 , n3189 , n682 );
    and g6081 ( n4762 , n4759 , n2665 );
    not g6082 ( n5409 , n8684 );
    or g6083 ( n5542 , n4995 , n9792 );
    xnor g6084 ( n10930 , n3880 , n11670 );
    and g6085 ( n1558 , n2994 , n10713 );
    not g6086 ( n2473 , n10343 );
    xnor g6087 ( n10042 , n7369 , n7808 );
    not g6088 ( n2688 , n817 );
    or g6089 ( n608 , n10580 , n815 );
    xnor g6090 ( n105 , n4038 , n4424 );
    or g6091 ( n6980 , n6479 , n1653 );
    or g6092 ( n12664 , n2175 , n7873 );
    and g6093 ( n4729 , n10682 , n10896 );
    xnor g6094 ( n3362 , n3633 , n12863 );
    not g6095 ( n9181 , n1636 );
    and g6096 ( n4186 , n139 , n3853 );
    nor g6097 ( n1079 , n3919 , n12108 );
    and g6098 ( n3909 , n5671 , n8290 );
    or g6099 ( n10997 , n4087 , n8686 );
    nor g6100 ( n11359 , n1815 , n3555 );
    and g6101 ( n12140 , n4104 , n8186 );
    xnor g6102 ( n1281 , n4589 , n11503 );
    xnor g6103 ( n6598 , n11378 , n1661 );
    xnor g6104 ( n5309 , n2186 , n92 );
    or g6105 ( n3781 , n5500 , n11475 );
    nor g6106 ( n7039 , n1809 , n4287 );
    or g6107 ( n1240 , n6721 , n1144 );
    xnor g6108 ( n6617 , n10584 , n9911 );
    not g6109 ( n821 , n6357 );
    xnor g6110 ( n5563 , n3333 , n7478 );
    or g6111 ( n889 , n5999 , n2599 );
    nor g6112 ( n3236 , n9042 , n10612 );
    or g6113 ( n4283 , n6486 , n4640 );
    not g6114 ( n9283 , n12373 );
    xnor g6115 ( n4613 , n12697 , n7640 );
    and g6116 ( n5291 , n12253 , n3486 );
    or g6117 ( n5896 , n9113 , n8490 );
    buf g6118 ( n12273 , n5550 );
    xnor g6119 ( n12867 , n4400 , n3994 );
    and g6120 ( n10904 , n934 , n6674 );
    and g6121 ( n6582 , n8085 , n4679 );
    or g6122 ( n6657 , n13168 , n12188 );
    not g6123 ( n7119 , n3076 );
    nor g6124 ( n10902 , n8986 , n11601 );
    xnor g6125 ( n2708 , n12355 , n12264 );
    not g6126 ( n9492 , n411 );
    and g6127 ( n11387 , n9718 , n5933 );
    or g6128 ( n4224 , n8672 , n12188 );
    and g6129 ( n7643 , n12130 , n12181 );
    xor g6130 ( n1280 , n6644 , n2547 );
    and g6131 ( n11531 , n10491 , n13180 );
    not g6132 ( n11365 , n1717 );
    or g6133 ( n5306 , n1671 , n7323 );
    xnor g6134 ( n7584 , n2219 , n7509 );
    or g6135 ( n10353 , n207 , n12290 );
    xor g6136 ( n12993 , n2762 , n11154 );
    xnor g6137 ( n1862 , n8690 , n6995 );
    or g6138 ( n5537 , n2228 , n1570 );
    or g6139 ( n519 , n8050 , n663 );
    and g6140 ( n8767 , n12667 , n1787 );
    or g6141 ( n11442 , n3071 , n341 );
    or g6142 ( n3122 , n6769 , n6265 );
    not g6143 ( n11972 , n11939 );
    or g6144 ( n13214 , n10681 , n12596 );
    xnor g6145 ( n5498 , n1603 , n3455 );
    not g6146 ( n5839 , n8311 );
    or g6147 ( n7181 , n3908 , n1144 );
    xnor g6148 ( n1731 , n10911 , n8201 );
    xnor g6149 ( n3540 , n4147 , n1981 );
    not g6150 ( n11354 , n10642 );
    or g6151 ( n10585 , n10586 , n12126 );
    or g6152 ( n6449 , n6753 , n8573 );
    xnor g6153 ( n11272 , n7398 , n8287 );
    xnor g6154 ( n11766 , n9341 , n2161 );
    and g6155 ( n30 , n554 , n3975 );
    xnor g6156 ( n3611 , n7767 , n10372 );
    or g6157 ( n11009 , n7780 , n10106 );
    and g6158 ( n12815 , n1070 , n12169 );
    or g6159 ( n7015 , n5972 , n4987 );
    not g6160 ( n7709 , n9515 );
    or g6161 ( n10460 , n106 , n1266 );
    not g6162 ( n5446 , n6707 );
    and g6163 ( n12116 , n1973 , n6302 );
    xnor g6164 ( n4632 , n12670 , n10971 );
    or g6165 ( n6707 , n1402 , n9223 );
    buf g6166 ( n8534 , n6596 );
    not g6167 ( n11540 , n8745 );
    or g6168 ( n8334 , n10924 , n2787 );
    xnor g6169 ( n8713 , n3796 , n5325 );
    xnor g6170 ( n11698 , n11733 , n9815 );
    xnor g6171 ( n3612 , n8814 , n9560 );
    not g6172 ( n4080 , n497 );
    xnor g6173 ( n8069 , n3810 , n4918 );
    xnor g6174 ( n6648 , n9331 , n4625 );
    and g6175 ( n822 , n7926 , n1334 );
    and g6176 ( n4196 , n1391 , n10967 );
    buf g6177 ( n12695 , n2278 );
    not g6178 ( n6533 , n4188 );
    xnor g6179 ( n6605 , n2312 , n12685 );
    or g6180 ( n11235 , n1402 , n2059 );
    and g6181 ( n2917 , n8751 , n8344 );
    xnor g6182 ( n4577 , n8366 , n7176 );
    not g6183 ( n9402 , n7896 );
    buf g6184 ( n5797 , n2278 );
    not g6185 ( n9586 , n12248 );
    or g6186 ( n2144 , n2538 , n3949 );
    or g6187 ( n13066 , n6908 , n5819 );
    and g6188 ( n3843 , n5900 , n9781 );
    and g6189 ( n5596 , n1332 , n11463 );
    or g6190 ( n9443 , n7068 , n9159 );
    not g6191 ( n12171 , n4651 );
    nor g6192 ( n4571 , n12981 , n6272 );
    xnor g6193 ( n5244 , n7869 , n754 );
    and g6194 ( n9106 , n12322 , n12374 );
    xnor g6195 ( n6213 , n7926 , n236 );
    not g6196 ( n8835 , n2577 );
    or g6197 ( n6951 , n12469 , n12273 );
    and g6198 ( n164 , n4761 , n6013 );
    or g6199 ( n12310 , n10775 , n9956 );
    xnor g6200 ( n8373 , n12073 , n8003 );
    not g6201 ( n3761 , n10288 );
    or g6202 ( n4279 , n7966 , n6404 );
    nor g6203 ( n1803 , n5399 , n7405 );
    and g6204 ( n9134 , n1652 , n10419 );
    not g6205 ( n10035 , n2212 );
    or g6206 ( n8559 , n6595 , n7935 );
    xnor g6207 ( n10192 , n12518 , n12024 );
    xor g6208 ( n9580 , n3365 , n11819 );
    nor g6209 ( n3733 , n3868 , n11143 );
    or g6210 ( n12311 , n5803 , n3193 );
    xnor g6211 ( n158 , n13050 , n5106 );
    or g6212 ( n3786 , n4451 , n5725 );
    not g6213 ( n8843 , n1302 );
    or g6214 ( n5867 , n11455 , n10374 );
    xnor g6215 ( n825 , n11562 , n12497 );
    nor g6216 ( n10443 , n12437 , n3799 );
    or g6217 ( n267 , n10314 , n12959 );
    and g6218 ( n2500 , n5207 , n3707 );
    and g6219 ( n10564 , n11014 , n4770 );
    or g6220 ( n4938 , n7283 , n12273 );
    nor g6221 ( n4388 , n4500 , n1 );
    or g6222 ( n2345 , n3619 , n13053 );
    not g6223 ( n10263 , n10162 );
    or g6224 ( n2370 , n1218 , n5242 );
    not g6225 ( n2387 , n6168 );
    or g6226 ( n5199 , n13063 , n5493 );
    not g6227 ( n10519 , n12078 );
    or g6228 ( n11194 , n7091 , n3438 );
    and g6229 ( n1417 , n11420 , n2363 );
    and g6230 ( n11817 , n3750 , n11399 );
    nor g6231 ( n2019 , n10496 , n5159 );
    and g6232 ( n5248 , n3325 , n4942 );
    xor g6233 ( n1068 , n10979 , n8875 );
    and g6234 ( n8642 , n11703 , n8853 );
    and g6235 ( n976 , n2717 , n6920 );
    nor g6236 ( n3484 , n10967 , n1391 );
    xnor g6237 ( n9351 , n11602 , n8100 );
    nor g6238 ( n11437 , n5621 , n5533 );
    nor g6239 ( n7203 , n6656 , n10036 );
    nor g6240 ( n13070 , n914 , n592 );
    and g6241 ( n2939 , n9253 , n7972 );
    or g6242 ( n3304 , n696 , n9352 );
    not g6243 ( n8111 , n1792 );
    or g6244 ( n408 , n5968 , n10179 );
    or g6245 ( n7457 , n1554 , n6133 );
    and g6246 ( n6565 , n9757 , n6131 );
    xnor g6247 ( n120 , n12035 , n2939 );
    xnor g6248 ( n10638 , n8487 , n10394 );
    xnor g6249 ( n8056 , n8061 , n6084 );
    xnor g6250 ( n9007 , n1282 , n11529 );
    xnor g6251 ( n10790 , n2650 , n3569 );
    nor g6252 ( n2796 , n6536 , n4866 );
    not g6253 ( n10666 , n594 );
    xnor g6254 ( n5143 , n8942 , n6632 );
    xnor g6255 ( n1414 , n5850 , n187 );
    and g6256 ( n2667 , n4205 , n1351 );
    xnor g6257 ( n9631 , n9708 , n684 );
    or g6258 ( n11210 , n13194 , n10319 );
    not g6259 ( n13183 , n2295 );
    and g6260 ( n1245 , n1018 , n764 );
    xnor g6261 ( n88 , n7583 , n6168 );
    or g6262 ( n10610 , n5944 , n7305 );
    not g6263 ( n8561 , n9093 );
    xnor g6264 ( n4894 , n7657 , n6795 );
    or g6265 ( n565 , n5588 , n10029 );
    or g6266 ( n10646 , n1434 , n3459 );
    not g6267 ( n156 , n6489 );
    xnor g6268 ( n10954 , n12622 , n6470 );
    not g6269 ( n12246 , n2765 );
    nor g6270 ( n9985 , n4368 , n7716 );
    xnor g6271 ( n10504 , n3122 , n6477 );
    or g6272 ( n5503 , n7532 , n6635 );
    nor g6273 ( n11261 , n6668 , n7812 );
    not g6274 ( n3222 , n4457 );
    and g6275 ( n2617 , n4929 , n12060 );
    xnor g6276 ( n1591 , n676 , n6432 );
    and g6277 ( n9252 , n3224 , n1888 );
    not g6278 ( n11471 , n5747 );
    xnor g6279 ( n1164 , n4313 , n12029 );
    xnor g6280 ( n9756 , n11160 , n8069 );
    xnor g6281 ( n10156 , n1380 , n5254 );
    or g6282 ( n10351 , n10587 , n9159 );
    and g6283 ( n11822 , n10136 , n3174 );
    or g6284 ( n5337 , n5558 , n13043 );
    not g6285 ( n10558 , n12579 );
    and g6286 ( n3186 , n2931 , n7313 );
    xnor g6287 ( n12991 , n331 , n11994 );
    nor g6288 ( n3075 , n12381 , n4589 );
    not g6289 ( n9033 , n5498 );
    not g6290 ( n10383 , n2174 );
    and g6291 ( n2938 , n10631 , n10329 );
    xnor g6292 ( n535 , n10327 , n10074 );
    xnor g6293 ( n2139 , n9945 , n3513 );
    nor g6294 ( n12907 , n6273 , n12145 );
    xnor g6295 ( n12034 , n9039 , n2775 );
    or g6296 ( n1970 , n513 , n9027 );
    xnor g6297 ( n11305 , n3834 , n9411 );
    xnor g6298 ( n8015 , n9870 , n1104 );
    or g6299 ( n7669 , n11781 , n902 );
    not g6300 ( n8644 , n9474 );
    and g6301 ( n7321 , n1126 , n13083 );
    not g6302 ( n493 , n12853 );
    and g6303 ( n4812 , n12569 , n7508 );
    and g6304 ( n10806 , n9619 , n5382 );
    and g6305 ( n2250 , n2753 , n7593 );
    not g6306 ( n5494 , n6043 );
    and g6307 ( n2023 , n2725 , n13228 );
    xnor g6308 ( n12776 , n7316 , n4510 );
    xnor g6309 ( n11303 , n2656 , n323 );
    not g6310 ( n1263 , n4789 );
    or g6311 ( n7420 , n1485 , n5931 );
    xnor g6312 ( n8813 , n11278 , n8482 );
    not g6313 ( n7013 , n4259 );
    or g6314 ( n4 , n11242 , n2133 );
    or g6315 ( n8825 , n2504 , n8563 );
    not g6316 ( n12812 , n10654 );
    xnor g6317 ( n2909 , n2069 , n9030 );
    xnor g6318 ( n7637 , n8358 , n3087 );
    not g6319 ( n10525 , n1988 );
    xnor g6320 ( n7764 , n10812 , n5074 );
    xnor g6321 ( n1121 , n6555 , n12338 );
    not g6322 ( n8654 , n9580 );
    xor g6323 ( n5998 , n5659 , n11988 );
    or g6324 ( n4145 , n8510 , n8702 );
    or g6325 ( n13009 , n10558 , n7723 );
    xnor g6326 ( n9553 , n7555 , n2864 );
    and g6327 ( n4389 , n11249 , n13207 );
    or g6328 ( n11115 , n5574 , n5604 );
    xnor g6329 ( n1583 , n6305 , n984 );
    and g6330 ( n2751 , n1905 , n2608 );
    not g6331 ( n8026 , n1498 );
    not g6332 ( n10988 , n13034 );
    xnor g6333 ( n3678 , n2431 , n11169 );
    not g6334 ( n2580 , n11671 );
    xnor g6335 ( n4626 , n7585 , n9947 );
    xnor g6336 ( n2888 , n4035 , n8902 );
    not g6337 ( n7771 , n12340 );
    and g6338 ( n1794 , n12230 , n4204 );
    or g6339 ( n8668 , n7000 , n10937 );
    xnor g6340 ( n8459 , n11899 , n2926 );
    or g6341 ( n2015 , n2031 , n10130 );
    or g6342 ( n3326 , n950 , n3257 );
    or g6343 ( n2613 , n10474 , n5782 );
    not g6344 ( n7700 , n13060 );
    and g6345 ( n7353 , n5883 , n7653 );
    nor g6346 ( n3179 , n10259 , n12454 );
    or g6347 ( n5441 , n5973 , n8563 );
    and g6348 ( n3995 , n103 , n10408 );
    or g6349 ( n5233 , n9606 , n12188 );
    and g6350 ( n3559 , n6135 , n4859 );
    not g6351 ( n3334 , n11386 );
    xnor g6352 ( n10074 , n6711 , n2523 );
    or g6353 ( n10096 , n6726 , n7530 );
    nor g6354 ( n9126 , n6431 , n8826 );
    xnor g6355 ( n4060 , n5098 , n3647 );
    or g6356 ( n1200 , n13181 , n1589 );
    or g6357 ( n7105 , n6658 , n7221 );
    and g6358 ( n3716 , n8471 , n6688 );
    and g6359 ( n9657 , n11313 , n883 );
    nor g6360 ( n3717 , n4710 , n3840 );
    not g6361 ( n9118 , n5962 );
    or g6362 ( n5139 , n6595 , n7903 );
    and g6363 ( n5722 , n10144 , n8545 );
    or g6364 ( n6739 , n3465 , n10222 );
    not g6365 ( n9765 , n4968 );
    nor g6366 ( n10576 , n12994 , n4422 );
    xnor g6367 ( n3748 , n9151 , n2664 );
    xnor g6368 ( n4240 , n1116 , n3670 );
    or g6369 ( n1868 , n8392 , n9159 );
    or g6370 ( n11361 , n1360 , n3531 );
    not g6371 ( n8834 , n90 );
    xnor g6372 ( n7212 , n7427 , n9203 );
    not g6373 ( n9697 , n2011 );
    not g6374 ( n12930 , n4470 );
    xnor g6375 ( n6413 , n2739 , n975 );
    xnor g6376 ( n1993 , n5025 , n523 );
    xnor g6377 ( n12650 , n9974 , n11747 );
    not g6378 ( n11242 , n12408 );
    and g6379 ( n3702 , n13163 , n2440 );
    not g6380 ( n8504 , n429 );
    or g6381 ( n2442 , n813 , n10029 );
    xnor g6382 ( n10271 , n6539 , n12257 );
    not g6383 ( n8039 , n5513 );
    xnor g6384 ( n4623 , n9168 , n9639 );
    xor g6385 ( n2630 , n11366 , n4269 );
    not g6386 ( n9265 , n10231 );
    not g6387 ( n11781 , n4470 );
    not g6388 ( n5713 , n12651 );
    or g6389 ( n7657 , n6733 , n1570 );
    nor g6390 ( n10957 , n8417 , n10011 );
    or g6391 ( n9025 , n7184 , n6635 );
    not g6392 ( n13242 , n11537 );
    not g6393 ( n4680 , n3447 );
    xor g6394 ( n7577 , n5544 , n10149 );
    or g6395 ( n11462 , n10429 , n252 );
    xnor g6396 ( n9817 , n12797 , n4726 );
    xnor g6397 ( n11882 , n8520 , n4329 );
    xnor g6398 ( n5384 , n8811 , n6932 );
    or g6399 ( n10851 , n2985 , n9704 );
    xnor g6400 ( n12040 , n8794 , n11814 );
    and g6401 ( n8001 , n7065 , n12180 );
    not g6402 ( n6768 , n4006 );
    nor g6403 ( n2531 , n12710 , n4193 );
    not g6404 ( n7346 , n5933 );
    and g6405 ( n6281 , n3363 , n2680 );
    xor g6406 ( n6197 , n10796 , n12058 );
    or g6407 ( n1136 , n10900 , n2449 );
    not g6408 ( n6421 , n7670 );
    not g6409 ( n585 , n1432 );
    xnor g6410 ( n6294 , n6130 , n8780 );
    and g6411 ( n9295 , n7269 , n9342 );
    or g6412 ( n7850 , n5595 , n2875 );
    not g6413 ( n5927 , n10004 );
    xnor g6414 ( n11604 , n11655 , n738 );
    or g6415 ( n3856 , n7941 , n4868 );
    or g6416 ( n5711 , n3697 , n7655 );
    xnor g6417 ( n4246 , n11987 , n3019 );
    xnor g6418 ( n1088 , n11998 , n6051 );
    not g6419 ( n617 , n8233 );
    xnor g6420 ( n12644 , n15 , n3056 );
    or g6421 ( n5411 , n2013 , n6484 );
    and g6422 ( n8566 , n11258 , n11967 );
    or g6423 ( n4753 , n7124 , n11550 );
    or g6424 ( n4965 , n13084 , n12501 );
    not g6425 ( n2943 , n13058 );
    and g6426 ( n4954 , n3128 , n3203 );
    xnor g6427 ( n6476 , n3627 , n13212 );
    xnor g6428 ( n8269 , n10999 , n10342 );
    or g6429 ( n8618 , n4584 , n4373 );
    xnor g6430 ( n415 , n9261 , n11977 );
    not g6431 ( n12335 , n12003 );
    nor g6432 ( n11208 , n1205 , n2649 );
    xnor g6433 ( n3952 , n12362 , n3987 );
    nor g6434 ( n7983 , n1395 , n8781 );
    xnor g6435 ( n3482 , n10371 , n13015 );
    and g6436 ( n2700 , n579 , n7977 );
    or g6437 ( n9884 , n7018 , n3016 );
    nor g6438 ( n1656 , n2107 , n8548 );
    or g6439 ( n452 , n216 , n7445 );
    not g6440 ( n241 , n9534 );
    or g6441 ( n13169 , n2711 , n9268 );
    nor g6442 ( n8004 , n12186 , n6163 );
    xor g6443 ( n12422 , n7919 , n11056 );
    not g6444 ( n4818 , n1612 );
    or g6445 ( n4927 , n5666 , n12273 );
    xnor g6446 ( n12923 , n8889 , n6022 );
    or g6447 ( n2792 , n5923 , n1026 );
    or g6448 ( n6835 , n3347 , n5036 );
    or g6449 ( n11142 , n4514 , n11244 );
    or g6450 ( n1888 , n1621 , n2133 );
    not g6451 ( n1152 , n10451 );
    or g6452 ( n10316 , n3587 , n9223 );
    xnor g6453 ( n7000 , n8028 , n4162 );
    xnor g6454 ( n3850 , n3628 , n9218 );
    not g6455 ( n2941 , n5066 );
    and g6456 ( n6012 , n11886 , n4025 );
    xnor g6457 ( n8839 , n4876 , n769 );
    and g6458 ( n8445 , n3732 , n7438 );
    and g6459 ( n7429 , n9332 , n5818 );
    or g6460 ( n6712 , n5890 , n8534 );
    or g6461 ( n11315 , n12514 , n514 );
    nor g6462 ( n3955 , n11306 , n8432 );
    not g6463 ( n11605 , n7326 );
    not g6464 ( n1536 , n8332 );
    xnor g6465 ( n1455 , n9236 , n5023 );
    and g6466 ( n10526 , n12517 , n7303 );
    xnor g6467 ( n11319 , n8800 , n7628 );
    or g6468 ( n12018 , n13061 , n1212 );
    not g6469 ( n7142 , n1198 );
    not g6470 ( n5923 , n5189 );
    not g6471 ( n7798 , n2339 );
    or g6472 ( n2900 , n8556 , n11772 );
    xor g6473 ( n12014 , n1268 , n3865 );
    and g6474 ( n9686 , n11943 , n2305 );
    and g6475 ( n581 , n4737 , n1785 );
    or g6476 ( n11192 , n2689 , n8702 );
    or g6477 ( n432 , n8141 , n11510 );
    and g6478 ( n8125 , n8183 , n5920 );
    and g6479 ( n6562 , n4905 , n10703 );
    or g6480 ( n2400 , n1406 , n5999 );
    not g6481 ( n5890 , n2737 );
    and g6482 ( n1782 , n3266 , n2224 );
    or g6483 ( n2096 , n5004 , n4314 );
    xnor g6484 ( n10554 , n10921 , n11675 );
    not g6485 ( n8836 , n3116 );
    and g6486 ( n3550 , n1669 , n1185 );
    xnor g6487 ( n2921 , n2439 , n1049 );
    xnor g6488 ( n12406 , n1655 , n10082 );
    nor g6489 ( n12505 , n12867 , n11079 );
    xnor g6490 ( n7717 , n6009 , n9055 );
    not g6491 ( n8664 , n7090 );
    or g6492 ( n4538 , n7142 , n2675 );
    or g6493 ( n6602 , n8697 , n10648 );
    or g6494 ( n4097 , n6988 , n11591 );
    xnor g6495 ( n9644 , n3848 , n7484 );
    xnor g6496 ( n7425 , n11189 , n6512 );
    or g6497 ( n11069 , n10954 , n4504 );
    xor g6498 ( n6484 , n6132 , n6094 );
    xnor g6499 ( n9183 , n4224 , n9864 );
    xnor g6500 ( n2561 , n6690 , n7141 );
    not g6501 ( n3908 , n6655 );
    and g6502 ( n10024 , n10800 , n8019 );
    nor g6503 ( n7422 , n744 , n12484 );
    not g6504 ( n8020 , n1709 );
    not g6505 ( n2723 , n8768 );
    or g6506 ( n11706 , n1387 , n4565 );
    not g6507 ( n12552 , n11891 );
    xnor g6508 ( n4319 , n9213 , n7651 );
    not g6509 ( n9828 , n1573 );
    xnor g6510 ( n6831 , n4146 , n4623 );
    xnor g6511 ( n10720 , n9519 , n6541 );
    nor g6512 ( n7063 , n4012 , n8189 );
    xnor g6513 ( n6192 , n978 , n11009 );
    or g6514 ( n5459 , n11718 , n5081 );
    xnor g6515 ( n10330 , n7763 , n5578 );
    not g6516 ( n10210 , n7637 );
    xnor g6517 ( n948 , n10795 , n12667 );
    or g6518 ( n4826 , n12441 , n4063 );
    and g6519 ( n1232 , n1420 , n8387 );
    xnor g6520 ( n137 , n3069 , n8365 );
    xnor g6521 ( n8807 , n12472 , n1926 );
    not g6522 ( n3041 , n9381 );
    xnor g6523 ( n5147 , n2814 , n12123 );
    or g6524 ( n5511 , n9422 , n1109 );
    xnor g6525 ( n11390 , n7002 , n7308 );
    or g6526 ( n10157 , n11903 , n5765 );
    or g6527 ( n3814 , n555 , n5677 );
    not g6528 ( n6645 , n3645 );
    not g6529 ( n1324 , n4233 );
    not g6530 ( n5243 , n741 );
    not g6531 ( n1406 , n9887 );
    or g6532 ( n400 , n2566 , n7624 );
    xor g6533 ( n8689 , n1495 , n4518 );
    xnor g6534 ( n3057 , n3394 , n12392 );
    nor g6535 ( n12053 , n672 , n2912 );
    or g6536 ( n1779 , n9767 , n8030 );
    nor g6537 ( n12456 , n8470 , n5469 );
    and g6538 ( n1361 , n10232 , n9520 );
    not g6539 ( n12099 , n9849 );
    or g6540 ( n3545 , n3369 , n6227 );
    xnor g6541 ( n70 , n7240 , n735 );
    or g6542 ( n5649 , n12834 , n2449 );
    and g6543 ( n5677 , n8663 , n6476 );
    and g6544 ( n12133 , n8466 , n7720 );
    xnor g6545 ( n1100 , n6842 , n86 );
    or g6546 ( n3439 , n7377 , n9075 );
    and g6547 ( n3481 , n12418 , n11713 );
    not g6548 ( n10492 , n12389 );
    or g6549 ( n12726 , n10772 , n11144 );
    xnor g6550 ( n1249 , n9056 , n7612 );
    xnor g6551 ( n1208 , n12824 , n6897 );
    not g6552 ( n3509 , n3112 );
    or g6553 ( n11156 , n7891 , n8048 );
    xnor g6554 ( n5178 , n3354 , n10367 );
    and g6555 ( n4700 , n12838 , n4479 );
    or g6556 ( n6159 , n6738 , n9486 );
    not g6557 ( n80 , n951 );
    or g6558 ( n4128 , n10281 , n206 );
    or g6559 ( n7568 , n8035 , n6565 );
    xnor g6560 ( n6310 , n4277 , n9908 );
    or g6561 ( n6453 , n7033 , n5521 );
    not g6562 ( n6219 , n841 );
    or g6563 ( n2826 , n79 , n4442 );
    or g6564 ( n6953 , n12000 , n4253 );
    or g6565 ( n6748 , n3892 , n12069 );
    xnor g6566 ( n11001 , n10918 , n3528 );
    xnor g6567 ( n7663 , n4772 , n12495 );
    xnor g6568 ( n8958 , n11064 , n5237 );
    and g6569 ( n1344 , n3602 , n6807 );
    or g6570 ( n2070 , n8950 , n6635 );
    or g6571 ( n13134 , n5520 , n10761 );
    or g6572 ( n10359 , n1706 , n4643 );
    and g6573 ( n356 , n8221 , n7261 );
    nor g6574 ( n276 , n9456 , n1754 );
    xnor g6575 ( n8089 , n10690 , n10095 );
    not g6576 ( n8285 , n6142 );
    not g6577 ( n8971 , n253 );
    not g6578 ( n6706 , n1486 );
    and g6579 ( n2195 , n13056 , n385 );
    and g6580 ( n2935 , n521 , n11039 );
    or g6581 ( n876 , n5125 , n12077 );
    xnor g6582 ( n12369 , n7889 , n2685 );
    not g6583 ( n11106 , n12784 );
    xnor g6584 ( n11894 , n2851 , n9121 );
    or g6585 ( n6890 , n11009 , n12387 );
    and g6586 ( n374 , n7017 , n1970 );
    xnor g6587 ( n11762 , n921 , n10650 );
    nor g6588 ( n7712 , n9448 , n6483 );
    xnor g6589 ( n6622 , n6208 , n352 );
    or g6590 ( n8620 , n6846 , n3703 );
    or g6591 ( n9854 , n12084 , n13054 );
    xnor g6592 ( n2719 , n13223 , n12822 );
    not g6593 ( n47 , n5551 );
    or g6594 ( n9716 , n1903 , n10931 );
    or g6595 ( n1460 , n7047 , n12783 );
    xnor g6596 ( n2928 , n6527 , n7278 );
    not g6597 ( n12848 , n13120 );
    and g6598 ( n325 , n5031 , n8506 );
    or g6599 ( n8683 , n2232 , n2958 );
    or g6600 ( n8344 , n1559 , n6919 );
    or g6601 ( n1683 , n1571 , n7530 );
    not g6602 ( n9069 , n6392 );
    or g6603 ( n38 , n6672 , n13238 );
    or g6604 ( n6723 , n5943 , n8730 );
    xnor g6605 ( n3876 , n3536 , n6857 );
    xnor g6606 ( n4553 , n10790 , n4083 );
    xnor g6607 ( n2202 , n12394 , n11863 );
    or g6608 ( n7861 , n7620 , n9195 );
    and g6609 ( n4320 , n7529 , n7772 );
    and g6610 ( n12694 , n231 , n8906 );
    not g6611 ( n8592 , n4008 );
    nor g6612 ( n2320 , n12260 , n11433 );
    or g6613 ( n5009 , n4184 , n12725 );
    xor g6614 ( n12742 , n8839 , n1281 );
    or g6615 ( n6806 , n11599 , n7892 );
    xnor g6616 ( n8409 , n3642 , n5196 );
    not g6617 ( n5176 , n8768 );
    not g6618 ( n2415 , n4740 );
    xor g6619 ( n4788 , n4803 , n256 );
    and g6620 ( n523 , n12918 , n5246 );
    nor g6621 ( n7487 , n10913 , n3746 );
    not g6622 ( n3498 , n4470 );
    and g6623 ( n12005 , n10851 , n3275 );
    and g6624 ( n5781 , n9509 , n357 );
    xnor g6625 ( n8991 , n9448 , n7389 );
    xnor g6626 ( n8403 , n4654 , n1958 );
    nor g6627 ( n3891 , n7474 , n4068 );
    xnor g6628 ( n4417 , n9554 , n3849 );
    or g6629 ( n440 , n12871 , n12388 );
    or g6630 ( n3087 , n6769 , n1026 );
    and g6631 ( n10079 , n7331 , n5204 );
    not g6632 ( n8436 , n12603 );
    and g6633 ( n4835 , n13215 , n150 );
    xnor g6634 ( n11725 , n9523 , n11656 );
    or g6635 ( n7706 , n6724 , n7723 );
    xnor g6636 ( n3370 , n4251 , n3079 );
    not g6637 ( n10986 , n11445 );
    xnor g6638 ( n4614 , n4101 , n9357 );
    not g6639 ( n2207 , n8455 );
    and g6640 ( n5296 , n4667 , n10546 );
    or g6641 ( n3901 , n7884 , n12426 );
    and g6642 ( n9933 , n10228 , n3915 );
    not g6643 ( n9821 , n8036 );
    xnor g6644 ( n10399 , n10499 , n6893 );
    or g6645 ( n1763 , n3299 , n8301 );
    xnor g6646 ( n3324 , n6294 , n3034 );
    nor g6647 ( n13045 , n5505 , n13171 );
    not g6648 ( n8672 , n9669 );
    not g6649 ( n4361 , n1228 );
    and g6650 ( n1770 , n5314 , n188 );
    and g6651 ( n4687 , n9153 , n12001 );
    or g6652 ( n2266 , n8528 , n13237 );
    not g6653 ( n5105 , n4006 );
    and g6654 ( n11746 , n9928 , n9445 );
    not g6655 ( n7159 , n3064 );
    nor g6656 ( n12628 , n786 , n4428 );
    xnor g6657 ( n632 , n12637 , n2046 );
    not g6658 ( n3025 , n7316 );
    and g6659 ( n46 , n2826 , n10965 );
    xnor g6660 ( n1743 , n8689 , n6516 );
    not g6661 ( n1618 , n7720 );
    buf g6662 ( n10319 , n13005 );
    nor g6663 ( n833 , n2088 , n5851 );
    nor g6664 ( n6594 , n12707 , n5333 );
    not g6665 ( n3783 , n7360 );
    or g6666 ( n12771 , n11171 , n12273 );
    and g6667 ( n2152 , n3345 , n8112 );
    xnor g6668 ( n8818 , n10920 , n5975 );
    not g6669 ( n3132 , n3711 );
    nor g6670 ( n1856 , n10033 , n8669 );
    and g6671 ( n5071 , n2652 , n11369 );
    not g6672 ( n1226 , n1312 );
    and g6673 ( n7528 , n8146 , n169 );
    xor g6674 ( n485 , n2535 , n11741 );
    xnor g6675 ( n12956 , n11567 , n4999 );
    and g6676 ( n4093 , n10760 , n5330 );
    not g6677 ( n1750 , n8228 );
    and g6678 ( n504 , n3445 , n6581 );
    or g6679 ( n7213 , n7249 , n2836 );
    or g6680 ( n11989 , n10525 , n2212 );
    not g6681 ( n4143 , n7113 );
    and g6682 ( n323 , n508 , n6393 );
    xnor g6683 ( n7043 , n10743 , n6529 );
    or g6684 ( n7588 , n2858 , n8097 );
    or g6685 ( n3070 , n1571 , n12388 );
    xnor g6686 ( n10516 , n11893 , n6350 );
    xnor g6687 ( n11276 , n1547 , n466 );
    or g6688 ( n10940 , n1930 , n8348 );
    xnor g6689 ( n9542 , n4204 , n4241 );
    and g6690 ( n5311 , n4096 , n9072 );
    or g6691 ( n2302 , n4692 , n2351 );
    and g6692 ( n11846 , n9216 , n13058 );
    or g6693 ( n4433 , n6713 , n2989 );
    or g6694 ( n3227 , n9723 , n8030 );
    or g6695 ( n7112 , n4430 , n68 );
    xnor g6696 ( n6283 , n36 , n5219 );
    xnor g6697 ( n6794 , n1935 , n9587 );
    and g6698 ( n8627 , n1021 , n8628 );
    xnor g6699 ( n7740 , n2233 , n1421 );
    not g6700 ( n3681 , n8543 );
    or g6701 ( n3683 , n10481 , n9075 );
    xnor g6702 ( n637 , n382 , n3967 );
    xnor g6703 ( n6897 , n5188 , n13022 );
    and g6704 ( n7630 , n8396 , n11383 );
    nor g6705 ( n1322 , n8539 , n3525 );
    and g6706 ( n12672 , n7894 , n6300 );
    xnor g6707 ( n12457 , n3345 , n580 );
    or g6708 ( n7658 , n1571 , n8702 );
    or g6709 ( n5367 , n5810 , n3133 );
    not g6710 ( n10291 , n9667 );
    or g6711 ( n5144 , n3516 , n5547 );
    and g6712 ( n11796 , n4870 , n9487 );
    not g6713 ( n3963 , n3130 );
    or g6714 ( n2283 , n7223 , n3981 );
    and g6715 ( n10442 , n5644 , n7179 );
    xnor g6716 ( n6079 , n7669 , n10767 );
    not g6717 ( n1321 , n2630 );
    not g6718 ( n10877 , n4357 );
    and g6719 ( n12225 , n1797 , n9722 );
    and g6720 ( n12511 , n7771 , n3524 );
    not g6721 ( n11014 , n5777 );
    nor g6722 ( n3823 , n12675 , n3629 );
    not g6723 ( n7824 , n4543 );
    and g6724 ( n10436 , n993 , n6353 );
    xnor g6725 ( n750 , n1442 , n9967 );
    xnor g6726 ( n2966 , n877 , n12991 );
    xnor g6727 ( n2735 , n13172 , n2567 );
    not g6728 ( n7167 , n11634 );
    and g6729 ( n4560 , n4779 , n7832 );
    or g6730 ( n9743 , n9822 , n634 );
    or g6731 ( n10329 , n2914 , n655 );
    not g6732 ( n11297 , n10633 );
    not g6733 ( n9868 , n9570 );
    or g6734 ( n11433 , n6915 , n1710 );
    and g6735 ( n11267 , n4532 , n7279 );
    xnor g6736 ( n4262 , n6321 , n5780 );
    or g6737 ( n6095 , n3420 , n6123 );
    xnor g6738 ( n12459 , n12659 , n5351 );
    nor g6739 ( n12794 , n4112 , n4389 );
    xnor g6740 ( n8841 , n6384 , n13142 );
    nor g6741 ( n2251 , n11775 , n12139 );
    and g6742 ( n2319 , n8802 , n6235 );
    not g6743 ( n9431 , n3012 );
    not g6744 ( n2582 , n9887 );
    nor g6745 ( n4926 , n9624 , n4914 );
    xnor g6746 ( n8955 , n7264 , n1208 );
    and g6747 ( n7859 , n1680 , n451 );
    and g6748 ( n8435 , n2694 , n12528 );
    xnor g6749 ( n2934 , n8495 , n11048 );
    xnor g6750 ( n50 , n10695 , n12331 );
    or g6751 ( n3163 , n6774 , n10875 );
    nor g6752 ( n12946 , n3345 , n8112 );
    nor g6753 ( n6121 , n9548 , n1124 );
    and g6754 ( n1543 , n11174 , n13052 );
    xnor g6755 ( n8581 , n8652 , n658 );
    and g6756 ( n11016 , n3442 , n2191 );
    not g6757 ( n9268 , n9732 );
    nor g6758 ( n13131 , n833 , n12706 );
    xor g6759 ( n9515 , n841 , n6734 );
    or g6760 ( n11329 , n4022 , n206 );
    not g6761 ( n5947 , n8860 );
    not g6762 ( n3387 , n7436 );
    xnor g6763 ( n8750 , n12979 , n12589 );
    xnor g6764 ( n7097 , n8548 , n2107 );
    xnor g6765 ( n1801 , n3436 , n1157 );
    nor g6766 ( n4050 , n9629 , n6253 );
    and g6767 ( n2020 , n9158 , n6902 );
    and g6768 ( n129 , n7987 , n12556 );
    or g6769 ( n10698 , n12009 , n4947 );
    not g6770 ( n11545 , n3361 );
    xnor g6771 ( n6603 , n6654 , n5180 );
    or g6772 ( n9826 , n4620 , n6265 );
    xor g6773 ( n183 , n11473 , n2047 );
    or g6774 ( n6065 , n6332 , n2675 );
    xnor g6775 ( n8394 , n7822 , n9603 );
    or g6776 ( n8350 , n1816 , n10367 );
    not g6777 ( n6308 , n9394 );
    or g6778 ( n11630 , n11134 , n816 );
    xnor g6779 ( n5106 , n9859 , n5830 );
    and g6780 ( n12134 , n2330 , n7320 );
    xnor g6781 ( n6867 , n3289 , n8765 );
    or g6782 ( n329 , n10877 , n2675 );
    nor g6783 ( n5819 , n6647 , n6052 );
    xnor g6784 ( n7851 , n5273 , n8379 );
    or g6785 ( n8286 , n12264 , n12355 );
    nor g6786 ( n13130 , n11002 , n3930 );
    and g6787 ( n6473 , n4914 , n9624 );
    not g6788 ( n2689 , n2498 );
    and g6789 ( n4172 , n5597 , n5846 );
    xnor g6790 ( n12094 , n4554 , n8927 );
    xnor g6791 ( n9547 , n3404 , n7704 );
    xnor g6792 ( n4935 , n8737 , n1244 );
    not g6793 ( n11230 , n8616 );
    not g6794 ( n12159 , n12605 );
    and g6795 ( n990 , n6493 , n6517 );
    xnor g6796 ( n9779 , n2081 , n9681 );
    and g6797 ( n10531 , n3393 , n6812 );
    xnor g6798 ( n7365 , n1821 , n8298 );
    or g6799 ( n636 , n7900 , n4640 );
    not g6800 ( n13226 , n10733 );
    or g6801 ( n3596 , n7133 , n1043 );
    xnor g6802 ( n3607 , n6413 , n12562 );
    nor g6803 ( n360 , n10204 , n3876 );
    or g6804 ( n7179 , n11801 , n1901 );
    xnor g6805 ( n6736 , n5071 , n1133 );
    and g6806 ( n1742 , n6950 , n10002 );
    and g6807 ( n8150 , n9617 , n10359 );
    xnor g6808 ( n6516 , n9833 , n9544 );
    xnor g6809 ( n221 , n10745 , n5457 );
    not g6810 ( n11007 , n834 );
    xnor g6811 ( n11246 , n3308 , n2349 );
    and g6812 ( n2746 , n12911 , n2792 );
    not g6813 ( n11729 , n2737 );
    xnor g6814 ( n5928 , n4451 , n2308 );
    and g6815 ( n12963 , n8573 , n6753 );
    or g6816 ( n8785 , n11933 , n206 );
    not g6817 ( n9739 , n11734 );
    xnor g6818 ( n10614 , n5319 , n12005 );
    and g6819 ( n12379 , n9848 , n7807 );
    or g6820 ( n6236 , n691 , n2941 );
    not g6821 ( n11113 , n12065 );
    xnor g6822 ( n3086 , n4874 , n7692 );
    and g6823 ( n770 , n8905 , n12625 );
    nor g6824 ( n11964 , n12083 , n2478 );
    xnor g6825 ( n11585 , n3668 , n6560 );
    xnor g6826 ( n8087 , n8170 , n662 );
    and g6827 ( n3287 , n6187 , n4072 );
    nor g6828 ( n3308 , n8025 , n9865 );
    xnor g6829 ( n2519 , n7558 , n5682 );
    not g6830 ( n12625 , n9903 );
    not g6831 ( n11751 , n8768 );
    xnor g6832 ( n10952 , n12440 , n1541 );
    or g6833 ( n12708 , n9728 , n11555 );
    xnor g6834 ( n10307 , n6479 , n5315 );
    xnor g6835 ( n6570 , n5660 , n10562 );
    nor g6836 ( n9047 , n8914 , n7296 );
    or g6837 ( n6912 , n11168 , n590 );
    nor g6838 ( n9314 , n2294 , n12228 );
    not g6839 ( n7460 , n8031 );
    not g6840 ( n6469 , n4217 );
    and g6841 ( n7760 , n3492 , n8286 );
    xnor g6842 ( n5858 , n1534 , n3292 );
    or g6843 ( n10888 , n5086 , n12814 );
    not g6844 ( n9934 , n11634 );
    xnor g6845 ( n2488 , n9571 , n12149 );
    or g6846 ( n2947 , n10166 , n6497 );
    not g6847 ( n2404 , n1929 );
    or g6848 ( n10993 , n154 , n776 );
    or g6849 ( n3507 , n4880 , n10659 );
    and g6850 ( n10015 , n9353 , n834 );
    or g6851 ( n5893 , n8660 , n2938 );
    and g6852 ( n3144 , n10392 , n9655 );
    and g6853 ( n6317 , n1931 , n4666 );
    not g6854 ( n343 , n504 );
    nor g6855 ( n718 , n2307 , n9258 );
    nor g6856 ( n10130 , n3973 , n11185 );
    not g6857 ( n3565 , n7288 );
    xnor g6858 ( n1177 , n9050 , n10080 );
    or g6859 ( n7869 , n4944 , n12298 );
    or g6860 ( n3193 , n9632 , n8268 );
    or g6861 ( n4963 , n618 , n9858 );
    nor g6862 ( n8706 , n6072 , n10840 );
    xnor g6863 ( n10076 , n12699 , n11363 );
    and g6864 ( n4896 , n6578 , n6712 );
    and g6865 ( n7982 , n4527 , n9067 );
    not g6866 ( n448 , n13003 );
    xnor g6867 ( n5188 , n5574 , n5764 );
    and g6868 ( n12978 , n12283 , n11543 );
    nor g6869 ( n9423 , n10568 , n12520 );
    xnor g6870 ( n2467 , n3367 , n3938 );
    and g6871 ( n1756 , n4129 , n11862 );
    not g6872 ( n4149 , n397 );
    xnor g6873 ( n7841 , n498 , n9459 );
    nor g6874 ( n11214 , n1942 , n2115 );
    xnor g6875 ( n11050 , n7214 , n1237 );
    or g6876 ( n778 , n13036 , n4640 );
    not g6877 ( n3674 , n3411 );
    or g6878 ( n6510 , n7798 , n8268 );
    nor g6879 ( n11167 , n865 , n8055 );
    not g6880 ( n7780 , n10594 );
    or g6881 ( n8961 , n3660 , n8958 );
    xor g6882 ( n4591 , n9313 , n764 );
    or g6883 ( n8073 , n2913 , n12654 );
    nor g6884 ( n6010 , n12809 , n12066 );
    or g6885 ( n6640 , n4625 , n9331 );
    or g6886 ( n3620 , n8471 , n6688 );
    and g6887 ( n342 , n3163 , n286 );
    xnor g6888 ( n86 , n11831 , n10647 );
    xnor g6889 ( n426 , n4986 , n4626 );
    nor g6890 ( n3246 , n624 , n12752 );
    xnor g6891 ( n3074 , n9614 , n1581 );
    not g6892 ( n12145 , n11335 );
    xnor g6893 ( n12480 , n4309 , n8999 );
    and g6894 ( n997 , n4382 , n1724 );
    xnor g6895 ( n11412 , n1096 , n5575 );
    xnor g6896 ( n1304 , n11917 , n1339 );
    and g6897 ( n6344 , n10511 , n3360 );
    not g6898 ( n12243 , n9315 );
    or g6899 ( n3040 , n6056 , n9492 );
    nor g6900 ( n1454 , n1921 , n933 );
    xnor g6901 ( n2188 , n1340 , n9840 );
    or g6902 ( n6468 , n9228 , n12273 );
    and g6903 ( n12089 , n1842 , n6697 );
    and g6904 ( n9984 , n9659 , n395 );
    or g6905 ( n10640 , n10021 , n2222 );
    not g6906 ( n4058 , n8467 );
    not g6907 ( n204 , n9762 );
    or g6908 ( n8085 , n1089 , n8143 );
    xnor g6909 ( n5326 , n3571 , n3517 );
    or g6910 ( n8802 , n63 , n2544 );
    nor g6911 ( n13107 , n13008 , n4637 );
    or g6912 ( n12879 , n185 , n4431 );
    and g6913 ( n8795 , n7162 , n7769 );
    xnor g6914 ( n6415 , n7157 , n9742 );
    and g6915 ( n3433 , n5188 , n9637 );
    not g6916 ( n6171 , n7829 );
    or g6917 ( n7098 , n3643 , n6544 );
    or g6918 ( n4173 , n868 , n8269 );
    nor g6919 ( n4641 , n10762 , n1675 );
    or g6920 ( n12658 , n2606 , n11422 );
    not g6921 ( n11965 , n5320 );
    not g6922 ( n9444 , n6392 );
    or g6923 ( n7934 , n3460 , n6635 );
    or g6924 ( n12124 , n7074 , n5242 );
    not g6925 ( n11054 , n4006 );
    or g6926 ( n1050 , n13090 , n12415 );
    or g6927 ( n3415 , n3142 , n2320 );
    or g6928 ( n6503 , n7825 , n10029 );
    xnor g6929 ( n2992 , n13056 , n3021 );
    nor g6930 ( n10246 , n7712 , n7389 );
    xnor g6931 ( n13151 , n2602 , n13147 );
    or g6932 ( n4804 , n2854 , n2853 );
    not g6933 ( n3726 , n9887 );
    and g6934 ( n3831 , n9216 , n5920 );
    or g6935 ( n4634 , n8671 , n5796 );
    not g6936 ( n12663 , n8923 );
    not g6937 ( n4209 , n287 );
    xnor g6938 ( n624 , n12267 , n9495 );
    xor g6939 ( n12602 , n9061 , n5876 );
    or g6940 ( n8252 , n6958 , n12360 );
    and g6941 ( n5223 , n6634 , n7547 );
    and g6942 ( n194 , n1413 , n9398 );
    or g6943 ( n6576 , n4814 , n8584 );
    xnor g6944 ( n12937 , n5752 , n12827 );
    and g6945 ( n4392 , n168 , n1245 );
    nor g6946 ( n12396 , n4788 , n8122 );
    nor g6947 ( n10604 , n656 , n9514 );
    and g6948 ( n486 , n9653 , n1979 );
    not g6949 ( n1370 , n11734 );
    or g6950 ( n12921 , n354 , n12934 );
    and g6951 ( n4636 , n809 , n7404 );
    xnor g6952 ( n1939 , n10351 , n1788 );
    or g6953 ( n5687 , n9010 , n121 );
    xnor g6954 ( n7563 , n12774 , n6228 );
    or g6955 ( n5579 , n12124 , n7437 );
    xnor g6956 ( n5116 , n2665 , n7992 );
    xnor g6957 ( n4615 , n4102 , n8528 );
    and g6958 ( n8104 , n12419 , n790 );
    or g6959 ( n6198 , n1191 , n2544 );
    xnor g6960 ( n2426 , n4279 , n7348 );
    or g6961 ( n12558 , n3428 , n4230 );
    and g6962 ( n10254 , n5310 , n5630 );
    or g6963 ( n2353 , n186 , n7551 );
    and g6964 ( n316 , n7529 , n5729 );
    or g6965 ( n9133 , n2692 , n5242 );
    or g6966 ( n3330 , n13013 , n4454 );
    and g6967 ( n4474 , n7973 , n4963 );
    not g6968 ( n8578 , n1423 );
    xnor g6969 ( n3704 , n12756 , n9408 );
    xnor g6970 ( n12015 , n9927 , n10493 );
    xnor g6971 ( n8908 , n4025 , n11886 );
    xnor g6972 ( n5104 , n11445 , n3055 );
    not g6973 ( n6770 , n10408 );
    xnor g6974 ( n11855 , n2831 , n5826 );
    or g6975 ( n10571 , n11680 , n9195 );
    or g6976 ( n3688 , n2630 , n561 );
    and g6977 ( n11860 , n289 , n7934 );
    or g6978 ( n2634 , n2950 , n5945 );
    not g6979 ( n12086 , n5659 );
    not g6980 ( n6327 , n10105 );
    not g6981 ( n6186 , n9058 );
    xor g6982 ( n887 , n5731 , n2314 );
    and g6983 ( n3202 , n7253 , n8531 );
    or g6984 ( n9468 , n8575 , n12423 );
    or g6985 ( n9424 , n4778 , n11491 );
    or g6986 ( n5118 , n10202 , n8226 );
    not g6987 ( n3703 , n10642 );
    not g6988 ( n9885 , n2350 );
    xnor g6989 ( n2926 , n383 , n3177 );
    xnor g6990 ( n1600 , n2812 , n3207 );
    xnor g6991 ( n4291 , n5365 , n4892 );
    and g6992 ( n6390 , n636 , n9365 );
    or g6993 ( n1575 , n11114 , n1012 );
    not g6994 ( n4686 , n8139 );
    xnor g6995 ( n5486 , n1079 , n1616 );
    or g6996 ( n2950 , n10188 , n2958 );
    or g6997 ( n912 , n5430 , n9075 );
    and g6998 ( n3526 , n7130 , n5489 );
    xnor g6999 ( n2235 , n1543 , n426 );
    not g7000 ( n11152 , n2590 );
    nor g7001 ( n10579 , n7635 , n12087 );
    or g7002 ( n12445 , n10588 , n9744 );
    or g7003 ( n10668 , n10253 , n6703 );
    xnor g7004 ( n5254 , n6588 , n1115 );
    nor g7005 ( n8773 , n10069 , n5419 );
    xnor g7006 ( n10238 , n4837 , n8013 );
    and g7007 ( n9952 , n9552 , n5608 );
    and g7008 ( n7100 , n4377 , n10633 );
    nor g7009 ( n9393 , n4952 , n1133 );
    xnor g7010 ( n7189 , n8300 , n148 );
    xnor g7011 ( n1479 , n891 , n2082 );
    nor g7012 ( n9278 , n5879 , n13176 );
    or g7013 ( n3597 , n1571 , n1026 );
    xnor g7014 ( n9357 , n4306 , n4362 );
    xnor g7015 ( n2931 , n10984 , n9547 );
    nor g7016 ( n3882 , n4035 , n3912 );
    or g7017 ( n12646 , n1230 , n9699 );
    and g7018 ( n12575 , n5272 , n5194 );
    or g7019 ( n7412 , n8472 , n8563 );
    xnor g7020 ( n10297 , n11603 , n12776 );
    not g7021 ( n10535 , n7479 );
    and g7022 ( n8123 , n1912 , n12263 );
    and g7023 ( n10667 , n7410 , n8070 );
    xnor g7024 ( n12278 , n4233 , n8966 );
    buf g7025 ( n177 , n6210 );
    or g7026 ( n6363 , n4221 , n6769 );
    not g7027 ( n7135 , n10594 );
    xnor g7028 ( n12056 , n3444 , n838 );
    not g7029 ( n9162 , n8332 );
    and g7030 ( n4411 , n11701 , n11194 );
    nor g7031 ( n9456 , n382 , n3967 );
    or g7032 ( n8808 , n7680 , n12818 );
    or g7033 ( n993 , n3195 , n10470 );
    xnor g7034 ( n12669 , n11550 , n2458 );
    xnor g7035 ( n10080 , n1765 , n8393 );
    nor g7036 ( n1381 , n10148 , n8232 );
    or g7037 ( n3661 , n11080 , n10155 );
    xnor g7038 ( n2340 , n10609 , n13126 );
    or g7039 ( n9403 , n5853 , n5658 );
    or g7040 ( n2238 , n7672 , n7221 );
    xnor g7041 ( n6256 , n6951 , n3018 );
    or g7042 ( n9964 , n9700 , n4652 );
    or g7043 ( n4573 , n2504 , n2276 );
    not g7044 ( n6726 , n8859 );
    or g7045 ( n11937 , n3516 , n559 );
    not g7046 ( n8024 , n1364 );
    nor g7047 ( n3471 , n778 , n10704 );
    or g7048 ( n5039 , n11018 , n9159 );
    xnor g7049 ( n9425 , n13171 , n5555 );
    not g7050 ( n205 , n6484 );
    not g7051 ( n1652 , n2000 );
    not g7052 ( n11697 , n3352 );
    or g7053 ( n2225 , n8729 , n9159 );
    xnor g7054 ( n2336 , n6191 , n1894 );
    not g7055 ( n2412 , n9924 );
    not g7056 ( n3194 , n11709 );
    not g7057 ( n11323 , n13172 );
    or g7058 ( n599 , n9676 , n5817 );
    or g7059 ( n10184 , n10616 , n11578 );
    and g7060 ( n5984 , n4756 , n2901 );
    and g7061 ( n4728 , n6260 , n2918 );
    xnor g7062 ( n3088 , n11030 , n11488 );
    xnor g7063 ( n7437 , n6283 , n12779 );
    and g7064 ( n2053 , n5348 , n6523 );
    not g7065 ( n334 , n401 );
    xnor g7066 ( n2476 , n5649 , n1685 );
    nor g7067 ( n11520 , n7197 , n4447 );
    and g7068 ( n1465 , n10975 , n6352 );
    and g7069 ( n5432 , n5988 , n6992 );
    not g7070 ( n9809 , n12276 );
    not g7071 ( n12837 , n12482 );
    and g7072 ( n6286 , n10719 , n9454 );
    xnor g7073 ( n2724 , n7360 , n10818 );
    xnor g7074 ( n8942 , n7823 , n9875 );
    and g7075 ( n481 , n13066 , n4468 );
    and g7076 ( n11885 , n6772 , n8574 );
    xnor g7077 ( n6691 , n9391 , n9057 );
    xnor g7078 ( n10889 , n5816 , n6642 );
    nor g7079 ( n6799 , n12008 , n1863 );
    or g7080 ( n7650 , n10334 , n11668 );
    nor g7081 ( n8429 , n5599 , n6613 );
    xnor g7082 ( n3953 , n6114 , n4839 );
    not g7083 ( n3940 , n12651 );
    xnor g7084 ( n8328 , n12627 , n7079 );
    nor g7085 ( n10387 , n259 , n12138 );
    or g7086 ( n7949 , n2140 , n620 );
    xnor g7087 ( n1764 , n11684 , n2309 );
    and g7088 ( n1528 , n5214 , n3409 );
    xnor g7089 ( n5935 , n3013 , n11410 );
    or g7090 ( n281 , n9969 , n7732 );
    xnor g7091 ( n5396 , n3475 , n11932 );
    and g7092 ( n9549 , n11646 , n9976 );
    and g7093 ( n8034 , n9288 , n10006 );
    or g7094 ( n2310 , n2669 , n6635 );
    not g7095 ( n9017 , n11222 );
    or g7096 ( n4619 , n12926 , n8341 );
    xnor g7097 ( n6116 , n11059 , n13091 );
    and g7098 ( n3782 , n10241 , n10959 );
    xnor g7099 ( n5605 , n6518 , n557 );
    and g7100 ( n6589 , n5531 , n5602 );
    xnor g7101 ( n5329 , n3159 , n12507 );
    or g7102 ( n3241 , n9465 , n9772 );
    and g7103 ( n7252 , n8560 , n6365 );
    not g7104 ( n9712 , n3850 );
    not g7105 ( n1544 , n6570 );
    not g7106 ( n11157 , n7411 );
    or g7107 ( n8531 , n5095 , n2205 );
    xnor g7108 ( n9836 , n2485 , n12752 );
    or g7109 ( n11821 , n7446 , n5223 );
    not g7110 ( n7636 , n1384 );
    or g7111 ( n3316 , n481 , n10899 );
    and g7112 ( n708 , n6238 , n2137 );
    and g7113 ( n12424 , n4964 , n2339 );
    xnor g7114 ( n10853 , n9965 , n10831 );
    not g7115 ( n3598 , n12853 );
    xnor g7116 ( n4369 , n11401 , n6899 );
    or g7117 ( n11241 , n3496 , n6966 );
    or g7118 ( n10837 , n7809 , n13232 );
    not g7119 ( n5245 , n11064 );
    xnor g7120 ( n7265 , n9530 , n13057 );
    and g7121 ( n6903 , n4901 , n6403 );
    or g7122 ( n7229 , n7608 , n6404 );
    xnor g7123 ( n1581 , n9315 , n4399 );
    not g7124 ( n11171 , n1916 );
    or g7125 ( n8112 , n2942 , n1618 );
    not g7126 ( n3036 , n6075 );
    or g7127 ( n7625 , n1490 , n4904 );
    and g7128 ( n4658 , n3461 , n6259 );
    or g7129 ( n1878 , n7193 , n9933 );
    or g7130 ( n7810 , n12476 , n5184 );
    and g7131 ( n9270 , n4488 , n3036 );
    xnor g7132 ( n7673 , n3368 , n7576 );
    or g7133 ( n8479 , n8108 , n8702 );
    nor g7134 ( n5349 , n7326 , n3565 );
    xnor g7135 ( n6500 , n10423 , n3276 );
    or g7136 ( n9555 , n8849 , n5414 );
    xnor g7137 ( n6043 , n2482 , n10113 );
    or g7138 ( n7758 , n7133 , n12847 );
    xor g7139 ( n10733 , n10751 , n1032 );
    or g7140 ( n6649 , n2017 , n7692 );
    xnor g7141 ( n8725 , n11417 , n11019 );
    nor g7142 ( n961 , n10811 , n836 );
    or g7143 ( n1705 , n2144 , n12421 );
    and g7144 ( n11199 , n6308 , n6925 );
    xnor g7145 ( n4747 , n2516 , n5728 );
    or g7146 ( n6430 , n4355 , n8933 );
    and g7147 ( n74 , n2724 , n6455 );
    xnor g7148 ( n12283 , n10697 , n2366 );
    not g7149 ( n8898 , n1812 );
    and g7150 ( n8092 , n7450 , n7867 );
    or g7151 ( n7315 , n7409 , n2714 );
    not g7152 ( n11244 , n13058 );
    xnor g7153 ( n7030 , n3637 , n12047 );
    and g7154 ( n7224 , n6566 , n155 );
    not g7155 ( n3752 , n2392 );
    and g7156 ( n3502 , n4033 , n1503 );
    and g7157 ( n5292 , n3250 , n4117 );
    or g7158 ( n9477 , n4946 , n4139 );
    xnor g7159 ( n8633 , n11970 , n2502 );
    and g7160 ( n7648 , n9049 , n2827 );
    or g7161 ( n5572 , n12563 , n10029 );
    xnor g7162 ( n10205 , n28 , n253 );
    and g7163 ( n2955 , n6624 , n7575 );
    or g7164 ( n1413 , n6787 , n4669 );
    or g7165 ( n3656 , n3270 , n13143 );
    not g7166 ( n10057 , n5962 );
    not g7167 ( n10552 , n6668 );
    or g7168 ( n5704 , n1887 , n1043 );
    nor g7169 ( n2050 , n5798 , n9276 );
    xnor g7170 ( n5643 , n4781 , n8633 );
    not g7171 ( n9421 , n11574 );
    or g7172 ( n11363 , n161 , n10179 );
    not g7173 ( n4620 , n2295 );
    xnor g7174 ( n4705 , n5759 , n12038 );
    xnor g7175 ( n2584 , n2125 , n10118 );
    nor g7176 ( n7169 , n11530 , n4472 );
    and g7177 ( n9048 , n3545 , n13140 );
    and g7178 ( n4219 , n7055 , n6292 );
    or g7179 ( n4363 , n994 , n1433 );
    xnor g7180 ( n7808 , n6199 , n3147 );
    xnor g7181 ( n1758 , n4531 , n6077 );
    nor g7182 ( n3686 , n12468 , n2202 );
    and g7183 ( n9414 , n308 , n4302 );
    or g7184 ( n310 , n8392 , n8030 );
    xor g7185 ( n8919 , n8887 , n5270 );
    xnor g7186 ( n6698 , n1549 , n12611 );
    not g7187 ( n12563 , n12306 );
    or g7188 ( n2337 , n8335 , n6265 );
    not g7189 ( n1377 , n10424 );
    and g7190 ( n8903 , n12776 , n11603 );
    or g7191 ( n13119 , n318 , n10106 );
    not g7192 ( n9723 , n7659 );
    or g7193 ( n10225 , n9112 , n4947 );
    or g7194 ( n4045 , n1995 , n1081 );
    xnor g7195 ( n2073 , n9389 , n9551 );
    not g7196 ( n7950 , n9915 );
    xnor g7197 ( n8121 , n9436 , n3674 );
    xnor g7198 ( n11970 , n494 , n11329 );
    xnor g7199 ( n7838 , n7294 , n10111 );
    xnor g7200 ( n2828 , n10424 , n13076 );
    not g7201 ( n11800 , n3838 );
    and g7202 ( n5061 , n7523 , n7975 );
    not g7203 ( n1186 , n8227 );
    not g7204 ( n1725 , n6409 );
    or g7205 ( n12137 , n7372 , n11628 );
    xnor g7206 ( n6908 , n1313 , n3667 );
    and g7207 ( n5732 , n7529 , n10451 );
    or g7208 ( n5160 , n7283 , n7723 );
    and g7209 ( n10040 , n3987 , n12362 );
    or g7210 ( n3871 , n6975 , n7871 );
    or g7211 ( n160 , n9934 , n2675 );
    and g7212 ( n9247 , n2715 , n4265 );
    and g7213 ( n5024 , n4729 , n3204 );
    not g7214 ( n1255 , n2202 );
    xnor g7215 ( n7781 , n4337 , n10478 );
    xnor g7216 ( n7958 , n12716 , n9322 );
    xnor g7217 ( n4302 , n1849 , n5594 );
    xnor g7218 ( n10506 , n3741 , n9143 );
    not g7219 ( n3589 , n589 );
    xnor g7220 ( n6094 , n11561 , n8578 );
    xnor g7221 ( n1519 , n4356 , n10499 );
    or g7222 ( n6855 , n8400 , n13148 );
    not g7223 ( n930 , n12577 );
    or g7224 ( n2610 , n9945 , n2418 );
    or g7225 ( n9937 , n9892 , n10526 );
    or g7226 ( n12030 , n3259 , n80 );
    not g7227 ( n9465 , n4507 );
    not g7228 ( n1045 , n12443 );
    xnor g7229 ( n5756 , n10341 , n3636 );
    not g7230 ( n3516 , n3311 );
    nor g7231 ( n11916 , n3728 , n8537 );
    or g7232 ( n8250 , n12055 , n1285 );
    and g7233 ( n8763 , n12737 , n5956 );
    not g7234 ( n8658 , n13184 );
    not g7235 ( n2406 , n2458 );
    not g7236 ( n6543 , n12641 );
    and g7237 ( n4561 , n7924 , n2528 );
    and g7238 ( n4941 , n2412 , n5668 );
    and g7239 ( n5303 , n6690 , n12772 );
    xnor g7240 ( n7613 , n2514 , n13160 );
    or g7241 ( n4738 , n74 , n9278 );
    xor g7242 ( n12916 , n424 , n1698 );
    or g7243 ( n2509 , n8008 , n12113 );
    xnor g7244 ( n396 , n9292 , n11921 );
    xnor g7245 ( n3055 , n6446 , n4178 );
    or g7246 ( n52 , n6849 , n12526 );
    xnor g7247 ( n456 , n1546 , n2204 );
    not g7248 ( n11808 , n11324 );
    and g7249 ( n8826 , n2648 , n9829 );
    or g7250 ( n7192 , n5040 , n6370 );
    nor g7251 ( n3884 , n1676 , n10083 );
    and g7252 ( n7855 , n4595 , n11343 );
    and g7253 ( n1515 , n12139 , n11775 );
    xnor g7254 ( n2937 , n4175 , n3231 );
    or g7255 ( n197 , n10290 , n11668 );
    and g7256 ( n5815 , n8093 , n7019 );
    nor g7257 ( n10600 , n145 , n853 );
    nor g7258 ( n11265 , n12642 , n3291 );
    xnor g7259 ( n8287 , n4713 , n11441 );
    or g7260 ( n13178 , n11626 , n2891 );
    nor g7261 ( n3219 , n11488 , n1982 );
    and g7262 ( n3997 , n724 , n11163 );
    xnor g7263 ( n8195 , n7874 , n5922 );
    xnor g7264 ( n8484 , n12610 , n13067 );
    nor g7265 ( n367 , n5556 , n13198 );
    or g7266 ( n9918 , n1320 , n2671 );
    or g7267 ( n5365 , n5423 , n2133 );
    or g7268 ( n12058 , n4622 , n11214 );
    not g7269 ( n6595 , n13060 );
    or g7270 ( n2177 , n1883 , n6732 );
    and g7271 ( n8560 , n1522 , n3483 );
    or g7272 ( n2922 , n6035 , n11146 );
    or g7273 ( n747 , n626 , n7887 );
    xnor g7274 ( n2813 , n1256 , n1619 );
    and g7275 ( n3973 , n2198 , n193 );
    and g7276 ( n11712 , n11690 , n12743 );
    xnor g7277 ( n2439 , n1803 , n7587 );
    or g7278 ( n8901 , n11320 , n6293 );
    and g7279 ( n2335 , n2747 , n8762 );
    xnor g7280 ( n3863 , n9371 , n8323 );
    and g7281 ( n3251 , n9828 , n10804 );
    nor g7282 ( n5221 , n4968 , n11700 );
    xnor g7283 ( n11603 , n2513 , n11578 );
    xnor g7284 ( n13020 , n3878 , n7248 );
    xnor g7285 ( n10217 , n5407 , n2708 );
    buf g7286 ( n1144 , n8569 );
    nor g7287 ( n449 , n3764 , n2888 );
    nor g7288 ( n12587 , n232 , n3580 );
    or g7289 ( n6240 , n683 , n4144 );
    xnor g7290 ( n7148 , n13193 , n2642 );
    or g7291 ( n12530 , n154 , n9962 );
    xnor g7292 ( n7121 , n6184 , n2115 );
    not g7293 ( n11986 , n12417 );
    and g7294 ( n9242 , n1582 , n5706 );
    or g7295 ( n9535 , n660 , n1530 );
    xnor g7296 ( n1141 , n880 , n2856 );
    xnor g7297 ( n6809 , n11518 , n10337 );
    xnor g7298 ( n441 , n12737 , n10009 );
    or g7299 ( n8699 , n6726 , n206 );
    or g7300 ( n7174 , n9094 , n6605 );
    xnor g7301 ( n8921 , n565 , n10445 );
    and g7302 ( n10362 , n1539 , n12633 );
    or g7303 ( n13062 , n1296 , n8702 );
    xnor g7304 ( n3904 , n1461 , n2303 );
    and g7305 ( n5834 , n2482 , n12289 );
    not g7306 ( n1337 , n11254 );
    nor g7307 ( n3080 , n6805 , n7691 );
    nor g7308 ( n10270 , n1744 , n315 );
    xnor g7309 ( n6984 , n10134 , n183 );
    not g7310 ( n2329 , n7974 );
    or g7311 ( n3767 , n11291 , n7530 );
    and g7312 ( n1326 , n3473 , n8337 );
    nor g7313 ( n1287 , n5402 , n5149 );
    or g7314 ( n11877 , n10263 , n12695 );
    or g7315 ( n12712 , n5365 , n8749 );
    not g7316 ( n1538 , n12418 );
    or g7317 ( n8127 , n5667 , n5242 );
    not g7318 ( n2118 , n12408 );
    xnor g7319 ( n13143 , n10409 , n741 );
    or g7320 ( n8047 , n9450 , n6968 );
    and g7321 ( n9092 , n2458 , n9669 );
    nor g7322 ( n9208 , n5702 , n7866 );
    not g7323 ( n5697 , n13098 );
    not g7324 ( n3870 , n825 );
    not g7325 ( n1741 , n10606 );
    or g7326 ( n2204 , n7158 , n2059 );
    not g7327 ( n8863 , n3409 );
    and g7328 ( n10004 , n4964 , n11222 );
    xnor g7329 ( n10971 , n12812 , n2983 );
    and g7330 ( n10191 , n545 , n1849 );
    and g7331 ( n5237 , n5118 , n6806 );
    xnor g7332 ( n2120 , n2807 , n10355 );
    nor g7333 ( n11843 , n11673 , n42 );
    and g7334 ( n1987 , n7869 , n3606 );
    or g7335 ( n3310 , n10871 , n1463 );
    not g7336 ( n6178 , n11537 );
    and g7337 ( n4427 , n4708 , n12550 );
    and g7338 ( n394 , n12902 , n1684 );
    and g7339 ( n4001 , n433 , n9224 );
    xnor g7340 ( n2665 , n10483 , n6782 );
    or g7341 ( n7680 , n10143 , n12847 );
    and g7342 ( n336 , n93 , n7772 );
    and g7343 ( n11439 , n6164 , n413 );
    and g7344 ( n12760 , n1030 , n4243 );
    or g7345 ( n5366 , n5926 , n10884 );
    and g7346 ( n12341 , n11985 , n5435 );
    nor g7347 ( n13111 , n6179 , n5674 );
    or g7348 ( n8292 , n11548 , n9159 );
    or g7349 ( n11795 , n6010 , n11746 );
    and g7350 ( n5262 , n9646 , n12984 );
    xnor g7351 ( n10663 , n10053 , n12087 );
    xnor g7352 ( n8678 , n5114 , n3506 );
    or g7353 ( n9995 , n6498 , n258 );
    or g7354 ( n4648 , n10290 , n6265 );
    xnor g7355 ( n5951 , n5935 , n8181 );
    xnor g7356 ( n54 , n5438 , n5070 );
    or g7357 ( n4903 , n12397 , n5235 );
    or g7358 ( n703 , n10990 , n13032 );
    xnor g7359 ( n12215 , n3296 , n5458 );
    nor g7360 ( n13150 , n10163 , n4344 );
    and g7361 ( n13121 , n855 , n2047 );
    and g7362 ( n11652 , n8940 , n5536 );
    not g7363 ( n10384 , n9895 );
    not g7364 ( n9282 , n8139 );
    not g7365 ( n5650 , n5302 );
    nor g7366 ( n10515 , n149 , n8152 );
    and g7367 ( n10703 , n5270 , n5383 );
    and g7368 ( n7144 , n4848 , n4984 );
    not g7369 ( n3450 , n6700 );
    and g7370 ( n4799 , n4114 , n8506 );
    not g7371 ( n8907 , n9610 );
    and g7372 ( n2583 , n12592 , n3085 );
    xnor g7373 ( n9090 , n2630 , n2561 );
    nor g7374 ( n13019 , n10048 , n12842 );
    and g7375 ( n7761 , n8183 , n9475 );
    and g7376 ( n1917 , n3998 , n4486 );
    or g7377 ( n7561 , n4411 , n11135 );
    nor g7378 ( n969 , n3263 , n12045 );
    xnor g7379 ( n529 , n4264 , n6287 );
    or g7380 ( n132 , n9567 , n7429 );
    not g7381 ( n7074 , n469 );
    or g7382 ( n4929 , n9553 , n6278 );
    xnor g7383 ( n444 , n11433 , n12214 );
    not g7384 ( n12490 , n9475 );
    nor g7385 ( n7520 , n6800 , n13236 );
    not g7386 ( n2614 , n1302 );
    or g7387 ( n4976 , n9181 , n5740 );
    or g7388 ( n7012 , n5890 , n2133 );
    nor g7389 ( n3491 , n13094 , n8218 );
    and g7390 ( n13040 , n4618 , n1232 );
    and g7391 ( n6080 , n6421 , n13088 );
    not g7392 ( n4412 , n1753 );
    or g7393 ( n12788 , n12855 , n9088 );
    or g7394 ( n4321 , n2877 , n7903 );
    and g7395 ( n4047 , n3342 , n8606 );
    not g7396 ( n6488 , n3076 );
    nor g7397 ( n10990 , n2431 , n10178 );
    and g7398 ( n972 , n12043 , n1005 );
    or g7399 ( n8244 , n189 , n11929 );
    or g7400 ( n5210 , n1331 , n4455 );
    xnor g7401 ( n5211 , n4021 , n6863 );
    or g7402 ( n3172 , n11582 , n3801 );
    and g7403 ( n10651 , n233 , n11539 );
    xnor g7404 ( n4011 , n7277 , n5378 );
    or g7405 ( n4942 , n5377 , n12491 );
    xnor g7406 ( n6288 , n1092 , n1479 );
    xnor g7407 ( n4601 , n10802 , n10684 );
    or g7408 ( n1933 , n8532 , n12273 );
    nor g7409 ( n185 , n6264 , n11458 );
    nor g7410 ( n12111 , n2063 , n12586 );
    or g7411 ( n4784 , n2130 , n8465 );
    or g7412 ( n2802 , n6768 , n9195 );
    or g7413 ( n3444 , n7228 , n1383 );
    nor g7414 ( n8364 , n6765 , n10744 );
    xnor g7415 ( n378 , n12374 , n12322 );
    xnor g7416 ( n7399 , n11763 , n8021 );
    not g7417 ( n7388 , n6417 );
    and g7418 ( n10417 , n10708 , n9588 );
    not g7419 ( n9606 , n4748 );
    nor g7420 ( n8513 , n6902 , n9158 );
    not g7421 ( n7817 , n720 );
    or g7422 ( n6335 , n5897 , n159 );
    not g7423 ( n1082 , n12564 );
    nor g7424 ( n5392 , n2334 , n3468 );
    not g7425 ( n4139 , n5753 );
    xnor g7426 ( n6785 , n3951 , n5896 );
    xnor g7427 ( n12319 , n4369 , n9805 );
    not g7428 ( n9992 , n1521 );
    not g7429 ( n6846 , n12482 );
    or g7430 ( n3284 , n10761 , n12388 );
    not g7431 ( n3890 , n9620 );
    nor g7432 ( n10308 , n12230 , n4204 );
    or g7433 ( n6146 , n1359 , n2438 );
    xnor g7434 ( n9792 , n2011 , n9483 );
    nor g7435 ( n4386 , n6097 , n11416 );
    xnor g7436 ( n11454 , n10500 , n6542 );
    or g7437 ( n505 , n5107 , n1571 );
    and g7438 ( n2631 , n7011 , n7117 );
    not g7439 ( n10916 , n3395 );
    not g7440 ( n12478 , n4318 );
    and g7441 ( n7240 , n10948 , n9137 );
    xnor g7442 ( n9081 , n6242 , n10276 );
    not g7443 ( n7075 , n6168 );
    or g7444 ( n5212 , n3159 , n9507 );
    or g7445 ( n9892 , n12748 , n12188 );
    or g7446 ( n3750 , n6172 , n7610 );
    not g7447 ( n11122 , n7720 );
    xnor g7448 ( n10073 , n5299 , n13072 );
    and g7449 ( n9115 , n3435 , n11697 );
    and g7450 ( n13139 , n8835 , n8521 );
    or g7451 ( n978 , n652 , n5076 );
    not g7452 ( n8936 , n28 );
    xnor g7453 ( n363 , n1675 , n4573 );
    or g7454 ( n13011 , n6590 , n1985 );
    or g7455 ( n7547 , n6509 , n9590 );
    and g7456 ( n9199 , n4736 , n5256 );
    or g7457 ( n9240 , n9489 , n5242 );
    nor g7458 ( n4057 , n4840 , n5887 );
    or g7459 ( n10172 , n4495 , n8499 );
    and g7460 ( n11583 , n8026 , n9623 );
    xnor g7461 ( n9818 , n11599 , n8226 );
    not g7462 ( n13052 , n5965 );
    or g7463 ( n2098 , n7418 , n11744 );
    not g7464 ( n6630 , n497 );
    and g7465 ( n8983 , n4164 , n5441 );
    not g7466 ( n5974 , n9212 );
    or g7467 ( n10155 , n12552 , n8030 );
    or g7468 ( n4883 , n5370 , n5983 );
    or g7469 ( n5993 , n8646 , n177 );
    not g7470 ( n9910 , n7671 );
    and g7471 ( n7452 , n6533 , n427 );
    not g7472 ( n5522 , n7919 );
    xnor g7473 ( n5358 , n6254 , n4367 );
    xnor g7474 ( n3693 , n3770 , n10758 );
    xnor g7475 ( n11895 , n9578 , n213 );
    and g7476 ( n10146 , n10388 , n10700 );
    not g7477 ( n3063 , n5576 );
    and g7478 ( n3987 , n11596 , n11721 );
    and g7479 ( n5346 , n6943 , n3637 );
    and g7480 ( n8660 , n5776 , n924 );
    nor g7481 ( n1614 , n2379 , n690 );
    xnor g7482 ( n7516 , n3138 , n7058 );
    not g7483 ( n7872 , n11109 );
    not g7484 ( n10882 , n4528 );
    or g7485 ( n3579 , n3564 , n10871 );
    and g7486 ( n10288 , n6194 , n2721 );
    or g7487 ( n3984 , n2889 , n10319 );
    or g7488 ( n2663 , n9695 , n8305 );
    not g7489 ( n12859 , n12670 );
    and g7490 ( n7885 , n11878 , n7390 );
    nor g7491 ( n3295 , n5742 , n12170 );
    xnor g7492 ( n3357 , n7751 , n750 );
    or g7493 ( n10446 , n9017 , n8534 );
    or g7494 ( n1072 , n8131 , n1985 );
    or g7495 ( n4189 , n11033 , n2126 );
    not g7496 ( n4714 , n2856 );
    and g7497 ( n6036 , n8248 , n7155 );
    xnor g7498 ( n2374 , n7496 , n9981 );
    or g7499 ( n844 , n1715 , n8313 );
    not g7500 ( n9272 , n10063 );
    and g7501 ( n1138 , n10142 , n13058 );
    not g7502 ( n1051 , n7113 );
    and g7503 ( n4358 , n5592 , n4607 );
    or g7504 ( n12037 , n10410 , n4073 );
    xnor g7505 ( n6251 , n3145 , n1583 );
    and g7506 ( n9014 , n10943 , n6511 );
    or g7507 ( n8396 , n6129 , n4947 );
    xnor g7508 ( n2873 , n5926 , n10884 );
    not g7509 ( n3257 , n194 );
    not g7510 ( n4808 , n4335 );
    not g7511 ( n812 , n3431 );
    and g7512 ( n9585 , n7772 , n7411 );
    and g7513 ( n12709 , n6605 , n9094 );
    or g7514 ( n12775 , n10421 , n12388 );
    xnor g7515 ( n87 , n2658 , n10396 );
    not g7516 ( n2674 , n5998 );
    and g7517 ( n6577 , n9691 , n217 );
    and g7518 ( n1003 , n5097 , n8002 );
    or g7519 ( n4876 , n3301 , n1415 );
    xnor g7520 ( n12313 , n11560 , n10646 );
    xnor g7521 ( n3849 , n4252 , n12666 );
    not g7522 ( n10794 , n13087 );
    or g7523 ( n8444 , n5720 , n8502 );
    or g7524 ( n10189 , n6148 , n11494 );
    or g7525 ( n3184 , n2528 , n7924 );
    buf g7526 ( n8760 , n11123 );
    not g7527 ( n5654 , n8308 );
    xnor g7528 ( n5032 , n589 , n7217 );
    or g7529 ( n6480 , n5266 , n3380 );
    not g7530 ( n8728 , n1495 );
    and g7531 ( n7655 , n6480 , n6835 );
    or g7532 ( n12990 , n3225 , n7530 );
    xnor g7533 ( n1409 , n4760 , n12516 );
    and g7534 ( n9285 , n8389 , n7192 );
    xnor g7535 ( n3198 , n4042 , n2271 );
    nor g7536 ( n7124 , n2458 , n8230 );
    not g7537 ( n7473 , n8357 );
    xnor g7538 ( n8184 , n6961 , n1527 );
    xnor g7539 ( n11410 , n5353 , n4456 );
    or g7540 ( n5514 , n7234 , n12718 );
    xnor g7541 ( n9312 , n9883 , n8404 );
    not g7542 ( n13154 , n287 );
    xnor g7543 ( n11298 , n12816 , n8037 );
    and g7544 ( n2149 , n10908 , n6937 );
    and g7545 ( n11963 , n3503 , n11070 );
    xnor g7546 ( n11529 , n3593 , n1455 );
    and g7547 ( n4881 , n11235 , n6113 );
    or g7548 ( n8154 , n10158 , n1583 );
    and g7549 ( n8509 , n6119 , n4432 );
    xnor g7550 ( n9932 , n9407 , n1933 );
    or g7551 ( n12806 , n7532 , n4724 );
    or g7552 ( n9853 , n6215 , n4453 );
    or g7553 ( n5150 , n8030 , n4640 );
    or g7554 ( n842 , n1163 , n3920 );
    xnor g7555 ( n2525 , n8996 , n6592 );
    and g7556 ( n8997 , n10014 , n8235 );
    or g7557 ( n8766 , n12469 , n8534 );
    or g7558 ( n8610 , n3730 , n12302 );
    nor g7559 ( n11082 , n10850 , n1486 );
    and g7560 ( n3820 , n3956 , n13123 );
    not g7561 ( n1521 , n2690 );
    xnor g7562 ( n12232 , n8074 , n9615 );
    and g7563 ( n12909 , n4771 , n12332 );
    and g7564 ( n11026 , n3719 , n9958 );
    xnor g7565 ( n7534 , n4842 , n858 );
    xor g7566 ( n2595 , n2220 , n2198 );
    and g7567 ( n11204 , n4187 , n10512 );
    and g7568 ( n289 , n7927 , n7456 );
    and g7569 ( n11176 , n12227 , n11286 );
    or g7570 ( n7518 , n8583 , n11524 );
    or g7571 ( n11924 , n6112 , n12623 );
    xnor g7572 ( n3137 , n3283 , n4281 );
    not g7573 ( n9132 , n7115 );
    nor g7574 ( n8018 , n8297 , n13055 );
    or g7575 ( n5516 , n1939 , n8116 );
    and g7576 ( n1628 , n7516 , n1236 );
    or g7577 ( n615 , n6875 , n12847 );
    or g7578 ( n8388 , n3344 , n8609 );
    xnor g7579 ( n12865 , n6424 , n6884 );
    or g7580 ( n5135 , n6175 , n1192 );
    xnor g7581 ( n9857 , n3255 , n12672 );
    or g7582 ( n1959 , n1215 , n8511 );
    not g7583 ( n3243 , n11396 );
    or g7584 ( n11399 , n3636 , n10341 );
    xor g7585 ( n11567 , n12990 , n1024 );
    xnor g7586 ( n3796 , n4334 , n12958 );
    not g7587 ( n521 , n11873 );
    not g7588 ( n963 , n6611 );
    or g7589 ( n3827 , n12512 , n10249 );
    xnor g7590 ( n10450 , n2282 , n5940 );
    or g7591 ( n1213 , n12604 , n2449 );
    xnor g7592 ( n8608 , n7199 , n10924 );
    not g7593 ( n6944 , n834 );
    xnor g7594 ( n5431 , n9993 , n6275 );
    not g7595 ( n413 , n3623 );
    not g7596 ( n6524 , n7417 );
    xnor g7597 ( n1339 , n810 , n8138 );
    not g7598 ( n61 , n11091 );
    xnor g7599 ( n1537 , n12530 , n797 );
    xnor g7600 ( n9990 , n6614 , n6996 );
    not g7601 ( n5200 , n12589 );
    not g7602 ( n3634 , n8860 );
    nor g7603 ( n7200 , n82 , n2481 );
    or g7604 ( n12236 , n7234 , n206 );
    or g7605 ( n8426 , n11729 , n5797 );
    xnor g7606 ( n9532 , n10704 , n778 );
    nor g7607 ( n11034 , n9826 , n8261 );
    not g7608 ( n9055 , n11089 );
    nor g7609 ( n5648 , n6534 , n3474 );
    and g7610 ( n4193 , n7322 , n730 );
    not g7611 ( n2872 , n9531 );
    not g7612 ( n4198 , n3769 );
    xnor g7613 ( n3624 , n8311 , n6836 );
    or g7614 ( n4749 , n8665 , n12655 );
    or g7615 ( n12333 , n11157 , n8030 );
    xnor g7616 ( n2797 , n973 , n2281 );
    or g7617 ( n59 , n3531 , n4230 );
    xnor g7618 ( n9719 , n8429 , n11443 );
    and g7619 ( n11316 , n10215 , n5929 );
    not g7620 ( n2899 , n817 );
    not g7621 ( n5709 , n11974 );
    or g7622 ( n9567 , n2129 , n4373 );
    not g7623 ( n4371 , n7128 );
    and g7624 ( n3422 , n1496 , n5844 );
    or g7625 ( n10301 , n12166 , n1197 );
    and g7626 ( n11980 , n10931 , n1903 );
    or g7627 ( n3557 , n8362 , n6181 );
    xnor g7628 ( n2494 , n8004 , n2981 );
    and g7629 ( n4906 , n3507 , n5717 );
    not g7630 ( n53 , n761 );
    or g7631 ( n2299 , n7129 , n2617 );
    and g7632 ( n3303 , n10770 , n287 );
    or g7633 ( n10190 , n333 , n12967 );
    not g7634 ( n8529 , n5969 );
    xnor g7635 ( n4130 , n5934 , n12002 );
    and g7636 ( n11188 , n10849 , n7784 );
    or g7637 ( n9059 , n5947 , n12695 );
    and g7638 ( n1410 , n10642 , n7720 );
    buf g7639 ( n8268 , n765 );
    or g7640 ( n6354 , n7608 , n206 );
    xnor g7641 ( n2230 , n12141 , n12407 );
    xor g7642 ( n6362 , n4349 , n2419 );
    xnor g7643 ( n3250 , n1121 , n12125 );
    not g7644 ( n1767 , n12950 );
    nor g7645 ( n9235 , n12237 , n2512 );
    not g7646 ( n6264 , n2754 );
    or g7647 ( n4836 , n7719 , n275 );
    and g7648 ( n6325 , n13201 , n3085 );
    nor g7649 ( n6842 , n4684 , n12927 );
    or g7650 ( n8653 , n11103 , n5388 );
    nor g7651 ( n6207 , n8773 , n4345 );
    or g7652 ( n745 , n5569 , n7221 );
    and g7653 ( n6729 , n3517 , n3571 );
    or g7654 ( n7703 , n12416 , n9159 );
    or g7655 ( n13115 , n11450 , n4757 );
    not g7656 ( n5865 , n11835 );
    xnor g7657 ( n4951 , n5793 , n1990 );
    not g7658 ( n9772 , n1342 );
    and g7659 ( n2324 , n10565 , n5585 );
    or g7660 ( n810 , n12671 , n10430 );
    nor g7661 ( n7488 , n11883 , n9598 );
    not g7662 ( n2056 , n5451 );
    or g7663 ( n11055 , n379 , n2816 );
    and g7664 ( n928 , n4052 , n109 );
    xnor g7665 ( n1563 , n4509 , n875 );
    or g7666 ( n7546 , n6680 , n2890 );
    or g7667 ( n1593 , n8011 , n2772 );
    xnor g7668 ( n7034 , n94 , n6935 );
    xnor g7669 ( n10518 , n10671 , n1317 );
    or g7670 ( n8866 , n13013 , n0 );
    or g7671 ( n7874 , n3826 , n10106 );
    not g7672 ( n1073 , n7749 );
    and g7673 ( n11219 , n5113 , n9133 );
    xnor g7674 ( n5757 , n1077 , n11598 );
    or g7675 ( n8979 , n2484 , n10552 );
    or g7676 ( n9053 , n2391 , n2531 );
    and g7677 ( n6971 , n1107 , n10571 );
    and g7678 ( n12539 , n8153 , n11275 );
    buf g7679 ( n11668 , n9280 );
    or g7680 ( n238 , n1206 , n11490 );
    or g7681 ( n1879 , n8665 , n1720 );
    or g7682 ( n6945 , n3796 , n12724 );
    or g7683 ( n2812 , n9098 , n6002 );
    xnor g7684 ( n7724 , n1338 , n4471 );
    not g7685 ( n173 , n10906 );
    not g7686 ( n10039 , n7144 );
    and g7687 ( n4078 , n12348 , n5065 );
    and g7688 ( n4533 , n10078 , n11040 );
    not g7689 ( n2350 , n10301 );
    or g7690 ( n4829 , n12951 , n7988 );
    or g7691 ( n4885 , n9882 , n11300 );
    not g7692 ( n12183 , n6242 );
    and g7693 ( n4354 , n3982 , n752 );
    not g7694 ( n7072 , n4399 );
    xnor g7695 ( n148 , n10377 , n3608 );
    and g7696 ( n10350 , n5516 , n6976 );
    not g7697 ( n5097 , n7605 );
    and g7698 ( n2827 , n767 , n3832 );
    xnor g7699 ( n1806 , n10455 , n1147 );
    xnor g7700 ( n5487 , n4558 , n1811 );
    and g7701 ( n5656 , n5530 , n1068 );
    nor g7702 ( n10612 , n5391 , n9231 );
    not g7703 ( n1018 , n9313 );
    xnor g7704 ( n5003 , n953 , n8746 );
    xnor g7705 ( n12692 , n3607 , n2525 );
    or g7706 ( n1749 , n6913 , n9650 );
    or g7707 ( n208 , n11980 , n8375 );
    not g7708 ( n490 , n2869 );
    or g7709 ( n7106 , n8766 , n2647 );
    xnor g7710 ( n9105 , n1141 , n10521 );
    xor g7711 ( n7515 , n3613 , n12527 );
    not g7712 ( n6112 , n8332 );
    and g7713 ( n873 , n4173 , n7275 );
    nor g7714 ( n4817 , n3502 , n3857 );
    or g7715 ( n4467 , n3208 , n7221 );
    and g7716 ( n2126 , n4659 , n3151 );
    or g7717 ( n12792 , n3818 , n12040 );
    and g7718 ( n9611 , n2008 , n12318 );
    not g7719 ( n11284 , n11222 );
    xnor g7720 ( n3899 , n4568 , n2693 );
    or g7721 ( n2887 , n1416 , n4967 );
    or g7722 ( n7519 , n4478 , n1599 );
    or g7723 ( n2424 , n6769 , n7935 );
    not g7724 ( n3619 , n12661 );
    or g7725 ( n10277 , n2424 , n6729 );
    not g7726 ( n9558 , n12750 );
    nor g7727 ( n9173 , n9200 , n5471 );
    or g7728 ( n6719 , n12607 , n8041 );
    nor g7729 ( n11161 , n7375 , n10819 );
    xnor g7730 ( n9946 , n1871 , n10868 );
    or g7731 ( n2644 , n6488 , n6265 );
    xor g7732 ( n1022 , n10318 , n11196 );
    or g7733 ( n1679 , n10966 , n9075 );
    or g7734 ( n9042 , n9575 , n1500 );
    not g7735 ( n657 , n2841 );
    and g7736 ( n1 , n8430 , n10255 );
    xnor g7737 ( n4177 , n6292 , n10418 );
    xnor g7738 ( n8635 , n12815 , n3799 );
    and g7739 ( n2375 , n1759 , n11382 );
    and g7740 ( n4798 , n9239 , n487 );
    xnor g7741 ( n11112 , n2144 , n11001 );
    or g7742 ( n12210 , n6129 , n11144 );
    and g7743 ( n7016 , n3444 , n7652 );
    not g7744 ( n3058 , n2482 );
    or g7745 ( n9662 , n8992 , n541 );
    xnor g7746 ( n6154 , n1540 , n6221 );
    or g7747 ( n5133 , n5842 , n6033 );
    or g7748 ( n3869 , n12465 , n13086 );
    xnor g7749 ( n11090 , n12791 , n6666 );
    nor g7750 ( n3872 , n570 , n3366 );
    and g7751 ( n6950 , n103 , n854 );
    and g7752 ( n5186 , n7622 , n8815 );
    or g7753 ( n10674 , n4844 , n9075 );
    not g7754 ( n5136 , n7214 );
    or g7755 ( n12504 , n6476 , n8663 );
    and g7756 ( n11681 , n9417 , n256 );
    xnor g7757 ( n11036 , n8109 , n3515 );
    xnor g7758 ( n6261 , n2203 , n7623 );
    xnor g7759 ( n3306 , n11775 , n665 );
    or g7760 ( n10938 , n227 , n6635 );
    and g7761 ( n12824 , n8175 , n7616 );
    xor g7762 ( n2829 , n5786 , n1687 );
    and g7763 ( n10778 , n5217 , n12011 );
    not g7764 ( n11790 , n12134 );
    nor g7765 ( n5599 , n889 , n7897 );
    or g7766 ( n7230 , n4890 , n4936 );
    or g7767 ( n11825 , n7210 , n12499 );
    xnor g7768 ( n10825 , n6650 , n3390 );
    or g7769 ( n9814 , n11187 , n8517 );
    xnor g7770 ( n7550 , n4260 , n2093 );
    not g7771 ( n6881 , n12539 );
    xnor g7772 ( n607 , n4708 , n10644 );
    and g7773 ( n11443 , n6267 , n3400 );
    or g7774 ( n11119 , n8105 , n13204 );
    xnor g7775 ( n5763 , n5015 , n11380 );
    not g7776 ( n8719 , n3828 );
    not g7777 ( n2394 , n9536 );
    or g7778 ( n1777 , n2622 , n8268 );
    not g7779 ( n2452 , n3409 );
    and g7780 ( n11968 , n4791 , n11517 );
    xnor g7781 ( n11997 , n13134 , n3935 );
    or g7782 ( n10603 , n3225 , n2675 );
    or g7783 ( n3728 , n11114 , n11522 );
    xnor g7784 ( n9652 , n2294 , n13017 );
    not g7785 ( n12211 , n3756 );
    xnor g7786 ( n5463 , n7192 , n8389 );
    xnor g7787 ( n277 , n10323 , n1955 );
    or g7788 ( n7773 , n10462 , n4230 );
    and g7789 ( n3648 , n12264 , n12355 );
    not g7790 ( n8913 , n2354 );
    and g7791 ( n2490 , n12266 , n11625 );
    xnor g7792 ( n4027 , n369 , n5339 );
    xor g7793 ( n4387 , n12987 , n3141 );
    not g7794 ( n7925 , n443 );
    not g7795 ( n7533 , n9062 );
    and g7796 ( n4624 , n9132 , n770 );
    or g7797 ( n95 , n2416 , n8534 );
    xnor g7798 ( n3626 , n11098 , n4280 );
    xnor g7799 ( n1112 , n13211 , n8725 );
    not g7800 ( n1117 , n2591 );
    xnor g7801 ( n8054 , n5370 , n5983 );
    xnor g7802 ( n11445 , n8836 , n6953 );
    xnor g7803 ( n2567 , n9654 , n2866 );
    xnor g7804 ( n7511 , n3807 , n5624 );
    or g7805 ( n6735 , n6028 , n7723 );
    xnor g7806 ( n1615 , n2699 , n8946 );
    nor g7807 ( n5680 , n4400 , n12285 );
    xnor g7808 ( n11221 , n2237 , n9081 );
    not g7809 ( n8511 , n3845 );
    and g7810 ( n7336 , n879 , n12413 );
    or g7811 ( n9976 , n6354 , n8707 );
    and g7812 ( n3141 , n8259 , n12511 );
    xnor g7813 ( n12611 , n400 , n8596 );
    xnor g7814 ( n10216 , n5133 , n10020 );
    not g7815 ( n2416 , n9570 );
    nor g7816 ( n5734 , n20 , n732 );
    nor g7817 ( n3065 , n10191 , n9414 );
    not g7818 ( n12324 , n7720 );
    and g7819 ( n9543 , n684 , n8617 );
    xor g7820 ( n8884 , n2640 , n9983 );
    xnor g7821 ( n8851 , n10600 , n3897 );
    not g7822 ( n1847 , n4874 );
    xnor g7823 ( n4150 , n5140 , n6791 );
    or g7824 ( n12744 , n971 , n3981 );
    not g7825 ( n12748 , n12651 );
    buf g7826 ( n12188 , n9257 );
    or g7827 ( n7739 , n3127 , n3949 );
    and g7828 ( n2633 , n349 , n11283 );
    xnor g7829 ( n6384 , n10602 , n2771 );
    xor g7830 ( n11149 , n3544 , n10553 );
    not g7831 ( n3616 , n2341 );
    xnor g7832 ( n4043 , n10592 , n12502 );
    xnor g7833 ( n11962 , n8883 , n9479 );
    and g7834 ( n5274 , n4305 , n407 );
    not g7835 ( n4294 , n12990 );
    not g7836 ( n868 , n11663 );
    or g7837 ( n5456 , n6048 , n5919 );
    not g7838 ( n12316 , n10142 );
    nor g7839 ( n10089 , n12339 , n8342 );
    not g7840 ( n12425 , n1700 );
    not g7841 ( n119 , n3815 );
    and g7842 ( n5121 , n10908 , n5065 );
    not g7843 ( n1269 , n2388 );
    nor g7844 ( n7803 , n7613 , n12303 );
    xnor g7845 ( n7759 , n4858 , n6896 );
    xnor g7846 ( n10817 , n6694 , n11017 );
    xnor g7847 ( n4423 , n5424 , n3838 );
    or g7848 ( n7187 , n7263 , n12492 );
    xnor g7849 ( n7439 , n1048 , n378 );
    not g7850 ( n2330 , n8267 );
    and g7851 ( n1569 , n13147 , n2602 );
    xnor g7852 ( n11931 , n3533 , n4754 );
    xnor g7853 ( n8043 , n11386 , n1497 );
    and g7854 ( n12443 , n2273 , n1598 );
    nor g7855 ( n8130 , n1471 , n13033 );
    or g7856 ( n6518 , n5626 , n12291 );
    and g7857 ( n3581 , n9897 , n897 );
    xnor g7858 ( n12208 , n6521 , n7565 );
    nor g7859 ( n7134 , n4689 , n4705 );
    not g7860 ( n1820 , n8290 );
    and g7861 ( n11613 , n1965 , n11784 );
    not g7862 ( n10120 , n12477 );
    or g7863 ( n7607 , n10761 , n2675 );
    not g7864 ( n2848 , n11111 );
    xnor g7865 ( n12024 , n8432 , n8045 );
    not g7866 ( n1967 , n9481 );
    or g7867 ( n2027 , n9868 , n1043 );
    xnor g7868 ( n12139 , n12011 , n4897 );
    xnor g7869 ( n9794 , n8387 , n10333 );
    not g7870 ( n10508 , n7384 );
    and g7871 ( n7831 , n6880 , n5072 );
    and g7872 ( n11663 , n12478 , n13139 );
    or g7873 ( n8816 , n36 , n1703 );
    and g7874 ( n6248 , n372 , n12572 );
    not g7875 ( n7049 , n10606 );
    or g7876 ( n6923 , n7787 , n6878 );
    and g7877 ( n10269 , n12380 , n5082 );
    or g7878 ( n1751 , n6735 , n9791 );
    xnor g7879 ( n4383 , n897 , n4126 );
    and g7880 ( n3328 , n10771 , n1878 );
    not g7881 ( n5469 , n9847 );
    not g7882 ( n9436 , n11012 );
    not g7883 ( n4132 , n2339 );
    nor g7884 ( n11938 , n8996 , n3607 );
    not g7885 ( n12224 , n7659 );
    not g7886 ( n12254 , n2339 );
    not g7887 ( n2956 , n1344 );
    or g7888 ( n3966 , n1354 , n7723 );
    xnor g7889 ( n7822 , n13145 , n319 );
    and g7890 ( n5631 , n5236 , n9954 );
    or g7891 ( n10742 , n8598 , n4640 );
    or g7892 ( n3992 , n9113 , n10179 );
    and g7893 ( n2959 , n6241 , n1846 );
    and g7894 ( n5368 , n4379 , n2897 );
    not g7895 ( n10127 , n10876 );
    not g7896 ( n8492 , n6209 );
    xnor g7897 ( n5560 , n2766 , n7566 );
    xnor g7898 ( n11886 , n5161 , n6116 );
    nor g7899 ( n3162 , n6780 , n8855 );
    not g7900 ( n7544 , n11372 );
    or g7901 ( n11530 , n4620 , n2675 );
    or g7902 ( n10520 , n11392 , n9760 );
    nor g7903 ( n12733 , n8057 , n4415 );
    xor g7904 ( n8399 , n8954 , n11294 );
    not g7905 ( n9113 , n10874 );
    and g7906 ( n10100 , n2563 , n1509 );
    or g7907 ( n7508 , n7438 , n3732 );
    or g7908 ( n11288 , n7191 , n1144 );
    nor g7909 ( n12727 , n12333 , n12640 );
    not g7910 ( n10462 , n1916 );
    or g7911 ( n1673 , n8426 , n11754 );
    not g7912 ( n7614 , n9052 );
    xnor g7913 ( n8007 , n2804 , n10678 );
    and g7914 ( n1143 , n10425 , n10380 );
    xnor g7915 ( n9943 , n2618 , n11179 );
    and g7916 ( n2695 , n10493 , n9927 );
    or g7917 ( n5980 , n11864 , n7961 );
    not g7918 ( n12000 , n9591 );
    or g7919 ( n9748 , n2759 , n3653 );
    or g7920 ( n12999 , n5296 , n2277 );
    or g7921 ( n7674 , n6854 , n8268 );
    not g7922 ( n11398 , n13212 );
    or g7923 ( n1838 , n10784 , n10576 );
    xnor g7924 ( n7853 , n8682 , n9351 );
    xnor g7925 ( n1721 , n9579 , n7024 );
    or g7926 ( n11829 , n8091 , n10932 );
    nor g7927 ( n793 , n6965 , n1626 );
    or g7928 ( n4859 , n1150 , n6005 );
    not g7929 ( n11418 , n10416 );
    xnor g7930 ( n9753 , n8981 , n598 );
    not g7931 ( n4257 , n2012 );
    nor g7932 ( n9689 , n4233 , n5229 );
    or g7933 ( n5844 , n1335 , n3890 );
    xnor g7934 ( n3436 , n7321 , n11993 );
    and g7935 ( n10214 , n11074 , n8753 );
    and g7936 ( n5413 , n9403 , n4578 );
    not g7937 ( n1881 , n3910 );
    or g7938 ( n8264 , n1618 , n12273 );
    not g7939 ( n8877 , n1291 );
    and g7940 ( n245 , n761 , n5548 );
    nor g7941 ( n10899 , n5952 , n205 );
    or g7942 ( n9646 , n10501 , n4373 );
    and g7943 ( n517 , n5384 , n6118 );
    nor g7944 ( n2990 , n12928 , n2247 );
    not g7945 ( n2013 , n5952 );
    or g7946 ( n10536 , n10637 , n9234 );
    not g7947 ( n6724 , n12408 );
    or g7948 ( n6202 , n8904 , n10029 );
    or g7949 ( n1817 , n4038 , n9984 );
    xnor g7950 ( n835 , n344 , n6639 );
    nor g7951 ( n8933 , n2910 , n1430 );
    xnor g7952 ( n2839 , n12020 , n964 );
    or g7953 ( n7253 , n2097 , n2917 );
    xnor g7954 ( n7915 , n8805 , n11623 );
    and g7955 ( n12532 , n6369 , n13167 );
    and g7956 ( n764 , n8228 , n5920 );
    xnor g7957 ( n12950 , n1125 , n12488 );
    not g7958 ( n7730 , n5167 );
    nor g7959 ( n3864 , n5294 , n8289 );
    or g7960 ( n4167 , n9113 , n177 );
    and g7961 ( n3398 , n8877 , n11133 );
    xnor g7962 ( n7268 , n8923 , n7479 );
    or g7963 ( n973 , n13026 , n177 );
    and g7964 ( n7464 , n9303 , n11029 );
    or g7965 ( n944 , n9371 , n12016 );
    and g7966 ( n6550 , n1586 , n2253 );
    not g7967 ( n10437 , n1302 );
    or g7968 ( n4485 , n1529 , n604 );
    xnor g7969 ( n5418 , n9221 , n12344 );
    xnor g7970 ( n11716 , n6952 , n8149 );
    nor g7971 ( n12541 , n7349 , n12447 );
    xnor g7972 ( n6017 , n12821 , n9452 );
    xnor g7973 ( n12531 , n10088 , n12494 );
    and g7974 ( n1183 , n6168 , n12853 );
    and g7975 ( n9744 , n13041 , n3661 );
    or g7976 ( n7953 , n1261 , n177 );
    xnor g7977 ( n13142 , n9588 , n10708 );
    or g7978 ( n190 , n9983 , n8246 );
    nor g7979 ( n1690 , n11837 , n913 );
    and g7980 ( n5112 , n6100 , n10389 );
    not g7981 ( n13036 , n9187 );
    xnor g7982 ( n4449 , n3923 , n261 );
    and g7983 ( n2082 , n7990 , n3609 );
    xnor g7984 ( n6696 , n4988 , n9686 );
    or g7985 ( n12198 , n1947 , n8018 );
    or g7986 ( n9342 , n1334 , n7926 );
    not g7987 ( n128 , n13011 );
    not g7988 ( n881 , n10951 );
    or g7989 ( n8401 , n1727 , n8083 );
    xnor g7990 ( n717 , n475 , n10012 );
    and g7991 ( n9324 , n8948 , n8786 );
    nor g7992 ( n11234 , n10186 , n10206 );
    and g7993 ( n888 , n8295 , n6694 );
    not g7994 ( n1353 , n4748 );
    xnor g7995 ( n5901 , n3973 , n11389 );
    xnor g7996 ( n4570 , n1426 , n3751 );
    not g7997 ( n11352 , n7411 );
    or g7998 ( n12446 , n1068 , n5530 );
    not g7999 ( n9008 , n7164 );
    xnor g8000 ( n1835 , n175 , n9377 );
    nor g8001 ( n5253 , n625 , n9390 );
    and g8002 ( n3461 , n10676 , n1091 );
    xnor g8003 ( n6704 , n633 , n1000 );
    or g8004 ( n5744 , n9739 , n10106 );
    or g8005 ( n7219 , n11256 , n9657 );
    and g8006 ( n12394 , n1315 , n10174 );
    xnor g8007 ( n5023 , n3179 , n11465 );
    xnor g8008 ( n2647 , n8428 , n11341 );
    xnor g8009 ( n6730 , n6498 , n4246 );
    or g8010 ( n1507 , n734 , n10956 );
    xnor g8011 ( n8731 , n962 , n11405 );
    or g8012 ( n9389 , n11007 , n2675 );
    xnor g8013 ( n11556 , n9823 , n2704 );
    not g8014 ( n5420 , n3181 );
    and g8015 ( n11338 , n21 , n2740 );
    or g8016 ( n7777 , n2217 , n10871 );
    xor g8017 ( n9039 , n6068 , n5834 );
    and g8018 ( n10432 , n3161 , n3249 );
    nor g8019 ( n7627 , n9678 , n5171 );
    or g8020 ( n10731 , n992 , n7239 );
    not g8021 ( n8012 , n3283 );
    not g8022 ( n3816 , n5062 );
    not g8023 ( n8481 , n3939 );
    xnor g8024 ( n5702 , n7096 , n7458 );
    or g8025 ( n2963 , n9226 , n9521 );
    or g8026 ( n7972 , n10919 , n4765 );
    xnor g8027 ( n1449 , n12894 , n6459 );
    xnor g8028 ( n10968 , n11710 , n11702 );
    or g8029 ( n8703 , n7900 , n10106 );
    not g8030 ( n2430 , n10458 );
    and g8031 ( n11056 , n5400 , n4047 );
    xnor g8032 ( n3959 , n7542 , n3710 );
    or g8033 ( n9205 , n11965 , n4844 );
    and g8034 ( n9619 , n4382 , n11109 );
    or g8035 ( n2106 , n3327 , n926 );
    not g8036 ( n7672 , n12579 );
    and g8037 ( n10985 , n9135 , n12548 );
    and g8038 ( n5770 , n3311 , n6085 );
    nor g8039 ( n9524 , n4851 , n2998 );
    or g8040 ( n9153 , n4213 , n4255 );
    xnor g8041 ( n10119 , n6268 , n4358 );
    not g8042 ( n8400 , n11109 );
    or g8043 ( n8 , n8645 , n8563 );
    and g8044 ( n5378 , n11430 , n7519 );
    xnor g8045 ( n2364 , n8638 , n10679 );
    and g8046 ( n5978 , n818 , n6563 );
    xnor g8047 ( n10621 , n12851 , n13112 );
    or g8048 ( n2062 , n4198 , n4373 );
    not g8049 ( n8723 , n105 );
    not g8050 ( n6638 , n7374 );
    and g8051 ( n8433 , n325 , n3739 );
    not g8052 ( n2385 , n7802 );
    xnor g8053 ( n13231 , n4785 , n4120 );
    or g8054 ( n9318 , n6841 , n8129 );
    and g8055 ( n3372 , n4485 , n5936 );
    xnor g8056 ( n7604 , n3032 , n847 );
    and g8057 ( n11169 , n9707 , n8888 );
    not g8058 ( n8540 , n10787 );
    xnor g8059 ( n6148 , n11742 , n3098 );
    or g8060 ( n8833 , n3724 , n7959 );
    xor g8061 ( n6526 , n3395 , n11402 );
    and g8062 ( n2944 , n11592 , n4491 );
    xnor g8063 ( n3694 , n6176 , n13062 );
    or g8064 ( n9617 , n7069 , n1694 );
    or g8065 ( n2897 , n12758 , n5797 );
    not g8066 ( n5842 , n951 );
    nor g8067 ( n4545 , n12897 , n5133 );
    nor g8068 ( n9388 , n5323 , n4094 );
    or g8069 ( n9124 , n8082 , n1026 );
    xnor g8070 ( n10556 , n29 , n7029 );
    xnor g8071 ( n7345 , n10762 , n363 );
    and g8072 ( n6462 , n11702 , n11710 );
    xnor g8073 ( n10744 , n4232 , n5137 );
    nor g8074 ( n4983 , n2951 , n4369 );
    and g8075 ( n11785 , n2465 , n1868 );
    not g8076 ( n5875 , n5920 );
    and g8077 ( n5171 , n10727 , n1967 );
    and g8078 ( n2883 , n2068 , n12284 );
    or g8079 ( n8984 , n11102 , n2280 );
    not g8080 ( n1055 , n2791 );
    nor g8081 ( n3238 , n6892 , n9952 );
    xnor g8082 ( n13219 , n2370 , n13161 );
    xnor g8083 ( n6832 , n5627 , n9009 );
    not g8084 ( n4398 , n7059 );
    xnor g8085 ( n4797 , n6352 , n9616 );
    xnor g8086 ( n9508 , n12988 , n2012 );
    and g8087 ( n4482 , n3209 , n8760 );
    xnor g8088 ( n1412 , n3666 , n10218 );
    xnor g8089 ( n11976 , n12097 , n1375 );
    not g8090 ( n7073 , n3199 );
    xnor g8091 ( n9467 , n4602 , n11487 );
    xnor g8092 ( n8119 , n402 , n12679 );
    not g8093 ( n813 , n9528 );
    and g8094 ( n8326 , n7319 , n12764 );
    or g8095 ( n5474 , n5993 , n1298 );
    xnor g8096 ( n6535 , n2088 , n11731 );
    or g8097 ( n6929 , n7730 , n3825 );
    xor g8098 ( n8675 , n6522 , n11840 );
    buf g8099 ( n4640 , n12128 );
    and g8100 ( n9061 , n525 , n10753 );
    xnor g8101 ( n1092 , n7363 , n11216 );
    or g8102 ( n9326 , n2046 , n12637 );
    and g8103 ( n12784 , n5823 , n5381 );
    and g8104 ( n11666 , n5522 , n11056 );
    xnor g8105 ( n733 , n8424 , n2225 );
    xnor g8106 ( n2597 , n12590 , n4410 );
    or g8107 ( n6378 , n4983 , n553 );
    or g8108 ( n1821 , n8950 , n12695 );
    not g8109 ( n1366 , n10869 );
    or g8110 ( n7569 , n6749 , n7076 );
    or g8111 ( n5187 , n12458 , n4303 );
    xnor g8112 ( n9941 , n10312 , n4353 );
    or g8113 ( n1711 , n1158 , n1713 );
    or g8114 ( n5090 , n9913 , n11868 );
    nor g8115 ( n12826 , n7442 , n12464 );
    xnor g8116 ( n12061 , n7694 , n9438 );
    or g8117 ( n4827 , n2462 , n10319 );
    not g8118 ( n5460 , n3769 );
    or g8119 ( n2607 , n294 , n11164 );
    buf g8120 ( n11084 , n3527 );
    not g8121 ( n1134 , n2619 );
    or g8122 ( n8878 , n10332 , n1344 );
    or g8123 ( n671 , n3957 , n11273 );
    or g8124 ( n3213 , n9383 , n3981 );
    nor g8125 ( n13233 , n11973 , n12163 );
    or g8126 ( n3345 , n2723 , n4209 );
    or g8127 ( n7275 , n10999 , n10342 );
    nor g8128 ( n9500 , n4403 , n1828 );
    not g8129 ( n8259 , n2966 );
    and g8130 ( n4565 , n10920 , n5497 );
    xnor g8131 ( n7172 , n8606 , n3342 );
    and g8132 ( n6795 , n6136 , n8022 );
    xnor g8133 ( n10829 , n2995 , n2840 );
    not g8134 ( n8800 , n5722 );
    not g8135 ( n3116 , n2647 );
    not g8136 ( n7532 , n497 );
    nor g8137 ( n5849 , n13070 , n6840 );
    or g8138 ( n1997 , n7770 , n8066 );
    or g8139 ( n9020 , n10149 , n9413 );
    buf g8140 ( n5242 , n1750 );
    or g8141 ( n7468 , n719 , n290 );
    and g8142 ( n9773 , n1912 , n13060 );
    xnor g8143 ( n2704 , n10766 , n7287 );
    xnor g8144 ( n5364 , n10390 , n12034 );
    not g8145 ( n7784 , n13223 );
    nor g8146 ( n6963 , n5800 , n1624 );
    or g8147 ( n3571 , n9162 , n12328 );
    not g8148 ( n5533 , n3043 );
    not g8149 ( n2135 , n1982 );
    or g8150 ( n2380 , n5465 , n6861 );
    not g8151 ( n7191 , n12651 );
    and g8152 ( n11626 , n8584 , n4814 );
    xor g8153 ( n10769 , n8731 , n9437 );
    xnor g8154 ( n7107 , n8457 , n6903 );
    or g8155 ( n13085 , n2789 , n8029 );
    and g8156 ( n3615 , n12933 , n3526 );
    not g8157 ( n3118 , n12217 );
    or g8158 ( n10170 , n12202 , n2042 );
    or g8159 ( n6457 , n6614 , n6996 );
    not g8160 ( n2849 , n10395 );
    xnor g8161 ( n10721 , n4266 , n483 );
    or g8162 ( n7927 , n11407 , n4787 );
    or g8163 ( n5943 , n121 , n9118 );
    xnor g8164 ( n9371 , n454 , n1179 );
    or g8165 ( n12112 , n63 , n479 );
    xnor g8166 ( n4849 , n1508 , n4955 );
    or g8167 ( n4400 , n12295 , n10319 );
    xnor g8168 ( n7943 , n9498 , n6217 );
    and g8169 ( n4987 , n8680 , n222 );
    not g8170 ( n2822 , n11809 );
    xnor g8171 ( n12559 , n8497 , n10634 );
    and g8172 ( n5280 , n4042 , n1646 );
    or g8173 ( n2886 , n10550 , n6258 );
    and g8174 ( n12817 , n9174 , n9250 );
    not g8175 ( n10944 , n10850 );
    or g8176 ( n10530 , n10357 , n409 );
    not g8177 ( n11942 , n3014 );
    not g8178 ( n2579 , n12429 );
    and g8179 ( n3079 , n8378 , n12080 );
    or g8180 ( n7355 , n1320 , n9223 );
    or g8181 ( n4692 , n4465 , n8534 );
    not g8182 ( n5520 , n5758 );
    not g8183 ( n418 , n12622 );
    xnor g8184 ( n4845 , n914 , n6840 );
    xor g8185 ( n5938 , n1602 , n1612 );
    not g8186 ( n10929 , n9846 );
    xnor g8187 ( n3893 , n12199 , n13004 );
    and g8188 ( n293 , n2743 , n1620 );
    and g8189 ( n5967 , n3006 , n5729 );
    not g8190 ( n8458 , n12614 );
    xnor g8191 ( n3261 , n6016 , n8782 );
    or g8192 ( n4391 , n10877 , n4936 );
    not g8193 ( n1893 , n2882 );
    or g8194 ( n2413 , n4171 , n10516 );
    xnor g8195 ( n12827 , n2177 , n7571 );
    and g8196 ( n12428 , n5420 , n10980 );
    and g8197 ( n11743 , n2409 , n12026 );
    not g8198 ( n3429 , n13188 );
    nor g8199 ( n4924 , n10745 , n5457 );
    xnor g8200 ( n6222 , n5016 , n1238 );
    xnor g8201 ( n12852 , n4978 , n5236 );
    and g8202 ( n9707 , n3311 , n13058 );
    or g8203 ( n3621 , n6629 , n12188 );
    xnor g8204 ( n3150 , n4934 , n23 );
    nor g8205 ( n3857 , n1060 , n5860 );
    not g8206 ( n4256 , n1836 );
    and g8207 ( n1850 , n5009 , n7632 );
    not g8208 ( n10696 , n411 );
    xnor g8209 ( n8311 , n6744 , n5263 );
    not g8210 ( n2045 , n10751 );
    or g8211 ( n3627 , n11449 , n12847 );
    not g8212 ( n7481 , n4708 );
    or g8213 ( n9474 , n7068 , n2544 );
    xnor g8214 ( n5083 , n7418 , n3015 );
    xnor g8215 ( n12603 , n3695 , n4774 );
    or g8216 ( n6805 , n10045 , n2675 );
    not g8217 ( n9378 , n12850 );
    nor g8218 ( n3934 , n7368 , n11916 );
    not g8219 ( n6883 , n10606 );
    not g8220 ( n1191 , n1231 );
    xnor g8221 ( n5794 , n12479 , n2655 );
    or g8222 ( n7876 , n9112 , n2671 );
    or g8223 ( n5407 , n4366 , n2970 );
    xnor g8224 ( n11991 , n5207 , n1708 );
    not g8225 ( n5040 , n6826 );
    not g8226 ( n5521 , n11030 );
    or g8227 ( n1791 , n2940 , n11756 );
    or g8228 ( n4489 , n10798 , n6404 );
    xnor g8229 ( n7209 , n8517 , n6324 );
    or g8230 ( n6717 , n10137 , n8268 );
    and g8231 ( n1678 , n4701 , n10507 );
    not g8232 ( n7825 , n9093 );
    or g8233 ( n10660 , n10266 , n1695 );
    xnor g8234 ( n13205 , n11716 , n873 );
    nor g8235 ( n9851 , n6001 , n10866 );
    or g8236 ( n3156 , n5163 , n3981 );
    and g8237 ( n7060 , n8659 , n2153 );
    not g8238 ( n11165 , n5311 );
    or g8239 ( n2107 , n2296 , n2387 );
    xnor g8240 ( n1780 , n4417 , n12156 );
    and g8241 ( n9347 , n11509 , n1254 );
    xnor g8242 ( n7653 , n1169 , n10401 );
    or g8243 ( n12161 , n12109 , n206 );
    not g8244 ( n7567 , n11416 );
    nor g8245 ( n9759 , n13104 , n8566 );
    xnor g8246 ( n12546 , n8914 , n12231 );
    nor g8247 ( n7245 , n9347 , n13030 );
    xnor g8248 ( n11715 , n649 , n5691 );
    not g8249 ( n11002 , n9401 );
    not g8250 ( n9257 , n7772 );
    and g8251 ( n9390 , n11365 , n6531 );
    and g8252 ( n1627 , n4583 , n2925 );
    nor g8253 ( n225 , n11026 , n661 );
    and g8254 ( n13204 , n2613 , n12233 );
    nor g8255 ( n5567 , n5872 , n1170 );
    or g8256 ( n12336 , n9794 , n9681 );
    and g8257 ( n8331 , n8875 , n8491 );
    and g8258 ( n12975 , n5206 , n9789 );
    not g8259 ( n6166 , n11030 );
    xor g8260 ( n9236 , n4278 , n1879 );
    and g8261 ( n12415 , n2479 , n8292 );
    or g8262 ( n10429 , n2487 , n9075 );
    or g8263 ( n12270 , n6220 , n8225 );
    not g8264 ( n4841 , n9824 );
    or g8265 ( n8200 , n6231 , n5797 );
    or g8266 ( n3424 , n109 , n4052 );
    or g8267 ( n475 , n1893 , n206 );
    or g8268 ( n9670 , n98 , n10286 );
    not g8269 ( n9601 , n4423 );
    or g8270 ( n1800 , n8837 , n5100 );
    and g8271 ( n167 , n9330 , n11357 );
    or g8272 ( n720 , n785 , n4373 );
    or g8273 ( n3022 , n10412 , n5262 );
    nor g8274 ( n6053 , n13024 , n6887 );
    xnor g8275 ( n7423 , n10546 , n2277 );
    not g8276 ( n9019 , n1916 );
    or g8277 ( n6172 , n11781 , n8505 );
    not g8278 ( n10792 , n6409 );
    nor g8279 ( n2125 , n819 , n2324 );
    not g8280 ( n11212 , n7974 );
    or g8281 ( n12829 , n10830 , n7530 );
    or g8282 ( n82 , n8645 , n3981 );
    and g8283 ( n2611 , n8576 , n8825 );
    or g8284 ( n2444 , n1571 , n11668 );
    or g8285 ( n11558 , n11400 , n111 );
    xnor g8286 ( n7896 , n6382 , n5183 );
    and g8287 ( n1171 , n11132 , n1854 );
    or g8288 ( n6349 , n7805 , n11144 );
    not g8289 ( n12203 , n8468 );
    xnor g8290 ( n6277 , n5563 , n1118 );
    not g8291 ( n3091 , n2376 );
    and g8292 ( n925 , n4846 , n7678 );
    xnor g8293 ( n7449 , n5091 , n907 );
    xnor g8294 ( n8192 , n4445 , n6970 );
    xnor g8295 ( n8407 , n8385 , n3406 );
    xnor g8296 ( n7509 , n13053 , n1851 );
    and g8297 ( n2562 , n7557 , n3430 );
    or g8298 ( n6279 , n13106 , n6963 );
    or g8299 ( n4907 , n2118 , n4230 );
    or g8300 ( n11874 , n1323 , n13238 );
    or g8301 ( n2916 , n3026 , n13209 );
    not g8302 ( n2572 , n10744 );
    not g8303 ( n10830 , n8163 );
    not g8304 ( n12544 , n7428 );
    not g8305 ( n5968 , n11574 );
    and g8306 ( n7585 , n10041 , n11741 );
    or g8307 ( n1078 , n821 , n10904 );
    or g8308 ( n8926 , n7930 , n7935 );
    xnor g8309 ( n2979 , n2091 , n5580 );
    and g8310 ( n6834 , n3313 , n14 );
    xnor g8311 ( n8886 , n5250 , n11345 );
    xnor g8312 ( n11955 , n9254 , n5635 );
    or g8313 ( n12393 , n8325 , n12695 );
    xor g8314 ( n12863 , n9891 , n4997 );
    or g8315 ( n13103 , n1688 , n10871 );
    xnor g8316 ( n3090 , n3563 , n12460 );
    not g8317 ( n2711 , n11109 );
    not g8318 ( n11933 , n2341 );
    and g8319 ( n3821 , n319 , n13145 );
    or g8320 ( n5590 , n4132 , n7723 );
    nor g8321 ( n3759 , n3042 , n12403 );
    and g8322 ( n13189 , n9724 , n11956 );
    not g8323 ( n12620 , n11181 );
    and g8324 ( n4503 , n12017 , n2474 );
    xnor g8325 ( n1723 , n6948 , n4395 );
    and g8326 ( n2198 , n3178 , n834 );
    xnor g8327 ( n10942 , n9624 , n5710 );
    not g8328 ( n8384 , n4713 );
    and g8329 ( n3136 , n9345 , n4003 );
    or g8330 ( n2003 , n5321 , n1013 );
    xnor g8331 ( n11584 , n59 , n12209 );
    or g8332 ( n2563 , n8143 , n12328 );
    not g8333 ( n6580 , n6632 );
    or g8334 ( n11557 , n11237 , n8494 );
    or g8335 ( n4468 , n713 , n8319 );
    xnor g8336 ( n7274 , n10653 , n7397 );
    nor g8337 ( n5525 , n4896 , n7910 );
    not g8338 ( n93 , n7161 );
    nor g8339 ( n3668 , n9960 , n9393 );
    or g8340 ( n4153 , n2148 , n2133 );
    and g8341 ( n13091 , n5122 , n35 );
    and g8342 ( n3035 , n5586 , n2498 );
    or g8343 ( n9614 , n7966 , n177 );
    or g8344 ( n13243 , n5347 , n5373 );
    not g8345 ( n96 , n9039 );
    and g8346 ( n10876 , n2691 , n8363 );
    or g8347 ( n8266 , n1783 , n2757 );
    nor g8348 ( n7207 , n2987 , n2822 );
    or g8349 ( n13010 , n5704 , n10194 );
    or g8350 ( n6374 , n12212 , n3379 );
    xnor g8351 ( n1617 , n7064 , n11317 );
    xnor g8352 ( n5776 , n1722 , n12103 );
    or g8353 ( n7139 , n575 , n12870 );
    or g8354 ( n8917 , n5048 , n8702 );
    and g8355 ( n3003 , n11893 , n11705 );
    and g8356 ( n5914 , n7518 , n7112 );
    or g8357 ( n2687 , n12178 , n7840 );
    or g8358 ( n6135 , n2312 , n7820 );
    and g8359 ( n8657 , n5055 , n5593 );
    nor g8360 ( n4932 , n6757 , n11000 );
    and g8361 ( n10824 , n3595 , n9109 );
    and g8362 ( n634 , n1237 , n3216 );
    or g8363 ( n11996 , n9527 , n4469 );
    xnor g8364 ( n2137 , n4831 , n13034 );
    and g8365 ( n10325 , n10989 , n1226 );
    or g8366 ( n6676 , n6347 , n12377 );
    xnor g8367 ( n10828 , n8584 , n4119 );
    xnor g8368 ( n12238 , n310 , n6503 );
    xnor g8369 ( n1852 , n9695 , n8305 );
    and g8370 ( n7378 , n4516 , n5121 );
    or g8371 ( n11917 , n12834 , n7950 );
    or g8372 ( n2901 , n4566 , n8719 );
    or g8373 ( n6157 , n7564 , n11415 );
    not g8374 ( n5634 , n1084 );
    and g8375 ( n10867 , n3239 , n3037 );
    and g8376 ( n11146 , n9969 , n7732 );
    xnor g8377 ( n1604 , n12076 , n13162 );
    nor g8378 ( n7466 , n7250 , n1822 );
    and g8379 ( n9787 , n4619 , n5288 );
    xnor g8380 ( n6020 , n9094 , n431 );
    and g8381 ( n8521 , n3870 , n5584 );
    and g8382 ( n3576 , n7418 , n11744 );
    or g8383 ( n3101 , n1621 , n8534 );
    and g8384 ( n7734 , n4288 , n10503 );
    or g8385 ( n6612 , n1868 , n2465 );
    and g8386 ( n3485 , n940 , n568 );
    or g8387 ( n1539 , n5857 , n6177 );
    buf g8388 ( n1026 , n8160 );
    not g8389 ( n13148 , n8183 );
    and g8390 ( n7697 , n9639 , n9168 );
    xnor g8391 ( n10333 , n1163 , n5022 );
    or g8392 ( n4215 , n3940 , n8038 );
    xnor g8393 ( n10934 , n920 , n11282 );
    nor g8394 ( n2817 , n2350 , n1073 );
    nor g8395 ( n6915 , n1393 , n7708 );
    and g8396 ( n6958 , n11719 , n8158 );
    or g8397 ( n6291 , n12806 , n2589 );
    xnor g8398 ( n6071 , n2285 , n5304 );
    and g8399 ( n13225 , n5032 , n6426 );
    xnor g8400 ( n1391 , n387 , n10887 );
    not g8401 ( n10221 , n6794 );
    or g8402 ( n12230 , n12023 , n3698 );
    xnor g8403 ( n8258 , n7503 , n3794 );
    and g8404 ( n10800 , n937 , n3769 );
    or g8405 ( n880 , n7661 , n11668 );
    xnor g8406 ( n7280 , n10048 , n12842 );
    xnor g8407 ( n12739 , n6526 , n8066 );
    or g8408 ( n5829 , n7607 , n3501 );
    not g8409 ( n12617 , n3832 );
    or g8410 ( n2173 , n7167 , n12657 );
    xnor g8411 ( n9556 , n5335 , n3453 );
    not g8412 ( n278 , n8714 );
    or g8413 ( n9445 , n8243 , n11267 );
    and g8414 ( n8649 , n351 , n9764 );
    or g8415 ( n3265 , n9711 , n1463 );
    and g8416 ( n12143 , n6515 , n2393 );
    not g8417 ( n12595 , n9666 );
    and g8418 ( n5307 , n3995 , n9899 );
    nor g8419 ( n12896 , n1617 , n5596 );
    xnor g8420 ( n8557 , n12883 , n8441 );
    and g8421 ( n4505 , n6492 , n11464 );
    or g8422 ( n4668 , n114 , n121 );
    xnor g8423 ( n3262 , n1361 , n4849 );
    and g8424 ( n5716 , n8926 , n5736 );
    or g8425 ( n7190 , n710 , n11500 );
    xnor g8426 ( n580 , n8112 , n7940 );
    xnor g8427 ( n10121 , n8127 , n9298 );
    not g8428 ( n8173 , n12284 );
    not g8429 ( n1447 , n3076 );
    xnor g8430 ( n12028 , n4389 , n4746 );
    or g8431 ( n2973 , n829 , n5242 );
    or g8432 ( n9332 , n3013 , n2398 );
    nor g8433 ( n13237 , n7697 , n11172 );
    or g8434 ( n884 , n3096 , n12383 );
    or g8435 ( n10093 , n3584 , n376 );
    not g8436 ( n12778 , n7882 );
    and g8437 ( n7898 , n4653 , n2514 );
    xnor g8438 ( n6713 , n3385 , n6485 );
    not g8439 ( n10345 , n1148 );
    xnor g8440 ( n11129 , n2754 , n11458 );
    or g8441 ( n11481 , n740 , n4847 );
    or g8442 ( n524 , n5788 , n12811 );
    or g8443 ( n11954 , n445 , n121 );
    not g8444 ( n584 , n2771 );
    or g8445 ( n6669 , n1571 , n13086 );
    or g8446 ( n2740 , n3005 , n13017 );
    xnor g8447 ( n6498 , n8604 , n11030 );
    or g8448 ( n4494 , n6371 , n10071 );
    or g8449 ( n6856 , n12431 , n8385 );
    or g8450 ( n3385 , n1152 , n9195 );
    xnor g8451 ( n5635 , n2532 , n8140 );
    not g8452 ( n12082 , n32 );
    not g8453 ( n11333 , n772 );
    xnor g8454 ( n6445 , n8009 , n6628 );
    not g8455 ( n6293 , n2771 );
    and g8456 ( n1064 , n937 , n8233 );
    or g8457 ( n5007 , n10641 , n6635 );
    not g8458 ( n11914 , n5012 );
    or g8459 ( n11701 , n2546 , n8076 );
    not g8460 ( n7930 , n3085 );
    nor g8461 ( n4270 , n12047 , n5346 );
    or g8462 ( n1932 , n11910 , n4490 );
    not g8463 ( n9005 , n7087 );
    not g8464 ( n5261 , n12912 );
    not g8465 ( n8514 , n2071 );
    not g8466 ( n12952 , n10544 );
    and g8467 ( n3046 , n2518 , n5331 );
    nor g8468 ( n6106 , n11637 , n2432 );
    and g8469 ( n12426 , n11373 , n8829 );
    or g8470 ( n9740 , n10066 , n6690 );
    nor g8471 ( n10617 , n1233 , n13213 );
    not g8472 ( n1289 , n2656 );
    xnor g8473 ( n2925 , n12167 , n11586 );
    xnor g8474 ( n8072 , n505 , n3377 );
    not g8475 ( n5899 , n11561 );
    not g8476 ( n4260 , n6920 );
    xnor g8477 ( n12142 , n8745 , n919 );
    not g8478 ( n7154 , n3567 );
    or g8479 ( n10304 , n2868 , n10350 );
    or g8480 ( n2091 , n542 , n6404 );
    and g8481 ( n4337 , n2122 , n7388 );
    xnor g8482 ( n6424 , n3775 , n3756 );
    or g8483 ( n12533 , n2449 , n2675 );
    not g8484 ( n5251 , n3226 );
    or g8485 ( n4823 , n12795 , n4453 );
    or g8486 ( n6214 , n2456 , n13233 );
    or g8487 ( n1379 , n10920 , n5497 );
    xnor g8488 ( n6440 , n4154 , n898 );
    not g8489 ( n3514 , n1038 );
    and g8490 ( n234 , n6299 , n8064 );
    and g8491 ( n7615 , n11080 , n10155 );
    or g8492 ( n4945 , n1873 , n12074 );
    xnor g8493 ( n2857 , n4436 , n642 );
    nor g8494 ( n1947 , n10211 , n3734 );
    xnor g8495 ( n6155 , n4742 , n11084 );
    not g8496 ( n8029 , n12520 );
    xnor g8497 ( n12740 , n12720 , n12175 );
    or g8498 ( n1206 , n5595 , n12388 );
    or g8499 ( n5965 , n956 , n12188 );
    xnor g8500 ( n11117 , n1319 , n957 );
    and g8501 ( n6684 , n4364 , n12165 );
    not g8502 ( n2657 , n5920 );
    not g8503 ( n6133 , n4335 );
    or g8504 ( n9967 , n10929 , n6635 );
    xnor g8505 ( n10881 , n3753 , n6819 );
    xnor g8506 ( n5942 , n7984 , n12261 );
    xnor g8507 ( n8821 , n8474 , n1827 );
    or g8508 ( n6517 , n44 , n4947 );
    nor g8509 ( n9594 , n6473 , n10694 );
    xnor g8510 ( n9667 , n7931 , n915 );
    xnor g8511 ( n2381 , n3631 , n10841 );
    and g8512 ( n12356 , n2605 , n5245 );
    xnor g8513 ( n10992 , n1658 , n7233 );
    and g8514 ( n2311 , n1740 , n9881 );
    not g8515 ( n10017 , n5969 );
    not g8516 ( n10814 , n13060 );
    or g8517 ( n4605 , n9625 , n1767 );
    and g8518 ( n970 , n11236 , n6937 );
    not g8519 ( n12596 , n854 );
    xnor g8520 ( n7500 , n9996 , n1721 );
    or g8521 ( n454 , n3972 , n8534 );
    not g8522 ( n13170 , n3085 );
    and g8523 ( n7923 , n4885 , n585 );
    xnor g8524 ( n1217 , n8771 , n3842 );
    not g8525 ( n12241 , n6009 );
    not g8526 ( n8306 , n9906 );
    xnor g8527 ( n4777 , n4449 , n9077 );
    or g8528 ( n6911 , n4387 , n726 );
    not g8529 ( n9710 , n7208 );
    xnor g8530 ( n6296 , n12386 , n6261 );
    xnor g8531 ( n9348 , n3684 , n9189 );
    or g8532 ( n3171 , n795 , n12930 );
    and g8533 ( n5768 , n10770 , n6392 );
    nor g8534 ( n8103 , n4617 , n5162 );
    xor g8535 ( n11140 , n1344 , n3950 );
    or g8536 ( n6345 , n5176 , n3640 );
    or g8537 ( n6401 , n5841 , n542 );
    xnor g8538 ( n11930 , n2555 , n11479 );
    or g8539 ( n7235 , n11723 , n2893 );
    xnor g8540 ( n8794 , n10472 , n12148 );
    not g8541 ( n10474 , n11324 );
    and g8542 ( n3177 , n13068 , n7361 );
    or g8543 ( n4725 , n10023 , n11042 );
    or g8544 ( n9299 , n1989 , n7805 );
    xnor g8545 ( n4549 , n3592 , n11811 );
    not g8546 ( n9784 , n1364 );
    xnor g8547 ( n8923 , n3441 , n3277 );
    or g8548 ( n8372 , n9421 , n6732 );
    and g8549 ( n11866 , n5801 , n10408 );
    or g8550 ( n7350 , n2733 , n1272 );
    and g8551 ( n9909 , n24 , n1593 );
    or g8552 ( n13098 , n3646 , n6635 );
    or g8553 ( n10495 , n8518 , n11750 );
    xnor g8554 ( n4311 , n729 , n1071 );
    or g8555 ( n12227 , n7363 , n10 );
    or g8556 ( n5786 , n10814 , n2675 );
    xnor g8557 ( n9446 , n6483 , n8991 );
    or g8558 ( n8815 , n8529 , n8702 );
    xnor g8559 ( n8686 , n2283 , n3762 );
    or g8560 ( n6391 , n8390 , n2076 );
    xnor g8561 ( n6104 , n9320 , n10449 );
    xnor g8562 ( n7617 , n67 , n5587 );
    xnor g8563 ( n2317 , n6468 , n8599 );
    or g8564 ( n1874 , n2279 , n9126 );
    or g8565 ( n5558 , n2346 , n12695 );
    not g8566 ( n5992 , n10738 );
    xnor g8567 ( n11834 , n1642 , n12280 );
    xor g8568 ( n9316 , n2720 , n12645 );
    not g8569 ( n9311 , n1405 );
    xnor g8570 ( n5000 , n8710 , n10933 );
    or g8571 ( n13024 , n737 , n8702 );
    xnor g8572 ( n8735 , n5321 , n6351 );
    or g8573 ( n6465 , n3516 , n3126 );
    or g8574 ( n4923 , n10546 , n4667 );
    or g8575 ( n11718 , n3222 , n4925 );
    and g8576 ( n786 , n4758 , n6420 );
    not g8577 ( n9453 , n12842 );
    and g8578 ( n11655 , n12969 , n12686 );
    not g8579 ( n2660 , n8867 );
    not g8580 ( n13168 , n4330 );
    and g8581 ( n270 , n3241 , n601 );
    nor g8582 ( n4115 , n1343 , n11047 );
    nor g8583 ( n2706 , n3879 , n4115 );
    not g8584 ( n13021 , n4074 );
    and g8585 ( n10838 , n10762 , n1675 );
    nor g8586 ( n1853 , n13162 , n3883 );
    not g8587 ( n9154 , n8522 );
    and g8588 ( n738 , n9029 , n7679 );
    xnor g8589 ( n2588 , n12161 , n12455 );
    not g8590 ( n4396 , n4698 );
    or g8591 ( n10749 , n12448 , n7838 );
    nor g8592 ( n4127 , n5499 , n5363 );
    or g8593 ( n8708 , n6268 , n4358 );
    and g8594 ( n186 , n9792 , n4995 );
    and g8595 ( n13053 , n8508 , n13235 );
    xnor g8596 ( n9680 , n12928 , n2247 );
    not g8597 ( n3111 , n2431 );
    not g8598 ( n8234 , n10763 );
    xnor g8599 ( n1097 , n7716 , n7103 );
    xnor g8600 ( n4092 , n1968 , n9572 );
    nor g8601 ( n3331 , n7286 , n8798 );
    or g8602 ( n286 , n3767 , n11257 );
    xnor g8603 ( n11534 , n5199 , n2039 );
    or g8604 ( n10670 , n6289 , n1614 );
    xnor g8605 ( n611 , n610 , n1275 );
    or g8606 ( n7056 , n3268 , n6270 );
    nor g8607 ( n8968 , n120 , n12028 );
    or g8608 ( n7573 , n9627 , n12195 );
    not g8609 ( n7356 , n9750 );
    not g8610 ( n11121 , n691 );
    xnor g8611 ( n8395 , n1385 , n10554 );
    xnor g8612 ( n11802 , n13217 , n6550 );
    not g8613 ( n8510 , n817 );
    xnor g8614 ( n446 , n5075 , n1430 );
    or g8615 ( n5518 , n4473 , n7935 );
    or g8616 ( n1914 , n3273 , n1780 );
    xnor g8617 ( n658 , n2259 , n949 );
    and g8618 ( n12302 , n1933 , n9407 );
    or g8619 ( n6205 , n1783 , n2958 );
    not g8620 ( n6183 , n4591 );
    nor g8621 ( n512 , n10645 , n7583 );
    and g8622 ( n3285 , n12598 , n1003 );
    not g8623 ( n4515 , n9475 );
    xnor g8624 ( n11656 , n1805 , n8694 );
    and g8625 ( n10455 , n3729 , n11006 );
    or g8626 ( n7498 , n596 , n1825 );
    xnor g8627 ( n2984 , n3009 , n10488 );
    or g8628 ( n8412 , n11858 , n5873 );
    xnor g8629 ( n6334 , n10335 , n3966 );
    xnor g8630 ( n6548 , n3188 , n4002 );
    or g8631 ( n13207 , n5360 , n6601 );
    not g8632 ( n10903 , n4623 );
    nor g8633 ( n7826 , n5255 , n10436 );
    and g8634 ( n9416 , n9374 , n3389 );
    nor g8635 ( n12147 , n1003 , n12598 );
    or g8636 ( n11127 , n4793 , n10165 );
    not g8637 ( n4187 , n5827 );
    xnor g8638 ( n4592 , n12532 , n1330 );
    and g8639 ( n6513 , n11975 , n8408 );
    or g8640 ( n8356 , n6689 , n10049 );
    or g8641 ( n11661 , n13 , n2127 );
    xnor g8642 ( n8830 , n329 , n8479 );
    xor g8643 ( n9663 , n2791 , n4138 );
    and g8644 ( n2097 , n2205 , n5095 );
    and g8645 ( n3358 , n6808 , n1289 );
    and g8646 ( n1268 , n10768 , n10154 );
    and g8647 ( n2154 , n5872 , n1170 );
    or g8648 ( n13215 , n10895 , n9014 );
    and g8649 ( n12077 , n11060 , n5633 );
    xnor g8650 ( n8596 , n11903 , n5765 );
    xnor g8651 ( n6798 , n12805 , n4 );
    nor g8652 ( n3942 , n3230 , n10486 );
    xnor g8653 ( n6395 , n277 , n7050 );
    or g8654 ( n8316 , n9668 , n5242 );
    xor g8655 ( n10797 , n13011 , n13219 );
    and g8656 ( n2099 , n7037 , n5337 );
    or g8657 ( n7348 , n12109 , n6732 );
    or g8658 ( n12374 , n3243 , n206 );
    or g8659 ( n9395 , n8576 , n8825 );
    xnor g8660 ( n10546 , n3722 , n3903 );
    nor g8661 ( n7581 , n13152 , n5950 );
    and g8662 ( n7164 , n12722 , n2134 );
    or g8663 ( n1699 , n11680 , n2542 );
    and g8664 ( n3399 , n8892 , n4522 );
    not g8665 ( n2455 , n1774 );
    xnor g8666 ( n11289 , n4853 , n12337 );
    or g8667 ( n6877 , n4584 , n7723 );
    xnor g8668 ( n5632 , n1865 , n7922 );
    xnor g8669 ( n1340 , n12855 , n1670 );
    nor g8670 ( n9863 , n3471 , n11287 );
    or g8671 ( n3397 , n10830 , n6265 );
    or g8672 ( n8105 , n8759 , n9075 );
    or g8673 ( n243 , n9581 , n8348 );
    or g8674 ( n3922 , n1284 , n10885 );
    and g8675 ( n9714 , n9477 , n12611 );
    or g8676 ( n6137 , n7505 , n8278 );
    and g8677 ( n2514 , n4780 , n10623 );
    and g8678 ( n8218 , n2211 , n7772 );
    or g8679 ( n12098 , n7251 , n9229 );
    xnor g8680 ( n1411 , n11297 , n4100 );
    xnor g8681 ( n11057 , n2377 , n2147 );
    not g8682 ( n4179 , n411 );
    xnor g8683 ( n3610 , n11625 , n12266 );
    or g8684 ( n8993 , n12785 , n12900 );
    or g8685 ( n3473 , n6280 , n742 );
    or g8686 ( n12290 , n1113 , n8030 );
    or g8687 ( n9387 , n13181 , n9444 );
    or g8688 ( n1472 , n1035 , n8702 );
    or g8689 ( n4848 , n10223 , n2082 );
    and g8690 ( n10403 , n12105 , n10129 );
    not g8691 ( n11853 , n11968 );
    and g8692 ( n12941 , n11611 , n3985 );
    or g8693 ( n5602 , n5342 , n2609 );
    xnor g8694 ( n8564 , n390 , n6328 );
    xnor g8695 ( n1653 , n5757 , n10119 );
    or g8696 ( n1715 , n0 , n8348 );
    not g8697 ( n4333 , n851 );
    xnor g8698 ( n10647 , n2780 , n7314 );
    xnor g8699 ( n9260 , n5469 , n8470 );
    and g8700 ( n3739 , n8466 , n5536 );
    xnor g8701 ( n2205 , n10662 , n8303 );
    or g8702 ( n1739 , n12619 , n5344 );
    nor g8703 ( n6272 , n6363 , n6582 );
    not g8704 ( n10131 , n12845 );
    not g8705 ( n4584 , n11350 );
    xnor g8706 ( n7849 , n11188 , n7387 );
    not g8707 ( n6129 , n443 );
    not g8708 ( n2545 , n12267 );
    xnor g8709 ( n7051 , n11275 , n8459 );
    xnor g8710 ( n7687 , n3327 , n10729 );
    and g8711 ( n2729 , n9842 , n4275 );
    xnor g8712 ( n4331 , n2721 , n9343 );
    or g8713 ( n11187 , n4166 , n7530 );
    not g8714 ( n12889 , n11290 );
    xnor g8715 ( n10394 , n3174 , n10136 );
    not g8716 ( n10117 , n12005 );
    not g8717 ( n12330 , n11715 );
    not g8718 ( n11815 , n3378 );
    not g8719 ( n1089 , n3669 );
    xor g8720 ( n3411 , n6174 , n4003 );
    or g8721 ( n7694 , n6557 , n13108 );
    nor g8722 ( n7405 , n11938 , n6592 );
    not g8723 ( n6250 , n12651 );
    not g8724 ( n8858 , n5981 );
    xnor g8725 ( n2233 , n5160 , n6510 );
    not g8726 ( n583 , n962 );
    xnor g8727 ( n12201 , n13138 , n564 );
    xnor g8728 ( n5419 , n12866 , n9214 );
    nor g8729 ( n7870 , n5113 , n9133 );
    nor g8730 ( n12127 , n3642 , n11913 );
    xnor g8731 ( n8172 , n8543 , n582 );
    and g8732 ( n9608 , n2786 , n8972 );
    xnor g8733 ( n2654 , n5095 , n2917 );
    buf g8734 ( n10933 , n10301 );
    xnor g8735 ( n9073 , n8507 , n9852 );
    or g8736 ( n4617 , n8006 , n6178 );
    and g8737 ( n8152 , n1200 , n7645 );
    and g8738 ( n3276 , n9451 , n5366 );
    or g8739 ( n5120 , n6755 , n2556 );
    nor g8740 ( n7381 , n12147 , n4733 );
    not g8741 ( n7555 , n3303 );
    or g8742 ( n9244 , n12777 , n1034 );
    xnor g8743 ( n8583 , n11027 , n11693 );
    xnor g8744 ( n5912 , n739 , n11488 );
    and g8745 ( n2408 , n10208 , n8683 );
    xnor g8746 ( n1167 , n8512 , n7658 );
    xnor g8747 ( n1937 , n491 , n9680 );
    not g8748 ( n6120 , n9893 );
    xnor g8749 ( n8791 , n3785 , n12185 );
    not g8750 ( n3185 , n11058 );
    not g8751 ( n6238 , n342 );
    xnor g8752 ( n12499 , n10572 , n2703 );
    or g8753 ( n12843 , n1194 , n206 );
    or g8754 ( n5601 , n12102 , n2197 );
    and g8755 ( n1894 , n4811 , n8787 );
    and g8756 ( n10028 , n8355 , n2663 );
    nor g8757 ( n13033 , n2644 , n2803 );
    or g8758 ( n1585 , n45 , n9075 );
    xnor g8759 ( n268 , n7564 , n11415 );
    xnor g8760 ( n11836 , n5293 , n4409 );
    not g8761 ( n2504 , n12965 );
    and g8762 ( n7844 , n11175 , n6612 );
    or g8763 ( n9700 , n8562 , n1985 );
    not g8764 ( n7908 , n10538 );
    and g8765 ( n1180 , n8391 , n5762 );
    or g8766 ( n12855 , n12483 , n10573 );
    xor g8767 ( n7323 , n4293 , n7877 );
    and g8768 ( n253 , n9434 , n3466 );
    or g8769 ( n11266 , n3225 , n4936 );
    and g8770 ( n9989 , n7072 , n12243 );
    or g8771 ( n3907 , n8275 , n11712 );
    or g8772 ( n2268 , n2944 , n7733 );
    and g8773 ( n5710 , n5511 , n7913 );
    or g8774 ( n5922 , n6751 , n5076 );
    or g8775 ( n4663 , n6769 , n2675 );
    and g8776 ( n10173 , n9699 , n1230 );
    not g8777 ( n11745 , n4086 );
    not g8778 ( n6086 , n9747 );
    and g8779 ( n3097 , n5214 , n9669 );
    xnor g8780 ( n12810 , n568 , n7246 );
    or g8781 ( n9485 , n4750 , n2460 );
    not g8782 ( n12169 , n1494 );
    xnor g8783 ( n2241 , n5908 , n11469 );
    xnor g8784 ( n7138 , n3291 , n9198 );
    or g8785 ( n10324 , n11680 , n11078 );
    or g8786 ( n7836 , n2861 , n1026 );
    buf g8787 ( n12501 , n9257 );
    or g8788 ( n9780 , n6447 , n5987 );
    and g8789 ( n12830 , n8446 , n6413 );
    not g8790 ( n12758 , n6023 );
    or g8791 ( n508 , n4531 , n12909 );
    or g8792 ( n4943 , n10911 , n2181 );
    and g8793 ( n9078 , n1892 , n1679 );
    xnor g8794 ( n5362 , n1859 , n7816 );
    or g8795 ( n8337 , n9436 , n3411 );
    xnor g8796 ( n13232 , n1427 , n5591 );
    not g8797 ( n12403 , n10207 );
    and g8798 ( n7080 , n11015 , n7955 );
    xnor g8799 ( n7745 , n6170 , n11181 );
    nor g8800 ( n514 , n1625 , n1829 );
    and g8801 ( n2379 , n4396 , n6893 );
    not g8802 ( n8759 , n6826 );
    and g8803 ( n2249 , n8685 , n3780 );
    and g8804 ( n7250 , n504 , n7356 );
    xor g8805 ( n2354 , n11457 , n5991 );
    and g8806 ( n2627 , n4497 , n8619 );
    not g8807 ( n3928 , n11734 );
    not g8808 ( n8640 , n7529 );
    and g8809 ( n13089 , n10069 , n5419 );
    not g8810 ( n3531 , n510 );
    and g8811 ( n8914 , n8985 , n6585 );
    or g8812 ( n11674 , n10898 , n12695 );
    not g8813 ( n9919 , n4335 );
    not g8814 ( n12115 , n10497 );
    xnor g8815 ( n4281 , n4457 , n4925 );
    or g8816 ( n7104 , n1893 , n1570 );
    or g8817 ( n3280 , n7745 , n418 );
    xnor g8818 ( n12106 , n6812 , n6548 );
    not g8819 ( n13026 , n12263 );
    or g8820 ( n1775 , n8646 , n6404 );
    or g8821 ( n3159 , n121 , n2890 );
    or g8822 ( n11849 , n1835 , n8509 );
    or g8823 ( n5760 , n1700 , n11045 );
    or g8824 ( n4754 , n6743 , n8702 );
    and g8825 ( n4809 , n12039 , n8245 );
    xnor g8826 ( n9156 , n1760 , n8451 );
    or g8827 ( n7299 , n1601 , n10508 );
    xnor g8828 ( n10295 , n5846 , n5597 );
    nor g8829 ( n10420 , n6342 , n4093 );
    or g8830 ( n3700 , n8428 , n8530 );
    xnor g8831 ( n8765 , n9845 , n7800 );
    or g8832 ( n6167 , n12629 , n6732 );
    xnor g8833 ( n7536 , n95 , n4579 );
    and g8834 ( n9086 , n11570 , n4239 );
    or g8835 ( n10199 , n4628 , n12205 );
    and g8836 ( n12932 , n9216 , n10606 );
    nor g8837 ( n6069 , n9837 , n7290 );
    not g8838 ( n2141 , n3631 );
    not g8839 ( n5990 , n8290 );
    or g8840 ( n372 , n1281 , n2672 );
    and g8841 ( n9565 , n1857 , n9096 );
    not g8842 ( n12914 , n4113 );
    and g8843 ( n1646 , n2592 , n497 );
    or g8844 ( n12728 , n11920 , n237 );
    not g8845 ( n8630 , n4325 );
    and g8846 ( n1958 , n10894 , n2503 );
    nor g8847 ( n12869 , n8157 , n9086 );
    not g8848 ( n1188 , n11222 );
    nor g8849 ( n7941 , n7045 , n4069 );
    xnor g8850 ( n8507 , n7654 , n8555 );
    and g8851 ( n5712 , n390 , n9439 );
    or g8852 ( n13234 , n5013 , n84 );
    xnor g8853 ( n2629 , n3136 , n587 );
    and g8854 ( n5340 , n5528 , n11377 );
    xnor g8855 ( n1950 , n2603 , n10224 );
    xnor g8856 ( n2953 , n5192 , n722 );
    nor g8857 ( n4049 , n7609 , n11924 );
    not g8858 ( n10471 , n12965 );
    or g8859 ( n7416 , n189 , n5875 );
    not g8860 ( n8392 , n10594 );
    nor g8861 ( n6545 , n12880 , n8478 );
    xnor g8862 ( n10815 , n247 , n7995 );
    and g8863 ( n8969 , n4837 , n6740 );
    or g8864 ( n4402 , n11567 , n7526 );
    xnor g8865 ( n10406 , n335 , n10349 );
    or g8866 ( n1424 , n3965 , n8941 );
    xnor g8867 ( n10839 , n3579 , n6998 );
    and g8868 ( n3008 , n11236 , n10408 );
    xnor g8869 ( n6307 , n10415 , n6415 );
    not g8870 ( n3437 , n10928 );
    nor g8871 ( n12706 , n7413 , n8220 );
    nor g8872 ( n13018 , n5625 , n9539 );
    xnor g8873 ( n3249 , n12819 , n7960 );
    and g8874 ( n11780 , n2018 , n411 );
    not g8875 ( n5148 , n10162 );
    or g8876 ( n9331 , n2639 , n2675 );
    xnor g8877 ( n6531 , n6888 , n4671 );
    xnor g8878 ( n2739 , n6363 , n2328 );
    and g8879 ( n5881 , n4660 , n6633 );
    and g8880 ( n1173 , n12578 , n7163 );
    xnor g8881 ( n964 , n3939 , n9006 );
    or g8882 ( n4984 , n891 , n1092 );
    xnor g8883 ( n12381 , n10867 , n10648 );
    xnor g8884 ( n2121 , n8750 , n12481 );
    xnor g8885 ( n2659 , n12091 , n9752 );
    xnor g8886 ( n6646 , n5030 , n11547 );
    xnor g8887 ( n5192 , n4699 , n13101 );
    and g8888 ( n3183 , n6790 , n10398 );
    and g8889 ( n2698 , n7534 , n7427 );
    nor g8890 ( n9811 , n4609 , n2461 );
    or g8891 ( n1015 , n1427 , n5591 );
    and g8892 ( n1467 , n2636 , n7815 );
    and g8893 ( n8684 , n3781 , n9485 );
    xnor g8894 ( n7978 , n3735 , n8484 );
    and g8895 ( n10175 , n9025 , n11374 );
    and g8896 ( n5344 , n252 , n10429 );
    xnor g8897 ( n246 , n4562 , n1384 );
    not g8898 ( n2446 , n7012 );
    or g8899 ( n5624 , n4657 , n1605 );
    or g8900 ( n12025 , n2228 , n12604 );
    or g8901 ( n1599 , n1438 , n479 );
    and g8902 ( n1738 , n10724 , n9880 );
    or g8903 ( n572 , n9723 , n12501 );
    not g8904 ( n12384 , n5068 );
    nor g8905 ( n4838 , n4920 , n6049 );
    not g8906 ( n5502 , n5477 );
    nor g8907 ( n4160 , n12276 , n5244 );
    and g8908 ( n8869 , n6977 , n5007 );
    xnor g8909 ( n9755 , n359 , n7905 );
    not g8910 ( n3800 , n5570 );
    not g8911 ( n906 , n7569 );
    not g8912 ( n10059 , n3815 );
    xnor g8913 ( n4138 , n7728 , n12956 );
    xnor g8914 ( n32 , n6212 , n6406 );
    not g8915 ( n3537 , n1198 );
    xor g8916 ( n2977 , n5248 , n1689 );
    xnor g8917 ( n10687 , n6080 , n3463 );
    not g8918 ( n3173 , n10482 );
    and g8919 ( n2051 , n1029 , n10252 );
    not g8920 ( n5163 , n1392 );
    not g8921 ( n1883 , n9915 );
    not g8922 ( n11514 , n4452 );
    xor g8923 ( n6823 , n10599 , n5117 );
    or g8924 ( n11983 , n11514 , n7430 );
    xnor g8925 ( n10082 , n47 , n1728 );
    and g8926 ( n9418 , n11020 , n2727 );
    xnor g8927 ( n5546 , n11719 , n5629 );
    not g8928 ( n8081 , n4395 );
    not g8929 ( n1389 , n246 );
    not g8930 ( n785 , n12408 );
    not g8931 ( n6942 , n7285 );
    and g8932 ( n503 , n3008 , n9005 );
    not g8933 ( n9888 , n2062 );
    or g8934 ( n10132 , n5588 , n4640 );
    and g8935 ( n11282 , n613 , n4137 );
    xnor g8936 ( n11949 , n1762 , n11003 );
    or g8937 ( n8717 , n4453 , n3225 );
    xnor g8938 ( n724 , n10873 , n4512 );
    or g8939 ( n6520 , n8020 , n10179 );
    not g8940 ( n4779 , n9230 );
    not g8941 ( n4063 , n9732 );
    and g8942 ( n2618 , n8033 , n2949 );
    and g8943 ( n5620 , n6524 , n5380 );
    xnor g8944 ( n10344 , n10064 , n12549 );
    and g8945 ( n5785 , n7683 , n4592 );
    or g8946 ( n7386 , n8966 , n9689 );
    xnor g8947 ( n11389 , n1278 , n2031 );
    xnor g8948 ( n3718 , n7794 , n9114 );
    or g8949 ( n12444 , n5146 , n2958 );
    or g8950 ( n693 , n5199 , n2039 );
    not g8951 ( n8613 , n12936 );
    or g8952 ( n11092 , n10439 , n7530 );
    xnor g8953 ( n7492 , n11776 , n3290 );
    nor g8954 ( n6720 , n5907 , n5785 );
    or g8955 ( n11710 , n3616 , n10179 );
    not g8956 ( n10182 , n1330 );
    or g8957 ( n5996 , n8609 , n9919 );
    and g8958 ( n10163 , n11777 , n10774 );
    or g8959 ( n4736 , n371 , n5186 );
    nor g8960 ( n5282 , n535 , n8274 );
    or g8961 ( n12349 , n12199 , n9582 );
    or g8962 ( n8207 , n1051 , n5076 );
    not g8963 ( n1296 , n3815 );
    or g8964 ( n1926 , n11212 , n8702 );
    or g8965 ( n5445 , n75 , n4936 );
    and g8966 ( n10 , n11768 , n7836 );
    not g8967 ( n12441 , n1636 );
    xnor g8968 ( n12079 , n11777 , n12761 );
    or g8969 ( n2601 , n2434 , n2036 );
    nor g8970 ( n9360 , n4681 , n1313 );
    or g8971 ( n11998 , n6699 , n6265 );
    nor g8972 ( n6554 , n2665 , n4759 );
    and g8973 ( n5173 , n6981 , n1020 );
    and g8974 ( n3312 , n673 , n366 );
    and g8975 ( n170 , n7350 , n4180 );
    and g8976 ( n13055 , n7213 , n8961 );
    and g8977 ( n6096 , n11557 , n3375 );
    or g8978 ( n9288 , n12122 , n6091 );
    not g8979 ( n9837 , n336 );
    or g8980 ( n5748 , n8778 , n1999 );
    and g8981 ( n1935 , n6219 , n6734 );
    or g8982 ( n12911 , n3225 , n6404 );
    or g8983 ( n8676 , n6810 , n10871 );
    and g8984 ( n4594 , n2018 , n13058 );
    not g8985 ( n10331 , n13064 );
    and g8986 ( n8066 , n12349 , n8444 );
    and g8987 ( n11173 , n1850 , n8882 );
    or g8988 ( n1647 , n4999 , n5652 );
    nor g8989 ( n1166 , n6712 , n6578 );
    xnor g8990 ( n1911 , n11024 , n3156 );
    xnor g8991 ( n5913 , n5228 , n3330 );
    and g8992 ( n10019 , n1431 , n10856 );
    or g8993 ( n11005 , n11929 , n9268 );
    or g8994 ( n10999 , n6063 , n1463 );
    and g8995 ( n7551 , n1305 , n747 );
    or g8996 ( n8726 , n7134 , n8247 );
    xnor g8997 ( n6647 , n5584 , n825 );
    xnor g8998 ( n11216 , n7836 , n11768 );
    and g8999 ( n9448 , n909 , n4805 );
    xnor g9000 ( n6619 , n5702 , n12201 );
    xnor g9001 ( n7802 , n8549 , n5804 );
    xor g9002 ( n7779 , n11559 , n8542 );
    nor g9003 ( n5225 , n9037 , n7599 );
    not g9004 ( n9286 , n7 );
    not g9005 ( n1919 , n8290 );
    or g9006 ( n2661 , n7741 , n9159 );
    or g9007 ( n11213 , n718 , n12862 );
    or g9008 ( n12168 , n5565 , n1144 );
    xnor g9009 ( n7359 , n13031 , n3073 );
    xnor g9010 ( n6747 , n8 , n4401 );
    or g9011 ( n9277 , n1325 , n3825 );
    not g9012 ( n5740 , n8139 );
    or g9013 ( n11571 , n7819 , n2449 );
    xnor g9014 ( n9560 , n10431 , n9299 );
    nor g9015 ( n6761 , n2518 , n5331 );
    xnor g9016 ( n8544 , n5185 , n9650 );
    xnor g9017 ( n2957 , n5072 , n9289 );
    or g9018 ( n6446 , n10411 , n11239 );
    and g9019 ( n2074 , n6447 , n5987 );
    not g9020 ( n6988 , n10657 );
    not g9021 ( n11864 , n3832 );
    and g9022 ( n1187 , n6180 , n1862 );
    xnor g9023 ( n8217 , n11464 , n11651 );
    or g9024 ( n4034 , n11094 , n4936 );
    xnor g9025 ( n2929 , n10630 , n2690 );
    or g9026 ( n5153 , n11648 , n8805 );
    or g9027 ( n7517 , n6749 , n2943 );
    xnor g9028 ( n11736 , n12312 , n12239 );
    xnor g9029 ( n10722 , n223 , n1590 );
    and g9030 ( n7873 , n8915 , n12012 );
    xnor g9031 ( n4897 , n9138 , n11254 );
    or g9032 ( n8565 , n12254 , n4230 );
    xnor g9033 ( n9530 , n13171 , n7536 );
    xnor g9034 ( n1870 , n2388 , n4186 );
    not g9035 ( n4499 , n5603 );
    xnor g9036 ( n5728 , n13196 , n4727 );
    and g9037 ( n3506 , n1328 , n6741 );
    or g9038 ( n12354 , n6173 , n4116 );
    not g9039 ( n8650 , n7725 );
    xnor g9040 ( n3594 , n5324 , n3074 );
    or g9041 ( n12773 , n9580 , n486 );
    and g9042 ( n5995 , n5449 , n5855 );
    or g9043 ( n593 , n10351 , n8448 );
    xnor g9044 ( n8124 , n9247 , n2979 );
    xnor g9045 ( n11719 , n6926 , n746 );
    or g9046 ( n5964 , n6901 , n11670 );
    or g9047 ( n10252 , n745 , n982 );
    xnor g9048 ( n4843 , n1932 , n7850 );
    xnor g9049 ( n10827 , n3708 , n5496 );
    not g9050 ( n12986 , n8520 );
    or g9051 ( n7545 , n6086 , n5076 );
    or g9052 ( n7921 , n7862 , n9861 );
    or g9053 ( n11096 , n2416 , n8348 );
    nor g9054 ( n12864 , n9878 , n3030 );
    and g9055 ( n5096 , n10147 , n2564 );
    xnor g9056 ( n7445 , n5431 , n4429 );
    and g9057 ( n1254 , n8183 , n854 );
    and g9058 ( n6901 , n8953 , n3880 );
    or g9059 ( n9384 , n10509 , n11928 );
    or g9060 ( n9600 , n5233 , n9579 );
    xnor g9061 ( n7726 , n3161 , n251 );
    or g9062 ( n8177 , n6492 , n11464 );
    not g9063 ( n3344 , n10162 );
    and g9064 ( n12670 , n12615 , n7667 );
    xnor g9065 ( n2119 , n4187 , n2216 );
    xnor g9066 ( n3152 , n6607 , n7116 );
    and g9067 ( n12087 , n2194 , n5109 );
    not g9068 ( n11548 , n9093 );
    or g9069 ( n6479 , n10798 , n10179 );
    and g9070 ( n4787 , n8264 , n10834 );
    or g9071 ( n8443 , n12894 , n2969 );
    xnor g9072 ( n3988 , n12652 , n10076 );
    xnor g9073 ( n6351 , n615 , n8386 );
    or g9074 ( n11228 , n3928 , n12501 );
    xnor g9075 ( n4882 , n3886 , n8899 );
    or g9076 ( n1630 , n2823 , n566 );
    or g9077 ( n8959 , n11761 , n6874 );
    nor g9078 ( n12223 , n5615 , n805 );
    xnor g9079 ( n11134 , n3006 , n5568 );
    xnor g9080 ( n12468 , n5616 , n5332 );
    xnor g9081 ( n6059 , n11203 , n3926 );
    or g9082 ( n2265 , n11084 , n3479 );
    or g9083 ( n10489 , n5923 , n8188 );
    not g9084 ( n8082 , n2295 );
    xnor g9085 ( n8283 , n2437 , n691 );
    xnor g9086 ( n6553 , n1450 , n703 );
    and g9087 ( n8996 , n3903 , n3722 );
    xnor g9088 ( n2736 , n2137 , n342 );
    or g9089 ( n5738 , n9019 , n8348 );
    and g9090 ( n7854 , n5671 , n4335 );
    and g9091 ( n5333 , n11745 , n1920 );
    and g9092 ( n1133 , n13127 , n452 );
    not g9093 ( n11614 , n6857 );
    not g9094 ( n13159 , n6818 );
    xnor g9095 ( n10055 , n9384 , n2401 );
    not g9096 ( n7945 , n12391 );
    or g9097 ( n5771 , n5544 , n3372 );
    xor g9098 ( n10150 , n2062 , n6394 );
    or g9099 ( n1400 , n11928 , n2958 );
    or g9100 ( n14 , n6672 , n1043 );
    and g9101 ( n8321 , n1997 , n4054 );
    and g9102 ( n11434 , n11324 , n12284 );
    xnor g9103 ( n5501 , n2536 , n982 );
    not g9104 ( n9675 , n353 );
    and g9105 ( n3286 , n629 , n5153 );
    xnor g9106 ( n901 , n7545 , n4276 );
    xnor g9107 ( n5549 , n2569 , n4590 );
    xnor g9108 ( n5137 , n3974 , n11906 );
    and g9109 ( n13032 , n1009 , n8296 );
    and g9110 ( n6478 , n9032 , n3235 );
    xnor g9111 ( n6624 , n9190 , n9503 );
    or g9112 ( n8185 , n9776 , n8587 );
    nor g9113 ( n8238 , n6513 , n2475 );
    xnor g9114 ( n6771 , n6310 , n9950 );
    xnor g9115 ( n296 , n12649 , n11983 );
    not g9116 ( n7942 , n2043 );
    nor g9117 ( n1124 , n5649 , n8695 );
    and g9118 ( n2655 , n10168 , n3832 );
    and g9119 ( n4286 , n3413 , n9708 );
    or g9120 ( n2833 , n3062 , n542 );
    and g9121 ( n4169 , n4133 , n11915 );
    or g9122 ( n5250 , n2688 , n6265 );
    xnor g9123 ( n5458 , n3683 , n9832 );
    and g9124 ( n5817 , n12077 , n5125 );
    xor g9125 ( n12321 , n9474 , n11854 );
    not g9126 ( n8383 , n2771 );
    not g9127 ( n1345 , n2758 );
    or g9128 ( n4365 , n304 , n10079 );
    and g9129 ( n5044 , n13075 , n2390 );
    not g9130 ( n11696 , n12560 );
    and g9131 ( n5848 , n6543 , n13187 );
    xnor g9132 ( n12121 , n8242 , n10209 );
    not g9133 ( n991 , n12306 );
    nor g9134 ( n9865 , n8238 , n725 );
    and g9135 ( n6273 , n4888 , n6579 );
    nor g9136 ( n3221 , n8989 , n3 );
    or g9137 ( n6084 , n4462 , n8702 );
    not g9138 ( n3049 , n9732 );
    or g9139 ( n1559 , n10481 , n8563 );
    and g9140 ( n3799 , n3795 , n1736 );
    and g9141 ( n2448 , n11105 , n9355 );
    not g9142 ( n7791 , n3029 );
    or g9143 ( n9969 , n4536 , n10057 );
    or g9144 ( n2677 , n7291 , n5076 );
    xnor g9145 ( n6600 , n11587 , n2684 );
    and g9146 ( n10605 , n12235 , n12204 );
    not g9147 ( n11784 , n4703 );
    or g9148 ( n12935 , n10950 , n8268 );
    and g9149 ( n564 , n3867 , n442 );
    nor g9150 ( n12420 , n11501 , n7630 );
    or g9151 ( n1011 , n536 , n6834 );
    not g9152 ( n8206 , n5962 );
    and g9153 ( n1137 , n1428 , n9191 );
    or g9154 ( n1736 , n5447 , n4861 );
    xnor g9155 ( n1036 , n9958 , n12461 );
    or g9156 ( n11951 , n4716 , n6055 );
    or g9157 ( n1131 , n2449 , n7935 );
    nor g9158 ( n5006 , n11774 , n3828 );
    not g9159 ( n2166 , n4709 );
    buf g9160 ( n10343 , n7342 );
    xnor g9161 ( n7282 , n434 , n3787 );
    not g9162 ( n2131 , n8535 );
    or g9163 ( n12888 , n3265 , n2188 );
    not g9164 ( n2443 , n11553 );
    or g9165 ( n9304 , n1484 , n3432 );
    not g9166 ( n4077 , n3769 );
    or g9167 ( n12222 , n3459 , n3225 );
    xnor g9168 ( n4367 , n12764 , n7319 );
    nor g9169 ( n853 , n1523 , n9002 );
    or g9170 ( n4364 , n6803 , n8763 );
    xor g9171 ( n983 , n1876 , n9303 );
    not g9172 ( n683 , n7061 );
    and g9173 ( n1021 , n8308 , n3409 );
    xnor g9174 ( n5493 , n11184 , n8258 );
    or g9175 ( n12754 , n6769 , n1570 );
    or g9176 ( n4544 , n13080 , n4337 );
    xnor g9177 ( n12731 , n9004 , n11735 );
    xnor g9178 ( n6118 , n970 , n997 );
    not g9179 ( n12380 , n11814 );
    not g9180 ( n12955 , n103 );
    xnor g9181 ( n10635 , n6929 , n12664 );
    xnor g9182 ( n2776 , n163 , n3065 );
    and g9183 ( n4870 , n5238 , n5350 );
    or g9184 ( n4159 , n10270 , n9595 );
    xnor g9185 ( n10070 , n3603 , n1622 );
    xnor g9186 ( n2418 , n9792 , n11428 );
    or g9187 ( n7042 , n5547 , n3981 );
    or g9188 ( n7583 , n1480 , n905 );
    xnor g9189 ( n9065 , n3477 , n7861 );
    xnor g9190 ( n9550 , n10834 , n8264 );
    not g9191 ( n1308 , n13044 );
    xnor g9192 ( n9901 , n4830 , n10541 );
    not g9193 ( n715 , n11396 );
    or g9194 ( n10822 , n3288 , n5291 );
    and g9195 ( n962 , n8840 , n13157 );
    nor g9196 ( n10299 , n6574 , n7614 );
    or g9197 ( n4088 , n6960 , n4723 );
    xnor g9198 ( n743 , n11585 , n12094 );
    and g9199 ( n8305 , n9060 , n8722 );
    not g9200 ( n10041 , n2535 );
    xnor g9201 ( n9000 , n12411 , n4745 );
    xnor g9202 ( n11179 , n2896 , n1061 );
    or g9203 ( n1234 , n5973 , n9075 );
    or g9204 ( n7955 , n12481 , n8750 );
    or g9205 ( n5054 , n3296 , n3114 );
    nor g9206 ( n9562 , n1827 , n13059 );
    and g9207 ( n716 , n9144 , n6870 );
    not g9208 ( n1638 , n5729 );
    not g9209 ( n2463 , n12289 );
    and g9210 ( n10537 , n2045 , n1032 );
    xnor g9211 ( n9983 , n4152 , n2159 );
    or g9212 ( n10959 , n511 , n12162 );
    nor g9213 ( n6613 , n2495 , n2026 );
    not g9214 ( n1526 , n2813 );
    xnor g9215 ( n12 , n6593 , n2511 );
    xor g9216 ( n4719 , n3040 , n7761 );
    xnor g9217 ( n12276 , n7898 , n11285 );
    not g9218 ( n12174 , n6392 );
    xnor g9219 ( n1974 , n12736 , n1994 );
    xnor g9220 ( n9583 , n1304 , n4718 );
    and g9221 ( n1506 , n12348 , n469 );
    not g9222 ( n2484 , n10594 );
    and g9223 ( n5515 , n5138 , n8784 );
    or g9224 ( n3469 , n8324 , n8702 );
    xnor g9225 ( n10523 , n9914 , n697 );
    or g9226 ( n8148 , n3070 , n4930 );
    or g9227 ( n8943 , n6156 , n10207 );
    and g9228 ( n9699 , n1011 , n3350 );
    nor g9229 ( n4675 , n2010 , n10661 );
    or g9230 ( n12452 , n7608 , n12388 );
    not g9231 ( n1017 , n5881 );
    xnor g9232 ( n7527 , n3846 , n6277 );
    xor g9233 ( n10392 , n6209 , n11084 );
    not g9234 ( n5286 , n7573 );
    not g9235 ( n5 , n11511 );
    nor g9236 ( n9335 , n3988 , n2445 );
    and g9237 ( n6615 , n12390 , n1075 );
    or g9238 ( n6502 , n10150 , n9512 );
    xnor g9239 ( n10167 , n10746 , n4712 );
    or g9240 ( n6634 , n2230 , n12120 );
    xnor g9241 ( n7574 , n4391 , n6102 );
    and g9242 ( n11351 , n3420 , n6123 );
    or g9243 ( n2495 , n6755 , n8374 );
    xnor g9244 ( n5621 , n5391 , n9231 );
    and g9245 ( n4819 , n7947 , n12601 );
    or g9246 ( n2862 , n9484 , n2842 );
    xnor g9247 ( n11598 , n7227 , n5231 );
    not g9248 ( n3201 , n7713 );
    xnor g9249 ( n3740 , n11688 , n5374 );
    not g9250 ( n2157 , n11692 );
    nor g9251 ( n3855 , n8331 , n798 );
    or g9252 ( n1311 , n2933 , n13225 );
    or g9253 ( n3770 , n2041 , n1144 );
    or g9254 ( n1740 , n787 , n4947 );
    nor g9255 ( n10705 , n1321 , n3144 );
    nor g9256 ( n3383 , n6107 , n9988 );
    nor g9257 ( n12008 , n4754 , n3533 );
    or g9258 ( n8743 , n11291 , n1026 );
    or g9259 ( n12365 , n4227 , n3418 );
    xor g9260 ( n1790 , n8469 , n9473 );
    or g9261 ( n1274 , n4308 , n3820 );
    or g9262 ( n5904 , n9659 , n395 );
    and g9263 ( n702 , n8234 , n10820 );
    xnor g9264 ( n2743 , n6153 , n2392 );
    or g9265 ( n9830 , n5079 , n8030 );
    and g9266 ( n9149 , n1158 , n1713 );
    not g9267 ( n633 , n5309 );
    or g9268 ( n11022 , n361 , n3039 );
    and g9269 ( n265 , n3847 , n10065 );
    xnor g9270 ( n11048 , n12458 , n1151 );
    or g9271 ( n4771 , n1919 , n8348 );
    xnor g9272 ( n2843 , n11720 , n4045 );
    not g9273 ( n10565 , n8092 );
    not g9274 ( n7485 , n8518 );
    not g9275 ( n2757 , n9732 );
    not g9276 ( n4655 , n3188 );
    xor g9277 ( n10485 , n7040 , n3763 );
    nor g9278 ( n106 , n9592 , n2668 );
    nor g9279 ( n3347 , n9209 , n6528 );
    nor g9280 ( n6792 , n3749 , n46 );
    or g9281 ( n538 , n1141 , n8937 );
    xnor g9282 ( n773 , n172 , n4973 );
    or g9283 ( n5818 , n4456 , n5353 );
    xnor g9284 ( n8651 , n3558 , n11766 );
    nor g9285 ( n12719 , n9138 , n11254 );
    nor g9286 ( n3546 , n8867 , n9827 );
    xnor g9287 ( n520 , n3236 , n9197 );
    and g9288 ( n10935 , n1102 , n11908 );
    xnor g9289 ( n531 , n12135 , n6714 );
    xnor g9290 ( n2852 , n11881 , n6991 );
    and g9291 ( n5505 , n146 , n95 );
    xnor g9292 ( n1776 , n12056 , n446 );
    and g9293 ( n9735 , n9152 , n6457 );
    xnor g9294 ( n7160 , n12949 , n8818 );
    nor g9295 ( n9561 , n9220 , n8333 );
    xnor g9296 ( n1149 , n9496 , n8034 );
    and g9297 ( n3580 , n2838 , n2388 );
    and g9298 ( n1482 , n646 , n47 );
    xnor g9299 ( n6965 , n11279 , n11454 );
    xnor g9300 ( n601 , n8241 , n7462 );
    and g9301 ( n5535 , n3311 , n10606 );
    not g9302 ( n10381 , n8284 );
    not g9303 ( n8248 , n9825 );
    xnor g9304 ( n4039 , n5655 , n2206 );
    nor g9305 ( n10629 , n4199 , n6938 );
    xnor g9306 ( n12275 , n2173 , n3490 );
    or g9307 ( n5465 , n5433 , n4230 );
    or g9308 ( n10212 , n12832 , n1690 );
    or g9309 ( n9970 , n9723 , n10871 );
    nor g9310 ( n3608 , n4026 , n1243 );
    not g9311 ( n1168 , n10162 );
    xnor g9312 ( n8144 , n7578 , n6775 );
    xnor g9313 ( n12845 , n264 , n6500 );
    or g9314 ( n10682 , n856 , n8602 );
    or g9315 ( n11487 , n5226 , n8024 );
    xnor g9316 ( n11077 , n5073 , n12962 );
    and g9317 ( n9098 , n2932 , n11182 );
    or g9318 ( n3708 , n2346 , n8348 );
    or g9319 ( n6490 , n9066 , n7681 );
    or g9320 ( n10566 , n9444 , n4373 );
    xnor g9321 ( n13047 , n11338 , n6609 );
    and g9322 ( n3650 , n9864 , n4224 );
    buf g9323 ( n8702 , n4013 );
    xnor g9324 ( n12291 , n6583 , n1142 );
    and g9325 ( n9855 , n7673 , n1223 );
    or g9326 ( n5335 , n11404 , n12273 );
    not g9327 ( n9325 , n8827 );
    not g9328 ( n6223 , n4006 );
    and g9329 ( n5750 , n11969 , n4560 );
    or g9330 ( n6076 , n10220 , n12215 );
    and g9331 ( n1004 , n570 , n3366 );
    not g9332 ( n8295 , n11017 );
    and g9333 ( n2005 , n7828 , n3888 );
    xnor g9334 ( n12067 , n7734 , n1374 );
    xnor g9335 ( n2040 , n11722 , n7502 );
    not g9336 ( n12615 , n12961 );
    and g9337 ( n487 , n2590 , n7720 );
    xnor g9338 ( n1120 , n10160 , n10625 );
    xnor g9339 ( n4734 , n4094 , n5323 );
    or g9340 ( n4869 , n3095 , n2983 );
    or g9341 ( n9653 , n3480 , n3119 );
    xnor g9342 ( n8023 , n8801 , n12509 );
    xnor g9343 ( n5110 , n11456 , n7589 );
    xnor g9344 ( n7070 , n2065 , n1565 );
    xnor g9345 ( n9458 , n8547 , n416 );
    or g9346 ( n10500 , n5782 , n10319 );
    and g9347 ( n3883 , n12270 , n12076 );
    xnor g9348 ( n1726 , n6372 , n10624 );
    xnor g9349 ( n806 , n271 , n12647 );
    or g9350 ( n1170 , n5105 , n8505 );
    or g9351 ( n1691 , n385 , n13056 );
    xnor g9352 ( n6964 , n2564 , n10147 );
    or g9353 ( n4393 , n7748 , n2133 );
    and g9354 ( n12589 , n12705 , n9051 );
    xnor g9355 ( n9825 , n2677 , n6708 );
    xnor g9356 ( n687 , n2886 , n8854 );
    or g9357 ( n3275 , n9559 , n4690 );
    nor g9358 ( n9045 , n5439 , n10315 );
    xnor g9359 ( n6477 , n1509 , n2563 );
    or g9360 ( n1606 , n10498 , n10889 );
    xnor g9361 ( n5534 , n8825 , n8576 );
    xnor g9362 ( n5857 , n9625 , n12950 );
    not g9363 ( n602 , n2824 );
    xnor g9364 ( n2093 , n6697 , n1842 );
    or g9365 ( n5603 , n8941 , n5797 );
    and g9366 ( n13078 , n840 , n6667 );
    and g9367 ( n427 , n3006 , n4470 );
    not g9368 ( n12813 , n11897 );
    and g9369 ( n4789 , n8940 , n11222 );
    or g9370 ( n8028 , n9761 , n1570 );
    not g9371 ( n4305 , n10111 );
    or g9372 ( n8346 , n9502 , n2719 );
    and g9373 ( n3760 , n10908 , n10408 );
    xnor g9374 ( n11102 , n6426 , n5032 );
    xnor g9375 ( n6616 , n109 , n3287 );
    not g9376 ( n3232 , n62 );
    or g9377 ( n126 , n2488 , n793 );
    or g9378 ( n7227 , n2825 , n6404 );
    nor g9379 ( n4068 , n9630 , n12359 );
    or g9380 ( n12253 , n3333 , n6715 );
    xor g9381 ( n4102 , n1978 , n3168 );
    not g9382 ( n10977 , n2174 );
    and g9383 ( n11673 , n11236 , n854 );
    nor g9384 ( n9923 , n12389 , n7539 );
    xnor g9385 ( n3930 , n11913 , n8409 );
    xnor g9386 ( n3896 , n10969 , n2843 );
    or g9387 ( n9628 , n2625 , n4386 );
    nor g9388 ( n9754 , n7833 , n791 );
    and g9389 ( n2209 , n12141 , n10513 );
    not g9390 ( n3630 , n22 );
    not g9391 ( n3655 , n3123 );
    or g9392 ( n5705 , n8817 , n10106 );
    or g9393 ( n10391 , n898 , n4154 );
    and g9394 ( n4959 , n2860 , n10125 );
    or g9395 ( n1062 , n6038 , n1468 );
    xnor g9396 ( n1707 , n9248 , n6872 );
    xnor g9397 ( n1384 , n7201 , n11337 );
    not g9398 ( n2226 , n12605 );
    not g9399 ( n7283 , n1307 );
    or g9400 ( n8370 , n2444 , n11461 );
    or g9401 ( n2114 , n11094 , n7530 );
    and g9402 ( n6442 , n1452 , n5503 );
    nor g9403 ( n13030 , n4097 , n12876 );
    xnor g9404 ( n12279 , n6573 , n9671 );
    or g9405 ( n9420 , n3974 , n9018 );
    or g9406 ( n5353 , n8498 , n4373 );
    not g9407 ( n8609 , n11061 );
    and g9408 ( n9737 , n6024 , n4915 );
    not g9409 ( n9340 , n13161 );
    nor g9410 ( n8439 , n11444 , n12430 );
    or g9411 ( n5850 , n9679 , n9118 );
    xnor g9412 ( n5894 , n11332 , n4240 );
    xnor g9413 ( n11586 , n10316 , n12022 );
    not g9414 ( n12772 , n4293 );
    xnor g9415 ( n11126 , n7796 , n4829 );
    xnor g9416 ( n3391 , n6778 , n12110 );
    xnor g9417 ( n187 , n11005 , n1896 );
    not g9418 ( n8849 , n12482 );
    xnor g9419 ( n6969 , n155 , n9806 );
    xnor g9420 ( n9440 , n8536 , n3896 );
    or g9421 ( n9346 , n3425 , n1028 );
    and g9422 ( n11645 , n2888 , n3764 );
    and g9423 ( n10697 , n5483 , n6889 );
    or g9424 ( n1553 , n583 , n11405 );
    and g9425 ( n2927 , n12022 , n10316 );
    nor g9426 ( n2594 , n691 , n1874 );
    and g9427 ( n8196 , n1751 , n9801 );
    nor g9428 ( n1924 , n10054 , n10651 );
    xnor g9429 ( n1386 , n9944 , n1898 );
    and g9430 ( n8696 , n8124 , n4262 );
    xnor g9431 ( n10743 , n6943 , n7030 );
    xnor g9432 ( n9823 , n12021 , n11695 );
    or g9433 ( n4915 , n7597 , n6732 );
    or g9434 ( n596 , n10286 , n6944 );
    or g9435 ( n6305 , n10898 , n12847 );
    or g9436 ( n11095 , n9400 , n8030 );
    not g9437 ( n18 , n4357 );
    and g9438 ( n3566 , n13096 , n6146 );
    or g9439 ( n11566 , n8431 , n12666 );
    and g9440 ( n2116 , n7891 , n8048 );
    xnor g9441 ( n9574 , n6513 , n725 );
    nor g9442 ( n9734 , n3964 , n6879 );
    or g9443 ( n3453 , n0 , n4230 );
    and g9444 ( n1430 , n6444 , n11489 );
    or g9445 ( n12178 , n11171 , n12847 );
    not g9446 ( n8280 , n4368 );
    or g9447 ( n10241 , n12312 , n12781 );
    xnor g9448 ( n3925 , n4953 , n8119 );
    xnor g9449 ( n556 , n8313 , n1715 );
    not g9450 ( n13051 , n9669 );
    or g9451 ( n10232 , n7677 , n12048 );
    and g9452 ( n1044 , n11951 , n11936 );
    and g9453 ( n2985 , n4690 , n9559 );
    xnor g9454 ( n7397 , n11875 , n11755 );
    not g9455 ( n6575 , n4695 );
    and g9456 ( n5371 , n1183 , n7747 );
    xnor g9457 ( n6134 , n8867 , n2382 );
    and g9458 ( n10813 , n8208 , n12375 );
    xnor g9459 ( n4548 , n2208 , n3402 );
    not g9460 ( n9512 , n2334 );
    or g9461 ( n3393 , n4655 , n6924 );
    xnor g9462 ( n8049 , n10878 , n8308 );
    and g9463 ( n361 , n1510 , n12816 );
    or g9464 ( n2008 , n8090 , n11282 );
    not g9465 ( n8225 , n5729 );
    or g9466 ( n8924 , n4967 , n3981 );
    and g9467 ( n3567 , n1499 , n1210 );
    not g9468 ( n11427 , n12937 );
    and g9469 ( n4348 , n12003 , n11109 );
    xnor g9470 ( n9201 , n6131 , n9757 );
    and g9471 ( n4684 , n4977 , n6864 );
    and g9472 ( n3644 , n12920 , n9727 );
    or g9473 ( n7695 , n12477 , n8231 );
    not g9474 ( n3586 , n3263 );
    not g9475 ( n9429 , n9528 );
    or g9476 ( n36 , n3049 , n5264 );
    not g9477 ( n473 , n4459 );
    or g9478 ( n7125 , n11588 , n8748 );
    nor g9479 ( n12247 , n7671 , n8078 );
    or g9480 ( n430 , n10138 , n9386 );
    xnor g9481 ( n3289 , n8944 , n6567 );
    and g9482 ( n2803 , n7650 , n3657 );
    or g9483 ( n6329 , n345 , n1961 );
    xnor g9484 ( n1590 , n10294 , n13222 );
    xnor g9485 ( n4051 , n10992 , n8015 );
    or g9486 ( n7600 , n3564 , n10029 );
    xnor g9487 ( n8554 , n3204 , n4729 );
    nor g9488 ( n4699 , n7161 , n8030 );
    or g9489 ( n11704 , n2262 , n4865 );
    not g9490 ( n290 , n5457 );
    not g9491 ( n6366 , n3625 );
    xnor g9492 ( n10699 , n4086 , n1920 );
    and g9493 ( n2026 , n889 , n7897 );
    not g9494 ( n1329 , n11429 );
    not g9495 ( n1451 , n9906 );
    not g9496 ( n3318 , n6604 );
    xnor g9497 ( n763 , n1170 , n5872 );
    xnor g9498 ( n2196 , n5128 , n6200 );
    or g9499 ( n2783 , n987 , n10319 );
    xnor g9500 ( n2039 , n4467 , n12142 );
    not g9501 ( n482 , n2777 );
    xnor g9502 ( n6865 , n346 , n5755 );
    or g9503 ( n2528 , n3726 , n2133 );
    xnor g9504 ( n3494 , n8476 , n10689 );
    xnor g9505 ( n788 , n9892 , n10526 );
    xnor g9506 ( n3756 , n13 , n11687 );
    and g9507 ( n4579 , n5832 , n3303 );
    xnor g9508 ( n12436 , n4508 , n11432 );
    or g9509 ( n11947 , n4715 , n6561 );
    not g9510 ( n11926 , n9127 );
    not g9511 ( n7033 , n9093 );
    xnor g9512 ( n6985 , n11393 , n2997 );
    nor g9513 ( n1551 , n12247 , n10754 );
    xnor g9514 ( n12571 , n4525 , n7684 );
    and g9515 ( n979 , n4931 , n11084 );
    not g9516 ( n7846 , n2590 );
    xnor g9517 ( n3190 , n8747 , n10737 );
    not g9518 ( n11807 , n8359 );
    xnor g9519 ( n328 , n6525 , n8232 );
    and g9520 ( n12401 , n6995 , n8690 );
    not g9521 ( n2306 , n2979 );
    and g9522 ( n6062 , n11263 , n13081 );
    and g9523 ( n13192 , n6830 , n3786 );
    and g9524 ( n1297 , n8197 , n10245 );
    or g9525 ( n10413 , n13146 , n8564 );
    xnor g9526 ( n1811 , n6700 , n5277 );
    xnor g9527 ( n7162 , n9553 , n6059 );
    not g9528 ( n5679 , n6655 );
    xnor g9529 ( n11205 , n3699 , n4976 );
    and g9530 ( n4831 , n8111 , n2967 );
    xnor g9531 ( n370 , n12453 , n7766 );
    or g9532 ( n5228 , n1737 , n9638 );
    and g9533 ( n3155 , n925 , n8199 );
    not g9534 ( n3103 , n11332 );
    not g9535 ( n10681 , n3130 );
    not g9536 ( n12438 , n6251 );
    or g9537 ( n1766 , n12568 , n8534 );
    or g9538 ( n7811 , n829 , n9075 );
    or g9539 ( n4988 , n6986 , n10430 );
    or g9540 ( n123 , n991 , n12501 );
    and g9541 ( n4350 , n9662 , n10386 );
    or g9542 ( n4359 , n1536 , n2675 );
    and g9543 ( n5205 , n2044 , n12293 );
    xnor g9544 ( n12639 , n3542 , n5418 );
    and g9545 ( n9292 , n7434 , n8185 );
    and g9546 ( n7040 , n2163 , n2618 );
    xnor g9547 ( n9775 , n5689 , n2467 );
    not g9548 ( n12655 , n10408 );
    or g9549 ( n13174 , n2698 , n9203 );
    not g9550 ( n1621 , n10162 );
    not g9551 ( n11087 , n5470 );
    not g9552 ( n9790 , n9965 );
    and g9553 ( n2436 , n2407 , n2578 );
    or g9554 ( n8277 , n1571 , n7935 );
    and g9555 ( n3396 , n10884 , n5926 );
    xnor g9556 ( n9841 , n12074 , n11767 );
    and g9557 ( n7409 , n11490 , n1206 );
    or g9558 ( n6259 , n13182 , n1985 );
    or g9559 ( n2327 , n794 , n2980 );
    and g9560 ( n7182 , n3336 , n5685 );
    xnor g9561 ( n11177 , n752 , n3982 );
    not g9562 ( n13097 , n9049 );
    xnor g9563 ( n3887 , n3836 , n11892 );
    and g9564 ( n2676 , n7722 , n11485 );
    or g9565 ( n5843 , n1987 , n285 );
    xnor g9566 ( n13092 , n6712 , n12186 );
    and g9567 ( n10958 , n7010 , n2752 );
    xnor g9568 ( n8758 , n9609 , n3134 );
    xnor g9569 ( n2626 , n12942 , n717 );
    xnor g9570 ( n12182 , n10109 , n3232 );
    or g9571 ( n7231 , n560 , n8490 );
    or g9572 ( n3927 , n7231 , n6583 );
    nor g9573 ( n1352 , n12816 , n1510 );
    and g9574 ( n9684 , n3102 , n10385 );
    not g9575 ( n2083 , n791 );
    and g9576 ( n1342 , n6137 , n6379 );
    xnor g9577 ( n1944 , n3357 , n3012 );
    not g9578 ( n9281 , n11508 );
    xnor g9579 ( n886 , n8122 , n8995 );
    or g9580 ( n7303 , n5076 , n10106 );
    xnor g9581 ( n5532 , n1391 , n3737 );
    or g9582 ( n11958 , n12493 , n177 );
    or g9583 ( n6644 , n10761 , n206 );
    nor g9584 ( n6298 , n7161 , n5076 );
    and g9585 ( n3392 , n9353 , n10063 );
    xnor g9586 ( n1700 , n9074 , n4799 );
    xnor g9587 ( n414 , n9939 , n2356 );
    or g9588 ( n3366 , n8174 , n2958 );
    not g9589 ( n12732 , n12965 );
    nor g9590 ( n9870 , n6053 , n3080 );
    xnor g9591 ( n4765 , n6661 , n6675 );
    xnor g9592 ( n4581 , n14 , n3313 );
    or g9593 ( n7284 , n3505 , n6689 );
    not g9594 ( n6180 , n1283 );
    not g9595 ( n2453 , n11890 );
    xnor g9596 ( n380 , n8240 , n5373 );
    and g9597 ( n6433 , n1912 , n2498 );
    or g9598 ( n11060 , n12660 , n4881 );
    and g9599 ( n11873 , n5768 , n10563 );
    xnor g9600 ( n5682 , n8823 , n4434 );
    or g9601 ( n2782 , n1250 , n3113 );
    or g9602 ( n7011 , n12395 , n4960 );
    xnor g9603 ( n6701 , n8207 , n1106 );
    and g9604 ( n8963 , n8847 , n3007 );
    xnor g9605 ( n5979 , n12279 , n9210 );
    and g9606 ( n10140 , n848 , n10620 );
    and g9607 ( n7379 , n10196 , n10104 );
    not g9608 ( n8700 , n4813 );
    or g9609 ( n9764 , n5770 , n4312 );
    xnor g9610 ( n11541 , n4639 , n1457 );
    and g9611 ( n4919 , n7468 , n8442 );
    xnor g9612 ( n12347 , n7910 , n11358 );
    xnor g9613 ( n7115 , n5126 , n1363 );
    and g9614 ( n5870 , n4964 , n510 );
    not g9615 ( n13088 , n6537 );
    and g9616 ( n4413 , n5661 , n7174 );
    and g9617 ( n6786 , n5092 , n12462 );
    or g9618 ( n7738 , n2829 , n228 );
    xnor g9619 ( n10627 , n4661 , n8713 );
    xor g9620 ( n4874 , n11288 , n8408 );
    and g9621 ( n5084 , n2643 , n4629 );
    xor g9622 ( n7455 , n4828 , n8197 );
    not g9623 ( n11683 , n6937 );
    or g9624 ( n6070 , n10792 , n542 );
    and g9625 ( n8530 , n4863 , n243 );
    or g9626 ( n667 , n11239 , n8030 );
    or g9627 ( n7003 , n8240 , n9123 );
    xnor g9628 ( n141 , n7289 , n5463 );
    xnor g9629 ( n10484 , n1756 , n6380 );
    xnor g9630 ( n8456 , n9871 , n9350 );
    xnor g9631 ( n2036 , n5810 , n10720 );
    or g9632 ( n9407 , n2582 , n6635 );
    or g9633 ( n4053 , n4201 , n11144 );
    not g9634 ( n5433 , n9887 );
    not g9635 ( n8129 , n5962 );
    or g9636 ( n11238 , n1053 , n9491 );
    xnor g9637 ( n11004 , n9433 , n5628 );
    or g9638 ( n7222 , n6651 , n2658 );
    or g9639 ( n9659 , n8585 , n4640 );
    not g9640 ( n4116 , n3130 );
    or g9641 ( n13096 , n3069 , n8365 );
    xnor g9642 ( n7909 , n9602 , n2870 );
    and g9643 ( n3723 , n8900 , n5284 );
    xnor g9644 ( n85 , n8256 , n5582 );
    not g9645 ( n6405 , n124 );
    not g9646 ( n9245 , n9214 );
    not g9647 ( n2515 , n8924 );
    and g9648 ( n10725 , n12007 , n2066 );
    or g9649 ( n677 , n1558 , n1692 );
    not g9650 ( n13028 , n9732 );
    nor g9651 ( n12687 , n4458 , n9091 );
    or g9652 ( n4701 , n2214 , n10589 );
    or g9653 ( n395 , n11466 , n479 );
    nor g9654 ( n5258 , n6009 , n11089 );
    not g9655 ( n5372 , n6998 );
    not g9656 ( n10430 , n3130 );
    not g9657 ( n3970 , n11306 );
    xnor g9658 ( n2994 , n13144 , n4911 );
    xnor g9659 ( n12619 , n2767 , n6617 );
    xnor g9660 ( n8135 , n10623 , n1902 );
    xnor g9661 ( n1547 , n986 , n9471 );
    xnor g9662 ( n1882 , n8064 , n3843 );
    xnor g9663 ( n1573 , n7476 , n11948 );
    or g9664 ( n13241 , n11915 , n4133 );
    not g9665 ( n7586 , n8398 );
    and g9666 ( n6011 , n590 , n11168 );
    nor g9667 ( n6539 , n7100 , n9045 );
    nor g9668 ( n6145 , n10785 , n429 );
    xnor g9669 ( n12361 , n9901 , n1350 );
    xnor g9670 ( n6107 , n9344 , n5735 );
    not g9671 ( n11006 , n1065 );
    and g9672 ( n10809 , n864 , n8458 );
    xnor g9673 ( n1350 , n11801 , n6216 );
    not g9674 ( n11680 , n11891 );
    or g9675 ( n2763 , n1280 , n12907 );
    and g9676 ( n8718 , n1346 , n5839 );
    xnor g9677 ( n13015 , n1537 , n5464 );
    nor g9678 ( n8623 , n2323 , n183 );
    and g9679 ( n8046 , n937 , n287 );
    and g9680 ( n212 , n5257 , n8425 );
    xnor g9681 ( n11158 , n11108 , n887 );
    not g9682 ( n153 , n1721 );
    or g9683 ( n8022 , n5231 , n7227 );
    or g9684 ( n1445 , n3780 , n8685 );
    and g9685 ( n2186 , n3639 , n503 );
    xnor g9686 ( n9213 , n10540 , n8343 );
    not g9687 ( n3459 , n3669 );
    not g9688 ( n3906 , n11881 );
    or g9689 ( n6466 , n7604 , n4585 );
    xnor g9690 ( n6927 , n659 , n1591 );
    xnor g9691 ( n1802 , n5465 , n7760 );
    or g9692 ( n2755 , n7986 , n8540 );
    or g9693 ( n6859 , n8776 , n10761 );
    or g9694 ( n1979 , n10221 , n2977 );
    xor g9695 ( n8158 , n12953 , n6140 );
    not g9696 ( n2462 , n13058 );
    or g9697 ( n7194 , n6971 , n3798 );
    xnor g9698 ( n11274 , n3224 , n340 );
    and g9699 ( n8606 , n9353 , n9915 );
    not g9700 ( n13146 , n3868 );
    xnor g9701 ( n5014 , n9858 , n618 );
    not g9702 ( n6295 , n2758 );
    xnor g9703 ( n5124 , n10167 , n4643 );
    nor g9704 ( n5213 , n11572 , n1584 );
    xnor g9705 ( n10970 , n7887 , n626 );
    xnor g9706 ( n3964 , n9938 , n8184 );
    and g9707 ( n8577 , n9797 , n12584 );
    nor g9708 ( n9527 , n2541 , n11280 );
    or g9709 ( n12417 , n48 , n11144 );
    or g9710 ( n4206 , n3755 , n2845 );
    or g9711 ( n7933 , n13168 , n1985 );
    or g9712 ( n2466 , n2861 , n12388 );
    and g9713 ( n4414 , n12734 , n2441 );
    buf g9714 ( n10761 , n6405 );
    or g9715 ( n6379 , n5700 , n9975 );
    or g9716 ( n3527 , n12596 , n5242 );
    not g9717 ( n7900 , n9747 );
    and g9718 ( n1778 , n12745 , n1968 );
    or g9719 ( n11511 , n10343 , n6983 );
    xnor g9720 ( n11676 , n6296 , n11073 );
    not g9721 ( n7089 , n6286 );
    not g9722 ( n8621 , n9415 );
    xnor g9723 ( n7123 , n11004 , n5994 );
    xnor g9724 ( n12423 , n90 , n6262 );
    xnor g9725 ( n8377 , n5447 , n2367 );
    or g9726 ( n7226 , n6011 , n13105 );
    not g9727 ( n5035 , n13040 );
    xnor g9728 ( n474 , n11930 , n9316 );
    or g9729 ( n12766 , n595 , n3221 );
    xnor g9730 ( n7660 , n1490 , n54 );
    and g9731 ( n1854 , n3017 , n6921 );
    not g9732 ( n12969 , n7229 );
    or g9733 ( n7731 , n6638 , n1043 );
    or g9734 ( n2156 , n10000 , n10534 );
    not g9735 ( n1505 , n7779 );
    xor g9736 ( n7238 , n4957 , n8452 );
    nor g9737 ( n10441 , n17 , n11460 );
    xnor g9738 ( n12486 , n10502 , n7617 );
    xnor g9739 ( n8140 , n11765 , n8851 );
    not g9740 ( n12959 , n10770 );
    or g9741 ( n249 , n1680 , n451 );
    xnor g9742 ( n1415 , n3434 , n5211 );
    buf g9743 ( n4936 , n2623 );
    and g9744 ( n10923 , n1378 , n9835 );
    or g9745 ( n7689 , n12757 , n225 );
    not g9746 ( n6557 , n8332 );
    and g9747 ( n4908 , n6668 , n10451 );
    or g9748 ( n12433 , n7575 , n6624 );
    xnor g9749 ( n796 , n12506 , n4631 );
    and g9750 ( n10821 , n7857 , n1396 );
    nor g9751 ( n4763 , n9555 , n1830 );
    nor g9752 ( n1224 , n2166 , n3862 );
    not g9753 ( n899 , n9187 );
    not g9754 ( n467 , n10572 );
    or g9755 ( n7269 , n822 , n11176 );
    xor g9756 ( n1278 , n5334 , n9215 );
    not g9757 ( n4980 , n11634 );
    and g9758 ( n2615 , n11051 , n7953 );
    and g9759 ( n13132 , n1682 , n1306 );
    and g9760 ( n10360 , n3302 , n8133 );
    or g9761 ( n2920 , n12814 , n5740 );
    nor g9762 ( n8930 , n484 , n7618 );
    xnor g9763 ( n9599 , n9853 , n12044 );
    nor g9764 ( n2933 , n3589 , n7217 );
    not g9765 ( n4253 , n10770 );
    nor g9766 ( n335 , n688 , n9816 );
    xnor g9767 ( n769 , n10919 , n4765 );
    or g9768 ( n9409 , n5441 , n4164 );
    or g9769 ( n11041 , n7769 , n7162 );
    nor g9770 ( n4032 , n6530 , n4950 );
    nor g9771 ( n12476 , n10499 , n12269 );
    not g9772 ( n1963 , n9204 );
    or g9773 ( n9334 , n11381 , n1848 );
    nor g9774 ( n11081 , n4800 , n2089 );
    not g9775 ( n578 , n7959 );
    and g9776 ( n4111 , n7772 , n12853 );
    and g9777 ( n10249 , n944 , n1673 );
    not g9778 ( n3588 , n6831 );
    xnor g9779 ( n1272 , n4325 , n1743 );
    and g9780 ( n2754 , n2411 , n757 );
    not g9781 ( n10112 , n10594 );
    and g9782 ( n3104 , n11108 , n5731 );
    nor g9783 ( n9227 , n9166 , n4284 );
    xor g9784 ( n6143 , n1609 , n8544 );
    nor g9785 ( n9009 , n8215 , n270 );
    xnor g9786 ( n9665 , n7843 , n5151 );
    or g9787 ( n12647 , n12316 , n11960 );
    not g9788 ( n7342 , n9249 );
    not g9789 ( n2104 , n1202 );
    nor g9790 ( n10901 , n6559 , n8071 );
    not g9791 ( n8142 , n1731 );
    xnor g9792 ( n12564 , n6338 , n9644 );
    and g9793 ( n11141 , n759 , n12035 );
    not g9794 ( n1367 , n3558 );
    or g9795 ( n2100 , n9931 , n8348 );
    xnor g9796 ( n3672 , n7769 , n2959 );
    or g9797 ( n8938 , n7201 , n10725 );
    or g9798 ( n6323 , n9378 , n2632 );
    xnor g9799 ( n8427 , n7514 , n10305 );
    xnor g9800 ( n10317 , n1148 , n13003 );
    xnor g9801 ( n8227 , n7973 , n5014 );
    or g9802 ( n7862 , n10256 , n9159 );
    or g9803 ( n11123 , n1869 , n3981 );
    not g9804 ( n11950 , n13058 );
    xnor g9805 ( n12690 , n12449 , n7104 );
    xnor g9806 ( n11631 , n3109 , n5275 );
    or g9807 ( n6300 , n2767 , n10584 );
    nor g9808 ( n2171 , n8847 , n3007 );
    buf g9809 ( n6404 , n5041 );
    xnor g9810 ( n9616 , n1669 , n4820 );
    xnor g9811 ( n8369 , n12771 , n5813 );
    or g9812 ( n4916 , n12411 , n4745 );
    xnor g9813 ( n8937 , n4690 , n11435 );
    not g9814 ( n13117 , n9531 );
    xnor g9815 ( n3994 , n12285 , n82 );
    not g9816 ( n8486 , n12987 );
    or g9817 ( n7340 , n10929 , n12273 );
    xnor g9818 ( n5453 , n1245 , n6386 );
    not g9819 ( n8485 , n4798 );
    and g9820 ( n91 , n6796 , n8984 );
    not g9821 ( n6210 , n13201 );
    and g9822 ( n12267 , n5554 , n11321 );
    not g9823 ( n10105 , n9125 );
    and g9824 ( n9062 , n12626 , n1562 );
    not g9825 ( n12212 , n3448 );
    nor g9826 ( n6 , n5791 , n2517 );
    xnor g9827 ( n1341 , n8654 , n2457 );
    or g9828 ( n13072 , n10977 , n4230 );
    nor g9829 ( n12608 , n4649 , n10866 );
    nor g9830 ( n5345 , n5206 , n9789 );
    xnor g9831 ( n6872 , n3828 , n4566 );
    xnor g9832 ( n358 , n530 , n1022 );
    or g9833 ( n3279 , n2474 , n12017 );
    or g9834 ( n12762 , n785 , n8534 );
    and g9835 ( n8359 , n6341 , n9244 );
    xnor g9836 ( n4477 , n9824 , n13078 );
    or g9837 ( n11343 , n11929 , n2958 );
    and g9838 ( n1830 , n6873 , n7555 );
    xnor g9839 ( n6682 , n3599 , n773 );
    not g9840 ( n3508 , n7702 );
    xnor g9841 ( n5594 , n7296 , n12546 );
    not g9842 ( n958 , n13065 );
    and g9843 ( n698 , n4114 , n510 );
    and g9844 ( n7383 , n1672 , n6321 );
    or g9845 ( n6611 , n12324 , n4724 );
    and g9846 ( n2841 , n11771 , n128 );
    xnor g9847 ( n7246 , n8055 , n712 );
    not g9848 ( n5667 , n9906 );
    and g9849 ( n1623 , n6228 , n12774 );
    or g9850 ( n8170 , n6630 , n8005 );
    nor g9851 ( n5612 , n5140 , n6791 );
    not g9852 ( n10447 , n4006 );
    xnor g9853 ( n5276 , n11301 , n5444 );
    or g9854 ( n4898 , n12465 , n644 );
    xnor g9855 ( n12562 , n5052 , n11325 );
    xor g9856 ( n4156 , n5044 , n1444 );
    xnor g9857 ( n12409 , n3905 , n9111 );
    not g9858 ( n6274 , n10560 );
    and g9859 ( n11684 , n9148 , n282 );
    not g9860 ( n464 , n11448 );
    or g9861 ( n9645 , n18 , n6732 );
    xnor g9862 ( n12898 , n5558 , n9941 );
    and g9863 ( n3133 , n6541 , n9519 );
    and g9864 ( n6643 , n153 , n9996 );
    and g9865 ( n8590 , n2057 , n1198 );
    and g9866 ( n4259 , n5559 , n1526 );
    or g9867 ( n1305 , n9318 , n10532 );
    and g9868 ( n10671 , n8925 , n2930 );
    or g9869 ( n9104 , n11170 , n5575 );
    not g9870 ( n2080 , n7812 );
    not g9871 ( n3208 , n9846 );
    nor g9872 ( n2780 , n8338 , n4200 );
    not g9873 ( n2441 , n3097 );
    and g9874 ( n9812 , n13009 , n7105 );
    nor g9875 ( n6002 , n10133 , n8052 );
    and g9876 ( n639 , n1050 , n11728 );
    or g9877 ( n3560 , n9868 , n7846 );
    and g9878 ( n5647 , n11807 , n1366 );
    or g9879 ( n3938 , n8720 , n1554 );
    not g9880 ( n947 , n11324 );
    and g9881 ( n10563 , n10770 , n3769 );
    or g9882 ( n5639 , n495 , n6853 );
    or g9883 ( n2090 , n947 , n11950 );
    xnor g9884 ( n11622 , n8994 , n6847 );
    nor g9885 ( n1694 , n10167 , n11158 );
    or g9886 ( n5855 , n7852 , n1449 );
    or g9887 ( n5238 , n3032 , n12244 );
    or g9888 ( n1550 , n9867 , n5076 );
    xnor g9889 ( n4476 , n3358 , n5927 );
    nor g9890 ( n1429 , n8180 , n2667 );
    xnor g9891 ( n11658 , n2248 , n462 );
    or g9892 ( n619 , n8919 , n8549 );
    not g9893 ( n10258 , n9875 );
    xnor g9894 ( n9189 , n10945 , n3969 );
    or g9895 ( n3245 , n4491 , n11592 );
    and g9896 ( n8965 , n2773 , n6380 );
    or g9897 ( n9529 , n11864 , n8079 );
    or g9898 ( n12130 , n6968 , n10761 );
    xnor g9899 ( n12836 , n13037 , n12865 );
    nor g9900 ( n6779 , n1839 , n7182 );
    not g9901 ( n8755 , n2393 );
    or g9902 ( n5956 , n8249 , n7723 );
    or g9903 ( n8430 , n1082 , n12258 );
    or g9904 ( n12580 , n12837 , n4230 );
    not g9905 ( n6731 , n10809 );
    or g9906 ( n457 , n2941 , n9822 );
    xnor g9907 ( n2138 , n1068 , n11538 );
    xnor g9908 ( n3548 , n9775 , n4282 );
    and g9909 ( n4250 , n2284 , n8770 );
    not g9910 ( n848 , n1569 );
    xnor g9911 ( n9726 , n2359 , n4871 );
    or g9912 ( n7319 , n3805 , n2675 );
    nor g9913 ( n4109 , n9838 , n12943 );
    xnor g9914 ( n12591 , n10310 , n12414 );
    nor g9915 ( n2733 , n12272 , n10455 );
    xnor g9916 ( n11280 , n8285 , n5481 );
    or g9917 ( n7096 , n3572 , n9080 );
    or g9918 ( n9955 , n5306 , n12544 );
    nor g9919 ( n7631 , n7648 , n11208 );
    not g9920 ( n8941 , n4335 );
    or g9921 ( n11240 , n9035 , n3794 );
    or g9922 ( n1745 , n3104 , n11093 );
    or g9923 ( n8956 , n8277 , n2337 );
    and g9924 ( n9232 , n2136 , n13069 );
    xnor g9925 ( n1201 , n2925 , n4583 );
    xnor g9926 ( n2016 , n10152 , n8810 );
    and g9927 ( n7834 , n4530 , n7256 );
    xnor g9928 ( n957 , n3984 , n12964 );
    and g9929 ( n9367 , n1064 , n12952 );
    or g9930 ( n7897 , n6271 , n8754 );
    xnor g9931 ( n12488 , n1535 , n5775 );
    or g9932 ( n1747 , n542 , n1570 );
    or g9933 ( n8406 , n2705 , n5387 );
    or g9934 ( n13212 , n7396 , n7723 );
    not g9935 ( n1659 , n11327 );
    xnor g9936 ( n5747 , n6537 , n7670 );
    not g9937 ( n2536 , n6917 );
    or g9938 ( n10611 , n10795 , n5992 );
    and g9939 ( n2707 , n3684 , n11672 );
    and g9940 ( n7562 , n5696 , n538 );
    and g9941 ( n11425 , n6512 , n11189 );
    and g9942 ( n919 , n11240 , n2322 );
    and g9943 ( n6547 , n7098 , n9349 );
    not g9944 ( n9538 , n5995 );
    not g9945 ( n6439 , n8233 );
    and g9946 ( n10030 , n12455 , n12161 );
    and g9947 ( n10582 , n5343 , n2821 );
    xnor g9948 ( n1960 , n7340 , n9287 );
    or g9949 ( n3617 , n3255 , n6823 );
    and g9950 ( n9011 , n368 , n10839 );
    and g9951 ( n5504 , n7772 , n9093 );
    or g9952 ( n5231 , n3225 , n1570 );
    not g9953 ( n7152 , n3815 );
    not g9954 ( n2669 , n2174 );
    xnor g9955 ( n10688 , n3191 , n8588 );
    or g9956 ( n3343 , n4961 , n7292 );
    and g9957 ( n10253 , n126 , n5783 );
    not g9958 ( n6606 , n10785 );
    or g9959 ( n8457 , n6846 , n8534 );
    or g9960 ( n7108 , n12711 , n11259 );
    and g9961 ( n8452 , n8228 , n5962 );
    or g9962 ( n3647 , n10761 , n7935 );
    not g9963 ( n8754 , n2590 );
    xnor g9964 ( n606 , n5441 , n4164 );
    xnor g9965 ( n915 , n1028 , n3425 );
    or g9966 ( n12326 , n12558 , n11397 );
    and g9967 ( n2513 , n12304 , n12574 );
    xnor g9968 ( n4526 , n10317 , n3023 );
    and g9969 ( n3176 , n2402 , n12451 );
    or g9970 ( n11597 , n1634 , n12997 );
    and g9971 ( n1458 , n5452 , n12681 );
    xnor g9972 ( n2906 , n13110 , n5005 );
    xnor g9973 ( n6075 , n11500 , n4769 );
    xnor g9974 ( n7237 , n3776 , n1551 );
    not g9975 ( n146 , n4579 );
    not g9976 ( n8631 , n12091 );
    or g9977 ( n10491 , n5839 , n1346 );
    or g9978 ( n352 , n7621 , n2077 );
    not g9979 ( n11400 , n12260 );
    xnor g9980 ( n8774 , n6436 , n6735 );
    buf g9981 ( n4947 , n9709 );
    nor g9982 ( n11770 , n9621 , n7888 );
    or g9983 ( n7300 , n11210 , n2116 );
    and g9984 ( n1426 , n12371 , n12297 );
    xnor g9985 ( n10084 , n10358 , n3574 );
    not g9986 ( n4481 , n3579 );
    xnor g9987 ( n3252 , n8369 , n3286 );
    xnor g9988 ( n9979 , n6233 , n5598 );
    xnor g9989 ( n1266 , n1797 , n4676 );
    and g9990 ( n627 , n5134 , n6311 );
    nor g9991 ( n2245 , n9763 , n11812 );
    and g9992 ( n5615 , n6639 , n12031 );
    and g9993 ( n10601 , n9484 , n2842 );
    xnor g9994 ( n8241 , n9597 , n7531 );
    or g9995 ( n8881 , n2095 , n2599 );
    or g9996 ( n10368 , n5395 , n7915 );
    xnor g9997 ( n10779 , n7378 , n3202 );
    and g9998 ( n863 , n7263 , n12492 );
    xnor g9999 ( n10802 , n13231 , n7644 );
    and g10000 ( n6326 , n1456 , n11610 );
    or g10001 ( n11827 , n12090 , n2611 );
    or g10002 ( n10857 , n6590 , n10029 );
    or g10003 ( n768 , n633 , n1600 );
    xnor g10004 ( n8320 , n7355 , n9259 );
    or g10005 ( n1892 , n8129 , n10319 );
    nor g10006 ( n4228 , n4015 , n7465 );
    nor g10007 ( n12268 , n2403 , n11348 );
    or g10008 ( n1645 , n6110 , n5691 );
    xnor g10009 ( n7173 , n6165 , n2448 );
    or g10010 ( n5305 , n863 , n7559 );
    not g10011 ( n4815 , n6017 );
    or g10012 ( n2778 , n2955 , n8145 );
    or g10013 ( n674 , n8325 , n7221 );
    not g10014 ( n6063 , n6655 );
    xnor g10015 ( n1969 , n10406 , n11126 );
    xnor g10016 ( n13236 , n88 , n11411 );
    and g10017 ( n8602 , n7917 , n2049 );
    xnor g10018 ( n5302 , n661 , n1036 );
    not g10019 ( n13235 , n2948 );
    xnor g10020 ( n2775 , n3977 , n7175 );
    not g10021 ( n10974 , n1916 );
    not g10022 ( n7819 , n12352 );
    not g10023 ( n12508 , n9151 );
    xnor g10024 ( n7477 , n7091 , n10440 );
    xnor g10025 ( n9368 , n10876 , n6645 );
    xnor g10026 ( n7384 , n4586 , n1431 );
    xnor g10027 ( n4647 , n9997 , n9387 );
    nor g10028 ( n8367 , n3511 , n11738 );
    and g10029 ( n10034 , n10230 , n8525 );
    xnor g10030 ( n5064 , n930 , n2055 );
    not g10031 ( n321 , n6826 );
    or g10032 ( n568 , n6190 , n1861 );
    xnor g10033 ( n7646 , n7399 , n11984 );
    or g10034 ( n6614 , n4980 , n10179 );
    and g10035 ( n11890 , n7772 , n4470 );
    not g10036 ( n13063 , n3499 );
    and g10037 ( n9749 , n5752 , n2177 );
    and g10038 ( n6170 , n5697 , n10636 );
    not g10039 ( n9129 , n817 );
    xnor g10040 ( n4037 , n12889 , n171 );
    nor g10041 ( n9713 , n5112 , n1180 );
    xnor g10042 ( n3542 , n8901 , n11552 );
    not g10043 ( n4830 , n6920 );
    not g10044 ( n3259 , n5969 );
    or g10045 ( n7801 , n10571 , n1107 );
    and g10046 ( n12781 , n511 , n12162 );
    or g10047 ( n248 , n8349 , n12823 );
    and g10048 ( n11178 , n2590 , n6392 );
    xnor g10049 ( n8362 , n495 , n461 );
    and g10050 ( n8600 , n8263 , n2988 );
    and g10051 ( n9621 , n12348 , n854 );
    not g10052 ( n9882 , n5536 );
    or g10053 ( n12213 , n766 , n129 );
    or g10054 ( n4600 , n787 , n9223 );
    and g10055 ( n12802 , n4832 , n820 );
    not g10056 ( n11920 , n8506 );
    not g10057 ( n12698 , n2389 );
    not g10058 ( n3505 , n12965 );
    not g10059 ( n9016 , n8332 );
    or g10060 ( n8182 , n2449 , n6265 );
    and g10061 ( n4509 , n5671 , n510 );
    or g10062 ( n8223 , n6245 , n2449 );
    xnor g10063 ( n7236 , n8418 , n1260 );
    xnor g10064 ( n6620 , n1752 , n12367 );
    xnor g10065 ( n5778 , n7725 , n13023 );
    xnor g10066 ( n9876 , n216 , n3772 );
    xnor g10067 ( n2286 , n1409 , n5657 );
    not g10068 ( n338 , n12853 );
    or g10069 ( n4041 , n8079 , n542 );
    and g10070 ( n11828 , n2478 , n10715 );
    or g10071 ( n4306 , n8254 , n12789 );
    not g10072 ( n6499 , n7270 );
    xnor g10073 ( n5798 , n3183 , n11445 );
    and g10074 ( n12519 , n12689 , n4103 );
    nor g10075 ( n12299 , n11189 , n6512 );
    xnor g10076 ( n2845 , n1365 , n11162 );
    xnor g10077 ( n4126 , n10366 , n12474 );
    and g10078 ( n3918 , n8168 , n12944 );
    nor g10079 ( n3877 , n8689 , n8630 );
    or g10080 ( n8680 , n6957 , n9370 );
    not g10081 ( n1354 , n6023 );
    or g10082 ( n4939 , n8796 , n10214 );
    and g10083 ( n7335 , n4108 , n3554 );
    and g10084 ( n2506 , n10908 , n411 );
    not g10085 ( n9913 , n7812 );
    xnor g10086 ( n4035 , n11812 , n1066 );
    or g10087 ( n10599 , n8463 , n12655 );
    nor g10088 ( n7995 , n5622 , n10531 );
    nor g10089 ( n2347 , n2653 , n13111 );
    xnor g10090 ( n10559 , n12993 , n6589 );
    xnor g10091 ( n1909 , n4245 , n5866 );
    xnor g10092 ( n2258 , n8953 , n10930 );
    not g10093 ( n8598 , n499 );
    xnor g10094 ( n7367 , n3612 , n9312 );
    xnor g10095 ( n1397 , n8349 , n10121 );
    xnor g10096 ( n678 , n5056 , n2819 );
    not g10097 ( n8720 , n10162 );
    xnor g10098 ( n11667 , n11826 , n8353 );
    nor g10099 ( n5410 , n6108 , n4091 );
    nor g10100 ( n11486 , n4049 , n11161 );
    xnor g10101 ( n2836 , n3660 , n8958 );
    or g10102 ( n6130 , n10143 , n13238 );
    not g10103 ( n10730 , n9528 );
    and g10104 ( n7147 , n6825 , n6467 );
    xnor g10105 ( n9139 , n5774 , n2236 );
    xnor g10106 ( n11335 , n11652 , n1446 );
    xnor g10107 ( n2646 , n3310 , n4909 );
    or g10108 ( n6738 , n202 , n10106 );
    or g10109 ( n307 , n5520 , n542 );
    xnor g10110 ( n2328 , n4679 , n8085 );
    xnor g10111 ( n3788 , n1475 , n12489 );
    xnor g10112 ( n9322 , n4810 , n3936 );
    and g10113 ( n1687 , n2057 , n2295 );
    or g10114 ( n7151 , n1136 , n716 );
    xnor g10115 ( n10553 , n12936 , n7312 );
    or g10116 ( n3423 , n119 , n6404 );
    and g10117 ( n7866 , n6764 , n13138 );
    not g10118 ( n4420 , n10642 );
    xnor g10119 ( n10061 , n11820 , n9979 );
    xnor g10120 ( n751 , n5868 , n5805 );
    and g10121 ( n10909 , n12775 , n4359 );
    nor g10122 ( n10580 , n9856 , n6101 );
    and g10123 ( n5181 , n8858 , n8194 );
    and g10124 ( n12250 , n8557 , n12756 );
    xnor g10125 ( n6458 , n1087 , n9546 );
    xnor g10126 ( n4263 , n10853 , n1311 );
    or g10127 ( n4791 , n5028 , n2735 );
    not g10128 ( n8153 , n8459 );
    nor g10129 ( n12366 , n9833 , n5746 );
    xor g10130 ( n9805 , n10034 , n2951 );
    or g10131 ( n11191 , n11677 , n2572 );
    xnor g10132 ( n4031 , n12984 , n9646 );
    not g10133 ( n10470 , n11885 );
    or g10134 ( n7277 , n1331 , n11107 );
    or g10135 ( n2464 , n3854 , n11668 );
    xnor g10136 ( n4511 , n4552 , n3324 );
    and g10137 ( n3968 , n9940 , n8397 );
    not g10138 ( n4028 , n7792 );
    or g10139 ( n9365 , n13084 , n479 );
    or g10140 ( n10700 , n5794 , n3512 );
    not g10141 ( n4161 , n287 );
    or g10142 ( n5669 , n5168 , n11107 );
    or g10143 ( n73 , n3129 , n3143 );
    not g10144 ( n5954 , n1978 );
    xnor g10145 ( n6221 , n1745 , n3349 );
    xnor g10146 ( n10709 , n368 , n5891 );
    xnor g10147 ( n506 , n3314 , n9583 );
    xnor g10148 ( n2142 , n5621 , n3043 );
    or g10149 ( n1907 , n10835 , n10843 );
    xnor g10150 ( n9359 , n8627 , n12694 );
    xnor g10151 ( n6597 , n8573 , n12096 );
    and g10152 ( n9076 , n7506 , n10543 );
    and g10153 ( n9049 , n10626 , n8271 );
    not g10154 ( n5688 , n4748 );
    and g10155 ( n12360 , n11115 , n2509 );
    not g10156 ( n11331 , n2751 );
    not g10157 ( n789 , n9216 );
    nor g10158 ( n11277 , n12577 , n2055 );
    not g10159 ( n7805 , n13058 );
    xnor g10160 ( n12214 , n12260 , n3142 );
    or g10161 ( n1096 , n9668 , n10886 );
    or g10162 ( n1256 , n1058 , n3817 );
    not g10163 ( n13080 , n5556 );
    xnor g10164 ( n8151 , n6964 , n4539 );
    or g10165 ( n6685 , n10263 , n7221 );
    xnor g10166 ( n4347 , n1306 , n7753 );
    or g10167 ( n4376 , n6040 , n10179 );
    xor g10168 ( n8805 , n8410 , n10800 );
    and g10169 ( n6758 , n8308 , n4330 );
    not g10170 ( n2670 , n10103 );
    xnor g10171 ( n6759 , n2638 , n415 );
    or g10172 ( n4096 , n2527 , n2030 );
    xnor g10173 ( n12473 , n7299 , n4082 );
    or g10174 ( n12682 , n3225 , n6041 );
    or g10175 ( n626 , n2889 , n121 );
    or g10176 ( n8240 , n6419 , n11107 );
    or g10177 ( n1639 , n3982 , n752 );
    or g10178 ( n7310 , n9383 , n2958 );
    or g10179 ( n7271 , n10400 , n8348 );
    or g10180 ( n13068 , n1235 , n8673 );
    or g10181 ( n11552 , n12416 , n10029 );
    xnor g10182 ( n9087 , n2948 , n8155 );
    or g10183 ( n12150 , n3866 , n2675 );
    or g10184 ( n10160 , n6438 , n7530 );
    xnor g10185 ( n7431 , n4304 , n11885 );
    not g10186 ( n11842 , n10615 );
    xnor g10187 ( n6027 , n11896 , n7120 );
    or g10188 ( n8216 , n3302 , n8133 );
    not g10189 ( n13181 , n937 );
    nor g10190 ( n244 , n13093 , n4338 );
    or g10191 ( n349 , n9919 , n6635 );
    and g10192 ( n4523 , n2520 , n255 );
    or g10193 ( n934 , n5914 , n3356 );
    or g10194 ( n10208 , n11628 , n8563 );
    xnor g10195 ( n5316 , n5943 , n12929 );
    nor g10196 ( n5019 , n12422 , n10198 );
    or g10197 ( n7390 , n1214 , n9418 );
    not g10198 ( n6968 , n3669 );
    not g10199 ( n5971 , n11766 );
    or g10200 ( n3282 , n11319 , n4067 );
    buf g10201 ( n9195 , n11418 );
    not g10202 ( n8131 , n2252 );
    and g10203 ( n84 , n6503 , n310 );
    or g10204 ( n136 , n9339 , n10029 );
    or g10205 ( n7261 , n10136 , n3174 );
    or g10206 ( n2267 , n5835 , n3488 );
    and g10207 ( n3903 , n5586 , n3832 );
    nor g10208 ( n8371 , n229 , n651 );
    not g10209 ( n11975 , n11288 );
    xnor g10210 ( n5735 , n6566 , n6969 );
    xor g10211 ( n6451 , n13106 , n7447 );
    xnor g10212 ( n9219 , n3711 , n8294 );
    nor g10213 ( n11268 , n10254 , n4730 );
    xnor g10214 ( n1034 , n1835 , n11349 );
    nor g10215 ( n10953 , n12259 , n3048 );
    or g10216 ( n10228 , n122 , n6062 );
    xor g10217 ( n11893 , n12614 , n864 );
    xnor g10218 ( n3991 , n404 , n6759 );
    and g10219 ( n8418 , n8790 , n10312 );
    and g10220 ( n8235 , n5954 , n3168 );
    and g10221 ( n11375 , n2677 , n10912 );
    nor g10222 ( n2878 , n9387 , n9997 );
    not g10223 ( n6721 , n11891 );
    and g10224 ( n6853 , n1779 , n10132 );
    or g10225 ( n1087 , n7234 , n8702 );
    not g10226 ( n530 , n4987 );
    or g10227 ( n12793 , n6191 , n1894 );
    not g10228 ( n8339 , n11559 );
    xnor g10229 ( n2864 , n2100 , n12220 );
    and g10230 ( n670 , n1220 , n3878 );
    xnor g10231 ( n12038 , n664 , n3968 );
    xnor g10232 ( n6955 , n3265 , n1433 );
    xnor g10233 ( n7818 , n9065 , n3332 );
    and g10234 ( n1239 , n12281 , n1698 );
    not g10235 ( n5959 , n7806 );
    and g10236 ( n10002 , n9732 , n854 );
    and g10237 ( n3732 , n6414 , n12770 );
    or g10238 ( n7946 , n8327 , n3374 );
    and g10239 ( n13023 , n7022 , n3656 );
    xnor g10240 ( n9746 , n10395 , n102 );
    xnor g10241 ( n8357 , n10294 , n8283 );
    xnor g10242 ( n10613 , n10549 , n3693 );
    or g10243 ( n10949 , n406 , n7998 );
    or g10244 ( n7281 , n11218 , n2059 );
    xnor g10245 ( n2697 , n10475 , n7021 );
    xnor g10246 ( n6340 , n10718 , n10124 );
    buf g10247 ( n9223 , n12954 );
    nor g10248 ( n10723 , n12152 , n7735 );
    or g10249 ( n2224 , n12754 , n11714 );
    not g10250 ( n10849 , n12822 );
    xnor g10251 ( n10767 , n9101 , n2214 );
    or g10252 ( n125 , n9039 , n10466 );
    xor g10253 ( n2465 , n3361 , n4908 );
    xnor g10254 ( n1146 , n5727 , n13175 );
    or g10255 ( n3983 , n11352 , n10029 );
    and g10256 ( n1466 , n12613 , n375 );
    xnor g10257 ( n13158 , n12296 , n10096 );
    or g10258 ( n4438 , n12493 , n11668 );
    xnor g10259 ( n10027 , n6992 , n10297 );
    xnor g10260 ( n7308 , n9240 , n10659 );
    not g10261 ( n3911 , n11180 );
    or g10262 ( n12913 , n121 , n4960 );
    not g10263 ( n8498 , n10162 );
    xnor g10264 ( n3244 , n1524 , n6873 );
    or g10265 ( n6509 , n13168 , n2544 );
    nor g10266 ( n12981 , n8085 , n4679 );
    or g10267 ( n3028 , n75 , n8024 );
    or g10268 ( n11249 , n7970 , n3075 );
    xnor g10269 ( n4329 , n8273 , n4156 );
    and g10270 ( n11606 , n9199 , n11192 );
    or g10271 ( n12938 , n3489 , n3715 );
    and g10272 ( n10364 , n9987 , n7901 );
    xnor g10273 ( n10917 , n6240 , n7211 );
    or g10274 ( n11024 , n11514 , n8777 );
    xnor g10275 ( n984 , n3123 , n9212 );
    or g10276 ( n2182 , n1515 , n7004 );
    xnor g10277 ( n4233 , n11133 , n1291 );
    xnor g10278 ( n707 , n2811 , n11250 );
    and g10279 ( n13210 , n11704 , n2348 );
    and g10280 ( n7610 , n3636 , n10341 );
    nor g10281 ( n8342 , n2476 , n2510 );
    not g10282 ( n6182 , n6937 );
    nor g10283 ( n1450 , n2616 , n5285 );
    not g10284 ( n1058 , n510 );
    not g10285 ( n1030 , n4017 );
    not g10286 ( n9160 , n12892 );
    xnor g10287 ( n2460 , n9099 , n245 );
    and g10288 ( n11202 , n11236 , n411 );
    not g10289 ( n1936 , n3566 );
    or g10290 ( n7634 , n5733 , n10474 );
    or g10291 ( n2960 , n7038 , n1833 );
    or g10292 ( n13090 , n10112 , n5076 );
    xnor g10293 ( n8282 , n11804 , n4548 );
    xnor g10294 ( n6328 , n2659 , n2736 );
    and g10295 ( n11086 , n1747 , n11423 );
    xnor g10296 ( n12118 , n7637 , n5038 );
    or g10297 ( n11493 , n10857 , n8793 );
    nor g10298 ( n9002 , n10796 , n12058 );
    xnor g10299 ( n5078 , n8292 , n13090 );
    not g10300 ( n9238 , n469 );
    xnor g10301 ( n2684 , n12974 , n10038 );
    and g10302 ( n3862 , n5490 , n10740 );
    xnor g10303 ( n5075 , n9324 , n4090 );
    nor g10304 ( n1840 , n12873 , n8756 );
    or g10305 ( n6844 , n1323 , n12062 );
    and g10306 ( n258 , n3019 , n11987 );
    or g10307 ( n1990 , n2899 , n11910 );
    xnor g10308 ( n4631 , n1276 , n184 );
    and g10309 ( n507 , n2243 , n4311 );
    and g10310 ( n2546 , n7056 , n7432 );
    or g10311 ( n6688 , n12032 , n8490 );
    not g10312 ( n7223 , n3677 );
    and g10313 ( n8352 , n2530 , n12473 );
    or g10314 ( n6422 , n6881 , n10702 );
    or g10315 ( n9146 , n13190 , n206 );
    xor g10316 ( n1875 , n4135 , n12612 );
    or g10317 ( n11330 , n9698 , n4023 );
    not g10318 ( n10989 , n12939 );
    or g10319 ( n10013 , n9429 , n4640 );
    and g10320 ( n1371 , n6934 , n3871 );
    not g10321 ( n2875 , n11537 );
    or g10322 ( n12525 , n7566 , n2766 );
    not g10323 ( n1885 , n3977 );
    not g10324 ( n11172 , n4102 );
    not g10325 ( n5970 , n5786 );
    and g10326 ( n10823 , n3957 , n11273 );
    or g10327 ( n11372 , n2449 , n8490 );
    not g10328 ( n7158 , n6085 );
    and g10329 ( n4508 , n8974 , n10726 );
    xnor g10330 ( n2981 , n1373 , n10721 );
    and g10331 ( n7153 , n7073 , n1477 );
    or g10332 ( n5132 , n10527 , n11107 );
    not g10333 ( n12624 , n10238 );
    xnor g10334 ( n2976 , n9502 , n2719 );
    not g10335 ( n8374 , n510 );
    xnor g10336 ( n5686 , n4171 , n5173 );
    nor g10337 ( n7077 , n8279 , n802 );
    and g10338 ( n145 , n12058 , n10796 );
    and g10339 ( n9575 , n11996 , n12650 );
    xnor g10340 ( n7670 , n2006 , n6325 );
    or g10341 ( n10741 , n12775 , n4359 );
    xnor g10342 ( n12715 , n10671 , n1927 );
    and g10343 ( n12934 , n1791 , n1886 );
    and g10344 ( n9067 , n11614 , n3536 );
    not g10345 ( n7247 , n5470 );
    or g10346 ( n373 , n10824 , n9923 );
    and g10347 ( n7137 , n4361 , n4563 );
    and g10348 ( n11021 , n3458 , n4475 );
    nor g10349 ( n8643 , n8923 , n7479 );
    not g10350 ( n9804 , n11567 );
    not g10351 ( n1438 , n10594 );
    or g10352 ( n2162 , n1513 , n2298 );
    not g10353 ( n5489 , n5590 );
    or g10354 ( n7886 , n12353 , n8316 );
    or g10355 ( n10370 , n6231 , n12273 );
    xnor g10356 ( n4120 , n10155 , n11080 );
    xnor g10357 ( n2459 , n2854 , n2853 );
    or g10358 ( n8541 , n10897 , n1856 );
    and g10359 ( n10502 , n8664 , n10161 );
    nor g10360 ( n3474 , n4538 , n12450 );
    not g10361 ( n1145 , n4681 );
    or g10362 ( n10555 , n2614 , n5076 );
    and g10363 ( n4044 , n6823 , n3255 );
    and g10364 ( n5753 , n11515 , n1542 );
    nor g10365 ( n3574 , n3131 , n7627 );
    xnor g10366 ( n1734 , n4706 , n7851 );
    not g10367 ( n10305 , n7778 );
    or g10368 ( n7037 , n10608 , n3618 );
    nor g10369 ( n11935 , n10282 , n5859 );
    not g10370 ( n6160 , n3774 );
    or g10371 ( n11476 , n8384 , n10098 );
    nor g10372 ( n11912 , n10328 , n10366 );
    and g10373 ( n5889 , n5773 , n12600 );
    and g10374 ( n5524 , n8120 , n9334 );
    xor g10375 ( n12102 , n3110 , n7083 );
    and g10376 ( n6607 , n6046 , n2333 );
    nor g10377 ( n4637 , n6844 , n11085 );
    or g10378 ( n7612 , n845 , n9075 );
    or g10379 ( n3699 , n6506 , n7865 );
    xnor g10380 ( n10463 , n12850 , n2632 );
    nor g10381 ( n9179 , n3387 , n12115 );
    and g10382 ( n2501 , n10997 , n3996 );
    xnor g10383 ( n9982 , n6075 , n10821 );
    not g10384 ( n11379 , n8291 );
    not g10385 ( n10948 , n10172 );
    or g10386 ( n12660 , n11982 , n10764 );
    xnor g10387 ( n1753 , n4489 , n10968 );
    or g10388 ( n8932 , n2757 , n6001 );
    or g10389 ( n6254 , n6769 , n12388 );
    not g10390 ( n12713 , n10378 );
    xnor g10391 ( n9950 , n5371 , n2441 );
    nor g10392 ( n5836 , n7527 , n8913 );
    not g10393 ( n11910 , n951 );
    xnor g10394 ( n6105 , n544 , n6025 );
    xnor g10395 ( n5975 , n5497 , n1387 );
    nor g10396 ( n10404 , n5998 , n3173 );
    and g10397 ( n7656 , n7415 , n3436 );
    or g10398 ( n337 , n3647 , n5098 );
    xnor g10399 ( n8031 , n2798 , n4670 );
    or g10400 ( n1842 , n4808 , n8534 );
    and g10401 ( n2280 , n10422 , n12773 );
    or g10402 ( n12659 , n10471 , n5242 );
    or g10403 ( n3056 , n3900 , n5443 );
    xnor g10404 ( n4712 , n7534 , n7212 );
    not g10405 ( n7086 , n8824 );
    and g10406 ( n2891 , n2471 , n165 );
    xnor g10407 ( n11348 , n2475 , n9574 );
    or g10408 ( n5963 , n1261 , n7935 );
    or g10409 ( n1735 , n6770 , n10319 );
    not g10410 ( n5853 , n5140 );
    xnor g10411 ( n7948 , n1368 , n10042 );
    nor g10412 ( n12588 , n215 , n10629 );
    xnor g10413 ( n2577 , n11845 , n7057 );
    xnor g10414 ( n7858 , n3480 , n2859 );
    and g10415 ( n1046 , n3539 , n12446 );
    xnor g10416 ( n2565 , n3980 , n3714 );
    or g10417 ( n297 , n6517 , n6493 );
    or g10418 ( n12720 , n4166 , n1570 );
    nor g10419 ( n215 , n2024 , n6508 );
    or g10420 ( n10994 , n1989 , n6770 );
    and g10421 ( n1986 , n10889 , n10498 );
    or g10422 ( n4720 , n9637 , n5188 );
    or g10423 ( n12184 , n7783 , n6265 );
    xnor g10424 ( n7393 , n4345 , n12570 );
    not g10425 ( n11237 , n6701 );
    not g10426 ( n2287 , n8230 );
    xnor g10427 ( n5232 , n7896 , n851 );
    not g10428 ( n4498 , n5546 );
    and g10429 ( n9151 , n4638 , n7453 );
    not g10430 ( n1434 , n8332 );
    and g10431 ( n9704 , n867 , n9326 );
    or g10432 ( n1876 , n11548 , n1985 );
    not g10433 ( n3817 , n2590 );
    xnor g10434 ( n3455 , n4600 , n1723 );
    nor g10435 ( n12631 , n7439 , n10963 );
    xnor g10436 ( n6819 , n12845 , n13087 );
    or g10437 ( n6880 , n13039 , n2133 );
    or g10438 ( n5976 , n1875 , n12366 );
    not g10439 ( n2403 , n13121 );
    nor g10440 ( n12400 , n1774 , n8413 );
    xnor g10441 ( n13155 , n10547 , n7689 );
    not g10442 ( n9897 , n4126 );
    and g10443 ( n12832 , n3662 , n6664 );
    or g10444 ( n12427 , n3091 , n2083 );
    not g10445 ( n1579 , n10075 );
    not g10446 ( n12838 , n10582 );
    not g10447 ( n7377 , n5962 );
    or g10448 ( n3692 , n13025 , n2059 );
    not g10449 ( n10872 , n4906 );
    or g10450 ( n12179 , n11779 , n7254 );
    xnor g10451 ( n11306 , n5357 , n3887 );
    not g10452 ( n713 , n6647 );
    or g10453 ( n5577 , n9564 , n5029 );
    xnor g10454 ( n6007 , n6388 , n6243 );
    xnor g10455 ( n236 , n1334 , n11176 );
    xnor g10456 ( n1309 , n9066 , n7681 );
    not g10457 ( n9172 , n2073 );
    or g10458 ( n5072 , n9069 , n8268 );
    xor g10459 ( n4349 , n4376 , n11813 );
    xnor g10460 ( n1844 , n7754 , n775 );
    xnor g10461 ( n12598 , n9922 , n6031 );
    xnor g10462 ( n12439 , n9083 , n4390 );
    not g10463 ( n5554 , n748 );
    not g10464 ( n5001 , n8559 );
    or g10465 ( n5693 , n12573 , n4640 );
    xnor g10466 ( n9579 , n6079 , n1293 );
    xnor g10467 ( n11353 , n7067 , n5979 );
    or g10468 ( n6976 , n6657 , n265 );
    xnor g10469 ( n8897 , n5693 , n667 );
    not g10470 ( n12535 , n4042 );
    xnor g10471 ( n384 , n12933 , n6158 );
    and g10472 ( n1452 , n8610 , n12521 );
    nor g10473 ( n7004 , n2251 , n665 );
    or g10474 ( n932 , n5655 , n2206 );
    not g10475 ( n5666 , n6392 );
    not g10476 ( n1035 , n353 );
    and g10477 ( n1603 , n3570 , n7898 );
    not g10478 ( n10281 , n1650 );
    xnor g10479 ( n4535 , n300 , n10619 );
    xor g10480 ( n6677 , n6956 , n2583 );
    or g10481 ( n451 , n11779 , n4640 );
    xnor g10482 ( n11031 , n5421 , n11806 );
    xnor g10483 ( n11405 , n3747 , n999 );
    or g10484 ( n8093 , n3550 , n5059 );
    not g10485 ( n13133 , n7465 );
    and g10486 ( n4353 , n1867 , n1448 );
    or g10487 ( n11459 , n161 , n12328 );
    xnor g10488 ( n557 , n12448 , n7838 );
    not g10489 ( n6652 , n4645 );
    not g10490 ( n3861 , n3913 );
    and g10491 ( n10551 , n10094 , n147 );
    not g10492 ( n5645 , n10805 );
    nor g10493 ( n2087 , n9797 , n12584 );
    xnor g10494 ( n3296 , n7891 , n6693 );
    and g10495 ( n315 , n12585 , n6315 );
    xnor g10496 ( n6678 , n12235 , n1253 );
    xnor g10497 ( n9800 , n5933 , n6670 );
    or g10498 ( n12953 , n1035 , n6732 );
    or g10499 ( n4261 , n4974 , n5076 );
    or g10500 ( n1654 , n3587 , n4947 );
    and g10501 ( n7279 , n8139 , n10606 );
    and g10502 ( n8520 , n3316 , n5411 );
    or g10503 ( n11273 , n2639 , n8490 );
    or g10504 ( n5206 , n9131 , n10871 );
    or g10505 ( n8165 , n2109 , n488 );
    not g10506 ( n6716 , n68 );
    or g10507 ( n4180 , n983 , n9177 );
    not g10508 ( n7914 , n8818 );
    or g10509 ( n4930 , n8335 , n2675 );
    xnor g10510 ( n1282 , n11556 , n3745 );
    or g10511 ( n6664 , n12241 , n9055 );
    xnor g10512 ( n9136 , n9565 , n4597 );
    not g10513 ( n735 , n1528 );
    or g10514 ( n4314 , n4610 , n479 );
    not g10515 ( n12166 , n11324 );
    nor g10516 ( n6443 , n12167 , n2927 );
    xor g10517 ( n7290 , n72 , n9250 );
    or g10518 ( n3113 , n7780 , n1144 );
    nor g10519 ( n8099 , n5327 , n4421 );
    and g10520 ( n11959 , n1311 , n10853 );
    xnor g10521 ( n67 , n3899 , n4195 );
    buf g10522 ( n7935 , n9558 );
    or g10523 ( n1373 , n8727 , n6824 );
    or g10524 ( n8829 , n2236 , n5774 );
    or g10525 ( n10577 , n13028 , n6173 );
    not g10526 ( n1695 , n7720 );
    xnor g10527 ( n10151 , n13188 , n1288 );
    nor g10528 ( n2042 , n2486 , n979 );
    not g10529 ( n7480 , n11129 );
    not g10530 ( n10021 , n11891 );
    or g10531 ( n5564 , n11099 , n10689 );
    or g10532 ( n9152 , n10688 , n10759 );
    not g10533 ( n2890 , n13058 );
    or g10534 ( n11366 , n6751 , n1463 );
    nor g10535 ( n6078 , n8476 , n10027 );
    not g10536 ( n3999 , n5962 );
    nor g10537 ( n5690 , n7457 , n3117 );
    not g10538 ( n10586 , n11411 );
    xnor g10539 ( n11971 , n11199 , n4601 );
    and g10540 ( n7244 , n5166 , n10536 );
    or g10541 ( n1601 , n5616 , n4055 );
    xnor g10542 ( n3810 , n5763 , n459 );
    xnor g10543 ( n4670 , n7265 , n12100 );
    xor g10544 ( n12054 , n8715 , n6921 );
    or g10545 ( n8873 , n3802 , n12189 );
    not g10546 ( n1493 , n2169 );
    xor g10547 ( n5556 , n9904 , n12915 );
    and g10548 ( n8090 , n9079 , n920 );
    and g10549 ( n8537 , n5090 , n7638 );
    xnor g10550 ( n7744 , n1262 , n5235 );
    not g10551 ( n10941 , n8422 );
    not g10552 ( n12573 , n11891 );
    not g10553 ( n12377 , n8798 );
    xnor g10554 ( n10478 , n5556 , n6073 );
    or g10555 ( n272 , n9399 , n13031 );
    or g10556 ( n3060 , n11790 , n7574 );
    not g10557 ( n9681 , n12810 );
    xnor g10558 ( n1369 , n2289 , n4569 );
    or g10559 ( n10145 , n8457 , n9972 );
    or g10560 ( n9287 , n6922 , n6635 );
    or g10561 ( n8171 , n10287 , n12847 );
    or g10562 ( n12652 , n1447 , n6404 );
    xnor g10563 ( n4586 , n1233 , n10632 );
    xnor g10564 ( n1291 , n941 , n4071 );
    or g10565 ( n6302 , n6383 , n1570 );
    not g10566 ( n4203 , n9841 );
    xnor g10567 ( n1334 , n6167 , n5981 );
    nor g10568 ( n11695 , n1742 , n8475 );
    and g10569 ( n11813 , n8466 , n8506 );
    xnor g10570 ( n13120 , n7752 , n9274 );
    or g10571 ( n4795 , n5561 , n2315 );
    or g10572 ( n3687 , n3331 , n952 );
    xnor g10573 ( n5266 , n13040 , n859 );
    or g10574 ( n12309 , n10492 , n6138 );
    or g10575 ( n8769 , n9298 , n8127 );
    or g10576 ( n4542 , n10929 , n7723 );
    and g10577 ( n8437 , n204 , n5572 );
    xnor g10578 ( n8752 , n5546 , n13044 );
    or g10579 ( n8780 , n8329 , n5797 );
    and g10580 ( n10315 , n980 , n11297 );
    not g10581 ( n2717 , n10541 );
    and g10582 ( n5387 , n842 , n4274 );
    or g10583 ( n3515 , n946 , n12501 );
    xnor g10584 ( n6282 , n1206 , n2714 );
    nor g10585 ( n612 , n2743 , n1620 );
    and g10586 ( n7320 , n8142 , n4443 );
    or g10587 ( n12047 , n8759 , n13148 );
    and g10588 ( n4112 , n6495 , n12315 );
    xnor g10589 ( n6174 , n12151 , n12540 );
    or g10590 ( n9924 , n5271 , n6404 );
    or g10591 ( n3001 , n10411 , n4208 );
    not g10592 ( n1194 , n8163 );
    xnor g10593 ( n5464 , n12638 , n736 );
    nor g10594 ( n7578 , n8538 , n12200 );
    not g10595 ( n7188 , n510 );
    xnor g10596 ( n11472 , n5913 , n10379 );
    and g10597 ( n13173 , n761 , n3085 );
    not g10598 ( n8693 , n5307 );
    or g10599 ( n5793 , n5107 , n119 );
    and g10600 ( n12756 , n8123 , n3373 );
    xnor g10601 ( n8945 , n3578 , n4766 );
    nor g10602 ( n4633 , n12127 , n5196 );
    buf g10603 ( n6732 , n8160 );
    xnor g10604 ( n8483 , n3397 , n11459 );
    or g10605 ( n7361 , n6205 , n425 );
    or g10606 ( n891 , n12629 , n4936 );
    and g10607 ( n1306 , n12576 , n7817 );
    not g10608 ( n7084 , n817 );
    xnor g10609 ( n8573 , n12485 , n1309 );
    or g10610 ( n9690 , n11499 , n10909 );
    or g10611 ( n9584 , n9499 , n1381 );
    not g10612 ( n1437 , n11376 );
    or g10613 ( n2331 , n5809 , n9759 );
    not g10614 ( n7883 , n10620 );
    or g10615 ( n3256 , n3295 , n4751 );
    buf g10616 ( n1463 , n3058 );
    xnor g10617 ( n1403 , n10324 , n7202 );
    xnor g10618 ( n13050 , n9863 , n11128 );
    not g10619 ( n11628 , n5920 );
    xnor g10620 ( n134 , n68 , n6246 );
    xnor g10621 ( n669 , n8972 , n6125 );
    xnor g10622 ( n7698 , n2340 , n1386 );
    and g10623 ( n6496 , n7629 , n3197 );
    or g10624 ( n5361 , n11705 , n11893 );
    or g10625 ( n9994 , n10714 , n10319 );
    xnor g10626 ( n6427 , n2372 , n9785 );
    xnor g10627 ( n823 , n12660 , n6435 );
    not g10628 ( n8317 , n3379 );
    xnor g10629 ( n11992 , n9037 , n7599 );
    not g10630 ( n12998 , n10873 );
    not g10631 ( n757 , n4417 );
    xnor g10632 ( n10475 , n11676 , n2483 );
    not g10633 ( n11143 , n8564 );
    or g10634 ( n9140 , n6384 , n10417 );
    or g10635 ( n5452 , n12786 , n8268 );
    and g10636 ( n8387 , n10590 , n10483 );
    not g10637 ( n956 , n10451 );
    and g10638 ( n8762 , n8728 , n4518 );
    xnor g10639 ( n10630 , n9466 , n13120 );
    xnor g10640 ( n10728 , n12356 , n3734 );
    and g10641 ( n9986 , n3172 , n1773 );
    or g10642 ( n4135 , n4465 , n4373 );
    and g10643 ( n6119 , n7215 , n249 );
    and g10644 ( n2115 , n692 , n12676 );
    not g10645 ( n2129 , n8860 );
    and g10646 ( n11641 , n7772 , n9531 );
    xnor g10647 ( n11572 , n8180 , n4872 );
    xnor g10648 ( n9872 , n259 , n10227 );
    or g10649 ( n5736 , n2581 , n12328 );
    or g10650 ( n12448 , n11757 , n8490 );
    not g10651 ( n8585 , n2758 );
    xnor g10652 ( n3142 , n1608 , n12398 );
    or g10653 ( n331 , n11054 , n12188 );
    and g10654 ( n4326 , n8599 , n6468 );
    or g10655 ( n9559 , n6112 , n7935 );
    xnor g10656 ( n2502 , n11022 , n3343 );
    xnor g10657 ( n1473 , n12390 , n1300 );
    and g10658 ( n7676 , n4991 , n10066 );
    xnor g10659 ( n774 , n10949 , n7122 );
    xnor g10660 ( n3947 , n9956 , n10775 );
    or g10661 ( n5523 , n4080 , n11300 );
    xnor g10662 ( n11861 , n4866 , n908 );
    xnor g10663 ( n3268 , n112 , n10003 );
    and g10664 ( n6352 , n12114 , n2186 );
    xnor g10665 ( n7296 , n12601 , n9036 );
    nor g10666 ( n766 , n9992 , n10630 );
    not g10667 ( n5714 , n7183 );
    nor g10668 ( n4504 , n8137 , n4740 );
    or g10669 ( n11650 , n10381 , n7824 );
    or g10670 ( n730 , n7272 , n3918 );
    and g10671 ( n11555 , n5953 , n12712 );
    nor g10672 ( n10840 , n6797 , n3294 );
    and g10673 ( n7501 , n9304 , n6475 );
    and g10674 ( n12176 , n1440 , n8741 );
    xnor g10675 ( n7863 , n888 , n2765 );
    not g10676 ( n10512 , n3412 );
    and g10677 ( n3447 , n1520 , n10145 );
    not g10678 ( n6052 , n8319 );
    xor g10679 ( n8811 , n10577 , n3995 );
    not g10680 ( n10898 , n1307 );
    and g10681 ( n1798 , n11030 , n9531 );
    xnor g10682 ( n5585 , n5234 , n11201 );
    xnor g10683 ( n7842 , n10973 , n2761 );
    or g10684 ( n8310 , n9626 , n130 );
    not g10685 ( n13084 , n5884 );
    xnor g10686 ( n5273 , n12442 , n9839 );
    or g10687 ( n3662 , n8102 , n5258 );
    and g10688 ( n6670 , n1138 , n8125 );
    or g10689 ( n9102 , n10545 , n11639 );
    xnor g10690 ( n12074 , n6823 , n9857 );
    or g10691 ( n8999 , n3758 , n164 );
    not g10692 ( n1113 , n4006 );
    nor g10693 ( n4554 , n1877 , n1429 );
    or g10694 ( n8975 , n6305 , n984 );
    and g10695 ( n5472 , n9150 , n8743 );
    and g10696 ( n7305 , n7566 , n2766 );
    and g10697 ( n630 , n5307 , n4036 );
    not g10698 ( n4618 , n10946 );
    xnor g10699 ( n8916 , n9648 , n955 );
    or g10700 ( n8853 , n7523 , n7975 );
    and g10701 ( n2651 , n9605 , n1054 );
    and g10702 ( n2377 , n10260 , n5916 );
    and g10703 ( n6714 , n1257 , n6845 );
    or g10704 ( n7969 , n4875 , n12328 );
    xnor g10705 ( n2874 , n4578 , n4150 );
    and g10706 ( n4708 , n906 , n2056 );
    or g10707 ( n4178 , n12552 , n10213 );
    xnor g10708 ( n5380 , n10023 , n11042 );
    xnor g10709 ( n1204 , n5918 , n811 );
    not g10710 ( n11700 , n7491 );
    or g10711 ( n7797 , n11751 , n617 );
    xnor g10712 ( n4247 , n12321 , n5781 );
    or g10713 ( n6659 , n8009 , n6628 );
    or g10714 ( n3528 , n7049 , n8563 );
    or g10715 ( n11945 , n3307 , n5566 );
    xnor g10716 ( n11064 , n2451 , n9034 );
    and g10717 ( n8118 , n3822 , n3339 );
    or g10718 ( n9819 , n8817 , n9159 );
    not g10719 ( n13082 , n2174 );
    xnor g10720 ( n1362 , n4968 , n756 );
    or g10721 ( n4475 , n13183 , n177 );
    xnor g10722 ( n3666 , n9269 , n515 );
    nor g10723 ( n4887 , n12606 , n7020 );
    or g10724 ( n5508 , n10452 , n6243 );
    not g10725 ( n8491 , n10979 );
    nor g10726 ( n2489 , n3959 , n4286 );
    xnor g10727 ( n9077 , n6852 , n6307 );
    and g10728 ( n11494 , n9546 , n1087 );
    nor g10729 ( n3990 , n3606 , n7869 );
    and g10730 ( n6093 , n10351 , n8448 );
    not g10731 ( n803 , n11990 );
    or g10732 ( n9442 , n4855 , n10319 );
    not g10733 ( n3418 , n3319 );
    and g10734 ( n9847 , n8139 , n12965 );
    or g10735 ( n10584 , n1741 , n9537 );
    not g10736 ( n9668 , n6826 );
    and g10737 ( n9114 , n7498 , n4225 );
    not g10738 ( n6290 , n1421 );
    not g10739 ( n12808 , n6607 );
    xnor g10740 ( n927 , n12784 , n6620 );
    or g10741 ( n4158 , n1663 , n2415 );
    xnor g10742 ( n6153 , n5274 , n11296 );
    not g10743 ( n10798 , n2295 );
    not g10744 ( n8900 , n818 );
    xnor g10745 ( n11326 , n11414 , n12354 );
    not g10746 ( n7847 , n10575 );
    not g10747 ( n10587 , n5729 );
    xnor g10748 ( n9777 , n9796 , n2040 );
    xnor g10749 ( n1399 , n11125 , n10249 );
    xnor g10750 ( n3746 , n5711 , n6895 );
    xnor g10751 ( n12193 , n1137 , n6899 );
    nor g10752 ( n3148 , n2053 , n7834 );
    xnor g10753 ( n10538 , n5509 , n12875 );
    or g10754 ( n12257 , n8732 , n3882 );
    xnor g10755 ( n11062 , n10640 , n3382 );
    or g10756 ( n12679 , n1634 , n9745 );
    not g10757 ( n4792 , n10451 );
    xnor g10758 ( n5764 , n8008 , n12113 );
    and g10759 ( n9215 , n5031 , n510 );
    not g10760 ( n1624 , n5796 );
    and g10761 ( n5055 , n5568 , n5729 );
    or g10762 ( n3117 , n2582 , n2816 );
    or g10763 ( n9411 , n6416 , n9075 );
    not g10764 ( n8739 , n4978 );
    or g10765 ( n9612 , n7748 , n4373 );
    xnor g10766 ( n11561 , n5306 , n7428 );
    xnor g10767 ( n9196 , n4263 , n11816 );
    or g10768 ( n7156 , n8776 , n6769 );
    xnor g10769 ( n2560 , n2049 , n7917 );
    or g10770 ( n4103 , n12236 , n4835 );
    or g10771 ( n4629 , n6215 , n10433 );
    not g10772 ( n4013 , n2057 );
    and g10773 ( n2255 , n10248 , n5369 );
    and g10774 ( n12725 , n5826 , n2831 );
    not g10775 ( n7719 , n7439 );
    xnor g10776 ( n5060 , n9048 , n6105 );
    or g10777 ( n3204 , n3634 , n1043 );
    or g10778 ( n12569 , n11117 , n8445 );
    or g10779 ( n3878 , n3176 , n10652 );
    not g10780 ( n3696 , n1432 );
    or g10781 ( n3937 , n4475 , n3458 );
    or g10782 ( n5252 , n10153 , n3650 );
    xnor g10783 ( n4711 , n9955 , n3562 );
    xor g10784 ( n4303 , n1719 , n2423 );
    and g10785 ( n2006 , n5671 , n8506 );
    and g10786 ( n11995 , n3922 , n2428 );
    xnor g10787 ( n1086 , n31 , n8872 );
    or g10788 ( n12964 , n11960 , n9075 );
    xnor g10789 ( n2044 , n5451 , n7569 );
    nor g10790 ( n9874 , n6151 , n5033 );
    xnor g10791 ( n6904 , n11692 , n7309 );
    or g10792 ( n7743 , n1087 , n9546 );
    or g10793 ( n1002 , n1909 , n3955 );
    or g10794 ( n7987 , n4739 , n4675 );
    xnor g10795 ( n3923 , n7875 , n4856 );
    not g10796 ( n9131 , n1302 );
    nor g10797 ( n1865 , n9423 , n3206 );
    or g10798 ( n11786 , n7062 , n12273 );
    xnor g10799 ( n12977 , n11168 , n13105 );
    or g10800 ( n6414 , n7042 , n9078 );
    and g10801 ( n6525 , n803 , n8558 );
    xnor g10802 ( n3889 , n5678 , n8684 );
    not g10803 ( n7009 , n10457 );
    not g10804 ( n1697 , n1938 );
    not g10805 ( n8428 , n10398 );
    nor g10806 ( n2574 , n7529 , n7715 );
    or g10807 ( n931 , n4564 , n3949 );
    xnor g10808 ( n10071 , n9903 , n3644 );
    or g10809 ( n7309 , n542 , n11668 );
    xnor g10810 ( n10995 , n4057 , n10994 );
    and g10811 ( n4450 , n6029 , n2179 );
    not g10812 ( n10465 , n7659 );
    xnor g10813 ( n11474 , n7330 , n11760 );
    or g10814 ( n5428 , n7142 , n6265 );
    and g10815 ( n7556 , n812 , n9717 );
    not g10816 ( n16 , n12348 );
    xnor g10817 ( n7540 , n8827 , n6378 );
    xnor g10818 ( n3123 , n10828 , n5651 );
    xnor g10819 ( n807 , n3274 , n49 );
    and g10820 ( n6515 , n4908 , n11545 );
    buf g10821 ( n2544 , n8640 );
    and g10822 ( n6034 , n1453 , n8216 );
    xnor g10823 ( n10218 , n2054 , n4575 );
    and g10824 ( n10038 , n5893 , n3124 );
    not g10825 ( n6407 , n834 );
    xnor g10826 ( n4048 , n8483 , n3881 );
    and g10827 ( n10482 , n13071 , n2419 );
    or g10828 ( n1864 , n6967 , n12328 );
    or g10829 ( n8008 , n1511 , n1026 );
    and g10830 ( n2146 , n1544 , n7611 );
    nor g10831 ( n8450 , n5568 , n8308 );
    or g10832 ( n13067 , n8020 , n7530 );
    xnor g10833 ( n6891 , n8141 , n11510 );
    xnor g10834 ( n6695 , n8559 , n1623 );
    or g10835 ( n7618 , n80 , n1571 );
    xnor g10836 ( n9433 , n8224 , n7449 );
    and g10837 ( n2234 , n2155 , n6291 );
    or g10838 ( n6813 , n6587 , n2675 );
    and g10839 ( n994 , n2188 , n3265 );
    xnor g10840 ( n3434 , n7038 , n10621 );
    xnor g10841 ( n7398 , n4210 , n1473 );
    or g10842 ( n1497 , n7146 , n8030 );
    or g10843 ( n6475 , n6244 , n9043 );
    not g10844 ( n12747 , n11518 );
    xnor g10845 ( n12103 , n4393 , n4073 );
    xnor g10846 ( n3402 , n2360 , n9128 );
    nor g10847 ( n8575 , n5494 , n9578 );
    or g10848 ( n11672 , n3969 , n10945 );
    or g10849 ( n2503 , n6566 , n155 );
    xnor g10850 ( n11961 , n2887 , n8244 );
    not g10851 ( n5359 , n5030 );
    xnor g10852 ( n11012 , n3549 , n11151 );
    nor g10853 ( n9385 , n3152 , n4815 );
    xnor g10854 ( n397 , n3401 , n1555 );
    not g10855 ( n7415 , n1157 );
    nor g10856 ( n9306 , n5292 , n8213 );
    or g10857 ( n9180 , n6740 , n4837 );
    not g10858 ( n5540 , n9777 );
    xnor g10859 ( n3242 , n1277 , n11627 );
    or g10860 ( n3032 , n2449 , n12388 );
    xnor g10861 ( n2511 , n3223 , n1518 );
    not g10862 ( n10109 , n13220 );
    or g10863 ( n4588 , n5466 , n11025 );
    or g10864 ( n5109 , n6118 , n5384 );
    or g10865 ( n9660 , n13128 , n10858 );
    nor g10866 ( n11720 , n3414 , n5708 );
    and g10867 ( n9981 , n6602 , n9255 );
    nor g10868 ( n6233 , n4579 , n4763 );
    or g10869 ( n12825 , n5854 , n13172 );
    not g10870 ( n11300 , n10770 );
    nor g10871 ( n5473 , n7289 , n9285 );
    or g10872 ( n9987 , n1208 , n7264 );
    and g10873 ( n9717 , n5341 , n9108 );
    or g10874 ( n3706 , n8696 , n12351 );
    xnor g10875 ( n3401 , n12090 , n5534 );
    xnor g10876 ( n4435 , n10469 , n4404 );
    xnor g10877 ( n8870 , n1753 , n1915 );
    xor g10878 ( n5480 , n11582 , n751 );
    or g10879 ( n3609 , n10533 , n12919 );
    and g10880 ( n10655 , n2506 , n5093 );
    not g10881 ( n740 , n3511 );
    or g10882 ( n11859 , n3208 , n8268 );
    or g10883 ( n1972 , n7188 , n5797 );
    xnor g10884 ( n4437 , n1003 , n4733 );
    not g10885 ( n2541 , n10343 );
    or g10886 ( n6540 , n6733 , n8702 );
    and g10887 ( n10012 , n2168 , n1445 );
    or g10888 ( n12051 , n10604 , n1516 );
    and g10889 ( n1209 , n10670 , n5172 );
    xnor g10890 ( n7118 , n13136 , n702 );
    and g10891 ( n7979 , n8940 , n8233 );
    or g10892 ( n10152 , n1188 , n8348 );
    xnor g10893 ( n7294 , n4052 , n6616 );
    not g10894 ( n3639 , n9820 );
    not g10895 ( n10727 , n10024 );
    nor g10896 ( n1730 , n12946 , n2508 );
    and g10897 ( n3464 , n2272 , n4704 );
    xnor g10898 ( n2366 , n6476 , n555 );
    and g10899 ( n890 , n3456 , n5355 );
    xnor g10900 ( n6641 , n7094 , n1086 );
    or g10901 ( n4755 , n9557 , n2958 );
    xnor g10902 ( n10766 , n948 , n9211 );
    xnor g10903 ( n6683 , n2697 , n12160 );
    or g10904 ( n10631 , n10001 , n5209 );
    xnor g10905 ( n11076 , n9193 , n2797 );
    nor g10906 ( n700 , n13188 , n1288 );
    and g10907 ( n2169 , n11165 , n3201 );
    and g10908 ( n3067 , n13151 , n2598 );
    or g10909 ( n11872 , n80 , n542 );
    and g10910 ( n7830 , n10170 , n12221 );
    xnor g10911 ( n366 , n141 , n607 );
    and g10912 ( n7753 , n2702 , n5057 );
    nor g10913 ( n8057 , n2774 , n67 );
    or g10914 ( n629 , n6126 , n2627 );
    nor g10915 ( n11011 , n9664 , n6047 );
    nor g10916 ( n3803 , n1048 , n9106 );
    and g10917 ( n10750 , n7510 , n3812 );
    xnor g10918 ( n10983 , n3267 , n33 );
    not g10919 ( n1349 , n3682 );
    or g10920 ( n1984 , n4385 , n7930 );
    or g10921 ( n7570 , n7355 , n9259 );
    xnor g10922 ( n11401 , n9829 , n423 );
    or g10923 ( n7078 , n973 , n2281 );
    or g10924 ( n6436 , n11122 , n8268 );
    or g10925 ( n2696 , n946 , n479 );
    or g10926 ( n11414 , n1422 , n2059 );
    nor g10927 ( n214 , n32 , n4020 );
    and g10928 ( n12574 , n12211 , n3775 );
    not g10929 ( n1957 , n744 );
    xnor g10930 ( n11907 , n12650 , n11996 );
    or g10931 ( n3910 , n1638 , n12188 );
    or g10932 ( n1495 , n10057 , n4947 );
    xnor g10933 ( n2892 , n8310 , n3081 );
    xnor g10934 ( n5300 , n11597 , n1483 );
    xnor g10935 ( n3346 , n5590 , n12935 );
    xnor g10936 ( n1275 , n8144 , n1666 );
    or g10937 ( n12167 , n12203 , n3949 );
    and g10938 ( n2995 , n5177 , n8098 );
    not g10939 ( n7903 , n9620 );
    nor g10940 ( n8929 , n4331 , n1151 );
    not g10941 ( n5348 , n9241 );
    xnor g10942 ( n2172 , n12233 , n8105 );
    and g10943 ( n9953 , n8580 , n6242 );
    or g10944 ( n10835 , n11446 , n3949 );
    and g10945 ( n7579 , n6728 , n2027 );
    and g10946 ( n130 , n7433 , n9107 );
    xnor g10947 ( n4123 , n3113 , n1250 );
    not g10948 ( n3445 , n9362 );
    xnor g10949 ( n3680 , n4388 , n11246 );
    and g10950 ( n13079 , n8517 , n11187 );
    xnor g10951 ( n1518 , n9524 , n2947 );
    or g10952 ( n2520 , n6865 , n5792 );
    or g10953 ( n6591 , n6686 , n6786 );
    xnor g10954 ( n13114 , n6679 , n9573 );
    xnor g10955 ( n3763 , n3016 , n4501 );
    or g10956 ( n11517 , n12916 , n657 );
    or g10957 ( n3160 , n11979 , n9360 );
    xnor g10958 ( n4861 , n7924 , n7994 );
    and g10959 ( n5324 , n958 , n11681 );
    and g10960 ( n8036 , n10903 , n5215 );
    and g10961 ( n10273 , n10276 , n12183 );
    buf g10962 ( n479 , n917 );
    not g10963 ( n4536 , n8183 );
    nor g10964 ( n8656 , n12947 , n9568 );
    not g10965 ( n1070 , n9297 );
    buf g10966 ( n11144 , n6274 );
    and g10967 ( n10418 , n11308 , n9321 );
    xnor g10968 ( n6124 , n1892 , n4297 );
    xnor g10969 ( n8603 , n989 , n11575 );
    nor g10970 ( n9886 , n11844 , n9076 );
    xnor g10971 ( n12942 , n6686 , n2760 );
    or g10972 ( n7867 , n8890 , n5955 );
    and g10973 ( n10686 , n10802 , n2785 );
    or g10974 ( n6772 , n11310 , n6827 );
    and g10975 ( n3129 , n5945 , n2950 );
    and g10976 ( n3977 , n7847 , n5170 );
    not g10977 ( n2213 , n6532 );
    xnor g10978 ( n8742 , n4563 , n1228 );
    xnor g10979 ( n11349 , n4432 , n6119 );
    xnor g10980 ( n12962 , n9095 , n11103 );
    xnor g10981 ( n10118 , n7633 , n77 );
    xnor g10982 ( n1203 , n2495 , n9246 );
    or g10983 ( n7940 , n6854 , n8754 );
    or g10984 ( n152 , n12882 , n8268 );
    and g10985 ( n1899 , n2912 , n672 );
    or g10986 ( n5944 , n8499 , n1144 );
    xnor g10987 ( n5477 , n6337 , n10881 );
    or g10988 ( n11451 , n10293 , n2038 );
    and g10989 ( n2181 , n3622 , n7230 );
    and g10990 ( n3664 , n2176 , n881 );
    and g10991 ( n10186 , n1437 , n10200 );
    and g10992 ( n11133 , n9145 , n6036 );
    nor g10993 ( n12891 , n1227 , n4024 );
    xnor g10994 ( n3403 , n4821 , n4268 );
    not g10995 ( n4237 , n11324 );
    not g10996 ( n6841 , n8139 );
    xnor g10997 ( n3495 , n4735 , n2972 );
    and g10998 ( n6285 , n5803 , n3193 );
    and g10999 ( n2058 , n10117 , n10005 );
    xnor g11000 ( n2043 , n3135 , n4989 );
    or g11001 ( n7991 , n3727 , n118 );
    xnor g11002 ( n8745 , n5776 , n9457 );
    not g11003 ( n3419 , n9134 );
    or g11004 ( n7018 , n10977 , n5797 );
    and g11005 ( n9960 , n10861 , n5071 );
    or g11006 ( n2818 , n13082 , n8534 );
    not g11007 ( n4566 , n11774 );
    or g11008 ( n5385 , n9917 , n2943 );
    or g11009 ( n2243 , n436 , n9453 );
    or g11010 ( n9671 , n9335 , n8524 );
    nor g11011 ( n3912 , n1411 , n476 );
    nor g11012 ( n2784 , n954 , n1996 );
    nor g11013 ( n5906 , n630 , n12753 );
    or g11014 ( n2124 , n7230 , n3622 );
    or g11015 ( n8885 , n4143 , n9195 );
    not g11016 ( n9043 , n2820 );
    not g11017 ( n1783 , n12284 );
    nor g11018 ( n7140 , n2094 , n738 );
    and g11019 ( n11325 , n7315 , n238 );
    or g11020 ( n4099 , n3401 , n9233 );
    xnor g11021 ( n2690 , n2676 , n6868 );
    and g11022 ( n3488 , n8405 , n936 );
    xnor g11023 ( n12453 , n2365 , n9007 );
    or g11024 ( n34 , n7842 , n176 );
    or g11025 ( n2988 , n1327 , n9375 );
    not g11026 ( n2880 , n2762 );
    nor g11027 ( n5283 , n3382 , n10640 );
    and g11028 ( n9012 , n5901 , n12119 );
    and g11029 ( n8467 , n9382 , n10361 );
    or g11030 ( n4985 , n5565 , n9195 );
    xnor g11031 ( n10185 , n13104 , n8566 );
    xnor g11032 ( n9194 , n2409 , n6358 );
    and g11033 ( n5997 , n2158 , n11271 );
    or g11034 ( n9750 , n7700 , n1570 );
    not g11035 ( n12940 , n9981 );
    and g11036 ( n2333 , n6942 , n13240 );
    and g11037 ( n11432 , n6501 , n272 );
    or g11038 ( n6742 , n7277 , n5378 );
    or g11039 ( n5661 , n12709 , n431 );
    and g11040 ( n2989 , n4652 , n9700 );
    xnor g11041 ( n8709 , n1230 , n9699 );
    nor g11042 ( n2140 , n9585 , n3766 );
    xnor g11043 ( n2247 , n6850 , n8553 );
    xnor g11044 ( n5866 , n12591 , n10047 );
    xnor g11045 ( n8588 , n3423 , n2357 );
    xnor g11046 ( n6642 , n136 , n9744 );
    and g11047 ( n339 , n7699 , n8703 );
    or g11048 ( n11787 , n10077 , n4994 );
    or g11049 ( n10928 , n6575 , n9504 );
    and g11050 ( n4899 , n2091 , n3597 );
    xnor g11051 ( n9261 , n4752 , n10561 );
    not g11052 ( n8904 , n12853 );
    and g11053 ( n6425 , n5161 , n9119 );
    nor g11054 ( n13153 , n11504 , n10262 );
    not g11055 ( n640 , n405 );
    not g11056 ( n5229 , n4315 );
    or g11057 ( n6571 , n11149 , n8352 );
    or g11058 ( n6522 , n10352 , n11107 );
    and g11059 ( n2285 , n1047 , n963 );
    and g11060 ( n9738 , n11829 , n6940 );
    not g11061 ( n5434 , n7726 );
    or g11062 ( n3051 , n45 , n8563 );
    buf g11063 ( n2958 , n12954 );
    or g11064 ( n6722 , n4564 , n6370 );
    and g11065 ( n1160 , n7044 , n12368 );
    not g11066 ( n6983 , n9885 );
    not g11067 ( n10380 , n465 );
    xnor g11068 ( n11776 , n9205 , n5425 );
    not g11069 ( n12092 , n12715 );
    or g11070 ( n5440 , n899 , n11107 );
    and g11071 ( n665 , n8252 , n3120 );
    xnor g11072 ( n11691 , n6927 , n3107 );
    xnor g11073 ( n5689 , n4912 , n7773 );
    and g11074 ( n8538 , n5961 , n4244 );
    not g11075 ( n9795 , n12269 );
    and g11076 ( n8838 , n8460 , n2291 );
    or g11077 ( n10480 , n5351 , n12659 );
    not g11078 ( n9489 , n8468 );
    or g11079 ( n4418 , n9450 , n1570 );
    not g11080 ( n3412 , n11248 );
    and g11081 ( n11200 , n695 , n7483 );
    and g11082 ( n9898 , n1246 , n10597 );
    or g11083 ( n3501 , n12795 , n8702 );
    xnor g11084 ( n7992 , n9207 , n12207 );
    and g11085 ( n2277 , n500 , n13241 );
    xor g11086 ( n6209 , n1972 , n10015 );
    xnor g11087 ( n1262 , n4805 , n909 );
    not g11088 ( n4487 , n9904 );
    xnor g11089 ( n12961 , n10511 , n706 );
    nor g11090 ( n779 , n8731 , n3175 );
    nor g11091 ( n7198 , n6717 , n9812 );
    and g11092 ( n10036 , n489 , n12206 );
    nor g11093 ( n3440 , n3309 , n4513 );
    and g11094 ( n6996 , n2292 , n2362 );
    or g11095 ( n5085 , n7774 , n11355 );
    not g11096 ( n4495 , n6168 );
    nor g11097 ( n5831 , n4924 , n4919 );
    or g11098 ( n7665 , n3978 , n8270 );
    not g11099 ( n5611 , n7659 );
    and g11100 ( n4518 , n8228 , n6085 );
    or g11101 ( n1065 , n1152 , n1463 );
    xnor g11102 ( n8814 , n12608 , n7310 );
    and g11103 ( n8986 , n5159 , n10496 );
    xnor g11104 ( n8549 , n1107 , n9541 );
    or g11105 ( n12044 , n12741 , n13086 );
    and g11106 ( n7701 , n12754 , n11714 );
    nor g11107 ( n5652 , n7728 , n9804 );
    not g11108 ( n189 , n103 );
    or g11109 ( n3583 , n1017 , n8281 );
    and g11110 ( n543 , n9348 , n4271 );
    not g11111 ( n3894 , n7436 );
    xnor g11112 ( n2709 , n6987 , n6646 );
    and g11113 ( n7440 , n2090 , n3834 );
    not g11114 ( n7620 , n4748 );
    xnor g11115 ( n4569 , n3417 , n12432 );
    xnor g11116 ( n4264 , n7023 , n11497 );
    and g11117 ( n9147 , n4358 , n6268 );
    or g11118 ( n12633 , n9385 , n670 );
    not g11119 ( n6960 , n6535 );
    or g11120 ( n12132 , n5666 , n2133 );
    or g11121 ( n8982 , n10208 , n8683 );
    or g11122 ( n8296 , n3111 , n11169 );
    or g11123 ( n3851 , n9411 , n7440 );
    or g11124 ( n5592 , n8028 , n2746 );
    or g11125 ( n8133 , n2183 , n12695 );
    not g11126 ( n560 , n353 );
    or g11127 ( n1681 , n136 , n5816 );
    xnor g11128 ( n3305 , n6203 , n763 );
    or g11129 ( n11104 , n4948 , n11362 );
    xnor g11130 ( n5691 , n1034 , n12925 );
    or g11131 ( n12382 , n2090 , n3834 );
    not g11132 ( n12623 , n9620 );
    or g11133 ( n7453 , n1508 , n5454 );
    or g11134 ( n6111 , n115 , n479 );
    xnor g11135 ( n3787 , n6213 , n7144 );
    or g11136 ( n2066 , n11519 , n5242 );
    or g11137 ( n6947 , n700 , n6284 );
    nor g11138 ( n5622 , n3188 , n4002 );
    nor g11139 ( n11573 , n9500 , n1492 );
    nor g11140 ( n4018 , n11715 , n5289 );
    and g11141 ( n1961 , n5983 , n5370 );
    and g11142 ( n6864 , n4714 , n3690 );
    nor g11143 ( n5792 , n8357 , n8134 );
    and g11144 ( n10202 , n7892 , n11599 );
    xnor g11145 ( n5272 , n6453 , n11647 );
    xnor g11146 ( n7513 , n3868 , n8564 );
    nor g11147 ( n4868 , n11230 , n799 );
    or g11148 ( n122 , n5423 , n8348 );
    buf g11149 ( n2059 , n11148 );
    xnor g11150 ( n5101 , n547 , n8676 );
    or g11151 ( n8167 , n7299 , n4082 );
    and g11152 ( n10407 , n6374 , n3933 );
    xnor g11153 ( n1992 , n6014 , n5754 );
    not g11154 ( n6889 , n828 );
    and g11155 ( n3106 , n10113 , n2252 );
    and g11156 ( n2705 , n12215 , n10220 );
    xnor g11157 ( n12035 , n5027 , n9446 );
    xnor g11158 ( n11327 , n8550 , n1114 );
    and g11159 ( n1013 , n8386 , n615 );
    and g11160 ( n7400 , n1538 , n641 );
    or g11161 ( n2518 , n13117 , n2387 );
    and g11162 ( n8278 , n7461 , n8148 );
    not g11163 ( n9596 , n13138 );
    and g11164 ( n13037 , n13216 , n6502 );
    and g11165 ( n7491 , n9978 , n4322 );
    xnor g11166 ( n10393 , n3845 , n1215 );
    xnor g11167 ( n10799 , n549 , n4441 );
    and g11168 ( n2798 , n4744 , n10244 );
    and g11169 ( n2304 , n13047 , n8394 );
    and g11170 ( n2679 , n1319 , n3984 );
    and g11171 ( n3642 , n4440 , n8846 );
    not g11172 ( n6590 , n4470 );
    or g11173 ( n1504 , n871 , n8514 );
    xnor g11174 ( n7066 , n11725 , n3052 );
    or g11175 ( n11915 , n12617 , n8702 );
    and g11176 ( n2965 , n6918 , n4061 );
    not g11177 ( n8002 , n2310 );
    xnor g11178 ( n3873 , n9601 , n8934 );
    or g11179 ( n7414 , n10402 , n3981 );
    or g11180 ( n8952 , n4827 , n2240 );
    xor g11181 ( n5808 , n11990 , n8558 );
    xnor g11182 ( n9197 , n9084 , n12744 );
    not g11183 ( n10010 , n11266 );
    xnor g11184 ( n3771 , n4867 , n10995 );
    nor g11185 ( n11730 , n12022 , n10316 );
    not g11186 ( n1976 , n1190 );
    and g11187 ( n3416 , n618 , n9858 );
    or g11188 ( n8946 , n9696 , n11011 );
    not g11189 ( n4657 , n8332 );
    or g11190 ( n8447 , n13137 , n5130 );
    or g11191 ( n11125 , n11242 , n5797 );
    and g11192 ( n4315 , n6320 , n127 );
    or g11193 ( n8488 , n75 , n7530 );
    and g11194 ( n10458 , n12921 , n9600 );
    nor g11195 ( n9243 , n7126 , n2227 );
    xnor g11196 ( n2903 , n8461 , n6007 );
    not g11197 ( n2055 , n10463 );
    not g11198 ( n11612 , n817 );
    or g11199 ( n12472 , n1194 , n2675 );
    not g11200 ( n12258 , n295 );
    not g11201 ( n320 , n8432 );
    xnor g11202 ( n941 , n2230 , n11726 );
    xnor g11203 ( n4000 , n8931 , n10416 );
    not g11204 ( n10892 , n1313 );
    not g11205 ( n11232 , n10442 );
    or g11206 ( n12897 , n12023 , n2449 );
    and g11207 ( n12237 , n7963 , n3334 );
    and g11208 ( n13209 , n8443 , n132 );
    xnor g11209 ( n10209 , n1491 , n1109 );
    xnor g11210 ( n3593 , n257 , n4190 );
    and g11211 ( n4469 , n910 , n178 );
    or g11212 ( n3657 , n11212 , n206 );
    not g11213 ( n4642 , n11666 );
    xnor g11214 ( n251 , n3249 , n10403 );
    nor g11215 ( n10257 , n13018 , n355 );
    or g11216 ( n4893 , n11514 , n11244 );
    xnor g11217 ( n12460 , n2076 , n8390 );
    or g11218 ( n1442 , n6922 , n4724 );
    or g11219 ( n6226 , n12997 , n5797 );
    and g11220 ( n13145 , n9008 , n3118 );
    not g11221 ( n4488 , n10821 );
    not g11222 ( n7839 , n4033 );
    nor g11223 ( n4416 , n8605 , n112 );
    or g11224 ( n11722 , n5806 , n3981 );
    or g11225 ( n203 , n6337 , n10881 );
    xnor g11226 ( n2369 , n11671 , n9062 );
    nor g11227 ( n1804 , n1134 , n3283 );
    nor g11228 ( n7800 , n11304 , n4463 );
    nor g11229 ( n4200 , n9494 , n2996 );
    or g11230 ( n1846 , n3530 , n5676 );
    not g11231 ( n755 , n8820 );
    not g11232 ( n2773 , n1756 );
    nor g11233 ( n9056 , n4641 , n6817 );
    xnor g11234 ( n4986 , n5504 , n5732 );
    and g11235 ( n1192 , n12027 , n11502 );
    not g11236 ( n10287 , n4075 );
    or g11237 ( n12613 , n1224 , n7781 );
    not g11238 ( n5921 , n925 );
    nor g11239 ( n7626 , n7806 , n11290 );
    xnor g11240 ( n10357 , n9293 , n6400 );
    xnor g11241 ( n13048 , n12293 , n2907 );
    or g11242 ( n9517 , n12599 , n941 );
    and g11243 ( n12566 , n6073 , n4544 );
    xnor g11244 ( n31 , n1789 , n2908 );
    xnor g11245 ( n8536 , n8205 , n11834 );
    nor g11246 ( n10486 , n4328 , n12320 );
    xnor g11247 ( n1205 , n7156 , n4843 );
    and g11248 ( n4300 , n3820 , n4308 );
    not g11249 ( n7837 , n2771 );
    or g11250 ( n4750 , n11612 , n7935 );
    and g11251 ( n6827 , n5301 , n422 );
    or g11252 ( n11258 , n11431 , n4435 );
    or g11253 ( n2134 , n383 , n11899 );
    and g11254 ( n1075 , n767 , n2498 );
    xnor g11255 ( n3042 , n1917 , n9777 );
    and g11256 ( n12358 , n2722 , n2146 );
    xnor g11257 ( n1277 , n8799 , n1665 );
    or g11258 ( n13126 , n11226 , n4640 );
    and g11259 ( n11549 , n11450 , n4757 );
    xnor g11260 ( n7993 , n7876 , n3692 );
    not g11261 ( n12378 , n5161 );
    not g11262 ( n7312 , n12538 );
    and g11263 ( n4516 , n10560 , n1636 );
    xnor g11264 ( n9024 , n6867 , n2454 );
    and g11265 ( n2391 , n8527 , n2143 );
    xnor g11266 ( n3458 , n11159 , n3952 );
    nor g11267 ( n11883 , n11702 , n11710 );
    not g11268 ( n9761 , n834 );
    and g11269 ( n12873 , n10876 , n3645 );
    or g11270 ( n495 , n2701 , n10029 );
    and g11271 ( n5275 , n6723 , n2327 );
    and g11272 ( n4981 , n10047 , n12591 );
    and g11273 ( n3168 , n13201 , n3815 );
    or g11274 ( n2854 , n10814 , n11668 );
    xnor g11275 ( n12277 , n12765 , n11346 );
    xnor g11276 ( n7373 , n437 , n10028 );
    and g11277 ( n952 , n6676 , n9869 );
    nor g11278 ( n10693 , n11798 , n551 );
    xnor g11279 ( n11013 , n1531 , n2001 );
    or g11280 ( n1582 , n9490 , n9618 );
    and g11281 ( n10390 , n12095 , n6464 );
    not g11282 ( n10016 , n10642 );
    not g11283 ( n5683 , n6085 );
    not g11284 ( n1216 , n4957 );
    and g11285 ( n5034 , n9762 , n3038 );
    or g11286 ( n12590 , n8414 , n4124 );
    and g11287 ( n11854 , n7715 , n9669 );
    not g11288 ( n5382 , n7419 );
    xnor g11289 ( n4338 , n12559 , n6026 );
    not g11290 ( n8161 , n1356 );
    nor g11291 ( n10784 , n7025 , n6994 );
    not g11292 ( n13012 , n5715 );
    or g11293 ( n4199 , n715 , n4936 );
    xnor g11294 ( n8442 , n6754 , n4009 );
    xnor g11295 ( n10789 , n122 , n10303 );
    not g11296 ( n4464 , n4330 );
    not g11297 ( n488 , n6085 );
    and g11298 ( n7054 , n11600 , n2610 );
    xnor g11299 ( n9902 , n12541 , n3680 );
    xnor g11300 ( n6032 , n11139 , n10393 );
    and g11301 ( n10452 , n8461 , n6388 );
    xnor g11302 ( n2847 , n8567 , n12176 );
    or g11303 ( n8911 , n6967 , n11871 );
    not g11304 ( n5467 , n3627 );
    xnor g11305 ( n12872 , n2888 , n11066 );
    xnor g11306 ( n11788 , n10807 , n12656 );
    xnor g11307 ( n11447 , n6669 , n11872 );
    xnor g11308 ( n9896 , n11270 , n6899 );
    and g11309 ( n72 , n7949 , n3215 );
    not g11310 ( n7526 , n7728 );
    xnor g11311 ( n4163 , n9306 , n6430 );
    nor g11312 ( n12653 , n6930 , n377 );
    nor g11313 ( n6342 , n1753 , n1915 );
    and g11314 ( n749 , n8500 , n3860 );
    and g11315 ( n9192 , n7681 , n9066 );
    xnor g11316 ( n9218 , n1173 , n8347 );
    xnor g11317 ( n10058 , n4308 , n3820 );
    or g11318 ( n3721 , n2048 , n121 );
    xnor g11319 ( n8067 , n5096 , n9536 );
    or g11320 ( n9938 , n10730 , n5076 );
    or g11321 ( n4241 , n392 , n6041 );
    or g11322 ( n9729 , n8131 , n4640 );
    xnor g11323 ( n975 , n13069 , n1130 );
    nor g11324 ( n9498 , n2102 , n4838 );
    and g11325 ( n11052 , n4588 , n1914 );
    xnor g11326 ( n8035 , n4316 , n3573 );
    xnor g11327 ( n11182 , n2949 , n10789 );
    nor g11328 ( n3811 , n3664 , n6408 );
    or g11329 ( n8887 , n813 , n10871 );
    xnor g11330 ( n10139 , n8998 , n4076 );
    or g11331 ( n10313 , n10439 , n1026 );
    nor g11332 ( n2065 , n11730 , n6443 );
    not g11333 ( n5565 , n2252 );
    and g11334 ( n10268 , n7529 , n2252 );
    or g11335 ( n3543 , n6630 , n4230 );
    nor g11336 ( n6885 , n10925 , n4256 );
    and g11337 ( n13213 , n563 , n9677 );
    or g11338 ( n1828 , n9421 , n8490 );
    nor g11339 ( n7989 , n2087 , n10557 );
    and g11340 ( n4751 , n5934 , n4461 );
    xnor g11341 ( n1142 , n7231 , n12519 );
    xnor g11342 ( n3153 , n5139 , n5518 );
    nor g11343 ( n5028 , n8626 , n2841 );
    xor g11344 ( n2072 , n912 , n3831 );
    xnor g11345 ( n11724 , n1172 , n6681 );
    or g11346 ( n1077 , n12069 , n9761 );
    xnor g11347 ( n10925 , n12539 , n10702 );
    not g11348 ( n9711 , n9528 );
    or g11349 ( n5869 , n3586 , n1771 );
    or g11350 ( n11647 , n1012 , n956 );
    xnor g11351 ( n923 , n2013 , n205 );
    xnor g11352 ( n11903 , n12134 , n7574 );
    not g11353 ( n10991 , n772 );
    not g11354 ( n9921 , n7572 );
    xnor g11355 ( n7782 , n11499 , n6784 );
    nor g11356 ( n2187 , n8717 , n3869 );
    xnor g11357 ( n6411 , n7483 , n4332 );
    or g11358 ( n3367 , n2226 , n9622 );
    and g11359 ( n2273 , n3311 , n411 );
    not g11360 ( n2130 , n12567 );
    not g11361 ( n1238 , n5768 );
    xnor g11362 ( n5049 , n9842 , n12803 );
    xnor g11363 ( n8527 , n11015 , n2121 );
    and g11364 ( n1698 , n2482 , n2758 );
    not g11365 ( n2671 , n3130 );
    xnor g11366 ( n7654 , n901 , n4775 );
    and g11367 ( n9481 , n2777 , n8860 );
    xor g11368 ( n726 , n12475 , n5488 );
    or g11369 ( n6866 , n10733 , n10331 );
    xor g11370 ( n7085 , n11553 , n11641 );
    not g11371 ( n1215 , n6445 );
    and g11372 ( n3837 , n1579 , n11307 );
    or g11373 ( n5851 , n3784 , n9075 );
    not g11374 ( n11045 , n600 );
    xnor g11375 ( n4953 , n10660 , n7351 );
    or g11376 ( n9094 , n7620 , n1985 );
    or g11377 ( n1968 , n5733 , n5242 );
    xnor g11378 ( n8589 , n11541 , n3742 );
    xnor g11379 ( n1114 , n13119 , n5499 );
    or g11380 ( n8548 , n4610 , n5169 );
    xnor g11381 ( n6361 , n12857 , n7804 );
    not g11382 ( n8335 , n5969 );
    and g11383 ( n6507 , n490 , n6389 );
    or g11384 ( n6382 , n11284 , n12273 );
    xnor g11385 ( n11510 , n7359 , n3199 );
    xnor g11386 ( n4800 , n5120 , n8821 );
    xnor g11387 ( n3790 , n10897 , n4996 );
    and g11388 ( n13125 , n3284 , n6813 );
    xnor g11389 ( n3021 , n385 , n3523 );
    or g11390 ( n10768 , n4001 , n12177 );
    and g11391 ( n9929 , n4818 , n1602 );
    or g11392 ( n12992 , n10638 , n8983 );
    nor g11393 ( n10349 , n10578 , n5282 );
    not g11394 ( n2163 , n11179 );
    and g11395 ( n8179 , n870 , n11655 );
    xnor g11396 ( n3868 , n7382 , n10461 );
    xnor g11397 ( n359 , n8967 , n12163 );
    or g11398 ( n1259 , n3090 , n990 );
    and g11399 ( n2351 , n1715 , n8313 );
    xnor g11400 ( n6165 , n4645 , n2447 );
    xnor g11401 ( n5629 , n8158 , n12360 );
    or g11402 ( n869 , n5902 , n11606 );
    not g11403 ( n9592 , n7085 );
    and g11404 ( n9233 , n10289 , n4755 );
    xnor g11405 ( n8690 , n13121 , n11348 );
    not g11406 ( n987 , n12065 );
    or g11407 ( n11229 , n11751 , n1820 );
    or g11408 ( n1499 , n10962 , n10473 );
    not g11409 ( n513 , n229 );
    or g11410 ( n4727 , n1101 , n10871 );
    xnor g11411 ( n8612 , n690 , n6893 );
    nor g11412 ( n4952 , n5071 , n10861 );
    not g11413 ( n2718 , n9620 );
    or g11414 ( n7971 , n9515 , n2569 );
    not g11415 ( n10654 , n3095 );
    not g11416 ( n3157 , n103 );
    not g11417 ( n5673 , n7153 );
    xor g11418 ( n4824 , n5965 , n485 );
    or g11419 ( n570 , n7925 , n8563 );
    and g11420 ( n1395 , n10479 , n11434 );
    xnor g11421 ( n7815 , n9989 , n12692 );
    nor g11422 ( n2450 , n9235 , n9506 );
    xnor g11423 ( n4713 , n9150 , n2397 );
    or g11424 ( n9482 , n11845 , n4658 );
    xnor g11425 ( n13193 , n11361 , n13016 );
    or g11426 ( n12765 , n10085 , n1570 );
    and g11427 ( n10595 , n8717 , n3869 );
    not g11428 ( n2893 , n8230 );
    and g11429 ( n6789 , n6066 , n3706 );
    xnor g11430 ( n1385 , n10446 , n10939 );
    and g11431 ( n3145 , n7443 , n12442 );
    xnor g11432 ( n9028 , n10046 , n5259 );
    or g11433 ( n2079 , n7872 , n8744 );
    or g11434 ( n4737 , n3348 , n11748 );
    nor g11435 ( n1995 , n2440 , n13163 );
    or g11436 ( n3842 , n3733 , n11426 );
    not g11437 ( n8005 , n2590 );
    xnor g11438 ( n7166 , n9861 , n1207 );
    or g11439 ( n5846 , n1168 , n8348 );
    and g11440 ( n7276 , n1757 , n4330 );
    xnor g11441 ( n11211 , n2261 , n7061 );
    or g11442 ( n7901 , n1633 , n5524 );
    xnor g11443 ( n10911 , n12754 , n7451 );
    nor g11444 ( n10454 , n705 , n9208 );
    xnor g11445 ( n11072 , n2730 , n11440 );
    not g11446 ( n12471 , n767 );
    not g11447 ( n9679 , n5320 );
    not g11448 ( n10411 , n1982 );
    not g11449 ( n6164 , n8917 );
    not g11450 ( n1346 , n6836 );
    or g11451 ( n2795 , n6054 , n5290 );
    or g11452 ( n12185 , n8670 , n2707 );
    xnor g11453 ( n388 , n6195 , n12886 );
    not g11454 ( n11270 , n691 );
    and g11455 ( n11569 , n8642 , n8488 );
    xnor g11456 ( n7664 , n7671 , n8078 );
    nor g11457 ( n9916 , n8718 , n11531 );
    xnor g11458 ( n10846 , n7593 , n10701 );
    and g11459 ( n8543 , n104 , n6911 );
    nor g11460 ( n11833 , n7500 , n3681 );
    or g11461 ( n9150 , n4166 , n6404 );
    and g11462 ( n9225 , n12361 , n10317 );
    xnor g11463 ( n2923 , n12217 , n7164 );
    or g11464 ( n6850 , n4966 , n9714 );
    xnor g11465 ( n10987 , n4750 , n11475 );
    xnor g11466 ( n9267 , n3309 , n11534 );
    and g11467 ( n4440 , n11665 , n8860 );
    and g11468 ( n4669 , n8736 , n7081 );
    not g11469 ( n8852 , n5214 );
    xnor g11470 ( n2293 , n6722 , n7416 );
    or g11471 ( n8909 , n9634 , n12029 );
    xnor g11472 ( n10816 , n10331 , n13226 );
    not g11473 ( n7068 , n9528 );
    and g11474 ( n2089 , n5268 , n7012 );
    nor g11475 ( n9275 , n7715 , n2458 );
    and g11476 ( n1710 , n5442 , n181 );
    xnor g11477 ( n10785 , n10804 , n1573 );
    or g11478 ( n3288 , n11320 , n10871 );
    not g11479 ( n1920 , n6064 );
    or g11480 ( n2781 , n12565 , n5067 );
    xnor g11481 ( n13029 , n6780 , n2111 );
    nor g11482 ( n11602 , n2058 , n6907 );
    xnor g11483 ( n4059 , n2731 , n5880 );
    or g11484 ( n3191 , n2449 , n1570 );
    or g11485 ( n4461 , n4348 , n7813 );
    or g11486 ( n8009 , n3025 , n4510 );
    and g11487 ( n4733 , n5129 , n9180 );
    xnor g11488 ( n9206 , n7118 , n12480 );
    xor g11489 ( n6861 , n10544 , n1064 );
    not g11490 ( n12667 , n6950 );
    xnor g11491 ( n4832 , n2821 , n5343 );
    not g11492 ( n7980 , n6277 );
    nor g11493 ( n1877 , n4205 , n1351 );
    or g11494 ( n6871 , n12522 , n5775 );
    buf g11495 ( n3981 , n789 );
    not g11496 ( n2824 , n5833 );
    or g11497 ( n9451 , n2384 , n3396 );
    and g11498 ( n11085 , n7797 , n5996 );
    or g11499 ( n3818 , n6086 , n12188 );
    xnor g11500 ( n800 , n8587 , n4707 );
    not g11501 ( n2768 , n4335 );
    xor g11502 ( n4739 , n5784 , n7722 );
    xnor g11503 ( n8137 , n2361 , n11897 );
    not g11504 ( n4890 , n3832 );
    and g11505 ( n12949 , n2583 , n10673 );
    and g11506 ( n1762 , n2472 , n11593 );
    and g11507 ( n7960 , n11665 , n9570 );
    xnor g11508 ( n7932 , n3739 , n325 );
    not g11509 ( n8778 , n3988 );
    not g11510 ( n9736 , n11474 );
    or g11511 ( n10469 , n4855 , n2958 );
    xnor g11512 ( n11355 , n52 , n11923 );
    xnor g11513 ( n2014 , n8411 , n807 );
    or g11514 ( n6981 , n7177 , n10551 );
    and g11515 ( n4587 , n6884 , n6424 );
    nor g11516 ( n6737 , n10047 , n12591 );
    buf g11517 ( n4724 , n3858 );
    not g11518 ( n2678 , n11734 );
    or g11519 ( n8239 , n2576 , n8262 );
    or g11520 ( n12833 , n13190 , n6265 );
    not g11521 ( n1480 , n11734 );
    not g11522 ( n10711 , n3715 );
    or g11523 ( n10771 , n2896 , n10311 );
    or g11524 ( n9361 , n7878 , n10552 );
    or g11525 ( n10650 , n4649 , n2059 );
    or g11526 ( n12716 , n11965 , n10764 );
    or g11527 ( n10624 , n5645 , n6732 );
    or g11528 ( n11867 , n12648 , n8561 );
    and g11529 ( n12231 , n417 , n7109 );
    or g11530 ( n13099 , n881 , n2176 );
    xnor g11531 ( n11083 , n11572 , n1584 );
    or g11532 ( n4322 , n12020 , n3210 );
    and g11533 ( n10658 , n12010 , n11451 );
    not g11534 ( n12315 , n2374 );
    xnor g11535 ( n12187 , n3862 , n571 );
    xnor g11536 ( n6434 , n824 , n1318 );
    xnor g11537 ( n13144 , n5874 , n10468 );
    nor g11538 ( n4752 , n3615 , n5507 );
    xnor g11539 ( n4721 , n9645 , n10056 );
    not g11540 ( n4778 , n382 );
    xnor g11541 ( n7924 , n4217 , n3029 );
    or g11542 ( n10561 , n1360 , n9511 );
    not g11543 ( n11340 , n11199 );
    or g11544 ( n2396 , n9593 , n8806 );
    not g11545 ( n1554 , n937 );
    not g11546 ( n5222 , n299 );
    or g11547 ( n11105 , n9341 , n2594 );
    xnor g11548 ( n6572 , n3802 , n2459 );
    or g11549 ( n12431 , n9339 , n9159 );
    xnor g11550 ( n710 , n4576 , n9773 );
    xnor g11551 ( n8323 , n8426 , n11754 );
    xnor g11552 ( n8515 , n9534 , n3268 );
    not g11553 ( n10459 , n9901 );
    or g11554 ( n8107 , n13205 , n4310 );
    and g11555 ( n3967 , n7470 , n3020 );
    not g11556 ( n4290 , n9531 );
    xnor g11557 ( n2548 , n6067 , n1076 );
    nor g11558 ( n8756 , n3305 , n5662 );
    not g11559 ( n845 , n7729 );
    or g11560 ( n723 , n3429 , n4030 );
    and g11561 ( n7785 , n3936 , n4810 );
    xnor g11562 ( n2382 , n9535 , n2852 );
    xnor g11563 ( n5796 , n9107 , n4520 );
    or g11564 ( n11408 , n10593 , n3063 );
    nor g11565 ( n12561 , n5309 , n1000 );
    xnor g11566 ( n1228 , n2128 , n8403 );
    not g11567 ( n2832 , n12422 );
    or g11568 ( n6039 , n9252 , n3464 );
    xnor g11569 ( n8027 , n10913 , n3746 );
    not g11570 ( n1789 , n3253 );
    or g11571 ( n8314 , n53 , n6769 );
    not g11572 ( n2825 , n5189 );
    or g11573 ( n11919 , n6043 , n327 );
    xnor g11574 ( n9951 , n10514 , n7293 );
    xnor g11575 ( n11413 , n1991 , n8603 );
    not g11576 ( n7362 , n13128 );
    and g11577 ( n12543 , n12992 , n9409 );
    or g11578 ( n9539 , n4665 , n1985 );
    or g11579 ( n5695 , n1511 , n11668 );
    not g11580 ( n10879 , n5031 );
    or g11581 ( n10092 , n7258 , n12234 );
    xnor g11582 ( n5617 , n9874 , n6397 );
    or g11583 ( n5491 , n10354 , n12763 );
    xnor g11584 ( n8584 , n487 , n9239 );
    or g11585 ( n6218 , n11318 , n8880 );
    and g11586 ( n9752 , n3583 , n13010 );
    or g11587 ( n2348 , n300 , n10619 );
    not g11588 ( n4744 , n1595 );
    and g11589 ( n5036 , n10346 , n2534 );
    and g11590 ( n11362 , n11415 , n7564 );
    or g11591 ( n5966 , n7984 , n11470 );
    not g11592 ( n2067 , n7137 );
    xnor g11593 ( n4802 , n11142 , n11762 );
    or g11594 ( n7419 , n10188 , n4947 );
    or g11595 ( n7887 , n5667 , n11144 );
    and g11596 ( n5676 , n3022 , n12807 );
    or g11597 ( n12344 , n12224 , n4979 );
    xnor g11598 ( n12011 , n12081 , n9936 );
    or g11599 ( n11633 , n1265 , n2552 );
    not g11600 ( n2673 , n1552 );
    or g11601 ( n9877 , n5079 , n1144 );
    and g11602 ( n9661 , n898 , n4154 );
    nor g11603 ( n11649 , n244 , n2436 );
    or g11604 ( n9313 , n4796 , n4947 );
    or g11605 ( n7751 , n2118 , n12273 );
    nor g11606 ( n12735 , n4508 , n7686 );
    and g11607 ( n10339 , n11339 , n1080 );
    xnor g11608 ( n9198 , n12061 , n753 );
    or g11609 ( n12375 , n8934 , n4423 );
    or g11610 ( n1351 , n3898 , n9223 );
    nor g11611 ( n10690 , n3254 , n3979 );
    and g11612 ( n1292 , n581 , n8957 );
    or g11613 ( n11742 , n12242 , n5087 );
    nor g11614 ( n5285 , n3138 , n11316 );
    and g11615 ( n3643 , n2451 , n2799 );
    not g11616 ( n11771 , n13219 );
    xnor g11617 ( n12928 , n10197 , n10615 );
    or g11618 ( n9520 , n278 , n11968 );
    or g11619 ( n11987 , n12748 , n10871 );
    xnor g11620 ( n6287 , n11229 , n7758 );
    or g11621 ( n13221 , n10761 , n13242 );
    nor g11622 ( n9269 , n9683 , n5849 );
    or g11623 ( n2034 , n97 , n4373 );
    xnor g11624 ( n12831 , n11653 , n13042 );
    and g11625 ( n5379 , n12129 , n10960 );
    nor g11626 ( n6494 , n3518 , n1069 );
    and g11627 ( n3860 , n11986 , n10376 );
    nor g11628 ( n4567 , n4568 , n3353 );
    xnor g11629 ( n4837 , n6861 , n1802 );
    and g11630 ( n6269 , n2590 , n8290 );
    not g11631 ( n9827 , n6317 );
    and g11632 ( n11898 , n11994 , n331 );
    xnor g11633 ( n1532 , n12584 , n3045 );
    xnor g11634 ( n4409 , n7788 , n8007 );
    and g11635 ( n6426 , n11819 , n8775 );
    or g11636 ( n6775 , n6710 , n5782 );
    and g11637 ( n11402 , n5568 , n4748 );
    or g11638 ( n10426 , n4235 , n3576 );
    not g11639 ( n5177 , n12557 );
    or g11640 ( n10891 , n9011 , n3559 );
    xnor g11641 ( n841 , n12796 , n8308 );
    and g11642 ( n8523 , n3944 , n3541 );
    not g11643 ( n10402 , n1636 );
    xnor g11644 ( n4772 , n7849 , n5543 );
    xnor g11645 ( n7558 , n8830 , n10181 );
    xnor g11646 ( n171 , n7806 , n11377 );
    xnor g11647 ( n9317 , n5744 , n7715 );
    xor g11648 ( n12172 , n13006 , n10268 );
    nor g11649 ( n6569 , n250 , n2492 );
    nor g11650 ( n7233 , n9543 , n2489 );
    xnor g11651 ( n5544 , n4559 , n5675 );
    nor g11652 ( n6817 , n4573 , n10838 );
    or g11653 ( n714 , n8324 , n2675 );
    or g11654 ( n4471 , n2405 , n8614 );
    xnor g11655 ( n4459 , n5197 , n6600 );
    xnor g11656 ( n5030 , n8657 , n9127 );
    nor g11657 ( n10166 , n7560 , n6600 );
    and g11658 ( n6239 , n1607 , n9780 );
    xnor g11659 ( n12345 , n4768 , n3943 );
    or g11660 ( n11660 , n6183 , n3977 );
    xnor g11661 ( n8804 , n3501 , n7607 );
    xnor g11662 ( n9214 , n536 , n4581 );
    not g11663 ( n6438 , n1165 );
    or g11664 ( n5381 , n6314 , n2354 );
    or g11665 ( n1125 , n10558 , n4724 );
    xor g11666 ( n9117 , n4211 , n10485 );
    or g11667 ( n5151 , n1101 , n2387 );
    not g11668 ( n11449 , n6392 );
    and g11669 ( n10652 , n1460 , n5506 );
    buf g11670 ( n12328 , n9280 );
    xnor g11671 ( n2368 , n11035 , n1439 );
    and g11672 ( n9920 , n100 , n9725 );
    or g11673 ( n3417 , n10128 , n11107 );
    or g11674 ( n11407 , n935 , n4230 );
    not g11675 ( n6314 , n7527 );
    not g11676 ( n8995 , n4788 );
    not g11677 ( n11707 , n2409 );
    xnor g11678 ( n9505 , n12769 , n2909 );
    or g11679 ( n8474 , n8912 , n2622 );
    and g11680 ( n10623 , n12915 , n4487 );
    and g11681 ( n4231 , n1024 , n4294 );
    not g11682 ( n6854 , n12482 );
    not g11683 ( n5787 , n7240 );
    xnor g11684 ( n12745 , n6816 , n7332 );
    xnor g11685 ( n10669 , n8317 , n12212 );
    xnor g11686 ( n10861 , n6353 , n7431 );
    xnor g11687 ( n4351 , n2830 , n10833 );
    nor g11688 ( n10086 , n7416 , n6722 );
    not g11689 ( n2472 , n3390 );
    or g11690 ( n1098 , n9489 , n2059 );
    or g11691 ( n6725 , n2662 , n6863 );
    xnor g11692 ( n8582 , n696 , n9000 );
    xnor g11693 ( n9999 , n10024 , n1967 );
    xnor g11694 ( n6812 , n7345 , n8895 );
    and g11695 ( n3353 , n9460 , n12452 );
    or g11696 ( n1132 , n715 , n11668 );
    not g11697 ( n10286 , n9620 );
    buf g11698 ( n3949 , n6274 );
    xnor g11699 ( n11467 , n9843 , n6528 );
    xnor g11700 ( n7347 , n6720 , n2584 );
    xnor g11701 ( n4507 , n4538 , n8667 );
    and g11702 ( n11473 , n8350 , n6000 );
    nor g11703 ( n660 , n4630 , n5312 );
    not g11704 ( n428 , n10599 );
    xnor g11705 ( n6169 , n9926 , n5175 );
    and g11706 ( n6949 , n7476 , n2301 );
    or g11707 ( n2811 , n9478 , n1144 );
    xnor g11708 ( n1714 , n9975 , n7482 );
    nor g11709 ( n4693 , n3885 , n6499 );
    xnor g11710 ( n10468 , n9122 , n7674 );
    not g11711 ( n12416 , n2252 );
    xnor g11712 ( n4069 , n12598 , n4437 );
    nor g11713 ( n11711 , n4081 , n9186 );
    not g11714 ( n5360 , n12381 );
    xnor g11715 ( n11579 , n4065 , n3226 );
    not g11716 ( n6587 , n10805 );
    or g11717 ( n5830 , n13202 , n7016 );
    or g11718 ( n11263 , n6133 , n4373 );
    not g11719 ( n10883 , n5920 );
    or g11720 ( n9191 , n11121 , n6899 );
    nor g11721 ( n8771 , n4992 , n2399 );
    xor g11722 ( n322 , n2546 , n7477 );
    xnor g11723 ( n13104 , n2700 , n3575 );
    and g11724 ( n7497 , n6670 , n7346 );
    xnor g11725 ( n2656 , n1954 , n1488 );
    or g11726 ( n9107 , n5008 , n4110 );
    or g11727 ( n4871 , n9383 , n5242 );
    and g11728 ( n4213 , n6014 , n6359 );
    not g11729 ( n5312 , n376 );
    or g11730 ( n3441 , n9711 , n8030 );
    or g11731 ( n2322 , n7503 , n11184 );
    xnor g11732 ( n11332 , n8070 , n8735 );
    and g11733 ( n9873 , n248 , n8769 );
    not g11734 ( n9962 , n5729 );
    and g11735 ( n1809 , n12229 , n4941 );
    xnor g11736 ( n10836 , n8130 , n3190 );
    nor g11737 ( n330 , n8866 , n8620 );
    xnor g11738 ( n4676 , n25 , n5901 );
    xnor g11739 ( n6201 , n4922 , n365 );
    xnor g11740 ( n12903 , n12558 , n12426 );
    or g11741 ( n9940 , n8104 , n7528 );
    or g11742 ( n9320 , n4519 , n7080 );
    and g11743 ( n8340 , n11504 , n10262 );
    and g11744 ( n1703 , n8594 , n12804 );
    and g11745 ( n7770 , n1951 , n6526 );
    and g11746 ( n4691 , n1630 , n5807 );
    not g11747 ( n8324 , n9300 );
    xnor g11748 ( n12749 , n12301 , n2180 );
    nor g11749 ( n10372 , n7676 , n1209 );
    or g11750 ( n7232 , n175 , n9369 );
    and g11751 ( n2315 , n10712 , n1864 );
    nor g11752 ( n11832 , n9855 , n7063 );
    xnor g11753 ( n10382 , n1841 , n10938 );
    or g11754 ( n4595 , n4967 , n8563 );
    not g11755 ( n4366 , n8233 );
    or g11756 ( n2559 , n7170 , n2631 );
    xor g11757 ( n8420 , n10225 , n10322 );
    or g11758 ( n4238 , n7783 , n12388 );
    not g11759 ( n9350 , n1826 );
    or g11760 ( n2480 , n9275 , n5744 );
    not g11761 ( n2581 , n10805 );
    or g11762 ( n3307 , n4063 , n1218 );
    xor g11763 ( n10680 , n1563 , n2951 );
    or g11764 ( n8525 , n423 , n9179 );
    not g11765 ( n2691 , n10190 );
    not g11766 ( n6358 , n12026 );
    not g11767 ( n10400 , n9846 );
    not g11768 ( n3804 , n1992 );
    or g11769 ( n8761 , n3726 , n7723 );
    or g11770 ( n11253 , n3911 , n9075 );
    or g11771 ( n1785 , n7658 , n8512 );
    or g11772 ( n11430 , n9648 , n8677 );
    and g11773 ( n3414 , n10258 , n7823 );
    nor g11774 ( n12782 , n11773 , n10116 );
    xnor g11775 ( n11257 , n3954 , n1792 );
    and g11776 ( n8431 , n9554 , n4252 );
    or g11777 ( n2952 , n10624 , n11708 );
    or g11778 ( n3192 , n3877 , n8874 );
    or g11779 ( n8740 , n12316 , n1422 );
    not g11780 ( n3534 , n1636 );
    or g11781 ( n347 , n8681 , n7723 );
    xnor g11782 ( n12002 , n7813 , n5742 );
    xnor g11783 ( n1555 , n4755 , n10289 );
    xnor g11784 ( n10831 , n2512 , n131 );
    and g11785 ( n8856 , n11068 , n9308 );
    xnor g11786 ( n3105 , n8380 , n7596 );
    xnor g11787 ( n8652 , n11295 , n1982 );
    xnor g11788 ( n11826 , n10983 , n12154 );
    or g11789 ( n11648 , n5148 , n4230 );
    xnor g11790 ( n9903 , n10516 , n5686 );
    and g11791 ( n8262 , n9169 , n1796 );
    xnor g11792 ( n8517 , n5902 , n6092 );
    or g11793 ( n3975 , n10650 , n921 );
    or g11794 ( n920 , n12254 , n1043 );
    or g11795 ( n12129 , n6828 , n11796 );
    and g11796 ( n12244 , n12150 , n4145 );
    not g11797 ( n1965 , n4557 );
    and g11798 ( n4346 , n1073 , n6983 );
    nor g11799 ( n6560 , n12470 , n7656 );
    xnor g11800 ( n180 , n5329 , n5701 );
    and g11801 ( n12850 , n3804 , n12941 );
    xor g11802 ( n11490 , n1202 , n10808 );
    xnor g11803 ( n2451 , n4719 , n11412 );
    or g11804 ( n7938 , n10977 , n8348 );
    xnor g11805 ( n5391 , n11907 , n12327 );
    not g11806 ( n11320 , n4330 );
    or g11807 ( n21 , n2255 , n9314 );
    xnor g11808 ( n7603 , n8331 , n1046 );
    or g11809 ( n1904 , n755 , n3598 );
    or g11810 ( n6900 , n12630 , n1240 );
    or g11811 ( n8906 , n10423 , n264 );
    or g11812 ( n10724 , n10854 , n837 );
    xor g11813 ( n12632 , n6633 , n11607 );
    or g11814 ( n8361 , n6630 , n4373 );
    nor g11815 ( n5043 , n6212 , n11219 );
    nor g11816 ( n314 , n12688 , n4270 );
    xnor g11817 ( n2505 , n12840 , n4611 );
    or g11818 ( n7973 , n305 , n5724 );
    or g11819 ( n37 , n7358 , n1571 );
    nor g11820 ( n3254 , n2284 , n8770 );
    nor g11821 ( n805 , n1716 , n11438 );
    or g11822 ( n10231 , n11910 , n2449 );
    not g11823 ( n8868 , n13058 );
    xor g11824 ( n66 , n2595 , n8760 );
    xnor g11825 ( n58 , n8766 , n6874 );
    not g11826 ( n11868 , n10451 );
    nor g11827 ( n10133 , n2932 , n11182 );
    xnor g11828 ( n12996 , n2417 , n4319 );
    nor g11829 ( n12108 , n2522 , n9998 );
    or g11830 ( n8954 , n6099 , n1043 );
    or g11831 ( n9355 , n11121 , n5802 );
    xnor g11832 ( n11731 , n5851 , n7413 );
    and g11833 ( n1154 , n8307 , n4940 );
    and g11834 ( n5510 , n8447 , n12292 );
    or g11835 ( n12790 , n3676 , n3640 );
    or g11836 ( n11773 , n10266 , n9745 );
    not g11837 ( n12537 , n4964 );
    not g11838 ( n3572 , n1982 );
    or g11839 ( n5499 , n6486 , n12501 );
    xnor g11840 ( n13002 , n11190 , n10740 );
    xnor g11841 ( n11863 , n740 , n11738 );
    xnor g11842 ( n2693 , n12452 , n9115 );
    xnor g11843 ( n7593 , n9124 , n7229 );
    xnor g11844 ( n10868 , n2710 , n541 );
    not g11845 ( n6875 , n9591 );
    or g11846 ( n8168 , n8876 , n12487 );
    xnor g11847 ( n8701 , n2280 , n2185 );
    xnor g11848 ( n4140 , n7999 , n8171 );
    and g11849 ( n690 , n10611 , n11307 );
    xnor g11850 ( n2312 , n6172 , n5756 );
    and g11851 ( n11259 , n1062 , n12310 );
    and g11852 ( n11639 , n6329 , n4883 );
    xnor g11853 ( n3844 , n8235 , n3100 );
    xnor g11854 ( n11160 , n5123 , n2029 );
    xnor g11855 ( n756 , n4759 , n5116 );
    xnor g11856 ( n5481 , n2651 , n10933 );
    not g11857 ( n312 , n12112 );
    xor g11858 ( n12367 , n8838 , n3494 );
    xnor g11859 ( n13161 , n7979 , n3392 );
    and g11860 ( n2978 , n2874 , n12815 );
    not g11861 ( n3126 , n12965 );
    xnor g11862 ( n3014 , n13014 , n12751 );
    or g11863 ( n11203 , n10143 , n4373 );
    or g11864 ( n8432 , n9171 , n6257 );
    not g11865 ( n10574 , n394 );
    nor g11866 ( n12376 , n7485 , n4889 );
    or g11867 ( n294 , n5157 , n12049 );
    xnor g11868 ( n5052 , n6065 , n1120 );
    and g11869 ( n7010 , n9497 , n6330 );
    xnor g11870 ( n6397 , n12879 , n2494 );
    or g11871 ( n8446 , n2022 , n1193 );
    xnor g11872 ( n8114 , n10915 , n10226 );
    xnor g11873 ( n9419 , n3088 , n7121 );
    and g11874 ( n8260 , n12738 , n3543 );
    or g11875 ( n10529 , n7953 , n11051 );
    and g11876 ( n9413 , n3372 , n5544 );
    or g11877 ( n1713 , n12465 , n11668 );
    not g11878 ( n6878 , n9293 );
    not g11879 ( n9607 , n5647 );
    and g11880 ( n76 , n11104 , n6157 );
    and g11881 ( n8614 , n3326 , n387 );
    xnor g11882 ( n2756 , n9522 , n10635 );
    and g11883 ( n8552 , n9930 , n3980 );
    xnor g11884 ( n11371 , n686 , n2885 );
    or g11885 ( n3599 , n2067 , n8096 );
    or g11886 ( n4558 , n8977 , n10179 );
    or g11887 ( n840 , n1778 , n9572 );
    xnor g11888 ( n4690 , n12025 , n8314 );
    not g11889 ( n5949 , n6392 );
    or g11890 ( n662 , n11225 , n2133 );
    xnor g11891 ( n6931 , n3101 , n2290 );
    xnor g11892 ( n12096 , n6753 , n4812 );
    and g11893 ( n6455 , n1333 , n8842 );
    xnor g11894 ( n5882 , n7379 , n9165 );
    or g11895 ( n11690 , n5498 , n8800 );
    or g11896 ( n12984 , n11404 , n5797 );
    xnor g11897 ( n2859 , n10221 , n5812 );
    nor g11898 ( n6656 , n9374 , n3389 );
    xnor g11899 ( n6820 , n1242 , n12173 );
    xnor g11900 ( n9956 , n4459 , n1662 );
    xnor g11901 ( n6030 , n8813 , n2470 );
    and g11902 ( n10740 , n3006 , n10451 );
    not g11903 ( n10641 , n2737 );
    not g11904 ( n3570 , n11285 );
    xnor g11905 ( n9875 , n11334 , n9359 );
    not g11906 ( n5550 , n11665 );
    or g11907 ( n6067 , n795 , n10135 );
    xnor g11908 ( n2316 , n10150 , n12054 );
    nor g11909 ( n6564 , n9526 , n10146 );
    and g11910 ( n7682 , n11345 , n5250 );
    xnor g11911 ( n3277 , n7776 , n518 );
    or g11912 ( n12878 , n10991 , n8268 );
    or g11913 ( n10220 , n12295 , n3981 );
    or g11914 ( n1665 , n11370 , n4724 );
    or g11915 ( n13177 , n398 , n10813 );
    not g11916 ( n3460 , n9570 );
    or g11917 ( n11497 , n10137 , n2133 );
    xnor g11918 ( n7332 , n1419 , n30 );
    nor g11919 ( n391 , n2072 , n8481 );
    not g11920 ( n8044 , n1762 );
    xnor g11921 ( n858 , n6975 , n7871 );
    xnor g11922 ( n10159 , n4033 , n3552 );
    and g11923 ( n496 , n9328 , n5948 );
    xnor g11924 ( n9185 , n10844 , n5042 );
    or g11925 ( n2358 , n12648 , n9962 );
    or g11926 ( n3408 , n3259 , n6732 );
    not g11927 ( n1358 , n976 );
    and g11928 ( n6636 , n10039 , n11110 );
    xnor g11929 ( n11763 , n1299 , n5397 );
    and g11930 ( n7988 , n4085 , n10348 );
    xnor g11931 ( n11953 , n6821 , n1369 );
    or g11932 ( n5774 , n69 , n12273 );
    xnor g11933 ( n7462 , n2466 , n11068 );
    xnor g11934 ( n12570 , n5419 , n10069 );
    and g11935 ( n9088 , n12630 , n1240 );
    and g11936 ( n3600 , n11818 , n10022 );
    xnor g11937 ( n12207 , n4284 , n9166 );
    xnor g11938 ( n1061 , n7193 , n9933 );
    nor g11939 ( n3776 , n242 , n6941 );
    not g11940 ( n11783 , n10025 );
    or g11941 ( n2357 , n9129 , n1026 );
    and g11942 ( n12567 , n12370 , n12824 );
    xnor g11943 ( n13163 , n3907 , n7513 );
    and g11944 ( n4534 , n7114 , n4192 );
    xnor g11945 ( n12146 , n9049 , n1577 );
    or g11946 ( n8208 , n7997 , n4959 );
    or g11947 ( n11803 , n3836 , n1103 );
    and g11948 ( n10328 , n5372 , n4481 );
    nor g11949 ( n1848 , n7952 , n9571 );
    nor g11950 ( n13206 , n8389 , n7192 );
    or g11951 ( n11692 , n1571 , n8490 );
    xnor g11952 ( n7435 , n6148 , n6458 );
    or g11953 ( n11642 , n10499 , n11843 );
    xnor g11954 ( n3368 , n10477 , n10484 );
    xnor g11955 ( n6396 , n9928 , n12314 );
    and g11956 ( n8094 , n7765 , n10906 );
    nor g11957 ( n10242 , n7156 , n1932 );
    and g11958 ( n11281 , n1489 , n10806 );
    and g11959 ( n2334 , n7544 , n198 );
    xnor g11960 ( n7053 , n3543 , n9367 );
    and g11961 ( n11988 , n9216 , n9475 );
    not g11962 ( n4967 , n6085 );
    or g11963 ( n11956 , n3249 , n3161 );
    and g11964 ( n12017 , n7475 , n8982 );
    or g11965 ( n8788 , n6367 , n10319 );
    nor g11966 ( n1108 , n7885 , n1187 );
    nor g11967 ( n8947 , n8567 , n6718 );
    xnor g11968 ( n8691 , n7136 , n10698 );
    xnor g11969 ( n12947 , n7375 , n12618 );
    not g11970 ( n6743 , n22 );
    not g11971 ( n6990 , n5475 );
    xnor g11972 ( n13160 , n5316 , n8320 );
    not g11973 ( n10527 , n10122 );
    not g11974 ( n12153 , n11411 );
    and g11975 ( n10589 , n7669 , n9101 );
    xnor g11976 ( n1119 , n8299 , n11752 );
    not g11977 ( n1052 , n6826 );
    not g11978 ( n6504 , n498 );
    or g11979 ( n7418 , n8615 , n8268 );
    xnor g11980 ( n12151 , n1977 , n849 );
    not g11981 ( n9339 , n11891 );
    xnor g11982 ( n4860 , n3148 , n4902 );
    not g11983 ( n4722 , n3677 );
    and g11984 ( n2071 , n5811 , n8202 );
    not g11985 ( n913 , n6561 );
    or g11986 ( n6566 , n11868 , n5076 );
    xnor g11987 ( n7928 , n4480 , n10598 );
    or g11988 ( n3442 , n567 , n11833 );
    xnor g11989 ( n437 , n720 , n5600 );
    xnor g11990 ( n12217 , n1456 , n9333 );
    or g11991 ( n3214 , n1367 , n5971 );
    not g11992 ( n13039 , n3769 );
    and g11993 ( n8493 , n8034 , n9496 );
    and g11994 ( n2308 , n2607 , n6640 );
    and g11995 ( n8016 , n9418 , n1214 );
    nor g11996 ( n4922 , n3872 , n9301 );
    and g11997 ( n12876 , n4441 , n2600 );
    and g11998 ( n4033 , n8046 , n1410 );
    not g11999 ( n12967 , n4470 );
    xnor g12000 ( n801 , n10965 , n2826 );
    xnor g12001 ( n5657 , n6494 , n4438 );
    xnor g12002 ( n5587 , n2774 , n4415 );
    xnor g12003 ( n5051 , n11039 , n11873 );
    not g12004 ( n1105 , n587 );
    and g12005 ( n792 , n4138 , n239 );
    xnor g12006 ( n3431 , n6206 , n2170 );
    not g12007 ( n11871 , n761 );
    xnor g12008 ( n8553 , n4271 , n9348 );
    not g12009 ( n12221 , n8156 );
    or g12010 ( n8042 , n2296 , n7254 );
    and g12011 ( n5209 , n655 , n2914 );
    nor g12012 ( n8075 , n4439 , n2956 );
    buf g12013 ( n12388 , n7424 );
    or g12014 ( n1684 , n5039 , n7821 );
    or g12015 ( n12516 , n1651 , n6265 );
    not g12016 ( n9068 , n3709 );
    and g12017 ( n12498 , n12013 , n1632 );
    xor g12018 ( n908 , n10293 , n5480 );
    nor g12019 ( n10222 , n12715 , n11027 );
    xnor g12020 ( n3100 , n12533 , n3694 );
    or g12021 ( n4962 , n2692 , n3981 );
    or g12022 ( n4277 , n734 , n493 );
    xnor g12023 ( n7092 , n1974 , n1595 );
    or g12024 ( n12874 , n5795 , n5510 );
    not g12025 ( n2352 , n10657 );
    xnor g12026 ( n1196 , n4651 , n12118 );
    not g12027 ( n8710 , n10343 );
    not g12028 ( n8892 , n10479 );
    or g12029 ( n6753 , n10018 , n3981 );
    or g12030 ( n8120 , n9350 , n10627 );
    or g12031 ( n3957 , n3225 , n11668 );
    xnor g12032 ( n12301 , n9516 , n11789 );
    xnor g12033 ( n8746 , n13205 , n4310 );
    or g12034 ( n11313 , n3696 , n447 );
    not g12035 ( n9635 , n1603 );
    not g12036 ( n9276 , n9685 );
    or g12037 ( n7289 , n1416 , n10696 );
    not g12038 ( n8360 , n6826 );
    xnor g12039 ( n10379 , n6412 , n12763 );
    or g12040 ( n6671 , n5749 , n8534 );
    or g12041 ( n8574 , n440 , n5431 );
    xnor g12042 ( n12160 , n7123 , n1119 );
    and g12043 ( n11079 , n5508 , n861 );
    xnor g12044 ( n7804 , n8276 , n2905 );
    nor g12045 ( n7489 , n11873 , n4529 );
    or g12046 ( n7947 , n12713 , n7082 );
    xnor g12047 ( n12305 , n10077 , n9229 );
    and g12048 ( n4583 , n2353 , n5542 );
    xor g12049 ( n12101 , n10575 , n5170 );
    nor g12050 ( n3462 , n10152 , n5368 );
    xnor g12051 ( n1612 , n590 , n12977 );
    xnor g12052 ( n6773 , n7645 , n1200 );
    not g12053 ( n11132 , n1273 );
    not g12054 ( n8212 , n7051 );
    or g12055 ( n11392 , n5271 , n8490 );
    or g12056 ( n9881 , n5634 , n5242 );
    and g12057 ( n10289 , n1705 , n2788 );
    xnor g12058 ( n9457 , n924 , n2938 );
    not g12059 ( n4796 , n13058 );
    or g12060 ( n12780 , n5581 , n5173 );
    xnor g12061 ( n6324 , n11187 , n6474 );
    xnor g12062 ( n10775 , n6809 , n11000 );
    or g12063 ( n8393 , n4022 , n177 );
    xnor g12064 ( n12703 , n733 , n2200 );
    and g12065 ( n3792 , n10650 , n921 );
    xnor g12066 ( n1535 , n11472 , n11949 );
    and g12067 ( n2918 , n3318 , n5714 );
    and g12068 ( n1564 , n11411 , n6168 );
    not g12069 ( n2109 , n10142 );
    or g12070 ( n7019 , n1185 , n1669 );
    and g12071 ( n11279 , n12086 , n11988 );
    xnor g12072 ( n11896 , n1205 , n12146 );
    or g12073 ( n4937 , n9080 , n9159 );
    xnor g12074 ( n827 , n9726 , n8962 );
    or g12075 ( n9927 , n13051 , n2544 );
    and g12076 ( n6973 , n7386 , n5745 );
    not g12077 ( n2278 , n8940 );
    xnor g12078 ( n5918 , n11961 , n12571 );
    and g12079 ( n13105 , n2713 , n7325 );
    not g12080 ( n2332 , n3076 );
    xnor g12081 ( n6994 , n10306 , n8678 );
    or g12082 ( n11168 , n13082 , n7221 );
    xnor g12083 ( n4834 , n1410 , n8046 );
    or g12084 ( n4627 , n5329 , n4503 );
    or g12085 ( n10260 , n756 , n5221 );
    nor g12086 ( n11186 , n6838 , n12587 );
    xnor g12087 ( n11043 , n1730 , n7077 );
    and g12088 ( n11290 , n10201 , n7204 );
    xnor g12089 ( n2001 , n4556 , n135 );
    or g12090 ( n12322 , n3630 , n12328 );
    or g12091 ( n4608 , n3986 , n5716 );
    not g12092 ( n3489 , n10613 );
    and g12093 ( n8874 , n6516 , n9085 );
    or g12094 ( n5659 , n10696 , n9075 );
    not g12095 ( n142 , n2370 );
    xnor g12096 ( n5207 , n7668 , n12232 );
    not g12097 ( n8864 , n9270 );
    and g12098 ( n10147 , n2057 , n10063 );
    or g12099 ( n9728 , n4080 , n7723 );
    or g12100 ( n5352 , n9309 , n8005 );
    or g12101 ( n5113 , n5694 , n4947 );
    nor g12102 ( n6437 , n2358 , n8462 );
    xor g12103 ( n11482 , n10928 , n4155 );
    and g12104 ( n1895 , n7301 , n1274 );
    and g12105 ( n4807 , n2800 , n2466 );
    and g12106 ( n1032 , n11815 , n191 );
    xnor g12107 ( n8737 , n9173 , n13100 );
    or g12108 ( n8064 , n6557 , n1570 );
    nor g12109 ( n10847 , n11384 , n11141 );
    or g12110 ( n2469 , n8639 , n10935 );
    and g12111 ( n3206 , n13085 , n12696 );
    or g12112 ( n9949 , n5358 , n5011 );
    xnor g12113 ( n10423 , n8628 , n1021 );
    or g12114 ( n11065 , n5757 , n9147 );
    or g12115 ( n4757 , n3158 , n4724 );
    or g12116 ( n9708 , n9934 , n12388 );
    or g12117 ( n5660 , n338 , n5076 );
    buf g12118 ( n7530 , n6210 );
    xnor g12119 ( n108 , n3841 , n1829 );
    nor g12120 ( n8215 , n4507 , n1342 );
    and g12121 ( n12526 , n8416 , n12590 );
    not g12122 ( n650 , n8233 );
    or g12123 ( n6388 , n7865 , n3149 );
    or g12124 ( n6793 , n1353 , n9159 );
    not g12125 ( n1357 , n3543 );
    and g12126 ( n12068 , n5676 , n3530 );
    nor g12127 ( n7922 , n2621 , n3220 );
    xnor g12128 ( n4996 , n11799 , n8669 );
    or g12129 ( n866 , n1248 , n10878 );
    nor g12130 ( n5541 , n966 , n7336 );
    not g12131 ( n7257 , n5277 );
    xnor g12132 ( n11608 , n12682 , n9362 );
    or g12133 ( n5301 , n11742 , n13125 );
    or g12134 ( n12510 , n5415 , n167 );
    not g12135 ( n5168 , n11734 );
    or g12136 ( n6338 , n4370 , n8348 );
    xnor g12137 ( n1502 , n4383 , n3566 );
    not g12138 ( n11723 , n4330 );
    xnor g12139 ( n7531 , n5224 , n37 );
    nor g12140 ( n9427 , n9879 , n12983 );
    xnor g12141 ( n10803 , n5100 , n10185 );
    or g12142 ( n7807 , n8064 , n6299 );
    not g12143 ( n11635 , n7161 );
    or g12144 ( n1376 , n2301 , n7476 );
    and g12145 ( n11841 , n6139 , n6490 );
    or g12146 ( n2553 , n1067 , n1195 );
    or g12147 ( n12528 , n5265 , n10871 );
    xnor g12148 ( n9613 , n10219 , n11411 );
    nor g12149 ( n8738 , n3357 , n3012 );
    or g12150 ( n3377 , n6726 , n10179 );
    xnor g12151 ( n2180 , n2395 , n1615 );
    not g12152 ( n10032 , n11734 );
    or g12153 ( n1359 , n318 , n1985 );
    and g12154 ( n4004 , n6572 , n5888 );
    or g12155 ( n10717 , n4000 , n4223 );
    not g12156 ( n4098 , n11640 );
    or g12157 ( n13149 , n4161 , n2970 );
    or g12158 ( n11250 , n4665 , n10871 );
    xnor g12159 ( n4142 , n1575 , n8622 );
    not g12160 ( n3493 , n10860 );
    not g12161 ( n6025 , n322 );
    not g12162 ( n1320 , n11109 );
    or g12163 ( n231 , n4969 , n3276 );
    or g12164 ( n10180 , n6518 , n557 );
    and g12165 ( n7069 , n654 , n230 );
    not g12166 ( n2747 , n1397 );
    not g12167 ( n13122 , n4376 );
    nor g12168 ( n10735 , n2297 , n3421 );
    xnor g12169 ( n2585 , n3941 , n12658 );
    and g12170 ( n13007 , n12846 , n12486 );
    and g12171 ( n10278 , n11232 , n7243 );
    or g12172 ( n6393 , n4771 , n12332 );
    or g12173 ( n2356 , n12249 , n8563 );
    or g12174 ( n5773 , n11010 , n9046 );
    and g12175 ( n1774 , n11294 , n10748 );
    xnor g12176 ( n1443 , n4825 , n7165 );
    xnor g12177 ( n2170 , n12236 , n4835 );
    not g12178 ( n882 , n6965 );
    or g12179 ( n10248 , n8600 , n1804 );
    xnor g12180 ( n10864 , n5130 , n10113 );
    buf g12181 ( n9159 , n2406 );
    or g12182 ( n3933 , n4587 , n9251 );
    or g12183 ( n13102 , n9416 , n7203 );
    not g12184 ( n5265 , n9669 );
    or g12185 ( n6242 , n9934 , n1570 );
    nor g12186 ( n10358 , n2878 , n12891 );
    or g12187 ( n12556 , n5404 , n5721 );
    not g12188 ( n2726 , n9475 );
    or g12189 ( n11286 , n7836 , n11768 );
    xnor g12190 ( n12197 , n314 , n11253 );
    nor g12191 ( n1461 , n5567 , n11563 );
    and g12192 ( n1609 , n8449 , n1533 );
    or g12193 ( n9071 , n12843 , n8988 );
    not g12194 ( n4066 , n7745 );
    or g12195 ( n175 , n2041 , n584 );
    nor g12196 ( n3793 , n10765 , n852 );
    nor g12197 ( n1898 , n5861 , n7548 );
    or g12198 ( n4934 , n3364 , n11007 );
    not g12199 ( n6402 , n11339 );
    or g12200 ( n1091 , n4108 , n3554 );
    or g12201 ( n3986 , n10761 , n6265 );
    and g12202 ( n2002 , n5725 , n4451 );
    and g12203 ( n2392 , n10180 , n10749 );
    not g12204 ( n2485 , n624 );
    or g12205 ( n3730 , n8615 , n4230 );
    not g12206 ( n10616 , n2513 );
    and g12207 ( n12064 , n12342 , n9977 );
    nor g12208 ( n4007 , n976 , n260 );
    and g12209 ( n11457 , n2570 , n6923 );
    xnor g12210 ( n12314 , n12809 , n11267 );
    or g12211 ( n1509 , n9016 , n206 );
    or g12212 ( n11512 , n12859 , n10971 );
    xnor g12213 ( n4977 , n1470 , n10614 );
    and g12214 ( n4405 , n10598 , n4480 );
    not g12215 ( n12957 , n937 );
    or g12216 ( n1264 , n11799 , n3187 );
    xnor g12217 ( n6177 , n6196 , n12831 );
    and g12218 ( n8408 , n10113 , n7411 );
    not g12219 ( n4955 , n5454 );
    xnor g12220 ( n8889 , n4692 , n556 );
    or g12221 ( n11502 , n544 , n322 );
    or g12222 ( n7131 , n3522 , n8086 );
    or g12223 ( n3009 , n2226 , n9309 );
    and g12224 ( n10926 , n6027 , n6898 );
    and g12225 ( n625 , n5638 , n6888 );
    xnor g12226 ( n1214 , n1297 , n6984 );
    xnor g12227 ( n11944 , n903 , n12197 );
    xnor g12228 ( n8178 , n2936 , n9356 );
    and g12229 ( n6060 , n1238 , n3819 );
    and g12230 ( n2609 , n5613 , n12555 );
    not g12231 ( n967 , n5322 );
    xnor g12232 ( n12218 , n2101 , n4794 );
    xnor g12233 ( n11769 , n11971 , n12102 );
    or g12234 ( n3602 , n8980 , n7509 );
    or g12235 ( n8378 , n8862 , n12072 );
    xnor g12236 ( n11993 , n10861 , n6736 );
    or g12237 ( n4853 , n1725 , n12948 );
    and g12238 ( n2117 , n3837 , n6327 );
    not g12239 ( n406 , n10657 );
    nor g12240 ( n12152 , n7929 , n12106 );
    xnor g12241 ( n11819 , n783 , n8893 );
    xnor g12242 ( n10776 , n8135 , n11536 );
    not g12243 ( n8645 , n11835 );
    and g12244 ( n9486 , n7951 , n7921 );
    xnor g12245 ( n5022 , n7414 , n8845 );
    not g12246 ( n237 , n10642 );
    or g12247 ( n2240 , n10883 , n9075 );
    xor g12248 ( n9437 , n10419 , n2000 );
    xnor g12249 ( n1669 , n9676 , n11367 );
    or g12250 ( n6191 , n202 , n1985 );
    not g12251 ( n3690 , n880 );
    or g12252 ( n8880 , n10591 , n7723 );
    nor g12253 ( n1658 , n11496 , n7893 );
    not g12254 ( n3866 , n3815 );
    xnor g12255 ( n11536 , n12140 , n3989 );
    or g12256 ( n434 , n1651 , n4936 );
    xor g12257 ( n10101 , n10392 , n9655 );
    or g12258 ( n6961 , n9154 , n12501 );
    xnor g12259 ( n13022 , n9637 , n3649 );
    and g12260 ( n4074 , n3335 , n11178 );
    xnor g12261 ( n2432 , n4521 , n2497 );
    xnor g12262 ( n7553 , n2841 , n11528 );
    xnor g12263 ( n3181 , n11592 , n4656 );
    nor g12264 ( n1462 , n7552 , n10793 );
    or g12265 ( n2088 , n6375 , n10319 );
    xnor g12266 ( n11484 , n12581 , n12905 );
    not g12267 ( n5037 , n4413 );
    or g12268 ( n17 , n11683 , n10319 );
    and g12269 ( n4888 , n9353 , n3085 );
    xnor g12270 ( n5219 , n12804 , n8594 );
    xnor g12271 ( n11151 , n1758 , n6034 );
    xnor g12272 ( n7967 , n1810 , n1755 );
    not g12273 ( n11664 , n5375 );
    xnor g12274 ( n9034 , n2799 , n6544 );
    not g12275 ( n2183 , n9591 );
    and g12276 ( n4164 , n1906 , n6095 );
    or g12277 ( n10683 , n9917 , n11446 );
    or g12278 ( n9835 , n4370 , n4724 );
    nor g12279 ( n3039 , n1352 , n8037 );
    not g12280 ( n5782 , n411 );
    not g12281 ( n12357 , n4015 );
    or g12282 ( n250 , n11356 , n8702 );
    and g12283 ( n10897 , n5456 , n8833 );
    and g12284 ( n4695 , n1889 , n4320 );
    or g12285 ( n4607 , n12911 , n2792 );
    xnor g12286 ( n10511 , n10217 , n2837 );
    nor g12287 ( n1824 , n8067 , n10817 );
    or g12288 ( n9954 , n8739 , n8036 );
    xnor g12289 ( n8201 , n7230 , n3622 );
    or g12290 ( n11374 , n12758 , n4724 );
    xnor g12291 ( n6765 , n1601 , n7384 );
    or g12292 ( n9161 , n12768 , n1570 );
    or g12293 ( n3266 , n1772 , n7701 );
    xnor g12294 ( n6702 , n7852 , n1770 );
    or g12295 ( n1546 , n6381 , n4947 );
    and g12296 ( n12609 , n4891 , n6360 );
    or g12297 ( n11183 , n1638 , n10029 );
    xnor g12298 ( n5095 , n5121 , n4516 );
    or g12299 ( n7354 , n542 , n6265 );
    nor g12300 ( n7912 , n11709 , n3447 );
    xnor g12301 ( n6400 , n5453 , n12836 );
    or g12302 ( n3492 , n5407 , n3648 );
    nor g12303 ( n8417 , n6535 , n4064 );
    nor g12304 ( n9254 , n12467 , n9561 );
    and g12305 ( n5277 , n6894 , n6980 );
    or g12306 ( n4810 , n5182 , n11521 );
    and g12307 ( n4249 , n5526 , n1691 );
    or g12308 ( n12449 , n12617 , n9808 );
    xnor g12309 ( n10342 , n7802 , n5336 );
    xnor g12310 ( n2101 , n267 , n12762 );
    nor g12311 ( n8727 , n5251 , n4065 );
    xnor g12312 ( n3606 , n890 , n7209 );
    or g12313 ( n968 , n11113 , n9223 );
    not g12314 ( n3784 , n12065 );
    nor g12315 ( n176 , n1349 , n4259 );
    xnor g12316 ( n2206 , n6371 , n10071 );
    or g12317 ( n3530 , n3460 , n12695 );
    and g12318 ( n6047 , n7554 , n591 );
    not g12319 ( n719 , n10745 );
    not g12320 ( n10900 , n1364 );
    and g12321 ( n2102 , n7514 , n7778 );
    nor g12322 ( n12467 , n5005 , n13110 );
    buf g12323 ( n8348 , n3671 );
    not g12324 ( n9310 , n5470 );
    xnor g12325 ( n6447 , n7256 , n832 );
    not g12326 ( n651 , n9027 );
    not g12327 ( n3633 , n6973 );
    not g12328 ( n3854 , n353 );
    or g12329 ( n5784 , n3225 , n8490 );
    nor g12330 ( n8275 , n9033 , n5722 );
    not g12331 ( n5847 , n6820 );
    or g12332 ( n4756 , n9248 , n5006 );
    xnor g12333 ( n1613 , n3339 , n12878 );
    not g12334 ( n3336 , n6189 );
    and g12335 ( n4378 , n5911 , n3603 );
    xnor g12336 ( n9839 , n2994 , n8110 );
    or g12337 ( n5531 , n10139 , n8101 );
    not g12338 ( n4430 , n1225 );
    xnor g12339 ( n11913 , n11936 , n3252 );
    nor g12340 ( n10706 , n1640 , n1704 );
    and g12341 ( n10075 , n10738 , n11673 );
    xnor g12342 ( n11416 , n10385 , n3863 );
    not g12343 ( n1258 , n6597 );
    or g12344 ( n2806 , n872 , n7252 );
    or g12345 ( n11943 , n7546 , n2490 );
    xnor g12346 ( n9166 , n10325 , n1929 );
    not g12347 ( n445 , n5065 );
    not g12348 ( n4716 , n8369 );
    and g12349 ( n6150 , n11927 , n1300 );
    or g12350 ( n3915 , n11263 , n13081 );
    nor g12351 ( n6752 , n3171 , n5154 );
    not g12352 ( n5694 , n3677 );
    and g12353 ( n3143 , n3359 , n7570 );
    or g12354 ( n784 , n930 , n10463 );
    nor g12355 ( n5255 , n4304 , n11885 );
    and g12356 ( n7155 , n316 , n4084 );
    xnor g12357 ( n12414 , n11793 , n11177 );
    nor g12358 ( n1468 , n11534 , n3440 );
    not g12359 ( n1402 , n10606 );
    xnor g12360 ( n7736 , n12013 , n8222 );
    or g12361 ( n9807 , n6672 , n4420 );
    and g12362 ( n875 , n13201 , n834 );
    buf g12363 ( n3225 , n6193 );
    not g12364 ( n8950 , n11429 );
    or g12365 ( n3563 , n13028 , n8777 );
    xnor g12366 ( n3438 , n11900 , n10816 );
    xnor g12367 ( n3808 , n2286 , n647 );
    or g12368 ( n8068 , n7637 , n12171 );
    and g12369 ( n6082 , n3800 , n10269 );
    and g12370 ( n13176 , n11408 , n7911 );
    or g12371 ( n9293 , n8865 , n8819 );
    or g12372 ( n5719 , n5932 , n2633 );
    and g12373 ( n351 , n4537 , n5962 );
    or g12374 ( n4251 , n48 , n3981 );
    not g12375 ( n4689 , n3797 );
    or g12376 ( n12337 , n332 , n12733 );
    or g12377 ( n1560 , n787 , n2059 );
    or g12378 ( n3273 , n987 , n5242 );
    nor g12379 ( n10054 , n11070 , n3503 );
    xnor g12380 ( n9858 , n8616 , n799 );
    not g12381 ( n4484 , n919 );
    not g12382 ( n11779 , n7659 );
    xnor g12383 ( n8473 , n2347 , n12346 );
    and g12384 ( n5184 , n4356 , n4010 );
    not g12385 ( n12069 , n11537 );
    nor g12386 ( n2748 , n6750 , n7572 );
    and g12387 ( n6141 , n11247 , n2812 );
    not g12388 ( n1587 , n2498 );
    not g12389 ( n9497 , n1563 );
    or g12390 ( n12340 , n3498 , n10106 );
    nor g12391 ( n9405 , n11215 , n2375 );
    xnor g12392 ( n10955 , n7882 , n1923 );
    and g12393 ( n3551 , n6731 , n11901 );
    and g12394 ( n6821 , n11513 , n312 );
    or g12395 ( n9487 , n98 , n8702 );
    or g12396 ( n1786 , n1645 , n6169 );
    and g12397 ( n6467 , n3760 , n5446 );
    and g12398 ( n4024 , n9387 , n9997 );
    xnor g12399 ( n8080 , n12270 , n1604 );
    not g12400 ( n7127 , n7452 );
    not g12401 ( n2022 , n5052 );
    or g12402 ( n5529 , n7176 , n8366 );
    or g12403 ( n12256 , n8891 , n3961 );
    not g12404 ( n4208 , n12289 );
    xor g12405 ( n2159 , n7272 , n195 );
    xnor g12406 ( n1845 , n6322 , n10649 );
    nor g12407 ( n3388 , n10829 , n6071 );
    and g12408 ( n4662 , n11 , n8956 );
    xnor g12409 ( n12905 , n6314 , n8913 );
    and g12410 ( n7696 , n10212 , n11947 );
    not g12411 ( n7710 , n7906 );
    and g12412 ( n4546 , n2795 , n11654 );
    and g12413 ( n2421 , n4836 , n12883 );
    or g12414 ( n3255 , n3505 , n9537 );
    or g12415 ( n500 , n7782 , n4169 );
    and g12416 ( n528 , n8940 , n8290 );
    and g12417 ( n605 , n11914 , n12760 );
    and g12418 ( n4121 , n3006 , n12853 );
    or g12419 ( n3605 , n13154 , n6635 );
    or g12420 ( n3679 , n5478 , n6293 );
    or g12421 ( n1439 , n10974 , n8534 );
    nor g12422 ( n242 , n7699 , n8703 );
    and g12423 ( n8480 , n12942 , n475 );
    xnor g12424 ( n12286 , n9642 , n714 );
    not g12425 ( n2264 , n10606 );
    xnor g12426 ( n7754 , n27 , n11353 );
    or g12427 ( n1765 , n4221 , n3225 );
    not g12428 ( n4696 , n4114 );
    xnor g12429 ( n12524 , n12829 , n6461 );
    not g12430 ( n2910 , n5075 );
    or g12431 ( n10097 , n12024 , n8568 );
    and g12432 ( n3231 , n6168 , n4470 );
    or g12433 ( n10497 , n11218 , n2958 );
    xnor g12434 ( n5102 , n8807 , n12275 );
    or g12435 ( n1427 , n5679 , n11107 );
    xnor g12436 ( n2009 , n2533 , n8042 );
    not g12437 ( n1151 , n4303 );
    and g12438 ( n5218 , n6926 , n4418 );
    or g12439 ( n5872 , n10893 , n6364 );
    or g12440 ( n385 , n12032 , n12388 );
    xnor g12441 ( n12039 , n6828 , n4917 );
    and g12442 ( n12390 , n7371 , n8438 );
    nor g12443 ( n6941 , n4965 , n339 );
    or g12444 ( n2850 , n877 , n11898 );
    xnor g12445 ( n7094 , n707 , n4307 );
    not g12446 ( n8848 , n6021 );
    xnor g12447 ( n11830 , n11584 , n9738 );
    nor g12448 ( n11532 , n7236 , n2099 );
    xnor g12449 ( n960 , n7618 , n4617 );
    and g12450 ( n638 , n1896 , n11005 );
    or g12451 ( n3124 , n924 , n5776 );
    xnor g12452 ( n775 , n11046 , n6030 );
    not g12453 ( n8661 , n7161 );
    or g12454 ( n3847 , n572 , n11375 );
    or g12455 ( n6348 , n12878 , n8118 );
    or g12456 ( n5911 , n12082 , n4786 );
    or g12457 ( n6778 , n8681 , n5797 );
    or g12458 ( n13196 , n11054 , n1463 );
    not g12459 ( n12383 , n834 );
    or g12460 ( n10753 , n9674 , n1255 );
    or g12461 ( n4480 , n2487 , n5242 );
    xnor g12462 ( n3332 , n3139 , n9470 );
    nor g12463 ( n9463 , n5737 , n7643 );
    and g12464 ( n9290 , n9259 , n7355 );
    or g12465 ( n10895 , n12768 , n6265 );
    not g12466 ( n3044 , n10102 );
    not g12467 ( n1795 , n7500 );
    and g12468 ( n256 , n2394 , n5096 );
    xnor g12469 ( n12440 , n7403 , n4034 );
    or g12470 ( n35 , n3707 , n5207 );
    or g12471 ( n9605 , n549 , n5 );
    not g12472 ( n1155 , n1910 );
    and g12473 ( n6368 , n10828 , n3346 );
    xnor g12474 ( n11875 , n8302 , n7366 );
    and g12475 ( n8502 , n11493 , n5529 );
    xnor g12476 ( n1090 , n371 , n439 );
    xnor g12477 ( n7671 , n7699 , n874 );
    xor g12478 ( n11397 , n11055 , n139 );
    and g12479 ( n11870 , n8390 , n2076 );
    nor g12480 ( n4181 , n1166 , n5525 );
    or g12481 ( n9625 , n12808 , n8857 );
    or g12482 ( n12674 , n10217 , n6442 );
    and g12483 ( n11851 , n12084 , n13054 );
    xnor g12484 ( n6353 , n1716 , n835 );
    xnor g12485 ( n13054 , n12941 , n1992 );
    or g12486 ( n1626 , n10404 , n3997 );
    nor g12487 ( n6339 , n3388 , n12140 );
    not g12488 ( n9400 , n2252 );
    not g12489 ( n9396 , n4797 );
    and g12490 ( n9833 , n2809 , n9013 );
    not g12491 ( n2487 , n1724 );
    or g12492 ( n11260 , n968 , n2923 );
    and g12493 ( n3037 , n9160 , n2335 );
    not g12494 ( n9618 , n9952 );
    or g12495 ( n7450 , n5313 , n12973 );
    not g12496 ( n8905 , n3644 );
    not g12497 ( n6710 , n4452 );
    or g12498 ( n2132 , n4600 , n1723 );
    or g12499 ( n12918 , n1425 , n11689 );
    and g12500 ( n8347 , n9003 , n1606 );
    nor g12501 ( n11966 , n3427 , n3949 );
    not g12502 ( n8935 , n12553 );
    and g12503 ( n12421 , n3528 , n10918 );
    xnor g12504 ( n9852 , n11206 , n1845 );
    or g12505 ( n11120 , n2538 , n2059 );
    not g12506 ( n11404 , n12482 );
    or g12507 ( n11015 , n4228 , n12684 );
    xnor g12508 ( n8224 , n9860 , n1761 );
    xnor g12509 ( n4195 , n3061 , n13192 );
    xnor g12510 ( n6031 , n12603 , n1910 );
    not g12511 ( n3719 , n12461 );
    not g12512 ( n10005 , n5319 );
    nor g12513 ( n3452 , n11964 , n10766 );
    xnor g12514 ( n1285 , n11736 , n12015 );
    not g12515 ( n10421 , n9915 );
    or g12516 ( n6936 , n3822 , n3339 );
    xnor g12517 ( n369 , n5514 , n7916 );
    xnor g12518 ( n659 , n12690 , n7511 );
    and g12519 ( n4086 , n93 , n10113 );
    and g12520 ( n11581 , n3016 , n7018 );
    not g12521 ( n1989 , n9041 );
    and g12522 ( n7823 , n10794 , n10131 );
    not g12523 ( n4194 , n8230 );
    or g12524 ( n2834 , n10731 , n5485 );
    xnor g12525 ( n1253 , n5475 , n974 );
    xnor g12526 ( n5263 , n347 , n6797 );
    or g12527 ( n12435 , n6970 , n4445 );
    not g12528 ( n2437 , n1055 );
    not g12529 ( n6370 , n9732 );
    and g12530 ( n1530 , n4380 , n10093 );
    and g12531 ( n8639 , n9190 , n3532 );
    or g12532 ( n9398 , n12580 , n4834 );
    xnor g12533 ( n12020 , n4084 , n316 );
    or g12534 ( n12192 , n3281 , n4116 );
    or g12535 ( n1918 , n8926 , n5736 );
    and g12536 ( n5114 , n4371 , n4078 );
    xnor g12537 ( n924 , n7706 , n679 );
    or g12538 ( n6131 , n5271 , n1026 );
    or g12539 ( n11811 , n10274 , n11527 );
    or g12540 ( n3109 , n7872 , n8563 );
    or g12541 ( n3522 , n5482 , n1303 );
    or g12542 ( n7370 , n6106 , n5986 );
    xnor g12543 ( n11299 , n11832 , n4040 );
    or g12544 ( n2407 , n10517 , n11735 );
    or g12545 ( n10428 , n10029 , n8030 );
    or g12546 ( n8687 , n1975 , n6454 );
    xnor g12547 ( n6852 , n2519 , n8591 );
    and g12548 ( n10457 , n2458 , n12306 );
    not g12549 ( n9177 , n10455 );
    or g12550 ( n8973 , n9635 , n3455 );
    not g12551 ( n4107 , n5962 );
    nor g12552 ( n9593 , n11783 , n12079 );
    and g12553 ( n4023 , n4580 , n12844 );
    or g12554 ( n7301 , n9364 , n4300 );
    not g12555 ( n7966 , n4357 );
    or g12556 ( n11376 , n6769 , n177 );
    or g12557 ( n8634 , n5679 , n8030 );
    not g12558 ( n787 , n6818 );
    xnor g12559 ( n12976 , n3375 , n480 );
    xnor g12560 ( n362 , n6930 , n9031 );
    xnor g12561 ( n6083 , n13227 , n2770 );
    or g12562 ( n7891 , n2276 , n5430 );
    and g12563 ( n12767 , n8593 , n565 );
    or g12564 ( n4005 , n6438 , n11668 );
    and g12565 ( n11339 , n1963 , n1008 );
    xnor g12566 ( n2805 , n6831 , n5967 );
    nor g12567 ( n2410 , n3705 , n13177 );
    not g12568 ( n2793 , n102 );
    or g12569 ( n9914 , n7647 , n10387 );
    xnor g12570 ( n12513 , n9807 , n12790 );
    xnor g12571 ( n2343 , n2146 , n9163 );
    xor g12572 ( n1871 , n7792 , n6851 );
    nor g12573 ( n11619 , n1169 , n5620 );
    xnor g12574 ( n2658 , n3696 , n4885 );
    or g12575 ( n782 , n4480 , n10598 );
    or g12576 ( n2086 , n4772 , n12495 );
    or g12577 ( n10618 , n7313 , n2931 );
    xnor g12578 ( n8156 , n577 , n780 );
    or g12579 ( n2914 , n11729 , n7723 );
    and g12580 ( n9074 , n5671 , n5536 );
    xnor g12581 ( n143 , n562 , n6398 );
    and g12582 ( n10493 , n5103 , n3768 );
    xnor g12583 ( n9961 , n12989 , n7143 );
    or g12584 ( n410 , n7205 , n9985 );
    xnor g12585 ( n12515 , n8647 , n4168 );
    not g12586 ( n1625 , n3841 );
    or g12587 ( n8313 , n9931 , n4373 );
    or g12588 ( n1759 , n5679 , n10871 );
    and g12589 ( n4312 , n8139 , n9906 );
    or g12590 ( n7293 , n5261 , n9223 );
    and g12591 ( n832 , n6659 , n9071 );
    xnor g12592 ( n1541 , n2182 , n5278 );
    not g12593 ( n235 , n8742 );
    or g12594 ( n5091 , n13026 , n7961 );
    xnor g12595 ( n5156 , n2598 , n10985 );
    or g12596 ( n10346 , n9843 , n11394 );
    nor g12597 ( n41 , n12771 , n5538 );
    xnor g12598 ( n9036 , n10378 , n4249 );
    or g12599 ( n3024 , n11328 , n3763 );
    xnor g12600 ( n4856 , n10639 , n2921 );
    nor g12601 ( n3027 , n12222 , n4336 );
    xnor g12602 ( n7263 , n9294 , n212 );
    nor g12603 ( n10193 , n4978 , n9821 );
    and g12604 ( n1484 , n10060 , n6866 );
    not g12605 ( n10978 , n9609 );
    or g12606 ( n2049 , n5148 , n4724 );
    xnor g12607 ( n6997 , n3934 , n2414 );
    or g12608 ( n527 , n6245 , n6769 );
    not g12609 ( n13239 , n6487 );
    or g12610 ( n12292 , n1144 , n10871 );
    and g12611 ( n6126 , n8805 , n11648 );
    not g12612 ( n4243 , n2258 );
    xnor g12613 ( n9459 , n870 , n11604 );
    xnor g12614 ( n12797 , n8546 , n1585 );
    xnor g12615 ( n955 , n1599 , n4478 );
    or g12616 ( n6371 , n8757 , n8490 );
    nor g12617 ( n10282 , n518 , n7776 );
    and g12618 ( n139 , n937 , n8506 );
    and g12619 ( n11824 , n4065 , n5251 );
    or g12620 ( n5010 , n12475 , n3759 );
    xnor g12621 ( n831 , n3953 , n796 );
    nor g12622 ( n262 , n6993 , n3506 );
    xnor g12623 ( n3108 , n1067 , n12303 );
    and g12624 ( n7044 , n11061 , n8506 );
    not g12625 ( n6232 , n12255 );
    or g12626 ( n9217 , n10705 , n2561 );
    or g12627 ( n11283 , n97 , n1043 );
    not g12628 ( n12043 , n10091 );
    xnor g12629 ( n12729 , n5158 , n3861 );
    not g12630 ( n11226 , n5884 );
    and g12631 ( n6905 , n8196 , n11269 );
    not g12632 ( n1577 , n2827 );
    nor g12633 ( n9370 , n5062 , n7262 );
    xnor g12634 ( n11939 , n1653 , n10307 );
    xor g12635 ( n109 , n2464 , n8123 );
    or g12636 ( n10533 , n2689 , n10179 );
    not g12637 ( n3858 , n5671 );
    xnor g12638 ( n5675 , n336 , n7290 );
    xnor g12639 ( n12085 , n5738 , n7365 );
    xnor g12640 ( n8281 , n5704 , n10194 );
    not g12641 ( n591 , n140 );
    and g12642 ( n4559 , n4155 , n3437 );
    nor g12643 ( n12714 , n10873 , n8419 );
    xnor g12644 ( n1110 , n5452 , n12307 );
    not g12645 ( n12657 , n1364 );
    or g12646 ( n7295 , n3194 , n4680 );
    xnor g12647 ( n1983 , n7772 , n7529 );
    or g12648 ( n5321 , n4454 , n8268 );
    not g12649 ( n12297 , n11589 );
    or g12650 ( n654 , n1719 , n2686 );
    buf g12651 ( n691 , n11966 );
    and g12652 ( n819 , n10203 , n5234 );
    not g12653 ( n10240 , n5548 );
    xnor g12654 ( n1147 , n983 , n1272 );
    xnor g12655 ( n3073 , n9399 , n11841 );
    nor g12656 ( n10645 , n6168 , n11411 );
    not g12657 ( n2175 , n40 );
    buf g12658 ( n12847 , n11940 );
    and g12659 ( n341 , n52 , n144 );
    and g12660 ( n10708 , n866 , n10428 );
    nor g12661 ( n2804 , n11659 , n12945 );
    nor g12662 ( n6163 , n38 , n7923 );
    xnor g12663 ( n2876 , n2991 , n9440 );
    xnor g12664 ( n791 , n9684 , n12691 );
    xnor g12665 ( n3578 , n5789 , n5437 );
    xnor g12666 ( n11506 , n2982 , n11764 );
    and g12667 ( n12816 , n9773 , n4576 );
    xnor g12668 ( n6115 , n10429 , n252 );
    or g12669 ( n5561 , n542 , n7935 );
    and g12670 ( n12884 , n12897 , n5133 );
    not g12671 ( n9638 , n10642 );
    xnor g12672 ( n11792 , n4188 , n427 );
    and g12673 ( n5357 , n11202 , n1117 );
    xnor g12674 ( n9495 , n5018 , n4477 );
    or g12675 ( n10608 , n10978 , n11008 );
    not g12676 ( n154 , n8820 );
    xnor g12677 ( n3134 , n11303 , n8572 );
    xnor g12678 ( n2846 , n5440 , n2244 );
    xnor g12679 ( n8931 , n2298 , n1757 );
    not g12680 ( n3427 , n854 );
    xnor g12681 ( n7755 , n9769 , n11388 );
    not g12682 ( n3102 , n3863 );
    or g12683 ( n7828 , n7825 , n1144 );
    xnor g12684 ( n11019 , n7759 , n3200 );
    nor g12685 ( n11304 , n10395 , n102 );
    xnor g12686 ( n1860 , n3144 , n9090 );
    or g12687 ( n6803 , n8315 , n12847 );
    xnor g12688 ( n5304 , n4317 , n5405 );
    or g12689 ( n3638 , n5191 , n4070 );
    and g12690 ( n10852 , n10625 , n10160 );
    xnor g12691 ( n10745 , n11215 , n8214 );
    xnor g12692 ( n6365 , n6954 , n1556 );
    not g12693 ( n5462 , n873 );
    not g12694 ( n8122 , n7863 );
    or g12695 ( n6887 , n2329 , n177 );
    xnor g12696 ( n10675 , n6123 , n3420 );
    or g12697 ( n11247 , n2832 , n9943 );
    not g12698 ( n3082 , n1466 );
    xnor g12699 ( n3762 , n9841 , n12219 );
    xnor g12700 ( n3224 , n11178 , n3335 );
    or g12701 ( n6674 , n5158 , n3913 );
    xnor g12702 ( n11687 , n11877 , n10566 );
    and g12703 ( n5977 , n8909 , n3004 );
    or g12704 ( n8109 , n2080 , n13117 );
    xnor g12705 ( n3745 , n3611 , n13155 );
    not g12706 ( n8817 , n7113 );
    xnor g12707 ( n731 , n1424 , n1693 );
    or g12708 ( n13027 , n6416 , n121 );
    xnor g12709 ( n12419 , n11397 , n12903 );
    or g12710 ( n2767 , n4536 , n7430 );
    or g12711 ( n5220 , n8188 , n2738 );
    and g12712 ( n10223 , n1092 , n891 );
    xnor g12713 ( n2753 , n11608 , n4894 );
    nor g12714 ( n8475 , n9211 , n8767 );
    xnor g12715 ( n4671 , n12730 , n328 );
    or g12716 ( n7580 , n11723 , n2222 );
    or g12717 ( n12702 , n12765 , n11447 );
    not g12718 ( n6757 , n6809 );
    xnor g12719 ( n675 , n8779 , n5828 );
    xnor g12720 ( n3670 , n6229 , n6263 );
    and g12721 ( n10932 , n10938 , n1841 );
    xnor g12722 ( n3226 , n11129 , n11052 );
    or g12723 ( n7026 , n6202 , n721 );
    or g12724 ( n10375 , n5016 , n4172 );
    xnor g12725 ( n12862 , n8036 , n12852 );
    xor g12726 ( n4774 , n602 , n10654 );
    or g12727 ( n8074 , n12732 , n121 );
    and g12728 ( n12359 , n12780 , n2413 );
    xnor g12729 ( n3449 , n12078 , n4798 );
    not g12730 ( n10509 , n10142 );
    or g12731 ( n494 , n7819 , n12383 );
    or g12732 ( n7317 , n10195 , n12691 );
    nor g12733 ( n6044 , n6811 , n11364 );
    and g12734 ( n2602 , n8230 , n12289 );
    or g12735 ( n4828 , n10068 , n12173 );
    or g12736 ( n11625 , n6986 , n2059 );
    xnor g12737 ( n9866 , n12341 , n8027 );
    xnor g12738 ( n12506 , n2865 , n3548 );
    xor g12739 ( n8155 , n7541 , n1953 );
    or g12740 ( n2856 , n4890 , n6265 );
    or g12741 ( n10760 , n4412 , n8679 );
    or g12742 ( n10880 , n8802 , n6235 );
    or g12743 ( n5437 , n9501 , n1044 );
    xnor g12744 ( n11812 , n3317 , n7812 );
    or g12745 ( n7401 , n4107 , n11144 );
    nor g12746 ( n8519 , n1610 , n10605 );
    not g12747 ( n7407 , n12746 );
    or g12748 ( n7606 , n10941 , n12746 );
    not g12749 ( n11110 , n6213 );
    xnor g12750 ( n12890 , n12019 , n620 );
    xnor g12751 ( n4895 , n10815 , n8791 );
    xnor g12752 ( n11755 , n6785 , n8691 );
    xnor g12753 ( n11852 , n7711 , n9756 );
    or g12754 ( n7329 , n5328 , n1463 );
    nor g12755 ( n8276 , n3405 , n6752 );
    not g12756 ( n8143 , n9915 );
    buf g12757 ( n6265 , n138 );
    xnor g12758 ( n9504 , n2974 , n788 );
    and g12759 ( n13200 , n6189 , n9092 );
    xnor g12760 ( n12429 , n5384 , n4296 );
    xnor g12761 ( n1260 , n8203 , n315 );
    and g12762 ( n7504 , n1250 , n3113 );
    not g12763 ( n10334 , n8163 );
    and g12764 ( n11685 , n8533 , n2515 );
    or g12765 ( n3216 , n11091 , n12665 );
    or g12766 ( n4466 , n5808 , n3135 );
    xnor g12767 ( n3463 , n9856 , n313 );
    or g12768 ( n5436 , n1747 , n11423 );
    or g12769 ( n11345 , n2738 , n7935 );
    or g12770 ( n6584 , n4937 , n978 );
    nor g12771 ( n1081 , n8647 , n3702 );
    or g12772 ( n11215 , n813 , n1144 );
    xnor g12773 ( n7343 , n8043 , n814 );
    or g12774 ( n5833 , n3509 , n6635 );
    nor g12775 ( n5471 , n7751 , n7093 );
    or g12776 ( n5512 , n12135 , n6714 );
    xnor g12777 ( n2300 , n6747 , n6553 );
    not g12778 ( n198 , n1667 );
    and g12779 ( n6456 , n6428 , n839 );
    and g12780 ( n305 , n3594 , n4632 );
    not g12781 ( n7395 , n10567 );
    xnor g12782 ( n10921 , n5982 , n10827 );
    and g12783 ( n11689 , n7640 , n12697 );
    or g12784 ( n9072 , n5892 , n5942 );
    xnor g12785 ( n2760 , n12462 , n5092 );
    or g12786 ( n5883 , n2734 , n9921 );
    or g12787 ( n11322 , n6837 , n11166 );
    or g12788 ( n6916 , n13227 , n11028 );
    not g12789 ( n13190 , n4357 );
    xnor g12790 ( n10326 , n3725 , n263 );
    not g12791 ( n8050 , n10782 );
    not g12792 ( n4621 , n5920 );
    xnor g12793 ( n4374 , n8433 , n441 );
    xnor g12794 ( n28 , n6624 , n4993 );
    and g12795 ( n10444 , n5100 , n8837 );
    or g12796 ( n11749 , n8053 , n7935 );
    and g12797 ( n420 , n11488 , n12853 );
    or g12798 ( n11705 , n8529 , n7935 );
    xnor g12799 ( n11623 , n11648 , n2627 );
    not g12800 ( n656 , n3713 );
    or g12801 ( n3554 , n12573 , n1463 );
    xnor g12802 ( n7685 , n5404 , n4739 );
    xnor g12803 ( n8497 , n2358 , n2009 );
    or g12804 ( n6018 , n3158 , n12957 );
    or g12805 ( n11957 , n640 , n1808 );
    xnor g12806 ( n12331 , n13208 , n7070 );
    xnor g12807 ( n1063 , n9271 , n3925 );
    or g12808 ( n7404 , n1290 , n9151 );
    or g12809 ( n2769 , n10825 , n6869 );
    xnor g12810 ( n9111 , n9488 , n2114 );
    not g12811 ( n8925 , n209 );
    not g12812 ( n8251 , n9452 );
    not g12813 ( n11218 , n854 );
    xnor g12814 ( n5955 , n12429 , n5815 );
    or g12815 ( n2318 , n4191 , n5074 );
    not g12816 ( n7471 , n6644 );
    or g12817 ( n1938 , n5562 , n9075 );
    and g12818 ( n1038 , n3164 , n8928 );
    xnor g12819 ( n4568 , n4710 , n2313 );
    not g12820 ( n3195 , n4304 );
    not g12821 ( n9280 , n6333 );
    nor g12822 ( n3675 , n11082 , n627 );
    xnor g12823 ( n10791 , n451 , n1680 );
    nor g12824 ( n8806 , n8650 , n13023 );
    nor g12825 ( n4323 , n5203 , n309 );
    or g12826 ( n4217 , n6225 , n12717 );
    nor g12827 ( n2635 , n11363 , n10539 );
    or g12828 ( n371 , n542 , n12388 );
    not g12829 ( n10178 , n11169 );
    or g12830 ( n7087 , n2264 , n5242 );
    not g12831 ( n12088 , n13069 );
    xnor g12832 ( n5325 , n2971 , n6684 );
    or g12833 ( n8405 , n2968 , n4018 );
    and g12834 ( n3919 , n3002 , n11223 );
    or g12835 ( n13049 , n4317 , n11549 );
    nor g12836 ( n4408 , n7364 , n219 );
    xnor g12837 ( n3487 , n4994 , n12305 );
    not g12838 ( n6689 , n3130 );
    xor g12839 ( n1900 , n1484 , n9771 );
    and g12840 ( n6493 , n12597 , n9834 );
    xnor g12841 ( n13057 , n11709 , n3447 );
    and g12842 ( n5457 , n7194 , n7801 );
    nor g12843 ( n8692 , n11577 , n9408 );
    xnor g12844 ( n9640 , n9467 , n13158 );
    or g12845 ( n4356 , n10075 , n7737 );
    or g12846 ( n7679 , n7593 , n2753 );
    and g12847 ( n7954 , n10336 , n6771 );
    xnor g12848 ( n11417 , n7066 , n9156 );
    or g12849 ( n9926 , n9478 , n479 );
    not g12850 ( n7718 , n9475 );
    xnor g12851 ( n1221 , n6864 , n7562 );
    and g12852 ( n13076 , n12098 , n11787 );
    xnor g12853 ( n9246 , n7897 , n889 );
    and g12854 ( n4265 , n3178 , n1007 );
    and g12855 ( n7641 , n1649 , n4263 );
    not g12856 ( n2622 , n5536 );
    not g12857 ( n42 , n3527 );
    nor g12858 ( n8797 , n8908 , n8376 );
    not g12859 ( n7443 , n9839 );
    xnor g12860 ( n7766 , n7380 , n10156 );
    or g12861 ( n5862 , n1888 , n3224 );
    not g12862 ( n8243 , n12809 );
    or g12863 ( n1314 , n11651 , n4505 );
    xnor g12864 ( n9922 , n3659 , n7053 );
    or g12865 ( n6423 , n12496 , n6093 );
    or g12866 ( n2305 , n12266 , n11625 );
    or g12867 ( n151 , n9193 , n12287 );
    xor g12868 ( n2447 , n9358 , n3720 );
    xnor g12869 ( n5421 , n992 , n12319 );
    and g12870 ( n10539 , n12652 , n12699 );
    xnor g12871 ( n10787 , n1326 , n11406 );
    and g12872 ( n11000 , n4784 , n4493 );
    xnor g12873 ( n5288 , n5403 , n9800 );
    not g12874 ( n9889 , n13078 );
    xnor g12875 ( n465 , n2903 , n10922 );
    or g12876 ( n254 , n9926 , n5175 );
    xnor g12877 ( n8422 , n12117 , n12594 );
    or g12878 ( n5892 , n7661 , n4936 );
    or g12879 ( n8464 , n6223 , n10871 );
    xnor g12880 ( n13179 , n5881 , n8281 );
    xnor g12881 ( n483 , n12826 , n5761 );
    xnor g12882 ( n3351 , n1592 , n3850 );
    xnor g12883 ( n6930 , n8230 , n6668 );
    or g12884 ( n1631 , n5541 , n6234 );
    and g12885 ( n1686 , n7871 , n6975 );
    or g12886 ( n5025 , n3564 , n11107 );
    xnor g12887 ( n4009 , n10906 , n9905 );
    or g12888 ( n8307 , n13144 , n6905 );
    xnor g12889 ( n3375 , n10765 , n6662 );
    not g12890 ( n10501 , n7720 );
    or g12891 ( n344 , n2877 , n12388 );
    not g12892 ( n4030 , n1288 );
    not g12893 ( n5638 , n4671 );
    xnor g12894 ( n261 , n9222 , n1348 );
    or g12895 ( n9015 , n1262 , n2986 );
    xnor g12896 ( n7376 , n6611 , n3605 );
    not g12897 ( n2838 , n4186 );
    or g12898 ( n3164 , n1872 , n11995 );
    or g12899 ( n4216 , n1480 , n902 );
    not g12900 ( n13017 , n12228 );
    nor g12901 ( n13136 , n2749 , n10515 );
    or g12902 ( n11378 , n1930 , n8268 );
    xnor g12903 ( n13188 , n5428 , n9774 );
    xnor g12904 ( n33 , n6395 , n7148 );
    not g12905 ( n6330 , n11544 );
    not g12906 ( n1080 , n9918 );
    or g12907 ( n12063 , n137 , n4636 );
    xnor g12908 ( n3711 , n503 , n9820 );
    not g12909 ( n2623 , n3178 );
    nor g12910 ( n7796 , n1033 , n4127 );
    nor g12911 ( n7136 , n3993 , n2007 );
    or g12912 ( n5164 , n2657 , n3949 );
    and g12913 ( n5197 , n4484 , n11540 );
    xor g12914 ( n211 , n10680 , n4121 );
    not g12915 ( n1135 , n9041 );
    not g12916 ( n2217 , n1231 );
    nor g12917 ( n11456 , n4954 , n8162 );
    xnor g12918 ( n3170 , n10855 , n3547 );
    xnor g12919 ( n10568 , n668 , n2543 );
    or g12920 ( n518 , n3908 , n4640 );
    not g12921 ( n7062 , n7374 );
    or g12922 ( n8764 , n5660 , n2319 );
    not g12923 ( n5279 , n7514 );
    xnor g12924 ( n9127 , n8060 , n10169 );
    or g12925 ( n11386 , n8729 , n4640 );
    or g12926 ( n2823 , n11941 , n2133 );
    or g12927 ( n3360 , n10383 , n4724 );
    xnor g12928 ( n291 , n7105 , n13009 );
    or g12929 ( n12353 , n7718 , n4947 );
    xnor g12930 ( n9449 , n11289 , n13114 );
    or g12931 ( n12288 , n9496 , n8034 );
    xnor g12932 ( n11694 , n6965 , n2488 );
    xnor g12933 ( n9774 , n1828 , n4403 );
    nor g12934 ( n10115 , n2643 , n4629 );
    and g12935 ( n6902 , n3035 , n8590 );
    or g12936 ( n10490 , n9131 , n1144 );
    xor g12937 ( n4188 , n9849 , n11866 );
    xnor g12938 ( n9844 , n7594 , n7512 );
    not g12939 ( n6245 , n4419 );
    xnor g12940 ( n3838 , n4291 , n2256 );
    not g12941 ( n333 , n11488 );
    xnor g12942 ( n6862 , n12051 , n7663 );
    or g12943 ( n11463 , n12293 , n2044 );
    or g12944 ( n13140 , n4339 , n170 );
    xnor g12945 ( n4273 , n3535 , n393 );
    and g12946 ( n11905 , n8385 , n12431 );
    xnor g12947 ( n184 , n13197 , n8945 );
    xnor g12948 ( n7288 , n3933 , n10669 );
    or g12949 ( n8048 , n2657 , n3149 );
    not g12950 ( n6041 , n11537 );
    not g12951 ( n7675 , n7411 );
    not g12952 ( n12717 , n2590 );
    xnor g12953 ( n3015 , n11744 , n4235 );
    or g12954 ( n4822 , n8113 , n7032 );
    or g12955 ( n12392 , n12441 , n6814 );
    or g12956 ( n8741 , n8420 , n1866 );
    xnor g12957 ( n12084 , n11508 , n6623 );
    xnor g12958 ( n12091 , n7829 , n5532 );
    xnor g12959 ( n3735 , n781 , n4582 );
    not g12960 ( n8569 , n1757 );
    nor g12961 ( n6208 , n9243 , n2245 );
    xnor g12962 ( n3754 , n12484 , n1957 );
    xnor g12963 ( n4867 , n5539 , n12444 );
    xnor g12964 ( n3072 , n3389 , n9374 );
    and g12965 ( n11097 , n4835 , n12236 );
    xnor g12966 ( n12269 , n4396 , n8612 );
    and g12967 ( n1949 , n4754 , n3533 );
    or g12968 ( n7566 , n8561 , n10871 );
    or g12969 ( n8899 , n13130 , n8828 );
    or g12970 ( n3120 , n8158 , n11719 );
    not g12971 ( n4517 , n10113 );
    xnor g12972 ( n10702 , n968 , n2923 );
    and g12973 ( n3900 , n2892 , n108 );
    not g12974 ( n8985 , n160 );
    not g12975 ( n10890 , n9324 );
    and g12976 ( n10873 , n13122 , n11813 );
    or g12977 ( n6501 , n7327 , n11841 );
    not g12978 ( n8669 , n3187 );
    or g12979 ( n8257 , n10313 , n1782 );
    xnor g12980 ( n5591 , n2750 , n8824 );
    xnor g12981 ( n5576 , n2238 , n12248 );
    not g12982 ( n3712 , n3973 );
    and g12983 ( n10483 , n5527 , n3831 );
    and g12984 ( n8102 , n10668 , n5141 );
    or g12985 ( n1596 , n7427 , n7534 );
    and g12986 ( n11925 , n7159 , n4928 );
    not g12987 ( n8744 , n8139 );
    xnor g12988 ( n8966 , n2534 , n11467 );
    and g12989 ( n9715 , n10891 , n5653 );
    and g12990 ( n10967 , n7960 , n12819 );
    and g12991 ( n3920 , n8845 , n7414 );
    nor g12992 ( n9200 , n9967 , n1442 );
    nor g12993 ( n10226 , n7937 , n7721 );
    not g12994 ( n5527 , n912 );
    not g12995 ( n8175 , n6083 );
    or g12996 ( n5323 , n5713 , n10029 );
    not g12997 ( n5310 , n13047 );
    xnor g12998 ( n7178 , n9701 , n7009 );
    or g12999 ( n12868 , n5044 , n12860 );
    and g13000 ( n2510 , n3493 , n1085 );
    not g13001 ( n2294 , n3005 );
    not g13002 ( n12858 , n4350 );
endmodule
