module top( n2 , n11 , n13 , n16 , n21 , n44 , n45 , n46 , n55 , n74 , n75 , n81 , n84 , n85 , n87 , n93 , n96 , n98 , n101 , n105 , n111 , n123 , n128 , n131 , n134 , n139 , n148 , n153 , n159 , n163 , n177 , n191 , n196 , n199 , n206 , n211 , n216 , n223 , n226 , n240 , n243 , n254 , n260 , n264 , n266 , n280 , n282 , n283 , n287 , n290 , n291 , n299 , n309 , n336 , n346 , n349 , n360 , n368 , n369 , n377 , n388 , n394 , n409 , n428 , n435 , n442 , n447 , n449 , n454 , n457 , n468 , n471 , n481 , n484 , n494 , n500 , n507 , n511 , n518 , n519 , n525 , n534 , n542 , n547 , n557 , n561 , n568 , n569 , n571 , n575 , n581 , n582 , n583 , n587 , n600 , n603 , n609 , n613 , n614 , n616 , n627 , n635 , n646 , n659 , n661 , n664 , n672 , n673 );
    input n2 , n11 , n13 , n16 , n21 , n45 , n46 , n55 , n74 , n75 , n81 , n84 , n85 , n93 , n96 , n98 , n101 , n111 , n128 , n131 , n134 , n139 , n153 , n159 , n177 , n199 , n206 , n211 , n216 , n223 , n243 , n264 , n266 , n280 , n282 , n287 , n290 , n309 , n336 , n346 , n349 , n360 , n368 , n369 , n377 , n388 , n394 , n409 , n428 , n435 , n447 , n454 , n457 , n468 , n471 , n481 , n494 , n500 , n507 , n511 , n519 , n525 , n557 , n561 , n569 , n571 , n575 , n581 , n582 , n583 , n587 , n600 , n603 , n609 , n613 , n614 , n616 , n646 , n659 , n661 , n664 , n673 ;
    output n44 , n87 , n105 , n123 , n148 , n163 , n191 , n196 , n226 , n240 , n254 , n260 , n283 , n291 , n299 , n442 , n449 , n484 , n518 , n534 , n542 , n547 , n568 , n627 , n635 , n672 ;
    wire n0 , n1 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , n12 , n14 , n15 , n17 , n18 , n19 , n20 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n76 , n77 , n78 , n79 , n80 , n82 , n83 , n86 , n88 , n89 , n90 , n91 , n92 , n94 , n95 , n97 , n99 , n100 , n102 , n103 , n104 , n106 , n107 , n108 , n109 , n110 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n124 , n125 , n126 , n127 , n129 , n130 , n132 , n133 , n135 , n136 , n137 , n138 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n149 , n150 , n151 , n152 , n154 , n155 , n156 , n157 , n158 , n160 , n161 , n162 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n192 , n193 , n194 , n195 , n197 , n198 , n200 , n201 , n202 , n203 , n204 , n205 , n207 , n208 , n209 , n210 , n212 , n213 , n214 , n215 , n217 , n218 , n219 , n220 , n221 , n222 , n224 , n225 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n241 , n242 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n255 , n256 , n257 , n258 , n259 , n261 , n262 , n263 , n265 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n281 , n284 , n285 , n286 , n288 , n289 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n347 , n348 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n389 , n390 , n391 , n392 , n393 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n429 , n430 , n431 , n432 , n433 , n434 , n436 , n437 , n438 , n439 , n440 , n441 , n443 , n444 , n445 , n446 , n448 , n450 , n451 , n452 , n453 , n455 , n456 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n469 , n470 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n482 , n483 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n495 , n496 , n497 , n498 , n499 , n501 , n502 , n503 , n504 , n505 , n506 , n508 , n509 , n510 , n512 , n513 , n514 , n515 , n516 , n517 , n520 , n521 , n522 , n523 , n524 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n543 , n544 , n545 , n546 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n558 , n559 , n560 , n562 , n563 , n564 , n565 , n566 , n567 , n570 , n572 , n573 , n574 , n576 , n577 , n578 , n579 , n580 , n584 , n585 , n586 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n601 , n602 , n604 , n605 , n606 , n607 , n608 , n610 , n611 , n612 , n615 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n660 , n662 , n663 , n665 , n666 , n667 , n668 , n669 , n670 , n671 ;
assign n657 = n356 & n451;
assign n203 = n224 & n349;
assign n660 = n340 & n25;
assign n347 = ~(n468 | n417);
assign n253 = ~n54;
assign n6 = n48 | n383;
assign n291 = ~(n339 ^ n668);
assign n308 = n515 & n168;
assign n629 = n253 | n652;
assign n187 = ~(n2 | n159);
assign n585 = ~n434;
assign n570 = n389;
assign n47 = ~(n414 | n467);
assign n393 = ~(n444 ^ n216);
assign n391 = ~n531;
assign n443 = ~n176;
assign n76 = ~(n556 ^ n16);
assign n390 = ~(n598 ^ n290);
assign n38 = ~n499;
assign n426 = n524 | n62;
assign n117 = ~(n93 | n396);
assign n89 = n9 & n72;
assign n628 = ~(n107 ^ n531);
assign n550 = ~n159;
assign n365 = n321 & n253;
assign n163 = ~(n0 ^ n479);
assign n61 = ~(n7 ^ n613);
assign n648 = n127 & n125;
assign n283 = ~(n31 ^ n648);
assign n608 = ~n31;
assign n327 = n638 & n367;
assign n444 = n285 | n412;
assign n373 = ~n639;
assign n602 = n570 & n101;
assign n251 = ~n75;
assign n107 = ~n520;
assign n427 = n608 | n125;
assign n480 = ~(n349 | n322);
assign n359 = n137 & n604;
assign n95 = ~(n13 | n2);
assign n118 = ~(n623 | n540);
assign n474 = ~n613;
assign n115 = ~(n93 | n37);
assign n398 = ~n0;
assign n289 = ~(n280 ^ n287);
assign n543 = n390 & n266;
assign n60 = ~(n624 ^ n464);
assign n141 = n538 | n452;
assign n572 = ~n466;
assign n339 = n5 | n492;
assign n31 = n559 | n424;
assign n514 = ~n206;
assign n234 = n198 & n326;
assign n258 = n19 & n266;
assign n300 = ~n428;
assign n651 = n526 & n570;
assign n197 = ~n138;
assign n351 = ~n508;
assign n649 = ~n225;
assign n100 = n413 | n179;
assign n670 = ~(n203 | n611);
assign n30 = n318 | n342;
assign n144 = n385 | n445;
assign n453 = n539 | n344;
assign n78 = ~n365;
assign n496 = n233 & n93;
assign n179 = ~(n570 | n330);
assign n39 = ~(n490 | n480);
assign n149 = ~n144;
assign n182 = ~(n183 | n370);
assign n9 = n513 & n551;
assign n152 = ~(n356 ^ n616);
assign n576 = ~n100;
assign n662 = n580 & n264;
assign n123 = ~(n182 ^ n463);
assign n65 = n201 | n439;
assign n259 = n58 | n1;
assign n591 = ~(n590 | n275);
assign n200 = n136 & n266;
assign n399 = ~n573;
assign n558 = n64 | n453;
assign n434 = n450 | n86;
assign n618 = n537 | n18;
assign n140 = n333 & n654;
assign n553 = ~(n6 ^ n432);
assign n34 = n375 | n116;
assign n5 = n570 & n500;
assign n530 = ~(n472 | n327);
assign n626 = n384 | n642;
assign n401 = ~(n582 ^ n2);
assign n450 = n190 | n307;
assign n106 = n465 & n608;
assign n40 = n421 & n93;
assign n520 = ~n248;
assign n299 = ~(n395 ^ n175);
assign n501 = ~n171;
assign n420 = ~n45;
assign n169 = n319 | n629;
assign n637 = n124 & n335;
assign n621 = ~n380;
assign n267 = ~(n570 | n140);
assign n105 = ~(n54 ^ n615);
assign n533 = n331 | n52;
assign n355 = n71 | n591;
assign n260 = ~(n508 ^ n669);
assign n594 = n514 | n516;
assign n395 = ~(n431 | n663);
assign n302 = ~(n453 ^ n336);
assign n363 = n526 | n239;
assign n238 = n42 & n93;
assign n424 = n61 & n266;
assign n567 = n77 & n569;
assign n79 = n29 & n266;
assign n598 = n298 | n460;
assign n620 = ~(n632 ^ n392);
assign n479 = ~(n185 | n425);
assign n143 = ~n339;
assign n77 = n389;
assign n624 = n285 | n305;
assign n218 = n249 & n266;
assign n3 = n147 & n266;
assign n88 = ~(n199 | n85);
assign n249 = ~(n426 ^ n282);
assign n380 = n358 | n597;
assign n654 = n58 | n562;
assign n165 = n201 | n660;
assign n212 = ~(n75 | n131);
assign n623 = ~n577;
assign n7 = n636 | n477;
assign n340 = ~(n170 | n418);
assign n114 = n482 | n444;
assign n560 = ~n209;
assign n580 = n666 & n43;
assign n274 = n570 & n603;
assign n1 = ~n381;
assign n484 = ~(n180 ^ n584);
assign n592 = n606 | n503;
assign n222 = n26 & n436;
assign n335 = n397 | n517;
assign n461 = ~n13;
assign n650 = ~(n665 | n15);
assign n552 = n220 | n461;
assign n475 = n227 | n637;
assign n386 = n231 | n323;
assign n130 = n440 | n548;
assign n312 = ~(n77 | n637);
assign n463 = n566 | n543;
assign n497 = n538 | n278;
assign n655 = n470 | n324;
assign n257 = n387 | n200;
assign n110 = n65 & n601;
assign n478 = n570 & n153;
assign n90 = n653 | n459;
assign n658 = n302 & n266;
assign n262 = ~(n177 ^ n75);
assign n155 = ~n521;
assign n383 = ~n468;
assign n167 = n359 | n219;
assign n15 = ~n373;
assign n247 = n662 | n404;
assign n640 = n284 & n552;
assign n201 = ~n352;
assign n415 = ~(n194 | n133);
assign n367 = n625 | n209;
assign n635 = ~(n12 ^ n4);
assign n207 = ~n641;
assign n344 = n429 | n353;
assign n192 = ~(n34 | n517);
assign n189 = n235 & n487;
assign n261 = n428 | n48;
assign n389 = ~n266;
assign n148 = ~(n36 ^ n17);
assign n372 = n57 & n266;
assign n579 = n586 | n78;
assign n374 = n393 & n206;
assign n124 = n334 | n140;
assign n174 = ~n51;
assign n4 = n434 & n52;
assign n588 = ~n388;
assign n269 = n564 & n126;
assign n156 = n63 | n495;
assign n286 = n455 & n482;
assign n161 = ~(n657 | n438);
assign n483 = ~n6;
assign n509 = ~n368;
assign n541 = ~(n472 | n39);
assign n43 = ~n93;
assign n64 = ~n336;
assign n284 = n95 | n294;
assign n328 = ~n631;
assign n464 = ~(n511 ^ n454);
assign n433 = n158 & n441;
assign n563 = ~n511;
assign n71 = n2 & n582;
assign n67 = n94 & n35;
assign n456 = n251 | n8;
assign n217 = ~(n135 | n419);
assign n448 = ~n595;
assign n310 = ~n533;
assign n265 = ~(n289 | n316);
assign n151 = n286 | n408;
assign n281 = n221 | n593;
assign n568 = ~(n217 ^ n406);
assign n644 = n570 & n614;
assign n73 = ~n450;
assign n154 = ~(n459 ^ n583);
assign n532 = n475 & n167;
assign n607 = ~(n355 ^ n97);
assign n256 = n553 & n93;
assign n150 = n570 & n519;
assign n304 = ~(n107 | n219);
assign n80 = ~n352;
assign n667 = n639 & n174;
assign n248 = ~n359;
assign n87 = ~(n156 ^ n49);
assign n168 = n359 | n271;
assign n403 = n451 | n295;
assign n324 = ~n560;
assign n593 = n546 & n527;
assign n215 = ~n235;
assign n32 = n659 & n93;
assign n458 = ~(n294 ^ n112);
assign n513 = n187 | n632;
assign n467 = n206 | n509;
assign n385 = n237 | n129;
assign n72 = n251 | n121;
assign n517 = ~n197;
assign n8 = ~n177;
assign n482 = ~n216;
assign n337 = ~(n443 | n269);
assign n476 = n650 | n50;
assign n638 = ~(n229 | n265);
assign n319 = ~n586;
assign n157 = n212 | n89;
assign n240 = ~(n341 ^ n402);
assign n24 = ~n491;
assign n295 = n493 | n114;
assign n627 = ~(n130 ^ n366);
assign n625 = ~n664;
assign n178 = n616 | n66;
assign n642 = n505 | n90;
assign n311 = n228 | n363;
assign n33 = ~(n620 | n623);
assign n18 = ~(n77 | n60);
assign n171 = n351 | n169;
assign n341 = n343 | n345;
assign n68 = n570 & n581;
assign n556 = n102 | n329;
assign n437 = ~(n119 | n293);
assign n606 = ~n646;
assign n565 = ~n624;
assign n412 = ~n454;
assign n473 = ~n432;
assign n462 = ~n381;
assign n503 = n315 | n426;
assign n48 = ~n409;
assign n285 = ~n659;
assign n27 = ~(n119 | n356);
assign n263 = ~(n626 ^ n388);
assign n430 = ~n579;
assign n112 = ~(n13 ^ n2);
assign n536 = ~n561;
assign n527 = n478 | n574;
assign n358 = ~(n20 | n43);
assign n632 = n276 | n120;
assign n505 = ~n55;
assign n313 = n386 & n259;
assign n104 = n511 | n659;
assign n296 = ~(n435 | n75);
assign n146 = n454 & n511;
assign n307 = n272 & n266;
assign n321 = ~n656;
assign n554 = ~n555;
assign n276 = ~n287;
assign n442 = ~(n172 ^ n382);
assign n619 = ~(n6 | n473);
assign n396 = n165 & n522;
assign n566 = n77 & n74;
assign n22 = ~n425;
assign n120 = ~n96;
assign n323 = ~(n306 | n562);
assign n224 = n275 ^ n401;
assign n315 = ~n282;
assign n23 = n596 & n155;
assign n172 = n274 | n325;
assign n306 = ~n576;
assign n241 = n506 | n592;
assign n528 = n405 | n427;
assign n63 = n570 & n139;
assign n183 = n242 & n555;
assign n378 = ~(n292 | n193);
assign n20 = ~(n428 ^ n454);
assign n666 = ~(n80 | n209);
assign n669 = n579 & n169;
assign n353 = n634 | n612;
assign n126 = ~n350;
assign n548 = n622 & n266;
assign n42 = ~(n10 ^ n202);
assign n508 = n166 | n258;
assign n488 = n279 & n77;
assign n498 = ~(n423 ^ n45);
assign n116 = ~(n77 | n76);
assign n489 = n437 | n10;
assign n37 = n273 & n594;
assign n510 = ~n211;
assign n278 = ~n38;
assign n460 = n230 | n558;
assign n226 = ~(n213 ^ n245);
assign n397 = ~n448;
assign n559 = n77 & n609;
assign n371 = n77 & n11;
assign n405 = ~n172;
assign n555 = n486 | n647;
assign n268 = ~n629;
assign n589 = n106 & n405;
assign n205 = n422 | n241;
assign n665 = ~n51;
assign n421 = ~(n455 ^ n103);
assign n186 = n580 & n21;
assign n417 = n409 & n428;
assign n209 = n85 | n349;
assign n293 = ~(n261 ^ n468);
assign n516 = ~(n214 ^ n114);
assign n135 = n231 & n77;
assign n518 = ~(n555 ^ n195);
assign n633 = n624 & n104;
assign n438 = n489 & n178;
assign n663 = ~(n570 | n532);
assign n12 = n602 | n3;
assign n82 = ~(n160 | n312);
assign n504 = ~(n296 | n91);
assign n250 = ~(n177 | n75);
assign n384 = ~n128;
assign n142 = n236 & n497;
assign n599 = ~n216;
assign n645 = n59 | n228;
assign n436 = n485 | n23;
assign n564 = ~n132;
assign n162 = ~(n514 | n643);
assign n108 = n210 & n85;
assign n173 = n317 & n266;
assign n596 = n32 | n332;
assign n50 = ~(n667 | n532);
assign n230 = ~n494;
assign n305 = ~n511;
assign n298 = ~n223;
assign n350 = n68 | n529;
assign n160 = n67 & n77;
assign n326 = n599 | n305;
assign n366 = n144 & n184;
assign n485 = ~n618;
assign n577 = ~n467;
assign n109 = ~n527;
assign n522 = ~(n374 | n118);
assign n615 = n656 & n652;
assign n537 = n77 & n46;
assign n431 = n308 & n570;
assign n254 = n411 | n281;
assign n597 = ~(n93 | n110);
assign n147 = ~(n344 ^ n369);
assign n499 = n40 | n117;
assign n121 = ~n131;
assign n601 = ~(n33 | n162);
assign n127 = ~n465;
assign n26 = n380 | n354;
assign n17 = ~(n448 ^ n138);
assign n231 = n181 & n141;
assign n198 = ~n288;
assign n387 = n570 & n457;
assign n653 = ~n583;
assign n590 = ~(n582 | n2);
assign n361 = n28 & n53;
assign n136 = ~(n288 ^ n113);
assign n652 = n266 | n415;
assign n531 = n186 | n256;
assign n166 = n570 & n571;
assign n610 = ~n138;
assign n297 = n498 & n266;
assign n94 = n192 | n313;
assign n145 = ~n130;
assign n193 = n47 | n530;
assign n232 = ~n377;
assign n342 = n145 | n184;
assign n138 = n247 | n496;
assign n470 = ~n525;
assign n213 = ~(n488 | n362);
assign n325 = n154 & n266;
assign n382 = n446 & n427;
assign n429 = ~n575;
assign n538 = ~n207;
assign n449 = ~(n155 ^ n596);
assign n418 = n607 & n349;
assign n176 = n126 | n30;
assign n605 = n570 & n84;
assign n70 = n143 | n171;
assign n370 = n411 & n554;
assign n86 = ~n269;
assign n119 = ~n616;
assign n273 = ~(n502 | n541);
assign n441 = ~n239;
assign n316 = n349 | n92;
assign n630 = n149 & n145;
assign n294 = n276 | n545;
assign n318 = ~n341;
assign n219 = ~n391;
assign n604 = n266 | n232;
assign n402 = ~(n416 | n630);
assign n672 = ~(n385 ^ n400);
assign n208 = ~n528;
assign n272 = ~(n353 ^ n575);
assign n320 = ~n600;
assign n376 = ~(n511 ^ n616);
assign n52 = n73 | n176;
assign n314 = ~n109;
assign n92 = ~n85;
assign n611 = ~(n458 | n316);
assign n181 = n122 | n279;
assign n53 = ~n180;
assign n338 = n75 & n435;
assign n245 = ~(n207 ^ n499);
assign n244 = ~(n558 ^ n494);
assign n521 = ~n526;
assign n14 = ~n23;
assign n540 = ~(n9 ^ n164);
assign n574 = n244 & n266;
assign n303 = n77 & n346;
assign n132 = n341 | n56;
assign n422 = ~n557;
assign n529 = n469 & n266;
assign n671 = n313 & n77;
assign n419 = ~(n77 | n142);
assign n354 = ~(n618 | n14);
assign n255 = n563 | n348;
assign n221 = ~(n527 | n225);
assign n54 = n605 | n79;
assign n102 = ~(n563 | n214);
assign n25 = n510 | n324;
assign n204 = ~(n257 | n452);
assign n362 = ~(n570 | n222);
assign n636 = ~n471;
assign n252 = n599 | n455;
assign n356 = n483 | n347;
assign n524 = ~n111;
assign n413 = n77 & n507;
assign n292 = ~(n659 | n493);
assign n357 = ~(n241 ^ n557);
assign n133 = ~(n99 | n308);
assign n647 = n410 & n266;
assign n639 = n277 | n549;
assign n495 = n357 & n266;
assign n36 = ~(n671 | n267);
assign n329 = ~n234;
assign n35 = n397 | n610;
assign n526 = n24 & n270;
assign n0 = n303 | n173;
assign n379 = ~n156;
assign n586 = n371 | n218;
assign n28 = n585 & n331;
assign n57 = ~(n477 ^ n471);
assign n472 = n368 | n206;
assign n180 = n567 | n658;
assign n535 = ~(n90 ^ n55);
assign n656 = n77 | n476;
assign n91 = ~(n338 | n355);
assign n44 = ~(n466 ^ n189);
assign n41 = ~n16;
assign n381 = n238 | n115;
assign n56 = ~n630;
assign n451 = ~n616;
assign n99 = n373 & n174;
assign n348 = ~n423;
assign n322 = n88 | n108;
assign n233 = ~(n438 ^ n152);
assign n220 = ~n2;
assign n506 = ~n243;
assign n235 = n0 | n22;
assign n184 = n69 | n528;
assign n539 = ~n369;
assign n270 = n266 | n83;
assign n551 = n220 | n550;
assign n188 = ~(n268 | n365);
assign n465 = n215 & n572;
assign n410 = ~(n460 ^ n223);
assign n195 = ~(n242 | n411);
assign n122 = ~(n257 | n278);
assign n288 = n146 | n565;
assign n408 = ~(n428 ^ n409);
assign n49 = n573 & n70;
assign n578 = n640 & n456;
assign n547 = ~(n82 ^ n628);
assign n493 = ~n206;
assign n331 = ~n12;
assign n400 = ~(n208 | n589);
assign n66 = ~n293;
assign n51 = n150 | n297;
assign n631 = n430 & n351;
assign n214 = ~n616;
assign n236 = n204 | n222;
assign n343 = n77 & n360;
assign n668 = ~(n501 | n631);
assign n137 = n77 | n255;
assign n406 = ~(n306 ^ n381);
assign n185 = ~n544;
assign n641 = ~n257;
assign n62 = n420 | n423;
assign n246 = ~(n640 ^ n262);
assign n229 = n364 & n349;
assign n59 = n491 | n651;
assign n271 = ~n531;
assign n227 = ~(n248 | n271);
assign n158 = n407 | n621;
assign n242 = n649 & n314;
assign n277 = n580 & n98;
assign n29 = ~(n62 ^ n111);
assign n190 = n570 & n134;
assign n491 = n633 & n266;
assign n549 = n619 & n93;
assign n634 = ~n661;
assign n333 = n617 | n142;
assign n202 = ~(n293 ^ n616);
assign n196 = ~(n645 ^ n433);
assign n58 = ~n100;
assign n459 = n474 | n7;
assign n364 = n600 ^ n287;
assign n622 = ~(n642 ^ n128);
assign n643 = ~(n659 ^ n454);
assign n486 = n77 & n309;
assign n515 = n304 | n67;
assign n414 = ~(n287 ^ n96);
assign n194 = n15 & n51;
assign n490 = n504 & n349;
assign n584 = ~(n310 | n28);
assign n446 = ~n106;
assign n191 = ~(n350 ^ n523);
assign n125 = n572 | n487;
assign n103 = ~(n408 ^ n216);
assign n469 = ~(n612 ^ n661);
assign n228 = ~n596;
assign n332 = ~(n93 | n378);
assign n502 = ~(n467 | n157);
assign n10 = n151 & n252;
assign n512 = ~n556;
assign n237 = n570 & n447;
assign n573 = n339 | n328;
assign n164 = ~(n75 ^ n131);
assign n69 = ~n385;
assign n225 = n53 | n533;
assign n239 = n621 & n407;
assign n466 = n644 | n372;
assign n407 = ~n618;
assign n523 = n132 & n30;
assign n175 = n99 | n194;
assign n440 = n570 & n394;
assign n544 = n379 | n70;
assign n487 = n398 | n544;
assign n545 = ~n280;
assign n534 = ~(n586 ^ n188);
assign n210 = n250 | n578;
assign n542 = ~(n450 ^ n337);
assign n279 = n311 & n158;
assign n275 = n276 | n320;
assign n330 = ~(n234 ^ n376);
assign n416 = ~n342;
assign n546 = ~(n649 | n361);
assign n477 = n536 | n205;
assign n411 = n361 & n109;
assign n352 = ~n472;
assign n612 = n588 | n626;
assign n452 = ~n499;
assign n423 = n41 | n512;
assign n375 = n77 & n81;
assign n492 = n301 & n266;
assign n392 = ~(n2 ^ n159);
assign n129 = n535 & n266;
assign n562 = ~n462;
assign n334 = ~(n34 | n610);
assign n113 = ~(n511 ^ n216);
assign n439 = n670 & n655;
assign n455 = n300 | n412;
assign n345 = n263 & n266;
assign n617 = ~(n100 | n1);
assign n97 = ~(n435 ^ n75);
assign n425 = n399 & n379;
assign n432 = n27 | n161;
assign n301 = ~(n592 ^ n243);
assign n445 = ~n589;
assign n317 = ~(n205 ^ n561);
assign n19 = ~(n503 ^ n646);
assign n595 = ~n34;
assign n404 = ~(n93 | n403);
assign n170 = ~(n316 | n246);
assign n83 = ~n673;
endmodule
