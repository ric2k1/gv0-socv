module top( n1 , n3 , n4 , n15 , n21 , n23 , n28 , n32 , n37 , 
n38 , n40 , n45 , n47 , n50 , n52 , n53 , n54 , n60 , n72 , 
n75 , n79 , n81 , n83 , n86 , n87 , n91 , n95 , n97 , n99 , 
n105 , n111 , n114 , n117 , n122 , n139 , n152 , n154 , n155 , n160 , 
n162 , n168 , n176 , n183 , n185 , n187 , n191 , n194 , n197 , n198 , 
n200 , n205 , n206 , n208 , n211 , n214 , n215 , n218 , n220 , n227 , 
n228 , n231 , n242 , n243 , n248 , n254 , n262 , n265 , n269 , n273 , 
n276 , n278 , n280 , n283 );
    input n1 , n4 , n15 , n21 , n23 , n28 , n37 , n38 , n45 , 
n52 , n53 , n60 , n75 , n79 , n83 , n87 , n95 , n105 , n114 , 
n117 , n122 , n152 , n155 , n160 , n162 , n168 , n183 , n187 , n194 , 
n198 , n206 , n215 , n218 , n227 , n228 , n231 , n242 , n269 , n276 , 
n278 , n280 ;
    output n3 , n32 , n40 , n47 , n50 , n54 , n72 , n81 , n86 , 
n91 , n97 , n99 , n111 , n139 , n154 , n176 , n185 , n191 , n197 , 
n200 , n205 , n208 , n211 , n214 , n220 , n243 , n248 , n254 , n262 , 
n265 , n273 , n283 ;
    wire n0 , n2 , n5 , n6 , n7 , n8 , n9 , n10 , n11 , 
n12 , n13 , n14 , n16 , n17 , n18 , n19 , n20 , n22 , n24 , 
n25 , n26 , n27 , n29 , n30 , n31 , n33 , n34 , n35 , n36 , 
n39 , n41 , n42 , n43 , n44 , n46 , n48 , n49 , n51 , n55 , 
n56 , n57 , n58 , n59 , n61 , n62 , n63 , n64 , n65 , n66 , 
n67 , n68 , n69 , n70 , n71 , n73 , n74 , n76 , n77 , n78 , 
n80 , n82 , n84 , n85 , n88 , n89 , n90 , n92 , n93 , n94 , 
n96 , n98 , n100 , n101 , n102 , n103 , n104 , n106 , n107 , n108 , 
n109 , n110 , n112 , n113 , n115 , n116 , n118 , n119 , n120 , n121 , 
n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , 
n133 , n134 , n135 , n136 , n137 , n138 , n140 , n141 , n142 , n143 , 
n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n153 , n156 , 
n157 , n158 , n159 , n161 , n163 , n164 , n165 , n166 , n167 , n169 , 
n170 , n171 , n172 , n173 , n174 , n175 , n177 , n178 , n179 , n180 , 
n181 , n182 , n184 , n186 , n188 , n189 , n190 , n192 , n193 , n195 , 
n196 , n199 , n201 , n202 , n203 , n204 , n207 , n209 , n210 , n212 , 
n213 , n216 , n217 , n219 , n221 , n222 , n223 , n224 , n225 , n226 , 
n229 , n230 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , 
n240 , n241 , n244 , n245 , n246 , n247 , n249 , n250 , n251 , n252 , 
n253 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n263 , n264 , 
n266 , n267 , n268 , n270 , n271 , n272 , n274 , n275 , n277 , n279 , 
n281 , n282 , n284 , n285 ;
    and g0 ( n140 , n247 , n201 );
    xnor g1 ( n72 , n126 , n162 );
    or g2 ( n244 , n173 , n230 );
    or g3 ( n18 , n141 , n136 );
    not g4 ( n43 , n4 );
    not g5 ( n177 , n198 );
    xnor g6 ( n16 , n215 , n206 );
    or g7 ( n80 , n237 , n252 );
    xnor g8 ( n81 , n216 , n194 );
    not g9 ( n261 , n193 );
    not g10 ( n55 , n172 );
    not g11 ( n148 , n168 );
    xnor g12 ( n136 , n209 , n77 );
    xnor g13 ( n263 , n206 , n183 );
    xnor g14 ( n257 , n280 , n21 );
    xnor g15 ( n159 , n285 , n24 );
    xor g16 ( n254 , n0 , n28 );
    or g17 ( n33 , n115 , n256 );
    or g18 ( n110 , n55 , n18 );
    xnor g19 ( n68 , n227 , n21 );
    xnor g20 ( n181 , n187 , n45 );
    not g21 ( n49 , n26 );
    or g22 ( n126 , n90 , n235 );
    not g23 ( n225 , n12 );
    or g24 ( n202 , n103 , n235 );
    xnor g25 ( n200 , n186 , n23 );
    or g26 ( n30 , n78 , n101 );
    not g27 ( n123 , n137 );
    or g28 ( n281 , n193 , n169 );
    xnor g29 ( n50 , n179 , n87 );
    xnor g30 ( n164 , n28 , n15 );
    xor g31 ( n47 , n272 , n38 );
    not g32 ( n137 , n35 );
    or g33 ( n27 , n142 , n5 );
    not g34 ( n175 , n128 );
    or g35 ( n277 , n223 , n108 );
    and g36 ( n149 , n2 , n240 );
    xnor g37 ( n213 , n89 , n165 );
    not g38 ( n66 , n275 );
    not g39 ( n103 , n224 );
    or g40 ( n190 , n226 , n281 );
    not g41 ( n115 , n224 );
    or g42 ( n42 , n137 , n222 );
    not g43 ( n56 , n114 );
    xnor g44 ( n283 , n48 , n105 );
    or g45 ( n259 , n59 , n43 );
    or g46 ( n48 , n195 , n157 );
    not g47 ( n11 , n199 );
    or g48 ( n104 , n7 , n232 );
    xnor g49 ( n209 , n170 , n188 );
    not g50 ( n78 , n250 );
    or g51 ( n174 , n55 , n150 );
    not g52 ( n239 , n2 );
    xnor g53 ( n176 , n33 , n95 );
    or g54 ( n17 , n173 , n235 );
    xnor g55 ( n219 , n112 , n16 );
    not g56 ( n249 , n60 );
    xnor g57 ( n40 , n147 , n183 );
    or g58 ( n134 , n203 , n43 );
    and g59 ( n274 , n65 , n239 );
    or g60 ( n41 , n107 , n266 );
    xnor g61 ( n236 , n228 , n95 );
    xnor g62 ( n77 , n279 , n258 );
    or g63 ( n119 , n49 , n88 );
    xnor g64 ( n74 , n278 , n52 );
    and g65 ( n270 , n161 , n7 );
    or g66 ( n163 , n78 , n19 );
    xnor g67 ( n100 , n82 , n74 );
    xnor g68 ( n284 , n271 , n20 );
    xnor g69 ( n241 , n75 , n45 );
    or g70 ( n131 , n249 , n127 );
    xnor g71 ( n97 , n27 , n53 );
    xnor g72 ( n94 , n138 , n212 );
    xnor g73 ( n54 , n124 , n160 );
    not g74 ( n224 , n104 );
    not g75 ( n237 , n149 );
    xnor g76 ( n31 , n152 , n280 );
    not g77 ( n203 , n218 );
    xnor g78 ( n165 , n152 , n227 );
    nor g79 ( n129 , n237 , n190 );
    xnor g80 ( n193 , n71 , n62 );
    not g81 ( n166 , n26 );
    not g82 ( n256 , n247 );
    not g83 ( n107 , n136 );
    or g84 ( n144 , n166 , n163 );
    xnor g85 ( n2 , n245 , n217 );
    not g86 ( n240 , n65 );
    xnor g87 ( n153 , n276 , n95 );
    xnor g88 ( n111 , n264 , n83 );
    or g89 ( n268 , n173 , n36 );
    xnor g90 ( n29 , n28 , n1 );
    xnor g91 ( n125 , n8 , n31 );
    or g92 ( n51 , n180 , n196 );
    nor g93 ( n272 , n182 , n190 );
    or g94 ( n19 , n121 , n260 );
    not g95 ( n141 , n266 );
    not g96 ( n118 , n210 );
    or g97 ( n5 , n252 , n275 );
    xnor g98 ( n212 , n23 , n83 );
    or g99 ( n179 , n115 , n230 );
    or g100 ( n88 , n174 , n196 );
    xnor g101 ( n245 , n9 , n68 );
    xnor g102 ( n91 , n119 , n152 );
    and g103 ( n92 , n26 , n46 );
    xnor g104 ( n71 , n8 , n178 );
    and g105 ( n26 , n6 , n35 );
    xnor g106 ( n82 , n242 , n87 );
    or g107 ( n143 , n226 , n36 );
    xnor g108 ( n20 , n219 , n134 );
    xnor g109 ( n170 , n167 , n257 );
    or g110 ( n196 , n261 , n96 );
    or g111 ( n169 , n192 , n123 );
    not g112 ( n7 , n225 );
    not g113 ( n172 , n58 );
    xnor g114 ( n204 , n135 , n73 );
    or g115 ( n246 , n169 , n19 );
    not g116 ( n161 , n41 );
    or g117 ( n147 , n260 , n143 );
    not g118 ( n69 , n210 );
    xnor g119 ( n138 , n53 , n155 );
    or g120 ( n130 , n103 , n282 );
    xor g121 ( n265 , n238 , n79 );
    xor g122 ( n262 , n129 , n1 );
    not g123 ( n90 , n270 );
    xnor g124 ( n3 , n130 , n278 );
    xnor g125 ( n22 , n100 , n263 );
    xnor g126 ( n234 , n83 , n52 );
    or g127 ( n145 , n275 , n19 );
    xnor g128 ( n208 , n63 , n52 );
    or g129 ( n184 , n177 , n108 );
    or g130 ( n73 , n148 , n127 );
    xnor g131 ( n207 , n105 , n194 );
    xnor g132 ( n98 , n1 , n38 );
    xnor g133 ( n135 , n153 , n102 );
    xnor g134 ( n217 , n234 , n76 );
    xnor g135 ( n85 , n162 , n183 );
    or g136 ( n93 , n180 , n101 );
    xnor g137 ( n112 , n122 , n187 );
    or g138 ( n267 , n69 , n80 );
    or g139 ( n157 , n128 , n174 );
    or g140 ( n106 , n56 , n221 );
    xnor g141 ( n271 , n23 , n278 );
    and g142 ( n199 , n92 , n149 );
    or g143 ( n84 , n173 , n80 );
    not g144 ( n142 , n158 );
    or g145 ( n61 , n222 , n123 );
    xnor g146 ( n191 , n133 , n215 );
    not g147 ( n101 , n92 );
    not g148 ( n158 , n233 );
    xnor g149 ( n243 , n202 , n45 );
    not g150 ( n222 , n192 );
    or g151 ( n235 , n182 , n128 );
    xnor g152 ( n279 , n79 , n276 );
    or g153 ( n230 , n142 , n281 );
    not g154 ( n201 , n110 );
    xnor g155 ( n12 , n116 , n151 );
    not g156 ( n156 , n231 );
    not g157 ( n260 , n274 );
    not g158 ( n180 , n66 );
    xnor g159 ( n24 , n9 , n277 );
    xnor g160 ( n197 , n44 , n242 );
    xnor g161 ( n39 , n170 , n259 );
    xnor g162 ( n57 , n98 , n39 );
    xnor g163 ( n109 , n213 , n184 );
    or g164 ( n133 , n90 , n80 );
    or g165 ( n25 , n156 , n221 );
    and g166 ( n238 , n199 , n201 );
    not g167 ( n250 , n174 );
    xnor g168 ( n8 , n13 , n29 );
    xnor g169 ( n89 , n105 , n160 );
    or g170 ( n275 , n12 , n41 );
    not g171 ( n96 , n149 );
    xnor g172 ( n178 , n160 , n37 );
    xnor g173 ( n285 , n53 , n242 );
    or g174 ( n233 , n240 , n239 );
    xnor g175 ( n9 , n241 , n85 );
    not g176 ( n210 , n104 );
    not g177 ( n70 , n233 );
    not g178 ( n221 , n4 );
    or g179 ( n132 , n118 , n11 );
    or g180 ( n226 , n58 , n232 );
    not g181 ( n58 , n12 );
    xnor g182 ( n151 , n236 , n10 );
    or g183 ( n128 , n121 , n42 );
    or g184 ( n186 , n166 , n51 );
    not g185 ( n59 , n269 );
    xnor g186 ( n86 , n244 , n37 );
    xnor g187 ( n171 , n155 , n87 );
    xnor g188 ( n62 , n171 , n204 );
    xnor g189 ( n6 , n146 , n159 );
    not g190 ( n223 , n117 );
    or g191 ( n264 , n49 , n145 );
    xnor g192 ( n113 , n215 , n162 );
    xnor g193 ( n167 , n194 , n37 );
    not g194 ( n127 , n4 );
    xnor g195 ( n258 , n213 , n131 );
    xnor g196 ( n13 , n79 , n228 );
    not g197 ( n108 , n4 );
    xor g198 ( n139 , n189 , n155 );
    xnor g199 ( n220 , n144 , n227 );
    or g200 ( n44 , n195 , n251 );
    xnor g201 ( n65 , n125 , n284 );
    and g202 ( n247 , n92 , n274 );
    xnor g203 ( n102 , n15 , n38 );
    not g204 ( n252 , n175 );
    xnor g205 ( n255 , n94 , n113 );
    or g206 ( n150 , n136 , n266 );
    not g207 ( n229 , n70 );
    and g208 ( n0 , n199 , n270 );
    not g209 ( n182 , n274 );
    xnor g210 ( n67 , n164 , n109 );
    buf g211 ( n173 , n110 );
    xnor g212 ( n214 , n267 , n187 );
    not g213 ( n121 , n34 );
    xnor g214 ( n188 , n122 , n75 );
    xnor g215 ( n116 , n100 , n181 );
    or g216 ( n216 , n229 , n268 );
    or g217 ( n14 , n173 , n282 );
    not g218 ( n192 , n6 );
    xnor g219 ( n146 , n219 , n207 );
    or g220 ( n36 , n261 , n61 );
    xnor g221 ( n154 , n64 , n206 );
    and g222 ( n120 , n247 , n270 );
    xnor g223 ( n32 , n132 , n228 );
    nor g224 ( n189 , n233 , n93 );
    xnor g225 ( n205 , n253 , n21 );
    xnor g226 ( n266 , n255 , n67 );
    xnor g227 ( n35 , n22 , n57 );
    xor g228 ( n185 , n140 , n276 );
    xnor g229 ( n211 , n84 , n122 );
    not g230 ( n46 , n193 );
    or g231 ( n64 , n96 , n143 );
    or g232 ( n253 , n173 , n246 );
    not g233 ( n195 , n158 );
    not g234 ( n34 , n46 );
    or g235 ( n124 , n229 , n30 );
    or g236 ( n232 , n107 , n141 );
    xnor g237 ( n10 , n94 , n106 );
    or g238 ( n63 , n69 , n246 );
    xnor g239 ( n273 , n17 , n75 );
    or g240 ( n251 , n36 , n118 );
    xor g241 ( n248 , n120 , n15 );
    xnor g242 ( n76 , n135 , n25 );
    or g243 ( n282 , n169 , n196 );
    xnor g244 ( n99 , n14 , n280 );
endmodule
