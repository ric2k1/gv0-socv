module top( n5 , n13 , n17 , n20 , n27 , n36 , n37 , n53 , n62 , n75 , n80 , n86 , n93 , n105 , n106 , n111 , n117 , n139 , n145 , n147 , n157 , n161 , n175 , n176 , n182 , n190 , n198 , n204 , n208 , n214 , n217 , n219 , n224 , n225 , n226 , n229 , n235 , n241 , n244 , n249 , n256 , n281 , n287 , n289 , n294 , n300 , n303 , n319 , n345 , n346 , n364 , n365 , n368 , n384 , n387 , n389 , n393 , n403 , n409 , n410 , n417 , n430 , n439 , n442 , n457 , n465 , n473 , n477 , n489 , n491 , n493 , n503 , n506 , n511 , n515 , n518 , n521 , n532 , n537 , n587 , n588 , n593 , n594 , n595 , n606 , n618 , n630 , n642 , n648 , n656 , n671 , n680 , n684 , n690 , n691 , n693 , n699 , n702 , n703 , n704 , n706 , n716 , n741 , n742 , n743 , n746 , n753 , n756 , n765 , n777 , n782 , n788 );
    input n5 , n13 , n17 , n20 , n36 , n37 , n53 , n75 , n80 , n86 , n93 , n105 , n106 , n111 , n117 , n139 , n147 , n157 , n161 , n182 , n190 , n198 , n204 , n208 , n214 , n217 , n219 , n224 , n226 , n229 , n235 , n244 , n249 , n281 , n287 , n289 , n300 , n303 , n319 , n346 , n364 , n365 , n368 , n384 , n393 , n403 , n409 , n410 , n417 , n439 , n457 , n465 , n473 , n477 , n503 , n506 , n511 , n518 , n521 , n532 , n537 , n587 , n588 , n593 , n594 , n595 , n606 , n642 , n648 , n656 , n671 , n680 , n684 , n690 , n693 , n699 , n702 , n706 , n716 , n741 , n742 , n743 , n746 , n777 , n782 , n788 ;
    output n27 , n62 , n145 , n175 , n176 , n225 , n241 , n256 , n294 , n345 , n387 , n389 , n430 , n442 , n489 , n491 , n493 , n515 , n618 , n630 , n691 , n703 , n704 , n753 , n756 , n765 ;
    wire n0 , n1 , n2 , n3 , n4 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n14 , n15 , n16 , n18 , n19 , n21 , n22 , n23 , n24 , n25 , n26 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n76 , n77 , n78 , n79 , n81 , n82 , n83 , n84 , n85 , n87 , n88 , n89 , n90 , n91 , n92 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n107 , n108 , n109 , n110 , n112 , n113 , n114 , n115 , n116 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n140 , n141 , n142 , n143 , n144 , n146 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n158 , n159 , n160 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n177 , n178 , n179 , n180 , n181 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n199 , n200 , n201 , n202 , n203 , n205 , n206 , n207 , n209 , n210 , n211 , n212 , n213 , n215 , n216 , n218 , n220 , n221 , n222 , n223 , n227 , n228 , n230 , n231 , n232 , n233 , n234 , n236 , n237 , n238 , n239 , n240 , n242 , n243 , n245 , n246 , n247 , n248 , n250 , n251 , n252 , n253 , n254 , n255 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n282 , n283 , n284 , n285 , n286 , n288 , n290 , n291 , n292 , n293 , n295 , n296 , n297 , n298 , n299 , n301 , n302 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n366 , n367 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n385 , n386 , n388 , n390 , n391 , n392 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n404 , n405 , n406 , n407 , n408 , n411 , n412 , n413 , n414 , n415 , n416 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n440 , n441 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n474 , n475 , n476 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n490 , n492 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n504 , n505 , n507 , n508 , n509 , n510 , n512 , n513 , n514 , n516 , n517 , n519 , n520 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n533 , n534 , n535 , n536 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n589 , n590 , n591 , n592 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n643 , n644 , n645 , n646 , n647 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n681 , n682 , n683 , n685 , n686 , n687 , n688 , n689 , n692 , n694 , n695 , n696 , n697 , n698 , n700 , n701 , n705 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n744 , n745 , n747 , n748 , n749 , n750 , n751 , n752 , n754 , n755 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n778 , n779 , n780 , n781 , n783 , n784 , n785 , n786 , n787 , n789 ;
assign n8 = n559 | n136;
assign n676 = n578 & n778;
assign n683 = ~(n403 | n783);
assign n213 = n293 | n774;
assign n273 = ~(n300 | n250);
assign n34 = ~(n196 | n40);
assign n109 = n787 & n405;
assign n122 = n114 & n600;
assign n645 = ~(n452 | n488);
assign n621 = n433 | n106;
assign n312 = n381 | n296;
assign n534 = ~n226;
assign n657 = n341 | n59;
assign n6 = ~(n393 | n447);
assign n778 = ~n268;
assign n673 = n717 | n737;
assign n634 = n692 & n597;
assign n719 = ~(n452 | n655);
assign n644 = ~(n475 ^ n716);
assign n323 = ~(n648 | n223);
assign n646 = ~n5;
assign n369 = n46 & n230;
assign n681 = ~n521;
assign n411 = n760 & n88;
assign n600 = ~(n656 | n155);
assign n698 = ~(n452 | n552);
assign n774 = n656 & n695;
assign n311 = ~(n751 ^ n680);
assign n586 = n391 | n652;
assign n206 = n165 | n153;
assign n760 = ~n202;
assign n628 = ~n157;
assign n91 = n165 & n153;
assign n493 = n309 | n12;
assign n203 = n38 | n697;
assign n375 = n686 | n772;
assign n288 = n150 | n598;
assign n268 = n522 & n443;
assign n31 = n459 | n656;
assign n415 = ~(n98 | n363);
assign n685 = n546 | n276;
assign n63 = n131 & n627;
assign n764 = n656 & n135;
assign n707 = n452 | n761;
assign n450 = n666 & n257;
assign n52 = n391 & n767;
assign n772 = n452 | n270;
assign n252 = ~(n166 | n189);
assign n466 = n75 & n452;
assign n399 = ~n603;
assign n16 = n42 & n29;
assign n207 = ~(n537 | n212);
assign n277 = n581 & n248;
assign n407 = ~n749;
assign n574 = n607 | n264;
assign n383 = ~n520;
assign n169 = ~n236;
assign n97 = n537 | n300;
assign n559 = ~n393;
assign n14 = ~(n440 ^ n19);
assign n762 = ~(n484 | n635);
assign n589 = ~(n656 | n568);
assign n462 = n42 | n29;
assign n110 = ~(n403 | n590);
assign n258 = n331 | n121;
assign n257 = n546 & n757;
assign n639 = n16 | n752;
assign n661 = ~n351;
assign n127 = ~n106;
assign n655 = ~(n749 ^ n163);
assign n48 = ~(n656 | n674);
assign n678 = ~(n417 | n550);
assign n381 = ~n439;
assign n65 = ~(n582 ^ n788);
assign n153 = n609 & n81;
assign n615 = ~(n409 ^ n642);
assign n264 = ~n584;
assign n452 = ~n656;
assign n177 = ~(n643 ^ n780);
assign n200 = n728 | n694;
assign n42 = n591 & n288;
assign n173 = n330 & n599;
assign n533 = ~(n452 | n676);
assign n269 = ~(n439 | n117);
assign n233 = n559 | n779;
assign n167 = ~n300;
assign n552 = ~(n228 ^ n487);
assign n76 = n766 | n158;
assign n664 = ~n642;
assign n471 = n559 | n436;
assign n186 = ~n713;
assign n456 = n300 | n106;
assign n604 = ~(n656 | n3);
assign n557 = n37 & n501;
assign n643 = n460 | n7;
assign n56 = ~(n656 | n140);
assign n688 = ~n700;
assign n519 = ~n17;
assign n199 = n362 & n397;
assign n602 = ~n786;
assign n251 = n127 | n74;
assign n766 = n503 & n182;
assign n126 = ~n657;
assign n185 = n660 & n441;
assign n755 = n202 | n560;
assign n154 = ~(n384 | n129);
assign n133 = ~(n693 | n17);
assign n659 = n746 & n127;
assign n163 = n152 & n596;
assign n274 = n656 & n776;
assign n733 = ~(n214 | n69);
assign n514 = ~(n355 | n536);
assign n77 = n656 & n71;
assign n336 = ~(n228 | n372);
assign n115 = ~(n452 | n544);
assign n376 = n656 | n563;
assign n222 = ~n148;
assign n597 = n393 | n454;
assign n360 = n356 | n299;
assign n228 = n535 | n274;
assign n391 = ~n680;
assign n636 = n626 | n641;
assign n350 = n458 | n613;
assign n170 = ~(n649 | n376);
assign n461 = ~(n350 | n0);
assign n181 = n595 & n452;
assign n526 = n767 ^ n453;
assign n316 = n393 | n508;
assign n516 = ~(n439 ^ n742);
assign n686 = ~(n513 | n28);
assign n50 = n218 & n396;
assign n168 = n656 & n444;
assign n480 = ~n592;
assign n70 = ~(n656 | n631);
assign n441 = ~n19;
assign n549 = n628 | n340;
assign n490 = n228 & n372;
assign n497 = n656 & n408;
assign n267 = n403 & n311;
assign n174 = n23 | n520;
assign n581 = ~n159;
assign n30 = n519 | n423;
assign n143 = n366 & n369;
assign n502 = ~(n705 | n251);
assign n582 = n125 | n353;
assign n380 = n462 & n639;
assign n529 = ~(n656 | n388);
assign n736 = n621 | n553;
assign n540 = ~(n759 | n246);
assign n607 = n690 & n217;
assign n58 = n687 | n148;
assign n404 = ~(n189 ^ n61);
assign n618 = n589 | n576;
assign n763 = ~(n300 | n789);
assign n753 = n47 | n395;
assign n561 = n547 & n260;
assign n102 = ~(n452 | n385);
assign n29 = ~n68;
assign n39 = ~(n452 | n33);
assign n292 = ~n287;
assign n573 = ~(n440 | n441);
assign n354 = ~n330;
assign n262 = n525 | n524;
assign n197 = ~(n157 | n303);
assign n332 = n174 & n509;
assign n396 = n549 | n374;
assign n114 = n297 | n60;
assign n520 = ~(n574 ^ n690);
assign n339 = ~(n527 | n667);
assign n25 = ~(n537 | n286);
assign n494 = ~(n724 | n35);
assign n592 = n506 & n169;
assign n155 = ~(n495 | n556);
assign n241 = n731 | n698;
assign n130 = ~(n76 ^ n777);
assign n270 = n513 & n28;
assign n221 = n518 & n452;
assign n717 = n352 & n516;
assign n507 = ~(n726 | n193);
assign n726 = n754 | n497;
assign n230 = n608 & n237;
assign n385 = ~(n213 ^ n230);
assign n555 = ~(n17 ^ n13);
assign n340 = ~n303;
assign n756 = n386 | n172;
assign n560 = n688 & n314;
assign n98 = ~(n78 | n470);
assign n322 = n656 & n344;
assign n697 = n403 | n537;
assign n565 = n73 | n446;
assign n119 = ~(n787 | n405);
assign n663 = n735 | n200;
assign n370 = ~(n185 | n727);
assign n256 = n160 | n321;
assign n749 = n632 | n476;
assign n694 = ~n76;
assign n327 = n127 | n714;
assign n735 = ~n281;
assign n486 = ~(n452 | n432);
assign n132 = ~n200;
assign n296 = ~n742;
assign n525 = ~n648;
assign n499 = ~(n300 | n485);
assign n227 = n15 | n668;
assign n695 = ~(n236 ^ n506);
assign n725 = n373 & n101;
assign n331 = ~n417;
assign n438 = n368 & n452;
assign n547 = ~n549;
assign n400 = n292 | n656;
assign n246 = ~(n355 ^ n141);
assign n701 = n660 | n19;
assign n189 = n32 | n658;
assign n476 = n656 & n770;
assign n583 = n44 | n380;
assign n566 = ~n636;
assign n131 = n412 | n787;
assign n530 = ~n299;
assign n687 = ~n672;
assign n789 = n137 & n327;
assign n239 = n608 | n636;
assign n348 = n20 & n57;
assign n669 = n666 | n685;
assign n46 = ~n213;
assign n341 = n161 & n452;
assign n286 = ~(n313 | n763);
assign n108 = ~(n350 ^ n369);
assign n771 = n78 & n470;
assign n430 = n494 | n307;
assign n609 = n688 | n164;
assign n148 = n407 | n232;
assign n775 = ~(n5 ^ n157);
assign n692 = n559 | n418;
assign n32 = n439 & n117;
assign n263 = ~(n258 ^ n20);
assign n454 = ~(n358 | n482);
assign n479 = ~n606;
assign n255 = ~n490;
assign n62 = n604 | n87;
assign n489 = n56 | n102;
assign n142 = n559 | n722;
assign n193 = n687 & n392;
assign n548 = ~(n759 | n615);
assign n278 = ~(n64 | n625);
assign n470 = n495 | n778;
assign n202 = n700 & n164;
assign n55 = n244 & n452;
assign n469 = n656 & n65;
assign n247 = n547 | n197;
assign n144 = ~(n656 | n496);
assign n553 = n272 | n97;
assign n750 = n24 & n193;
assign n329 = n532 & n452;
assign n632 = n743 & n452;
assign n611 = n715 & n623;
assign n220 = n702 & n452;
assign n405 = ~(n184 ^ n422);
assign n759 = ~n537;
assign n343 = n116 | n603;
assign n483 = ~(n159 ^ n248);
assign n345 = n144 | n696;
assign n712 = n14 & n173;
assign n95 = n429 | n539;
assign n183 = ~n706;
assign n458 = n224 & n452;
assign n783 = ~(n577 | n207);
assign n603 = n24 | n58;
assign n758 = ~n384;
assign n211 = ~(n94 | n169);
assign n652 = ~n594;
assign n382 = n455 | n747;
assign n569 = ~(n452 | n10);
assign n429 = n235 & n452;
assign n721 = n46 | n239;
assign n242 = ~(n540 | n191);
assign n492 = n300 & n404;
assign n445 = ~(n439 ^ n117);
assign n435 = ~(n700 ^ n314);
assign n640 = n412 & n787;
assign n41 = n662 | n480;
assign n402 = n400 & n375;
assign n201 = ~(n377 | n647);
assign n421 = ~(n284 | n380);
assign n724 = n617 & n638;
assign n428 = n184 & n240;
assign n413 = ~(n349 ^ n445);
assign n243 = n452 | n379;
assign n660 = ~n440;
assign n424 = n620 | n178;
assign n146 = ~n190;
assign n704 = n624 | n533;
assign n362 = n472 | n335;
assign n158 = ~(n720 | n28);
assign n614 = ~n582;
assign n123 = ~(n217 ^ n365);
assign n770 = ~(n154 | n661);
assign n718 = ~n663;
assign n576 = n206 & n134;
assign n527 = ~n382;
assign n45 = ~(n298 | n718);
assign n24 = ~n726;
assign n658 = ~(n349 | n269);
assign n769 = n610 | n650;
assign n113 = ~n685;
assign n28 = n586 & n781;
assign n1 = ~(n452 | n177);
assign n596 = n185 | n173;
assign n196 = ~(n741 | n713);
assign n440 = n221 | n261;
assign n408 = ~(n323 | n390);
assign n612 = ~(n36 | n348);
assign n460 = n587 & n452;
assign n482 = ~(n403 | n242);
assign n103 = ~n669;
assign n238 = n249 & n439;
assign n394 = ~n564;
assign n558 = ~n214;
assign n500 = n120 & n748;
assign n578 = n522 | n443;
assign n156 = n336 | n490;
assign n554 = ~n741;
assign n416 = ~(n367 | n171);
assign n0 = ~n721;
assign n101 = n478 | n290;
assign n727 = ~n152;
assign n314 = n481 & n85;
assign n129 = n699 & n718;
assign n512 = n364 & n452;
assign n508 = ~(n267 | n110);
assign n317 = ~(n619 ^ n503);
assign n149 = ~(n656 | n538);
assign n23 = ~n503;
assign n682 = ~(n700 | n314);
assign n544 = ~(n505 ^ n257);
assign n635 = n656 | n2;
assign n517 = ~(n359 | n128);
assign n780 = n179 & n487;
assign n89 = n628 | n739;
assign n225 = n271 | n531;
assign n351 = n758 | n320;
assign n356 = ~n245;
assign n309 = ~(n461 | n670);
assign n218 = n646 | n107;
assign n231 = ~n402;
assign n412 = ~n184;
assign n324 = ~n69;
assign n371 = ~(n657 ^ n567);
assign n732 = n537 & n304;
assign n359 = n473 & n127;
assign n484 = n435 & n285;
assign n54 = ~(n495 ^ n268);
assign n118 = ~(n749 ^ n49);
assign n605 = n428 | n580;
assign n487 = n116 & n750;
assign n398 = n416 | n113;
assign n357 = ~(n334 | n354);
assign n740 = n157 & n393;
assign n84 = n343 & n529;
assign n307 = ~(n452 | n26);
assign n786 = n558 | n324;
assign n776 = ~(n678 | n57);
assign n297 = ~n495;
assign n443 = n356 & n143;
assign n590 = ~(n732 | n572);
assign n510 = n229 & n452;
assign n260 = n5 ^ n671;
assign n531 = ~(n452 | n679);
assign n501 = n53 & n602;
assign n74 = n30 & n729;
assign n620 = n503 & n611;
assign n389 = n72 | n543;
assign n321 = ~(n452 | n483);
assign n768 = ~n240;
assign n22 = n55 | n708;
assign n236 = n681 | n4;
assign n378 = n14 | n173;
assign n349 = n664 | n479;
assign n495 = n310 | n83;
assign n641 = ~n446;
assign n67 = ~(n284 | n420);
assign n172 = ~(n452 | n371);
assign n432 = ~(n629 ^ n755);
assign n81 = n682 | n21;
assign n474 = ~(n78 ^ n114);
assign n747 = ~(n452 | n247);
assign n290 = n51 & n504;
assign n209 = ~(n672 | n222);
assign n73 = ~(n159 | n318);
assign n406 = ~(n663 ^ n699);
assign n3 = ~(n290 ^ n67);
assign n59 = n656 & n644;
assign n505 = n512 | n469;
assign n308 = ~(n672 ^ n392);
assign n444 = ~(n612 | n614);
assign n35 = n656 | n11;
assign n546 = ~n367;
assign n737 = n127 | n315;
assign n386 = n419 & n434;
assign n330 = n472 | n677;
assign n134 = ~(n452 | n91);
assign n730 = ~n41;
assign n773 = ~(n452 | n130);
assign n467 = ~(n657 | n563);
assign n622 = ~(n452 | n712);
assign n223 = n457 & n661;
assign n591 = n183 | n656;
assign n691 = n9 | n415;
assign n302 = n42 & n68;
assign n434 = ~(n656 | n467);
assign n138 = n656 | n556;
assign n145 = n84 | n39;
assign n675 = ~(n505 ^ n113);
assign n433 = ~n319;
assign n472 = ~n283;
assign n563 = ~n333;
assign n51 = n42 | n68;
assign n187 = n220 | n99;
assign n668 = n347 | n266;
assign n723 = ~(n95 ^ n450);
assign n535 = n465 & n452;
assign n9 = ~(n656 | n474);
assign n191 = ~(n537 | n431);
assign n387 = n170 | n637;
assign n475 = n554 | n186;
assign n513 = ~(n503 ^ n182);
assign n528 = ~n574;
assign n192 = ~(n167 | n413);
assign n667 = n740 | n295;
assign n250 = n90 & n673;
assign n66 = n534 | n656;
assign n305 = n522 & n360;
assign n100 = n785 & n424;
assign n585 = n656 & n45;
assign n254 = ~(n187 | n566);
assign n333 = n275 | n669;
assign n104 = ~(n680 ^ n594);
assign n551 = ~(n786 ^ n53);
assign n754 = n588 & n452;
assign n152 = n660 | n441;
assign n69 = n208 & n730;
assign n784 = ~n111;
assign n447 = ~(n403 | n18);
assign n64 = n693 & n17;
assign n781 = n280 | n50;
assign n194 = ~n210;
assign n373 = n402 | n210;
assign n463 = ~(n367 ^ n757);
assign n175 = n768 | n339;
assign n377 = ~(n17 | n782);
assign n610 = ~(n37 | n501);
assign n779 = ~(n332 ^ n43);
assign n26 = ~(n605 ^ n616);
assign n488 = n44 & n380;
assign n99 = n656 & n211;
assign n347 = n393 | n403;
assign n283 = n151 | n585;
assign n353 = ~n348;
assign n703 = n48 | n1;
assign n729 = n312 & n326;
assign n291 = ~(n642 ^ n606);
assign n638 = ~(n42 ^ n29);
assign n448 = ~(n283 | n677);
assign n248 = n126 & n567;
assign n679 = ~(n245 ^ n143);
assign n395 = ~(n452 | n451);
assign n625 = n238 | n514;
assign n71 = ~(n162 ^ n147);
assign n731 = ~(n656 | n156);
assign n38 = ~n93;
assign n363 = n452 | n771;
assign n124 = ~(n739 | n279);
assign n374 = ~(n5 | n671);
assign n538 = ~(n188 ^ n446);
assign n426 = ~(n555 | n729);
assign n579 = n656 | n109;
assign n295 = n89 & n6;
assign n584 = n449 | n265;
assign n650 = n452 | n557;
assign n15 = n711 | n106;
assign n313 = ~(n167 | n291);
assign n82 = ~(n184 | n240);
assign n536 = ~(n249 | n439);
assign n710 = ~(n633 | n730);
assign n361 = n573 | n199;
assign n564 = n716 & n40;
assign n392 = n407 & n163;
assign n121 = ~n550;
assign n491 = n70 | n498;
assign n179 = ~n228;
assign n562 = ~(n452 | n54);
assign n623 = n52 | n123;
assign n33 = ~(n22 ^ n750);
assign n180 = n147 & n523;
assign n285 = ~n725;
assign n68 = n112 & n316;
assign n478 = ~(n231 | n194);
assign n498 = ~(n507 | n243);
assign n715 = n391 | n767;
assign n320 = ~n129;
assign n677 = ~n335;
assign n92 = ~n511;
assign n79 = n104 & n50;
assign n212 = ~(n201 | n499);
assign n575 = ~(n188 ^ n277);
assign n326 = n352 | n216;
assign n713 = n788 & n614;
assign n709 = ~n643;
assign n437 = n393 | n651;
assign n379 = n726 & n193;
assign n275 = ~n95;
assign n116 = ~n22;
assign n388 = ~(n22 | n399);
assign n310 = n410 & n452;
assign n556 = ~n60;
assign n651 = ~(n601 | n683);
assign n601 = n403 & n317;
assign n335 = n736 & n233;
assign n739 = ~n403;
assign n276 = n709 | n255;
assign n515 = n653 | n719;
assign n481 = n393 | n427;
assign n571 = n656 & n195;
assign n617 = ~n63;
assign n696 = n378 & n622;
assign n464 = ~(n452 | n575);
assign n245 = n466 | n571;
assign n672 = n438 | n322;
assign n504 = n302 | n63;
assign n176 = n762 | n486;
assign n271 = ~(n656 | n541);
assign n419 = n126 | n333;
assign n522 = n31 & n707;
assign n165 = ~(n283 ^ n335);
assign n670 = n656 | n530;
assign n11 = ~(n617 | n638);
assign n261 = n656 & n406;
assign n568 = ~(n411 ^ n357);
assign n150 = ~(n104 | n50);
assign n141 = ~(n249 ^ n439);
assign n662 = ~n86;
assign n734 = ~n58;
assign n40 = ~n475;
assign n401 = ~(n262 ^ n204);
assign n397 = n448 | n411;
assign n112 = n559 | n526;
assign n334 = n472 & n677;
assign n567 = n275 & n450;
assign n572 = ~(n537 | n328);
assign n171 = ~n276;
assign n294 = n342 | n115;
assign n748 = ~(n452 | n561);
assign n509 = n205 | n100;
assign n159 = n329 | n764;
assign n272 = n393 | n403;
assign n352 = n664 | n784;
assign n282 = ~(n456 | n203);
assign n19 = n227 & n142;
assign n94 = ~(n521 | n180);
assign n580 = ~(n82 | n422);
assign n279 = n23 | n619;
assign n280 = ~(n680 | n594);
assign n7 = n656 & n263;
assign n616 = ~(n42 ^ n68);
assign n265 = ~n365;
assign n423 = ~n13;
assign n751 = n646 | n628;
assign n523 = ~n162;
assign n425 = ~(n452 | n463);
assign n125 = ~n36;
assign n372 = ~n343;
assign n253 = n346 & n452;
assign n665 = ~(n693 ^ n17);
assign n160 = ~(n656 | n565);
assign n633 = ~(n86 | n592);
assign n627 = n640 | n634;
assign n195 = ~(n41 ^ n208);
assign n390 = ~n262;
assign n446 = n159 & n318;
assign n631 = ~(n726 ^ n734);
assign n542 = ~n239;
assign n711 = ~n139;
assign n577 = ~(n133 | n325);
assign n87 = n583 & n645;
assign n708 = n656 & n401;
assign n744 = ~(n178 ^ n503);
assign n599 = n334 | n153;
assign n598 = n452 | n79;
assign n43 = n215 | n528;
assign n761 = n733 | n602;
assign n422 = ~n634;
assign n78 = n66 & n769;
assign n366 = ~n350;
assign n757 = n709 & n780;
assign n418 = ~(n5 ^ n365);
assign n649 = ~(n95 | n103);
assign n284 = n402 & n194;
assign n215 = ~n690;
assign n414 = ~n409;
assign n720 = ~(n503 | n182);
assign n451 = ~(n240 ^ n405);
assign n442 = n122 | n562;
assign n325 = n759 | n278;
assign n745 = ~(n300 | n517);
assign n107 = ~n671;
assign n626 = ~n188;
assign n240 = n382 | n689;
assign n420 = n231 & n210;
assign n135 = ~(n545 | n523);
assign n301 = n127 | n738;
assign n674 = ~(n643 ^ n490);
assign n44 = ~(n231 ^ n210);
assign n96 = ~(n306 | n100);
assign n205 = ~(n503 | n383);
assign n315 = ~(n352 | n516);
assign n367 = n181 | n168;
assign n57 = ~n258;
assign n705 = ~(n17 | n13);
assign n61 = ~(n17 ^ n782);
assign n550 = n204 & n390;
assign n624 = ~(n305 | n138);
assign n164 = ~n314;
assign n714 = ~(n642 ^ n111);
assign n468 = ~n289;
assign n47 = ~(n119 | n579);
assign n608 = ~n187;
assign n647 = n167 | n252;
assign n629 = n420 | n421;
assign n700 = n253 | n773;
assign n630 = n234 | n425;
assign n654 = ~(n209 | n734);
assign n216 = ~(n439 | n742);
assign n293 = n80 & n452;
assign n266 = n537 | n300;
assign n728 = ~n777;
assign n128 = ~(n426 | n301);
assign n449 = ~n217;
assign n689 = ~n667;
assign n337 = n593 & n452;
assign n2 = ~(n435 | n285);
assign n765 = n338 | n569;
assign n162 = n146 | n394;
assign n140 = ~(n213 ^ n542);
assign n436 = n306 & n100;
assign n338 = ~(n656 | n570);
assign n237 = n626 & n277;
assign n136 = ~(n611 ^ n744);
assign n752 = ~n605;
assign n619 = n391 | n751;
assign n18 = n548 | n25;
assign n485 = ~(n659 | n502);
assign n543 = ~(n452 | n308);
assign n342 = ~(n656 | n675);
assign n4 = ~n180;
assign n539 = n656 & n34;
assign n431 = ~(n192 | n273);
assign n455 = n684 & n452;
assign n90 = n92 | n106;
assign n137 = n468 | n106;
assign n304 = ~(n625 ^ n665);
assign n232 = n701 & n361;
assign n85 = n96 | n471;
assign n785 = n503 | n611;
assign n27 = n149 | n464;
assign n666 = ~n505;
assign n210 = n437 & n8;
assign n358 = ~(n739 | n775);
assign n496 = ~(n199 ^ n370);
assign n21 = ~n629;
assign n184 = n337 | n500;
assign n259 = ~(n584 ^ n217);
assign n541 = ~(n245 ^ n530);
assign n298 = ~(n281 | n132);
assign n49 = ~n232;
assign n10 = ~(n187 ^ n237);
assign n299 = n366 | n721;
assign n722 = n43 | n332;
assign n88 = n560 | n725;
assign n344 = ~(n351 ^ n457);
assign n12 = ~(n452 | n108);
assign n188 = n510 | n77;
assign n653 = ~(n656 | n118);
assign n459 = ~n105;
assign n178 = ~(n259 ^ n690);
assign n427 = ~(n124 | n282);
assign n328 = ~(n492 | n745);
assign n355 = n414 | n664;
assign n545 = ~(n190 | n564);
assign n767 = n646 | n265;
assign n613 = n656 & n710;
assign n120 = n547 | n260;
assign n570 = n254 | n542;
assign n318 = ~n419;
assign n151 = n219 & n452;
assign n637 = ~(n452 | n723);
assign n306 = ~(n383 ^ n503);
assign n453 = ~(n123 ^ n680);
assign n524 = ~n223;
assign n787 = n527 | n689;
assign n72 = n452 & n654;
assign n234 = ~(n656 | n398);
assign n166 = n17 & n782;
assign n60 = n522 | n360;
assign n738 = n555 & n729;
assign n83 = n656 & n551;
endmodule
