module top(in1, in2, in3, out1, out2);
  input [15:0] in1, in2, in3;
  output [31:0] out1, out2;
  wire [15:0] in1, in2, in3;
  wire [31:0] out1, out2;
  wire csa_tree_add_7_27_groupi_n_0, csa_tree_add_7_27_groupi_n_1, csa_tree_add_7_27_groupi_n_2, csa_tree_add_7_27_groupi_n_3, csa_tree_add_7_27_groupi_n_6, csa_tree_add_7_27_groupi_n_7, csa_tree_add_7_27_groupi_n_8, csa_tree_add_7_27_groupi_n_9;
  wire csa_tree_add_7_27_groupi_n_10, csa_tree_add_7_27_groupi_n_11, csa_tree_add_7_27_groupi_n_12, csa_tree_add_7_27_groupi_n_13, csa_tree_add_7_27_groupi_n_14, csa_tree_add_7_27_groupi_n_15, csa_tree_add_7_27_groupi_n_16, csa_tree_add_7_27_groupi_n_17;
  wire csa_tree_add_7_27_groupi_n_18, csa_tree_add_7_27_groupi_n_19, csa_tree_add_7_27_groupi_n_20, csa_tree_add_7_27_groupi_n_21, csa_tree_add_7_27_groupi_n_22, csa_tree_add_7_27_groupi_n_23, csa_tree_add_7_27_groupi_n_24, csa_tree_add_7_27_groupi_n_25;
  wire csa_tree_add_7_27_groupi_n_26, csa_tree_add_7_27_groupi_n_27, csa_tree_add_7_27_groupi_n_28, csa_tree_add_7_27_groupi_n_29, csa_tree_add_7_27_groupi_n_30, csa_tree_add_7_27_groupi_n_31, csa_tree_add_7_27_groupi_n_32, csa_tree_add_7_27_groupi_n_33;
  wire csa_tree_add_7_27_groupi_n_34, csa_tree_add_7_27_groupi_n_35, csa_tree_add_7_27_groupi_n_36, csa_tree_add_7_27_groupi_n_37, csa_tree_add_7_27_groupi_n_38, csa_tree_add_7_27_groupi_n_39, csa_tree_add_7_27_groupi_n_40, csa_tree_add_7_27_groupi_n_41;
  wire csa_tree_add_7_27_groupi_n_42, csa_tree_add_7_27_groupi_n_43, csa_tree_add_7_27_groupi_n_44, csa_tree_add_7_27_groupi_n_45, csa_tree_add_7_27_groupi_n_46, csa_tree_add_7_27_groupi_n_47, csa_tree_add_7_27_groupi_n_48, csa_tree_add_7_27_groupi_n_49;
  wire csa_tree_add_7_27_groupi_n_50, csa_tree_add_7_27_groupi_n_51, csa_tree_add_7_27_groupi_n_52, csa_tree_add_7_27_groupi_n_53, csa_tree_add_7_27_groupi_n_54, csa_tree_add_7_27_groupi_n_55, csa_tree_add_7_27_groupi_n_56, csa_tree_add_7_27_groupi_n_57;
  wire csa_tree_add_7_27_groupi_n_58, csa_tree_add_7_27_groupi_n_59, csa_tree_add_7_27_groupi_n_60, csa_tree_add_7_27_groupi_n_61, csa_tree_add_7_27_groupi_n_62, csa_tree_add_7_27_groupi_n_63, csa_tree_add_7_27_groupi_n_64, csa_tree_add_7_27_groupi_n_65;
  wire csa_tree_add_7_27_groupi_n_66, csa_tree_add_7_27_groupi_n_67, csa_tree_add_7_27_groupi_n_68, csa_tree_add_7_27_groupi_n_69, csa_tree_add_7_27_groupi_n_70, csa_tree_add_7_27_groupi_n_71, csa_tree_add_7_27_groupi_n_72, csa_tree_add_7_27_groupi_n_73;
  wire csa_tree_add_7_27_groupi_n_74, csa_tree_add_7_27_groupi_n_75, csa_tree_add_7_27_groupi_n_76, csa_tree_add_7_27_groupi_n_77, csa_tree_add_7_27_groupi_n_78, csa_tree_add_7_27_groupi_n_79, csa_tree_add_7_27_groupi_n_80, csa_tree_add_7_27_groupi_n_81;
  wire csa_tree_add_7_27_groupi_n_82, csa_tree_add_7_27_groupi_n_83, csa_tree_add_7_27_groupi_n_84, csa_tree_add_7_27_groupi_n_85, csa_tree_add_7_27_groupi_n_86, csa_tree_add_7_27_groupi_n_87, csa_tree_add_7_27_groupi_n_88, csa_tree_add_7_27_groupi_n_89;
  wire csa_tree_add_7_27_groupi_n_90, csa_tree_add_7_27_groupi_n_91, csa_tree_add_7_27_groupi_n_92, csa_tree_add_7_27_groupi_n_93, csa_tree_add_7_27_groupi_n_94, csa_tree_add_7_27_groupi_n_95, csa_tree_add_7_27_groupi_n_96, csa_tree_add_7_27_groupi_n_97;
  wire csa_tree_add_7_27_groupi_n_98, csa_tree_add_7_27_groupi_n_99, csa_tree_add_7_27_groupi_n_100, csa_tree_add_7_27_groupi_n_101, csa_tree_add_7_27_groupi_n_102, csa_tree_add_7_27_groupi_n_103, csa_tree_add_7_27_groupi_n_104, csa_tree_add_7_27_groupi_n_105;
  wire csa_tree_add_7_27_groupi_n_106, csa_tree_add_7_27_groupi_n_107, csa_tree_add_7_27_groupi_n_108, csa_tree_add_7_27_groupi_n_109, csa_tree_add_7_27_groupi_n_110, csa_tree_add_7_27_groupi_n_111, csa_tree_add_7_27_groupi_n_112, csa_tree_add_7_27_groupi_n_113;
  wire csa_tree_add_7_27_groupi_n_114, csa_tree_add_7_27_groupi_n_115, csa_tree_add_7_27_groupi_n_116, csa_tree_add_7_27_groupi_n_117, csa_tree_add_7_27_groupi_n_118, csa_tree_add_7_27_groupi_n_119, csa_tree_add_7_27_groupi_n_120, csa_tree_add_7_27_groupi_n_121;
  wire csa_tree_add_7_27_groupi_n_122, csa_tree_add_7_27_groupi_n_123, csa_tree_add_7_27_groupi_n_124, csa_tree_add_7_27_groupi_n_125, csa_tree_add_7_27_groupi_n_126, csa_tree_add_7_27_groupi_n_127, csa_tree_add_7_27_groupi_n_128, csa_tree_add_7_27_groupi_n_129;
  wire csa_tree_add_7_27_groupi_n_130, csa_tree_add_7_27_groupi_n_131, csa_tree_add_7_27_groupi_n_132, csa_tree_add_7_27_groupi_n_133, csa_tree_add_7_27_groupi_n_134, csa_tree_add_7_27_groupi_n_135, csa_tree_add_7_27_groupi_n_136, csa_tree_add_7_27_groupi_n_137;
  wire csa_tree_add_7_27_groupi_n_138, csa_tree_add_7_27_groupi_n_139, csa_tree_add_7_27_groupi_n_140, csa_tree_add_7_27_groupi_n_141, csa_tree_add_7_27_groupi_n_142, csa_tree_add_7_27_groupi_n_143, csa_tree_add_7_27_groupi_n_144, csa_tree_add_7_27_groupi_n_145;
  wire csa_tree_add_7_27_groupi_n_146, csa_tree_add_7_27_groupi_n_147, csa_tree_add_7_27_groupi_n_148, csa_tree_add_7_27_groupi_n_149, csa_tree_add_7_27_groupi_n_150, csa_tree_add_7_27_groupi_n_151, csa_tree_add_7_27_groupi_n_152, csa_tree_add_7_27_groupi_n_153;
  wire csa_tree_add_7_27_groupi_n_154, csa_tree_add_7_27_groupi_n_155, csa_tree_add_7_27_groupi_n_156, csa_tree_add_7_27_groupi_n_157, csa_tree_add_7_27_groupi_n_158, csa_tree_add_7_27_groupi_n_159, csa_tree_add_7_27_groupi_n_160, csa_tree_add_7_27_groupi_n_161;
  wire csa_tree_add_7_27_groupi_n_162, csa_tree_add_7_27_groupi_n_163, csa_tree_add_7_27_groupi_n_164, csa_tree_add_7_27_groupi_n_165, csa_tree_add_7_27_groupi_n_166, csa_tree_add_7_27_groupi_n_167, csa_tree_add_7_27_groupi_n_168, csa_tree_add_7_27_groupi_n_169;
  wire csa_tree_add_7_27_groupi_n_170, csa_tree_add_7_27_groupi_n_171, csa_tree_add_7_27_groupi_n_172, csa_tree_add_7_27_groupi_n_173, csa_tree_add_7_27_groupi_n_174, csa_tree_add_7_27_groupi_n_175, csa_tree_add_7_27_groupi_n_176, csa_tree_add_7_27_groupi_n_177;
  wire csa_tree_add_7_27_groupi_n_178, csa_tree_add_7_27_groupi_n_179, csa_tree_add_7_27_groupi_n_180, csa_tree_add_7_27_groupi_n_181, csa_tree_add_7_27_groupi_n_182, csa_tree_add_7_27_groupi_n_183, csa_tree_add_7_27_groupi_n_184, csa_tree_add_7_27_groupi_n_185;
  wire csa_tree_add_7_27_groupi_n_186, csa_tree_add_7_27_groupi_n_187, csa_tree_add_7_27_groupi_n_188, csa_tree_add_7_27_groupi_n_189, csa_tree_add_7_27_groupi_n_190, csa_tree_add_7_27_groupi_n_191, csa_tree_add_7_27_groupi_n_192, csa_tree_add_7_27_groupi_n_193;
  wire csa_tree_add_7_27_groupi_n_194, csa_tree_add_7_27_groupi_n_195, csa_tree_add_7_27_groupi_n_196, csa_tree_add_7_27_groupi_n_197, csa_tree_add_7_27_groupi_n_198, csa_tree_add_7_27_groupi_n_199, csa_tree_add_7_27_groupi_n_200, csa_tree_add_7_27_groupi_n_201;
  wire csa_tree_add_7_27_groupi_n_202, csa_tree_add_7_27_groupi_n_203, csa_tree_add_7_27_groupi_n_204, csa_tree_add_7_27_groupi_n_205, csa_tree_add_7_27_groupi_n_206, csa_tree_add_7_27_groupi_n_207, csa_tree_add_7_27_groupi_n_208, csa_tree_add_7_27_groupi_n_209;
  wire csa_tree_add_7_27_groupi_n_210, csa_tree_add_7_27_groupi_n_211, csa_tree_add_7_27_groupi_n_212, csa_tree_add_7_27_groupi_n_213, csa_tree_add_7_27_groupi_n_214, csa_tree_add_7_27_groupi_n_215, csa_tree_add_7_27_groupi_n_216, csa_tree_add_7_27_groupi_n_217;
  wire csa_tree_add_7_27_groupi_n_218, csa_tree_add_7_27_groupi_n_219, csa_tree_add_7_27_groupi_n_220, csa_tree_add_7_27_groupi_n_221, csa_tree_add_7_27_groupi_n_222, csa_tree_add_7_27_groupi_n_223, csa_tree_add_7_27_groupi_n_224, csa_tree_add_7_27_groupi_n_225;
  wire csa_tree_add_7_27_groupi_n_226, csa_tree_add_7_27_groupi_n_227, csa_tree_add_7_27_groupi_n_228, csa_tree_add_7_27_groupi_n_229, csa_tree_add_7_27_groupi_n_230, csa_tree_add_7_27_groupi_n_231, csa_tree_add_7_27_groupi_n_232, csa_tree_add_7_27_groupi_n_233;
  wire csa_tree_add_7_27_groupi_n_234, csa_tree_add_7_27_groupi_n_235, csa_tree_add_7_27_groupi_n_236, csa_tree_add_7_27_groupi_n_237, csa_tree_add_7_27_groupi_n_238, csa_tree_add_7_27_groupi_n_239, csa_tree_add_7_27_groupi_n_240, csa_tree_add_7_27_groupi_n_241;
  wire csa_tree_add_7_27_groupi_n_242, csa_tree_add_7_27_groupi_n_243, csa_tree_add_7_27_groupi_n_244, csa_tree_add_7_27_groupi_n_245, csa_tree_add_7_27_groupi_n_246, csa_tree_add_7_27_groupi_n_247, csa_tree_add_7_27_groupi_n_248, csa_tree_add_7_27_groupi_n_249;
  wire csa_tree_add_7_27_groupi_n_250, csa_tree_add_7_27_groupi_n_251, csa_tree_add_7_27_groupi_n_252, csa_tree_add_7_27_groupi_n_253, csa_tree_add_7_27_groupi_n_254, csa_tree_add_7_27_groupi_n_255, csa_tree_add_7_27_groupi_n_256, csa_tree_add_7_27_groupi_n_257;
  wire csa_tree_add_7_27_groupi_n_258, csa_tree_add_7_27_groupi_n_259, csa_tree_add_7_27_groupi_n_260, csa_tree_add_7_27_groupi_n_261, csa_tree_add_7_27_groupi_n_262, csa_tree_add_7_27_groupi_n_263, csa_tree_add_7_27_groupi_n_264, csa_tree_add_7_27_groupi_n_265;
  wire csa_tree_add_7_27_groupi_n_266, csa_tree_add_7_27_groupi_n_267, csa_tree_add_7_27_groupi_n_268, csa_tree_add_7_27_groupi_n_269, csa_tree_add_7_27_groupi_n_270, csa_tree_add_7_27_groupi_n_271, csa_tree_add_7_27_groupi_n_272, csa_tree_add_7_27_groupi_n_273;
  wire csa_tree_add_7_27_groupi_n_274, csa_tree_add_7_27_groupi_n_275, csa_tree_add_7_27_groupi_n_276, csa_tree_add_7_27_groupi_n_277, csa_tree_add_7_27_groupi_n_278, csa_tree_add_7_27_groupi_n_279, csa_tree_add_7_27_groupi_n_280, csa_tree_add_7_27_groupi_n_281;
  wire csa_tree_add_7_27_groupi_n_282, csa_tree_add_7_27_groupi_n_283, csa_tree_add_7_27_groupi_n_284, csa_tree_add_7_27_groupi_n_285, csa_tree_add_7_27_groupi_n_286, csa_tree_add_7_27_groupi_n_287, csa_tree_add_7_27_groupi_n_288, csa_tree_add_7_27_groupi_n_289;
  wire csa_tree_add_7_27_groupi_n_290, csa_tree_add_7_27_groupi_n_291, csa_tree_add_7_27_groupi_n_292, csa_tree_add_7_27_groupi_n_293, csa_tree_add_7_27_groupi_n_294, csa_tree_add_7_27_groupi_n_295, csa_tree_add_7_27_groupi_n_296, csa_tree_add_7_27_groupi_n_297;
  wire csa_tree_add_7_27_groupi_n_298, csa_tree_add_7_27_groupi_n_299, csa_tree_add_7_27_groupi_n_300, csa_tree_add_7_27_groupi_n_301, csa_tree_add_7_27_groupi_n_302, csa_tree_add_7_27_groupi_n_303, csa_tree_add_7_27_groupi_n_304, csa_tree_add_7_27_groupi_n_305;
  wire csa_tree_add_7_27_groupi_n_306, csa_tree_add_7_27_groupi_n_307, csa_tree_add_7_27_groupi_n_308, csa_tree_add_7_27_groupi_n_309, csa_tree_add_7_27_groupi_n_310, csa_tree_add_7_27_groupi_n_311, csa_tree_add_7_27_groupi_n_312, csa_tree_add_7_27_groupi_n_313;
  wire csa_tree_add_7_27_groupi_n_314, csa_tree_add_7_27_groupi_n_315, csa_tree_add_7_27_groupi_n_316, csa_tree_add_7_27_groupi_n_317, csa_tree_add_7_27_groupi_n_318, csa_tree_add_7_27_groupi_n_319, csa_tree_add_7_27_groupi_n_320, csa_tree_add_7_27_groupi_n_321;
  wire csa_tree_add_7_27_groupi_n_322, csa_tree_add_7_27_groupi_n_323, csa_tree_add_7_27_groupi_n_324, csa_tree_add_7_27_groupi_n_325, csa_tree_add_7_27_groupi_n_326, csa_tree_add_7_27_groupi_n_327, csa_tree_add_7_27_groupi_n_328, csa_tree_add_7_27_groupi_n_329;
  wire csa_tree_add_7_27_groupi_n_330, csa_tree_add_7_27_groupi_n_331, csa_tree_add_7_27_groupi_n_332, csa_tree_add_7_27_groupi_n_333, csa_tree_add_7_27_groupi_n_334, csa_tree_add_7_27_groupi_n_335, csa_tree_add_7_27_groupi_n_336, csa_tree_add_7_27_groupi_n_337;
  wire csa_tree_add_7_27_groupi_n_338, csa_tree_add_7_27_groupi_n_339, csa_tree_add_7_27_groupi_n_340, csa_tree_add_7_27_groupi_n_341, csa_tree_add_7_27_groupi_n_342, csa_tree_add_7_27_groupi_n_343, csa_tree_add_7_27_groupi_n_344, csa_tree_add_7_27_groupi_n_345;
  wire csa_tree_add_7_27_groupi_n_346, csa_tree_add_7_27_groupi_n_347, csa_tree_add_7_27_groupi_n_348, csa_tree_add_7_27_groupi_n_349, csa_tree_add_7_27_groupi_n_350, csa_tree_add_7_27_groupi_n_351, csa_tree_add_7_27_groupi_n_352, csa_tree_add_7_27_groupi_n_353;
  wire csa_tree_add_7_27_groupi_n_354, csa_tree_add_7_27_groupi_n_355, csa_tree_add_7_27_groupi_n_356, csa_tree_add_7_27_groupi_n_357, csa_tree_add_7_27_groupi_n_358, csa_tree_add_7_27_groupi_n_359, csa_tree_add_7_27_groupi_n_360, csa_tree_add_7_27_groupi_n_361;
  wire csa_tree_add_7_27_groupi_n_362, csa_tree_add_7_27_groupi_n_363, csa_tree_add_7_27_groupi_n_364, csa_tree_add_7_27_groupi_n_365, csa_tree_add_7_27_groupi_n_366, csa_tree_add_7_27_groupi_n_367, csa_tree_add_7_27_groupi_n_368, csa_tree_add_7_27_groupi_n_369;
  wire csa_tree_add_7_27_groupi_n_370, csa_tree_add_7_27_groupi_n_371, csa_tree_add_7_27_groupi_n_372, csa_tree_add_7_27_groupi_n_373, csa_tree_add_7_27_groupi_n_374, csa_tree_add_7_27_groupi_n_375, csa_tree_add_7_27_groupi_n_376, csa_tree_add_7_27_groupi_n_377;
  wire csa_tree_add_7_27_groupi_n_378, csa_tree_add_7_27_groupi_n_379, csa_tree_add_7_27_groupi_n_380, csa_tree_add_7_27_groupi_n_381, csa_tree_add_7_27_groupi_n_382, csa_tree_add_7_27_groupi_n_383, csa_tree_add_7_27_groupi_n_384, csa_tree_add_7_27_groupi_n_385;
  wire csa_tree_add_7_27_groupi_n_386, csa_tree_add_7_27_groupi_n_387, csa_tree_add_7_27_groupi_n_388, csa_tree_add_7_27_groupi_n_389, csa_tree_add_7_27_groupi_n_390, csa_tree_add_7_27_groupi_n_391, csa_tree_add_7_27_groupi_n_392, csa_tree_add_7_27_groupi_n_393;
  wire csa_tree_add_7_27_groupi_n_394, csa_tree_add_7_27_groupi_n_395, csa_tree_add_7_27_groupi_n_396, csa_tree_add_7_27_groupi_n_397, csa_tree_add_7_27_groupi_n_398, csa_tree_add_7_27_groupi_n_399, csa_tree_add_7_27_groupi_n_400, csa_tree_add_7_27_groupi_n_401;
  wire csa_tree_add_7_27_groupi_n_402, csa_tree_add_7_27_groupi_n_403, csa_tree_add_7_27_groupi_n_404, csa_tree_add_7_27_groupi_n_405, csa_tree_add_7_27_groupi_n_406, csa_tree_add_7_27_groupi_n_407, csa_tree_add_7_27_groupi_n_408, csa_tree_add_7_27_groupi_n_409;
  wire csa_tree_add_7_27_groupi_n_410, csa_tree_add_7_27_groupi_n_411, csa_tree_add_7_27_groupi_n_412, csa_tree_add_7_27_groupi_n_413, csa_tree_add_7_27_groupi_n_414, csa_tree_add_7_27_groupi_n_415, csa_tree_add_7_27_groupi_n_416, csa_tree_add_7_27_groupi_n_417;
  wire csa_tree_add_7_27_groupi_n_418, csa_tree_add_7_27_groupi_n_419, csa_tree_add_7_27_groupi_n_420, csa_tree_add_7_27_groupi_n_421, csa_tree_add_7_27_groupi_n_422, csa_tree_add_7_27_groupi_n_423, csa_tree_add_7_27_groupi_n_424, csa_tree_add_7_27_groupi_n_425;
  wire csa_tree_add_7_27_groupi_n_426, csa_tree_add_7_27_groupi_n_427, csa_tree_add_7_27_groupi_n_428, csa_tree_add_7_27_groupi_n_429, csa_tree_add_7_27_groupi_n_430, csa_tree_add_7_27_groupi_n_431, csa_tree_add_7_27_groupi_n_432, csa_tree_add_7_27_groupi_n_433;
  wire csa_tree_add_7_27_groupi_n_434, csa_tree_add_7_27_groupi_n_435, csa_tree_add_7_27_groupi_n_436, csa_tree_add_7_27_groupi_n_437, csa_tree_add_7_27_groupi_n_438, csa_tree_add_7_27_groupi_n_439, csa_tree_add_7_27_groupi_n_440, csa_tree_add_7_27_groupi_n_441;
  wire csa_tree_add_7_27_groupi_n_442, csa_tree_add_7_27_groupi_n_443, csa_tree_add_7_27_groupi_n_444, csa_tree_add_7_27_groupi_n_445, csa_tree_add_7_27_groupi_n_446, csa_tree_add_7_27_groupi_n_447, csa_tree_add_7_27_groupi_n_448, csa_tree_add_7_27_groupi_n_449;
  wire csa_tree_add_7_27_groupi_n_450, csa_tree_add_7_27_groupi_n_451, csa_tree_add_7_27_groupi_n_452, csa_tree_add_7_27_groupi_n_453, csa_tree_add_7_27_groupi_n_454, csa_tree_add_7_27_groupi_n_455, csa_tree_add_7_27_groupi_n_456, csa_tree_add_7_27_groupi_n_457;
  wire csa_tree_add_7_27_groupi_n_458, csa_tree_add_7_27_groupi_n_459, csa_tree_add_7_27_groupi_n_460, csa_tree_add_7_27_groupi_n_461, csa_tree_add_7_27_groupi_n_462, csa_tree_add_7_27_groupi_n_463, csa_tree_add_7_27_groupi_n_464, csa_tree_add_7_27_groupi_n_465;
  wire csa_tree_add_7_27_groupi_n_466, csa_tree_add_7_27_groupi_n_467, csa_tree_add_7_27_groupi_n_468, csa_tree_add_7_27_groupi_n_469, csa_tree_add_7_27_groupi_n_470, csa_tree_add_7_27_groupi_n_471, csa_tree_add_7_27_groupi_n_472, csa_tree_add_7_27_groupi_n_473;
  wire csa_tree_add_7_27_groupi_n_474, csa_tree_add_7_27_groupi_n_475, csa_tree_add_7_27_groupi_n_476, csa_tree_add_7_27_groupi_n_477, csa_tree_add_7_27_groupi_n_478, csa_tree_add_7_27_groupi_n_479, csa_tree_add_7_27_groupi_n_480, csa_tree_add_7_27_groupi_n_481;
  wire csa_tree_add_7_27_groupi_n_482, csa_tree_add_7_27_groupi_n_483, csa_tree_add_7_27_groupi_n_484, csa_tree_add_7_27_groupi_n_485, csa_tree_add_7_27_groupi_n_486, csa_tree_add_7_27_groupi_n_487, csa_tree_add_7_27_groupi_n_488, csa_tree_add_7_27_groupi_n_489;
  wire csa_tree_add_7_27_groupi_n_490, csa_tree_add_7_27_groupi_n_491, csa_tree_add_7_27_groupi_n_492, csa_tree_add_7_27_groupi_n_493, csa_tree_add_7_27_groupi_n_494, csa_tree_add_7_27_groupi_n_495, csa_tree_add_7_27_groupi_n_496, csa_tree_add_7_27_groupi_n_497;
  wire csa_tree_add_7_27_groupi_n_498, csa_tree_add_7_27_groupi_n_499, csa_tree_add_7_27_groupi_n_500, csa_tree_add_7_27_groupi_n_501, csa_tree_add_7_27_groupi_n_502, csa_tree_add_7_27_groupi_n_503, csa_tree_add_7_27_groupi_n_504, csa_tree_add_7_27_groupi_n_505;
  wire csa_tree_add_7_27_groupi_n_506, csa_tree_add_7_27_groupi_n_507, csa_tree_add_7_27_groupi_n_508, csa_tree_add_7_27_groupi_n_509, csa_tree_add_7_27_groupi_n_510, csa_tree_add_7_27_groupi_n_511, csa_tree_add_7_27_groupi_n_512, csa_tree_add_7_27_groupi_n_513;
  wire csa_tree_add_7_27_groupi_n_514, csa_tree_add_7_27_groupi_n_515, csa_tree_add_7_27_groupi_n_516, csa_tree_add_7_27_groupi_n_517, csa_tree_add_7_27_groupi_n_518, csa_tree_add_7_27_groupi_n_519, csa_tree_add_7_27_groupi_n_520, csa_tree_add_7_27_groupi_n_521;
  wire csa_tree_add_7_27_groupi_n_522, csa_tree_add_7_27_groupi_n_523, csa_tree_add_7_27_groupi_n_524, csa_tree_add_7_27_groupi_n_525, csa_tree_add_7_27_groupi_n_526, csa_tree_add_7_27_groupi_n_527, csa_tree_add_7_27_groupi_n_528, csa_tree_add_7_27_groupi_n_529;
  wire csa_tree_add_7_27_groupi_n_530, csa_tree_add_7_27_groupi_n_531, csa_tree_add_7_27_groupi_n_532, csa_tree_add_7_27_groupi_n_533, csa_tree_add_7_27_groupi_n_534, csa_tree_add_7_27_groupi_n_535, csa_tree_add_7_27_groupi_n_536, csa_tree_add_7_27_groupi_n_537;
  wire csa_tree_add_7_27_groupi_n_538, csa_tree_add_7_27_groupi_n_539, csa_tree_add_7_27_groupi_n_540, csa_tree_add_7_27_groupi_n_541, csa_tree_add_7_27_groupi_n_542, csa_tree_add_7_27_groupi_n_543, csa_tree_add_7_27_groupi_n_544, csa_tree_add_7_27_groupi_n_545;
  wire csa_tree_add_7_27_groupi_n_546, csa_tree_add_7_27_groupi_n_547, csa_tree_add_7_27_groupi_n_548, csa_tree_add_7_27_groupi_n_549, csa_tree_add_7_27_groupi_n_550, csa_tree_add_7_27_groupi_n_551, csa_tree_add_7_27_groupi_n_552, csa_tree_add_7_27_groupi_n_553;
  wire csa_tree_add_7_27_groupi_n_554, csa_tree_add_7_27_groupi_n_555, csa_tree_add_7_27_groupi_n_556, csa_tree_add_7_27_groupi_n_557, csa_tree_add_7_27_groupi_n_558, csa_tree_add_7_27_groupi_n_559, csa_tree_add_7_27_groupi_n_560, csa_tree_add_7_27_groupi_n_561;
  wire csa_tree_add_7_27_groupi_n_562, csa_tree_add_7_27_groupi_n_563, csa_tree_add_7_27_groupi_n_564, csa_tree_add_7_27_groupi_n_565, csa_tree_add_7_27_groupi_n_566, csa_tree_add_7_27_groupi_n_567, csa_tree_add_7_27_groupi_n_568, csa_tree_add_7_27_groupi_n_569;
  wire csa_tree_add_7_27_groupi_n_570, csa_tree_add_7_27_groupi_n_571, csa_tree_add_7_27_groupi_n_572, csa_tree_add_7_27_groupi_n_573, csa_tree_add_7_27_groupi_n_574, csa_tree_add_7_27_groupi_n_575, csa_tree_add_7_27_groupi_n_576, csa_tree_add_7_27_groupi_n_577;
  wire csa_tree_add_7_27_groupi_n_578, csa_tree_add_7_27_groupi_n_579, csa_tree_add_7_27_groupi_n_580, csa_tree_add_7_27_groupi_n_581, csa_tree_add_7_27_groupi_n_582, csa_tree_add_7_27_groupi_n_583, csa_tree_add_7_27_groupi_n_584, csa_tree_add_7_27_groupi_n_585;
  wire csa_tree_add_7_27_groupi_n_586, csa_tree_add_7_27_groupi_n_587, csa_tree_add_7_27_groupi_n_588, csa_tree_add_7_27_groupi_n_589, csa_tree_add_7_27_groupi_n_590, csa_tree_add_7_27_groupi_n_591, csa_tree_add_7_27_groupi_n_592, csa_tree_add_7_27_groupi_n_593;
  wire csa_tree_add_7_27_groupi_n_594, csa_tree_add_7_27_groupi_n_595, csa_tree_add_7_27_groupi_n_596, csa_tree_add_7_27_groupi_n_597, csa_tree_add_7_27_groupi_n_598, csa_tree_add_7_27_groupi_n_599, csa_tree_add_7_27_groupi_n_600, csa_tree_add_7_27_groupi_n_601;
  wire csa_tree_add_7_27_groupi_n_602, csa_tree_add_7_27_groupi_n_603, csa_tree_add_7_27_groupi_n_604, csa_tree_add_7_27_groupi_n_605, csa_tree_add_7_27_groupi_n_606, csa_tree_add_7_27_groupi_n_607, csa_tree_add_7_27_groupi_n_608, csa_tree_add_7_27_groupi_n_609;
  wire csa_tree_add_7_27_groupi_n_610, csa_tree_add_7_27_groupi_n_611, csa_tree_add_7_27_groupi_n_612, csa_tree_add_7_27_groupi_n_613, csa_tree_add_7_27_groupi_n_614, csa_tree_add_7_27_groupi_n_615, csa_tree_add_7_27_groupi_n_616, csa_tree_add_7_27_groupi_n_617;
  wire csa_tree_add_7_27_groupi_n_618, csa_tree_add_7_27_groupi_n_619, csa_tree_add_7_27_groupi_n_620, csa_tree_add_7_27_groupi_n_621, csa_tree_add_7_27_groupi_n_622, csa_tree_add_7_27_groupi_n_623, csa_tree_add_7_27_groupi_n_624, csa_tree_add_7_27_groupi_n_625;
  wire csa_tree_add_7_27_groupi_n_626, csa_tree_add_7_27_groupi_n_627, csa_tree_add_7_27_groupi_n_628, csa_tree_add_7_27_groupi_n_629, csa_tree_add_7_27_groupi_n_630, csa_tree_add_7_27_groupi_n_631, csa_tree_add_7_27_groupi_n_632, csa_tree_add_7_27_groupi_n_633;
  wire csa_tree_add_7_27_groupi_n_634, csa_tree_add_7_27_groupi_n_635, csa_tree_add_7_27_groupi_n_636, csa_tree_add_7_27_groupi_n_637, csa_tree_add_7_27_groupi_n_638, csa_tree_add_7_27_groupi_n_639, csa_tree_add_7_27_groupi_n_640, csa_tree_add_7_27_groupi_n_641;
  wire csa_tree_add_7_27_groupi_n_642, csa_tree_add_7_27_groupi_n_643, csa_tree_add_7_27_groupi_n_644, csa_tree_add_7_27_groupi_n_645, csa_tree_add_7_27_groupi_n_646, csa_tree_add_7_27_groupi_n_647, csa_tree_add_7_27_groupi_n_648, csa_tree_add_7_27_groupi_n_649;
  wire csa_tree_add_7_27_groupi_n_656, csa_tree_add_7_27_groupi_n_657, csa_tree_add_7_27_groupi_n_658, csa_tree_add_7_27_groupi_n_659, csa_tree_add_7_27_groupi_n_660, csa_tree_add_7_27_groupi_n_661, csa_tree_add_7_27_groupi_n_662, csa_tree_add_7_27_groupi_n_663;
  wire csa_tree_add_7_27_groupi_n_664, csa_tree_add_7_27_groupi_n_665, csa_tree_add_7_27_groupi_n_666, csa_tree_add_7_27_groupi_n_667, csa_tree_add_7_27_groupi_n_668, csa_tree_add_7_27_groupi_n_669, csa_tree_add_7_27_groupi_n_670, csa_tree_add_7_27_groupi_n_671;
  wire csa_tree_add_7_27_groupi_n_672, csa_tree_add_7_27_groupi_n_673, csa_tree_add_7_27_groupi_n_674, csa_tree_add_7_27_groupi_n_675, csa_tree_add_7_27_groupi_n_676, csa_tree_add_7_27_groupi_n_677, csa_tree_add_7_27_groupi_n_678, csa_tree_add_7_27_groupi_n_679;
  wire csa_tree_add_7_27_groupi_n_680, csa_tree_add_7_27_groupi_n_681, csa_tree_add_7_27_groupi_n_682, csa_tree_add_7_27_groupi_n_683, csa_tree_add_7_27_groupi_n_684, csa_tree_add_7_27_groupi_n_685, csa_tree_add_7_27_groupi_n_686, csa_tree_add_7_27_groupi_n_687;
  wire csa_tree_add_7_27_groupi_n_688, csa_tree_add_7_27_groupi_n_689, csa_tree_add_7_27_groupi_n_690, csa_tree_add_7_27_groupi_n_691, csa_tree_add_7_27_groupi_n_692, csa_tree_add_7_27_groupi_n_693, csa_tree_add_7_27_groupi_n_694, csa_tree_add_7_27_groupi_n_695;
  wire csa_tree_add_7_27_groupi_n_696, csa_tree_add_7_27_groupi_n_697, csa_tree_add_7_27_groupi_n_698, csa_tree_add_7_27_groupi_n_699, csa_tree_add_7_27_groupi_n_700, csa_tree_add_7_27_groupi_n_701, csa_tree_add_7_27_groupi_n_702, csa_tree_add_7_27_groupi_n_703;
  wire csa_tree_add_7_27_groupi_n_704, csa_tree_add_7_27_groupi_n_705, csa_tree_add_7_27_groupi_n_706, csa_tree_add_7_27_groupi_n_707, csa_tree_add_7_27_groupi_n_708, csa_tree_add_7_27_groupi_n_709, csa_tree_add_7_27_groupi_n_710, csa_tree_add_7_27_groupi_n_711;
  wire csa_tree_add_7_27_groupi_n_712, csa_tree_add_7_27_groupi_n_713, csa_tree_add_7_27_groupi_n_714, csa_tree_add_7_27_groupi_n_715, csa_tree_add_7_27_groupi_n_716, csa_tree_add_7_27_groupi_n_717, csa_tree_add_7_27_groupi_n_718, csa_tree_add_7_27_groupi_n_719;
  wire csa_tree_add_7_27_groupi_n_720, csa_tree_add_7_27_groupi_n_721, csa_tree_add_7_27_groupi_n_722, csa_tree_add_7_27_groupi_n_723, csa_tree_add_7_27_groupi_n_724, csa_tree_add_7_27_groupi_n_725, csa_tree_add_7_27_groupi_n_726, csa_tree_add_7_27_groupi_n_727;
  wire csa_tree_add_7_27_groupi_n_728, csa_tree_add_7_27_groupi_n_729, csa_tree_add_7_27_groupi_n_730, csa_tree_add_7_27_groupi_n_731, csa_tree_add_7_27_groupi_n_732, csa_tree_add_7_27_groupi_n_733, csa_tree_add_7_27_groupi_n_734, csa_tree_add_7_27_groupi_n_735;
  wire csa_tree_add_7_27_groupi_n_736, csa_tree_add_7_27_groupi_n_737, csa_tree_add_7_27_groupi_n_738, csa_tree_add_7_27_groupi_n_739, csa_tree_add_7_27_groupi_n_740, csa_tree_add_7_27_groupi_n_741, csa_tree_add_7_27_groupi_n_742, csa_tree_add_7_27_groupi_n_743;
  wire csa_tree_add_7_27_groupi_n_744, csa_tree_add_7_27_groupi_n_745, csa_tree_add_7_27_groupi_n_746, csa_tree_add_7_27_groupi_n_747, csa_tree_add_7_27_groupi_n_748, csa_tree_add_7_27_groupi_n_749, csa_tree_add_7_27_groupi_n_750, csa_tree_add_7_27_groupi_n_751;
  wire csa_tree_add_7_27_groupi_n_752, csa_tree_add_7_27_groupi_n_753, csa_tree_add_7_27_groupi_n_754, csa_tree_add_7_27_groupi_n_755, csa_tree_add_7_27_groupi_n_756, csa_tree_add_7_27_groupi_n_757, csa_tree_add_7_27_groupi_n_758, csa_tree_add_7_27_groupi_n_759;
  wire csa_tree_add_7_27_groupi_n_760, csa_tree_add_7_27_groupi_n_761, csa_tree_add_7_27_groupi_n_762, csa_tree_add_7_27_groupi_n_763, csa_tree_add_7_27_groupi_n_764, csa_tree_add_7_27_groupi_n_765, csa_tree_add_7_27_groupi_n_766, csa_tree_add_7_27_groupi_n_767;
  wire csa_tree_add_7_27_groupi_n_768, csa_tree_add_7_27_groupi_n_769, csa_tree_add_7_27_groupi_n_770, csa_tree_add_7_27_groupi_n_771, csa_tree_add_7_27_groupi_n_772, csa_tree_add_7_27_groupi_n_773, csa_tree_add_7_27_groupi_n_774, csa_tree_add_7_27_groupi_n_775;
  wire csa_tree_add_7_27_groupi_n_776, csa_tree_add_7_27_groupi_n_777, csa_tree_add_7_27_groupi_n_778, csa_tree_add_7_27_groupi_n_779, csa_tree_add_7_27_groupi_n_780, csa_tree_add_7_27_groupi_n_781, csa_tree_add_7_27_groupi_n_782, csa_tree_add_7_27_groupi_n_783;
  wire csa_tree_add_7_27_groupi_n_784, csa_tree_add_7_27_groupi_n_785, csa_tree_add_7_27_groupi_n_786, csa_tree_add_7_27_groupi_n_787, csa_tree_add_7_27_groupi_n_788, csa_tree_add_7_27_groupi_n_789, csa_tree_add_7_27_groupi_n_790, csa_tree_add_7_27_groupi_n_791;
  wire csa_tree_add_7_27_groupi_n_792, csa_tree_add_7_27_groupi_n_793, csa_tree_add_7_27_groupi_n_795, csa_tree_add_7_27_groupi_n_796, csa_tree_add_7_27_groupi_n_797, csa_tree_add_7_27_groupi_n_798, csa_tree_add_7_27_groupi_n_799, csa_tree_add_7_27_groupi_n_800;
  wire csa_tree_add_7_27_groupi_n_801, csa_tree_add_7_27_groupi_n_802, csa_tree_add_7_27_groupi_n_803, csa_tree_add_7_27_groupi_n_804, csa_tree_add_7_27_groupi_n_805, csa_tree_add_7_27_groupi_n_806, csa_tree_add_7_27_groupi_n_807, csa_tree_add_7_27_groupi_n_808;
  wire csa_tree_add_7_27_groupi_n_809, csa_tree_add_7_27_groupi_n_810, csa_tree_add_7_27_groupi_n_811, csa_tree_add_7_27_groupi_n_812, csa_tree_add_7_27_groupi_n_813, csa_tree_add_7_27_groupi_n_814, csa_tree_add_7_27_groupi_n_815, csa_tree_add_7_27_groupi_n_816;
  wire csa_tree_add_7_27_groupi_n_817, csa_tree_add_7_27_groupi_n_818, csa_tree_add_7_27_groupi_n_819, csa_tree_add_7_27_groupi_n_820, csa_tree_add_7_27_groupi_n_821, csa_tree_add_7_27_groupi_n_822, csa_tree_add_7_27_groupi_n_823, csa_tree_add_7_27_groupi_n_824;
  wire csa_tree_add_7_27_groupi_n_825, csa_tree_add_7_27_groupi_n_826, csa_tree_add_7_27_groupi_n_827, csa_tree_add_7_27_groupi_n_828, csa_tree_add_7_27_groupi_n_829, csa_tree_add_7_27_groupi_n_830, csa_tree_add_7_27_groupi_n_831, csa_tree_add_7_27_groupi_n_832;
  wire csa_tree_add_7_27_groupi_n_833, csa_tree_add_7_27_groupi_n_834, csa_tree_add_7_27_groupi_n_835, csa_tree_add_7_27_groupi_n_836, csa_tree_add_7_27_groupi_n_837, csa_tree_add_7_27_groupi_n_838, csa_tree_add_7_27_groupi_n_839, csa_tree_add_7_27_groupi_n_840;
  wire csa_tree_add_7_27_groupi_n_841, csa_tree_add_7_27_groupi_n_842, csa_tree_add_7_27_groupi_n_843, csa_tree_add_7_27_groupi_n_844, csa_tree_add_7_27_groupi_n_845, csa_tree_add_7_27_groupi_n_846, csa_tree_add_7_27_groupi_n_847, csa_tree_add_7_27_groupi_n_848;
  wire csa_tree_add_7_27_groupi_n_849, csa_tree_add_7_27_groupi_n_850, csa_tree_add_7_27_groupi_n_851, csa_tree_add_7_27_groupi_n_852, csa_tree_add_7_27_groupi_n_853, csa_tree_add_7_27_groupi_n_854, csa_tree_add_7_27_groupi_n_855, csa_tree_add_7_27_groupi_n_856;
  wire csa_tree_add_7_27_groupi_n_857, csa_tree_add_7_27_groupi_n_858, csa_tree_add_7_27_groupi_n_859, csa_tree_add_7_27_groupi_n_860, csa_tree_add_7_27_groupi_n_861, csa_tree_add_7_27_groupi_n_862, csa_tree_add_7_27_groupi_n_863, csa_tree_add_7_27_groupi_n_864;
  wire csa_tree_add_7_27_groupi_n_865, csa_tree_add_7_27_groupi_n_866, csa_tree_add_7_27_groupi_n_867, csa_tree_add_7_27_groupi_n_868, csa_tree_add_7_27_groupi_n_869, csa_tree_add_7_27_groupi_n_870, csa_tree_add_7_27_groupi_n_871, csa_tree_add_7_27_groupi_n_872;
  wire csa_tree_add_7_27_groupi_n_873, csa_tree_add_7_27_groupi_n_874, csa_tree_add_7_27_groupi_n_875, csa_tree_add_7_27_groupi_n_876, csa_tree_add_7_27_groupi_n_877, csa_tree_add_7_27_groupi_n_878, csa_tree_add_7_27_groupi_n_879, csa_tree_add_7_27_groupi_n_880;
  wire csa_tree_add_7_27_groupi_n_881, csa_tree_add_7_27_groupi_n_882, csa_tree_add_7_27_groupi_n_883, csa_tree_add_7_27_groupi_n_884, csa_tree_add_7_27_groupi_n_885, csa_tree_add_7_27_groupi_n_886, csa_tree_add_7_27_groupi_n_887, csa_tree_add_7_27_groupi_n_888;
  wire csa_tree_add_7_27_groupi_n_889, csa_tree_add_7_27_groupi_n_890, csa_tree_add_7_27_groupi_n_891, csa_tree_add_7_27_groupi_n_892, csa_tree_add_7_27_groupi_n_893, csa_tree_add_7_27_groupi_n_894, csa_tree_add_7_27_groupi_n_895, csa_tree_add_7_27_groupi_n_896;
  wire csa_tree_add_7_27_groupi_n_897, csa_tree_add_7_27_groupi_n_898, csa_tree_add_7_27_groupi_n_899, csa_tree_add_7_27_groupi_n_900, csa_tree_add_7_27_groupi_n_901, csa_tree_add_7_27_groupi_n_902, csa_tree_add_7_27_groupi_n_903, csa_tree_add_7_27_groupi_n_904;
  wire csa_tree_add_7_27_groupi_n_905, csa_tree_add_7_27_groupi_n_906, csa_tree_add_7_27_groupi_n_907, csa_tree_add_7_27_groupi_n_908, csa_tree_add_7_27_groupi_n_909, csa_tree_add_7_27_groupi_n_910, csa_tree_add_7_27_groupi_n_911, csa_tree_add_7_27_groupi_n_912;
  wire csa_tree_add_7_27_groupi_n_913, csa_tree_add_7_27_groupi_n_914, csa_tree_add_7_27_groupi_n_915, csa_tree_add_7_27_groupi_n_916, csa_tree_add_7_27_groupi_n_917, csa_tree_add_7_27_groupi_n_918, csa_tree_add_7_27_groupi_n_919, csa_tree_add_7_27_groupi_n_920;
  wire csa_tree_add_7_27_groupi_n_921, csa_tree_add_7_27_groupi_n_922, csa_tree_add_7_27_groupi_n_923, csa_tree_add_7_27_groupi_n_924, csa_tree_add_7_27_groupi_n_925, csa_tree_add_7_27_groupi_n_926, csa_tree_add_7_27_groupi_n_927, csa_tree_add_7_27_groupi_n_928;
  wire csa_tree_add_7_27_groupi_n_929, csa_tree_add_7_27_groupi_n_930, csa_tree_add_7_27_groupi_n_931, csa_tree_add_7_27_groupi_n_932, csa_tree_add_7_27_groupi_n_933, csa_tree_add_7_27_groupi_n_934, csa_tree_add_7_27_groupi_n_935, csa_tree_add_7_27_groupi_n_936;
  wire csa_tree_add_7_27_groupi_n_937, csa_tree_add_7_27_groupi_n_938, csa_tree_add_7_27_groupi_n_939, csa_tree_add_7_27_groupi_n_940, csa_tree_add_7_27_groupi_n_941, csa_tree_add_7_27_groupi_n_942, csa_tree_add_7_27_groupi_n_943, csa_tree_add_7_27_groupi_n_944;
  wire csa_tree_add_7_27_groupi_n_945, csa_tree_add_7_27_groupi_n_946, csa_tree_add_7_27_groupi_n_947, csa_tree_add_7_27_groupi_n_948, csa_tree_add_7_27_groupi_n_949, csa_tree_add_7_27_groupi_n_950, csa_tree_add_7_27_groupi_n_951, csa_tree_add_7_27_groupi_n_952;
  wire csa_tree_add_7_27_groupi_n_953, csa_tree_add_7_27_groupi_n_954, csa_tree_add_7_27_groupi_n_955, csa_tree_add_7_27_groupi_n_956, csa_tree_add_7_27_groupi_n_957, csa_tree_add_7_27_groupi_n_958, csa_tree_add_7_27_groupi_n_959, csa_tree_add_7_27_groupi_n_960;
  wire csa_tree_add_7_27_groupi_n_961, csa_tree_add_7_27_groupi_n_962, csa_tree_add_7_27_groupi_n_963, csa_tree_add_7_27_groupi_n_964, csa_tree_add_7_27_groupi_n_965, csa_tree_add_7_27_groupi_n_966, csa_tree_add_7_27_groupi_n_967, csa_tree_add_7_27_groupi_n_968;
  wire csa_tree_add_7_27_groupi_n_969, csa_tree_add_7_27_groupi_n_970, csa_tree_add_7_27_groupi_n_971, csa_tree_add_7_27_groupi_n_972, csa_tree_add_7_27_groupi_n_973, csa_tree_add_7_27_groupi_n_974, csa_tree_add_7_27_groupi_n_975, csa_tree_add_7_27_groupi_n_976;
  wire csa_tree_add_7_27_groupi_n_977, csa_tree_add_7_27_groupi_n_978, csa_tree_add_7_27_groupi_n_979, csa_tree_add_7_27_groupi_n_980, csa_tree_add_7_27_groupi_n_981, csa_tree_add_7_27_groupi_n_982, csa_tree_add_7_27_groupi_n_983, csa_tree_add_7_27_groupi_n_984;
  wire csa_tree_add_7_27_groupi_n_985, csa_tree_add_7_27_groupi_n_986, csa_tree_add_7_27_groupi_n_987, csa_tree_add_7_27_groupi_n_988, csa_tree_add_7_27_groupi_n_989, csa_tree_add_7_27_groupi_n_990, csa_tree_add_7_27_groupi_n_991, csa_tree_add_7_27_groupi_n_992;
  wire csa_tree_add_7_27_groupi_n_993, csa_tree_add_7_27_groupi_n_994, csa_tree_add_7_27_groupi_n_995, csa_tree_add_7_27_groupi_n_996, csa_tree_add_7_27_groupi_n_997, csa_tree_add_7_27_groupi_n_998, csa_tree_add_7_27_groupi_n_999, csa_tree_add_7_27_groupi_n_1000;
  wire csa_tree_add_7_27_groupi_n_1001, csa_tree_add_7_27_groupi_n_1002, csa_tree_add_7_27_groupi_n_1003, csa_tree_add_7_27_groupi_n_1004, csa_tree_add_7_27_groupi_n_1005, csa_tree_add_7_27_groupi_n_1006, csa_tree_add_7_27_groupi_n_1007, csa_tree_add_7_27_groupi_n_1008;
  wire csa_tree_add_7_27_groupi_n_1009, csa_tree_add_7_27_groupi_n_1010, csa_tree_add_7_27_groupi_n_1011, csa_tree_add_7_27_groupi_n_1012, csa_tree_add_7_27_groupi_n_1013, csa_tree_add_7_27_groupi_n_1014, csa_tree_add_7_27_groupi_n_1015, csa_tree_add_7_27_groupi_n_1016;
  wire csa_tree_add_7_27_groupi_n_1017, csa_tree_add_7_27_groupi_n_1018, csa_tree_add_7_27_groupi_n_1019, csa_tree_add_7_27_groupi_n_1020, csa_tree_add_7_27_groupi_n_1021, csa_tree_add_7_27_groupi_n_1022, csa_tree_add_7_27_groupi_n_1023, csa_tree_add_7_27_groupi_n_1024;
  wire csa_tree_add_7_27_groupi_n_1025, csa_tree_add_7_27_groupi_n_1026, csa_tree_add_7_27_groupi_n_1027, csa_tree_add_7_27_groupi_n_1028, csa_tree_add_7_27_groupi_n_1029, csa_tree_add_7_27_groupi_n_1030, csa_tree_add_7_27_groupi_n_1031, csa_tree_add_7_27_groupi_n_1032;
  wire csa_tree_add_7_27_groupi_n_1033, csa_tree_add_7_27_groupi_n_1034, csa_tree_add_7_27_groupi_n_1035, csa_tree_add_7_27_groupi_n_1036, csa_tree_add_7_27_groupi_n_1037, csa_tree_add_7_27_groupi_n_1038, csa_tree_add_7_27_groupi_n_1039, csa_tree_add_7_27_groupi_n_1040;
  wire csa_tree_add_7_27_groupi_n_1041, csa_tree_add_7_27_groupi_n_1042, csa_tree_add_7_27_groupi_n_1043, csa_tree_add_7_27_groupi_n_1044, csa_tree_add_7_27_groupi_n_1045, csa_tree_add_7_27_groupi_n_1046, csa_tree_add_7_27_groupi_n_1047, csa_tree_add_7_27_groupi_n_1048;
  wire csa_tree_add_7_27_groupi_n_1049, csa_tree_add_7_27_groupi_n_1050, csa_tree_add_7_27_groupi_n_1051, csa_tree_add_7_27_groupi_n_1052, csa_tree_add_7_27_groupi_n_1053, csa_tree_add_7_27_groupi_n_1054, csa_tree_add_7_27_groupi_n_1055, csa_tree_add_7_27_groupi_n_1056;
  wire csa_tree_add_7_27_groupi_n_1057, csa_tree_add_7_27_groupi_n_1058, csa_tree_add_7_27_groupi_n_1059, csa_tree_add_7_27_groupi_n_1060, csa_tree_add_7_27_groupi_n_1061, csa_tree_add_7_27_groupi_n_1062, csa_tree_add_7_27_groupi_n_1063, csa_tree_add_7_27_groupi_n_1064;
  wire csa_tree_add_7_27_groupi_n_1065, csa_tree_add_7_27_groupi_n_1066, csa_tree_add_7_27_groupi_n_1067, csa_tree_add_7_27_groupi_n_1068, csa_tree_add_7_27_groupi_n_1069, csa_tree_add_7_27_groupi_n_1070, csa_tree_add_7_27_groupi_n_1071, csa_tree_add_7_27_groupi_n_1072;
  wire csa_tree_add_7_27_groupi_n_1073, csa_tree_add_7_27_groupi_n_1074, csa_tree_add_7_27_groupi_n_1075, csa_tree_add_7_27_groupi_n_1076, csa_tree_add_7_27_groupi_n_1077, csa_tree_add_7_27_groupi_n_1078, csa_tree_add_7_27_groupi_n_1079, csa_tree_add_7_27_groupi_n_1080;
  wire csa_tree_add_7_27_groupi_n_1081, csa_tree_add_7_27_groupi_n_1082, csa_tree_add_7_27_groupi_n_1083, csa_tree_add_7_27_groupi_n_1084, csa_tree_add_7_27_groupi_n_1085, csa_tree_add_7_27_groupi_n_1086, csa_tree_add_7_27_groupi_n_1087, csa_tree_add_7_27_groupi_n_1088;
  wire csa_tree_add_7_27_groupi_n_1089, csa_tree_add_7_27_groupi_n_1090, csa_tree_add_7_27_groupi_n_1091, csa_tree_add_7_27_groupi_n_1092, csa_tree_add_7_27_groupi_n_1093, csa_tree_add_7_27_groupi_n_1094, csa_tree_add_7_27_groupi_n_1095, csa_tree_add_7_27_groupi_n_1096;
  wire csa_tree_add_7_27_groupi_n_1097, csa_tree_add_7_27_groupi_n_1098, csa_tree_add_7_27_groupi_n_1099, csa_tree_add_7_27_groupi_n_1100, csa_tree_add_7_27_groupi_n_1101, csa_tree_add_7_27_groupi_n_1102, csa_tree_add_7_27_groupi_n_1103, csa_tree_add_7_27_groupi_n_1104;
  wire csa_tree_add_7_27_groupi_n_1105, csa_tree_add_7_27_groupi_n_1106, csa_tree_add_7_27_groupi_n_1107, csa_tree_add_7_27_groupi_n_1108, csa_tree_add_7_27_groupi_n_1109, csa_tree_add_7_27_groupi_n_1110, csa_tree_add_7_27_groupi_n_1111, csa_tree_add_7_27_groupi_n_1112;
  wire csa_tree_add_7_27_groupi_n_1113, csa_tree_add_7_27_groupi_n_1114, csa_tree_add_7_27_groupi_n_1115, csa_tree_add_7_27_groupi_n_1116, csa_tree_add_7_27_groupi_n_1117, csa_tree_add_7_27_groupi_n_1118, csa_tree_add_7_27_groupi_n_1119, csa_tree_add_7_27_groupi_n_1120;
  wire csa_tree_add_7_27_groupi_n_1121, csa_tree_add_7_27_groupi_n_1122, csa_tree_add_7_27_groupi_n_1123, csa_tree_add_7_27_groupi_n_1124, csa_tree_add_7_27_groupi_n_1125, csa_tree_add_7_27_groupi_n_1126, csa_tree_add_7_27_groupi_n_1127, csa_tree_add_7_27_groupi_n_1128;
  wire csa_tree_add_7_27_groupi_n_1129, csa_tree_add_7_27_groupi_n_1130, csa_tree_add_7_27_groupi_n_1131, csa_tree_add_7_27_groupi_n_1132, csa_tree_add_7_27_groupi_n_1133, csa_tree_add_7_27_groupi_n_1134, csa_tree_add_7_27_groupi_n_1135, csa_tree_add_7_27_groupi_n_1136;
  wire csa_tree_add_7_27_groupi_n_1137, csa_tree_add_7_27_groupi_n_1138, csa_tree_add_7_27_groupi_n_1139, csa_tree_add_7_27_groupi_n_1140, csa_tree_add_7_27_groupi_n_1141, csa_tree_add_7_27_groupi_n_1142, csa_tree_add_7_27_groupi_n_1143, csa_tree_add_7_27_groupi_n_1144;
  wire csa_tree_add_7_27_groupi_n_1145, csa_tree_add_7_27_groupi_n_1146, csa_tree_add_7_27_groupi_n_1147, csa_tree_add_7_27_groupi_n_1148, csa_tree_add_7_27_groupi_n_1149, csa_tree_add_7_27_groupi_n_1150, csa_tree_add_7_27_groupi_n_1151, csa_tree_add_7_27_groupi_n_1152;
  wire csa_tree_add_7_27_groupi_n_1153, csa_tree_add_7_27_groupi_n_1154, csa_tree_add_7_27_groupi_n_1155, csa_tree_add_7_27_groupi_n_1156, csa_tree_add_7_27_groupi_n_1157, csa_tree_add_7_27_groupi_n_1158, csa_tree_add_7_27_groupi_n_1159, csa_tree_add_7_27_groupi_n_1160;
  wire csa_tree_add_7_27_groupi_n_1161, csa_tree_add_7_27_groupi_n_1162, csa_tree_add_7_27_groupi_n_1163, csa_tree_add_7_27_groupi_n_1164, csa_tree_add_7_27_groupi_n_1165, csa_tree_add_7_27_groupi_n_1166, csa_tree_add_7_27_groupi_n_1167, csa_tree_add_7_27_groupi_n_1168;
  wire csa_tree_add_7_27_groupi_n_1169, csa_tree_add_7_27_groupi_n_1170, csa_tree_add_7_27_groupi_n_1171, csa_tree_add_7_27_groupi_n_1172, csa_tree_add_7_27_groupi_n_1173, csa_tree_add_7_27_groupi_n_1174, csa_tree_add_7_27_groupi_n_1175, csa_tree_add_7_27_groupi_n_1176;
  wire csa_tree_add_7_27_groupi_n_1177, csa_tree_add_7_27_groupi_n_1178, csa_tree_add_7_27_groupi_n_1179, csa_tree_add_7_27_groupi_n_1180, csa_tree_add_7_27_groupi_n_1181, csa_tree_add_7_27_groupi_n_1182, csa_tree_add_7_27_groupi_n_1183, csa_tree_add_7_27_groupi_n_1184;
  wire csa_tree_add_7_27_groupi_n_1185, csa_tree_add_7_27_groupi_n_1186, csa_tree_add_7_27_groupi_n_1187, csa_tree_add_7_27_groupi_n_1188, csa_tree_add_7_27_groupi_n_1189, csa_tree_add_7_27_groupi_n_1190, csa_tree_add_7_27_groupi_n_1191, csa_tree_add_7_27_groupi_n_1192;
  wire csa_tree_add_7_27_groupi_n_1193, csa_tree_add_7_27_groupi_n_1194, csa_tree_add_7_27_groupi_n_1195, csa_tree_add_7_27_groupi_n_1196, csa_tree_add_7_27_groupi_n_1197, csa_tree_add_7_27_groupi_n_1198, csa_tree_add_7_27_groupi_n_1199, csa_tree_add_7_27_groupi_n_1200;
  wire csa_tree_add_7_27_groupi_n_1201, csa_tree_add_7_27_groupi_n_1202, csa_tree_add_7_27_groupi_n_1203, csa_tree_add_7_27_groupi_n_1204, csa_tree_add_7_27_groupi_n_1205, csa_tree_add_7_27_groupi_n_1206, csa_tree_add_7_27_groupi_n_1207, csa_tree_add_7_27_groupi_n_1208;
  wire csa_tree_add_7_27_groupi_n_1209, csa_tree_add_7_27_groupi_n_1210, csa_tree_add_7_27_groupi_n_1211, csa_tree_add_7_27_groupi_n_1212, csa_tree_add_7_27_groupi_n_1213, csa_tree_add_7_27_groupi_n_1214, csa_tree_add_7_27_groupi_n_1215, csa_tree_add_7_27_groupi_n_1216;
  wire csa_tree_add_7_27_groupi_n_1217, csa_tree_add_7_27_groupi_n_1218, csa_tree_add_7_27_groupi_n_1219, csa_tree_add_7_27_groupi_n_1220, csa_tree_add_7_27_groupi_n_1221, csa_tree_add_7_27_groupi_n_1222, csa_tree_add_7_27_groupi_n_1223, csa_tree_add_7_27_groupi_n_1224;
  wire csa_tree_add_7_27_groupi_n_1225, csa_tree_add_7_27_groupi_n_1226, csa_tree_add_7_27_groupi_n_1227, csa_tree_add_7_27_groupi_n_1228, csa_tree_add_7_27_groupi_n_1229, csa_tree_add_7_27_groupi_n_1230, csa_tree_add_7_27_groupi_n_1231, csa_tree_add_7_27_groupi_n_1232;
  wire csa_tree_add_7_27_groupi_n_1233, csa_tree_add_7_27_groupi_n_1234, csa_tree_add_7_27_groupi_n_1235, csa_tree_add_7_27_groupi_n_1236, csa_tree_add_7_27_groupi_n_1237, csa_tree_add_7_27_groupi_n_1238, csa_tree_add_7_27_groupi_n_1239, csa_tree_add_7_27_groupi_n_1240;
  wire csa_tree_add_7_27_groupi_n_1241, csa_tree_add_7_27_groupi_n_1242, csa_tree_add_7_27_groupi_n_1243, csa_tree_add_7_27_groupi_n_1244, csa_tree_add_7_27_groupi_n_1245, csa_tree_add_7_27_groupi_n_1246, csa_tree_add_7_27_groupi_n_1247, csa_tree_add_7_27_groupi_n_1248;
  wire csa_tree_add_7_27_groupi_n_1249, csa_tree_add_7_27_groupi_n_1250, csa_tree_add_7_27_groupi_n_1251, csa_tree_add_7_27_groupi_n_1252, csa_tree_add_7_27_groupi_n_1253, csa_tree_add_7_27_groupi_n_1254, csa_tree_add_7_27_groupi_n_1255, csa_tree_add_7_27_groupi_n_1256;
  wire csa_tree_add_7_27_groupi_n_1257, csa_tree_add_7_27_groupi_n_1258, csa_tree_add_7_27_groupi_n_1259, csa_tree_add_7_27_groupi_n_1260, csa_tree_add_7_27_groupi_n_1261, csa_tree_add_7_27_groupi_n_1262, csa_tree_add_7_27_groupi_n_1263, csa_tree_add_7_27_groupi_n_1264;
  wire csa_tree_add_7_27_groupi_n_1265, csa_tree_add_7_27_groupi_n_1266, csa_tree_add_7_27_groupi_n_1267, csa_tree_add_7_27_groupi_n_1268, csa_tree_add_7_27_groupi_n_1269, csa_tree_add_7_27_groupi_n_1270, csa_tree_add_7_27_groupi_n_1271, csa_tree_add_7_27_groupi_n_1272;
  wire csa_tree_add_7_27_groupi_n_1273, csa_tree_add_7_27_groupi_n_1274, csa_tree_add_7_27_groupi_n_1275, csa_tree_add_7_27_groupi_n_1276, csa_tree_add_7_27_groupi_n_1277, csa_tree_add_7_27_groupi_n_1278, csa_tree_add_7_27_groupi_n_1279, csa_tree_add_7_27_groupi_n_1280;
  wire csa_tree_add_7_27_groupi_n_1281, csa_tree_add_7_27_groupi_n_1282, csa_tree_add_7_27_groupi_n_1283, csa_tree_add_7_27_groupi_n_1284, csa_tree_add_7_27_groupi_n_1285, csa_tree_add_7_27_groupi_n_1286, csa_tree_add_7_27_groupi_n_1287, csa_tree_add_7_27_groupi_n_1288;
  wire csa_tree_add_7_27_groupi_n_1289, csa_tree_add_7_27_groupi_n_1290, csa_tree_add_7_27_groupi_n_1291, csa_tree_add_7_27_groupi_n_1292, csa_tree_add_7_27_groupi_n_1293, csa_tree_add_7_27_groupi_n_1294, csa_tree_add_7_27_groupi_n_1295, csa_tree_add_7_27_groupi_n_1296;
  wire csa_tree_add_7_27_groupi_n_1297, csa_tree_add_7_27_groupi_n_1298, csa_tree_add_7_27_groupi_n_1299, csa_tree_add_7_27_groupi_n_1300, csa_tree_add_7_27_groupi_n_1301, csa_tree_add_7_27_groupi_n_1302, csa_tree_add_7_27_groupi_n_1303, csa_tree_add_7_27_groupi_n_1304;
  wire csa_tree_add_7_27_groupi_n_1305, csa_tree_add_7_27_groupi_n_1306, csa_tree_add_7_27_groupi_n_1307, csa_tree_add_7_27_groupi_n_1308, csa_tree_add_7_27_groupi_n_1309, csa_tree_add_7_27_groupi_n_1310, csa_tree_add_7_27_groupi_n_1311, csa_tree_add_7_27_groupi_n_1312;
  wire csa_tree_add_7_27_groupi_n_1313, csa_tree_add_7_27_groupi_n_1314, csa_tree_add_7_27_groupi_n_1315, csa_tree_add_7_27_groupi_n_1316, csa_tree_add_7_27_groupi_n_1317, csa_tree_add_7_27_groupi_n_1318, csa_tree_add_7_27_groupi_n_1319, csa_tree_add_7_27_groupi_n_1320;
  wire csa_tree_add_7_27_groupi_n_1321, csa_tree_add_7_27_groupi_n_1322, csa_tree_add_7_27_groupi_n_1323, csa_tree_add_7_27_groupi_n_1324, csa_tree_add_7_27_groupi_n_1325, csa_tree_add_7_27_groupi_n_1326, csa_tree_add_7_27_groupi_n_1327, csa_tree_add_7_27_groupi_n_1328;
  wire csa_tree_add_7_27_groupi_n_1329, csa_tree_add_7_27_groupi_n_1330, csa_tree_add_7_27_groupi_n_1331, csa_tree_add_7_27_groupi_n_1332, csa_tree_add_7_27_groupi_n_1333, csa_tree_add_7_27_groupi_n_1334, csa_tree_add_7_27_groupi_n_1335, csa_tree_add_7_27_groupi_n_1336;
  wire csa_tree_add_7_27_groupi_n_1337, csa_tree_add_7_27_groupi_n_1338, csa_tree_add_7_27_groupi_n_1339, csa_tree_add_7_27_groupi_n_1340, csa_tree_add_7_27_groupi_n_1341, csa_tree_add_7_27_groupi_n_1342, csa_tree_add_7_27_groupi_n_1343, csa_tree_add_7_27_groupi_n_1344;
  wire csa_tree_add_7_27_groupi_n_1345, csa_tree_add_7_27_groupi_n_1346, csa_tree_add_7_27_groupi_n_1347, csa_tree_add_7_27_groupi_n_1348, csa_tree_add_7_27_groupi_n_1349, csa_tree_add_7_27_groupi_n_1350, csa_tree_add_7_27_groupi_n_1351, csa_tree_add_7_27_groupi_n_1352;
  wire csa_tree_add_7_27_groupi_n_1353, csa_tree_add_7_27_groupi_n_1354, csa_tree_add_7_27_groupi_n_1355, csa_tree_add_7_27_groupi_n_1356, csa_tree_add_7_27_groupi_n_1357, csa_tree_add_7_27_groupi_n_1358, csa_tree_add_7_27_groupi_n_1359, csa_tree_add_7_27_groupi_n_1360;
  wire csa_tree_add_7_27_groupi_n_1361, csa_tree_add_7_27_groupi_n_1362, csa_tree_add_7_27_groupi_n_1363, csa_tree_add_7_27_groupi_n_1364, csa_tree_add_7_27_groupi_n_1365, csa_tree_add_7_27_groupi_n_1366, csa_tree_add_7_27_groupi_n_1367, csa_tree_add_7_27_groupi_n_1368;
  wire csa_tree_add_7_27_groupi_n_1369, csa_tree_add_7_27_groupi_n_1370, csa_tree_add_7_27_groupi_n_1371, csa_tree_add_7_27_groupi_n_1372, csa_tree_add_7_27_groupi_n_1373, csa_tree_add_7_27_groupi_n_1374, csa_tree_add_7_27_groupi_n_1375, csa_tree_add_7_27_groupi_n_1376;
  wire csa_tree_add_7_27_groupi_n_1377, csa_tree_add_7_27_groupi_n_1378, csa_tree_add_7_27_groupi_n_1379, csa_tree_add_7_27_groupi_n_1380, csa_tree_add_7_27_groupi_n_1381, csa_tree_add_7_27_groupi_n_1382, csa_tree_add_7_27_groupi_n_1383, csa_tree_add_7_27_groupi_n_1384;
  wire csa_tree_add_7_27_groupi_n_1385, csa_tree_add_7_27_groupi_n_1386, csa_tree_add_7_27_groupi_n_1387, csa_tree_add_7_27_groupi_n_1388, csa_tree_add_7_27_groupi_n_1389, csa_tree_add_7_27_groupi_n_1390, csa_tree_add_7_27_groupi_n_1391, csa_tree_add_7_27_groupi_n_1392;
  wire csa_tree_add_7_27_groupi_n_1393, csa_tree_add_7_27_groupi_n_1394, csa_tree_add_7_27_groupi_n_1395, csa_tree_add_7_27_groupi_n_1396, csa_tree_add_7_27_groupi_n_1397, csa_tree_add_7_27_groupi_n_1398, csa_tree_add_7_27_groupi_n_1399, csa_tree_add_7_27_groupi_n_1400;
  wire csa_tree_add_7_27_groupi_n_1401, csa_tree_add_7_27_groupi_n_1402, csa_tree_add_7_27_groupi_n_1403, csa_tree_add_7_27_groupi_n_1404, csa_tree_add_7_27_groupi_n_1405, csa_tree_add_7_27_groupi_n_1406, csa_tree_add_7_27_groupi_n_1407, csa_tree_add_7_27_groupi_n_1408;
  wire csa_tree_add_7_27_groupi_n_1409, csa_tree_add_7_27_groupi_n_1410, csa_tree_add_7_27_groupi_n_1411, csa_tree_add_7_27_groupi_n_1412, csa_tree_add_7_27_groupi_n_1413, csa_tree_add_7_27_groupi_n_1414, csa_tree_add_7_27_groupi_n_1415, csa_tree_add_7_27_groupi_n_1416;
  wire csa_tree_add_7_27_groupi_n_1417, csa_tree_add_7_27_groupi_n_1418, csa_tree_add_7_27_groupi_n_1419, csa_tree_add_7_27_groupi_n_1420, csa_tree_add_7_27_groupi_n_1421, csa_tree_add_7_27_groupi_n_1422, csa_tree_add_7_27_groupi_n_1423, csa_tree_add_7_27_groupi_n_1424;
  wire csa_tree_add_7_27_groupi_n_1425, csa_tree_add_7_27_groupi_n_1426, csa_tree_add_7_27_groupi_n_1427, csa_tree_add_7_27_groupi_n_1428, csa_tree_add_7_27_groupi_n_1429, csa_tree_add_7_27_groupi_n_1430, csa_tree_add_7_27_groupi_n_1431, csa_tree_add_7_27_groupi_n_1432;
  wire csa_tree_add_7_27_groupi_n_1433, csa_tree_add_7_27_groupi_n_1434, csa_tree_add_7_27_groupi_n_1435, csa_tree_add_7_27_groupi_n_1436, csa_tree_add_7_27_groupi_n_1437, csa_tree_add_7_27_groupi_n_1438, csa_tree_add_7_27_groupi_n_1439, csa_tree_add_7_27_groupi_n_1440;
  wire csa_tree_add_7_27_groupi_n_1441, csa_tree_add_7_27_groupi_n_1442, csa_tree_add_7_27_groupi_n_1443, csa_tree_add_7_27_groupi_n_1444, csa_tree_add_7_27_groupi_n_1445, csa_tree_add_7_27_groupi_n_1446, csa_tree_add_7_27_groupi_n_1447, csa_tree_add_7_27_groupi_n_1448;
  wire csa_tree_add_7_27_groupi_n_1449, csa_tree_add_7_27_groupi_n_1450, csa_tree_add_7_27_groupi_n_1451, csa_tree_add_7_27_groupi_n_1452, csa_tree_add_7_27_groupi_n_1453, csa_tree_add_7_27_groupi_n_1454, csa_tree_add_7_27_groupi_n_1455, csa_tree_add_7_27_groupi_n_1456;
  wire csa_tree_add_7_27_groupi_n_1457, csa_tree_add_7_27_groupi_n_1458, csa_tree_add_7_27_groupi_n_1459, csa_tree_add_7_27_groupi_n_1460, csa_tree_add_7_27_groupi_n_1461, csa_tree_add_7_27_groupi_n_1462, csa_tree_add_7_27_groupi_n_1463, csa_tree_add_7_27_groupi_n_1464;
  wire csa_tree_add_7_27_groupi_n_1465, csa_tree_add_7_27_groupi_n_1466, csa_tree_add_7_27_groupi_n_1467, csa_tree_add_7_27_groupi_n_1468, csa_tree_add_7_27_groupi_n_1469, csa_tree_add_7_27_groupi_n_1470, csa_tree_add_7_27_groupi_n_1471, csa_tree_add_7_27_groupi_n_1472;
  wire csa_tree_add_7_27_groupi_n_1473, csa_tree_add_7_27_groupi_n_1474, csa_tree_add_7_27_groupi_n_1475, csa_tree_add_7_27_groupi_n_1476, csa_tree_add_7_27_groupi_n_1477, csa_tree_add_7_27_groupi_n_1478, csa_tree_add_7_27_groupi_n_1479, csa_tree_add_7_27_groupi_n_1480;
  wire csa_tree_add_7_27_groupi_n_1481, csa_tree_add_7_27_groupi_n_1482, csa_tree_add_7_27_groupi_n_1483, csa_tree_add_7_27_groupi_n_1484, csa_tree_add_7_27_groupi_n_1485, csa_tree_add_7_27_groupi_n_1486, csa_tree_add_7_27_groupi_n_1487, csa_tree_add_7_27_groupi_n_1488;
  wire csa_tree_add_7_27_groupi_n_1489, csa_tree_add_7_27_groupi_n_1490, csa_tree_add_7_27_groupi_n_1491, csa_tree_add_7_27_groupi_n_1492, csa_tree_add_7_27_groupi_n_1493, csa_tree_add_7_27_groupi_n_1494, csa_tree_add_7_27_groupi_n_1495, csa_tree_add_7_27_groupi_n_1496;
  wire csa_tree_add_7_27_groupi_n_1497, csa_tree_add_7_27_groupi_n_1498, csa_tree_add_7_27_groupi_n_1499, csa_tree_add_7_27_groupi_n_1500, csa_tree_add_7_27_groupi_n_1501, csa_tree_add_7_27_groupi_n_1502, csa_tree_add_7_27_groupi_n_1503, csa_tree_add_7_27_groupi_n_1504;
  wire csa_tree_add_7_27_groupi_n_1505, csa_tree_add_7_27_groupi_n_1506, csa_tree_add_7_27_groupi_n_1507, csa_tree_add_7_27_groupi_n_1508, csa_tree_add_7_27_groupi_n_1509, csa_tree_add_7_27_groupi_n_1510, csa_tree_add_7_27_groupi_n_1511, csa_tree_add_7_27_groupi_n_1512;
  wire csa_tree_add_7_27_groupi_n_1513, csa_tree_add_7_27_groupi_n_1514, csa_tree_add_7_27_groupi_n_1515, csa_tree_add_7_27_groupi_n_1516, csa_tree_add_7_27_groupi_n_1517, csa_tree_add_7_27_groupi_n_1518, csa_tree_add_7_27_groupi_n_1519, csa_tree_add_7_27_groupi_n_1520;
  wire csa_tree_add_7_27_groupi_n_1521, csa_tree_add_7_27_groupi_n_1522, csa_tree_add_7_27_groupi_n_1523, csa_tree_add_7_27_groupi_n_1524, csa_tree_add_7_27_groupi_n_1525, csa_tree_add_7_27_groupi_n_1526, csa_tree_add_7_27_groupi_n_1527, csa_tree_add_7_27_groupi_n_1528;
  wire csa_tree_add_7_27_groupi_n_1529, csa_tree_add_7_27_groupi_n_1530, csa_tree_add_7_27_groupi_n_1531, csa_tree_add_7_27_groupi_n_1532, csa_tree_add_7_27_groupi_n_1533, csa_tree_add_7_27_groupi_n_1534, csa_tree_add_7_27_groupi_n_1535, csa_tree_add_7_27_groupi_n_1536;
  wire csa_tree_add_7_27_groupi_n_1537, csa_tree_add_7_27_groupi_n_1538, csa_tree_add_7_27_groupi_n_1539, csa_tree_add_7_27_groupi_n_1540, csa_tree_add_7_27_groupi_n_1541, csa_tree_add_7_27_groupi_n_1542, csa_tree_add_7_27_groupi_n_1543, csa_tree_add_7_27_groupi_n_1544;
  wire csa_tree_add_7_27_groupi_n_1545, csa_tree_add_7_27_groupi_n_1546, csa_tree_add_7_27_groupi_n_1547, csa_tree_add_7_27_groupi_n_1548, csa_tree_add_7_27_groupi_n_1549, csa_tree_add_7_27_groupi_n_1550, csa_tree_add_7_27_groupi_n_1551, csa_tree_add_7_27_groupi_n_1552;
  wire csa_tree_add_7_27_groupi_n_1553, csa_tree_add_7_27_groupi_n_1554, csa_tree_add_7_27_groupi_n_1555, csa_tree_add_7_27_groupi_n_1556, csa_tree_add_7_27_groupi_n_1557, csa_tree_add_7_27_groupi_n_1558, csa_tree_add_7_27_groupi_n_1559, csa_tree_add_7_27_groupi_n_1561;
  wire csa_tree_add_7_27_groupi_n_1562, csa_tree_add_7_27_groupi_n_1563, csa_tree_add_7_27_groupi_n_1564, csa_tree_add_7_27_groupi_n_1565, csa_tree_add_7_27_groupi_n_1566, csa_tree_add_7_27_groupi_n_1567, csa_tree_add_7_27_groupi_n_1568, csa_tree_add_7_27_groupi_n_1569;
  wire csa_tree_add_7_27_groupi_n_1570, csa_tree_add_7_27_groupi_n_1571, csa_tree_add_7_27_groupi_n_1572, csa_tree_add_7_27_groupi_n_1573, csa_tree_add_7_27_groupi_n_1574, csa_tree_add_7_27_groupi_n_1575, csa_tree_add_7_27_groupi_n_1576, csa_tree_add_7_27_groupi_n_1577;
  wire csa_tree_add_7_27_groupi_n_1578, csa_tree_add_7_27_groupi_n_1579, csa_tree_add_7_27_groupi_n_1580, csa_tree_add_7_27_groupi_n_1581, csa_tree_add_7_27_groupi_n_1582, csa_tree_add_7_27_groupi_n_1583, csa_tree_add_7_27_groupi_n_1584, csa_tree_add_7_27_groupi_n_1585;
  wire csa_tree_add_7_27_groupi_n_1586, csa_tree_add_7_27_groupi_n_1587, csa_tree_add_7_27_groupi_n_1588, csa_tree_add_7_27_groupi_n_1589, csa_tree_add_7_27_groupi_n_1590, csa_tree_add_7_27_groupi_n_1591, csa_tree_add_7_27_groupi_n_1592, csa_tree_add_7_27_groupi_n_1593;
  wire csa_tree_add_7_27_groupi_n_1594, csa_tree_add_7_27_groupi_n_1595, csa_tree_add_7_27_groupi_n_1596, csa_tree_add_7_27_groupi_n_1597, csa_tree_add_7_27_groupi_n_1598, csa_tree_add_7_27_groupi_n_1599, csa_tree_add_7_27_groupi_n_1600, csa_tree_add_7_27_groupi_n_1601;
  wire csa_tree_add_7_27_groupi_n_1602, csa_tree_add_7_27_groupi_n_1603, csa_tree_add_7_27_groupi_n_1604, csa_tree_add_7_27_groupi_n_1605, csa_tree_add_7_27_groupi_n_1606, csa_tree_add_7_27_groupi_n_1607, csa_tree_add_7_27_groupi_n_1608, csa_tree_add_7_27_groupi_n_1609;
  wire csa_tree_add_7_27_groupi_n_1610, csa_tree_add_7_27_groupi_n_1611, csa_tree_add_7_27_groupi_n_1612, csa_tree_add_7_27_groupi_n_1613, csa_tree_add_7_27_groupi_n_1614, csa_tree_add_7_27_groupi_n_1615, csa_tree_add_7_27_groupi_n_1616, csa_tree_add_7_27_groupi_n_1617;
  wire csa_tree_add_7_27_groupi_n_1619, csa_tree_add_7_27_groupi_n_1620, csa_tree_add_7_27_groupi_n_1621, csa_tree_add_7_27_groupi_n_1622, csa_tree_add_7_27_groupi_n_1623, csa_tree_add_7_27_groupi_n_1624, csa_tree_add_7_27_groupi_n_1625, csa_tree_add_7_27_groupi_n_1626;
  wire csa_tree_add_7_27_groupi_n_1627, csa_tree_add_7_27_groupi_n_1628, csa_tree_add_7_27_groupi_n_1629, csa_tree_add_7_27_groupi_n_1630, csa_tree_add_7_27_groupi_n_1631, csa_tree_add_7_27_groupi_n_1632, csa_tree_add_7_27_groupi_n_1633, csa_tree_add_7_27_groupi_n_1634;
  wire csa_tree_add_7_27_groupi_n_1635, csa_tree_add_7_27_groupi_n_1636, csa_tree_add_7_27_groupi_n_1637, csa_tree_add_7_27_groupi_n_1638, csa_tree_add_7_27_groupi_n_1639, csa_tree_add_7_27_groupi_n_1640, csa_tree_add_7_27_groupi_n_1641, csa_tree_add_7_27_groupi_n_1642;
  wire csa_tree_add_7_27_groupi_n_1643, csa_tree_add_7_27_groupi_n_1644, csa_tree_add_7_27_groupi_n_1645, csa_tree_add_7_27_groupi_n_1646, csa_tree_add_7_27_groupi_n_1647, csa_tree_add_7_27_groupi_n_1648, csa_tree_add_7_27_groupi_n_1649, csa_tree_add_7_27_groupi_n_1650;
  wire csa_tree_add_7_27_groupi_n_1651, csa_tree_add_7_27_groupi_n_1652, csa_tree_add_7_27_groupi_n_1653, csa_tree_add_7_27_groupi_n_1654, csa_tree_add_7_27_groupi_n_1655, csa_tree_add_7_27_groupi_n_1656, csa_tree_add_7_27_groupi_n_1657, csa_tree_add_7_27_groupi_n_1658;
  wire csa_tree_add_7_27_groupi_n_1659, csa_tree_add_7_27_groupi_n_1660, csa_tree_add_7_27_groupi_n_1661, csa_tree_add_7_27_groupi_n_1662, csa_tree_add_7_27_groupi_n_1663, csa_tree_add_7_27_groupi_n_1664, csa_tree_add_7_27_groupi_n_1665, csa_tree_add_7_27_groupi_n_1666;
  wire csa_tree_add_7_27_groupi_n_1668, csa_tree_add_7_27_groupi_n_1669, csa_tree_add_7_27_groupi_n_1670, csa_tree_add_7_27_groupi_n_1671, csa_tree_add_7_27_groupi_n_1672, csa_tree_add_7_27_groupi_n_1673, csa_tree_add_7_27_groupi_n_1674, csa_tree_add_7_27_groupi_n_1675;
  wire csa_tree_add_7_27_groupi_n_1676, csa_tree_add_7_27_groupi_n_1677, csa_tree_add_7_27_groupi_n_1678, csa_tree_add_7_27_groupi_n_1679, csa_tree_add_7_27_groupi_n_1680, csa_tree_add_7_27_groupi_n_1681, csa_tree_add_7_27_groupi_n_1682, csa_tree_add_7_27_groupi_n_1683;
  wire csa_tree_add_7_27_groupi_n_1684, csa_tree_add_7_27_groupi_n_1685, csa_tree_add_7_27_groupi_n_1686, csa_tree_add_7_27_groupi_n_1687, csa_tree_add_7_27_groupi_n_1688, csa_tree_add_7_27_groupi_n_1689, csa_tree_add_7_27_groupi_n_1690, csa_tree_add_7_27_groupi_n_1691;
  wire csa_tree_add_7_27_groupi_n_1692, csa_tree_add_7_27_groupi_n_1693, csa_tree_add_7_27_groupi_n_1694, csa_tree_add_7_27_groupi_n_1695, csa_tree_add_7_27_groupi_n_1696, csa_tree_add_7_27_groupi_n_1697, csa_tree_add_7_27_groupi_n_1698, csa_tree_add_7_27_groupi_n_1699;
  wire csa_tree_add_7_27_groupi_n_1700, csa_tree_add_7_27_groupi_n_1701, csa_tree_add_7_27_groupi_n_1702, csa_tree_add_7_27_groupi_n_1703, csa_tree_add_7_27_groupi_n_1704, csa_tree_add_7_27_groupi_n_1705, csa_tree_add_7_27_groupi_n_1706, csa_tree_add_7_27_groupi_n_1707;
  wire csa_tree_add_7_27_groupi_n_1708, csa_tree_add_7_27_groupi_n_1709, csa_tree_add_7_27_groupi_n_1710, csa_tree_add_7_27_groupi_n_1711, csa_tree_add_7_27_groupi_n_1712, csa_tree_add_7_27_groupi_n_1713, csa_tree_add_7_27_groupi_n_1714, csa_tree_add_7_27_groupi_n_1715;
  wire csa_tree_add_7_27_groupi_n_1716, csa_tree_add_7_27_groupi_n_1717, csa_tree_add_7_27_groupi_n_1718, csa_tree_add_7_27_groupi_n_1719, csa_tree_add_7_27_groupi_n_1720, csa_tree_add_7_27_groupi_n_1721, csa_tree_add_7_27_groupi_n_1723, csa_tree_add_7_27_groupi_n_1724;
  wire csa_tree_add_7_27_groupi_n_1725, csa_tree_add_7_27_groupi_n_1726, csa_tree_add_7_27_groupi_n_1727, csa_tree_add_7_27_groupi_n_1728, csa_tree_add_7_27_groupi_n_1729, csa_tree_add_7_27_groupi_n_1730, csa_tree_add_7_27_groupi_n_1731, csa_tree_add_7_27_groupi_n_1732;
  wire csa_tree_add_7_27_groupi_n_1733, csa_tree_add_7_27_groupi_n_1734, csa_tree_add_7_27_groupi_n_1735, csa_tree_add_7_27_groupi_n_1736, csa_tree_add_7_27_groupi_n_1737, csa_tree_add_7_27_groupi_n_1738, csa_tree_add_7_27_groupi_n_1739, csa_tree_add_7_27_groupi_n_1740;
  wire csa_tree_add_7_27_groupi_n_1741, csa_tree_add_7_27_groupi_n_1742, csa_tree_add_7_27_groupi_n_1743, csa_tree_add_7_27_groupi_n_1744, csa_tree_add_7_27_groupi_n_1745, csa_tree_add_7_27_groupi_n_1746, csa_tree_add_7_27_groupi_n_1747, csa_tree_add_7_27_groupi_n_1748;
  wire csa_tree_add_7_27_groupi_n_1749, csa_tree_add_7_27_groupi_n_1750, csa_tree_add_7_27_groupi_n_1751, csa_tree_add_7_27_groupi_n_1752, csa_tree_add_7_27_groupi_n_1753, csa_tree_add_7_27_groupi_n_1754, csa_tree_add_7_27_groupi_n_1755, csa_tree_add_7_27_groupi_n_1756;
  wire csa_tree_add_7_27_groupi_n_1757, csa_tree_add_7_27_groupi_n_1758, csa_tree_add_7_27_groupi_n_1759, csa_tree_add_7_27_groupi_n_1760, csa_tree_add_7_27_groupi_n_1761, csa_tree_add_7_27_groupi_n_1762, csa_tree_add_7_27_groupi_n_1763, csa_tree_add_7_27_groupi_n_1764;
  wire csa_tree_add_7_27_groupi_n_1765, csa_tree_add_7_27_groupi_n_1766, csa_tree_add_7_27_groupi_n_1767, csa_tree_add_7_27_groupi_n_1768, csa_tree_add_7_27_groupi_n_1769, csa_tree_add_7_27_groupi_n_1770, csa_tree_add_7_27_groupi_n_1771, csa_tree_add_7_27_groupi_n_1772;
  wire csa_tree_add_7_27_groupi_n_1773, csa_tree_add_7_27_groupi_n_1774, csa_tree_add_7_27_groupi_n_1775, csa_tree_add_7_27_groupi_n_1776, csa_tree_add_7_27_groupi_n_1777, csa_tree_add_7_27_groupi_n_1778, csa_tree_add_7_27_groupi_n_1779, csa_tree_add_7_27_groupi_n_1780;
  wire csa_tree_add_7_27_groupi_n_1781, csa_tree_add_7_27_groupi_n_1782, csa_tree_add_7_27_groupi_n_1783, csa_tree_add_7_27_groupi_n_1784, csa_tree_add_7_27_groupi_n_1785, csa_tree_add_7_27_groupi_n_1786, csa_tree_add_7_27_groupi_n_1787, csa_tree_add_7_27_groupi_n_1788;
  wire csa_tree_add_7_27_groupi_n_1789, csa_tree_add_7_27_groupi_n_1790, csa_tree_add_7_27_groupi_n_1791, csa_tree_add_7_27_groupi_n_1792, csa_tree_add_7_27_groupi_n_1793, csa_tree_add_7_27_groupi_n_1794, csa_tree_add_7_27_groupi_n_1795, csa_tree_add_7_27_groupi_n_1796;
  wire csa_tree_add_7_27_groupi_n_1797, csa_tree_add_7_27_groupi_n_1798, csa_tree_add_7_27_groupi_n_1799, csa_tree_add_7_27_groupi_n_1800, csa_tree_add_7_27_groupi_n_1801, csa_tree_add_7_27_groupi_n_1802, csa_tree_add_7_27_groupi_n_1803, csa_tree_add_7_27_groupi_n_1804;
  wire csa_tree_add_7_27_groupi_n_1805, csa_tree_add_7_27_groupi_n_1806, csa_tree_add_7_27_groupi_n_1807, csa_tree_add_7_27_groupi_n_1808, csa_tree_add_7_27_groupi_n_1809, csa_tree_add_7_27_groupi_n_1810, csa_tree_add_7_27_groupi_n_1811, csa_tree_add_7_27_groupi_n_1812;
  wire csa_tree_add_7_27_groupi_n_1813, csa_tree_add_7_27_groupi_n_1814, csa_tree_add_7_27_groupi_n_1815, csa_tree_add_7_27_groupi_n_1816, csa_tree_add_7_27_groupi_n_1817, csa_tree_add_7_27_groupi_n_1818, csa_tree_add_7_27_groupi_n_1819, csa_tree_add_7_27_groupi_n_1820;
  wire csa_tree_add_7_27_groupi_n_1821, csa_tree_add_7_27_groupi_n_1822, csa_tree_add_7_27_groupi_n_1823, csa_tree_add_7_27_groupi_n_1824, csa_tree_add_7_27_groupi_n_1825, csa_tree_add_7_27_groupi_n_1826, csa_tree_add_7_27_groupi_n_1827, csa_tree_add_7_27_groupi_n_1828;
  wire csa_tree_add_7_27_groupi_n_1829, csa_tree_add_7_27_groupi_n_1831, csa_tree_add_7_27_groupi_n_1832, csa_tree_add_7_27_groupi_n_1833, csa_tree_add_7_27_groupi_n_1834, csa_tree_add_7_27_groupi_n_1835, csa_tree_add_7_27_groupi_n_1836, csa_tree_add_7_27_groupi_n_1837;
  wire csa_tree_add_7_27_groupi_n_1838, csa_tree_add_7_27_groupi_n_1839, csa_tree_add_7_27_groupi_n_1840, csa_tree_add_7_27_groupi_n_1841, csa_tree_add_7_27_groupi_n_1842, csa_tree_add_7_27_groupi_n_1843, csa_tree_add_7_27_groupi_n_1844, csa_tree_add_7_27_groupi_n_1845;
  wire csa_tree_add_7_27_groupi_n_1846, csa_tree_add_7_27_groupi_n_1847, csa_tree_add_7_27_groupi_n_1848, csa_tree_add_7_27_groupi_n_1849, csa_tree_add_7_27_groupi_n_1850, csa_tree_add_7_27_groupi_n_1851, csa_tree_add_7_27_groupi_n_1852, csa_tree_add_7_27_groupi_n_1853;
  wire csa_tree_add_7_27_groupi_n_1854, csa_tree_add_7_27_groupi_n_1855, csa_tree_add_7_27_groupi_n_1856, csa_tree_add_7_27_groupi_n_1857, csa_tree_add_7_27_groupi_n_1858, csa_tree_add_7_27_groupi_n_1859, csa_tree_add_7_27_groupi_n_1860, csa_tree_add_7_27_groupi_n_1861;
  wire csa_tree_add_7_27_groupi_n_1862, csa_tree_add_7_27_groupi_n_1863, csa_tree_add_7_27_groupi_n_1864, csa_tree_add_7_27_groupi_n_1865, csa_tree_add_7_27_groupi_n_1866, csa_tree_add_7_27_groupi_n_1867, csa_tree_add_7_27_groupi_n_1868, csa_tree_add_7_27_groupi_n_1869;
  wire csa_tree_add_7_27_groupi_n_1870, csa_tree_add_7_27_groupi_n_1871, csa_tree_add_7_27_groupi_n_1872, csa_tree_add_7_27_groupi_n_1873, csa_tree_add_7_27_groupi_n_1875, csa_tree_add_7_27_groupi_n_1876, csa_tree_add_7_27_groupi_n_1877, csa_tree_add_7_27_groupi_n_1878;
  wire csa_tree_add_7_27_groupi_n_1879, csa_tree_add_7_27_groupi_n_1880, csa_tree_add_7_27_groupi_n_1881, csa_tree_add_7_27_groupi_n_1882, csa_tree_add_7_27_groupi_n_1883, csa_tree_add_7_27_groupi_n_1884, csa_tree_add_7_27_groupi_n_1885, csa_tree_add_7_27_groupi_n_1886;
  wire csa_tree_add_7_27_groupi_n_1887, csa_tree_add_7_27_groupi_n_1888, csa_tree_add_7_27_groupi_n_1889, csa_tree_add_7_27_groupi_n_1890, csa_tree_add_7_27_groupi_n_1891, csa_tree_add_7_27_groupi_n_1892, csa_tree_add_7_27_groupi_n_1893, csa_tree_add_7_27_groupi_n_1894;
  wire csa_tree_add_7_27_groupi_n_1895, csa_tree_add_7_27_groupi_n_1896, csa_tree_add_7_27_groupi_n_1897, csa_tree_add_7_27_groupi_n_1898, csa_tree_add_7_27_groupi_n_1899, csa_tree_add_7_27_groupi_n_1900, csa_tree_add_7_27_groupi_n_1901, csa_tree_add_7_27_groupi_n_1902;
  wire csa_tree_add_7_27_groupi_n_1903, csa_tree_add_7_27_groupi_n_1904, csa_tree_add_7_27_groupi_n_1905, csa_tree_add_7_27_groupi_n_1906, csa_tree_add_7_27_groupi_n_1907, csa_tree_add_7_27_groupi_n_1908, csa_tree_add_7_27_groupi_n_1909, csa_tree_add_7_27_groupi_n_1910;
  wire csa_tree_add_7_27_groupi_n_1911, csa_tree_add_7_27_groupi_n_1912, csa_tree_add_7_27_groupi_n_1913, csa_tree_add_7_27_groupi_n_1914, csa_tree_add_7_27_groupi_n_1915, csa_tree_add_7_27_groupi_n_1916, csa_tree_add_7_27_groupi_n_1917, csa_tree_add_7_27_groupi_n_1918;
  wire csa_tree_add_7_27_groupi_n_1919, csa_tree_add_7_27_groupi_n_1920, csa_tree_add_7_27_groupi_n_1922, csa_tree_add_7_27_groupi_n_1923, csa_tree_add_7_27_groupi_n_1924, csa_tree_add_7_27_groupi_n_1925, csa_tree_add_7_27_groupi_n_1926, csa_tree_add_7_27_groupi_n_1927;
  wire csa_tree_add_7_27_groupi_n_1928, csa_tree_add_7_27_groupi_n_1929, csa_tree_add_7_27_groupi_n_1930, csa_tree_add_7_27_groupi_n_1931, csa_tree_add_7_27_groupi_n_1932, csa_tree_add_7_27_groupi_n_1933, csa_tree_add_7_27_groupi_n_1934, csa_tree_add_7_27_groupi_n_1935;
  wire csa_tree_add_7_27_groupi_n_1936, csa_tree_add_7_27_groupi_n_1937, csa_tree_add_7_27_groupi_n_1938, csa_tree_add_7_27_groupi_n_1939, csa_tree_add_7_27_groupi_n_1940, csa_tree_add_7_27_groupi_n_1941, csa_tree_add_7_27_groupi_n_1942, csa_tree_add_7_27_groupi_n_1943;
  wire csa_tree_add_7_27_groupi_n_1944, csa_tree_add_7_27_groupi_n_1945, csa_tree_add_7_27_groupi_n_1946, csa_tree_add_7_27_groupi_n_1947, csa_tree_add_7_27_groupi_n_1948, csa_tree_add_7_27_groupi_n_1949, csa_tree_add_7_27_groupi_n_1950, csa_tree_add_7_27_groupi_n_1951;
  wire csa_tree_add_7_27_groupi_n_1952, csa_tree_add_7_27_groupi_n_1953, csa_tree_add_7_27_groupi_n_1954, csa_tree_add_7_27_groupi_n_1955, csa_tree_add_7_27_groupi_n_1956, csa_tree_add_7_27_groupi_n_1957, csa_tree_add_7_27_groupi_n_1958, csa_tree_add_7_27_groupi_n_1959;
  wire csa_tree_add_7_27_groupi_n_1960, csa_tree_add_7_27_groupi_n_1961, csa_tree_add_7_27_groupi_n_1962, csa_tree_add_7_27_groupi_n_1963, csa_tree_add_7_27_groupi_n_1964, csa_tree_add_7_27_groupi_n_1965, csa_tree_add_7_27_groupi_n_1966, csa_tree_add_7_27_groupi_n_1967;
  wire csa_tree_add_7_27_groupi_n_1968, csa_tree_add_7_27_groupi_n_1969, csa_tree_add_7_27_groupi_n_1970, csa_tree_add_7_27_groupi_n_1971, csa_tree_add_7_27_groupi_n_1972, csa_tree_add_7_27_groupi_n_1973, csa_tree_add_7_27_groupi_n_1974, csa_tree_add_7_27_groupi_n_1975;
  wire csa_tree_add_7_27_groupi_n_1976, csa_tree_add_7_27_groupi_n_1977, csa_tree_add_7_27_groupi_n_1978, csa_tree_add_7_27_groupi_n_1979, csa_tree_add_7_27_groupi_n_1980, csa_tree_add_7_27_groupi_n_1981, csa_tree_add_7_27_groupi_n_1982, csa_tree_add_7_27_groupi_n_1983;
  wire csa_tree_add_7_27_groupi_n_1984, csa_tree_add_7_27_groupi_n_1985, csa_tree_add_7_27_groupi_n_1986, csa_tree_add_7_27_groupi_n_1987, csa_tree_add_7_27_groupi_n_1988, csa_tree_add_7_27_groupi_n_1989, csa_tree_add_7_27_groupi_n_1990, csa_tree_add_7_27_groupi_n_1991;
  wire csa_tree_add_7_27_groupi_n_1992, csa_tree_add_7_27_groupi_n_1993, csa_tree_add_7_27_groupi_n_1994, csa_tree_add_7_27_groupi_n_1995, csa_tree_add_7_27_groupi_n_1996, csa_tree_add_7_27_groupi_n_1997, csa_tree_add_7_27_groupi_n_1998, csa_tree_add_7_27_groupi_n_1999;
  wire csa_tree_add_7_27_groupi_n_2000, csa_tree_add_7_27_groupi_n_2001, csa_tree_add_7_27_groupi_n_2002, csa_tree_add_7_27_groupi_n_2003, csa_tree_add_7_27_groupi_n_2004, csa_tree_add_7_27_groupi_n_2005, csa_tree_add_7_27_groupi_n_2006, csa_tree_add_7_27_groupi_n_2007;
  wire csa_tree_add_7_27_groupi_n_2008, csa_tree_add_7_27_groupi_n_2009, csa_tree_add_7_27_groupi_n_2010, csa_tree_add_7_27_groupi_n_2011, csa_tree_add_7_27_groupi_n_2012, csa_tree_add_7_27_groupi_n_2013, csa_tree_add_7_27_groupi_n_2014, csa_tree_add_7_27_groupi_n_2015;
  wire csa_tree_add_7_27_groupi_n_2016, csa_tree_add_7_27_groupi_n_2018, csa_tree_add_7_27_groupi_n_2019, csa_tree_add_7_27_groupi_n_2020, csa_tree_add_7_27_groupi_n_2021, csa_tree_add_7_27_groupi_n_2022, csa_tree_add_7_27_groupi_n_2023, csa_tree_add_7_27_groupi_n_2024;
  wire csa_tree_add_7_27_groupi_n_2025, csa_tree_add_7_27_groupi_n_2026, csa_tree_add_7_27_groupi_n_2027, csa_tree_add_7_27_groupi_n_2028, csa_tree_add_7_27_groupi_n_2029, csa_tree_add_7_27_groupi_n_2030, csa_tree_add_7_27_groupi_n_2031, csa_tree_add_7_27_groupi_n_2032;
  wire csa_tree_add_7_27_groupi_n_2033, csa_tree_add_7_27_groupi_n_2034, csa_tree_add_7_27_groupi_n_2035, csa_tree_add_7_27_groupi_n_2036, csa_tree_add_7_27_groupi_n_2037, csa_tree_add_7_27_groupi_n_2038, csa_tree_add_7_27_groupi_n_2039, csa_tree_add_7_27_groupi_n_2040;
  wire csa_tree_add_7_27_groupi_n_2041, csa_tree_add_7_27_groupi_n_2042, csa_tree_add_7_27_groupi_n_2043, csa_tree_add_7_27_groupi_n_2044, csa_tree_add_7_27_groupi_n_2045, csa_tree_add_7_27_groupi_n_2046, csa_tree_add_7_27_groupi_n_2047, csa_tree_add_7_27_groupi_n_2048;
  wire csa_tree_add_7_27_groupi_n_2049, csa_tree_add_7_27_groupi_n_2050, csa_tree_add_7_27_groupi_n_2051, csa_tree_add_7_27_groupi_n_2052, csa_tree_add_7_27_groupi_n_2053, csa_tree_add_7_27_groupi_n_2054, csa_tree_add_7_27_groupi_n_2055, csa_tree_add_7_27_groupi_n_2056;
  wire csa_tree_add_7_27_groupi_n_2057, csa_tree_add_7_27_groupi_n_2058, csa_tree_add_7_27_groupi_n_2059, csa_tree_add_7_27_groupi_n_2060, csa_tree_add_7_27_groupi_n_2061, csa_tree_add_7_27_groupi_n_2062, csa_tree_add_7_27_groupi_n_2063, csa_tree_add_7_27_groupi_n_2064;
  wire csa_tree_add_7_27_groupi_n_2065, csa_tree_add_7_27_groupi_n_2066, csa_tree_add_7_27_groupi_n_2067, csa_tree_add_7_27_groupi_n_2068, csa_tree_add_7_27_groupi_n_2069, csa_tree_add_7_27_groupi_n_2070, csa_tree_add_7_27_groupi_n_2071, csa_tree_add_7_27_groupi_n_2072;
  wire csa_tree_add_7_27_groupi_n_2074, csa_tree_add_7_27_groupi_n_2075, csa_tree_add_7_27_groupi_n_2076, csa_tree_add_7_27_groupi_n_2077, csa_tree_add_7_27_groupi_n_2078, csa_tree_add_7_27_groupi_n_2079, csa_tree_add_7_27_groupi_n_2080, csa_tree_add_7_27_groupi_n_2081;
  wire csa_tree_add_7_27_groupi_n_2082, csa_tree_add_7_27_groupi_n_2083, csa_tree_add_7_27_groupi_n_2084, csa_tree_add_7_27_groupi_n_2085, csa_tree_add_7_27_groupi_n_2086, csa_tree_add_7_27_groupi_n_2087, csa_tree_add_7_27_groupi_n_2088, csa_tree_add_7_27_groupi_n_2089;
  wire csa_tree_add_7_27_groupi_n_2090, csa_tree_add_7_27_groupi_n_2091, csa_tree_add_7_27_groupi_n_2092, csa_tree_add_7_27_groupi_n_2093, csa_tree_add_7_27_groupi_n_2094, csa_tree_add_7_27_groupi_n_2095, csa_tree_add_7_27_groupi_n_2096, csa_tree_add_7_27_groupi_n_2097;
  wire csa_tree_add_7_27_groupi_n_2098, csa_tree_add_7_27_groupi_n_2099, csa_tree_add_7_27_groupi_n_2100, csa_tree_add_7_27_groupi_n_2101, csa_tree_add_7_27_groupi_n_2102, csa_tree_add_7_27_groupi_n_2103, csa_tree_add_7_27_groupi_n_2104, csa_tree_add_7_27_groupi_n_2105;
  wire csa_tree_add_7_27_groupi_n_2106, csa_tree_add_7_27_groupi_n_2107, csa_tree_add_7_27_groupi_n_2108, csa_tree_add_7_27_groupi_n_2109, csa_tree_add_7_27_groupi_n_2110, csa_tree_add_7_27_groupi_n_2111, csa_tree_add_7_27_groupi_n_2112, csa_tree_add_7_27_groupi_n_2113;
  wire csa_tree_add_7_27_groupi_n_2114, csa_tree_add_7_27_groupi_n_2115, csa_tree_add_7_27_groupi_n_2116, csa_tree_add_7_27_groupi_n_2117, csa_tree_add_7_27_groupi_n_2118, csa_tree_add_7_27_groupi_n_2119, csa_tree_add_7_27_groupi_n_2120, csa_tree_add_7_27_groupi_n_2121;
  wire csa_tree_add_7_27_groupi_n_2122, csa_tree_add_7_27_groupi_n_2123, csa_tree_add_7_27_groupi_n_2124, csa_tree_add_7_27_groupi_n_2125, csa_tree_add_7_27_groupi_n_2126, csa_tree_add_7_27_groupi_n_2127, csa_tree_add_7_27_groupi_n_2128, csa_tree_add_7_27_groupi_n_2129;
  wire csa_tree_add_7_27_groupi_n_2130, csa_tree_add_7_27_groupi_n_2131, csa_tree_add_7_27_groupi_n_2132, csa_tree_add_7_27_groupi_n_2133, csa_tree_add_7_27_groupi_n_2134, csa_tree_add_7_27_groupi_n_2135, csa_tree_add_7_27_groupi_n_2136, csa_tree_add_7_27_groupi_n_2137;
  wire csa_tree_add_7_27_groupi_n_2138, csa_tree_add_7_27_groupi_n_2139, csa_tree_add_7_27_groupi_n_2140, csa_tree_add_7_27_groupi_n_2141, csa_tree_add_7_27_groupi_n_2142, csa_tree_add_7_27_groupi_n_2143, csa_tree_add_7_27_groupi_n_2144, csa_tree_add_7_27_groupi_n_2145;
  wire csa_tree_add_7_27_groupi_n_2146, csa_tree_add_7_27_groupi_n_2147, csa_tree_add_7_27_groupi_n_2148, csa_tree_add_7_27_groupi_n_2149, csa_tree_add_7_27_groupi_n_2150, csa_tree_add_7_27_groupi_n_2151, csa_tree_add_7_27_groupi_n_2152, csa_tree_add_7_27_groupi_n_2154;
  wire csa_tree_add_7_27_groupi_n_2155, csa_tree_add_7_27_groupi_n_2156, csa_tree_add_7_27_groupi_n_2157, csa_tree_add_7_27_groupi_n_2158, csa_tree_add_7_27_groupi_n_2159, csa_tree_add_7_27_groupi_n_2160, csa_tree_add_7_27_groupi_n_2161, csa_tree_add_7_27_groupi_n_2162;
  wire csa_tree_add_7_27_groupi_n_2163, csa_tree_add_7_27_groupi_n_2164, csa_tree_add_7_27_groupi_n_2165, csa_tree_add_7_27_groupi_n_2166, csa_tree_add_7_27_groupi_n_2167, csa_tree_add_7_27_groupi_n_2168, csa_tree_add_7_27_groupi_n_2169, csa_tree_add_7_27_groupi_n_2170;
  wire csa_tree_add_7_27_groupi_n_2171, csa_tree_add_7_27_groupi_n_2172, csa_tree_add_7_27_groupi_n_2173, csa_tree_add_7_27_groupi_n_2174, csa_tree_add_7_27_groupi_n_2175, csa_tree_add_7_27_groupi_n_2176, csa_tree_add_7_27_groupi_n_2177, csa_tree_add_7_27_groupi_n_2178;
  wire csa_tree_add_7_27_groupi_n_2179, csa_tree_add_7_27_groupi_n_2180, csa_tree_add_7_27_groupi_n_2181, csa_tree_add_7_27_groupi_n_2182, csa_tree_add_7_27_groupi_n_2183, csa_tree_add_7_27_groupi_n_2184, csa_tree_add_7_27_groupi_n_2185, csa_tree_add_7_27_groupi_n_2186;
  wire csa_tree_add_7_27_groupi_n_2187, csa_tree_add_7_27_groupi_n_2188, csa_tree_add_7_27_groupi_n_2189, csa_tree_add_7_27_groupi_n_2190, csa_tree_add_7_27_groupi_n_2191, csa_tree_add_7_27_groupi_n_2192, csa_tree_add_7_27_groupi_n_2193, csa_tree_add_7_27_groupi_n_2194;
  wire csa_tree_add_7_27_groupi_n_2195, csa_tree_add_7_27_groupi_n_2196, csa_tree_add_7_27_groupi_n_2197, csa_tree_add_7_27_groupi_n_2198, csa_tree_add_7_27_groupi_n_2199, csa_tree_add_7_27_groupi_n_2200, csa_tree_add_7_27_groupi_n_2201, csa_tree_add_7_27_groupi_n_2202;
  wire csa_tree_add_7_27_groupi_n_2203, csa_tree_add_7_27_groupi_n_2204, csa_tree_add_7_27_groupi_n_2206, csa_tree_add_7_27_groupi_n_2207, csa_tree_add_7_27_groupi_n_2208, csa_tree_add_7_27_groupi_n_2209, csa_tree_add_7_27_groupi_n_2210, csa_tree_add_7_27_groupi_n_2211;
  wire csa_tree_add_7_27_groupi_n_2212, csa_tree_add_7_27_groupi_n_2213, csa_tree_add_7_27_groupi_n_2214, csa_tree_add_7_27_groupi_n_2215, csa_tree_add_7_27_groupi_n_2216, csa_tree_add_7_27_groupi_n_2217, csa_tree_add_7_27_groupi_n_2218, csa_tree_add_7_27_groupi_n_2219;
  wire csa_tree_add_7_27_groupi_n_2220, csa_tree_add_7_27_groupi_n_2221, csa_tree_add_7_27_groupi_n_2222, csa_tree_add_7_27_groupi_n_2223, csa_tree_add_7_27_groupi_n_2224, csa_tree_add_7_27_groupi_n_2225, csa_tree_add_7_27_groupi_n_2226, csa_tree_add_7_27_groupi_n_2227;
  wire csa_tree_add_7_27_groupi_n_2228, csa_tree_add_7_27_groupi_n_2229, csa_tree_add_7_27_groupi_n_2230, csa_tree_add_7_27_groupi_n_2231, csa_tree_add_7_27_groupi_n_2232, csa_tree_add_7_27_groupi_n_2233, csa_tree_add_7_27_groupi_n_2234, csa_tree_add_7_27_groupi_n_2235;
  wire csa_tree_add_7_27_groupi_n_2236, csa_tree_add_7_27_groupi_n_2237, csa_tree_add_7_27_groupi_n_2238, csa_tree_add_7_27_groupi_n_2239, csa_tree_add_7_27_groupi_n_2240, csa_tree_add_7_27_groupi_n_2241, csa_tree_add_7_27_groupi_n_2242, csa_tree_add_7_27_groupi_n_2243;
  wire csa_tree_add_7_27_groupi_n_2244, csa_tree_add_7_27_groupi_n_2245, csa_tree_add_7_27_groupi_n_2246, csa_tree_add_7_27_groupi_n_2247, csa_tree_add_7_27_groupi_n_2248, csa_tree_add_7_27_groupi_n_2249, csa_tree_add_7_27_groupi_n_2250, csa_tree_add_7_27_groupi_n_2251;
  wire csa_tree_add_7_27_groupi_n_2252, csa_tree_add_7_27_groupi_n_2253, csa_tree_add_7_27_groupi_n_2255, csa_tree_add_7_27_groupi_n_2256, csa_tree_add_7_27_groupi_n_2257, csa_tree_add_7_27_groupi_n_2258, csa_tree_add_7_27_groupi_n_2259, csa_tree_add_7_27_groupi_n_2260;
  wire csa_tree_add_7_27_groupi_n_2261, csa_tree_add_7_27_groupi_n_2262, csa_tree_add_7_27_groupi_n_2263, csa_tree_add_7_27_groupi_n_2264, csa_tree_add_7_27_groupi_n_2265, csa_tree_add_7_27_groupi_n_2266, csa_tree_add_7_27_groupi_n_2267, csa_tree_add_7_27_groupi_n_2268;
  wire csa_tree_add_7_27_groupi_n_2269, csa_tree_add_7_27_groupi_n_2270, csa_tree_add_7_27_groupi_n_2271, csa_tree_add_7_27_groupi_n_2272, csa_tree_add_7_27_groupi_n_2273, csa_tree_add_7_27_groupi_n_2274, csa_tree_add_7_27_groupi_n_2275, csa_tree_add_7_27_groupi_n_2276;
  wire csa_tree_add_7_27_groupi_n_2277, csa_tree_add_7_27_groupi_n_2278, csa_tree_add_7_27_groupi_n_2279, csa_tree_add_7_27_groupi_n_2280, csa_tree_add_7_27_groupi_n_2281, csa_tree_add_7_27_groupi_n_2282, csa_tree_add_7_27_groupi_n_2283, csa_tree_add_7_27_groupi_n_2284;
  wire csa_tree_add_7_27_groupi_n_2285, csa_tree_add_7_27_groupi_n_2286, csa_tree_add_7_27_groupi_n_2287, csa_tree_add_7_27_groupi_n_2288, csa_tree_add_7_27_groupi_n_2289, csa_tree_add_7_27_groupi_n_2290, csa_tree_add_7_27_groupi_n_2291, csa_tree_add_7_27_groupi_n_2292;
  wire csa_tree_add_7_27_groupi_n_2293, csa_tree_add_7_27_groupi_n_2294, csa_tree_add_7_27_groupi_n_2295, csa_tree_add_7_27_groupi_n_2296, csa_tree_add_7_27_groupi_n_2297, csa_tree_add_7_27_groupi_n_2298, csa_tree_add_7_27_groupi_n_2299, csa_tree_add_7_27_groupi_n_2300;
  wire csa_tree_add_7_27_groupi_n_2301, csa_tree_add_7_27_groupi_n_2302, csa_tree_add_7_27_groupi_n_2303, csa_tree_add_7_27_groupi_n_2304, csa_tree_add_7_27_groupi_n_2305, csa_tree_add_7_27_groupi_n_2306, csa_tree_add_7_27_groupi_n_2307, csa_tree_add_7_27_groupi_n_2308;
  wire csa_tree_add_7_27_groupi_n_2309, csa_tree_add_7_27_groupi_n_2311, csa_tree_add_7_27_groupi_n_2312, csa_tree_add_7_27_groupi_n_2314, csa_tree_add_7_27_groupi_n_2315, csa_tree_add_7_27_groupi_n_2317, csa_tree_add_7_27_groupi_n_2318, csa_tree_add_7_27_groupi_n_2320;
  wire csa_tree_add_7_27_groupi_n_2321, csa_tree_add_7_27_groupi_n_2323, csa_tree_add_7_27_groupi_n_2324, csa_tree_add_7_27_groupi_n_2325, csa_tree_add_7_27_groupi_n_2327, csa_tree_add_7_27_groupi_n_2328, csa_tree_add_7_27_groupi_n_2329, csa_tree_add_7_27_groupi_n_2330;
  wire csa_tree_add_7_27_groupi_n_2331, csa_tree_add_7_27_groupi_n_2332, csa_tree_add_7_27_groupi_n_2333, csa_tree_add_7_27_groupi_n_2334, csa_tree_add_7_27_groupi_n_2335, csa_tree_add_7_27_groupi_n_2337, csa_tree_add_7_27_groupi_n_2338, csa_tree_add_7_27_groupi_n_2340;
  wire csa_tree_add_7_27_groupi_n_2341, csa_tree_add_7_27_groupi_n_2342, csa_tree_add_7_27_groupi_n_2343, csa_tree_add_7_27_groupi_n_2344, csa_tree_add_7_27_groupi_n_2345, csa_tree_add_7_27_groupi_n_2347, csa_tree_add_7_27_groupi_n_2348, csa_tree_add_7_27_groupi_n_2350;
  wire csa_tree_add_7_27_groupi_n_2351, csa_tree_add_7_27_groupi_n_2353, dec_sub_8_33_n_3, dec_sub_8_33_n_6, dec_sub_8_33_n_7, dec_sub_8_33_n_8, dec_sub_8_33_n_9, dec_sub_8_33_n_10;
  wire dec_sub_8_33_n_11, dec_sub_8_33_n_12, dec_sub_8_33_n_13, dec_sub_8_33_n_14, dec_sub_8_33_n_15, dec_sub_8_33_n_16, dec_sub_8_33_n_17, dec_sub_8_33_n_18;
  wire dec_sub_8_33_n_19, dec_sub_8_33_n_20, dec_sub_8_33_n_21, dec_sub_8_33_n_22, dec_sub_8_33_n_23, dec_sub_8_33_n_24, dec_sub_8_33_n_25, dec_sub_8_33_n_26;
  wire dec_sub_8_33_n_27, dec_sub_8_33_n_28, dec_sub_8_33_n_29, dec_sub_8_33_n_30, dec_sub_8_33_n_31, dec_sub_8_33_n_32, dec_sub_8_33_n_33, dec_sub_8_33_n_34;
  wire dec_sub_8_33_n_35, dec_sub_8_33_n_36, dec_sub_8_33_n_37, dec_sub_8_33_n_38, dec_sub_8_33_n_39, dec_sub_8_33_n_40, dec_sub_8_33_n_41, dec_sub_8_33_n_42;
  wire dec_sub_8_33_n_43, dec_sub_8_33_n_44, dec_sub_8_33_n_45, dec_sub_8_33_n_46, dec_sub_8_33_n_47, dec_sub_8_33_n_48, dec_sub_8_33_n_49, dec_sub_8_33_n_50;
  wire dec_sub_8_33_n_51, dec_sub_8_33_n_52, dec_sub_8_33_n_53, dec_sub_8_33_n_54, dec_sub_8_33_n_55, dec_sub_8_33_n_56, dec_sub_8_33_n_57, dec_sub_8_33_n_58;
  wire dec_sub_8_33_n_59, dec_sub_8_33_n_60, dec_sub_8_33_n_61, dec_sub_8_33_n_62, dec_sub_8_33_n_63, dec_sub_8_33_n_64, dec_sub_8_33_n_65, dec_sub_8_33_n_66;
  wire dec_sub_8_33_n_67, dec_sub_8_33_n_68, dec_sub_8_33_n_69, dec_sub_8_33_n_70, dec_sub_8_33_n_71, dec_sub_8_33_n_72, dec_sub_8_33_n_73, dec_sub_8_33_n_74;
  wire dec_sub_8_33_n_75, dec_sub_8_33_n_76, dec_sub_8_33_n_77, dec_sub_8_33_n_79, dec_sub_8_33_n_80, dec_sub_8_33_n_81, dec_sub_8_33_n_82, dec_sub_8_33_n_84;
  wire dec_sub_8_33_n_85, dec_sub_8_33_n_86, dec_sub_8_33_n_87, dec_sub_8_33_n_88, dec_sub_8_33_n_90, dec_sub_8_33_n_91, dec_sub_8_33_n_92, dec_sub_8_33_n_93;
  wire dec_sub_8_33_n_96, dec_sub_8_33_n_97, dec_sub_8_33_n_99, dec_sub_8_33_n_100, dec_sub_8_33_n_101, dec_sub_8_33_n_102, dec_sub_8_33_n_104, dec_sub_8_33_n_105;
  wire dec_sub_8_33_n_106, dec_sub_8_33_n_110, dec_sub_8_33_n_113, dec_sub_8_33_n_114, dec_sub_8_33_n_115, dec_sub_8_33_n_117, dec_sub_8_33_n_118, dec_sub_8_33_n_119;
  wire dec_sub_8_33_n_120, dec_sub_8_33_n_122, dec_sub_8_33_n_123, dec_sub_8_33_n_124, dec_sub_8_33_n_128, dec_sub_8_33_n_131, dec_sub_8_33_n_132, dec_sub_8_33_n_133;
  wire dec_sub_8_33_n_135, dec_sub_8_33_n_136, dec_sub_8_33_n_137, dec_sub_8_33_n_138, dec_sub_8_33_n_140, dec_sub_8_33_n_141, dec_sub_8_33_n_143, dec_sub_8_33_n_144;
  wire dec_sub_8_33_n_146, dec_sub_8_33_n_147, dec_sub_8_33_n_148, dec_sub_8_33_n_150, inc_add_7_33_n_15, inc_add_7_33_n_16, inc_add_7_33_n_17, inc_add_7_33_n_18;
  wire inc_add_7_33_n_19, inc_add_7_33_n_20, inc_add_7_33_n_21, inc_add_7_33_n_22, inc_add_7_33_n_23, inc_add_7_33_n_24, inc_add_7_33_n_25, inc_add_7_33_n_26;
  wire inc_add_7_33_n_27, inc_add_7_33_n_28, inc_add_7_33_n_29, inc_add_7_33_n_30, inc_add_7_33_n_31, inc_add_7_33_n_32, inc_add_7_33_n_33, inc_add_7_33_n_34;
  wire inc_add_7_33_n_35, inc_add_7_33_n_36, inc_add_7_33_n_37, inc_add_7_33_n_38, inc_add_7_33_n_39, inc_add_7_33_n_40, inc_add_7_33_n_41, inc_add_7_33_n_42;
  wire inc_add_7_33_n_43, inc_add_7_33_n_44, inc_add_7_33_n_45, inc_add_7_33_n_46, inc_add_7_33_n_47, inc_add_7_33_n_48, inc_add_7_33_n_49, inc_add_7_33_n_50;
  wire inc_add_7_33_n_51, inc_add_7_33_n_52, inc_add_7_33_n_53, inc_add_7_33_n_54, inc_add_7_33_n_55, inc_add_7_33_n_56, inc_add_7_33_n_57, inc_add_7_33_n_58;
  wire inc_add_7_33_n_59, inc_add_7_33_n_60, inc_add_7_33_n_61, inc_add_7_33_n_62, inc_add_7_33_n_63, inc_add_7_33_n_64, inc_add_7_33_n_65, inc_add_7_33_n_66;
  wire inc_add_7_33_n_67, inc_add_7_33_n_68, inc_add_7_33_n_69, inc_add_7_33_n_70, inc_add_7_33_n_71, inc_add_7_33_n_72, inc_add_7_33_n_73, inc_add_7_33_n_74;
  wire inc_add_7_33_n_75, inc_add_7_33_n_76, inc_add_7_33_n_77, inc_add_7_33_n_78, inc_add_7_33_n_79, inc_add_7_33_n_80, inc_add_7_33_n_81, inc_add_7_33_n_82;
  wire inc_add_7_33_n_84, inc_add_7_33_n_85, inc_add_7_33_n_86, inc_add_7_33_n_87, inc_add_7_33_n_89, inc_add_7_33_n_90, inc_add_7_33_n_91, inc_add_7_33_n_92;
  wire inc_add_7_33_n_93, inc_add_7_33_n_94, inc_add_7_33_n_95, inc_add_7_33_n_96, inc_add_7_33_n_97, inc_add_7_33_n_100, inc_add_7_33_n_101, inc_add_7_33_n_102;
  wire inc_add_7_33_n_103, inc_add_7_33_n_104, inc_add_7_33_n_105, inc_add_7_33_n_106, inc_add_7_33_n_108, inc_add_7_33_n_109, inc_add_7_33_n_110, inc_add_7_33_n_113;
  wire inc_add_7_33_n_114, inc_add_7_33_n_116, inc_add_7_33_n_117, inc_add_7_33_n_119, inc_add_7_33_n_120, inc_add_7_33_n_121, inc_add_7_33_n_122, inc_add_7_33_n_123;
  wire inc_add_7_33_n_125, inc_add_7_33_n_126, inc_add_7_33_n_127, inc_add_7_33_n_130, inc_add_7_33_n_131, inc_add_7_33_n_132, inc_add_7_33_n_133, inc_add_7_33_n_134;
  wire inc_add_7_33_n_135, inc_add_7_33_n_137, inc_add_7_33_n_138, inc_add_7_33_n_139, inc_add_7_33_n_140, inc_add_7_33_n_141, inc_add_7_33_n_144, inc_add_7_33_n_145;
  wire inc_add_7_33_n_146, inc_add_7_33_n_147, n_2, n_3, n_4, n_5, n_6, n_7;
  wire n_8, n_9, n_10, n_11, n_12, n_13, n_14, n_15;
  wire n_16, n_17, n_18, n_19, n_20, n_21, n_22, n_23;
  wire n_24, n_25, n_26, n_27, n_28, n_29, n_30, n_31;
  wire n_32, n_33;
  buf constbuf_n1(out2[0], out1[0]);
  not g17(out1[0] ,n_2);
  xnor csa_tree_add_7_27_groupi_g4832__2398(n_33 ,csa_tree_add_7_27_groupi_n_2353 ,csa_tree_add_7_27_groupi_n_1431);
  or csa_tree_add_7_27_groupi_g4833__5107(csa_tree_add_7_27_groupi_n_2353 ,csa_tree_add_7_27_groupi_n_2224 ,csa_tree_add_7_27_groupi_n_2351);
  xnor csa_tree_add_7_27_groupi_g4834__6260(n_32 ,csa_tree_add_7_27_groupi_n_2350 ,csa_tree_add_7_27_groupi_n_2253);
  and csa_tree_add_7_27_groupi_g4835__4319(csa_tree_add_7_27_groupi_n_2351 ,csa_tree_add_7_27_groupi_n_2225 ,csa_tree_add_7_27_groupi_n_2350);
  or csa_tree_add_7_27_groupi_g4836__8428(csa_tree_add_7_27_groupi_n_2350 ,csa_tree_add_7_27_groupi_n_2270 ,csa_tree_add_7_27_groupi_n_2348);
  xnor csa_tree_add_7_27_groupi_g4837__5526(n_31 ,csa_tree_add_7_27_groupi_n_2347 ,csa_tree_add_7_27_groupi_n_2278);
  and csa_tree_add_7_27_groupi_g4838__6783(csa_tree_add_7_27_groupi_n_2348 ,csa_tree_add_7_27_groupi_n_2275 ,csa_tree_add_7_27_groupi_n_2347);
  or csa_tree_add_7_27_groupi_g4839__3680(csa_tree_add_7_27_groupi_n_2347 ,csa_tree_add_7_27_groupi_n_2271 ,csa_tree_add_7_27_groupi_n_2345);
  xnor csa_tree_add_7_27_groupi_g4840__1617(n_30 ,csa_tree_add_7_27_groupi_n_2344 ,csa_tree_add_7_27_groupi_n_2280);
  nor csa_tree_add_7_27_groupi_g4841__2802(csa_tree_add_7_27_groupi_n_2345 ,csa_tree_add_7_27_groupi_n_2276 ,csa_tree_add_7_27_groupi_n_2344);
  and csa_tree_add_7_27_groupi_g4842__1705(csa_tree_add_7_27_groupi_n_2344 ,csa_tree_add_7_27_groupi_n_2343 ,csa_tree_add_7_27_groupi_n_2295);
  or csa_tree_add_7_27_groupi_g4844__5122(csa_tree_add_7_27_groupi_n_2343 ,csa_tree_add_7_27_groupi_n_2290 ,csa_tree_add_7_27_groupi_n_2342);
  and csa_tree_add_7_27_groupi_g4846__8246(csa_tree_add_7_27_groupi_n_2342 ,csa_tree_add_7_27_groupi_n_2298 ,csa_tree_add_7_27_groupi_n_2341);
  or csa_tree_add_7_27_groupi_g4848__7098(csa_tree_add_7_27_groupi_n_2341 ,csa_tree_add_7_27_groupi_n_2291 ,csa_tree_add_7_27_groupi_n_2340);
  and csa_tree_add_7_27_groupi_g4850__6131(csa_tree_add_7_27_groupi_n_2340 ,csa_tree_add_7_27_groupi_n_2266 ,csa_tree_add_7_27_groupi_n_2338);
  xnor csa_tree_add_7_27_groupi_g4851__1881(n_27 ,csa_tree_add_7_27_groupi_n_2337 ,csa_tree_add_7_27_groupi_n_2282);
  or csa_tree_add_7_27_groupi_g4852__5115(csa_tree_add_7_27_groupi_n_2338 ,csa_tree_add_7_27_groupi_n_2265 ,csa_tree_add_7_27_groupi_n_2337);
  and csa_tree_add_7_27_groupi_g4853__7482(csa_tree_add_7_27_groupi_n_2337 ,csa_tree_add_7_27_groupi_n_2335 ,csa_tree_add_7_27_groupi_n_2296);
  xnor csa_tree_add_7_27_groupi_g4854__4733(n_26 ,csa_tree_add_7_27_groupi_n_2333 ,csa_tree_add_7_27_groupi_n_2301);
  or csa_tree_add_7_27_groupi_g4855__6161(csa_tree_add_7_27_groupi_n_2335 ,csa_tree_add_7_27_groupi_n_2289 ,csa_tree_add_7_27_groupi_n_2334);
  not csa_tree_add_7_27_groupi_g4856(csa_tree_add_7_27_groupi_n_2334 ,csa_tree_add_7_27_groupi_n_2333);
  or csa_tree_add_7_27_groupi_g4857__9315(csa_tree_add_7_27_groupi_n_2333 ,csa_tree_add_7_27_groupi_n_2294 ,csa_tree_add_7_27_groupi_n_2331);
  xnor csa_tree_add_7_27_groupi_g4858__9945(csa_tree_add_7_27_groupi_n_2332 ,csa_tree_add_7_27_groupi_n_2330 ,csa_tree_add_7_27_groupi_n_2300);
  and csa_tree_add_7_27_groupi_g4859__2883(csa_tree_add_7_27_groupi_n_2331 ,csa_tree_add_7_27_groupi_n_2330 ,csa_tree_add_7_27_groupi_n_2297);
  or csa_tree_add_7_27_groupi_g4860__2346(csa_tree_add_7_27_groupi_n_2330 ,csa_tree_add_7_27_groupi_n_2328 ,csa_tree_add_7_27_groupi_n_2269);
  xnor csa_tree_add_7_27_groupi_g4861__1666(csa_tree_add_7_27_groupi_n_2329 ,csa_tree_add_7_27_groupi_n_2327 ,csa_tree_add_7_27_groupi_n_2281);
  nor csa_tree_add_7_27_groupi_g4862__7410(csa_tree_add_7_27_groupi_n_2328 ,csa_tree_add_7_27_groupi_n_2267 ,csa_tree_add_7_27_groupi_n_2327);
  and csa_tree_add_7_27_groupi_g4863__6417(csa_tree_add_7_27_groupi_n_2327 ,csa_tree_add_7_27_groupi_n_2325 ,csa_tree_add_7_27_groupi_n_2283);
  xnor csa_tree_add_7_27_groupi_g4864__5477(n_23 ,csa_tree_add_7_27_groupi_n_2323 ,csa_tree_add_7_27_groupi_n_2305);
  or csa_tree_add_7_27_groupi_g4865__2398(csa_tree_add_7_27_groupi_n_2325 ,csa_tree_add_7_27_groupi_n_2288 ,csa_tree_add_7_27_groupi_n_2324);
  not csa_tree_add_7_27_groupi_g4866(csa_tree_add_7_27_groupi_n_2324 ,csa_tree_add_7_27_groupi_n_2323);
  or csa_tree_add_7_27_groupi_g4867__5107(csa_tree_add_7_27_groupi_n_2323 ,csa_tree_add_7_27_groupi_n_2321 ,csa_tree_add_7_27_groupi_n_2293);
  xnor csa_tree_add_7_27_groupi_g4868__6260(n_22 ,csa_tree_add_7_27_groupi_n_2320 ,csa_tree_add_7_27_groupi_n_2304);
  and csa_tree_add_7_27_groupi_g4869__4319(csa_tree_add_7_27_groupi_n_2321 ,csa_tree_add_7_27_groupi_n_2292 ,csa_tree_add_7_27_groupi_n_2320);
  or csa_tree_add_7_27_groupi_g4870__8428(csa_tree_add_7_27_groupi_n_2320 ,csa_tree_add_7_27_groupi_n_2318 ,csa_tree_add_7_27_groupi_n_2268);
  xnor csa_tree_add_7_27_groupi_g4871__5526(n_21 ,csa_tree_add_7_27_groupi_n_2317 ,csa_tree_add_7_27_groupi_n_2279);
  and csa_tree_add_7_27_groupi_g4872__6783(csa_tree_add_7_27_groupi_n_2318 ,csa_tree_add_7_27_groupi_n_2317 ,csa_tree_add_7_27_groupi_n_2255);
  or csa_tree_add_7_27_groupi_g4873__3680(csa_tree_add_7_27_groupi_n_2317 ,csa_tree_add_7_27_groupi_n_2315 ,csa_tree_add_7_27_groupi_n_2284);
  xnor csa_tree_add_7_27_groupi_g4874__1617(n_20 ,csa_tree_add_7_27_groupi_n_2314 ,csa_tree_add_7_27_groupi_n_2307);
  and csa_tree_add_7_27_groupi_g4875__2802(csa_tree_add_7_27_groupi_n_2315 ,csa_tree_add_7_27_groupi_n_2285 ,csa_tree_add_7_27_groupi_n_2314);
  or csa_tree_add_7_27_groupi_g4876__1705(csa_tree_add_7_27_groupi_n_2314 ,csa_tree_add_7_27_groupi_n_2287 ,csa_tree_add_7_27_groupi_n_2312);
  xnor csa_tree_add_7_27_groupi_g4877__5122(n_19 ,csa_tree_add_7_27_groupi_n_2311 ,csa_tree_add_7_27_groupi_n_2306);
  and csa_tree_add_7_27_groupi_g4878__8246(csa_tree_add_7_27_groupi_n_2312 ,csa_tree_add_7_27_groupi_n_2286 ,csa_tree_add_7_27_groupi_n_2311);
  or csa_tree_add_7_27_groupi_g4879__7098(csa_tree_add_7_27_groupi_n_2311 ,csa_tree_add_7_27_groupi_n_2309 ,csa_tree_add_7_27_groupi_n_2272);
  xnor csa_tree_add_7_27_groupi_g4880__6131(n_18 ,csa_tree_add_7_27_groupi_n_2299 ,csa_tree_add_7_27_groupi_n_2277);
  and csa_tree_add_7_27_groupi_g4881__1881(csa_tree_add_7_27_groupi_n_2309 ,csa_tree_add_7_27_groupi_n_2274 ,csa_tree_add_7_27_groupi_n_2299);
  xnor csa_tree_add_7_27_groupi_g4882__5115(csa_tree_add_7_27_groupi_n_2308 ,csa_tree_add_7_27_groupi_n_2251 ,csa_tree_add_7_27_groupi_n_2252);
  xnor csa_tree_add_7_27_groupi_g4883__7482(csa_tree_add_7_27_groupi_n_2307 ,csa_tree_add_7_27_groupi_n_2264 ,csa_tree_add_7_27_groupi_n_2235);
  xnor csa_tree_add_7_27_groupi_g4884__4733(csa_tree_add_7_27_groupi_n_2306 ,csa_tree_add_7_27_groupi_n_2248 ,csa_tree_add_7_27_groupi_n_2262);
  xnor csa_tree_add_7_27_groupi_g4885__6161(csa_tree_add_7_27_groupi_n_2305 ,csa_tree_add_7_27_groupi_n_2258 ,csa_tree_add_7_27_groupi_n_2233);
  xnor csa_tree_add_7_27_groupi_g4886__9315(csa_tree_add_7_27_groupi_n_2304 ,csa_tree_add_7_27_groupi_n_2232 ,csa_tree_add_7_27_groupi_n_2263);
  xnor csa_tree_add_7_27_groupi_g4887__9945(csa_tree_add_7_27_groupi_n_2303 ,csa_tree_add_7_27_groupi_n_2259 ,csa_tree_add_7_27_groupi_n_2234);
  xnor csa_tree_add_7_27_groupi_g4888__2883(csa_tree_add_7_27_groupi_n_2302 ,csa_tree_add_7_27_groupi_n_2244 ,csa_tree_add_7_27_groupi_n_2257);
  xnor csa_tree_add_7_27_groupi_g4889__2346(csa_tree_add_7_27_groupi_n_2301 ,csa_tree_add_7_27_groupi_n_2260 ,csa_tree_add_7_27_groupi_n_2236);
  xnor csa_tree_add_7_27_groupi_g4890__1666(csa_tree_add_7_27_groupi_n_2300 ,csa_tree_add_7_27_groupi_n_2245 ,csa_tree_add_7_27_groupi_n_2261);
  or csa_tree_add_7_27_groupi_g4891__7410(csa_tree_add_7_27_groupi_n_2298 ,csa_tree_add_7_27_groupi_n_2243 ,csa_tree_add_7_27_groupi_n_2256);
  or csa_tree_add_7_27_groupi_g4892__6417(csa_tree_add_7_27_groupi_n_2297 ,csa_tree_add_7_27_groupi_n_2245 ,csa_tree_add_7_27_groupi_n_2261);
  or csa_tree_add_7_27_groupi_g4893__5477(csa_tree_add_7_27_groupi_n_2296 ,csa_tree_add_7_27_groupi_n_2236 ,csa_tree_add_7_27_groupi_n_2260);
  or csa_tree_add_7_27_groupi_g4894__2398(csa_tree_add_7_27_groupi_n_2295 ,csa_tree_add_7_27_groupi_n_2234 ,csa_tree_add_7_27_groupi_n_2259);
  and csa_tree_add_7_27_groupi_g4895__5107(csa_tree_add_7_27_groupi_n_2294 ,csa_tree_add_7_27_groupi_n_2245 ,csa_tree_add_7_27_groupi_n_2261);
  and csa_tree_add_7_27_groupi_g4896__6260(csa_tree_add_7_27_groupi_n_2293 ,csa_tree_add_7_27_groupi_n_2232 ,csa_tree_add_7_27_groupi_n_2263);
  or csa_tree_add_7_27_groupi_g4897__4319(csa_tree_add_7_27_groupi_n_2292 ,csa_tree_add_7_27_groupi_n_2232 ,csa_tree_add_7_27_groupi_n_2263);
  nor csa_tree_add_7_27_groupi_g4898__8428(csa_tree_add_7_27_groupi_n_2291 ,csa_tree_add_7_27_groupi_n_2244 ,csa_tree_add_7_27_groupi_n_2257);
  and csa_tree_add_7_27_groupi_g4899__5526(csa_tree_add_7_27_groupi_n_2290 ,csa_tree_add_7_27_groupi_n_2234 ,csa_tree_add_7_27_groupi_n_2259);
  and csa_tree_add_7_27_groupi_g4900__6783(csa_tree_add_7_27_groupi_n_2289 ,csa_tree_add_7_27_groupi_n_2236 ,csa_tree_add_7_27_groupi_n_2260);
  or csa_tree_add_7_27_groupi_g4901__3680(csa_tree_add_7_27_groupi_n_2299 ,csa_tree_add_7_27_groupi_n_2273 ,csa_tree_add_7_27_groupi_n_2237);
  and csa_tree_add_7_27_groupi_g4902__1617(csa_tree_add_7_27_groupi_n_2288 ,csa_tree_add_7_27_groupi_n_2233 ,csa_tree_add_7_27_groupi_n_2258);
  and csa_tree_add_7_27_groupi_g4903__2802(csa_tree_add_7_27_groupi_n_2287 ,csa_tree_add_7_27_groupi_n_2248 ,csa_tree_add_7_27_groupi_n_2262);
  or csa_tree_add_7_27_groupi_g4904__1705(csa_tree_add_7_27_groupi_n_2286 ,csa_tree_add_7_27_groupi_n_2248 ,csa_tree_add_7_27_groupi_n_2262);
  or csa_tree_add_7_27_groupi_g4905__5122(csa_tree_add_7_27_groupi_n_2285 ,csa_tree_add_7_27_groupi_n_2264 ,csa_tree_add_7_27_groupi_n_2235);
  and csa_tree_add_7_27_groupi_g4906__8246(csa_tree_add_7_27_groupi_n_2284 ,csa_tree_add_7_27_groupi_n_2264 ,csa_tree_add_7_27_groupi_n_2235);
  or csa_tree_add_7_27_groupi_g4907__7098(csa_tree_add_7_27_groupi_n_2283 ,csa_tree_add_7_27_groupi_n_2233 ,csa_tree_add_7_27_groupi_n_2258);
  xnor csa_tree_add_7_27_groupi_g4908__6131(csa_tree_add_7_27_groupi_n_2282 ,csa_tree_add_7_27_groupi_n_2240 ,csa_tree_add_7_27_groupi_n_2227);
  xnor csa_tree_add_7_27_groupi_g4909__1881(csa_tree_add_7_27_groupi_n_2281 ,csa_tree_add_7_27_groupi_n_2241 ,csa_tree_add_7_27_groupi_n_2228);
  xnor csa_tree_add_7_27_groupi_g4910__5115(csa_tree_add_7_27_groupi_n_2280 ,csa_tree_add_7_27_groupi_n_2229 ,csa_tree_add_7_27_groupi_n_2246);
  xnor csa_tree_add_7_27_groupi_g4911__7482(csa_tree_add_7_27_groupi_n_2279 ,csa_tree_add_7_27_groupi_n_2249 ,csa_tree_add_7_27_groupi_n_2230);
  xnor csa_tree_add_7_27_groupi_g4912__4733(csa_tree_add_7_27_groupi_n_2278 ,csa_tree_add_7_27_groupi_n_2250 ,csa_tree_add_7_27_groupi_n_2208);
  xnor csa_tree_add_7_27_groupi_g4913__6161(csa_tree_add_7_27_groupi_n_2277 ,csa_tree_add_7_27_groupi_n_2221 ,csa_tree_add_7_27_groupi_n_2231);
  and csa_tree_add_7_27_groupi_g4914__9315(csa_tree_add_7_27_groupi_n_2276 ,csa_tree_add_7_27_groupi_n_2229 ,csa_tree_add_7_27_groupi_n_2247);
  or csa_tree_add_7_27_groupi_g4915__9945(csa_tree_add_7_27_groupi_n_2275 ,csa_tree_add_7_27_groupi_n_2250 ,csa_tree_add_7_27_groupi_n_2208);
  or csa_tree_add_7_27_groupi_g4916__2883(csa_tree_add_7_27_groupi_n_2274 ,csa_tree_add_7_27_groupi_n_2221 ,csa_tree_add_7_27_groupi_n_2231);
  and csa_tree_add_7_27_groupi_g4917__2346(csa_tree_add_7_27_groupi_n_2273 ,csa_tree_add_7_27_groupi_n_2251 ,csa_tree_add_7_27_groupi_n_2238);
  and csa_tree_add_7_27_groupi_g4918__1666(csa_tree_add_7_27_groupi_n_2272 ,csa_tree_add_7_27_groupi_n_2221 ,csa_tree_add_7_27_groupi_n_2231);
  nor csa_tree_add_7_27_groupi_g4919__7410(csa_tree_add_7_27_groupi_n_2271 ,csa_tree_add_7_27_groupi_n_2229 ,csa_tree_add_7_27_groupi_n_2247);
  and csa_tree_add_7_27_groupi_g4920__6417(csa_tree_add_7_27_groupi_n_2270 ,csa_tree_add_7_27_groupi_n_2250 ,csa_tree_add_7_27_groupi_n_2208);
  nor csa_tree_add_7_27_groupi_g4921__5477(csa_tree_add_7_27_groupi_n_2269 ,csa_tree_add_7_27_groupi_n_2242 ,csa_tree_add_7_27_groupi_n_2228);
  and csa_tree_add_7_27_groupi_g4922__2398(csa_tree_add_7_27_groupi_n_2268 ,csa_tree_add_7_27_groupi_n_2249 ,csa_tree_add_7_27_groupi_n_2230);
  and csa_tree_add_7_27_groupi_g4923__5107(csa_tree_add_7_27_groupi_n_2267 ,csa_tree_add_7_27_groupi_n_2242 ,csa_tree_add_7_27_groupi_n_2228);
  or csa_tree_add_7_27_groupi_g4924__6260(csa_tree_add_7_27_groupi_n_2266 ,csa_tree_add_7_27_groupi_n_2239 ,csa_tree_add_7_27_groupi_n_2227);
  nor csa_tree_add_7_27_groupi_g4925__4319(csa_tree_add_7_27_groupi_n_2265 ,csa_tree_add_7_27_groupi_n_2240 ,csa_tree_add_7_27_groupi_n_2226);
  not csa_tree_add_7_27_groupi_g4926(csa_tree_add_7_27_groupi_n_2256 ,csa_tree_add_7_27_groupi_n_2257);
  or csa_tree_add_7_27_groupi_g4927__8428(csa_tree_add_7_27_groupi_n_2255 ,csa_tree_add_7_27_groupi_n_2249 ,csa_tree_add_7_27_groupi_n_2230);
  xnor csa_tree_add_7_27_groupi_g4928__5526(n_16 ,csa_tree_add_7_27_groupi_n_2194 ,csa_tree_add_7_27_groupi_n_2203);
  xnor csa_tree_add_7_27_groupi_g4929__6783(csa_tree_add_7_27_groupi_n_2253 ,csa_tree_add_7_27_groupi_n_2223 ,csa_tree_add_7_27_groupi_n_1402);
  xnor csa_tree_add_7_27_groupi_g4930__3680(csa_tree_add_7_27_groupi_n_2252 ,csa_tree_add_7_27_groupi_n_2155 ,csa_tree_add_7_27_groupi_n_2207);
  xnor csa_tree_add_7_27_groupi_g4931__1617(csa_tree_add_7_27_groupi_n_2264 ,csa_tree_add_7_27_groupi_n_2165 ,csa_tree_add_7_27_groupi_n_2197);
  xnor csa_tree_add_7_27_groupi_g4932__2802(csa_tree_add_7_27_groupi_n_2263 ,csa_tree_add_7_27_groupi_n_2145 ,csa_tree_add_7_27_groupi_n_2196);
  xnor csa_tree_add_7_27_groupi_g4933__1705(csa_tree_add_7_27_groupi_n_2262 ,csa_tree_add_7_27_groupi_n_2141 ,csa_tree_add_7_27_groupi_n_2195);
  xnor csa_tree_add_7_27_groupi_g4934__5122(csa_tree_add_7_27_groupi_n_2261 ,csa_tree_add_7_27_groupi_n_2143 ,csa_tree_add_7_27_groupi_n_2200);
  xnor csa_tree_add_7_27_groupi_g4935__8246(csa_tree_add_7_27_groupi_n_2260 ,csa_tree_add_7_27_groupi_n_2167 ,csa_tree_add_7_27_groupi_n_2202);
  xnor csa_tree_add_7_27_groupi_g4936__7098(csa_tree_add_7_27_groupi_n_2259 ,csa_tree_add_7_27_groupi_n_2164 ,csa_tree_add_7_27_groupi_n_2201);
  xnor csa_tree_add_7_27_groupi_g4937__6131(csa_tree_add_7_27_groupi_n_2258 ,csa_tree_add_7_27_groupi_n_2166 ,csa_tree_add_7_27_groupi_n_2198);
  xnor csa_tree_add_7_27_groupi_g4938__1881(csa_tree_add_7_27_groupi_n_2257 ,csa_tree_add_7_27_groupi_n_2147 ,csa_tree_add_7_27_groupi_n_2199);
  not csa_tree_add_7_27_groupi_g4939(csa_tree_add_7_27_groupi_n_2247 ,csa_tree_add_7_27_groupi_n_2246);
  not csa_tree_add_7_27_groupi_g4940(csa_tree_add_7_27_groupi_n_2243 ,csa_tree_add_7_27_groupi_n_2244);
  not csa_tree_add_7_27_groupi_g4941(csa_tree_add_7_27_groupi_n_2242 ,csa_tree_add_7_27_groupi_n_2241);
  not csa_tree_add_7_27_groupi_g4942(csa_tree_add_7_27_groupi_n_2239 ,csa_tree_add_7_27_groupi_n_2240);
  or csa_tree_add_7_27_groupi_g4943__5115(csa_tree_add_7_27_groupi_n_2238 ,csa_tree_add_7_27_groupi_n_2155 ,csa_tree_add_7_27_groupi_n_2207);
  and csa_tree_add_7_27_groupi_g4944__7482(csa_tree_add_7_27_groupi_n_2237 ,csa_tree_add_7_27_groupi_n_2155 ,csa_tree_add_7_27_groupi_n_2207);
  or csa_tree_add_7_27_groupi_g4945__4733(csa_tree_add_7_27_groupi_n_2251 ,csa_tree_add_7_27_groupi_n_2217 ,csa_tree_add_7_27_groupi_n_2187);
  or csa_tree_add_7_27_groupi_g4946__6161(csa_tree_add_7_27_groupi_n_2250 ,csa_tree_add_7_27_groupi_n_1423 ,csa_tree_add_7_27_groupi_n_2215);
  or csa_tree_add_7_27_groupi_g4947__9315(csa_tree_add_7_27_groupi_n_2249 ,csa_tree_add_7_27_groupi_n_2216 ,csa_tree_add_7_27_groupi_n_2193);
  or csa_tree_add_7_27_groupi_g4948__9945(csa_tree_add_7_27_groupi_n_2248 ,csa_tree_add_7_27_groupi_n_2132 ,csa_tree_add_7_27_groupi_n_2219);
  or csa_tree_add_7_27_groupi_g4949__2883(csa_tree_add_7_27_groupi_n_2246 ,csa_tree_add_7_27_groupi_n_2185 ,csa_tree_add_7_27_groupi_n_2214);
  or csa_tree_add_7_27_groupi_g4950__2346(csa_tree_add_7_27_groupi_n_2245 ,csa_tree_add_7_27_groupi_n_2116 ,csa_tree_add_7_27_groupi_n_2212);
  or csa_tree_add_7_27_groupi_g4951__1666(csa_tree_add_7_27_groupi_n_2244 ,csa_tree_add_7_27_groupi_n_2124 ,csa_tree_add_7_27_groupi_n_2210);
  or csa_tree_add_7_27_groupi_g4952__7410(csa_tree_add_7_27_groupi_n_2241 ,csa_tree_add_7_27_groupi_n_2175 ,csa_tree_add_7_27_groupi_n_2211);
  or csa_tree_add_7_27_groupi_g4953__6417(csa_tree_add_7_27_groupi_n_2240 ,csa_tree_add_7_27_groupi_n_2173 ,csa_tree_add_7_27_groupi_n_2209);
  not csa_tree_add_7_27_groupi_g4954(csa_tree_add_7_27_groupi_n_2226 ,csa_tree_add_7_27_groupi_n_2227);
  or csa_tree_add_7_27_groupi_g4955__5477(csa_tree_add_7_27_groupi_n_2225 ,csa_tree_add_7_27_groupi_n_1401 ,csa_tree_add_7_27_groupi_n_2222);
  nor csa_tree_add_7_27_groupi_g4956__2398(csa_tree_add_7_27_groupi_n_2224 ,csa_tree_add_7_27_groupi_n_1402 ,csa_tree_add_7_27_groupi_n_2223);
  and csa_tree_add_7_27_groupi_g4957__5107(csa_tree_add_7_27_groupi_n_2236 ,csa_tree_add_7_27_groupi_n_2170 ,csa_tree_add_7_27_groupi_n_2220);
  or csa_tree_add_7_27_groupi_g4958__6260(csa_tree_add_7_27_groupi_n_2235 ,csa_tree_add_7_27_groupi_n_2206 ,csa_tree_add_7_27_groupi_n_2176);
  and csa_tree_add_7_27_groupi_g4959__4319(csa_tree_add_7_27_groupi_n_2234 ,csa_tree_add_7_27_groupi_n_2183 ,csa_tree_add_7_27_groupi_n_2218);
  and csa_tree_add_7_27_groupi_g4960__8428(csa_tree_add_7_27_groupi_n_2233 ,csa_tree_add_7_27_groupi_n_2172 ,csa_tree_add_7_27_groupi_n_2204);
  or csa_tree_add_7_27_groupi_g4961__5526(csa_tree_add_7_27_groupi_n_2232 ,csa_tree_add_7_27_groupi_n_2117 ,csa_tree_add_7_27_groupi_n_2213);
  xnor csa_tree_add_7_27_groupi_g4962__6783(csa_tree_add_7_27_groupi_n_2231 ,csa_tree_add_7_27_groupi_n_2179 ,csa_tree_add_7_27_groupi_n_2140);
  xnor csa_tree_add_7_27_groupi_g4963__3680(csa_tree_add_7_27_groupi_n_2230 ,csa_tree_add_7_27_groupi_n_2180 ,csa_tree_add_7_27_groupi_n_2138);
  xnor csa_tree_add_7_27_groupi_g4964__1617(csa_tree_add_7_27_groupi_n_2229 ,csa_tree_add_7_27_groupi_n_2177 ,csa_tree_add_7_27_groupi_n_1432);
  xnor csa_tree_add_7_27_groupi_g4965__2802(csa_tree_add_7_27_groupi_n_2228 ,csa_tree_add_7_27_groupi_n_2181 ,csa_tree_add_7_27_groupi_n_2137);
  xnor csa_tree_add_7_27_groupi_g4966__1705(csa_tree_add_7_27_groupi_n_2227 ,csa_tree_add_7_27_groupi_n_2178 ,csa_tree_add_7_27_groupi_n_2139);
  not csa_tree_add_7_27_groupi_g4967(csa_tree_add_7_27_groupi_n_2222 ,csa_tree_add_7_27_groupi_n_2223);
  or csa_tree_add_7_27_groupi_g4968__5122(csa_tree_add_7_27_groupi_n_2220 ,csa_tree_add_7_27_groupi_n_2182 ,csa_tree_add_7_27_groupi_n_2148);
  and csa_tree_add_7_27_groupi_g4969__8246(csa_tree_add_7_27_groupi_n_2219 ,csa_tree_add_7_27_groupi_n_2179 ,csa_tree_add_7_27_groupi_n_2133);
  or csa_tree_add_7_27_groupi_g4970__7098(csa_tree_add_7_27_groupi_n_2218 ,csa_tree_add_7_27_groupi_n_2186 ,csa_tree_add_7_27_groupi_n_2149);
  and csa_tree_add_7_27_groupi_g4971__6131(csa_tree_add_7_27_groupi_n_2217 ,csa_tree_add_7_27_groupi_n_2189 ,csa_tree_add_7_27_groupi_n_2194);
  and csa_tree_add_7_27_groupi_g4972__1881(csa_tree_add_7_27_groupi_n_2216 ,csa_tree_add_7_27_groupi_n_2165 ,csa_tree_add_7_27_groupi_n_2192);
  and csa_tree_add_7_27_groupi_g4973__5115(csa_tree_add_7_27_groupi_n_2215 ,csa_tree_add_7_27_groupi_n_1426 ,csa_tree_add_7_27_groupi_n_2177);
  and csa_tree_add_7_27_groupi_g4974__7482(csa_tree_add_7_27_groupi_n_2214 ,csa_tree_add_7_27_groupi_n_2164 ,csa_tree_add_7_27_groupi_n_2184);
  and csa_tree_add_7_27_groupi_g4975__4733(csa_tree_add_7_27_groupi_n_2213 ,csa_tree_add_7_27_groupi_n_2180 ,csa_tree_add_7_27_groupi_n_2121);
  and csa_tree_add_7_27_groupi_g4976__6161(csa_tree_add_7_27_groupi_n_2212 ,csa_tree_add_7_27_groupi_n_2181 ,csa_tree_add_7_27_groupi_n_2115);
  and csa_tree_add_7_27_groupi_g4977__9315(csa_tree_add_7_27_groupi_n_2211 ,csa_tree_add_7_27_groupi_n_2166 ,csa_tree_add_7_27_groupi_n_2174);
  and csa_tree_add_7_27_groupi_g4978__9945(csa_tree_add_7_27_groupi_n_2210 ,csa_tree_add_7_27_groupi_n_2178 ,csa_tree_add_7_27_groupi_n_2123);
  and csa_tree_add_7_27_groupi_g4979__2883(csa_tree_add_7_27_groupi_n_2209 ,csa_tree_add_7_27_groupi_n_2167 ,csa_tree_add_7_27_groupi_n_2171);
  and csa_tree_add_7_27_groupi_g4980__2346(csa_tree_add_7_27_groupi_n_2223 ,csa_tree_add_7_27_groupi_n_1273 ,csa_tree_add_7_27_groupi_n_2191);
  or csa_tree_add_7_27_groupi_g4981__1666(csa_tree_add_7_27_groupi_n_2221 ,csa_tree_add_7_27_groupi_n_2066 ,csa_tree_add_7_27_groupi_n_2190);
  nor csa_tree_add_7_27_groupi_g4982__7410(csa_tree_add_7_27_groupi_n_2206 ,csa_tree_add_7_27_groupi_n_2188 ,csa_tree_add_7_27_groupi_n_2152);
  xnor csa_tree_add_7_27_groupi_g4983__6417(n_15 ,csa_tree_add_7_27_groupi_n_2135 ,csa_tree_add_7_27_groupi_n_2136);
  or csa_tree_add_7_27_groupi_g4984__5477(csa_tree_add_7_27_groupi_n_2204 ,csa_tree_add_7_27_groupi_n_2169 ,csa_tree_add_7_27_groupi_n_2150);
  xnor csa_tree_add_7_27_groupi_g4985__2398(csa_tree_add_7_27_groupi_n_2203 ,csa_tree_add_7_27_groupi_n_2156 ,csa_tree_add_7_27_groupi_n_2108);
  xnor csa_tree_add_7_27_groupi_g4986__5107(csa_tree_add_7_27_groupi_n_2202 ,csa_tree_add_7_27_groupi_n_2159 ,csa_tree_add_7_27_groupi_n_2079);
  xnor csa_tree_add_7_27_groupi_g4987__6260(csa_tree_add_7_27_groupi_n_2201 ,csa_tree_add_7_27_groupi_n_1410 ,csa_tree_add_7_27_groupi_n_2163);
  xnor csa_tree_add_7_27_groupi_g4988__4319(csa_tree_add_7_27_groupi_n_2200 ,csa_tree_add_7_27_groupi_n_2112 ,csa_tree_add_7_27_groupi_n_2148);
  xnor csa_tree_add_7_27_groupi_g4989__8428(csa_tree_add_7_27_groupi_n_2199 ,csa_tree_add_7_27_groupi_n_2114 ,csa_tree_add_7_27_groupi_n_2149);
  xnor csa_tree_add_7_27_groupi_g4990__5526(csa_tree_add_7_27_groupi_n_2198 ,csa_tree_add_7_27_groupi_n_2161 ,csa_tree_add_7_27_groupi_n_2081);
  xnor csa_tree_add_7_27_groupi_g4991__6783(csa_tree_add_7_27_groupi_n_2197 ,csa_tree_add_7_27_groupi_n_2157 ,csa_tree_add_7_27_groupi_n_2087);
  xnor csa_tree_add_7_27_groupi_g4992__3680(csa_tree_add_7_27_groupi_n_2196 ,csa_tree_add_7_27_groupi_n_2110 ,csa_tree_add_7_27_groupi_n_2150);
  xnor csa_tree_add_7_27_groupi_g4993__1617(csa_tree_add_7_27_groupi_n_2195 ,csa_tree_add_7_27_groupi_n_2106 ,csa_tree_add_7_27_groupi_n_2152);
  xnor csa_tree_add_7_27_groupi_g4994__2802(csa_tree_add_7_27_groupi_n_2208 ,csa_tree_add_7_27_groupi_n_2151 ,csa_tree_add_7_27_groupi_n_1307);
  xnor csa_tree_add_7_27_groupi_g4995__1705(csa_tree_add_7_27_groupi_n_2207 ,csa_tree_add_7_27_groupi_n_2168 ,csa_tree_add_7_27_groupi_n_2071);
  and csa_tree_add_7_27_groupi_g4996__5122(csa_tree_add_7_27_groupi_n_2193 ,csa_tree_add_7_27_groupi_n_2157 ,csa_tree_add_7_27_groupi_n_2087);
  or csa_tree_add_7_27_groupi_g4997__8246(csa_tree_add_7_27_groupi_n_2192 ,csa_tree_add_7_27_groupi_n_2157 ,csa_tree_add_7_27_groupi_n_2087);
  or csa_tree_add_7_27_groupi_g4998__7098(csa_tree_add_7_27_groupi_n_2191 ,csa_tree_add_7_27_groupi_n_1278 ,csa_tree_add_7_27_groupi_n_2151);
  and csa_tree_add_7_27_groupi_g4999__6131(csa_tree_add_7_27_groupi_n_2190 ,csa_tree_add_7_27_groupi_n_2168 ,csa_tree_add_7_27_groupi_n_2064);
  or csa_tree_add_7_27_groupi_g5000__1881(csa_tree_add_7_27_groupi_n_2189 ,csa_tree_add_7_27_groupi_n_2156 ,csa_tree_add_7_27_groupi_n_2108);
  and csa_tree_add_7_27_groupi_g5001__5115(csa_tree_add_7_27_groupi_n_2188 ,csa_tree_add_7_27_groupi_n_2141 ,csa_tree_add_7_27_groupi_n_2107);
  and csa_tree_add_7_27_groupi_g5002__7482(csa_tree_add_7_27_groupi_n_2187 ,csa_tree_add_7_27_groupi_n_2156 ,csa_tree_add_7_27_groupi_n_2108);
  nor csa_tree_add_7_27_groupi_g5003__4733(csa_tree_add_7_27_groupi_n_2186 ,csa_tree_add_7_27_groupi_n_2146 ,csa_tree_add_7_27_groupi_n_2114);
  nor csa_tree_add_7_27_groupi_g5004__6161(csa_tree_add_7_27_groupi_n_2185 ,csa_tree_add_7_27_groupi_n_1410 ,csa_tree_add_7_27_groupi_n_2162);
  or csa_tree_add_7_27_groupi_g5005__9315(csa_tree_add_7_27_groupi_n_2184 ,csa_tree_add_7_27_groupi_n_1409 ,csa_tree_add_7_27_groupi_n_2163);
  or csa_tree_add_7_27_groupi_g5006__9945(csa_tree_add_7_27_groupi_n_2183 ,csa_tree_add_7_27_groupi_n_2147 ,csa_tree_add_7_27_groupi_n_2113);
  nor csa_tree_add_7_27_groupi_g5007__2883(csa_tree_add_7_27_groupi_n_2182 ,csa_tree_add_7_27_groupi_n_2142 ,csa_tree_add_7_27_groupi_n_2112);
  or csa_tree_add_7_27_groupi_g5008__2346(csa_tree_add_7_27_groupi_n_2194 ,csa_tree_add_7_27_groupi_n_2154 ,csa_tree_add_7_27_groupi_n_2134);
  nor csa_tree_add_7_27_groupi_g5009__1666(csa_tree_add_7_27_groupi_n_2176 ,csa_tree_add_7_27_groupi_n_2141 ,csa_tree_add_7_27_groupi_n_2107);
  nor csa_tree_add_7_27_groupi_g5010__7410(csa_tree_add_7_27_groupi_n_2175 ,csa_tree_add_7_27_groupi_n_2160 ,csa_tree_add_7_27_groupi_n_2081);
  or csa_tree_add_7_27_groupi_g5011__6417(csa_tree_add_7_27_groupi_n_2174 ,csa_tree_add_7_27_groupi_n_2161 ,csa_tree_add_7_27_groupi_n_2080);
  nor csa_tree_add_7_27_groupi_g5012__5477(csa_tree_add_7_27_groupi_n_2173 ,csa_tree_add_7_27_groupi_n_2158 ,csa_tree_add_7_27_groupi_n_2079);
  or csa_tree_add_7_27_groupi_g5013__2398(csa_tree_add_7_27_groupi_n_2172 ,csa_tree_add_7_27_groupi_n_2145 ,csa_tree_add_7_27_groupi_n_2109);
  or csa_tree_add_7_27_groupi_g5014__5107(csa_tree_add_7_27_groupi_n_2171 ,csa_tree_add_7_27_groupi_n_2159 ,csa_tree_add_7_27_groupi_n_2078);
  or csa_tree_add_7_27_groupi_g5015__6260(csa_tree_add_7_27_groupi_n_2170 ,csa_tree_add_7_27_groupi_n_2143 ,csa_tree_add_7_27_groupi_n_2111);
  nor csa_tree_add_7_27_groupi_g5016__4319(csa_tree_add_7_27_groupi_n_2169 ,csa_tree_add_7_27_groupi_n_2144 ,csa_tree_add_7_27_groupi_n_2110);
  xnor csa_tree_add_7_27_groupi_g5017__8428(csa_tree_add_7_27_groupi_n_2181 ,csa_tree_add_7_27_groupi_n_2126 ,in2[8]);
  xnor csa_tree_add_7_27_groupi_g5018__5526(csa_tree_add_7_27_groupi_n_2180 ,csa_tree_add_7_27_groupi_n_2127 ,in2[5]);
  xnor csa_tree_add_7_27_groupi_g5019__6783(csa_tree_add_7_27_groupi_n_2179 ,csa_tree_add_7_27_groupi_n_2130 ,in2[2]);
  xnor csa_tree_add_7_27_groupi_g5020__3680(csa_tree_add_7_27_groupi_n_2178 ,csa_tree_add_7_27_groupi_n_2128 ,in2[11]);
  xnor csa_tree_add_7_27_groupi_g5021__1617(csa_tree_add_7_27_groupi_n_2177 ,csa_tree_add_7_27_groupi_n_2129 ,in2[14]);
  not csa_tree_add_7_27_groupi_g5022(csa_tree_add_7_27_groupi_n_2162 ,csa_tree_add_7_27_groupi_n_2163);
  not csa_tree_add_7_27_groupi_g5023(csa_tree_add_7_27_groupi_n_2160 ,csa_tree_add_7_27_groupi_n_2161);
  not csa_tree_add_7_27_groupi_g5024(csa_tree_add_7_27_groupi_n_2158 ,csa_tree_add_7_27_groupi_n_2159);
  and csa_tree_add_7_27_groupi_g5025__2802(csa_tree_add_7_27_groupi_n_2154 ,csa_tree_add_7_27_groupi_n_2135 ,csa_tree_add_7_27_groupi_n_2131);
  xnor csa_tree_add_7_27_groupi_g5026__1705(n_14 ,csa_tree_add_7_27_groupi_n_2069 ,csa_tree_add_7_27_groupi_n_2070);
  xnor csa_tree_add_7_27_groupi_g5027__5122(csa_tree_add_7_27_groupi_n_2168 ,csa_tree_add_7_27_groupi_n_2101 ,in2[2]);
  or csa_tree_add_7_27_groupi_g5028__8246(csa_tree_add_7_27_groupi_n_2167 ,csa_tree_add_7_27_groupi_n_1990 ,csa_tree_add_7_27_groupi_n_2118);
  or csa_tree_add_7_27_groupi_g5029__7098(csa_tree_add_7_27_groupi_n_2166 ,csa_tree_add_7_27_groupi_n_1984 ,csa_tree_add_7_27_groupi_n_2119);
  or csa_tree_add_7_27_groupi_g5030__6131(csa_tree_add_7_27_groupi_n_2165 ,csa_tree_add_7_27_groupi_n_1988 ,csa_tree_add_7_27_groupi_n_2125);
  or csa_tree_add_7_27_groupi_g5031__1881(csa_tree_add_7_27_groupi_n_2164 ,csa_tree_add_7_27_groupi_n_1176 ,csa_tree_add_7_27_groupi_n_2122);
  xnor csa_tree_add_7_27_groupi_g5032__5115(csa_tree_add_7_27_groupi_n_2163 ,csa_tree_add_7_27_groupi_n_2099 ,in2[14]);
  xnor csa_tree_add_7_27_groupi_g5033__7482(csa_tree_add_7_27_groupi_n_2161 ,csa_tree_add_7_27_groupi_n_2102 ,in2[8]);
  xnor csa_tree_add_7_27_groupi_g5034__4733(csa_tree_add_7_27_groupi_n_2159 ,csa_tree_add_7_27_groupi_n_2098 ,in2[11]);
  xnor csa_tree_add_7_27_groupi_g5035__6161(csa_tree_add_7_27_groupi_n_2157 ,csa_tree_add_7_27_groupi_n_2096 ,in2[5]);
  xnor csa_tree_add_7_27_groupi_g5036__9315(csa_tree_add_7_27_groupi_n_2156 ,csa_tree_add_7_27_groupi_n_2090 ,csa_tree_add_7_27_groupi_n_2015);
  or csa_tree_add_7_27_groupi_g5037__9945(csa_tree_add_7_27_groupi_n_2155 ,csa_tree_add_7_27_groupi_n_1999 ,csa_tree_add_7_27_groupi_n_2120);
  not csa_tree_add_7_27_groupi_g5038(csa_tree_add_7_27_groupi_n_2146 ,csa_tree_add_7_27_groupi_n_2147);
  not csa_tree_add_7_27_groupi_g5039(csa_tree_add_7_27_groupi_n_2144 ,csa_tree_add_7_27_groupi_n_2145);
  not csa_tree_add_7_27_groupi_g5040(csa_tree_add_7_27_groupi_n_2142 ,csa_tree_add_7_27_groupi_n_2143);
  xnor csa_tree_add_7_27_groupi_g5041__2883(csa_tree_add_7_27_groupi_n_2140 ,csa_tree_add_7_27_groupi_n_2042 ,csa_tree_add_7_27_groupi_n_2077);
  xnor csa_tree_add_7_27_groupi_g5042__2346(csa_tree_add_7_27_groupi_n_2139 ,csa_tree_add_7_27_groupi_n_2085 ,csa_tree_add_7_27_groupi_n_2055);
  xnor csa_tree_add_7_27_groupi_g5043__1666(csa_tree_add_7_27_groupi_n_2138 ,csa_tree_add_7_27_groupi_n_2068 ,csa_tree_add_7_27_groupi_n_2086);
  xnor csa_tree_add_7_27_groupi_g5044__7410(csa_tree_add_7_27_groupi_n_2137 ,csa_tree_add_7_27_groupi_n_2057 ,csa_tree_add_7_27_groupi_n_2083);
  xnor csa_tree_add_7_27_groupi_g5045__6417(csa_tree_add_7_27_groupi_n_2136 ,csa_tree_add_7_27_groupi_n_2076 ,csa_tree_add_7_27_groupi_n_2043);
  xnor csa_tree_add_7_27_groupi_g5046__5477(csa_tree_add_7_27_groupi_n_2152 ,csa_tree_add_7_27_groupi_n_2089 ,csa_tree_add_7_27_groupi_n_2012);
  xnor csa_tree_add_7_27_groupi_g5047__2398(csa_tree_add_7_27_groupi_n_2151 ,csa_tree_add_7_27_groupi_n_2097 ,in2[14]);
  xnor csa_tree_add_7_27_groupi_g5048__5107(csa_tree_add_7_27_groupi_n_2150 ,csa_tree_add_7_27_groupi_n_2088 ,csa_tree_add_7_27_groupi_n_2011);
  xnor csa_tree_add_7_27_groupi_g5049__6260(csa_tree_add_7_27_groupi_n_2149 ,csa_tree_add_7_27_groupi_n_2091 ,csa_tree_add_7_27_groupi_n_1301);
  xnor csa_tree_add_7_27_groupi_g5050__4319(csa_tree_add_7_27_groupi_n_2148 ,csa_tree_add_7_27_groupi_n_2092 ,csa_tree_add_7_27_groupi_n_2010);
  xnor csa_tree_add_7_27_groupi_g5051__8428(csa_tree_add_7_27_groupi_n_2147 ,csa_tree_add_7_27_groupi_n_2093 ,in2[11]);
  xnor csa_tree_add_7_27_groupi_g5052__5526(csa_tree_add_7_27_groupi_n_2145 ,csa_tree_add_7_27_groupi_n_2095 ,in2[5]);
  xnor csa_tree_add_7_27_groupi_g5053__6783(csa_tree_add_7_27_groupi_n_2143 ,csa_tree_add_7_27_groupi_n_2094 ,in2[8]);
  xnor csa_tree_add_7_27_groupi_g5054__3680(csa_tree_add_7_27_groupi_n_2141 ,csa_tree_add_7_27_groupi_n_2100 ,in2[2]);
  and csa_tree_add_7_27_groupi_g5055__1617(csa_tree_add_7_27_groupi_n_2134 ,csa_tree_add_7_27_groupi_n_2076 ,csa_tree_add_7_27_groupi_n_2043);
  or csa_tree_add_7_27_groupi_g5056__2802(csa_tree_add_7_27_groupi_n_2133 ,csa_tree_add_7_27_groupi_n_2042 ,csa_tree_add_7_27_groupi_n_2077);
  and csa_tree_add_7_27_groupi_g5057__1705(csa_tree_add_7_27_groupi_n_2132 ,csa_tree_add_7_27_groupi_n_2042 ,csa_tree_add_7_27_groupi_n_2077);
  or csa_tree_add_7_27_groupi_g5058__5122(csa_tree_add_7_27_groupi_n_2131 ,csa_tree_add_7_27_groupi_n_2076 ,csa_tree_add_7_27_groupi_n_2043);
  nor csa_tree_add_7_27_groupi_g5059__8246(csa_tree_add_7_27_groupi_n_2130 ,csa_tree_add_7_27_groupi_n_1135 ,csa_tree_add_7_27_groupi_n_2104);
  nor csa_tree_add_7_27_groupi_g5060__7098(csa_tree_add_7_27_groupi_n_2129 ,csa_tree_add_7_27_groupi_n_1344 ,csa_tree_add_7_27_groupi_n_2072);
  nor csa_tree_add_7_27_groupi_g5061__6131(csa_tree_add_7_27_groupi_n_2128 ,csa_tree_add_7_27_groupi_n_1349 ,csa_tree_add_7_27_groupi_n_2075);
  nor csa_tree_add_7_27_groupi_g5062__1881(csa_tree_add_7_27_groupi_n_2127 ,csa_tree_add_7_27_groupi_n_1366 ,csa_tree_add_7_27_groupi_n_2105);
  nor csa_tree_add_7_27_groupi_g5063__5115(csa_tree_add_7_27_groupi_n_2126 ,csa_tree_add_7_27_groupi_n_1347 ,csa_tree_add_7_27_groupi_n_2074);
  or csa_tree_add_7_27_groupi_g5064__7482(csa_tree_add_7_27_groupi_n_2135 ,csa_tree_add_7_27_groupi_n_2067 ,csa_tree_add_7_27_groupi_n_2103);
  and csa_tree_add_7_27_groupi_g5065__4733(csa_tree_add_7_27_groupi_n_2125 ,csa_tree_add_7_27_groupi_n_2089 ,csa_tree_add_7_27_groupi_n_1987);
  nor csa_tree_add_7_27_groupi_g5066__6161(csa_tree_add_7_27_groupi_n_2124 ,csa_tree_add_7_27_groupi_n_2085 ,csa_tree_add_7_27_groupi_n_2054);
  or csa_tree_add_7_27_groupi_g5067__9315(csa_tree_add_7_27_groupi_n_2123 ,csa_tree_add_7_27_groupi_n_2084 ,csa_tree_add_7_27_groupi_n_2055);
  and csa_tree_add_7_27_groupi_g5068__9945(csa_tree_add_7_27_groupi_n_2122 ,csa_tree_add_7_27_groupi_n_1177 ,csa_tree_add_7_27_groupi_n_2091);
  or csa_tree_add_7_27_groupi_g5069__2883(csa_tree_add_7_27_groupi_n_2121 ,csa_tree_add_7_27_groupi_n_2068 ,csa_tree_add_7_27_groupi_n_2086);
  and csa_tree_add_7_27_groupi_g5070__2346(csa_tree_add_7_27_groupi_n_2120 ,csa_tree_add_7_27_groupi_n_2090 ,csa_tree_add_7_27_groupi_n_2002);
  and csa_tree_add_7_27_groupi_g5071__1666(csa_tree_add_7_27_groupi_n_2119 ,csa_tree_add_7_27_groupi_n_2088 ,csa_tree_add_7_27_groupi_n_1983);
  and csa_tree_add_7_27_groupi_g5072__7410(csa_tree_add_7_27_groupi_n_2118 ,csa_tree_add_7_27_groupi_n_2092 ,csa_tree_add_7_27_groupi_n_1989);
  and csa_tree_add_7_27_groupi_g5073__6417(csa_tree_add_7_27_groupi_n_2117 ,csa_tree_add_7_27_groupi_n_2068 ,csa_tree_add_7_27_groupi_n_2086);
  nor csa_tree_add_7_27_groupi_g5074__5477(csa_tree_add_7_27_groupi_n_2116 ,csa_tree_add_7_27_groupi_n_2056 ,csa_tree_add_7_27_groupi_n_2083);
  or csa_tree_add_7_27_groupi_g5075__2398(csa_tree_add_7_27_groupi_n_2115 ,csa_tree_add_7_27_groupi_n_2057 ,csa_tree_add_7_27_groupi_n_2082);
  not csa_tree_add_7_27_groupi_g5076(csa_tree_add_7_27_groupi_n_2113 ,csa_tree_add_7_27_groupi_n_2114);
  not csa_tree_add_7_27_groupi_g5077(csa_tree_add_7_27_groupi_n_2111 ,csa_tree_add_7_27_groupi_n_2112);
  not csa_tree_add_7_27_groupi_g5078(csa_tree_add_7_27_groupi_n_2109 ,csa_tree_add_7_27_groupi_n_2110);
  not csa_tree_add_7_27_groupi_g5079(csa_tree_add_7_27_groupi_n_2107 ,csa_tree_add_7_27_groupi_n_2106);
  nor csa_tree_add_7_27_groupi_g5080__5107(csa_tree_add_7_27_groupi_n_2105 ,csa_tree_add_7_27_groupi_n_465 ,csa_tree_add_7_27_groupi_n_509);
  nor csa_tree_add_7_27_groupi_g5081__6260(csa_tree_add_7_27_groupi_n_2104 ,csa_tree_add_7_27_groupi_n_462 ,csa_tree_add_7_27_groupi_n_2053);
  and csa_tree_add_7_27_groupi_g5082__4319(csa_tree_add_7_27_groupi_n_2103 ,csa_tree_add_7_27_groupi_n_2060 ,csa_tree_add_7_27_groupi_n_2069);
  nor csa_tree_add_7_27_groupi_g5083__8428(csa_tree_add_7_27_groupi_n_2102 ,csa_tree_add_7_27_groupi_n_1328 ,csa_tree_add_7_27_groupi_n_2065);
  nor csa_tree_add_7_27_groupi_g5084__5526(csa_tree_add_7_27_groupi_n_2101 ,csa_tree_add_7_27_groupi_n_1118 ,csa_tree_add_7_27_groupi_n_2047);
  or csa_tree_add_7_27_groupi_g5085__6783(csa_tree_add_7_27_groupi_n_2100 ,csa_tree_add_7_27_groupi_n_957 ,csa_tree_add_7_27_groupi_n_2052);
  nor csa_tree_add_7_27_groupi_g5086__3680(csa_tree_add_7_27_groupi_n_2099 ,csa_tree_add_7_27_groupi_n_1321 ,csa_tree_add_7_27_groupi_n_2059);
  nor csa_tree_add_7_27_groupi_g5087__1617(csa_tree_add_7_27_groupi_n_2098 ,csa_tree_add_7_27_groupi_n_1330 ,csa_tree_add_7_27_groupi_n_2063);
  or csa_tree_add_7_27_groupi_g5088__2802(csa_tree_add_7_27_groupi_n_2097 ,csa_tree_add_7_27_groupi_n_1253 ,csa_tree_add_7_27_groupi_n_2044);
  nor csa_tree_add_7_27_groupi_g5089__1705(csa_tree_add_7_27_groupi_n_2096 ,csa_tree_add_7_27_groupi_n_1293 ,csa_tree_add_7_27_groupi_n_2058);
  or csa_tree_add_7_27_groupi_g5090__5122(csa_tree_add_7_27_groupi_n_2095 ,csa_tree_add_7_27_groupi_n_1249 ,csa_tree_add_7_27_groupi_n_2045);
  or csa_tree_add_7_27_groupi_g5091__8246(csa_tree_add_7_27_groupi_n_2094 ,csa_tree_add_7_27_groupi_n_1254 ,csa_tree_add_7_27_groupi_n_2048);
  or csa_tree_add_7_27_groupi_g5092__7098(csa_tree_add_7_27_groupi_n_2093 ,csa_tree_add_7_27_groupi_n_1256 ,csa_tree_add_7_27_groupi_n_2051);
  or csa_tree_add_7_27_groupi_g5093__6131(csa_tree_add_7_27_groupi_n_2114 ,csa_tree_add_7_27_groupi_n_1424 ,csa_tree_add_7_27_groupi_n_2046);
  or csa_tree_add_7_27_groupi_g5094__1881(csa_tree_add_7_27_groupi_n_2112 ,csa_tree_add_7_27_groupi_n_1926 ,csa_tree_add_7_27_groupi_n_2050);
  or csa_tree_add_7_27_groupi_g5095__5115(csa_tree_add_7_27_groupi_n_2110 ,csa_tree_add_7_27_groupi_n_1924 ,csa_tree_add_7_27_groupi_n_2049);
  or csa_tree_add_7_27_groupi_g5096__7482(csa_tree_add_7_27_groupi_n_2108 ,csa_tree_add_7_27_groupi_n_1935 ,csa_tree_add_7_27_groupi_n_2062);
  or csa_tree_add_7_27_groupi_g5097__4733(csa_tree_add_7_27_groupi_n_2106 ,csa_tree_add_7_27_groupi_n_1940 ,csa_tree_add_7_27_groupi_n_2061);
  not csa_tree_add_7_27_groupi_g5098(csa_tree_add_7_27_groupi_n_2084 ,csa_tree_add_7_27_groupi_n_2085);
  not csa_tree_add_7_27_groupi_g5099(csa_tree_add_7_27_groupi_n_2082 ,csa_tree_add_7_27_groupi_n_2083);
  not csa_tree_add_7_27_groupi_g5100(csa_tree_add_7_27_groupi_n_2080 ,csa_tree_add_7_27_groupi_n_2081);
  not csa_tree_add_7_27_groupi_g5101(csa_tree_add_7_27_groupi_n_2078 ,csa_tree_add_7_27_groupi_n_2079);
  nor csa_tree_add_7_27_groupi_g5102__6161(csa_tree_add_7_27_groupi_n_2075 ,csa_tree_add_7_27_groupi_n_456 ,csa_tree_add_7_27_groupi_n_509);
  nor csa_tree_add_7_27_groupi_g5103__9315(csa_tree_add_7_27_groupi_n_2074 ,csa_tree_add_7_27_groupi_n_459 ,csa_tree_add_7_27_groupi_n_2053);
  xnor csa_tree_add_7_27_groupi_g5104__9945(n_13 ,csa_tree_add_7_27_groupi_n_2006 ,csa_tree_add_7_27_groupi_n_2014);
  nor csa_tree_add_7_27_groupi_g5105__2883(csa_tree_add_7_27_groupi_n_2072 ,csa_tree_add_7_27_groupi_n_468 ,csa_tree_add_7_27_groupi_n_508);
  xnor csa_tree_add_7_27_groupi_g5106__2346(csa_tree_add_7_27_groupi_n_2071 ,csa_tree_add_7_27_groupi_n_1977 ,csa_tree_add_7_27_groupi_n_2020);
  xnor csa_tree_add_7_27_groupi_g5107__1666(csa_tree_add_7_27_groupi_n_2070 ,csa_tree_add_7_27_groupi_n_1978 ,csa_tree_add_7_27_groupi_n_2019);
  xnor csa_tree_add_7_27_groupi_g5108__7410(csa_tree_add_7_27_groupi_n_2092 ,csa_tree_add_7_27_groupi_n_2028 ,in2[11]);
  xnor csa_tree_add_7_27_groupi_g5109__6417(csa_tree_add_7_27_groupi_n_2091 ,csa_tree_add_7_27_groupi_n_2029 ,in2[14]);
  xnor csa_tree_add_7_27_groupi_g5110__5477(csa_tree_add_7_27_groupi_n_2090 ,csa_tree_add_7_27_groupi_n_2027 ,in2[2]);
  xnor csa_tree_add_7_27_groupi_g5111__2398(csa_tree_add_7_27_groupi_n_2089 ,csa_tree_add_7_27_groupi_n_2030 ,in2[5]);
  xnor csa_tree_add_7_27_groupi_g5112__5107(csa_tree_add_7_27_groupi_n_2088 ,csa_tree_add_7_27_groupi_n_2026 ,in2[8]);
  xnor csa_tree_add_7_27_groupi_g5113__6260(csa_tree_add_7_27_groupi_n_2087 ,csa_tree_add_7_27_groupi_n_1980 ,csa_tree_add_7_27_groupi_n_2013);
  xnor csa_tree_add_7_27_groupi_g5114__4319(csa_tree_add_7_27_groupi_n_2086 ,csa_tree_add_7_27_groupi_n_2021 ,csa_tree_add_7_27_groupi_n_1946);
  xnor csa_tree_add_7_27_groupi_g5115__8428(csa_tree_add_7_27_groupi_n_2085 ,csa_tree_add_7_27_groupi_n_2022 ,csa_tree_add_7_27_groupi_n_1434);
  xnor csa_tree_add_7_27_groupi_g5116__5526(csa_tree_add_7_27_groupi_n_2083 ,csa_tree_add_7_27_groupi_n_2023 ,csa_tree_add_7_27_groupi_n_1945);
  xnor csa_tree_add_7_27_groupi_g5117__6783(csa_tree_add_7_27_groupi_n_2081 ,csa_tree_add_7_27_groupi_n_1981 ,csa_tree_add_7_27_groupi_n_2016);
  xnor csa_tree_add_7_27_groupi_g5118__3680(csa_tree_add_7_27_groupi_n_2079 ,csa_tree_add_7_27_groupi_n_1979 ,csa_tree_add_7_27_groupi_n_2009);
  xnor csa_tree_add_7_27_groupi_g5119__1617(csa_tree_add_7_27_groupi_n_2077 ,csa_tree_add_7_27_groupi_n_2025 ,csa_tree_add_7_27_groupi_n_1948);
  xnor csa_tree_add_7_27_groupi_g5120__2802(csa_tree_add_7_27_groupi_n_2076 ,csa_tree_add_7_27_groupi_n_2024 ,csa_tree_add_7_27_groupi_n_1949);
  and csa_tree_add_7_27_groupi_g5121__1705(csa_tree_add_7_27_groupi_n_2067 ,csa_tree_add_7_27_groupi_n_1978 ,csa_tree_add_7_27_groupi_n_2019);
  and csa_tree_add_7_27_groupi_g5122__5122(csa_tree_add_7_27_groupi_n_2066 ,csa_tree_add_7_27_groupi_n_1977 ,csa_tree_add_7_27_groupi_n_2020);
  or csa_tree_add_7_27_groupi_g5123__8246(csa_tree_add_7_27_groupi_n_2065 ,csa_tree_add_7_27_groupi_n_1137 ,csa_tree_add_7_27_groupi_n_2036);
  or csa_tree_add_7_27_groupi_g5124__7098(csa_tree_add_7_27_groupi_n_2064 ,csa_tree_add_7_27_groupi_n_1977 ,csa_tree_add_7_27_groupi_n_2020);
  or csa_tree_add_7_27_groupi_g5125__6131(csa_tree_add_7_27_groupi_n_2063 ,csa_tree_add_7_27_groupi_n_1123 ,csa_tree_add_7_27_groupi_n_2018);
  and csa_tree_add_7_27_groupi_g5126__1881(csa_tree_add_7_27_groupi_n_2062 ,csa_tree_add_7_27_groupi_n_2024 ,csa_tree_add_7_27_groupi_n_1934);
  and csa_tree_add_7_27_groupi_g5127__5115(csa_tree_add_7_27_groupi_n_2061 ,csa_tree_add_7_27_groupi_n_2025 ,csa_tree_add_7_27_groupi_n_1937);
  or csa_tree_add_7_27_groupi_g5128__7482(csa_tree_add_7_27_groupi_n_2060 ,csa_tree_add_7_27_groupi_n_1978 ,csa_tree_add_7_27_groupi_n_2019);
  or csa_tree_add_7_27_groupi_g5129__4733(csa_tree_add_7_27_groupi_n_2059 ,csa_tree_add_7_27_groupi_n_995 ,csa_tree_add_7_27_groupi_n_2031);
  or csa_tree_add_7_27_groupi_g5130__6161(csa_tree_add_7_27_groupi_n_2058 ,csa_tree_add_7_27_groupi_n_1244 ,csa_tree_add_7_27_groupi_n_2034);
  or csa_tree_add_7_27_groupi_g5131__9315(csa_tree_add_7_27_groupi_n_2069 ,csa_tree_add_7_27_groupi_n_2003 ,csa_tree_add_7_27_groupi_n_2038);
  or csa_tree_add_7_27_groupi_g5132__9945(csa_tree_add_7_27_groupi_n_2068 ,csa_tree_add_7_27_groupi_n_1998 ,csa_tree_add_7_27_groupi_n_2037);
  not csa_tree_add_7_27_groupi_g5133(csa_tree_add_7_27_groupi_n_2056 ,csa_tree_add_7_27_groupi_n_2057);
  not csa_tree_add_7_27_groupi_g5134(csa_tree_add_7_27_groupi_n_2054 ,csa_tree_add_7_27_groupi_n_2055);
  nor csa_tree_add_7_27_groupi_g5135__2883(csa_tree_add_7_27_groupi_n_2052 ,csa_tree_add_7_27_groupi_n_311 ,csa_tree_add_7_27_groupi_n_540);
  nor csa_tree_add_7_27_groupi_g5136__2346(csa_tree_add_7_27_groupi_n_2051 ,csa_tree_add_7_27_groupi_n_329 ,csa_tree_add_7_27_groupi_n_543);
  and csa_tree_add_7_27_groupi_g5137__1666(csa_tree_add_7_27_groupi_n_2050 ,csa_tree_add_7_27_groupi_n_2023 ,csa_tree_add_7_27_groupi_n_1928);
  and csa_tree_add_7_27_groupi_g5138__7410(csa_tree_add_7_27_groupi_n_2049 ,csa_tree_add_7_27_groupi_n_2021 ,csa_tree_add_7_27_groupi_n_1923);
  nor csa_tree_add_7_27_groupi_g5139__6417(csa_tree_add_7_27_groupi_n_2048 ,csa_tree_add_7_27_groupi_n_299 ,csa_tree_add_7_27_groupi_n_2040);
  or csa_tree_add_7_27_groupi_g5140__5477(csa_tree_add_7_27_groupi_n_2047 ,csa_tree_add_7_27_groupi_n_1051 ,csa_tree_add_7_27_groupi_n_2039);
  and csa_tree_add_7_27_groupi_g5141__2398(csa_tree_add_7_27_groupi_n_2046 ,csa_tree_add_7_27_groupi_n_1428 ,csa_tree_add_7_27_groupi_n_2022);
  nor csa_tree_add_7_27_groupi_g5142__5107(csa_tree_add_7_27_groupi_n_2045 ,csa_tree_add_7_27_groupi_n_356 ,csa_tree_add_7_27_groupi_n_541);
  nor csa_tree_add_7_27_groupi_g5143__6260(csa_tree_add_7_27_groupi_n_2044 ,csa_tree_add_7_27_groupi_n_278 ,csa_tree_add_7_27_groupi_n_543);
  or csa_tree_add_7_27_groupi_g5144__4319(csa_tree_add_7_27_groupi_n_2057 ,csa_tree_add_7_27_groupi_n_1986 ,csa_tree_add_7_27_groupi_n_2032);
  or csa_tree_add_7_27_groupi_g5145__8428(csa_tree_add_7_27_groupi_n_2055 ,csa_tree_add_7_27_groupi_n_1992 ,csa_tree_add_7_27_groupi_n_2033);
  or csa_tree_add_7_27_groupi_g5146__5526(csa_tree_add_7_27_groupi_n_2053 ,csa_tree_add_7_27_groupi_n_2041 ,csa_tree_add_7_27_groupi_n_2035);
  not csa_tree_add_7_27_groupi_g5147(csa_tree_add_7_27_groupi_n_2041 ,csa_tree_add_7_27_groupi_n_541);
  nor csa_tree_add_7_27_groupi_g5148__6783(csa_tree_add_7_27_groupi_n_2039 ,csa_tree_add_7_27_groupi_n_310 ,csa_tree_add_7_27_groupi_n_521);
  and csa_tree_add_7_27_groupi_g5149__3680(csa_tree_add_7_27_groupi_n_2038 ,csa_tree_add_7_27_groupi_n_2006 ,csa_tree_add_7_27_groupi_n_1997);
  and csa_tree_add_7_27_groupi_g5150__1617(csa_tree_add_7_27_groupi_n_2037 ,csa_tree_add_7_27_groupi_n_1980 ,csa_tree_add_7_27_groupi_n_1996);
  nor csa_tree_add_7_27_groupi_g5151__2802(csa_tree_add_7_27_groupi_n_2036 ,csa_tree_add_7_27_groupi_n_298 ,csa_tree_add_7_27_groupi_n_1994);
  nor csa_tree_add_7_27_groupi_g5152__1705(csa_tree_add_7_27_groupi_n_2035 ,in1[15] ,csa_tree_add_7_27_groupi_n_2008);
  nor csa_tree_add_7_27_groupi_g5153__5122(csa_tree_add_7_27_groupi_n_2034 ,csa_tree_add_7_27_groupi_n_355 ,csa_tree_add_7_27_groupi_n_521);
  and csa_tree_add_7_27_groupi_g5154__8246(csa_tree_add_7_27_groupi_n_2033 ,csa_tree_add_7_27_groupi_n_1979 ,csa_tree_add_7_27_groupi_n_1991);
  and csa_tree_add_7_27_groupi_g5155__7098(csa_tree_add_7_27_groupi_n_2032 ,csa_tree_add_7_27_groupi_n_1981 ,csa_tree_add_7_27_groupi_n_1985);
  nor csa_tree_add_7_27_groupi_g5156__6131(csa_tree_add_7_27_groupi_n_2031 ,csa_tree_add_7_27_groupi_n_277 ,csa_tree_add_7_27_groupi_n_1994);
  nor csa_tree_add_7_27_groupi_g5157__1881(csa_tree_add_7_27_groupi_n_2030 ,csa_tree_add_7_27_groupi_n_1269 ,csa_tree_add_7_27_groupi_n_1993);
  nor csa_tree_add_7_27_groupi_g5158__5115(csa_tree_add_7_27_groupi_n_2029 ,csa_tree_add_7_27_groupi_n_1360 ,csa_tree_add_7_27_groupi_n_2001);
  nor csa_tree_add_7_27_groupi_g5159__7482(csa_tree_add_7_27_groupi_n_2028 ,csa_tree_add_7_27_groupi_n_1350 ,csa_tree_add_7_27_groupi_n_2000);
  nor csa_tree_add_7_27_groupi_g5160__4733(csa_tree_add_7_27_groupi_n_2027 ,csa_tree_add_7_27_groupi_n_1146 ,csa_tree_add_7_27_groupi_n_1982);
  nor csa_tree_add_7_27_groupi_g5161__6161(csa_tree_add_7_27_groupi_n_2026 ,csa_tree_add_7_27_groupi_n_1320 ,csa_tree_add_7_27_groupi_n_2004);
  or csa_tree_add_7_27_groupi_g5162__9315(csa_tree_add_7_27_groupi_n_2043 ,csa_tree_add_7_27_groupi_n_1841 ,csa_tree_add_7_27_groupi_n_1995);
  or csa_tree_add_7_27_groupi_g5163__9945(csa_tree_add_7_27_groupi_n_2042 ,csa_tree_add_7_27_groupi_n_1844 ,csa_tree_add_7_27_groupi_n_2005);
  or csa_tree_add_7_27_groupi_g5164__2883(csa_tree_add_7_27_groupi_n_2040 ,csa_tree_add_7_27_groupi_n_10 ,csa_tree_add_7_27_groupi_n_2007);
  nor csa_tree_add_7_27_groupi_g5165__2346(csa_tree_add_7_27_groupi_n_2018 ,csa_tree_add_7_27_groupi_n_328 ,csa_tree_add_7_27_groupi_n_520);
  xnor csa_tree_add_7_27_groupi_g5166__1666(n_12 ,csa_tree_add_7_27_groupi_n_1944 ,csa_tree_add_7_27_groupi_n_1947);
  xnor csa_tree_add_7_27_groupi_g5167__7410(csa_tree_add_7_27_groupi_n_2016 ,csa_tree_add_7_27_groupi_n_1955 ,csa_tree_add_7_27_groupi_n_1894);
  xnor csa_tree_add_7_27_groupi_g5168__6417(csa_tree_add_7_27_groupi_n_2015 ,csa_tree_add_7_27_groupi_n_1916 ,csa_tree_add_7_27_groupi_n_1953);
  xnor csa_tree_add_7_27_groupi_g5169__5477(csa_tree_add_7_27_groupi_n_2014 ,csa_tree_add_7_27_groupi_n_1913 ,csa_tree_add_7_27_groupi_n_1956);
  xnor csa_tree_add_7_27_groupi_g5170__2398(csa_tree_add_7_27_groupi_n_2013 ,csa_tree_add_7_27_groupi_n_1961 ,csa_tree_add_7_27_groupi_n_1854);
  xnor csa_tree_add_7_27_groupi_g5171__5107(csa_tree_add_7_27_groupi_n_2012 ,csa_tree_add_7_27_groupi_n_1915 ,csa_tree_add_7_27_groupi_n_1963);
  xnor csa_tree_add_7_27_groupi_g5172__6260(csa_tree_add_7_27_groupi_n_2011 ,csa_tree_add_7_27_groupi_n_1918 ,csa_tree_add_7_27_groupi_n_1960);
  xnor csa_tree_add_7_27_groupi_g5173__4319(csa_tree_add_7_27_groupi_n_2010 ,csa_tree_add_7_27_groupi_n_1920 ,csa_tree_add_7_27_groupi_n_1958);
  xnor csa_tree_add_7_27_groupi_g5174__8428(csa_tree_add_7_27_groupi_n_2009 ,csa_tree_add_7_27_groupi_n_1412 ,csa_tree_add_7_27_groupi_n_1952);
  xnor csa_tree_add_7_27_groupi_g5175__5526(csa_tree_add_7_27_groupi_n_2025 ,csa_tree_add_7_27_groupi_n_1970 ,in2[5]);
  xnor csa_tree_add_7_27_groupi_g5176__6783(csa_tree_add_7_27_groupi_n_2024 ,csa_tree_add_7_27_groupi_n_1966 ,in2[2]);
  xnor csa_tree_add_7_27_groupi_g5177__3680(csa_tree_add_7_27_groupi_n_2023 ,csa_tree_add_7_27_groupi_n_1967 ,in2[11]);
  xnor csa_tree_add_7_27_groupi_g5178__1617(csa_tree_add_7_27_groupi_n_2022 ,csa_tree_add_7_27_groupi_n_1968 ,in2[14]);
  xnor csa_tree_add_7_27_groupi_g5179__2802(csa_tree_add_7_27_groupi_n_2021 ,csa_tree_add_7_27_groupi_n_1969 ,in2[8]);
  xnor csa_tree_add_7_27_groupi_g5180__1705(csa_tree_add_7_27_groupi_n_2020 ,csa_tree_add_7_27_groupi_n_1965 ,csa_tree_add_7_27_groupi_n_1848);
  xnor csa_tree_add_7_27_groupi_g5181__5122(csa_tree_add_7_27_groupi_n_2019 ,csa_tree_add_7_27_groupi_n_1964 ,csa_tree_add_7_27_groupi_n_1847);
  not csa_tree_add_7_27_groupi_g5182(csa_tree_add_7_27_groupi_n_2008 ,csa_tree_add_7_27_groupi_n_2007);
  and csa_tree_add_7_27_groupi_g5183__8246(csa_tree_add_7_27_groupi_n_2005 ,csa_tree_add_7_27_groupi_n_1965 ,csa_tree_add_7_27_groupi_n_1843);
  or csa_tree_add_7_27_groupi_g5184__7098(csa_tree_add_7_27_groupi_n_2004 ,csa_tree_add_7_27_groupi_n_1085 ,csa_tree_add_7_27_groupi_n_1974);
  and csa_tree_add_7_27_groupi_g5185__6131(csa_tree_add_7_27_groupi_n_2003 ,csa_tree_add_7_27_groupi_n_1913 ,csa_tree_add_7_27_groupi_n_1956);
  or csa_tree_add_7_27_groupi_g5186__1881(csa_tree_add_7_27_groupi_n_2002 ,csa_tree_add_7_27_groupi_n_1916 ,csa_tree_add_7_27_groupi_n_1953);
  or csa_tree_add_7_27_groupi_g5187__5115(csa_tree_add_7_27_groupi_n_2001 ,csa_tree_add_7_27_groupi_n_1112 ,csa_tree_add_7_27_groupi_n_1976);
  or csa_tree_add_7_27_groupi_g5188__7482(csa_tree_add_7_27_groupi_n_2000 ,csa_tree_add_7_27_groupi_n_1152 ,csa_tree_add_7_27_groupi_n_1950);
  and csa_tree_add_7_27_groupi_g5189__4733(csa_tree_add_7_27_groupi_n_1999 ,csa_tree_add_7_27_groupi_n_1916 ,csa_tree_add_7_27_groupi_n_1953);
  and csa_tree_add_7_27_groupi_g5190__6161(csa_tree_add_7_27_groupi_n_1998 ,csa_tree_add_7_27_groupi_n_1961 ,csa_tree_add_7_27_groupi_n_1854);
  or csa_tree_add_7_27_groupi_g5191__9315(csa_tree_add_7_27_groupi_n_1997 ,csa_tree_add_7_27_groupi_n_1913 ,csa_tree_add_7_27_groupi_n_1956);
  or csa_tree_add_7_27_groupi_g5192__9945(csa_tree_add_7_27_groupi_n_1996 ,csa_tree_add_7_27_groupi_n_1961 ,csa_tree_add_7_27_groupi_n_1854);
  and csa_tree_add_7_27_groupi_g5193__2883(csa_tree_add_7_27_groupi_n_1995 ,csa_tree_add_7_27_groupi_n_1964 ,csa_tree_add_7_27_groupi_n_1842);
  and csa_tree_add_7_27_groupi_g5194__2346(csa_tree_add_7_27_groupi_n_2007 ,csa_tree_add_7_27_groupi_n_773 ,csa_tree_add_7_27_groupi_n_1975);
  or csa_tree_add_7_27_groupi_g5195__1666(csa_tree_add_7_27_groupi_n_2006 ,csa_tree_add_7_27_groupi_n_1971 ,csa_tree_add_7_27_groupi_n_1930);
  or csa_tree_add_7_27_groupi_g5196__7410(csa_tree_add_7_27_groupi_n_1993 ,csa_tree_add_7_27_groupi_n_1216 ,csa_tree_add_7_27_groupi_n_1973);
  nor csa_tree_add_7_27_groupi_g5197__6417(csa_tree_add_7_27_groupi_n_1992 ,csa_tree_add_7_27_groupi_n_1412 ,csa_tree_add_7_27_groupi_n_1951);
  or csa_tree_add_7_27_groupi_g5198__5477(csa_tree_add_7_27_groupi_n_1991 ,csa_tree_add_7_27_groupi_n_1411 ,csa_tree_add_7_27_groupi_n_1952);
  nor csa_tree_add_7_27_groupi_g5199__2398(csa_tree_add_7_27_groupi_n_1990 ,csa_tree_add_7_27_groupi_n_1919 ,csa_tree_add_7_27_groupi_n_1958);
  or csa_tree_add_7_27_groupi_g5200__5107(csa_tree_add_7_27_groupi_n_1989 ,csa_tree_add_7_27_groupi_n_1920 ,csa_tree_add_7_27_groupi_n_1957);
  nor csa_tree_add_7_27_groupi_g5201__6260(csa_tree_add_7_27_groupi_n_1988 ,csa_tree_add_7_27_groupi_n_1914 ,csa_tree_add_7_27_groupi_n_1963);
  or csa_tree_add_7_27_groupi_g5202__4319(csa_tree_add_7_27_groupi_n_1987 ,csa_tree_add_7_27_groupi_n_1915 ,csa_tree_add_7_27_groupi_n_1962);
  nor csa_tree_add_7_27_groupi_g5203__8428(csa_tree_add_7_27_groupi_n_1986 ,csa_tree_add_7_27_groupi_n_1954 ,csa_tree_add_7_27_groupi_n_1894);
  or csa_tree_add_7_27_groupi_g5204__5526(csa_tree_add_7_27_groupi_n_1985 ,csa_tree_add_7_27_groupi_n_1955 ,csa_tree_add_7_27_groupi_n_1893);
  nor csa_tree_add_7_27_groupi_g5205__6783(csa_tree_add_7_27_groupi_n_1984 ,csa_tree_add_7_27_groupi_n_1917 ,csa_tree_add_7_27_groupi_n_1960);
  or csa_tree_add_7_27_groupi_g5206__3680(csa_tree_add_7_27_groupi_n_1983 ,csa_tree_add_7_27_groupi_n_1918 ,csa_tree_add_7_27_groupi_n_1959);
  or csa_tree_add_7_27_groupi_g5207__1617(csa_tree_add_7_27_groupi_n_1982 ,csa_tree_add_7_27_groupi_n_1006 ,csa_tree_add_7_27_groupi_n_1972);
  xnor csa_tree_add_7_27_groupi_g5208__2802(csa_tree_add_7_27_groupi_n_1994 ,csa_tree_add_7_27_groupi_n_1943 ,csa_tree_add_7_27_groupi_n_836);
  nor csa_tree_add_7_27_groupi_g5209__1705(csa_tree_add_7_27_groupi_n_1976 ,csa_tree_add_7_27_groupi_n_277 ,csa_tree_add_7_27_groupi_n_518);
  or csa_tree_add_7_27_groupi_g5210__5122(csa_tree_add_7_27_groupi_n_1975 ,csa_tree_add_7_27_groupi_n_782 ,csa_tree_add_7_27_groupi_n_1943);
  nor csa_tree_add_7_27_groupi_g5211__8246(csa_tree_add_7_27_groupi_n_1974 ,csa_tree_add_7_27_groupi_n_298 ,csa_tree_add_7_27_groupi_n_1932);
  nor csa_tree_add_7_27_groupi_g5212__7098(csa_tree_add_7_27_groupi_n_1973 ,csa_tree_add_7_27_groupi_n_355 ,csa_tree_add_7_27_groupi_n_518);
  nor csa_tree_add_7_27_groupi_g5213__6131(csa_tree_add_7_27_groupi_n_1972 ,csa_tree_add_7_27_groupi_n_310 ,csa_tree_add_7_27_groupi_n_1932);
  and csa_tree_add_7_27_groupi_g5214__1881(csa_tree_add_7_27_groupi_n_1971 ,csa_tree_add_7_27_groupi_n_1936 ,csa_tree_add_7_27_groupi_n_1944);
  nor csa_tree_add_7_27_groupi_g5215__5115(csa_tree_add_7_27_groupi_n_1970 ,csa_tree_add_7_27_groupi_n_1352 ,csa_tree_add_7_27_groupi_n_1938);
  nor csa_tree_add_7_27_groupi_g5216__7482(csa_tree_add_7_27_groupi_n_1969 ,csa_tree_add_7_27_groupi_n_1323 ,csa_tree_add_7_27_groupi_n_1925);
  nor csa_tree_add_7_27_groupi_g5217__4733(csa_tree_add_7_27_groupi_n_1968 ,csa_tree_add_7_27_groupi_n_1363 ,csa_tree_add_7_27_groupi_n_1941);
  nor csa_tree_add_7_27_groupi_g5218__6161(csa_tree_add_7_27_groupi_n_1967 ,csa_tree_add_7_27_groupi_n_1356 ,csa_tree_add_7_27_groupi_n_1929);
  nor csa_tree_add_7_27_groupi_g5219__9315(csa_tree_add_7_27_groupi_n_1966 ,csa_tree_add_7_27_groupi_n_1127 ,csa_tree_add_7_27_groupi_n_1922);
  or csa_tree_add_7_27_groupi_g5220__9945(csa_tree_add_7_27_groupi_n_1981 ,csa_tree_add_7_27_groupi_n_1828 ,csa_tree_add_7_27_groupi_n_1939);
  or csa_tree_add_7_27_groupi_g5221__2883(csa_tree_add_7_27_groupi_n_1980 ,csa_tree_add_7_27_groupi_n_1781 ,csa_tree_add_7_27_groupi_n_1931);
  or csa_tree_add_7_27_groupi_g5222__2346(csa_tree_add_7_27_groupi_n_1979 ,csa_tree_add_7_27_groupi_n_1179 ,csa_tree_add_7_27_groupi_n_1927);
  or csa_tree_add_7_27_groupi_g5223__1666(csa_tree_add_7_27_groupi_n_1978 ,csa_tree_add_7_27_groupi_n_1795 ,csa_tree_add_7_27_groupi_n_1933);
  or csa_tree_add_7_27_groupi_g5224__7410(csa_tree_add_7_27_groupi_n_1977 ,csa_tree_add_7_27_groupi_n_1791 ,csa_tree_add_7_27_groupi_n_1942);
  not csa_tree_add_7_27_groupi_g5225(csa_tree_add_7_27_groupi_n_1963 ,csa_tree_add_7_27_groupi_n_1962);
  not csa_tree_add_7_27_groupi_g5226(csa_tree_add_7_27_groupi_n_1959 ,csa_tree_add_7_27_groupi_n_1960);
  not csa_tree_add_7_27_groupi_g5227(csa_tree_add_7_27_groupi_n_1957 ,csa_tree_add_7_27_groupi_n_1958);
  not csa_tree_add_7_27_groupi_g5228(csa_tree_add_7_27_groupi_n_1954 ,csa_tree_add_7_27_groupi_n_1955);
  not csa_tree_add_7_27_groupi_g5229(csa_tree_add_7_27_groupi_n_1951 ,csa_tree_add_7_27_groupi_n_1952);
  nor csa_tree_add_7_27_groupi_g5230__6417(csa_tree_add_7_27_groupi_n_1950 ,csa_tree_add_7_27_groupi_n_328 ,csa_tree_add_7_27_groupi_n_517);
  xnor csa_tree_add_7_27_groupi_g5231__5477(csa_tree_add_7_27_groupi_n_1949 ,csa_tree_add_7_27_groupi_n_1798 ,csa_tree_add_7_27_groupi_n_1897);
  xnor csa_tree_add_7_27_groupi_g5232__2398(csa_tree_add_7_27_groupi_n_1948 ,csa_tree_add_7_27_groupi_n_1797 ,csa_tree_add_7_27_groupi_n_1898);
  xnor csa_tree_add_7_27_groupi_g5233__5107(csa_tree_add_7_27_groupi_n_1947 ,csa_tree_add_7_27_groupi_n_1796 ,csa_tree_add_7_27_groupi_n_1896);
  xnor csa_tree_add_7_27_groupi_g5234__6260(csa_tree_add_7_27_groupi_n_1946 ,csa_tree_add_7_27_groupi_n_1895 ,csa_tree_add_7_27_groupi_n_1871);
  xnor csa_tree_add_7_27_groupi_g5235__4319(csa_tree_add_7_27_groupi_n_1945 ,csa_tree_add_7_27_groupi_n_1892 ,csa_tree_add_7_27_groupi_n_1880);
  xnor csa_tree_add_7_27_groupi_g5236__8428(csa_tree_add_7_27_groupi_n_1965 ,csa_tree_add_7_27_groupi_n_1907 ,in2[5]);
  xnor csa_tree_add_7_27_groupi_g5237__5526(csa_tree_add_7_27_groupi_n_1964 ,csa_tree_add_7_27_groupi_n_1906 ,in2[2]);
  xnor csa_tree_add_7_27_groupi_g5238__6783(csa_tree_add_7_27_groupi_n_1962 ,csa_tree_add_7_27_groupi_n_1902 ,csa_tree_add_7_27_groupi_n_1801);
  xnor csa_tree_add_7_27_groupi_g5239__3680(csa_tree_add_7_27_groupi_n_1961 ,csa_tree_add_7_27_groupi_n_1908 ,in2[8]);
  xnor csa_tree_add_7_27_groupi_g5240__1617(csa_tree_add_7_27_groupi_n_1960 ,csa_tree_add_7_27_groupi_n_1901 ,csa_tree_add_7_27_groupi_n_1850);
  xnor csa_tree_add_7_27_groupi_g5241__2802(csa_tree_add_7_27_groupi_n_1958 ,csa_tree_add_7_27_groupi_n_1899 ,csa_tree_add_7_27_groupi_n_1306);
  xnor csa_tree_add_7_27_groupi_g5242__1705(csa_tree_add_7_27_groupi_n_1956 ,csa_tree_add_7_27_groupi_n_1903 ,csa_tree_add_7_27_groupi_n_1805);
  xnor csa_tree_add_7_27_groupi_g5243__5122(csa_tree_add_7_27_groupi_n_1955 ,csa_tree_add_7_27_groupi_n_1904 ,in2[11]);
  xnor csa_tree_add_7_27_groupi_g5244__8246(csa_tree_add_7_27_groupi_n_1953 ,csa_tree_add_7_27_groupi_n_1900 ,csa_tree_add_7_27_groupi_n_1804);
  xnor csa_tree_add_7_27_groupi_g5245__7098(csa_tree_add_7_27_groupi_n_1952 ,csa_tree_add_7_27_groupi_n_1905 ,in2[14]);
  and csa_tree_add_7_27_groupi_g5246__6131(csa_tree_add_7_27_groupi_n_1942 ,csa_tree_add_7_27_groupi_n_1900 ,csa_tree_add_7_27_groupi_n_1794);
  or csa_tree_add_7_27_groupi_g5247__1881(csa_tree_add_7_27_groupi_n_1941 ,csa_tree_add_7_27_groupi_n_1113 ,csa_tree_add_7_27_groupi_n_1889);
  and csa_tree_add_7_27_groupi_g5248__5115(csa_tree_add_7_27_groupi_n_1940 ,csa_tree_add_7_27_groupi_n_1797 ,csa_tree_add_7_27_groupi_n_1898);
  and csa_tree_add_7_27_groupi_g5249__7482(csa_tree_add_7_27_groupi_n_1939 ,csa_tree_add_7_27_groupi_n_1901 ,csa_tree_add_7_27_groupi_n_1827);
  or csa_tree_add_7_27_groupi_g5250__4733(csa_tree_add_7_27_groupi_n_1938 ,csa_tree_add_7_27_groupi_n_1101 ,csa_tree_add_7_27_groupi_n_1912);
  or csa_tree_add_7_27_groupi_g5251__6161(csa_tree_add_7_27_groupi_n_1937 ,csa_tree_add_7_27_groupi_n_1797 ,csa_tree_add_7_27_groupi_n_1898);
  or csa_tree_add_7_27_groupi_g5252__9315(csa_tree_add_7_27_groupi_n_1936 ,csa_tree_add_7_27_groupi_n_1796 ,csa_tree_add_7_27_groupi_n_1896);
  and csa_tree_add_7_27_groupi_g5253__9945(csa_tree_add_7_27_groupi_n_1935 ,csa_tree_add_7_27_groupi_n_1798 ,csa_tree_add_7_27_groupi_n_1897);
  or csa_tree_add_7_27_groupi_g5254__2883(csa_tree_add_7_27_groupi_n_1934 ,csa_tree_add_7_27_groupi_n_1798 ,csa_tree_add_7_27_groupi_n_1897);
  and csa_tree_add_7_27_groupi_g5255__2346(csa_tree_add_7_27_groupi_n_1933 ,csa_tree_add_7_27_groupi_n_1903 ,csa_tree_add_7_27_groupi_n_1790);
  or csa_tree_add_7_27_groupi_g5256__1666(csa_tree_add_7_27_groupi_n_1944 ,csa_tree_add_7_27_groupi_n_1839 ,csa_tree_add_7_27_groupi_n_1909);
  and csa_tree_add_7_27_groupi_g5257__7410(csa_tree_add_7_27_groupi_n_1943 ,csa_tree_add_7_27_groupi_n_792 ,csa_tree_add_7_27_groupi_n_1911);
  and csa_tree_add_7_27_groupi_g5258__6417(csa_tree_add_7_27_groupi_n_1931 ,csa_tree_add_7_27_groupi_n_1902 ,csa_tree_add_7_27_groupi_n_1780);
  and csa_tree_add_7_27_groupi_g5259__5477(csa_tree_add_7_27_groupi_n_1930 ,csa_tree_add_7_27_groupi_n_1796 ,csa_tree_add_7_27_groupi_n_1896);
  or csa_tree_add_7_27_groupi_g5260__2398(csa_tree_add_7_27_groupi_n_1929 ,csa_tree_add_7_27_groupi_n_987 ,csa_tree_add_7_27_groupi_n_1888);
  or csa_tree_add_7_27_groupi_g5261__5107(csa_tree_add_7_27_groupi_n_1928 ,csa_tree_add_7_27_groupi_n_1891 ,csa_tree_add_7_27_groupi_n_1880);
  and csa_tree_add_7_27_groupi_g5262__6260(csa_tree_add_7_27_groupi_n_1927 ,csa_tree_add_7_27_groupi_n_1180 ,csa_tree_add_7_27_groupi_n_1899);
  nor csa_tree_add_7_27_groupi_g5263__4319(csa_tree_add_7_27_groupi_n_1926 ,csa_tree_add_7_27_groupi_n_1892 ,csa_tree_add_7_27_groupi_n_1879);
  or csa_tree_add_7_27_groupi_g5264__8428(csa_tree_add_7_27_groupi_n_1925 ,csa_tree_add_7_27_groupi_n_1133 ,csa_tree_add_7_27_groupi_n_1890);
  and csa_tree_add_7_27_groupi_g5265__5526(csa_tree_add_7_27_groupi_n_1924 ,csa_tree_add_7_27_groupi_n_1895 ,csa_tree_add_7_27_groupi_n_1871);
  or csa_tree_add_7_27_groupi_g5266__6783(csa_tree_add_7_27_groupi_n_1923 ,csa_tree_add_7_27_groupi_n_1895 ,csa_tree_add_7_27_groupi_n_1871);
  or csa_tree_add_7_27_groupi_g5267__3680(csa_tree_add_7_27_groupi_n_1922 ,csa_tree_add_7_27_groupi_n_991 ,csa_tree_add_7_27_groupi_n_1910);
  xnor csa_tree_add_7_27_groupi_g5268__1617(n_11 ,csa_tree_add_7_27_groupi_n_1886 ,csa_tree_add_7_27_groupi_n_1851);
  xnor csa_tree_add_7_27_groupi_g5269__2802(csa_tree_add_7_27_groupi_n_1932 ,csa_tree_add_7_27_groupi_n_1887 ,csa_tree_add_7_27_groupi_n_840);
  not csa_tree_add_7_27_groupi_g5270(csa_tree_add_7_27_groupi_n_1919 ,csa_tree_add_7_27_groupi_n_1920);
  not csa_tree_add_7_27_groupi_g5271(csa_tree_add_7_27_groupi_n_1917 ,csa_tree_add_7_27_groupi_n_1918);
  not csa_tree_add_7_27_groupi_g5272(csa_tree_add_7_27_groupi_n_1914 ,csa_tree_add_7_27_groupi_n_1915);
  nor csa_tree_add_7_27_groupi_g5273__1705(csa_tree_add_7_27_groupi_n_1912 ,csa_tree_add_7_27_groupi_n_464 ,csa_tree_add_7_27_groupi_n_532);
  or csa_tree_add_7_27_groupi_g5274__5122(csa_tree_add_7_27_groupi_n_1911 ,csa_tree_add_7_27_groupi_n_793 ,csa_tree_add_7_27_groupi_n_1887);
  nor csa_tree_add_7_27_groupi_g5275__8246(csa_tree_add_7_27_groupi_n_1910 ,csa_tree_add_7_27_groupi_n_461 ,csa_tree_add_7_27_groupi_n_1878);
  and csa_tree_add_7_27_groupi_g5276__7098(csa_tree_add_7_27_groupi_n_1909 ,csa_tree_add_7_27_groupi_n_1838 ,csa_tree_add_7_27_groupi_n_1886);
  nor csa_tree_add_7_27_groupi_g5277__6131(csa_tree_add_7_27_groupi_n_1908 ,csa_tree_add_7_27_groupi_n_1294 ,csa_tree_add_7_27_groupi_n_1876);
  nor csa_tree_add_7_27_groupi_g5278__1881(csa_tree_add_7_27_groupi_n_1907 ,csa_tree_add_7_27_groupi_n_1346 ,csa_tree_add_7_27_groupi_n_1884);
  nor csa_tree_add_7_27_groupi_g5279__5115(csa_tree_add_7_27_groupi_n_1906 ,csa_tree_add_7_27_groupi_n_1150 ,csa_tree_add_7_27_groupi_n_1872);
  nor csa_tree_add_7_27_groupi_g5280__7482(csa_tree_add_7_27_groupi_n_1905 ,csa_tree_add_7_27_groupi_n_1348 ,csa_tree_add_7_27_groupi_n_1883);
  nor csa_tree_add_7_27_groupi_g5281__4733(csa_tree_add_7_27_groupi_n_1904 ,csa_tree_add_7_27_groupi_n_1286 ,csa_tree_add_7_27_groupi_n_1873);
  or csa_tree_add_7_27_groupi_g5282__6161(csa_tree_add_7_27_groupi_n_1920 ,csa_tree_add_7_27_groupi_n_1429 ,csa_tree_add_7_27_groupi_n_1875);
  or csa_tree_add_7_27_groupi_g5283__9315(csa_tree_add_7_27_groupi_n_1918 ,csa_tree_add_7_27_groupi_n_1778 ,csa_tree_add_7_27_groupi_n_1877);
  or csa_tree_add_7_27_groupi_g5284__9945(csa_tree_add_7_27_groupi_n_1916 ,csa_tree_add_7_27_groupi_n_1733 ,csa_tree_add_7_27_groupi_n_1885);
  or csa_tree_add_7_27_groupi_g5285__2883(csa_tree_add_7_27_groupi_n_1915 ,csa_tree_add_7_27_groupi_n_1739 ,csa_tree_add_7_27_groupi_n_1881);
  or csa_tree_add_7_27_groupi_g5286__2346(csa_tree_add_7_27_groupi_n_1913 ,csa_tree_add_7_27_groupi_n_1735 ,csa_tree_add_7_27_groupi_n_1882);
  not csa_tree_add_7_27_groupi_g5287(csa_tree_add_7_27_groupi_n_1893 ,csa_tree_add_7_27_groupi_n_1894);
  not csa_tree_add_7_27_groupi_g5288(csa_tree_add_7_27_groupi_n_1891 ,csa_tree_add_7_27_groupi_n_1892);
  nor csa_tree_add_7_27_groupi_g5289__1666(csa_tree_add_7_27_groupi_n_1890 ,csa_tree_add_7_27_groupi_n_458 ,csa_tree_add_7_27_groupi_n_532);
  nor csa_tree_add_7_27_groupi_g5290__7410(csa_tree_add_7_27_groupi_n_1889 ,csa_tree_add_7_27_groupi_n_467 ,csa_tree_add_7_27_groupi_n_1878);
  nor csa_tree_add_7_27_groupi_g5291__6417(csa_tree_add_7_27_groupi_n_1888 ,csa_tree_add_7_27_groupi_n_455 ,csa_tree_add_7_27_groupi_n_531);
  xnor csa_tree_add_7_27_groupi_g5292__5477(csa_tree_add_7_27_groupi_n_1903 ,csa_tree_add_7_27_groupi_n_1863 ,in2[2]);
  xnor csa_tree_add_7_27_groupi_g5293__2398(csa_tree_add_7_27_groupi_n_1902 ,csa_tree_add_7_27_groupi_n_1864 ,in2[8]);
  xnor csa_tree_add_7_27_groupi_g5294__5107(csa_tree_add_7_27_groupi_n_1901 ,csa_tree_add_7_27_groupi_n_1862 ,in2[11]);
  xnor csa_tree_add_7_27_groupi_g5295__6260(csa_tree_add_7_27_groupi_n_1900 ,csa_tree_add_7_27_groupi_n_1860 ,in2[5]);
  xnor csa_tree_add_7_27_groupi_g5296__4319(csa_tree_add_7_27_groupi_n_1899 ,csa_tree_add_7_27_groupi_n_1861 ,in2[14]);
  xnor csa_tree_add_7_27_groupi_g5297__8428(csa_tree_add_7_27_groupi_n_1898 ,csa_tree_add_7_27_groupi_n_1857 ,csa_tree_add_7_27_groupi_n_1746);
  xnor csa_tree_add_7_27_groupi_g5298__5526(csa_tree_add_7_27_groupi_n_1897 ,csa_tree_add_7_27_groupi_n_1859 ,csa_tree_add_7_27_groupi_n_1747);
  xnor csa_tree_add_7_27_groupi_g5299__6783(csa_tree_add_7_27_groupi_n_1896 ,csa_tree_add_7_27_groupi_n_1856 ,csa_tree_add_7_27_groupi_n_1748);
  xnor csa_tree_add_7_27_groupi_g5300__3680(csa_tree_add_7_27_groupi_n_1895 ,csa_tree_add_7_27_groupi_n_1858 ,csa_tree_add_7_27_groupi_n_1802);
  xnor csa_tree_add_7_27_groupi_g5301__1617(csa_tree_add_7_27_groupi_n_1894 ,csa_tree_add_7_27_groupi_n_1826 ,csa_tree_add_7_27_groupi_n_1849);
  xnor csa_tree_add_7_27_groupi_g5302__2802(csa_tree_add_7_27_groupi_n_1892 ,csa_tree_add_7_27_groupi_n_1855 ,csa_tree_add_7_27_groupi_n_1433);
  and csa_tree_add_7_27_groupi_g5303__1705(csa_tree_add_7_27_groupi_n_1885 ,csa_tree_add_7_27_groupi_n_1859 ,csa_tree_add_7_27_groupi_n_1732);
  or csa_tree_add_7_27_groupi_g5304__5122(csa_tree_add_7_27_groupi_n_1884 ,csa_tree_add_7_27_groupi_n_1106 ,csa_tree_add_7_27_groupi_n_1868);
  or csa_tree_add_7_27_groupi_g5305__8246(csa_tree_add_7_27_groupi_n_1883 ,csa_tree_add_7_27_groupi_n_1111 ,csa_tree_add_7_27_groupi_n_1853);
  and csa_tree_add_7_27_groupi_g5306__7098(csa_tree_add_7_27_groupi_n_1882 ,csa_tree_add_7_27_groupi_n_1856 ,csa_tree_add_7_27_groupi_n_1737);
  and csa_tree_add_7_27_groupi_g5307__6131(csa_tree_add_7_27_groupi_n_1881 ,csa_tree_add_7_27_groupi_n_1857 ,csa_tree_add_7_27_groupi_n_1738);
  and csa_tree_add_7_27_groupi_g5308__1881(csa_tree_add_7_27_groupi_n_1887 ,csa_tree_add_7_27_groupi_n_796 ,csa_tree_add_7_27_groupi_n_1865);
  or csa_tree_add_7_27_groupi_g5309__5115(csa_tree_add_7_27_groupi_n_1886 ,csa_tree_add_7_27_groupi_n_1776 ,csa_tree_add_7_27_groupi_n_1870);
  not csa_tree_add_7_27_groupi_g5310(csa_tree_add_7_27_groupi_n_1879 ,csa_tree_add_7_27_groupi_n_1880);
  and csa_tree_add_7_27_groupi_g5311__7482(csa_tree_add_7_27_groupi_n_1877 ,csa_tree_add_7_27_groupi_n_1858 ,csa_tree_add_7_27_groupi_n_1777);
  or csa_tree_add_7_27_groupi_g5312__4733(csa_tree_add_7_27_groupi_n_1876 ,csa_tree_add_7_27_groupi_n_1226 ,csa_tree_add_7_27_groupi_n_1852);
  and csa_tree_add_7_27_groupi_g5313__6161(csa_tree_add_7_27_groupi_n_1875 ,csa_tree_add_7_27_groupi_n_1395 ,csa_tree_add_7_27_groupi_n_1855);
  xnor csa_tree_add_7_27_groupi_g5314__9315(n_10 ,csa_tree_add_7_27_groupi_n_1836 ,csa_tree_add_7_27_groupi_n_1803);
  or csa_tree_add_7_27_groupi_g5315__9945(csa_tree_add_7_27_groupi_n_1873 ,csa_tree_add_7_27_groupi_n_1234 ,csa_tree_add_7_27_groupi_n_1869);
  or csa_tree_add_7_27_groupi_g5316__2883(csa_tree_add_7_27_groupi_n_1872 ,csa_tree_add_7_27_groupi_n_1005 ,csa_tree_add_7_27_groupi_n_1867);
  or csa_tree_add_7_27_groupi_g5317__2346(csa_tree_add_7_27_groupi_n_1880 ,csa_tree_add_7_27_groupi_n_1831 ,csa_tree_add_7_27_groupi_n_1866);
  xnor csa_tree_add_7_27_groupi_g5318__1666(csa_tree_add_7_27_groupi_n_1878 ,csa_tree_add_7_27_groupi_n_1846 ,csa_tree_add_7_27_groupi_n_834);
  and csa_tree_add_7_27_groupi_g5319__7410(csa_tree_add_7_27_groupi_n_1870 ,csa_tree_add_7_27_groupi_n_1788 ,csa_tree_add_7_27_groupi_n_1836);
  nor csa_tree_add_7_27_groupi_g5320__6417(csa_tree_add_7_27_groupi_n_1869 ,csa_tree_add_7_27_groupi_n_343 ,csa_tree_add_7_27_groupi_n_535);
  nor csa_tree_add_7_27_groupi_g5321__5477(csa_tree_add_7_27_groupi_n_1868 ,csa_tree_add_7_27_groupi_n_268 ,csa_tree_add_7_27_groupi_n_1835);
  nor csa_tree_add_7_27_groupi_g5322__2398(csa_tree_add_7_27_groupi_n_1867 ,csa_tree_add_7_27_groupi_n_304 ,csa_tree_add_7_27_groupi_n_535);
  and csa_tree_add_7_27_groupi_g5323__5107(csa_tree_add_7_27_groupi_n_1866 ,csa_tree_add_7_27_groupi_n_1826 ,csa_tree_add_7_27_groupi_n_1832);
  or csa_tree_add_7_27_groupi_g5324__6260(csa_tree_add_7_27_groupi_n_1865 ,csa_tree_add_7_27_groupi_n_785 ,csa_tree_add_7_27_groupi_n_1846);
  nor csa_tree_add_7_27_groupi_g5325__4319(csa_tree_add_7_27_groupi_n_1864 ,csa_tree_add_7_27_groupi_n_1288 ,csa_tree_add_7_27_groupi_n_1833);
  nor csa_tree_add_7_27_groupi_g5326__8428(csa_tree_add_7_27_groupi_n_1863 ,csa_tree_add_7_27_groupi_n_1142 ,csa_tree_add_7_27_groupi_n_1829);
  nor csa_tree_add_7_27_groupi_g5327__5526(csa_tree_add_7_27_groupi_n_1862 ,csa_tree_add_7_27_groupi_n_1353 ,csa_tree_add_7_27_groupi_n_1837);
  nor csa_tree_add_7_27_groupi_g5328__6783(csa_tree_add_7_27_groupi_n_1861 ,csa_tree_add_7_27_groupi_n_1258 ,csa_tree_add_7_27_groupi_n_1834);
  nor csa_tree_add_7_27_groupi_g5329__3680(csa_tree_add_7_27_groupi_n_1860 ,csa_tree_add_7_27_groupi_n_1340 ,csa_tree_add_7_27_groupi_n_1840);
  or csa_tree_add_7_27_groupi_g5330__1617(csa_tree_add_7_27_groupi_n_1871 ,csa_tree_add_7_27_groupi_n_1766 ,csa_tree_add_7_27_groupi_n_1845);
  nor csa_tree_add_7_27_groupi_g5331__2802(csa_tree_add_7_27_groupi_n_1853 ,csa_tree_add_7_27_groupi_n_316 ,csa_tree_add_7_27_groupi_n_1835);
  nor csa_tree_add_7_27_groupi_g5332__1705(csa_tree_add_7_27_groupi_n_1852 ,csa_tree_add_7_27_groupi_n_283 ,csa_tree_add_7_27_groupi_n_534);
  xnor csa_tree_add_7_27_groupi_g5333__5122(csa_tree_add_7_27_groupi_n_1851 ,csa_tree_add_7_27_groupi_n_1813 ,csa_tree_add_7_27_groupi_n_1785);
  xnor csa_tree_add_7_27_groupi_g5334__8246(csa_tree_add_7_27_groupi_n_1850 ,csa_tree_add_7_27_groupi_n_1773 ,csa_tree_add_7_27_groupi_n_1808);
  xnor csa_tree_add_7_27_groupi_g5335__7098(csa_tree_add_7_27_groupi_n_1849 ,csa_tree_add_7_27_groupi_n_1408 ,csa_tree_add_7_27_groupi_n_1810);
  xnor csa_tree_add_7_27_groupi_g5336__6131(csa_tree_add_7_27_groupi_n_1848 ,csa_tree_add_7_27_groupi_n_1812 ,csa_tree_add_7_27_groupi_n_1786);
  xnor csa_tree_add_7_27_groupi_g5337__1881(csa_tree_add_7_27_groupi_n_1847 ,csa_tree_add_7_27_groupi_n_1811 ,csa_tree_add_7_27_groupi_n_1787);
  xnor csa_tree_add_7_27_groupi_g5338__5115(csa_tree_add_7_27_groupi_n_1859 ,csa_tree_add_7_27_groupi_n_1819 ,in2[5]);
  xnor csa_tree_add_7_27_groupi_g5339__7482(csa_tree_add_7_27_groupi_n_1858 ,csa_tree_add_7_27_groupi_n_1818 ,in2[11]);
  xnor csa_tree_add_7_27_groupi_g5340__4733(csa_tree_add_7_27_groupi_n_1857 ,csa_tree_add_7_27_groupi_n_1815 ,in2[8]);
  xnor csa_tree_add_7_27_groupi_g5341__6161(csa_tree_add_7_27_groupi_n_1856 ,csa_tree_add_7_27_groupi_n_1817 ,in2[2]);
  xnor csa_tree_add_7_27_groupi_g5342__9315(csa_tree_add_7_27_groupi_n_1855 ,csa_tree_add_7_27_groupi_n_1816 ,in2[14]);
  xnor csa_tree_add_7_27_groupi_g5343__9945(csa_tree_add_7_27_groupi_n_1854 ,csa_tree_add_7_27_groupi_n_1814 ,csa_tree_add_7_27_groupi_n_1774);
  and csa_tree_add_7_27_groupi_g5344__2883(csa_tree_add_7_27_groupi_n_1845 ,csa_tree_add_7_27_groupi_n_1814 ,csa_tree_add_7_27_groupi_n_1765);
  and csa_tree_add_7_27_groupi_g5345__2346(csa_tree_add_7_27_groupi_n_1844 ,csa_tree_add_7_27_groupi_n_1812 ,csa_tree_add_7_27_groupi_n_1786);
  or csa_tree_add_7_27_groupi_g5346__1666(csa_tree_add_7_27_groupi_n_1843 ,csa_tree_add_7_27_groupi_n_1812 ,csa_tree_add_7_27_groupi_n_1786);
  or csa_tree_add_7_27_groupi_g5347__7410(csa_tree_add_7_27_groupi_n_1842 ,csa_tree_add_7_27_groupi_n_1811 ,csa_tree_add_7_27_groupi_n_1787);
  and csa_tree_add_7_27_groupi_g5348__6417(csa_tree_add_7_27_groupi_n_1841 ,csa_tree_add_7_27_groupi_n_1811 ,csa_tree_add_7_27_groupi_n_1787);
  or csa_tree_add_7_27_groupi_g5349__5477(csa_tree_add_7_27_groupi_n_1840 ,csa_tree_add_7_27_groupi_n_1103 ,csa_tree_add_7_27_groupi_n_1822);
  and csa_tree_add_7_27_groupi_g5350__2398(csa_tree_add_7_27_groupi_n_1839 ,csa_tree_add_7_27_groupi_n_1813 ,csa_tree_add_7_27_groupi_n_1785);
  or csa_tree_add_7_27_groupi_g5351__5107(csa_tree_add_7_27_groupi_n_1838 ,csa_tree_add_7_27_groupi_n_1813 ,csa_tree_add_7_27_groupi_n_1785);
  or csa_tree_add_7_27_groupi_g5352__6260(csa_tree_add_7_27_groupi_n_1837 ,csa_tree_add_7_27_groupi_n_1089 ,csa_tree_add_7_27_groupi_n_1821);
  and csa_tree_add_7_27_groupi_g5353__4319(csa_tree_add_7_27_groupi_n_1846 ,csa_tree_add_7_27_groupi_n_766 ,csa_tree_add_7_27_groupi_n_1825);
  or csa_tree_add_7_27_groupi_g5354__8428(csa_tree_add_7_27_groupi_n_1834 ,csa_tree_add_7_27_groupi_n_1220 ,csa_tree_add_7_27_groupi_n_1820);
  or csa_tree_add_7_27_groupi_g5355__5526(csa_tree_add_7_27_groupi_n_1833 ,csa_tree_add_7_27_groupi_n_1195 ,csa_tree_add_7_27_groupi_n_1806);
  or csa_tree_add_7_27_groupi_g5356__6783(csa_tree_add_7_27_groupi_n_1832 ,csa_tree_add_7_27_groupi_n_1407 ,csa_tree_add_7_27_groupi_n_1810);
  nor csa_tree_add_7_27_groupi_g5357__3680(csa_tree_add_7_27_groupi_n_1831 ,csa_tree_add_7_27_groupi_n_1408 ,csa_tree_add_7_27_groupi_n_1809);
  xnor csa_tree_add_7_27_groupi_g5358__1617(n_9 ,csa_tree_add_7_27_groupi_n_1799 ,csa_tree_add_7_27_groupi_n_1745);
  or csa_tree_add_7_27_groupi_g5359__2802(csa_tree_add_7_27_groupi_n_1829 ,csa_tree_add_7_27_groupi_n_1037 ,csa_tree_add_7_27_groupi_n_1823);
  nor csa_tree_add_7_27_groupi_g5360__1705(csa_tree_add_7_27_groupi_n_1828 ,csa_tree_add_7_27_groupi_n_1772 ,csa_tree_add_7_27_groupi_n_1808);
  or csa_tree_add_7_27_groupi_g5361__5122(csa_tree_add_7_27_groupi_n_1827 ,csa_tree_add_7_27_groupi_n_1773 ,csa_tree_add_7_27_groupi_n_1807);
  or csa_tree_add_7_27_groupi_g5362__8246(csa_tree_add_7_27_groupi_n_1836 ,csa_tree_add_7_27_groupi_n_1721 ,csa_tree_add_7_27_groupi_n_1824);
  xnor csa_tree_add_7_27_groupi_g5363__7098(csa_tree_add_7_27_groupi_n_1835 ,csa_tree_add_7_27_groupi_n_1800 ,csa_tree_add_7_27_groupi_n_847);
  or csa_tree_add_7_27_groupi_g5364__6131(csa_tree_add_7_27_groupi_n_1825 ,csa_tree_add_7_27_groupi_n_809 ,csa_tree_add_7_27_groupi_n_1800);
  and csa_tree_add_7_27_groupi_g5365__1881(csa_tree_add_7_27_groupi_n_1824 ,csa_tree_add_7_27_groupi_n_1720 ,csa_tree_add_7_27_groupi_n_1799);
  nor csa_tree_add_7_27_groupi_g5366__5115(csa_tree_add_7_27_groupi_n_1823 ,csa_tree_add_7_27_groupi_n_437 ,csa_tree_add_7_27_groupi_n_538);
  nor csa_tree_add_7_27_groupi_g5367__7482(csa_tree_add_7_27_groupi_n_1822 ,csa_tree_add_7_27_groupi_n_380 ,csa_tree_add_7_27_groupi_n_1784);
  nor csa_tree_add_7_27_groupi_g5368__4733(csa_tree_add_7_27_groupi_n_1821 ,csa_tree_add_7_27_groupi_n_453 ,csa_tree_add_7_27_groupi_n_538);
  nor csa_tree_add_7_27_groupi_g5369__6161(csa_tree_add_7_27_groupi_n_1820 ,csa_tree_add_7_27_groupi_n_407 ,csa_tree_add_7_27_groupi_n_1784);
  nor csa_tree_add_7_27_groupi_g5370__9315(csa_tree_add_7_27_groupi_n_1819 ,csa_tree_add_7_27_groupi_n_1345 ,csa_tree_add_7_27_groupi_n_1793);
  nor csa_tree_add_7_27_groupi_g5371__9945(csa_tree_add_7_27_groupi_n_1818 ,csa_tree_add_7_27_groupi_n_1364 ,csa_tree_add_7_27_groupi_n_1792);
  nor csa_tree_add_7_27_groupi_g5372__2883(csa_tree_add_7_27_groupi_n_1817 ,csa_tree_add_7_27_groupi_n_1121 ,csa_tree_add_7_27_groupi_n_1779);
  nor csa_tree_add_7_27_groupi_g5373__2346(csa_tree_add_7_27_groupi_n_1816 ,csa_tree_add_7_27_groupi_n_1329 ,csa_tree_add_7_27_groupi_n_1789);
  nor csa_tree_add_7_27_groupi_g5374__1666(csa_tree_add_7_27_groupi_n_1815 ,csa_tree_add_7_27_groupi_n_1290 ,csa_tree_add_7_27_groupi_n_1775);
  or csa_tree_add_7_27_groupi_g5375__7410(csa_tree_add_7_27_groupi_n_1826 ,csa_tree_add_7_27_groupi_n_1178 ,csa_tree_add_7_27_groupi_n_1782);
  not csa_tree_add_7_27_groupi_g5376(csa_tree_add_7_27_groupi_n_1809 ,csa_tree_add_7_27_groupi_n_1810);
  not csa_tree_add_7_27_groupi_g5377(csa_tree_add_7_27_groupi_n_1807 ,csa_tree_add_7_27_groupi_n_1808);
  nor csa_tree_add_7_27_groupi_g5378__6417(csa_tree_add_7_27_groupi_n_1806 ,csa_tree_add_7_27_groupi_n_425 ,csa_tree_add_7_27_groupi_n_537);
  xnor csa_tree_add_7_27_groupi_g5379__5477(csa_tree_add_7_27_groupi_n_1805 ,csa_tree_add_7_27_groupi_n_1756 ,csa_tree_add_7_27_groupi_n_1730);
  xnor csa_tree_add_7_27_groupi_g5380__2398(csa_tree_add_7_27_groupi_n_1804 ,csa_tree_add_7_27_groupi_n_1755 ,csa_tree_add_7_27_groupi_n_1729);
  xnor csa_tree_add_7_27_groupi_g5381__5107(csa_tree_add_7_27_groupi_n_1803 ,csa_tree_add_7_27_groupi_n_1754 ,csa_tree_add_7_27_groupi_n_1728);
  xnor csa_tree_add_7_27_groupi_g5382__6260(csa_tree_add_7_27_groupi_n_1802 ,csa_tree_add_7_27_groupi_n_1718 ,csa_tree_add_7_27_groupi_n_1753);
  xnor csa_tree_add_7_27_groupi_g5383__4319(csa_tree_add_7_27_groupi_n_1801 ,csa_tree_add_7_27_groupi_n_1757 ,csa_tree_add_7_27_groupi_n_1726);
  xnor csa_tree_add_7_27_groupi_g5384__8428(csa_tree_add_7_27_groupi_n_1814 ,csa_tree_add_7_27_groupi_n_1763 ,in2[11]);
  xnor csa_tree_add_7_27_groupi_g5385__5526(csa_tree_add_7_27_groupi_n_1813 ,csa_tree_add_7_27_groupi_n_1762 ,in2[2]);
  xnor csa_tree_add_7_27_groupi_g5386__6783(csa_tree_add_7_27_groupi_n_1812 ,csa_tree_add_7_27_groupi_n_1759 ,in2[8]);
  xnor csa_tree_add_7_27_groupi_g5387__3680(csa_tree_add_7_27_groupi_n_1811 ,csa_tree_add_7_27_groupi_n_1761 ,in2[5]);
  xnor csa_tree_add_7_27_groupi_g5388__1617(csa_tree_add_7_27_groupi_n_1810 ,csa_tree_add_7_27_groupi_n_1760 ,in2[14]);
  xnor csa_tree_add_7_27_groupi_g5389__2802(csa_tree_add_7_27_groupi_n_1808 ,csa_tree_add_7_27_groupi_n_1758 ,csa_tree_add_7_27_groupi_n_1300);
  and csa_tree_add_7_27_groupi_g5390__1705(csa_tree_add_7_27_groupi_n_1795 ,csa_tree_add_7_27_groupi_n_1756 ,csa_tree_add_7_27_groupi_n_1730);
  or csa_tree_add_7_27_groupi_g5391__5122(csa_tree_add_7_27_groupi_n_1794 ,csa_tree_add_7_27_groupi_n_1755 ,csa_tree_add_7_27_groupi_n_1729);
  or csa_tree_add_7_27_groupi_g5392__8246(csa_tree_add_7_27_groupi_n_1793 ,csa_tree_add_7_27_groupi_n_1102 ,csa_tree_add_7_27_groupi_n_1749);
  or csa_tree_add_7_27_groupi_g5393__7098(csa_tree_add_7_27_groupi_n_1792 ,csa_tree_add_7_27_groupi_n_1144 ,csa_tree_add_7_27_groupi_n_1751);
  and csa_tree_add_7_27_groupi_g5394__6131(csa_tree_add_7_27_groupi_n_1791 ,csa_tree_add_7_27_groupi_n_1755 ,csa_tree_add_7_27_groupi_n_1729);
  or csa_tree_add_7_27_groupi_g5395__1881(csa_tree_add_7_27_groupi_n_1790 ,csa_tree_add_7_27_groupi_n_1756 ,csa_tree_add_7_27_groupi_n_1730);
  or csa_tree_add_7_27_groupi_g5396__5115(csa_tree_add_7_27_groupi_n_1789 ,csa_tree_add_7_27_groupi_n_1092 ,csa_tree_add_7_27_groupi_n_1752);
  or csa_tree_add_7_27_groupi_g5397__7482(csa_tree_add_7_27_groupi_n_1788 ,csa_tree_add_7_27_groupi_n_1754 ,csa_tree_add_7_27_groupi_n_1728);
  and csa_tree_add_7_27_groupi_g5398__4733(csa_tree_add_7_27_groupi_n_1800 ,csa_tree_add_7_27_groupi_n_798 ,csa_tree_add_7_27_groupi_n_1768);
  or csa_tree_add_7_27_groupi_g5399__6161(csa_tree_add_7_27_groupi_n_1799 ,csa_tree_add_7_27_groupi_n_1681 ,csa_tree_add_7_27_groupi_n_1769);
  or csa_tree_add_7_27_groupi_g5400__9315(csa_tree_add_7_27_groupi_n_1798 ,csa_tree_add_7_27_groupi_n_1680 ,csa_tree_add_7_27_groupi_n_1767);
  or csa_tree_add_7_27_groupi_g5401__9945(csa_tree_add_7_27_groupi_n_1797 ,csa_tree_add_7_27_groupi_n_1686 ,csa_tree_add_7_27_groupi_n_1770);
  or csa_tree_add_7_27_groupi_g5402__2883(csa_tree_add_7_27_groupi_n_1796 ,csa_tree_add_7_27_groupi_n_1684 ,csa_tree_add_7_27_groupi_n_1764);
  xnor csa_tree_add_7_27_groupi_g5403__2346(csa_tree_add_7_27_groupi_n_1783 ,csa_tree_add_7_27_groupi_n_1731 ,csa_tree_add_7_27_groupi_n_1692);
  and csa_tree_add_7_27_groupi_g5404__1666(csa_tree_add_7_27_groupi_n_1782 ,csa_tree_add_7_27_groupi_n_1181 ,csa_tree_add_7_27_groupi_n_1758);
  and csa_tree_add_7_27_groupi_g5405__7410(csa_tree_add_7_27_groupi_n_1781 ,csa_tree_add_7_27_groupi_n_1757 ,csa_tree_add_7_27_groupi_n_1726);
  or csa_tree_add_7_27_groupi_g5406__6417(csa_tree_add_7_27_groupi_n_1780 ,csa_tree_add_7_27_groupi_n_1757 ,csa_tree_add_7_27_groupi_n_1726);
  or csa_tree_add_7_27_groupi_g5407__5477(csa_tree_add_7_27_groupi_n_1779 ,csa_tree_add_7_27_groupi_n_1011 ,csa_tree_add_7_27_groupi_n_1771);
  and csa_tree_add_7_27_groupi_g5408__2398(csa_tree_add_7_27_groupi_n_1778 ,csa_tree_add_7_27_groupi_n_1718 ,csa_tree_add_7_27_groupi_n_1753);
  or csa_tree_add_7_27_groupi_g5409__5107(csa_tree_add_7_27_groupi_n_1777 ,csa_tree_add_7_27_groupi_n_1718 ,csa_tree_add_7_27_groupi_n_1753);
  and csa_tree_add_7_27_groupi_g5410__6260(csa_tree_add_7_27_groupi_n_1776 ,csa_tree_add_7_27_groupi_n_1754 ,csa_tree_add_7_27_groupi_n_1728);
  or csa_tree_add_7_27_groupi_g5411__4319(csa_tree_add_7_27_groupi_n_1775 ,csa_tree_add_7_27_groupi_n_1204 ,csa_tree_add_7_27_groupi_n_1750);
  xnor csa_tree_add_7_27_groupi_g5412__8428(csa_tree_add_7_27_groupi_n_1774 ,csa_tree_add_7_27_groupi_n_1700 ,csa_tree_add_7_27_groupi_n_1727);
  xnor csa_tree_add_7_27_groupi_g5413__5526(csa_tree_add_7_27_groupi_n_1787 ,csa_tree_add_7_27_groupi_n_1742 ,csa_tree_add_7_27_groupi_n_1694);
  xnor csa_tree_add_7_27_groupi_g5414__6783(csa_tree_add_7_27_groupi_n_1786 ,csa_tree_add_7_27_groupi_n_1741 ,csa_tree_add_7_27_groupi_n_1693);
  xnor csa_tree_add_7_27_groupi_g5415__3680(csa_tree_add_7_27_groupi_n_1785 ,csa_tree_add_7_27_groupi_n_1743 ,csa_tree_add_7_27_groupi_n_1695);
  xnor csa_tree_add_7_27_groupi_g5416__1617(csa_tree_add_7_27_groupi_n_1784 ,csa_tree_add_7_27_groupi_n_1744 ,csa_tree_add_7_27_groupi_n_837);
  not csa_tree_add_7_27_groupi_g5417(csa_tree_add_7_27_groupi_n_1772 ,csa_tree_add_7_27_groupi_n_1773);
  nor csa_tree_add_7_27_groupi_g5418__2802(csa_tree_add_7_27_groupi_n_1771 ,csa_tree_add_7_27_groupi_n_305 ,csa_tree_add_7_27_groupi_n_527);
  and csa_tree_add_7_27_groupi_g5419__1705(csa_tree_add_7_27_groupi_n_1770 ,csa_tree_add_7_27_groupi_n_1685 ,csa_tree_add_7_27_groupi_n_1741);
  and csa_tree_add_7_27_groupi_g5420__5122(csa_tree_add_7_27_groupi_n_1769 ,csa_tree_add_7_27_groupi_n_1670 ,csa_tree_add_7_27_groupi_n_1731);
  or csa_tree_add_7_27_groupi_g5421__8246(csa_tree_add_7_27_groupi_n_1768 ,csa_tree_add_7_27_groupi_n_783 ,csa_tree_add_7_27_groupi_n_1744);
  and csa_tree_add_7_27_groupi_g5422__7098(csa_tree_add_7_27_groupi_n_1767 ,csa_tree_add_7_27_groupi_n_1679 ,csa_tree_add_7_27_groupi_n_1742);
  and csa_tree_add_7_27_groupi_g5423__6131(csa_tree_add_7_27_groupi_n_1766 ,csa_tree_add_7_27_groupi_n_1700 ,csa_tree_add_7_27_groupi_n_1727);
  or csa_tree_add_7_27_groupi_g5424__1881(csa_tree_add_7_27_groupi_n_1765 ,csa_tree_add_7_27_groupi_n_1700 ,csa_tree_add_7_27_groupi_n_1727);
  and csa_tree_add_7_27_groupi_g5425__5115(csa_tree_add_7_27_groupi_n_1764 ,csa_tree_add_7_27_groupi_n_1671 ,csa_tree_add_7_27_groupi_n_1743);
  nor csa_tree_add_7_27_groupi_g5426__7482(csa_tree_add_7_27_groupi_n_1763 ,csa_tree_add_7_27_groupi_n_1322 ,csa_tree_add_7_27_groupi_n_1734);
  nor csa_tree_add_7_27_groupi_g5427__4733(csa_tree_add_7_27_groupi_n_1762 ,csa_tree_add_7_27_groupi_n_1110 ,csa_tree_add_7_27_groupi_n_1719);
  nor csa_tree_add_7_27_groupi_g5428__6161(csa_tree_add_7_27_groupi_n_1761 ,csa_tree_add_7_27_groupi_n_1287 ,csa_tree_add_7_27_groupi_n_1724);
  nor csa_tree_add_7_27_groupi_g5429__9315(csa_tree_add_7_27_groupi_n_1760 ,csa_tree_add_7_27_groupi_n_1343 ,csa_tree_add_7_27_groupi_n_1740);
  nor csa_tree_add_7_27_groupi_g5430__9945(csa_tree_add_7_27_groupi_n_1759 ,csa_tree_add_7_27_groupi_n_1259 ,csa_tree_add_7_27_groupi_n_1723);
  or csa_tree_add_7_27_groupi_g5431__2883(csa_tree_add_7_27_groupi_n_1773 ,csa_tree_add_7_27_groupi_n_1316 ,csa_tree_add_7_27_groupi_n_1736);
  nor csa_tree_add_7_27_groupi_g5432__2346(csa_tree_add_7_27_groupi_n_1752 ,csa_tree_add_7_27_groupi_n_317 ,csa_tree_add_7_27_groupi_n_1725);
  nor csa_tree_add_7_27_groupi_g5433__1666(csa_tree_add_7_27_groupi_n_1751 ,csa_tree_add_7_27_groupi_n_344 ,csa_tree_add_7_27_groupi_n_527);
  nor csa_tree_add_7_27_groupi_g5434__7410(csa_tree_add_7_27_groupi_n_1750 ,csa_tree_add_7_27_groupi_n_284 ,csa_tree_add_7_27_groupi_n_1725);
  nor csa_tree_add_7_27_groupi_g5435__6417(csa_tree_add_7_27_groupi_n_1749 ,csa_tree_add_7_27_groupi_n_269 ,csa_tree_add_7_27_groupi_n_526);
  xnor csa_tree_add_7_27_groupi_g5436__5477(csa_tree_add_7_27_groupi_n_1748 ,csa_tree_add_7_27_groupi_n_1704 ,csa_tree_add_7_27_groupi_n_1675);
  xnor csa_tree_add_7_27_groupi_g5437__2398(csa_tree_add_7_27_groupi_n_1747 ,csa_tree_add_7_27_groupi_n_1703 ,csa_tree_add_7_27_groupi_n_1674);
  xnor csa_tree_add_7_27_groupi_g5438__5107(csa_tree_add_7_27_groupi_n_1746 ,csa_tree_add_7_27_groupi_n_1702 ,csa_tree_add_7_27_groupi_n_1673);
  xnor csa_tree_add_7_27_groupi_g5439__6260(csa_tree_add_7_27_groupi_n_1745 ,csa_tree_add_7_27_groupi_n_1701 ,csa_tree_add_7_27_groupi_n_1676);
  xnor csa_tree_add_7_27_groupi_g5440__4319(csa_tree_add_7_27_groupi_n_1758 ,csa_tree_add_7_27_groupi_n_1708 ,in2[14]);
  xnor csa_tree_add_7_27_groupi_g5441__8428(csa_tree_add_7_27_groupi_n_1757 ,csa_tree_add_7_27_groupi_n_1707 ,in2[11]);
  xnor csa_tree_add_7_27_groupi_g5442__5526(csa_tree_add_7_27_groupi_n_1756 ,csa_tree_add_7_27_groupi_n_1706 ,in2[5]);
  xnor csa_tree_add_7_27_groupi_g5443__6783(csa_tree_add_7_27_groupi_n_1755 ,csa_tree_add_7_27_groupi_n_1710 ,in2[8]);
  xnor csa_tree_add_7_27_groupi_g5444__3680(csa_tree_add_7_27_groupi_n_1754 ,csa_tree_add_7_27_groupi_n_1709 ,in2[2]);
  xnor csa_tree_add_7_27_groupi_g5445__1617(csa_tree_add_7_27_groupi_n_1753 ,csa_tree_add_7_27_groupi_n_1705 ,csa_tree_add_7_27_groupi_n_1372);
  or csa_tree_add_7_27_groupi_g5446__2802(csa_tree_add_7_27_groupi_n_1740 ,csa_tree_add_7_27_groupi_n_1130 ,csa_tree_add_7_27_groupi_n_1697);
  and csa_tree_add_7_27_groupi_g5447__1705(csa_tree_add_7_27_groupi_n_1739 ,csa_tree_add_7_27_groupi_n_1702 ,csa_tree_add_7_27_groupi_n_1673);
  or csa_tree_add_7_27_groupi_g5448__5122(csa_tree_add_7_27_groupi_n_1738 ,csa_tree_add_7_27_groupi_n_1702 ,csa_tree_add_7_27_groupi_n_1673);
  or csa_tree_add_7_27_groupi_g5449__8246(csa_tree_add_7_27_groupi_n_1737 ,csa_tree_add_7_27_groupi_n_1704 ,csa_tree_add_7_27_groupi_n_1675);
  and csa_tree_add_7_27_groupi_g5450__7098(csa_tree_add_7_27_groupi_n_1736 ,csa_tree_add_7_27_groupi_n_1317 ,csa_tree_add_7_27_groupi_n_1705);
  and csa_tree_add_7_27_groupi_g5451__6131(csa_tree_add_7_27_groupi_n_1735 ,csa_tree_add_7_27_groupi_n_1704 ,csa_tree_add_7_27_groupi_n_1675);
  or csa_tree_add_7_27_groupi_g5452__1881(csa_tree_add_7_27_groupi_n_1734 ,csa_tree_add_7_27_groupi_n_1134 ,csa_tree_add_7_27_groupi_n_1699);
  and csa_tree_add_7_27_groupi_g5453__5115(csa_tree_add_7_27_groupi_n_1733 ,csa_tree_add_7_27_groupi_n_1703 ,csa_tree_add_7_27_groupi_n_1674);
  or csa_tree_add_7_27_groupi_g5454__7482(csa_tree_add_7_27_groupi_n_1732 ,csa_tree_add_7_27_groupi_n_1703 ,csa_tree_add_7_27_groupi_n_1674);
  and csa_tree_add_7_27_groupi_g5455__4733(csa_tree_add_7_27_groupi_n_1744 ,csa_tree_add_7_27_groupi_n_768 ,csa_tree_add_7_27_groupi_n_1716);
  or csa_tree_add_7_27_groupi_g5456__6161(csa_tree_add_7_27_groupi_n_1743 ,csa_tree_add_7_27_groupi_n_1632 ,csa_tree_add_7_27_groupi_n_1713);
  or csa_tree_add_7_27_groupi_g5457__9315(csa_tree_add_7_27_groupi_n_1742 ,csa_tree_add_7_27_groupi_n_1629 ,csa_tree_add_7_27_groupi_n_1714);
  or csa_tree_add_7_27_groupi_g5458__9945(csa_tree_add_7_27_groupi_n_1741 ,csa_tree_add_7_27_groupi_n_1634 ,csa_tree_add_7_27_groupi_n_1711);
  or csa_tree_add_7_27_groupi_g5459__2883(csa_tree_add_7_27_groupi_n_1724 ,csa_tree_add_7_27_groupi_n_1197 ,csa_tree_add_7_27_groupi_n_1696);
  or csa_tree_add_7_27_groupi_g5460__2346(csa_tree_add_7_27_groupi_n_1723 ,csa_tree_add_7_27_groupi_n_1229 ,csa_tree_add_7_27_groupi_n_1698);
  xnor csa_tree_add_7_27_groupi_g5461__1666(n_7 ,csa_tree_add_7_27_groupi_n_1678 ,csa_tree_add_7_27_groupi_n_1644);
  and csa_tree_add_7_27_groupi_g5462__7410(csa_tree_add_7_27_groupi_n_1721 ,csa_tree_add_7_27_groupi_n_1701 ,csa_tree_add_7_27_groupi_n_1676);
  or csa_tree_add_7_27_groupi_g5463__6417(csa_tree_add_7_27_groupi_n_1720 ,csa_tree_add_7_27_groupi_n_1701 ,csa_tree_add_7_27_groupi_n_1676);
  or csa_tree_add_7_27_groupi_g5464__5477(csa_tree_add_7_27_groupi_n_1719 ,csa_tree_add_7_27_groupi_n_1019 ,csa_tree_add_7_27_groupi_n_1715);
  or csa_tree_add_7_27_groupi_g5465__2398(csa_tree_add_7_27_groupi_n_1731 ,csa_tree_add_7_27_groupi_n_1631 ,csa_tree_add_7_27_groupi_n_1712);
  xnor csa_tree_add_7_27_groupi_g5466__5107(csa_tree_add_7_27_groupi_n_1730 ,csa_tree_add_7_27_groupi_n_1689 ,csa_tree_add_7_27_groupi_n_1642);
  xnor csa_tree_add_7_27_groupi_g5467__6260(csa_tree_add_7_27_groupi_n_1729 ,csa_tree_add_7_27_groupi_n_1688 ,csa_tree_add_7_27_groupi_n_1643);
  xnor csa_tree_add_7_27_groupi_g5468__4319(csa_tree_add_7_27_groupi_n_1728 ,csa_tree_add_7_27_groupi_n_1677 ,csa_tree_add_7_27_groupi_n_1641);
  or csa_tree_add_7_27_groupi_g5469__8428(csa_tree_add_7_27_groupi_n_1727 ,csa_tree_add_7_27_groupi_n_1616 ,csa_tree_add_7_27_groupi_n_1717);
  xnor csa_tree_add_7_27_groupi_g5470__5526(csa_tree_add_7_27_groupi_n_1726 ,csa_tree_add_7_27_groupi_n_1690 ,csa_tree_add_7_27_groupi_n_1645);
  xnor csa_tree_add_7_27_groupi_g5471__6783(csa_tree_add_7_27_groupi_n_1725 ,csa_tree_add_7_27_groupi_n_1691 ,csa_tree_add_7_27_groupi_n_830);
  and csa_tree_add_7_27_groupi_g5472__3680(csa_tree_add_7_27_groupi_n_1717 ,csa_tree_add_7_27_groupi_n_1615 ,csa_tree_add_7_27_groupi_n_1690);
  or csa_tree_add_7_27_groupi_g5473__1617(csa_tree_add_7_27_groupi_n_1716 ,csa_tree_add_7_27_groupi_n_795 ,csa_tree_add_7_27_groupi_n_1691);
  nor csa_tree_add_7_27_groupi_g5474__2802(csa_tree_add_7_27_groupi_n_1715 ,csa_tree_add_7_27_groupi_n_98 ,csa_tree_add_7_27_groupi_n_555);
  and csa_tree_add_7_27_groupi_g5475__1705(csa_tree_add_7_27_groupi_n_1714 ,csa_tree_add_7_27_groupi_n_1628 ,csa_tree_add_7_27_groupi_n_1689);
  and csa_tree_add_7_27_groupi_g5476__5122(csa_tree_add_7_27_groupi_n_1713 ,csa_tree_add_7_27_groupi_n_1636 ,csa_tree_add_7_27_groupi_n_1677);
  and csa_tree_add_7_27_groupi_g5477__8246(csa_tree_add_7_27_groupi_n_1712 ,csa_tree_add_7_27_groupi_n_1619 ,csa_tree_add_7_27_groupi_n_1678);
  and csa_tree_add_7_27_groupi_g5478__7098(csa_tree_add_7_27_groupi_n_1711 ,csa_tree_add_7_27_groupi_n_1635 ,csa_tree_add_7_27_groupi_n_1688);
  nor csa_tree_add_7_27_groupi_g5479__6131(csa_tree_add_7_27_groupi_n_1710 ,csa_tree_add_7_27_groupi_n_1341 ,csa_tree_add_7_27_groupi_n_1683);
  nor csa_tree_add_7_27_groupi_g5480__1881(csa_tree_add_7_27_groupi_n_1709 ,csa_tree_add_7_27_groupi_n_1117 ,csa_tree_add_7_27_groupi_n_1666);
  nor csa_tree_add_7_27_groupi_g5481__5115(csa_tree_add_7_27_groupi_n_1708 ,csa_tree_add_7_27_groupi_n_1342 ,csa_tree_add_7_27_groupi_n_1687);
  nor csa_tree_add_7_27_groupi_g5482__7482(csa_tree_add_7_27_groupi_n_1707 ,csa_tree_add_7_27_groupi_n_1257 ,csa_tree_add_7_27_groupi_n_1668);
  nor csa_tree_add_7_27_groupi_g5483__4733(csa_tree_add_7_27_groupi_n_1706 ,csa_tree_add_7_27_groupi_n_1263 ,csa_tree_add_7_27_groupi_n_1669);
  or csa_tree_add_7_27_groupi_g5484__6161(csa_tree_add_7_27_groupi_n_1718 ,csa_tree_add_7_27_groupi_n_1390 ,csa_tree_add_7_27_groupi_n_1682);
  nor csa_tree_add_7_27_groupi_g5485__9315(csa_tree_add_7_27_groupi_n_1699 ,csa_tree_add_7_27_groupi_n_100 ,csa_tree_add_7_27_groupi_n_1672);
  nor csa_tree_add_7_27_groupi_g5486__9945(csa_tree_add_7_27_groupi_n_1698 ,csa_tree_add_7_27_groupi_n_102 ,csa_tree_add_7_27_groupi_n_555);
  nor csa_tree_add_7_27_groupi_g5487__2883(csa_tree_add_7_27_groupi_n_1697 ,csa_tree_add_7_27_groupi_n_106 ,csa_tree_add_7_27_groupi_n_1672);
  nor csa_tree_add_7_27_groupi_g5488__2346(csa_tree_add_7_27_groupi_n_1696 ,csa_tree_add_7_27_groupi_n_104 ,csa_tree_add_7_27_groupi_n_554);
  xnor csa_tree_add_7_27_groupi_g5489__1666(csa_tree_add_7_27_groupi_n_1695 ,csa_tree_add_7_27_groupi_n_1650 ,csa_tree_add_7_27_groupi_n_1621);
  xnor csa_tree_add_7_27_groupi_g5490__7410(csa_tree_add_7_27_groupi_n_1694 ,csa_tree_add_7_27_groupi_n_1651 ,csa_tree_add_7_27_groupi_n_1624);
  xnor csa_tree_add_7_27_groupi_g5491__6417(csa_tree_add_7_27_groupi_n_1693 ,csa_tree_add_7_27_groupi_n_1648 ,csa_tree_add_7_27_groupi_n_1623);
  xnor csa_tree_add_7_27_groupi_g5492__5477(csa_tree_add_7_27_groupi_n_1692 ,csa_tree_add_7_27_groupi_n_1649 ,csa_tree_add_7_27_groupi_n_1622);
  xnor csa_tree_add_7_27_groupi_g5493__2398(csa_tree_add_7_27_groupi_n_1705 ,csa_tree_add_7_27_groupi_n_1655 ,in2[14]);
  xnor csa_tree_add_7_27_groupi_g5494__5107(csa_tree_add_7_27_groupi_n_1704 ,csa_tree_add_7_27_groupi_n_1654 ,in2[5]);
  xnor csa_tree_add_7_27_groupi_g5495__6260(csa_tree_add_7_27_groupi_n_1703 ,csa_tree_add_7_27_groupi_n_1653 ,in2[8]);
  xnor csa_tree_add_7_27_groupi_g5496__4319(csa_tree_add_7_27_groupi_n_1702 ,csa_tree_add_7_27_groupi_n_1656 ,in2[11]);
  xnor csa_tree_add_7_27_groupi_g5497__8428(csa_tree_add_7_27_groupi_n_1701 ,csa_tree_add_7_27_groupi_n_1657 ,in2[2]);
  xnor csa_tree_add_7_27_groupi_g5498__5526(csa_tree_add_7_27_groupi_n_1700 ,csa_tree_add_7_27_groupi_n_1652 ,csa_tree_add_7_27_groupi_n_1394);
  or csa_tree_add_7_27_groupi_g5499__6783(csa_tree_add_7_27_groupi_n_1687 ,csa_tree_add_7_27_groupi_n_1091 ,csa_tree_add_7_27_groupi_n_1647);
  and csa_tree_add_7_27_groupi_g5500__3680(csa_tree_add_7_27_groupi_n_1686 ,csa_tree_add_7_27_groupi_n_1648 ,csa_tree_add_7_27_groupi_n_1623);
  or csa_tree_add_7_27_groupi_g5501__1617(csa_tree_add_7_27_groupi_n_1685 ,csa_tree_add_7_27_groupi_n_1648 ,csa_tree_add_7_27_groupi_n_1623);
  and csa_tree_add_7_27_groupi_g5502__2802(csa_tree_add_7_27_groupi_n_1684 ,csa_tree_add_7_27_groupi_n_1650 ,csa_tree_add_7_27_groupi_n_1621);
  or csa_tree_add_7_27_groupi_g5503__1705(csa_tree_add_7_27_groupi_n_1683 ,csa_tree_add_7_27_groupi_n_1114 ,csa_tree_add_7_27_groupi_n_1646);
  and csa_tree_add_7_27_groupi_g5504__5122(csa_tree_add_7_27_groupi_n_1682 ,csa_tree_add_7_27_groupi_n_1386 ,csa_tree_add_7_27_groupi_n_1652);
  and csa_tree_add_7_27_groupi_g5505__8246(csa_tree_add_7_27_groupi_n_1681 ,csa_tree_add_7_27_groupi_n_1649 ,csa_tree_add_7_27_groupi_n_1622);
  and csa_tree_add_7_27_groupi_g5506__7098(csa_tree_add_7_27_groupi_n_1680 ,csa_tree_add_7_27_groupi_n_1651 ,csa_tree_add_7_27_groupi_n_1624);
  or csa_tree_add_7_27_groupi_g5507__6131(csa_tree_add_7_27_groupi_n_1679 ,csa_tree_add_7_27_groupi_n_1651 ,csa_tree_add_7_27_groupi_n_1624);
  and csa_tree_add_7_27_groupi_g5508__1881(csa_tree_add_7_27_groupi_n_1691 ,csa_tree_add_7_27_groupi_n_787 ,csa_tree_add_7_27_groupi_n_1663);
  or csa_tree_add_7_27_groupi_g5509__5115(csa_tree_add_7_27_groupi_n_1690 ,csa_tree_add_7_27_groupi_n_1574 ,csa_tree_add_7_27_groupi_n_1662);
  or csa_tree_add_7_27_groupi_g5510__7482(csa_tree_add_7_27_groupi_n_1689 ,csa_tree_add_7_27_groupi_n_1576 ,csa_tree_add_7_27_groupi_n_1664);
  or csa_tree_add_7_27_groupi_g5511__4733(csa_tree_add_7_27_groupi_n_1688 ,csa_tree_add_7_27_groupi_n_1579 ,csa_tree_add_7_27_groupi_n_1661);
  or csa_tree_add_7_27_groupi_g5512__6161(csa_tree_add_7_27_groupi_n_1671 ,csa_tree_add_7_27_groupi_n_1650 ,csa_tree_add_7_27_groupi_n_1621);
  or csa_tree_add_7_27_groupi_g5513__9315(csa_tree_add_7_27_groupi_n_1670 ,csa_tree_add_7_27_groupi_n_1649 ,csa_tree_add_7_27_groupi_n_1622);
  or csa_tree_add_7_27_groupi_g5514__9945(csa_tree_add_7_27_groupi_n_1669 ,csa_tree_add_7_27_groupi_n_1214 ,csa_tree_add_7_27_groupi_n_1658);
  or csa_tree_add_7_27_groupi_g5515__2883(csa_tree_add_7_27_groupi_n_1668 ,csa_tree_add_7_27_groupi_n_1199 ,csa_tree_add_7_27_groupi_n_0);
  xnor csa_tree_add_7_27_groupi_g5516__2346(n_6 ,csa_tree_add_7_27_groupi_n_1625 ,csa_tree_add_7_27_groupi_n_1613);
  or csa_tree_add_7_27_groupi_g5517__1666(csa_tree_add_7_27_groupi_n_1666 ,csa_tree_add_7_27_groupi_n_1015 ,csa_tree_add_7_27_groupi_n_1659);
  or csa_tree_add_7_27_groupi_g5518__7410(csa_tree_add_7_27_groupi_n_1678 ,csa_tree_add_7_27_groupi_n_1605 ,csa_tree_add_7_27_groupi_n_1665);
  or csa_tree_add_7_27_groupi_g5519__6417(csa_tree_add_7_27_groupi_n_1677 ,csa_tree_add_7_27_groupi_n_1562 ,csa_tree_add_7_27_groupi_n_1660);
  xnor csa_tree_add_7_27_groupi_g5520__5477(csa_tree_add_7_27_groupi_n_1676 ,csa_tree_add_7_27_groupi_n_1626 ,csa_tree_add_7_27_groupi_n_1586);
  xnor csa_tree_add_7_27_groupi_g5521__2398(csa_tree_add_7_27_groupi_n_1675 ,csa_tree_add_7_27_groupi_n_1638 ,csa_tree_add_7_27_groupi_n_1588);
  xnor csa_tree_add_7_27_groupi_g5522__5107(csa_tree_add_7_27_groupi_n_1674 ,csa_tree_add_7_27_groupi_n_1637 ,csa_tree_add_7_27_groupi_n_1587);
  xnor csa_tree_add_7_27_groupi_g5523__6260(csa_tree_add_7_27_groupi_n_1673 ,csa_tree_add_7_27_groupi_n_1639 ,csa_tree_add_7_27_groupi_n_1589);
  xnor csa_tree_add_7_27_groupi_g5524__4319(csa_tree_add_7_27_groupi_n_1672 ,csa_tree_add_7_27_groupi_n_1640 ,csa_tree_add_7_27_groupi_n_838);
  and csa_tree_add_7_27_groupi_g5525__8428(csa_tree_add_7_27_groupi_n_1665 ,csa_tree_add_7_27_groupi_n_1606 ,csa_tree_add_7_27_groupi_n_1625);
  and csa_tree_add_7_27_groupi_g5526__5526(csa_tree_add_7_27_groupi_n_1664 ,csa_tree_add_7_27_groupi_n_1575 ,csa_tree_add_7_27_groupi_n_1638);
  or csa_tree_add_7_27_groupi_g5527__6783(csa_tree_add_7_27_groupi_n_1663 ,csa_tree_add_7_27_groupi_n_799 ,csa_tree_add_7_27_groupi_n_1640);
  and csa_tree_add_7_27_groupi_g5528__3680(csa_tree_add_7_27_groupi_n_1662 ,csa_tree_add_7_27_groupi_n_1573 ,csa_tree_add_7_27_groupi_n_1639);
  and csa_tree_add_7_27_groupi_g5529__1617(csa_tree_add_7_27_groupi_n_1661 ,csa_tree_add_7_27_groupi_n_1578 ,csa_tree_add_7_27_groupi_n_1637);
  and csa_tree_add_7_27_groupi_g5530__2802(csa_tree_add_7_27_groupi_n_1660 ,csa_tree_add_7_27_groupi_n_1563 ,csa_tree_add_7_27_groupi_n_1626);
  nor csa_tree_add_7_27_groupi_g5531__1705(csa_tree_add_7_27_groupi_n_1659 ,csa_tree_add_7_27_groupi_n_34 ,csa_tree_add_7_27_groupi_n_529);
  nor csa_tree_add_7_27_groupi_g5532__5122(csa_tree_add_7_27_groupi_n_1658 ,csa_tree_add_7_27_groupi_n_93 ,csa_tree_add_7_27_groupi_n_1620);
  nor csa_tree_add_7_27_groupi_g5533__8246(csa_tree_add_7_27_groupi_n_1657 ,csa_tree_add_7_27_groupi_n_1125 ,csa_tree_add_7_27_groupi_n_1614);
  nor csa_tree_add_7_27_groupi_g5534__7098(csa_tree_add_7_27_groupi_n_1656 ,csa_tree_add_7_27_groupi_n_1268 ,csa_tree_add_7_27_groupi_n_1617);
  nor csa_tree_add_7_27_groupi_g5535__6131(csa_tree_add_7_27_groupi_n_1655 ,csa_tree_add_7_27_groupi_n_1367 ,csa_tree_add_7_27_groupi_n_1633);
  nor csa_tree_add_7_27_groupi_g5536__1881(csa_tree_add_7_27_groupi_n_1654 ,csa_tree_add_7_27_groupi_n_1351 ,csa_tree_add_7_27_groupi_n_1627);
  nor csa_tree_add_7_27_groupi_g5537__5115(csa_tree_add_7_27_groupi_n_1653 ,csa_tree_add_7_27_groupi_n_1361 ,csa_tree_add_7_27_groupi_n_1630);
  nor csa_tree_add_7_27_groupi_g5538__7482(csa_tree_add_7_27_groupi_n_1647 ,csa_tree_add_7_27_groupi_n_65 ,csa_tree_add_7_27_groupi_n_529);
  nor csa_tree_add_7_27_groupi_g5539__4733(csa_tree_add_7_27_groupi_n_1646 ,csa_tree_add_7_27_groupi_n_47 ,csa_tree_add_7_27_groupi_n_1620);
  xnor csa_tree_add_7_27_groupi_g5541__6161(csa_tree_add_7_27_groupi_n_1645 ,csa_tree_add_7_27_groupi_n_3 ,csa_tree_add_7_27_groupi_n_1595);
  xnor csa_tree_add_7_27_groupi_g5542__9315(csa_tree_add_7_27_groupi_n_1644 ,csa_tree_add_7_27_groupi_n_1596 ,csa_tree_add_7_27_groupi_n_1569);
  xnor csa_tree_add_7_27_groupi_g5543__9945(csa_tree_add_7_27_groupi_n_1643 ,csa_tree_add_7_27_groupi_n_1599 ,csa_tree_add_7_27_groupi_n_1568);
  xnor csa_tree_add_7_27_groupi_g5544__2883(csa_tree_add_7_27_groupi_n_1642 ,csa_tree_add_7_27_groupi_n_1598 ,csa_tree_add_7_27_groupi_n_1571);
  xnor csa_tree_add_7_27_groupi_g5545__2346(csa_tree_add_7_27_groupi_n_1641 ,csa_tree_add_7_27_groupi_n_1597 ,csa_tree_add_7_27_groupi_n_1570);
  xnor csa_tree_add_7_27_groupi_g5546__1666(csa_tree_add_7_27_groupi_n_1652 ,csa_tree_add_7_27_groupi_n_1602 ,in2[14]);
  xnor csa_tree_add_7_27_groupi_g5547__7410(csa_tree_add_7_27_groupi_n_1651 ,csa_tree_add_7_27_groupi_n_1600 ,in2[8]);
  xnor csa_tree_add_7_27_groupi_g5548__6417(csa_tree_add_7_27_groupi_n_1650 ,csa_tree_add_7_27_groupi_n_1601 ,in2[5]);
  xnor csa_tree_add_7_27_groupi_g5549__5477(csa_tree_add_7_27_groupi_n_1649 ,csa_tree_add_7_27_groupi_n_1603 ,in2[2]);
  xnor csa_tree_add_7_27_groupi_g5550__2398(csa_tree_add_7_27_groupi_n_1648 ,csa_tree_add_7_27_groupi_n_1604 ,in2[11]);
  or csa_tree_add_7_27_groupi_g5551__5107(csa_tree_add_7_27_groupi_n_1636 ,csa_tree_add_7_27_groupi_n_1597 ,csa_tree_add_7_27_groupi_n_1570);
  or csa_tree_add_7_27_groupi_g5552__6260(csa_tree_add_7_27_groupi_n_1635 ,csa_tree_add_7_27_groupi_n_1599 ,csa_tree_add_7_27_groupi_n_1568);
  and csa_tree_add_7_27_groupi_g5553__4319(csa_tree_add_7_27_groupi_n_1634 ,csa_tree_add_7_27_groupi_n_1599 ,csa_tree_add_7_27_groupi_n_1568);
  or csa_tree_add_7_27_groupi_g5554__8428(csa_tree_add_7_27_groupi_n_1633 ,csa_tree_add_7_27_groupi_n_1082 ,csa_tree_add_7_27_groupi_n_1593);
  and csa_tree_add_7_27_groupi_g5555__5526(csa_tree_add_7_27_groupi_n_1632 ,csa_tree_add_7_27_groupi_n_1597 ,csa_tree_add_7_27_groupi_n_1570);
  and csa_tree_add_7_27_groupi_g5556__6783(csa_tree_add_7_27_groupi_n_1631 ,csa_tree_add_7_27_groupi_n_1596 ,csa_tree_add_7_27_groupi_n_1569);
  or csa_tree_add_7_27_groupi_g5557__3680(csa_tree_add_7_27_groupi_n_1630 ,csa_tree_add_7_27_groupi_n_1076 ,csa_tree_add_7_27_groupi_n_1591);
  and csa_tree_add_7_27_groupi_g5558__1617(csa_tree_add_7_27_groupi_n_1629 ,csa_tree_add_7_27_groupi_n_1598 ,csa_tree_add_7_27_groupi_n_1571);
  or csa_tree_add_7_27_groupi_g5559__2802(csa_tree_add_7_27_groupi_n_1628 ,csa_tree_add_7_27_groupi_n_1598 ,csa_tree_add_7_27_groupi_n_1571);
  or csa_tree_add_7_27_groupi_g5560__1705(csa_tree_add_7_27_groupi_n_1627 ,csa_tree_add_7_27_groupi_n_1107 ,csa_tree_add_7_27_groupi_n_1592);
  and csa_tree_add_7_27_groupi_g5561__5122(csa_tree_add_7_27_groupi_n_1640 ,csa_tree_add_7_27_groupi_n_770 ,csa_tree_add_7_27_groupi_n_1610);
  or csa_tree_add_7_27_groupi_g5562__8246(csa_tree_add_7_27_groupi_n_1639 ,csa_tree_add_7_27_groupi_n_1523 ,csa_tree_add_7_27_groupi_n_1609);
  or csa_tree_add_7_27_groupi_g5563__7098(csa_tree_add_7_27_groupi_n_1638 ,csa_tree_add_7_27_groupi_n_1519 ,csa_tree_add_7_27_groupi_n_1611);
  or csa_tree_add_7_27_groupi_g5564__6131(csa_tree_add_7_27_groupi_n_1637 ,csa_tree_add_7_27_groupi_n_1525 ,csa_tree_add_7_27_groupi_n_1608);
  or csa_tree_add_7_27_groupi_g5565__1881(csa_tree_add_7_27_groupi_n_1619 ,csa_tree_add_7_27_groupi_n_1596 ,csa_tree_add_7_27_groupi_n_1569);
  xnor csa_tree_add_7_27_groupi_g5566__5115(n_5 ,csa_tree_add_7_27_groupi_n_1582 ,csa_tree_add_7_27_groupi_n_1534);
  or csa_tree_add_7_27_groupi_g5567__7482(csa_tree_add_7_27_groupi_n_1617 ,csa_tree_add_7_27_groupi_n_1201 ,csa_tree_add_7_27_groupi_n_1594);
  and csa_tree_add_7_27_groupi_g5568__4733(csa_tree_add_7_27_groupi_n_1616 ,csa_tree_add_7_27_groupi_n_3 ,csa_tree_add_7_27_groupi_n_1595);
  or csa_tree_add_7_27_groupi_g5569__6161(csa_tree_add_7_27_groupi_n_1615 ,csa_tree_add_7_27_groupi_n_3 ,csa_tree_add_7_27_groupi_n_1595);
  or csa_tree_add_7_27_groupi_g5570__9315(csa_tree_add_7_27_groupi_n_1614 ,csa_tree_add_7_27_groupi_n_1033 ,csa_tree_add_7_27_groupi_n_1590);
  xnor csa_tree_add_7_27_groupi_g5571__9945(csa_tree_add_7_27_groupi_n_1613 ,csa_tree_add_7_27_groupi_n_1541 ,csa_tree_add_7_27_groupi_n_1567);
  or csa_tree_add_7_27_groupi_g5572__2883(csa_tree_add_7_27_groupi_n_1626 ,csa_tree_add_7_27_groupi_n_1521 ,csa_tree_add_7_27_groupi_n_1612);
  or csa_tree_add_7_27_groupi_g5573__2346(csa_tree_add_7_27_groupi_n_1625 ,csa_tree_add_7_27_groupi_n_1522 ,csa_tree_add_7_27_groupi_n_1607);
  xnor csa_tree_add_7_27_groupi_g5574__1666(csa_tree_add_7_27_groupi_n_1624 ,csa_tree_add_7_27_groupi_n_1583 ,csa_tree_add_7_27_groupi_n_1533);
  xnor csa_tree_add_7_27_groupi_g5575__7410(csa_tree_add_7_27_groupi_n_1623 ,csa_tree_add_7_27_groupi_n_1581 ,csa_tree_add_7_27_groupi_n_1530);
  xnor csa_tree_add_7_27_groupi_g5576__6417(csa_tree_add_7_27_groupi_n_1622 ,csa_tree_add_7_27_groupi_n_1572 ,csa_tree_add_7_27_groupi_n_1531);
  xnor csa_tree_add_7_27_groupi_g5577__5477(csa_tree_add_7_27_groupi_n_1621 ,csa_tree_add_7_27_groupi_n_1585 ,csa_tree_add_7_27_groupi_n_1532);
  xnor csa_tree_add_7_27_groupi_g5578__2398(csa_tree_add_7_27_groupi_n_1620 ,csa_tree_add_7_27_groupi_n_1584 ,csa_tree_add_7_27_groupi_n_832);
  and csa_tree_add_7_27_groupi_g5579__5107(csa_tree_add_7_27_groupi_n_1612 ,csa_tree_add_7_27_groupi_n_1526 ,csa_tree_add_7_27_groupi_n_1572);
  and csa_tree_add_7_27_groupi_g5580__6260(csa_tree_add_7_27_groupi_n_1611 ,csa_tree_add_7_27_groupi_n_1518 ,csa_tree_add_7_27_groupi_n_1585);
  or csa_tree_add_7_27_groupi_g5581__4319(csa_tree_add_7_27_groupi_n_1610 ,csa_tree_add_7_27_groupi_n_769 ,csa_tree_add_7_27_groupi_n_1584);
  and csa_tree_add_7_27_groupi_g5582__8428(csa_tree_add_7_27_groupi_n_1609 ,csa_tree_add_7_27_groupi_n_1517 ,csa_tree_add_7_27_groupi_n_1581);
  and csa_tree_add_7_27_groupi_g5583__5526(csa_tree_add_7_27_groupi_n_1608 ,csa_tree_add_7_27_groupi_n_1524 ,csa_tree_add_7_27_groupi_n_1583);
  and csa_tree_add_7_27_groupi_g5584__6783(csa_tree_add_7_27_groupi_n_1607 ,csa_tree_add_7_27_groupi_n_1516 ,csa_tree_add_7_27_groupi_n_1582);
  or csa_tree_add_7_27_groupi_g5585__3680(csa_tree_add_7_27_groupi_n_1606 ,csa_tree_add_7_27_groupi_n_1541 ,csa_tree_add_7_27_groupi_n_1567);
  and csa_tree_add_7_27_groupi_g5586__1617(csa_tree_add_7_27_groupi_n_1605 ,csa_tree_add_7_27_groupi_n_1541 ,csa_tree_add_7_27_groupi_n_1567);
  nor csa_tree_add_7_27_groupi_g5587__2802(csa_tree_add_7_27_groupi_n_1604 ,csa_tree_add_7_27_groupi_n_1289 ,csa_tree_add_7_27_groupi_n_1565);
  nor csa_tree_add_7_27_groupi_g5588__1705(csa_tree_add_7_27_groupi_n_1603 ,csa_tree_add_7_27_groupi_n_1128 ,csa_tree_add_7_27_groupi_n_1561);
  nor csa_tree_add_7_27_groupi_g5589__5122(csa_tree_add_7_27_groupi_n_1602 ,csa_tree_add_7_27_groupi_n_1271 ,csa_tree_add_7_27_groupi_n_1564);
  nor csa_tree_add_7_27_groupi_g5590__8246(csa_tree_add_7_27_groupi_n_1601 ,csa_tree_add_7_27_groupi_n_1338 ,csa_tree_add_7_27_groupi_n_1577);
  nor csa_tree_add_7_27_groupi_g5591__7098(csa_tree_add_7_27_groupi_n_1600 ,csa_tree_add_7_27_groupi_n_1362 ,csa_tree_add_7_27_groupi_n_1580);
  nor csa_tree_add_7_27_groupi_g5592__6131(csa_tree_add_7_27_groupi_n_1594 ,csa_tree_add_7_27_groupi_n_455 ,csa_tree_add_7_27_groupi_n_552);
  nor csa_tree_add_7_27_groupi_g5593__1881(csa_tree_add_7_27_groupi_n_1593 ,csa_tree_add_7_27_groupi_n_467 ,csa_tree_add_7_27_groupi_n_1566);
  nor csa_tree_add_7_27_groupi_g5594__5115(csa_tree_add_7_27_groupi_n_1592 ,csa_tree_add_7_27_groupi_n_464 ,csa_tree_add_7_27_groupi_n_552);
  nor csa_tree_add_7_27_groupi_g5595__7482(csa_tree_add_7_27_groupi_n_1591 ,csa_tree_add_7_27_groupi_n_458 ,csa_tree_add_7_27_groupi_n_1566);
  nor csa_tree_add_7_27_groupi_g5596__4733(csa_tree_add_7_27_groupi_n_1590 ,csa_tree_add_7_27_groupi_n_461 ,csa_tree_add_7_27_groupi_n_551);
  xnor csa_tree_add_7_27_groupi_g5597__6161(csa_tree_add_7_27_groupi_n_1589 ,csa_tree_add_7_27_groupi_n_2 ,csa_tree_add_7_27_groupi_n_1542);
  xnor csa_tree_add_7_27_groupi_g5598__9315(csa_tree_add_7_27_groupi_n_1588 ,csa_tree_add_7_27_groupi_n_1539 ,csa_tree_add_7_27_groupi_n_1544);
  xnor csa_tree_add_7_27_groupi_g5599__9945(csa_tree_add_7_27_groupi_n_1587 ,csa_tree_add_7_27_groupi_n_1540 ,csa_tree_add_7_27_groupi_n_1537);
  xnor csa_tree_add_7_27_groupi_g5600__2883(csa_tree_add_7_27_groupi_n_1586 ,csa_tree_add_7_27_groupi_n_1538 ,csa_tree_add_7_27_groupi_n_1543);
  xnor csa_tree_add_7_27_groupi_g5601__2346(csa_tree_add_7_27_groupi_n_1599 ,csa_tree_add_7_27_groupi_n_1547 ,in2[11]);
  xnor csa_tree_add_7_27_groupi_g5602__1666(csa_tree_add_7_27_groupi_n_1598 ,csa_tree_add_7_27_groupi_n_1545 ,in2[8]);
  xnor csa_tree_add_7_27_groupi_g5603__7410(csa_tree_add_7_27_groupi_n_1597 ,csa_tree_add_7_27_groupi_n_1546 ,in2[5]);
  xnor csa_tree_add_7_27_groupi_g5604__6417(csa_tree_add_7_27_groupi_n_1596 ,csa_tree_add_7_27_groupi_n_1549 ,in2[2]);
  xnor csa_tree_add_7_27_groupi_g5605__5477(csa_tree_add_7_27_groupi_n_1595 ,csa_tree_add_7_27_groupi_n_1548 ,in2[14]);
  or csa_tree_add_7_27_groupi_g5606__2398(csa_tree_add_7_27_groupi_n_1580 ,csa_tree_add_7_27_groupi_n_1120 ,csa_tree_add_7_27_groupi_n_1535);
  and csa_tree_add_7_27_groupi_g5607__5107(csa_tree_add_7_27_groupi_n_1579 ,csa_tree_add_7_27_groupi_n_1540 ,csa_tree_add_7_27_groupi_n_1537);
  or csa_tree_add_7_27_groupi_g5608__6260(csa_tree_add_7_27_groupi_n_1578 ,csa_tree_add_7_27_groupi_n_1540 ,csa_tree_add_7_27_groupi_n_1537);
  or csa_tree_add_7_27_groupi_g5609__4319(csa_tree_add_7_27_groupi_n_1577 ,csa_tree_add_7_27_groupi_n_1104 ,csa_tree_add_7_27_groupi_n_1552);
  and csa_tree_add_7_27_groupi_g5610__8428(csa_tree_add_7_27_groupi_n_1576 ,csa_tree_add_7_27_groupi_n_1539 ,csa_tree_add_7_27_groupi_n_1544);
  or csa_tree_add_7_27_groupi_g5611__5526(csa_tree_add_7_27_groupi_n_1575 ,csa_tree_add_7_27_groupi_n_1539 ,csa_tree_add_7_27_groupi_n_1544);
  and csa_tree_add_7_27_groupi_g5612__6783(csa_tree_add_7_27_groupi_n_1574 ,csa_tree_add_7_27_groupi_n_2 ,csa_tree_add_7_27_groupi_n_1542);
  or csa_tree_add_7_27_groupi_g5613__3680(csa_tree_add_7_27_groupi_n_1573 ,csa_tree_add_7_27_groupi_n_2 ,csa_tree_add_7_27_groupi_n_1542);
  or csa_tree_add_7_27_groupi_g5614__1617(csa_tree_add_7_27_groupi_n_1585 ,csa_tree_add_7_27_groupi_n_1491 ,csa_tree_add_7_27_groupi_n_1557);
  and csa_tree_add_7_27_groupi_g5615__2802(csa_tree_add_7_27_groupi_n_1584 ,csa_tree_add_7_27_groupi_n_779 ,csa_tree_add_7_27_groupi_n_1556);
  or csa_tree_add_7_27_groupi_g5616__1705(csa_tree_add_7_27_groupi_n_1583 ,csa_tree_add_7_27_groupi_n_1498 ,csa_tree_add_7_27_groupi_n_1559);
  or csa_tree_add_7_27_groupi_g5617__5122(csa_tree_add_7_27_groupi_n_1582 ,csa_tree_add_7_27_groupi_n_1495 ,csa_tree_add_7_27_groupi_n_1558);
  or csa_tree_add_7_27_groupi_g5618__8246(csa_tree_add_7_27_groupi_n_1581 ,csa_tree_add_7_27_groupi_n_1478 ,csa_tree_add_7_27_groupi_n_1554);
  or csa_tree_add_7_27_groupi_g5619__7098(csa_tree_add_7_27_groupi_n_1565 ,csa_tree_add_7_27_groupi_n_1235 ,csa_tree_add_7_27_groupi_n_1551);
  or csa_tree_add_7_27_groupi_g5620__6131(csa_tree_add_7_27_groupi_n_1564 ,csa_tree_add_7_27_groupi_n_1207 ,csa_tree_add_7_27_groupi_n_1550);
  or csa_tree_add_7_27_groupi_g5621__1881(csa_tree_add_7_27_groupi_n_1563 ,csa_tree_add_7_27_groupi_n_1538 ,csa_tree_add_7_27_groupi_n_1543);
  and csa_tree_add_7_27_groupi_g5622__5115(csa_tree_add_7_27_groupi_n_1562 ,csa_tree_add_7_27_groupi_n_1538 ,csa_tree_add_7_27_groupi_n_1543);
  or csa_tree_add_7_27_groupi_g5623__7482(csa_tree_add_7_27_groupi_n_1561 ,csa_tree_add_7_27_groupi_n_1029 ,csa_tree_add_7_27_groupi_n_1553);
  xnor csa_tree_add_7_27_groupi_g5624__4733(n_4 ,csa_tree_add_7_27_groupi_n_1515 ,csa_tree_add_7_27_groupi_n_1502);
  or csa_tree_add_7_27_groupi_g5625__6161(csa_tree_add_7_27_groupi_n_1572 ,csa_tree_add_7_27_groupi_n_1487 ,csa_tree_add_7_27_groupi_n_1555);
  xnor csa_tree_add_7_27_groupi_g5626__9315(csa_tree_add_7_27_groupi_n_1571 ,csa_tree_add_7_27_groupi_n_1527 ,csa_tree_add_7_27_groupi_n_1505);
  xnor csa_tree_add_7_27_groupi_g5627__9945(csa_tree_add_7_27_groupi_n_1570 ,csa_tree_add_7_27_groupi_n_1528 ,csa_tree_add_7_27_groupi_n_1504);
  xnor csa_tree_add_7_27_groupi_g5628__2883(csa_tree_add_7_27_groupi_n_1569 ,csa_tree_add_7_27_groupi_n_1514 ,csa_tree_add_7_27_groupi_n_1503);
  xnor csa_tree_add_7_27_groupi_g5629__2346(csa_tree_add_7_27_groupi_n_1568 ,csa_tree_add_7_27_groupi_n_1513 ,csa_tree_add_7_27_groupi_n_1501);
  xnor csa_tree_add_7_27_groupi_g5630__1666(csa_tree_add_7_27_groupi_n_1567 ,csa_tree_add_7_27_groupi_n_1406 ,csa_tree_add_7_27_groupi_n_1506);
  xnor csa_tree_add_7_27_groupi_g5631__7410(csa_tree_add_7_27_groupi_n_1566 ,csa_tree_add_7_27_groupi_n_1529 ,csa_tree_add_7_27_groupi_n_839);
  and csa_tree_add_7_27_groupi_g5632__6417(csa_tree_add_7_27_groupi_n_1559 ,csa_tree_add_7_27_groupi_n_1497 ,csa_tree_add_7_27_groupi_n_1527);
  and csa_tree_add_7_27_groupi_g5633__5477(csa_tree_add_7_27_groupi_n_1558 ,csa_tree_add_7_27_groupi_n_1493 ,csa_tree_add_7_27_groupi_n_1515);
  and csa_tree_add_7_27_groupi_g5634__2398(csa_tree_add_7_27_groupi_n_1557 ,csa_tree_add_7_27_groupi_n_1490 ,csa_tree_add_7_27_groupi_n_1528);
  or csa_tree_add_7_27_groupi_g5635__5107(csa_tree_add_7_27_groupi_n_1556 ,csa_tree_add_7_27_groupi_n_784 ,csa_tree_add_7_27_groupi_n_1529);
  and csa_tree_add_7_27_groupi_g5636__6260(csa_tree_add_7_27_groupi_n_1555 ,csa_tree_add_7_27_groupi_n_1494 ,csa_tree_add_7_27_groupi_n_1514);
  and csa_tree_add_7_27_groupi_g5637__4319(csa_tree_add_7_27_groupi_n_1554 ,csa_tree_add_7_27_groupi_n_1492 ,csa_tree_add_7_27_groupi_n_1513);
  nor csa_tree_add_7_27_groupi_g5638__8428(csa_tree_add_7_27_groupi_n_1553 ,csa_tree_add_7_27_groupi_n_437 ,csa_tree_add_7_27_groupi_n_546);
  nor csa_tree_add_7_27_groupi_g5639__5526(csa_tree_add_7_27_groupi_n_1552 ,csa_tree_add_7_27_groupi_n_380 ,csa_tree_add_7_27_groupi_n_1512);
  nor csa_tree_add_7_27_groupi_g5640__6783(csa_tree_add_7_27_groupi_n_1551 ,csa_tree_add_7_27_groupi_n_453 ,csa_tree_add_7_27_groupi_n_546);
  nor csa_tree_add_7_27_groupi_g5641__3680(csa_tree_add_7_27_groupi_n_1550 ,csa_tree_add_7_27_groupi_n_407 ,csa_tree_add_7_27_groupi_n_1512);
  nor csa_tree_add_7_27_groupi_g5642__1617(csa_tree_add_7_27_groupi_n_1549 ,csa_tree_add_7_27_groupi_n_1126 ,csa_tree_add_7_27_groupi_n_1510);
  nor csa_tree_add_7_27_groupi_g5643__2802(csa_tree_add_7_27_groupi_n_1548 ,csa_tree_add_7_27_groupi_n_1277 ,csa_tree_add_7_27_groupi_n_1509);
  nor csa_tree_add_7_27_groupi_g5644__1705(csa_tree_add_7_27_groupi_n_1547 ,csa_tree_add_7_27_groupi_n_1285 ,csa_tree_add_7_27_groupi_n_1507);
  nor csa_tree_add_7_27_groupi_g5645__5122(csa_tree_add_7_27_groupi_n_1546 ,csa_tree_add_7_27_groupi_n_1266 ,csa_tree_add_7_27_groupi_n_1508);
  nor csa_tree_add_7_27_groupi_g5646__8246(csa_tree_add_7_27_groupi_n_1545 ,csa_tree_add_7_27_groupi_n_1324 ,csa_tree_add_7_27_groupi_n_1520);
  xnor csa_tree_add_7_27_groupi_g5647__7098(csa_tree_add_7_27_groupi_n_1536 ,csa_tree_add_7_27_groupi_n_1460 ,csa_tree_add_7_27_groupi_n_1470);
  nor csa_tree_add_7_27_groupi_g5648__6131(csa_tree_add_7_27_groupi_n_1535 ,csa_tree_add_7_27_groupi_n_425 ,csa_tree_add_7_27_groupi_n_545);
  xnor csa_tree_add_7_27_groupi_g5649__1881(csa_tree_add_7_27_groupi_n_1534 ,csa_tree_add_7_27_groupi_n_1481 ,csa_tree_add_7_27_groupi_n_1444);
  xnor csa_tree_add_7_27_groupi_g5650__5115(csa_tree_add_7_27_groupi_n_1533 ,csa_tree_add_7_27_groupi_n_1447 ,csa_tree_add_7_27_groupi_n_1480);
  xnor csa_tree_add_7_27_groupi_g5651__7482(csa_tree_add_7_27_groupi_n_1532 ,csa_tree_add_7_27_groupi_n_1446 ,csa_tree_add_7_27_groupi_n_1479);
  xnor csa_tree_add_7_27_groupi_g5652__4733(csa_tree_add_7_27_groupi_n_1531 ,csa_tree_add_7_27_groupi_n_1445 ,csa_tree_add_7_27_groupi_n_1483);
  xnor csa_tree_add_7_27_groupi_g5653__6161(csa_tree_add_7_27_groupi_n_1530 ,csa_tree_add_7_27_groupi_n_1 ,csa_tree_add_7_27_groupi_n_1482);
  xnor csa_tree_add_7_27_groupi_g5654__9315(csa_tree_add_7_27_groupi_n_1544 ,csa_tree_add_7_27_groupi_n_1461 ,csa_tree_add_7_27_groupi_n_1468);
  xnor csa_tree_add_7_27_groupi_g5655__9945(csa_tree_add_7_27_groupi_n_1543 ,csa_tree_add_7_27_groupi_n_1465 ,csa_tree_add_7_27_groupi_n_1469);
  xnor csa_tree_add_7_27_groupi_g5656__2883(csa_tree_add_7_27_groupi_n_1542 ,csa_tree_add_7_27_groupi_n_1466 ,in2[14]);
  xnor csa_tree_add_7_27_groupi_g5657__2346(csa_tree_add_7_27_groupi_n_1541 ,csa_tree_add_7_27_groupi_n_1471 ,in2[2]);
  xnor csa_tree_add_7_27_groupi_g5658__1666(csa_tree_add_7_27_groupi_n_1540 ,csa_tree_add_7_27_groupi_n_1484 ,in2[11]);
  xnor csa_tree_add_7_27_groupi_g5659__7410(csa_tree_add_7_27_groupi_n_1539 ,csa_tree_add_7_27_groupi_n_1485 ,in2[8]);
  xnor csa_tree_add_7_27_groupi_g5660__6417(csa_tree_add_7_27_groupi_n_1538 ,csa_tree_add_7_27_groupi_n_1486 ,in2[5]);
  xnor csa_tree_add_7_27_groupi_g5661__5477(csa_tree_add_7_27_groupi_n_1537 ,csa_tree_add_7_27_groupi_n_1463 ,csa_tree_add_7_27_groupi_n_1467);
  or csa_tree_add_7_27_groupi_g5662__2398(csa_tree_add_7_27_groupi_n_1526 ,csa_tree_add_7_27_groupi_n_1445 ,csa_tree_add_7_27_groupi_n_1483);
  and csa_tree_add_7_27_groupi_g5663__5107(csa_tree_add_7_27_groupi_n_1525 ,csa_tree_add_7_27_groupi_n_1447 ,csa_tree_add_7_27_groupi_n_1480);
  or csa_tree_add_7_27_groupi_g5664__6260(csa_tree_add_7_27_groupi_n_1524 ,csa_tree_add_7_27_groupi_n_1447 ,csa_tree_add_7_27_groupi_n_1480);
  and csa_tree_add_7_27_groupi_g5665__4319(csa_tree_add_7_27_groupi_n_1523 ,csa_tree_add_7_27_groupi_n_1 ,csa_tree_add_7_27_groupi_n_1482);
  and csa_tree_add_7_27_groupi_g5666__8428(csa_tree_add_7_27_groupi_n_1522 ,csa_tree_add_7_27_groupi_n_1481 ,csa_tree_add_7_27_groupi_n_1444);
  and csa_tree_add_7_27_groupi_g5667__5526(csa_tree_add_7_27_groupi_n_1521 ,csa_tree_add_7_27_groupi_n_1445 ,csa_tree_add_7_27_groupi_n_1483);
  or csa_tree_add_7_27_groupi_g5668__6783(csa_tree_add_7_27_groupi_n_1520 ,csa_tree_add_7_27_groupi_n_1122 ,csa_tree_add_7_27_groupi_n_1472);
  and csa_tree_add_7_27_groupi_g5669__3680(csa_tree_add_7_27_groupi_n_1519 ,csa_tree_add_7_27_groupi_n_1446 ,csa_tree_add_7_27_groupi_n_1479);
  or csa_tree_add_7_27_groupi_g5670__1617(csa_tree_add_7_27_groupi_n_1518 ,csa_tree_add_7_27_groupi_n_1446 ,csa_tree_add_7_27_groupi_n_1479);
  or csa_tree_add_7_27_groupi_g5671__2802(csa_tree_add_7_27_groupi_n_1517 ,csa_tree_add_7_27_groupi_n_1 ,csa_tree_add_7_27_groupi_n_1482);
  or csa_tree_add_7_27_groupi_g5672__1705(csa_tree_add_7_27_groupi_n_1516 ,csa_tree_add_7_27_groupi_n_1481 ,csa_tree_add_7_27_groupi_n_1444);
  and csa_tree_add_7_27_groupi_g5673__5122(csa_tree_add_7_27_groupi_n_1529 ,csa_tree_add_7_27_groupi_n_778 ,csa_tree_add_7_27_groupi_n_1488);
  or csa_tree_add_7_27_groupi_g5674__8246(csa_tree_add_7_27_groupi_n_1528 ,csa_tree_add_7_27_groupi_n_1457 ,csa_tree_add_7_27_groupi_n_1489);
  or csa_tree_add_7_27_groupi_g5675__7098(csa_tree_add_7_27_groupi_n_1527 ,csa_tree_add_7_27_groupi_n_1449 ,csa_tree_add_7_27_groupi_n_1496);
  xnor csa_tree_add_7_27_groupi_g5676__6131(csa_tree_add_7_27_groupi_n_1511 ,csa_tree_add_7_27_groupi_n_1430 ,in3[0]);
  or csa_tree_add_7_27_groupi_g5677__1881(csa_tree_add_7_27_groupi_n_1510 ,csa_tree_add_7_27_groupi_n_1001 ,csa_tree_add_7_27_groupi_n_1475);
  or csa_tree_add_7_27_groupi_g5678__5115(csa_tree_add_7_27_groupi_n_1509 ,csa_tree_add_7_27_groupi_n_1246 ,csa_tree_add_7_27_groupi_n_1476);
  or csa_tree_add_7_27_groupi_g5679__7482(csa_tree_add_7_27_groupi_n_1508 ,csa_tree_add_7_27_groupi_n_1206 ,csa_tree_add_7_27_groupi_n_1474);
  or csa_tree_add_7_27_groupi_g5680__4733(csa_tree_add_7_27_groupi_n_1507 ,csa_tree_add_7_27_groupi_n_1198 ,csa_tree_add_7_27_groupi_n_1473);
  xnor csa_tree_add_7_27_groupi_g5681__6161(csa_tree_add_7_27_groupi_n_1506 ,csa_tree_add_7_27_groupi_n_1464 ,in3[4]);
  xnor csa_tree_add_7_27_groupi_g5682__9315(csa_tree_add_7_27_groupi_n_1505 ,csa_tree_add_7_27_groupi_n_1441 ,in3[11]);
  xnor csa_tree_add_7_27_groupi_g5683__9945(csa_tree_add_7_27_groupi_n_1504 ,csa_tree_add_7_27_groupi_n_1440 ,in3[8]);
  xnor csa_tree_add_7_27_groupi_g5684__2883(csa_tree_add_7_27_groupi_n_1503 ,csa_tree_add_7_27_groupi_n_1439 ,in3[5]);
  xnor csa_tree_add_7_27_groupi_g5685__2346(csa_tree_add_7_27_groupi_n_1502 ,csa_tree_add_7_27_groupi_n_1442 ,in3[2]);
  xnor csa_tree_add_7_27_groupi_g5686__1666(csa_tree_add_7_27_groupi_n_1501 ,csa_tree_add_7_27_groupi_n_1443 ,in3[14]);
  or csa_tree_add_7_27_groupi_g5687__7410(csa_tree_add_7_27_groupi_n_1515 ,csa_tree_add_7_27_groupi_n_1458 ,csa_tree_add_7_27_groupi_n_1477);
  or csa_tree_add_7_27_groupi_g5688__6417(csa_tree_add_7_27_groupi_n_1514 ,csa_tree_add_7_27_groupi_n_1455 ,csa_tree_add_7_27_groupi_n_1499);
  or csa_tree_add_7_27_groupi_g5689__5477(csa_tree_add_7_27_groupi_n_1513 ,csa_tree_add_7_27_groupi_n_1451 ,csa_tree_add_7_27_groupi_n_1500);
  xnor csa_tree_add_7_27_groupi_g5690__2398(csa_tree_add_7_27_groupi_n_1512 ,csa_tree_add_7_27_groupi_n_1462 ,csa_tree_add_7_27_groupi_n_846);
  and csa_tree_add_7_27_groupi_g5691__5107(csa_tree_add_7_27_groupi_n_1500 ,csa_tree_add_7_27_groupi_n_1463 ,csa_tree_add_7_27_groupi_n_1452);
  and csa_tree_add_7_27_groupi_g5692__6260(csa_tree_add_7_27_groupi_n_1499 ,csa_tree_add_7_27_groupi_n_1464 ,csa_tree_add_7_27_groupi_n_1454);
  and csa_tree_add_7_27_groupi_g5693__4319(csa_tree_add_7_27_groupi_n_1498 ,in3[11] ,csa_tree_add_7_27_groupi_n_1441);
  or csa_tree_add_7_27_groupi_g5694__8428(csa_tree_add_7_27_groupi_n_1497 ,in3[11] ,csa_tree_add_7_27_groupi_n_1441);
  and csa_tree_add_7_27_groupi_g5695__5526(csa_tree_add_7_27_groupi_n_1496 ,csa_tree_add_7_27_groupi_n_1461 ,csa_tree_add_7_27_groupi_n_1459);
  and csa_tree_add_7_27_groupi_g5696__6783(csa_tree_add_7_27_groupi_n_1495 ,in3[2] ,csa_tree_add_7_27_groupi_n_1442);
  or csa_tree_add_7_27_groupi_g5697__3680(csa_tree_add_7_27_groupi_n_1494 ,in3[5] ,csa_tree_add_7_27_groupi_n_1439);
  or csa_tree_add_7_27_groupi_g5698__1617(csa_tree_add_7_27_groupi_n_1493 ,in3[2] ,csa_tree_add_7_27_groupi_n_1442);
  or csa_tree_add_7_27_groupi_g5699__2802(csa_tree_add_7_27_groupi_n_1492 ,in3[14] ,csa_tree_add_7_27_groupi_n_1443);
  and csa_tree_add_7_27_groupi_g5700__1705(csa_tree_add_7_27_groupi_n_1491 ,in3[8] ,csa_tree_add_7_27_groupi_n_1440);
  or csa_tree_add_7_27_groupi_g5701__5122(csa_tree_add_7_27_groupi_n_1490 ,in3[8] ,csa_tree_add_7_27_groupi_n_1440);
  and csa_tree_add_7_27_groupi_g5702__8246(csa_tree_add_7_27_groupi_n_1489 ,csa_tree_add_7_27_groupi_n_1465 ,csa_tree_add_7_27_groupi_n_1456);
  or csa_tree_add_7_27_groupi_g5703__7098(csa_tree_add_7_27_groupi_n_1488 ,csa_tree_add_7_27_groupi_n_762 ,csa_tree_add_7_27_groupi_n_1462);
  and csa_tree_add_7_27_groupi_g5704__6131(csa_tree_add_7_27_groupi_n_1487 ,in3[5] ,csa_tree_add_7_27_groupi_n_1439);
  nor csa_tree_add_7_27_groupi_g5705__1881(csa_tree_add_7_27_groupi_n_1486 ,csa_tree_add_7_27_groupi_n_1339 ,csa_tree_add_7_27_groupi_n_1453);
  nor csa_tree_add_7_27_groupi_g5706__5115(csa_tree_add_7_27_groupi_n_1485 ,csa_tree_add_7_27_groupi_n_1357 ,csa_tree_add_7_27_groupi_n_1448);
  nor csa_tree_add_7_27_groupi_g5707__7482(csa_tree_add_7_27_groupi_n_1484 ,csa_tree_add_7_27_groupi_n_1292 ,csa_tree_add_7_27_groupi_n_1436);
  and csa_tree_add_7_27_groupi_g5708__4733(csa_tree_add_7_27_groupi_n_1478 ,in3[14] ,csa_tree_add_7_27_groupi_n_1443);
  and csa_tree_add_7_27_groupi_g5709__6161(csa_tree_add_7_27_groupi_n_1477 ,csa_tree_add_7_27_groupi_n_1460 ,csa_tree_add_7_27_groupi_n_1450);
  nor csa_tree_add_7_27_groupi_g5710__9315(csa_tree_add_7_27_groupi_n_1476 ,csa_tree_add_7_27_groupi_n_316 ,csa_tree_add_7_27_groupi_n_524);
  nor csa_tree_add_7_27_groupi_g5711__9945(csa_tree_add_7_27_groupi_n_1475 ,csa_tree_add_7_27_groupi_n_304 ,csa_tree_add_7_27_groupi_n_1438);
  nor csa_tree_add_7_27_groupi_g5712__2883(csa_tree_add_7_27_groupi_n_1474 ,csa_tree_add_7_27_groupi_n_268 ,csa_tree_add_7_27_groupi_n_524);
  nor csa_tree_add_7_27_groupi_g5713__2346(csa_tree_add_7_27_groupi_n_1473 ,csa_tree_add_7_27_groupi_n_343 ,csa_tree_add_7_27_groupi_n_1438);
  nor csa_tree_add_7_27_groupi_g5714__1666(csa_tree_add_7_27_groupi_n_1472 ,csa_tree_add_7_27_groupi_n_283 ,csa_tree_add_7_27_groupi_n_523);
  nor csa_tree_add_7_27_groupi_g5715__7410(csa_tree_add_7_27_groupi_n_1471 ,csa_tree_add_7_27_groupi_n_1129 ,csa_tree_add_7_27_groupi_n_1437);
  xnor csa_tree_add_7_27_groupi_g5716__6417(csa_tree_add_7_27_groupi_n_1470 ,csa_tree_add_7_27_groupi_n_1404 ,in3[1]);
  xnor csa_tree_add_7_27_groupi_g5717__5477(csa_tree_add_7_27_groupi_n_1469 ,csa_tree_add_7_27_groupi_n_1405 ,in3[7]);
  xnor csa_tree_add_7_27_groupi_g5718__2398(csa_tree_add_7_27_groupi_n_1468 ,csa_tree_add_7_27_groupi_n_1403 ,in3[10]);
  xnor csa_tree_add_7_27_groupi_g5719__5107(csa_tree_add_7_27_groupi_n_1467 ,csa_tree_add_7_27_groupi_n_1413 ,in3[13]);
  nor csa_tree_add_7_27_groupi_g5720__6260(csa_tree_add_7_27_groupi_n_1466 ,csa_tree_add_7_27_groupi_n_1270 ,csa_tree_add_7_27_groupi_n_1435);
  xnor csa_tree_add_7_27_groupi_g5721__4319(csa_tree_add_7_27_groupi_n_1483 ,csa_tree_add_7_27_groupi_n_1417 ,in2[5]);
  xnor csa_tree_add_7_27_groupi_g5722__8428(csa_tree_add_7_27_groupi_n_1482 ,csa_tree_add_7_27_groupi_n_1415 ,in2[14]);
  xnor csa_tree_add_7_27_groupi_g5723__5526(csa_tree_add_7_27_groupi_n_1481 ,csa_tree_add_7_27_groupi_n_1416 ,in2[2]);
  xnor csa_tree_add_7_27_groupi_g5724__6783(csa_tree_add_7_27_groupi_n_1480 ,csa_tree_add_7_27_groupi_n_1414 ,in2[11]);
  xnor csa_tree_add_7_27_groupi_g5725__3680(csa_tree_add_7_27_groupi_n_1479 ,csa_tree_add_7_27_groupi_n_1418 ,in2[8]);
  or csa_tree_add_7_27_groupi_g5726__1617(csa_tree_add_7_27_groupi_n_1459 ,in3[10] ,csa_tree_add_7_27_groupi_n_1403);
  and csa_tree_add_7_27_groupi_g5727__2802(csa_tree_add_7_27_groupi_n_1458 ,in3[1] ,csa_tree_add_7_27_groupi_n_1404);
  and csa_tree_add_7_27_groupi_g5728__1705(csa_tree_add_7_27_groupi_n_1457 ,in3[7] ,csa_tree_add_7_27_groupi_n_1405);
  or csa_tree_add_7_27_groupi_g5729__5122(csa_tree_add_7_27_groupi_n_1456 ,in3[7] ,csa_tree_add_7_27_groupi_n_1405);
  and csa_tree_add_7_27_groupi_g5730__8246(csa_tree_add_7_27_groupi_n_1455 ,in3[4] ,csa_tree_add_7_27_groupi_n_1406);
  or csa_tree_add_7_27_groupi_g5731__7098(csa_tree_add_7_27_groupi_n_1454 ,in3[4] ,csa_tree_add_7_27_groupi_n_1406);
  or csa_tree_add_7_27_groupi_g5732__6131(csa_tree_add_7_27_groupi_n_1453 ,csa_tree_add_7_27_groupi_n_1036 ,csa_tree_add_7_27_groupi_n_1399);
  or csa_tree_add_7_27_groupi_g5733__1881(csa_tree_add_7_27_groupi_n_1452 ,in3[13] ,csa_tree_add_7_27_groupi_n_1413);
  and csa_tree_add_7_27_groupi_g5734__5115(csa_tree_add_7_27_groupi_n_1451 ,in3[13] ,csa_tree_add_7_27_groupi_n_1413);
  or csa_tree_add_7_27_groupi_g5735__7482(csa_tree_add_7_27_groupi_n_1450 ,in3[1] ,csa_tree_add_7_27_groupi_n_1404);
  and csa_tree_add_7_27_groupi_g5736__4733(csa_tree_add_7_27_groupi_n_1449 ,in3[10] ,csa_tree_add_7_27_groupi_n_1403);
  or csa_tree_add_7_27_groupi_g5737__6161(csa_tree_add_7_27_groupi_n_1448 ,csa_tree_add_7_27_groupi_n_1014 ,csa_tree_add_7_27_groupi_n_1397);
  or csa_tree_add_7_27_groupi_g5738__9315(csa_tree_add_7_27_groupi_n_1465 ,csa_tree_add_7_27_groupi_n_765 ,csa_tree_add_7_27_groupi_n_1425);
  or csa_tree_add_7_27_groupi_g5739__9945(csa_tree_add_7_27_groupi_n_1464 ,csa_tree_add_7_27_groupi_n_801 ,csa_tree_add_7_27_groupi_n_1422);
  or csa_tree_add_7_27_groupi_g5740__2883(csa_tree_add_7_27_groupi_n_1463 ,csa_tree_add_7_27_groupi_n_763 ,csa_tree_add_7_27_groupi_n_1420);
  and csa_tree_add_7_27_groupi_g5741__2346(csa_tree_add_7_27_groupi_n_1462 ,csa_tree_add_7_27_groupi_n_776 ,csa_tree_add_7_27_groupi_n_1421);
  or csa_tree_add_7_27_groupi_g5742__1666(csa_tree_add_7_27_groupi_n_1461 ,csa_tree_add_7_27_groupi_n_761 ,csa_tree_add_7_27_groupi_n_1427);
  or csa_tree_add_7_27_groupi_g5743__7410(csa_tree_add_7_27_groupi_n_1460 ,csa_tree_add_7_27_groupi_n_774 ,csa_tree_add_7_27_groupi_n_1419);
  or csa_tree_add_7_27_groupi_g5744__6417(csa_tree_add_7_27_groupi_n_1437 ,csa_tree_add_7_27_groupi_n_1027 ,csa_tree_add_7_27_groupi_n_1400);
  or csa_tree_add_7_27_groupi_g5745__5477(csa_tree_add_7_27_groupi_n_1436 ,csa_tree_add_7_27_groupi_n_1247 ,csa_tree_add_7_27_groupi_n_1398);
  or csa_tree_add_7_27_groupi_g5746__2398(csa_tree_add_7_27_groupi_n_1435 ,csa_tree_add_7_27_groupi_n_1217 ,csa_tree_add_7_27_groupi_n_1396);
  xnor csa_tree_add_7_27_groupi_g5747__5107(csa_tree_add_7_27_groupi_n_1434 ,csa_tree_add_7_27_groupi_n_1392 ,csa_tree_add_7_27_groupi_n_669);
  xnor csa_tree_add_7_27_groupi_g5748__6260(csa_tree_add_7_27_groupi_n_1433 ,csa_tree_add_7_27_groupi_n_1393 ,csa_tree_add_7_27_groupi_n_671);
  xnor csa_tree_add_7_27_groupi_g5749__4319(csa_tree_add_7_27_groupi_n_1432 ,csa_tree_add_7_27_groupi_n_1391 ,csa_tree_add_7_27_groupi_n_1155);
  xnor csa_tree_add_7_27_groupi_g5750__8428(csa_tree_add_7_27_groupi_n_1431 ,csa_tree_add_7_27_groupi_n_873 ,csa_tree_add_7_27_groupi_n_1383);
  xnor csa_tree_add_7_27_groupi_g5751__5526(csa_tree_add_7_27_groupi_n_1430 ,csa_tree_add_7_27_groupi_n_1381 ,in2[2]);
  xnor csa_tree_add_7_27_groupi_g5752__6783(csa_tree_add_7_27_groupi_n_1447 ,csa_tree_add_7_27_groupi_n_1380 ,csa_tree_add_7_27_groupi_n_842);
  xnor csa_tree_add_7_27_groupi_g5753__3680(csa_tree_add_7_27_groupi_n_1446 ,csa_tree_add_7_27_groupi_n_1377 ,csa_tree_add_7_27_groupi_n_844);
  xnor csa_tree_add_7_27_groupi_g5754__1617(csa_tree_add_7_27_groupi_n_1445 ,csa_tree_add_7_27_groupi_n_1379 ,csa_tree_add_7_27_groupi_n_845);
  xnor csa_tree_add_7_27_groupi_g5755__2802(csa_tree_add_7_27_groupi_n_1444 ,csa_tree_add_7_27_groupi_n_1378 ,csa_tree_add_7_27_groupi_n_843);
  xnor csa_tree_add_7_27_groupi_g5756__1705(csa_tree_add_7_27_groupi_n_1443 ,csa_tree_add_7_27_groupi_n_1370 ,in2[14]);
  xnor csa_tree_add_7_27_groupi_g5757__5122(csa_tree_add_7_27_groupi_n_1442 ,csa_tree_add_7_27_groupi_n_1371 ,in2[2]);
  xnor csa_tree_add_7_27_groupi_g5758__8246(csa_tree_add_7_27_groupi_n_1441 ,csa_tree_add_7_27_groupi_n_1382 ,in2[11]);
  xnor csa_tree_add_7_27_groupi_g5759__7098(csa_tree_add_7_27_groupi_n_1440 ,csa_tree_add_7_27_groupi_n_1385 ,in2[8]);
  xnor csa_tree_add_7_27_groupi_g5760__6131(csa_tree_add_7_27_groupi_n_1439 ,csa_tree_add_7_27_groupi_n_1384 ,in2[5]);
  xnor csa_tree_add_7_27_groupi_g5761__1881(csa_tree_add_7_27_groupi_n_1438 ,csa_tree_add_7_27_groupi_n_1376 ,csa_tree_add_7_27_groupi_n_831);
  and csa_tree_add_7_27_groupi_g5762__5115(csa_tree_add_7_27_groupi_n_1429 ,csa_tree_add_7_27_groupi_n_659 ,csa_tree_add_7_27_groupi_n_1393);
  or csa_tree_add_7_27_groupi_g5763__7482(csa_tree_add_7_27_groupi_n_1428 ,csa_tree_add_7_27_groupi_n_657 ,csa_tree_add_7_27_groupi_n_1392);
  and csa_tree_add_7_27_groupi_g5764__4733(csa_tree_add_7_27_groupi_n_1427 ,csa_tree_add_7_27_groupi_n_786 ,csa_tree_add_7_27_groupi_n_1377);
  or csa_tree_add_7_27_groupi_g5765__6161(csa_tree_add_7_27_groupi_n_1426 ,csa_tree_add_7_27_groupi_n_488 ,csa_tree_add_7_27_groupi_n_1391);
  and csa_tree_add_7_27_groupi_g5766__9315(csa_tree_add_7_27_groupi_n_1425 ,csa_tree_add_7_27_groupi_n_772 ,csa_tree_add_7_27_groupi_n_1379);
  and csa_tree_add_7_27_groupi_g5767__9945(csa_tree_add_7_27_groupi_n_1424 ,csa_tree_add_7_27_groupi_n_657 ,csa_tree_add_7_27_groupi_n_1392);
  and csa_tree_add_7_27_groupi_g5768__2883(csa_tree_add_7_27_groupi_n_1423 ,csa_tree_add_7_27_groupi_n_488 ,csa_tree_add_7_27_groupi_n_1391);
  and csa_tree_add_7_27_groupi_g5769__2346(csa_tree_add_7_27_groupi_n_1422 ,csa_tree_add_7_27_groupi_n_789 ,csa_tree_add_7_27_groupi_n_1378);
  or csa_tree_add_7_27_groupi_g5770__1666(csa_tree_add_7_27_groupi_n_1421 ,csa_tree_add_7_27_groupi_n_771 ,csa_tree_add_7_27_groupi_n_1376);
  and csa_tree_add_7_27_groupi_g5771__7410(csa_tree_add_7_27_groupi_n_1420 ,csa_tree_add_7_27_groupi_n_764 ,csa_tree_add_7_27_groupi_n_1380);
  and csa_tree_add_7_27_groupi_g5772__6417(csa_tree_add_7_27_groupi_n_1419 ,csa_tree_add_7_27_groupi_n_775 ,csa_tree_add_7_27_groupi_n_1381);
  nor csa_tree_add_7_27_groupi_g5773__5477(csa_tree_add_7_27_groupi_n_1418 ,csa_tree_add_7_27_groupi_n_1359 ,csa_tree_add_7_27_groupi_n_1387);
  nor csa_tree_add_7_27_groupi_g5774__2398(csa_tree_add_7_27_groupi_n_1417 ,csa_tree_add_7_27_groupi_n_1325 ,csa_tree_add_7_27_groupi_n_1374);
  nor csa_tree_add_7_27_groupi_g5775__5107(csa_tree_add_7_27_groupi_n_1416 ,csa_tree_add_7_27_groupi_n_1147 ,csa_tree_add_7_27_groupi_n_1373);
  nor csa_tree_add_7_27_groupi_g5776__6260(csa_tree_add_7_27_groupi_n_1415 ,csa_tree_add_7_27_groupi_n_1264 ,csa_tree_add_7_27_groupi_n_1389);
  nor csa_tree_add_7_27_groupi_g5777__4319(csa_tree_add_7_27_groupi_n_1414 ,csa_tree_add_7_27_groupi_n_1265 ,csa_tree_add_7_27_groupi_n_1388);
  not csa_tree_add_7_27_groupi_g5778(csa_tree_add_7_27_groupi_n_1411 ,csa_tree_add_7_27_groupi_n_1412);
  not csa_tree_add_7_27_groupi_g5779(csa_tree_add_7_27_groupi_n_1409 ,csa_tree_add_7_27_groupi_n_1410);
  not csa_tree_add_7_27_groupi_g5780(csa_tree_add_7_27_groupi_n_1407 ,csa_tree_add_7_27_groupi_n_1408);
  not csa_tree_add_7_27_groupi_g5781(csa_tree_add_7_27_groupi_n_1402 ,csa_tree_add_7_27_groupi_n_1401);
  nor csa_tree_add_7_27_groupi_g5782__8428(csa_tree_add_7_27_groupi_n_1400 ,csa_tree_add_7_27_groupi_n_311 ,csa_tree_add_7_27_groupi_n_549);
  nor csa_tree_add_7_27_groupi_g5783__5526(csa_tree_add_7_27_groupi_n_1399 ,csa_tree_add_7_27_groupi_n_356 ,csa_tree_add_7_27_groupi_n_1375);
  nor csa_tree_add_7_27_groupi_g5784__6783(csa_tree_add_7_27_groupi_n_1398 ,csa_tree_add_7_27_groupi_n_329 ,csa_tree_add_7_27_groupi_n_549);
  nor csa_tree_add_7_27_groupi_g5785__3680(csa_tree_add_7_27_groupi_n_1397 ,csa_tree_add_7_27_groupi_n_299 ,csa_tree_add_7_27_groupi_n_1375);
  nor csa_tree_add_7_27_groupi_g5786__1617(csa_tree_add_7_27_groupi_n_1396 ,csa_tree_add_7_27_groupi_n_278 ,csa_tree_add_7_27_groupi_n_548);
  or csa_tree_add_7_27_groupi_g5787__2802(csa_tree_add_7_27_groupi_n_1395 ,csa_tree_add_7_27_groupi_n_659 ,csa_tree_add_7_27_groupi_n_1393);
  xnor csa_tree_add_7_27_groupi_g5788__1705(csa_tree_add_7_27_groupi_n_1394 ,csa_tree_add_7_27_groupi_n_1334 ,csa_tree_add_7_27_groupi_n_1369);
  xnor csa_tree_add_7_27_groupi_g5789__5122(csa_tree_add_7_27_groupi_n_1413 ,csa_tree_add_7_27_groupi_n_1308 ,in2[14]);
  xnor csa_tree_add_7_27_groupi_g5790__8246(csa_tree_add_7_27_groupi_n_1412 ,csa_tree_add_7_27_groupi_n_1303 ,csa_tree_add_7_27_groupi_n_1162);
  xnor csa_tree_add_7_27_groupi_g5791__7098(csa_tree_add_7_27_groupi_n_1410 ,csa_tree_add_7_27_groupi_n_1302 ,csa_tree_add_7_27_groupi_n_1159);
  xnor csa_tree_add_7_27_groupi_g5792__6131(csa_tree_add_7_27_groupi_n_1408 ,csa_tree_add_7_27_groupi_n_1304 ,csa_tree_add_7_27_groupi_n_1156);
  xnor csa_tree_add_7_27_groupi_g5793__1881(csa_tree_add_7_27_groupi_n_1406 ,csa_tree_add_7_27_groupi_n_1335 ,in2[5]);
  xnor csa_tree_add_7_27_groupi_g5794__5115(csa_tree_add_7_27_groupi_n_1405 ,csa_tree_add_7_27_groupi_n_1337 ,in2[8]);
  xnor csa_tree_add_7_27_groupi_g5795__7482(csa_tree_add_7_27_groupi_n_1404 ,csa_tree_add_7_27_groupi_n_1309 ,in2[2]);
  xnor csa_tree_add_7_27_groupi_g5796__4733(csa_tree_add_7_27_groupi_n_1403 ,csa_tree_add_7_27_groupi_n_1336 ,in2[11]);
  xnor csa_tree_add_7_27_groupi_g5797__6161(csa_tree_add_7_27_groupi_n_1401 ,csa_tree_add_7_27_groupi_n_1305 ,csa_tree_add_7_27_groupi_n_721);
  nor csa_tree_add_7_27_groupi_g5798__9315(csa_tree_add_7_27_groupi_n_1390 ,csa_tree_add_7_27_groupi_n_1334 ,csa_tree_add_7_27_groupi_n_1369);
  or csa_tree_add_7_27_groupi_g5799__9945(csa_tree_add_7_27_groupi_n_1389 ,csa_tree_add_7_27_groupi_n_1255 ,csa_tree_add_7_27_groupi_n_1311);
  or csa_tree_add_7_27_groupi_g5800__2883(csa_tree_add_7_27_groupi_n_1388 ,csa_tree_add_7_27_groupi_n_1250 ,csa_tree_add_7_27_groupi_n_1313);
  or csa_tree_add_7_27_groupi_g5801__2346(csa_tree_add_7_27_groupi_n_1387 ,csa_tree_add_7_27_groupi_n_1083 ,csa_tree_add_7_27_groupi_n_1312);
  or csa_tree_add_7_27_groupi_g5802__1666(csa_tree_add_7_27_groupi_n_1386 ,csa_tree_add_7_27_groupi_n_1333 ,csa_tree_add_7_27_groupi_n_1368);
  nor csa_tree_add_7_27_groupi_g5803__7410(csa_tree_add_7_27_groupi_n_1385 ,csa_tree_add_7_27_groupi_n_1331 ,csa_tree_add_7_27_groupi_n_1319);
  nor csa_tree_add_7_27_groupi_g5804__6417(csa_tree_add_7_27_groupi_n_1384 ,csa_tree_add_7_27_groupi_n_1272 ,csa_tree_add_7_27_groupi_n_1326);
  or csa_tree_add_7_27_groupi_g5805__5477(csa_tree_add_7_27_groupi_n_1383 ,csa_tree_add_7_27_groupi_n_1189 ,csa_tree_add_7_27_groupi_n_1355);
  nor csa_tree_add_7_27_groupi_g5806__2398(csa_tree_add_7_27_groupi_n_1382 ,csa_tree_add_7_27_groupi_n_1284 ,csa_tree_add_7_27_groupi_n_1354);
  or csa_tree_add_7_27_groupi_g5807__5107(csa_tree_add_7_27_groupi_n_1393 ,csa_tree_add_7_27_groupi_n_1183 ,csa_tree_add_7_27_groupi_n_1332);
  or csa_tree_add_7_27_groupi_g5808__6260(csa_tree_add_7_27_groupi_n_1392 ,csa_tree_add_7_27_groupi_n_1184 ,csa_tree_add_7_27_groupi_n_1327);
  or csa_tree_add_7_27_groupi_g5809__4319(csa_tree_add_7_27_groupi_n_1391 ,csa_tree_add_7_27_groupi_n_1187 ,csa_tree_add_7_27_groupi_n_1358);
  or csa_tree_add_7_27_groupi_g5810__8428(csa_tree_add_7_27_groupi_n_1374 ,csa_tree_add_7_27_groupi_n_1105 ,csa_tree_add_7_27_groupi_n_1314);
  or csa_tree_add_7_27_groupi_g5811__5526(csa_tree_add_7_27_groupi_n_1373 ,csa_tree_add_7_27_groupi_n_999 ,csa_tree_add_7_27_groupi_n_1315);
  xnor csa_tree_add_7_27_groupi_g5812__6783(csa_tree_add_7_27_groupi_n_1372 ,csa_tree_add_7_27_groupi_n_1297 ,csa_tree_add_7_27_groupi_n_501);
  nor csa_tree_add_7_27_groupi_g5813__3680(csa_tree_add_7_27_groupi_n_1371 ,csa_tree_add_7_27_groupi_n_1119 ,csa_tree_add_7_27_groupi_n_1318);
  nor csa_tree_add_7_27_groupi_g5814__1617(csa_tree_add_7_27_groupi_n_1370 ,csa_tree_add_7_27_groupi_n_1261 ,csa_tree_add_7_27_groupi_n_1310);
  xnor csa_tree_add_7_27_groupi_g5815__2802(csa_tree_add_7_27_groupi_n_1381 ,csa_tree_add_7_27_groupi_n_1237 ,in2[2]);
  xnor csa_tree_add_7_27_groupi_g5816__1705(csa_tree_add_7_27_groupi_n_1380 ,csa_tree_add_7_27_groupi_n_1240 ,in2[14]);
  xnor csa_tree_add_7_27_groupi_g5817__5122(csa_tree_add_7_27_groupi_n_1379 ,csa_tree_add_7_27_groupi_n_1239 ,in2[8]);
  xnor csa_tree_add_7_27_groupi_g5818__8246(csa_tree_add_7_27_groupi_n_1378 ,csa_tree_add_7_27_groupi_n_1238 ,in2[5]);
  xnor csa_tree_add_7_27_groupi_g5819__7098(csa_tree_add_7_27_groupi_n_1377 ,csa_tree_add_7_27_groupi_n_1241 ,in2[11]);
  and csa_tree_add_7_27_groupi_g5820__6131(csa_tree_add_7_27_groupi_n_1376 ,csa_tree_add_7_27_groupi_n_781 ,csa_tree_add_7_27_groupi_n_1365);
  xnor csa_tree_add_7_27_groupi_g5822__1881(csa_tree_add_7_27_groupi_n_1375 ,csa_tree_add_7_27_groupi_n_1298 ,csa_tree_add_7_27_groupi_n_833);
  not csa_tree_add_7_27_groupi_g5823(csa_tree_add_7_27_groupi_n_1369 ,csa_tree_add_7_27_groupi_n_1368);
  or csa_tree_add_7_27_groupi_g5824__5115(csa_tree_add_7_27_groupi_n_1367 ,csa_tree_add_7_27_groupi_n_1016 ,csa_tree_add_7_27_groupi_n_1233);
  or csa_tree_add_7_27_groupi_g5825__7482(csa_tree_add_7_27_groupi_n_1366 ,csa_tree_add_7_27_groupi_n_1047 ,csa_tree_add_7_27_groupi_n_1248);
  or csa_tree_add_7_27_groupi_g5826__4733(csa_tree_add_7_27_groupi_n_1365 ,csa_tree_add_7_27_groupi_n_797 ,csa_tree_add_7_27_groupi_n_1298);
  or csa_tree_add_7_27_groupi_g5827__6161(csa_tree_add_7_27_groupi_n_1364 ,csa_tree_add_7_27_groupi_n_1024 ,csa_tree_add_7_27_groupi_n_1245);
  or csa_tree_add_7_27_groupi_g5828__9315(csa_tree_add_7_27_groupi_n_1363 ,csa_tree_add_7_27_groupi_n_985 ,csa_tree_add_7_27_groupi_n_1243);
  or csa_tree_add_7_27_groupi_g5829__9945(csa_tree_add_7_27_groupi_n_1362 ,csa_tree_add_7_27_groupi_n_1040 ,csa_tree_add_7_27_groupi_n_1219);
  or csa_tree_add_7_27_groupi_g5830__2883(csa_tree_add_7_27_groupi_n_1361 ,csa_tree_add_7_27_groupi_n_1017 ,csa_tree_add_7_27_groupi_n_1213);
  or csa_tree_add_7_27_groupi_g5831__2346(csa_tree_add_7_27_groupi_n_1360 ,csa_tree_add_7_27_groupi_n_996 ,csa_tree_add_7_27_groupi_n_1215);
  or csa_tree_add_7_27_groupi_g5832__1666(csa_tree_add_7_27_groupi_n_1359 ,csa_tree_add_7_27_groupi_n_1044 ,csa_tree_add_7_27_groupi_n_1252);
  and csa_tree_add_7_27_groupi_g5833__7410(csa_tree_add_7_27_groupi_n_1358 ,csa_tree_add_7_27_groupi_n_1170 ,csa_tree_add_7_27_groupi_n_1186);
  or csa_tree_add_7_27_groupi_g5834__6417(csa_tree_add_7_27_groupi_n_1357 ,csa_tree_add_7_27_groupi_n_1013 ,csa_tree_add_7_27_groupi_n_1210);
  or csa_tree_add_7_27_groupi_g5835__5477(csa_tree_add_7_27_groupi_n_1356 ,csa_tree_add_7_27_groupi_n_1088 ,csa_tree_add_7_27_groupi_n_1175);
  and csa_tree_add_7_27_groupi_g5836__2398(csa_tree_add_7_27_groupi_n_1355 ,csa_tree_add_7_27_groupi_n_1167 ,csa_tree_add_7_27_groupi_n_1188);
  or csa_tree_add_7_27_groupi_g5837__5107(csa_tree_add_7_27_groupi_n_1354 ,csa_tree_add_7_27_groupi_n_1291 ,csa_tree_add_7_27_groupi_n_1192);
  or csa_tree_add_7_27_groupi_g5838__6260(csa_tree_add_7_27_groupi_n_1353 ,csa_tree_add_7_27_groupi_n_1020 ,csa_tree_add_7_27_groupi_n_1231);
  or csa_tree_add_7_27_groupi_g5839__4319(csa_tree_add_7_27_groupi_n_1352 ,csa_tree_add_7_27_groupi_n_1012 ,csa_tree_add_7_27_groupi_n_1208);
  or csa_tree_add_7_27_groupi_g5840__8428(csa_tree_add_7_27_groupi_n_1351 ,csa_tree_add_7_27_groupi_n_1038 ,csa_tree_add_7_27_groupi_n_1209);
  or csa_tree_add_7_27_groupi_g5841__5526(csa_tree_add_7_27_groupi_n_1350 ,csa_tree_add_7_27_groupi_n_989 ,csa_tree_add_7_27_groupi_n_1224);
  or csa_tree_add_7_27_groupi_g5842__6783(csa_tree_add_7_27_groupi_n_1349 ,csa_tree_add_7_27_groupi_n_1049 ,csa_tree_add_7_27_groupi_n_1200);
  or csa_tree_add_7_27_groupi_g5843__3680(csa_tree_add_7_27_groupi_n_1348 ,csa_tree_add_7_27_groupi_n_1000 ,csa_tree_add_7_27_groupi_n_1228);
  or csa_tree_add_7_27_groupi_g5844__1617(csa_tree_add_7_27_groupi_n_1347 ,csa_tree_add_7_27_groupi_n_1048 ,csa_tree_add_7_27_groupi_n_1211);
  or csa_tree_add_7_27_groupi_g5845__2802(csa_tree_add_7_27_groupi_n_1346 ,csa_tree_add_7_27_groupi_n_1021 ,csa_tree_add_7_27_groupi_n_1227);
  or csa_tree_add_7_27_groupi_g5846__1705(csa_tree_add_7_27_groupi_n_1345 ,csa_tree_add_7_27_groupi_n_1002 ,csa_tree_add_7_27_groupi_n_1225);
  or csa_tree_add_7_27_groupi_g5847__5122(csa_tree_add_7_27_groupi_n_1344 ,csa_tree_add_7_27_groupi_n_1053 ,csa_tree_add_7_27_groupi_n_1230);
  or csa_tree_add_7_27_groupi_g5848__8246(csa_tree_add_7_27_groupi_n_1343 ,csa_tree_add_7_27_groupi_n_1022 ,csa_tree_add_7_27_groupi_n_1212);
  or csa_tree_add_7_27_groupi_g5849__7098(csa_tree_add_7_27_groupi_n_1342 ,csa_tree_add_7_27_groupi_n_1045 ,csa_tree_add_7_27_groupi_n_1202);
  or csa_tree_add_7_27_groupi_g5850__6131(csa_tree_add_7_27_groupi_n_1341 ,csa_tree_add_7_27_groupi_n_1058 ,csa_tree_add_7_27_groupi_n_1223);
  or csa_tree_add_7_27_groupi_g5851__1881(csa_tree_add_7_27_groupi_n_1340 ,csa_tree_add_7_27_groupi_n_1042 ,csa_tree_add_7_27_groupi_n_1196);
  or csa_tree_add_7_27_groupi_g5852__5115(csa_tree_add_7_27_groupi_n_1339 ,csa_tree_add_7_27_groupi_n_1096 ,csa_tree_add_7_27_groupi_n_1279);
  or csa_tree_add_7_27_groupi_g5853__7482(csa_tree_add_7_27_groupi_n_1338 ,csa_tree_add_7_27_groupi_n_998 ,csa_tree_add_7_27_groupi_n_1232);
  nor csa_tree_add_7_27_groupi_g5854__4733(csa_tree_add_7_27_groupi_n_1337 ,csa_tree_add_7_27_groupi_n_1109 ,csa_tree_add_7_27_groupi_n_1267);
  nor csa_tree_add_7_27_groupi_g5855__6161(csa_tree_add_7_27_groupi_n_1336 ,csa_tree_add_7_27_groupi_n_975 ,csa_tree_add_7_27_groupi_n_1282);
  nor csa_tree_add_7_27_groupi_g5856__9315(csa_tree_add_7_27_groupi_n_1335 ,csa_tree_add_7_27_groupi_n_1139 ,csa_tree_add_7_27_groupi_n_1283);
  and csa_tree_add_7_27_groupi_g5857__9945(csa_tree_add_7_27_groupi_n_1368 ,csa_tree_add_7_27_groupi_n_1171 ,csa_tree_add_7_27_groupi_n_1299);
  not csa_tree_add_7_27_groupi_g5858(csa_tree_add_7_27_groupi_n_1333 ,csa_tree_add_7_27_groupi_n_1334);
  and csa_tree_add_7_27_groupi_g5859__2883(csa_tree_add_7_27_groupi_n_1332 ,csa_tree_add_7_27_groupi_n_1169 ,csa_tree_add_7_27_groupi_n_1182);
  or csa_tree_add_7_27_groupi_g5860__2346(csa_tree_add_7_27_groupi_n_1331 ,csa_tree_add_7_27_groupi_n_1055 ,csa_tree_add_7_27_groupi_n_1295);
  or csa_tree_add_7_27_groupi_g5861__1666(csa_tree_add_7_27_groupi_n_1330 ,csa_tree_add_7_27_groupi_n_997 ,csa_tree_add_7_27_groupi_n_1274);
  or csa_tree_add_7_27_groupi_g5862__7410(csa_tree_add_7_27_groupi_n_1329 ,csa_tree_add_7_27_groupi_n_1008 ,csa_tree_add_7_27_groupi_n_1222);
  or csa_tree_add_7_27_groupi_g5863__6417(csa_tree_add_7_27_groupi_n_1328 ,csa_tree_add_7_27_groupi_n_1035 ,csa_tree_add_7_27_groupi_n_1275);
  and csa_tree_add_7_27_groupi_g5864__5477(csa_tree_add_7_27_groupi_n_1327 ,csa_tree_add_7_27_groupi_n_1172 ,csa_tree_add_7_27_groupi_n_1185);
  or csa_tree_add_7_27_groupi_g5865__2398(csa_tree_add_7_27_groupi_n_1326 ,csa_tree_add_7_27_groupi_n_1276 ,csa_tree_add_7_27_groupi_n_1193);
  or csa_tree_add_7_27_groupi_g5866__5107(csa_tree_add_7_27_groupi_n_1325 ,csa_tree_add_7_27_groupi_n_1031 ,csa_tree_add_7_27_groupi_n_1251);
  or csa_tree_add_7_27_groupi_g5867__6260(csa_tree_add_7_27_groupi_n_1324 ,csa_tree_add_7_27_groupi_n_1007 ,csa_tree_add_7_27_groupi_n_1218);
  or csa_tree_add_7_27_groupi_g5868__4319(csa_tree_add_7_27_groupi_n_1323 ,csa_tree_add_7_27_groupi_n_1010 ,csa_tree_add_7_27_groupi_n_1205);
  or csa_tree_add_7_27_groupi_g5869__8428(csa_tree_add_7_27_groupi_n_1322 ,csa_tree_add_7_27_groupi_n_1009 ,csa_tree_add_7_27_groupi_n_1221);
  or csa_tree_add_7_27_groupi_g5870__5526(csa_tree_add_7_27_groupi_n_1321 ,csa_tree_add_7_27_groupi_n_1131 ,csa_tree_add_7_27_groupi_n_1203);
  or csa_tree_add_7_27_groupi_g5871__6783(csa_tree_add_7_27_groupi_n_1320 ,csa_tree_add_7_27_groupi_n_988 ,csa_tree_add_7_27_groupi_n_1242);
  or csa_tree_add_7_27_groupi_g5872__3680(csa_tree_add_7_27_groupi_n_1319 ,csa_tree_add_7_27_groupi_n_980 ,csa_tree_add_7_27_groupi_n_1191);
  or csa_tree_add_7_27_groupi_g5873__1617(csa_tree_add_7_27_groupi_n_1318 ,csa_tree_add_7_27_groupi_n_994 ,csa_tree_add_7_27_groupi_n_1194);
  or csa_tree_add_7_27_groupi_g5874__2802(csa_tree_add_7_27_groupi_n_1317 ,csa_tree_add_7_27_groupi_n_1158 ,csa_tree_add_7_27_groupi_n_1296);
  nor csa_tree_add_7_27_groupi_g5875__1705(csa_tree_add_7_27_groupi_n_1316 ,csa_tree_add_7_27_groupi_n_1157 ,csa_tree_add_7_27_groupi_n_1297);
  nor csa_tree_add_7_27_groupi_g5876__5122(csa_tree_add_7_27_groupi_n_1315 ,csa_tree_add_7_27_groupi_n_35 ,csa_tree_add_7_27_groupi_n_512);
  nor csa_tree_add_7_27_groupi_g5877__8246(csa_tree_add_7_27_groupi_n_1314 ,csa_tree_add_7_27_groupi_n_94 ,csa_tree_add_7_27_groupi_n_1236);
  nor csa_tree_add_7_27_groupi_g5878__7098(csa_tree_add_7_27_groupi_n_1313 ,csa_tree_add_7_27_groupi_n_17 ,csa_tree_add_7_27_groupi_n_512);
  nor csa_tree_add_7_27_groupi_g5879__6131(csa_tree_add_7_27_groupi_n_1312 ,csa_tree_add_7_27_groupi_n_48 ,csa_tree_add_7_27_groupi_n_1236);
  nor csa_tree_add_7_27_groupi_g5880__1881(csa_tree_add_7_27_groupi_n_1311 ,csa_tree_add_7_27_groupi_n_66 ,csa_tree_add_7_27_groupi_n_511);
  or csa_tree_add_7_27_groupi_g5881__5115(csa_tree_add_7_27_groupi_n_1310 ,csa_tree_add_7_27_groupi_n_1280 ,csa_tree_add_7_27_groupi_n_1190);
  nor csa_tree_add_7_27_groupi_g5882__7482(csa_tree_add_7_27_groupi_n_1309 ,csa_tree_add_7_27_groupi_n_1054 ,csa_tree_add_7_27_groupi_n_1260);
  nor csa_tree_add_7_27_groupi_g5883__4733(csa_tree_add_7_27_groupi_n_1308 ,csa_tree_add_7_27_groupi_n_976 ,csa_tree_add_7_27_groupi_n_1262);
  xnor csa_tree_add_7_27_groupi_g5884__6161(csa_tree_add_7_27_groupi_n_1307 ,csa_tree_add_7_27_groupi_n_1166 ,csa_tree_add_7_27_groupi_n_1155);
  xnor csa_tree_add_7_27_groupi_g5885(csa_tree_add_7_27_groupi_n_1306 ,csa_tree_add_7_27_groupi_n_484 ,csa_tree_add_7_27_groupi_n_1164);
  xnor csa_tree_add_7_27_groupi_g5886(csa_tree_add_7_27_groupi_n_1305 ,csa_tree_add_7_27_groupi_n_1167 ,in2[14]);
  xnor csa_tree_add_7_27_groupi_g5887(csa_tree_add_7_27_groupi_n_1304 ,csa_tree_add_7_27_groupi_n_1169 ,in2[5]);
  xnor csa_tree_add_7_27_groupi_g5888(csa_tree_add_7_27_groupi_n_1303 ,csa_tree_add_7_27_groupi_n_1172 ,in2[8]);
  xnor csa_tree_add_7_27_groupi_g5889(csa_tree_add_7_27_groupi_n_1302 ,csa_tree_add_7_27_groupi_n_1170 ,in2[11]);
  xnor csa_tree_add_7_27_groupi_g5890(csa_tree_add_7_27_groupi_n_1301 ,csa_tree_add_7_27_groupi_n_486 ,csa_tree_add_7_27_groupi_n_1161);
  xnor csa_tree_add_7_27_groupi_g5891(csa_tree_add_7_27_groupi_n_1300 ,csa_tree_add_7_27_groupi_n_485 ,csa_tree_add_7_27_groupi_n_1157);
  and csa_tree_add_7_27_groupi_g5893(csa_tree_add_7_27_groupi_n_1334 ,csa_tree_add_7_27_groupi_n_1281 ,csa_tree_add_7_27_groupi_n_1296);
  not csa_tree_add_7_27_groupi_g5895(csa_tree_add_7_27_groupi_n_1296 ,csa_tree_add_7_27_groupi_n_1297);
  and csa_tree_add_7_27_groupi_g5896(csa_tree_add_7_27_groupi_n_1295 ,in1[0] ,csa_tree_add_7_27_groupi_n_493);
  or csa_tree_add_7_27_groupi_g5897(csa_tree_add_7_27_groupi_n_1294 ,csa_tree_add_7_27_groupi_n_983 ,csa_tree_add_7_27_groupi_n_1136);
  or csa_tree_add_7_27_groupi_g5898(csa_tree_add_7_27_groupi_n_1293 ,csa_tree_add_7_27_groupi_n_1018 ,csa_tree_add_7_27_groupi_n_1145);
  or csa_tree_add_7_27_groupi_g5899(csa_tree_add_7_27_groupi_n_1292 ,csa_tree_add_7_27_groupi_n_1043 ,csa_tree_add_7_27_groupi_n_1086);
  and csa_tree_add_7_27_groupi_g5900(csa_tree_add_7_27_groupi_n_1291 ,in1[0] ,csa_tree_add_7_27_groupi_n_491);
  or csa_tree_add_7_27_groupi_g5901(csa_tree_add_7_27_groupi_n_1290 ,csa_tree_add_7_27_groupi_n_1025 ,csa_tree_add_7_27_groupi_n_1080);
  or csa_tree_add_7_27_groupi_g5902(csa_tree_add_7_27_groupi_n_1289 ,csa_tree_add_7_27_groupi_n_1026 ,csa_tree_add_7_27_groupi_n_1087);
  or csa_tree_add_7_27_groupi_g5903(csa_tree_add_7_27_groupi_n_1288 ,csa_tree_add_7_27_groupi_n_982 ,csa_tree_add_7_27_groupi_n_1081);
  or csa_tree_add_7_27_groupi_g5904(csa_tree_add_7_27_groupi_n_1287 ,csa_tree_add_7_27_groupi_n_1046 ,csa_tree_add_7_27_groupi_n_1108);
  or csa_tree_add_7_27_groupi_g5905(csa_tree_add_7_27_groupi_n_1286 ,csa_tree_add_7_27_groupi_n_992 ,csa_tree_add_7_27_groupi_n_1084);
  or csa_tree_add_7_27_groupi_g5906(csa_tree_add_7_27_groupi_n_1285 ,csa_tree_add_7_27_groupi_n_1030 ,csa_tree_add_7_27_groupi_n_1148);
  or csa_tree_add_7_27_groupi_g5907(csa_tree_add_7_27_groupi_n_1284 ,csa_tree_add_7_27_groupi_n_1052 ,csa_tree_add_7_27_groupi_n_1079);
  or csa_tree_add_7_27_groupi_g5908(csa_tree_add_7_27_groupi_n_1283 ,csa_tree_add_7_27_groupi_n_1138 ,csa_tree_add_7_27_groupi_n_974);
  or csa_tree_add_7_27_groupi_g5909(csa_tree_add_7_27_groupi_n_1282 ,csa_tree_add_7_27_groupi_n_1116 ,csa_tree_add_7_27_groupi_n_1143);
  or csa_tree_add_7_27_groupi_g5910(csa_tree_add_7_27_groupi_n_1281 ,in2[2] ,csa_tree_add_7_27_groupi_n_1174);
  and csa_tree_add_7_27_groupi_g5911(csa_tree_add_7_27_groupi_n_1280 ,in1[0] ,csa_tree_add_7_27_groupi_n_494);
  nor csa_tree_add_7_27_groupi_g5912(csa_tree_add_7_27_groupi_n_1279 ,csa_tree_add_7_27_groupi_n_91 ,csa_tree_add_7_27_groupi_n_691);
  nor csa_tree_add_7_27_groupi_g5913(csa_tree_add_7_27_groupi_n_1278 ,csa_tree_add_7_27_groupi_n_721 ,csa_tree_add_7_27_groupi_n_1166);
  or csa_tree_add_7_27_groupi_g5914(csa_tree_add_7_27_groupi_n_1277 ,csa_tree_add_7_27_groupi_n_1039 ,csa_tree_add_7_27_groupi_n_1078);
  and csa_tree_add_7_27_groupi_g5915(csa_tree_add_7_27_groupi_n_1276 ,in1[0] ,csa_tree_add_7_27_groupi_n_492);
  nor csa_tree_add_7_27_groupi_g5916(csa_tree_add_7_27_groupi_n_1275 ,csa_tree_add_7_27_groupi_n_358 ,csa_tree_add_7_27_groupi_n_682);
  nor csa_tree_add_7_27_groupi_g5917(csa_tree_add_7_27_groupi_n_1274 ,csa_tree_add_7_27_groupi_n_358 ,csa_tree_add_7_27_groupi_n_709);
  or csa_tree_add_7_27_groupi_g5918(csa_tree_add_7_27_groupi_n_1273 ,csa_tree_add_7_27_groupi_n_1165 ,csa_tree_add_7_27_groupi_n_1155);
  or csa_tree_add_7_27_groupi_g5919(csa_tree_add_7_27_groupi_n_1272 ,csa_tree_add_7_27_groupi_n_1050 ,csa_tree_add_7_27_groupi_n_1099);
  or csa_tree_add_7_27_groupi_g5920(csa_tree_add_7_27_groupi_n_1271 ,csa_tree_add_7_27_groupi_n_984 ,csa_tree_add_7_27_groupi_n_1094);
  or csa_tree_add_7_27_groupi_g5921(csa_tree_add_7_27_groupi_n_1270 ,csa_tree_add_7_27_groupi_n_986 ,csa_tree_add_7_27_groupi_n_1141);
  or csa_tree_add_7_27_groupi_g5922(csa_tree_add_7_27_groupi_n_1269 ,csa_tree_add_7_27_groupi_n_993 ,csa_tree_add_7_27_groupi_n_1097);
  or csa_tree_add_7_27_groupi_g5923(csa_tree_add_7_27_groupi_n_1268 ,csa_tree_add_7_27_groupi_n_1004 ,csa_tree_add_7_27_groupi_n_1057);
  or csa_tree_add_7_27_groupi_g5924(csa_tree_add_7_27_groupi_n_1267 ,csa_tree_add_7_27_groupi_n_1140 ,csa_tree_add_7_27_groupi_n_973);
  or csa_tree_add_7_27_groupi_g5925(csa_tree_add_7_27_groupi_n_1266 ,csa_tree_add_7_27_groupi_n_1041 ,csa_tree_add_7_27_groupi_n_1098);
  or csa_tree_add_7_27_groupi_g5926(csa_tree_add_7_27_groupi_n_1265 ,csa_tree_add_7_27_groupi_n_1034 ,csa_tree_add_7_27_groupi_n_1149);
  or csa_tree_add_7_27_groupi_g5927(csa_tree_add_7_27_groupi_n_1264 ,csa_tree_add_7_27_groupi_n_1028 ,csa_tree_add_7_27_groupi_n_1093);
  or csa_tree_add_7_27_groupi_g5928(csa_tree_add_7_27_groupi_n_1263 ,csa_tree_add_7_27_groupi_n_1003 ,csa_tree_add_7_27_groupi_n_1100);
  or csa_tree_add_7_27_groupi_g5929(csa_tree_add_7_27_groupi_n_1262 ,csa_tree_add_7_27_groupi_n_1151 ,csa_tree_add_7_27_groupi_n_1132);
  or csa_tree_add_7_27_groupi_g5930(csa_tree_add_7_27_groupi_n_1261 ,csa_tree_add_7_27_groupi_n_1056 ,csa_tree_add_7_27_groupi_n_1095);
  or csa_tree_add_7_27_groupi_g5931(csa_tree_add_7_27_groupi_n_1260 ,csa_tree_add_7_27_groupi_n_894 ,csa_tree_add_7_27_groupi_n_981);
  or csa_tree_add_7_27_groupi_g5932(csa_tree_add_7_27_groupi_n_1259 ,csa_tree_add_7_27_groupi_n_1032 ,csa_tree_add_7_27_groupi_n_1077);
  or csa_tree_add_7_27_groupi_g5933(csa_tree_add_7_27_groupi_n_1258 ,csa_tree_add_7_27_groupi_n_990 ,csa_tree_add_7_27_groupi_n_1124);
  or csa_tree_add_7_27_groupi_g5934(csa_tree_add_7_27_groupi_n_1257 ,csa_tree_add_7_27_groupi_n_1023 ,csa_tree_add_7_27_groupi_n_1090);
  nor csa_tree_add_7_27_groupi_g5935(csa_tree_add_7_27_groupi_n_1256 ,csa_tree_add_7_27_groupi_n_338 ,csa_tree_add_7_27_groupi_n_703);
  nor csa_tree_add_7_27_groupi_g5936(csa_tree_add_7_27_groupi_n_1255 ,csa_tree_add_7_27_groupi_n_349 ,csa_tree_add_7_27_groupi_n_700);
  nor csa_tree_add_7_27_groupi_g5937(csa_tree_add_7_27_groupi_n_1254 ,csa_tree_add_7_27_groupi_n_11 ,csa_tree_add_7_27_groupi_n_712);
  nor csa_tree_add_7_27_groupi_g5938(csa_tree_add_7_27_groupi_n_1253 ,csa_tree_add_7_27_groupi_n_377 ,csa_tree_add_7_27_groupi_n_694);
  nor csa_tree_add_7_27_groupi_g5939(csa_tree_add_7_27_groupi_n_1252 ,csa_tree_add_7_27_groupi_n_349 ,csa_tree_add_7_27_groupi_n_713);
  nor csa_tree_add_7_27_groupi_g5940(csa_tree_add_7_27_groupi_n_1251 ,csa_tree_add_7_27_groupi_n_451 ,csa_tree_add_7_27_groupi_n_685);
  nor csa_tree_add_7_27_groupi_g5941(csa_tree_add_7_27_groupi_n_1250 ,csa_tree_add_7_27_groupi_n_374 ,csa_tree_add_7_27_groupi_n_704);
  nor csa_tree_add_7_27_groupi_g5942(csa_tree_add_7_27_groupi_n_1249 ,csa_tree_add_7_27_groupi_n_367 ,csa_tree_add_7_27_groupi_n_686);
  nor csa_tree_add_7_27_groupi_g5943(csa_tree_add_7_27_groupi_n_1248 ,csa_tree_add_7_27_groupi_n_271 ,csa_tree_add_7_27_groupi_n_688);
  nor csa_tree_add_7_27_groupi_g5944(csa_tree_add_7_27_groupi_n_1247 ,csa_tree_add_7_27_groupi_n_320 ,csa_tree_add_7_27_groupi_n_706);
  nor csa_tree_add_7_27_groupi_g5945(csa_tree_add_7_27_groupi_n_1246 ,csa_tree_add_7_27_groupi_n_389 ,csa_tree_add_7_27_groupi_n_695);
  nor csa_tree_add_7_27_groupi_g5946(csa_tree_add_7_27_groupi_n_1245 ,csa_tree_add_7_27_groupi_n_322 ,csa_tree_add_7_27_groupi_n_710);
  nor csa_tree_add_7_27_groupi_g5947(csa_tree_add_7_27_groupi_n_1244 ,csa_tree_add_7_27_groupi_n_449 ,csa_tree_add_7_27_groupi_n_692);
  nor csa_tree_add_7_27_groupi_g5948(csa_tree_add_7_27_groupi_n_1243 ,csa_tree_add_7_27_groupi_n_346 ,csa_tree_add_7_27_groupi_n_697);
  nor csa_tree_add_7_27_groupi_g5949(csa_tree_add_7_27_groupi_n_1242 ,csa_tree_add_7_27_groupi_n_274 ,csa_tree_add_7_27_groupi_n_679);
  or csa_tree_add_7_27_groupi_g5950(csa_tree_add_7_27_groupi_n_1241 ,csa_tree_add_7_27_groupi_n_113 ,csa_tree_add_7_27_groupi_n_978);
  or csa_tree_add_7_27_groupi_g5951(csa_tree_add_7_27_groupi_n_1240 ,csa_tree_add_7_27_groupi_n_116 ,csa_tree_add_7_27_groupi_n_979);
  or csa_tree_add_7_27_groupi_g5952(csa_tree_add_7_27_groupi_n_1239 ,csa_tree_add_7_27_groupi_n_111 ,csa_tree_add_7_27_groupi_n_977);
  or csa_tree_add_7_27_groupi_g5953(csa_tree_add_7_27_groupi_n_1238 ,csa_tree_add_7_27_groupi_n_108 ,csa_tree_add_7_27_groupi_n_971);
  or csa_tree_add_7_27_groupi_g5954(csa_tree_add_7_27_groupi_n_1237 ,csa_tree_add_7_27_groupi_n_115 ,csa_tree_add_7_27_groupi_n_972);
  and csa_tree_add_7_27_groupi_g5955(csa_tree_add_7_27_groupi_n_1299 ,csa_tree_add_7_27_groupi_n_1168 ,csa_tree_add_7_27_groupi_n_1173);
  and csa_tree_add_7_27_groupi_g5956(csa_tree_add_7_27_groupi_n_1298 ,csa_tree_add_7_27_groupi_n_788 ,csa_tree_add_7_27_groupi_n_1115);
  and csa_tree_add_7_27_groupi_g5957(csa_tree_add_7_27_groupi_n_1297 ,in2[2] ,csa_tree_add_7_27_groupi_n_1174);
  nor csa_tree_add_7_27_groupi_g5958(csa_tree_add_7_27_groupi_n_1235 ,csa_tree_add_7_27_groupi_n_259 ,csa_tree_add_7_27_groupi_n_706);
  nor csa_tree_add_7_27_groupi_g5959(csa_tree_add_7_27_groupi_n_1234 ,csa_tree_add_7_27_groupi_n_325 ,csa_tree_add_7_27_groupi_n_707);
  nor csa_tree_add_7_27_groupi_g5960(csa_tree_add_7_27_groupi_n_1233 ,csa_tree_add_7_27_groupi_n_307 ,csa_tree_add_7_27_groupi_n_701);
  nor csa_tree_add_7_27_groupi_g5961(csa_tree_add_7_27_groupi_n_1232 ,csa_tree_add_7_27_groupi_n_259 ,csa_tree_add_7_27_groupi_n_688);
  nor csa_tree_add_7_27_groupi_g5962(csa_tree_add_7_27_groupi_n_1231 ,csa_tree_add_7_27_groupi_n_286 ,csa_tree_add_7_27_groupi_n_707);
  nor csa_tree_add_7_27_groupi_g5963(csa_tree_add_7_27_groupi_n_1230 ,csa_tree_add_7_27_groupi_n_271 ,csa_tree_add_7_27_groupi_n_697);
  nor csa_tree_add_7_27_groupi_g5964(csa_tree_add_7_27_groupi_n_1229 ,csa_tree_add_7_27_groupi_n_253 ,csa_tree_add_7_27_groupi_n_683);
  nor csa_tree_add_7_27_groupi_g5965(csa_tree_add_7_27_groupi_n_1228 ,csa_tree_add_7_27_groupi_n_325 ,csa_tree_add_7_27_groupi_n_698);
  nor csa_tree_add_7_27_groupi_g5966(csa_tree_add_7_27_groupi_n_1227 ,csa_tree_add_7_27_groupi_n_435 ,csa_tree_add_7_27_groupi_n_689);
  nor csa_tree_add_7_27_groupi_g5967(csa_tree_add_7_27_groupi_n_1226 ,csa_tree_add_7_27_groupi_n_443 ,csa_tree_add_7_27_groupi_n_679);
  nor csa_tree_add_7_27_groupi_g5968(csa_tree_add_7_27_groupi_n_1225 ,csa_tree_add_7_27_groupi_n_322 ,csa_tree_add_7_27_groupi_n_689);
  nor csa_tree_add_7_27_groupi_g5969(csa_tree_add_7_27_groupi_n_1224 ,csa_tree_add_7_27_groupi_n_274 ,csa_tree_add_7_27_groupi_n_710);
  nor csa_tree_add_7_27_groupi_g5970(csa_tree_add_7_27_groupi_n_1223 ,csa_tree_add_7_27_groupi_n_295 ,csa_tree_add_7_27_groupi_n_680);
  nor csa_tree_add_7_27_groupi_g5971(csa_tree_add_7_27_groupi_n_1222 ,csa_tree_add_7_27_groupi_n_430 ,csa_tree_add_7_27_groupi_n_698);
  nor csa_tree_add_7_27_groupi_g5972(csa_tree_add_7_27_groupi_n_1221 ,csa_tree_add_7_27_groupi_n_253 ,csa_tree_add_7_27_groupi_n_667);
  nor csa_tree_add_7_27_groupi_g5973(csa_tree_add_7_27_groupi_n_1220 ,csa_tree_add_7_27_groupi_n_286 ,csa_tree_add_7_27_groupi_n_701);
  nor csa_tree_add_7_27_groupi_g5974(csa_tree_add_7_27_groupi_n_1219 ,csa_tree_add_7_27_groupi_n_385 ,csa_tree_add_7_27_groupi_n_680);
  nor csa_tree_add_7_27_groupi_g5975(csa_tree_add_7_27_groupi_n_1218 ,csa_tree_add_7_27_groupi_n_340 ,csa_tree_add_7_27_groupi_n_683);
  nor csa_tree_add_7_27_groupi_g5976(csa_tree_add_7_27_groupi_n_1217 ,csa_tree_add_7_27_groupi_n_8 ,csa_tree_add_7_27_groupi_n_665);
  nor csa_tree_add_7_27_groupi_g5977(csa_tree_add_7_27_groupi_n_1216 ,csa_tree_add_7_27_groupi_n_405 ,csa_tree_add_7_27_groupi_n_692);
  nor csa_tree_add_7_27_groupi_g5978(csa_tree_add_7_27_groupi_n_1215 ,csa_tree_add_7_27_groupi_n_412 ,csa_tree_add_7_27_groupi_n_1070);
  nor csa_tree_add_7_27_groupi_g5979(csa_tree_add_7_27_groupi_n_1214 ,csa_tree_add_7_27_groupi_n_295 ,csa_tree_add_7_27_groupi_n_663);
  nor csa_tree_add_7_27_groupi_g5980(csa_tree_add_7_27_groupi_n_1213 ,csa_tree_add_7_27_groupi_n_307 ,csa_tree_add_7_27_groupi_n_661);
  nor csa_tree_add_7_27_groupi_g5981(csa_tree_add_7_27_groupi_n_1212 ,csa_tree_add_7_27_groupi_n_387 ,csa_tree_add_7_27_groupi_n_700);
  nor csa_tree_add_7_27_groupi_g5982(csa_tree_add_7_27_groupi_n_1211 ,csa_tree_add_7_27_groupi_n_395 ,csa_tree_add_7_27_groupi_n_1062);
  nor csa_tree_add_7_27_groupi_g5983(csa_tree_add_7_27_groupi_n_1210 ,csa_tree_add_7_27_groupi_n_382 ,csa_tree_add_7_27_groupi_n_682);
  nor csa_tree_add_7_27_groupi_g5984(csa_tree_add_7_27_groupi_n_1209 ,csa_tree_add_7_27_groupi_n_423 ,csa_tree_add_7_27_groupi_n_1066);
  nor csa_tree_add_7_27_groupi_g5985(csa_tree_add_7_27_groupi_n_1208 ,csa_tree_add_7_27_groupi_n_346 ,csa_tree_add_7_27_groupi_n_691);
  nor csa_tree_add_7_27_groupi_g5986(csa_tree_add_7_27_groupi_n_1207 ,csa_tree_add_7_27_groupi_n_392 ,csa_tree_add_7_27_groupi_n_695);
  nor csa_tree_add_7_27_groupi_g5987(csa_tree_add_7_27_groupi_n_1206 ,csa_tree_add_7_27_groupi_n_340 ,csa_tree_add_7_27_groupi_n_686);
  nor csa_tree_add_7_27_groupi_g5988(csa_tree_add_7_27_groupi_n_1205 ,csa_tree_add_7_27_groupi_n_441 ,csa_tree_add_7_27_groupi_n_713);
  nor csa_tree_add_7_27_groupi_g5989(csa_tree_add_7_27_groupi_n_1204 ,csa_tree_add_7_27_groupi_n_432 ,csa_tree_add_7_27_groupi_n_661);
  nor csa_tree_add_7_27_groupi_g5990(csa_tree_add_7_27_groupi_n_1203 ,csa_tree_add_7_27_groupi_n_371 ,csa_tree_add_7_27_groupi_n_665);
  nor csa_tree_add_7_27_groupi_g5991(csa_tree_add_7_27_groupi_n_1202 ,csa_tree_add_7_27_groupi_n_415 ,csa_tree_add_7_27_groupi_n_694);
  nor csa_tree_add_7_27_groupi_g5992(csa_tree_add_7_27_groupi_n_1201 ,csa_tree_add_7_27_groupi_n_427 ,csa_tree_add_7_27_groupi_n_1074);
  nor csa_tree_add_7_27_groupi_g5993(csa_tree_add_7_27_groupi_n_1200 ,csa_tree_add_7_27_groupi_n_400 ,csa_tree_add_7_27_groupi_n_709);
  nor csa_tree_add_7_27_groupi_g5994(csa_tree_add_7_27_groupi_n_1199 ,csa_tree_add_7_27_groupi_n_420 ,csa_tree_add_7_27_groupi_n_704);
  nor csa_tree_add_7_27_groupi_g5995(csa_tree_add_7_27_groupi_n_1198 ,csa_tree_add_7_27_groupi_n_439 ,csa_tree_add_7_27_groupi_n_667);
  nor csa_tree_add_7_27_groupi_g5996(csa_tree_add_7_27_groupi_n_1197 ,csa_tree_add_7_27_groupi_n_397 ,csa_tree_add_7_27_groupi_n_663);
  nor csa_tree_add_7_27_groupi_g5997(csa_tree_add_7_27_groupi_n_1196 ,csa_tree_add_7_27_groupi_n_403 ,csa_tree_add_7_27_groupi_n_685);
  nor csa_tree_add_7_27_groupi_g5998(csa_tree_add_7_27_groupi_n_1195 ,csa_tree_add_7_27_groupi_n_409 ,csa_tree_add_7_27_groupi_n_712);
  nor csa_tree_add_7_27_groupi_g5999(csa_tree_add_7_27_groupi_n_1194 ,csa_tree_add_7_27_groupi_n_305 ,csa_tree_add_7_27_groupi_n_515);
  nor csa_tree_add_7_27_groupi_g6000(csa_tree_add_7_27_groupi_n_1193 ,csa_tree_add_7_27_groupi_n_269 ,csa_tree_add_7_27_groupi_n_1075);
  nor csa_tree_add_7_27_groupi_g6001(csa_tree_add_7_27_groupi_n_1192 ,csa_tree_add_7_27_groupi_n_344 ,csa_tree_add_7_27_groupi_n_515);
  nor csa_tree_add_7_27_groupi_g6002(csa_tree_add_7_27_groupi_n_1191 ,csa_tree_add_7_27_groupi_n_284 ,csa_tree_add_7_27_groupi_n_1075);
  nor csa_tree_add_7_27_groupi_g6003(csa_tree_add_7_27_groupi_n_1190 ,csa_tree_add_7_27_groupi_n_317 ,csa_tree_add_7_27_groupi_n_514);
  nor csa_tree_add_7_27_groupi_g6004(csa_tree_add_7_27_groupi_n_1189 ,in2[14] ,csa_tree_add_7_27_groupi_n_489);
  or csa_tree_add_7_27_groupi_g6005(csa_tree_add_7_27_groupi_n_1188 ,csa_tree_add_7_27_groupi_n_730 ,csa_tree_add_7_27_groupi_n_1155);
  and csa_tree_add_7_27_groupi_g6006(csa_tree_add_7_27_groupi_n_1187 ,csa_tree_add_7_27_groupi_n_744 ,csa_tree_add_7_27_groupi_n_486);
  or csa_tree_add_7_27_groupi_g6007(csa_tree_add_7_27_groupi_n_1186 ,csa_tree_add_7_27_groupi_n_477 ,csa_tree_add_7_27_groupi_n_496);
  or csa_tree_add_7_27_groupi_g6008(csa_tree_add_7_27_groupi_n_1185 ,csa_tree_add_7_27_groupi_n_473 ,csa_tree_add_7_27_groupi_n_484);
  and csa_tree_add_7_27_groupi_g6009(csa_tree_add_7_27_groupi_n_1184 ,csa_tree_add_7_27_groupi_n_474 ,csa_tree_add_7_27_groupi_n_503);
  and csa_tree_add_7_27_groupi_g6010(csa_tree_add_7_27_groupi_n_1183 ,csa_tree_add_7_27_groupi_n_479 ,csa_tree_add_7_27_groupi_n_485);
  or csa_tree_add_7_27_groupi_g6011(csa_tree_add_7_27_groupi_n_1182 ,csa_tree_add_7_27_groupi_n_480 ,csa_tree_add_7_27_groupi_n_498);
  or csa_tree_add_7_27_groupi_g6012(csa_tree_add_7_27_groupi_n_1181 ,csa_tree_add_7_27_groupi_n_727 ,csa_tree_add_7_27_groupi_n_501);
  or csa_tree_add_7_27_groupi_g6013(csa_tree_add_7_27_groupi_n_1180 ,csa_tree_add_7_27_groupi_n_729 ,csa_tree_add_7_27_groupi_n_671);
  nor csa_tree_add_7_27_groupi_g6014(csa_tree_add_7_27_groupi_n_1179 ,csa_tree_add_7_27_groupi_n_1163 ,csa_tree_add_7_27_groupi_n_503);
  nor csa_tree_add_7_27_groupi_g6015(csa_tree_add_7_27_groupi_n_1178 ,csa_tree_add_7_27_groupi_n_1158 ,csa_tree_add_7_27_groupi_n_498);
  or csa_tree_add_7_27_groupi_g6016(csa_tree_add_7_27_groupi_n_1177 ,csa_tree_add_7_27_groupi_n_728 ,csa_tree_add_7_27_groupi_n_669);
  nor csa_tree_add_7_27_groupi_g6017(csa_tree_add_7_27_groupi_n_1176 ,csa_tree_add_7_27_groupi_n_1160 ,csa_tree_add_7_27_groupi_n_496);
  nor csa_tree_add_7_27_groupi_g6018(csa_tree_add_7_27_groupi_n_1175 ,csa_tree_add_7_27_groupi_n_446 ,csa_tree_add_7_27_groupi_n_703);
  xnor csa_tree_add_7_27_groupi_g6020(csa_tree_add_7_27_groupi_n_1236 ,csa_tree_add_7_27_groupi_n_970 ,csa_tree_add_7_27_groupi_n_841);
  not csa_tree_add_7_27_groupi_g6022(csa_tree_add_7_27_groupi_n_1165 ,csa_tree_add_7_27_groupi_n_1166);
  not csa_tree_add_7_27_groupi_g6023(csa_tree_add_7_27_groupi_n_1163 ,csa_tree_add_7_27_groupi_n_1164);
  not csa_tree_add_7_27_groupi_g6025(csa_tree_add_7_27_groupi_n_1160 ,csa_tree_add_7_27_groupi_n_1161);
  not csa_tree_add_7_27_groupi_g6027(csa_tree_add_7_27_groupi_n_1158 ,csa_tree_add_7_27_groupi_n_500);
  buf csa_tree_add_7_27_groupi_g6029(csa_tree_add_7_27_groupi_n_1155 ,csa_tree_add_7_27_groupi_n_1153);
  not csa_tree_add_7_27_groupi_g6030(csa_tree_add_7_27_groupi_n_1154 ,csa_tree_add_7_27_groupi_n_1153);
  nor csa_tree_add_7_27_groupi_g6031(csa_tree_add_7_27_groupi_n_1152 ,csa_tree_add_7_27_groupi_n_272 ,csa_tree_add_7_27_groupi_n_176);
  nor csa_tree_add_7_27_groupi_g6032(csa_tree_add_7_27_groupi_n_1151 ,csa_tree_add_7_27_groupi_n_242 ,csa_tree_add_7_27_groupi_n_108);
  or csa_tree_add_7_27_groupi_g6033(csa_tree_add_7_27_groupi_n_1150 ,csa_tree_add_7_27_groupi_n_877 ,csa_tree_add_7_27_groupi_n_959);
  nor csa_tree_add_7_27_groupi_g6034(csa_tree_add_7_27_groupi_n_1149 ,csa_tree_add_7_27_groupi_n_417 ,csa_tree_add_7_27_groupi_n_170);
  nor csa_tree_add_7_27_groupi_g6035(csa_tree_add_7_27_groupi_n_1148 ,csa_tree_add_7_27_groupi_n_308 ,csa_tree_add_7_27_groupi_n_175);
  or csa_tree_add_7_27_groupi_g6036(csa_tree_add_7_27_groupi_n_1147 ,csa_tree_add_7_27_groupi_n_880 ,csa_tree_add_7_27_groupi_n_956);
  or csa_tree_add_7_27_groupi_g6037(csa_tree_add_7_27_groupi_n_1146 ,csa_tree_add_7_27_groupi_n_852 ,csa_tree_add_7_27_groupi_n_961);
  nor csa_tree_add_7_27_groupi_g6038(csa_tree_add_7_27_groupi_n_1145 ,csa_tree_add_7_27_groupi_n_251 ,csa_tree_add_7_27_groupi_n_146);
  nor csa_tree_add_7_27_groupi_g6039(csa_tree_add_7_27_groupi_n_1144 ,csa_tree_add_7_27_groupi_n_326 ,csa_tree_add_7_27_groupi_n_128);
  nor csa_tree_add_7_27_groupi_g6040(csa_tree_add_7_27_groupi_n_1143 ,csa_tree_add_7_27_groupi_n_350 ,csa_tree_add_7_27_groupi_n_127);
  or csa_tree_add_7_27_groupi_g6041(csa_tree_add_7_27_groupi_n_1142 ,csa_tree_add_7_27_groupi_n_856 ,csa_tree_add_7_27_groupi_n_954);
  nor csa_tree_add_7_27_groupi_g6042(csa_tree_add_7_27_groupi_n_1141 ,csa_tree_add_7_27_groupi_n_260 ,csa_tree_add_7_27_groupi_n_143);
  nor csa_tree_add_7_27_groupi_g6043(csa_tree_add_7_27_groupi_n_1140 ,csa_tree_add_7_27_groupi_n_239 ,csa_tree_add_7_27_groupi_n_110);
  nor csa_tree_add_7_27_groupi_g6044(csa_tree_add_7_27_groupi_n_1139 ,csa_tree_add_7_27_groupi_n_362 ,csa_tree_add_7_27_groupi_n_230);
  nor csa_tree_add_7_27_groupi_g6045(csa_tree_add_7_27_groupi_n_1138 ,csa_tree_add_7_27_groupi_n_248 ,csa_tree_add_7_27_groupi_n_113);
  nor csa_tree_add_7_27_groupi_g6046(csa_tree_add_7_27_groupi_n_1137 ,csa_tree_add_7_27_groupi_n_338 ,csa_tree_add_7_27_groupi_n_194);
  nor csa_tree_add_7_27_groupi_g6047(csa_tree_add_7_27_groupi_n_1136 ,csa_tree_add_7_27_groupi_n_275 ,csa_tree_add_7_27_groupi_n_197);
  or csa_tree_add_7_27_groupi_g6048(csa_tree_add_7_27_groupi_n_1135 ,csa_tree_add_7_27_groupi_n_885 ,csa_tree_add_7_27_groupi_n_950);
  nor csa_tree_add_7_27_groupi_g6049(csa_tree_add_7_27_groupi_n_1134 ,csa_tree_add_7_27_groupi_n_287 ,csa_tree_add_7_27_groupi_n_176);
  nor csa_tree_add_7_27_groupi_g6050(csa_tree_add_7_27_groupi_n_1133 ,csa_tree_add_7_27_groupi_n_359 ,csa_tree_add_7_27_groupi_n_193);
  nor csa_tree_add_7_27_groupi_g6051(csa_tree_add_7_27_groupi_n_1132 ,csa_tree_add_7_27_groupi_n_19 ,csa_tree_add_7_27_groupi_n_215);
  nor csa_tree_add_7_27_groupi_g6052(csa_tree_add_7_27_groupi_n_1131 ,csa_tree_add_7_27_groupi_n_378 ,csa_tree_add_7_27_groupi_n_142);
  nor csa_tree_add_7_27_groupi_g6053(csa_tree_add_7_27_groupi_n_1130 ,csa_tree_add_7_27_groupi_n_293 ,csa_tree_add_7_27_groupi_n_131);
  or csa_tree_add_7_27_groupi_g6054(csa_tree_add_7_27_groupi_n_1129 ,csa_tree_add_7_27_groupi_n_881 ,csa_tree_add_7_27_groupi_n_955);
  or csa_tree_add_7_27_groupi_g6055(csa_tree_add_7_27_groupi_n_1128 ,csa_tree_add_7_27_groupi_n_850 ,csa_tree_add_7_27_groupi_n_932);
  or csa_tree_add_7_27_groupi_g6056(csa_tree_add_7_27_groupi_n_1127 ,csa_tree_add_7_27_groupi_n_851 ,csa_tree_add_7_27_groupi_n_945);
  or csa_tree_add_7_27_groupi_g6057(csa_tree_add_7_27_groupi_n_1126 ,csa_tree_add_7_27_groupi_n_858 ,csa_tree_add_7_27_groupi_n_935);
  or csa_tree_add_7_27_groupi_g6058(csa_tree_add_7_27_groupi_n_1125 ,csa_tree_add_7_27_groupi_n_862 ,csa_tree_add_7_27_groupi_n_916);
  nor csa_tree_add_7_27_groupi_g6059(csa_tree_add_7_27_groupi_n_1124 ,csa_tree_add_7_27_groupi_n_347 ,csa_tree_add_7_27_groupi_n_130);
  nor csa_tree_add_7_27_groupi_g6060(csa_tree_add_7_27_groupi_n_1123 ,csa_tree_add_7_27_groupi_n_250 ,csa_tree_add_7_27_groupi_n_175);
  nor csa_tree_add_7_27_groupi_g6061(csa_tree_add_7_27_groupi_n_1122 ,csa_tree_add_7_27_groupi_n_314 ,csa_tree_add_7_27_groupi_n_125);
  or csa_tree_add_7_27_groupi_g6062(csa_tree_add_7_27_groupi_n_1121 ,csa_tree_add_7_27_groupi_n_890 ,csa_tree_add_7_27_groupi_n_958);
  nor csa_tree_add_7_27_groupi_g6063(csa_tree_add_7_27_groupi_n_1120 ,csa_tree_add_7_27_groupi_n_296 ,csa_tree_add_7_27_groupi_n_124);
  or csa_tree_add_7_27_groupi_g6064(csa_tree_add_7_27_groupi_n_1119 ,csa_tree_add_7_27_groupi_n_884 ,csa_tree_add_7_27_groupi_n_953);
  or csa_tree_add_7_27_groupi_g6065(csa_tree_add_7_27_groupi_n_1118 ,csa_tree_add_7_27_groupi_n_859 ,csa_tree_add_7_27_groupi_n_949);
  or csa_tree_add_7_27_groupi_g6066(csa_tree_add_7_27_groupi_n_1117 ,csa_tree_add_7_27_groupi_n_861 ,csa_tree_add_7_27_groupi_n_960);
  nor csa_tree_add_7_27_groupi_g6067(csa_tree_add_7_27_groupi_n_1116 ,csa_tree_add_7_27_groupi_n_245 ,csa_tree_add_7_27_groupi_n_111);
  or csa_tree_add_7_27_groupi_g6068(csa_tree_add_7_27_groupi_n_1115 ,csa_tree_add_7_27_groupi_n_767 ,csa_tree_add_7_27_groupi_n_970);
  nor csa_tree_add_7_27_groupi_g6069(csa_tree_add_7_27_groupi_n_1114 ,csa_tree_add_7_27_groupi_n_323 ,csa_tree_add_7_27_groupi_n_194);
  nor csa_tree_add_7_27_groupi_g6070(csa_tree_add_7_27_groupi_n_1113 ,csa_tree_add_7_27_groupi_n_365 ,csa_tree_add_7_27_groupi_n_143);
  nor csa_tree_add_7_27_groupi_g6071(csa_tree_add_7_27_groupi_n_1112 ,csa_tree_add_7_27_groupi_n_281 ,csa_tree_add_7_27_groupi_n_142);
  nor csa_tree_add_7_27_groupi_g6072(csa_tree_add_7_27_groupi_n_1111 ,csa_tree_add_7_27_groupi_n_290 ,csa_tree_add_7_27_groupi_n_178);
  or csa_tree_add_7_27_groupi_g6073(csa_tree_add_7_27_groupi_n_1110 ,csa_tree_add_7_27_groupi_n_878 ,csa_tree_add_7_27_groupi_n_951);
  nor csa_tree_add_7_27_groupi_g6074(csa_tree_add_7_27_groupi_n_1109 ,csa_tree_add_7_27_groupi_n_375 ,csa_tree_add_7_27_groupi_n_193);
  nor csa_tree_add_7_27_groupi_g6075(csa_tree_add_7_27_groupi_n_1108 ,csa_tree_add_7_27_groupi_n_71 ,csa_tree_add_7_27_groupi_n_145);
  nor csa_tree_add_7_27_groupi_g6076(csa_tree_add_7_27_groupi_n_1107 ,csa_tree_add_7_27_groupi_n_254 ,csa_tree_add_7_27_groupi_n_119);
  nor csa_tree_add_7_27_groupi_g6077(csa_tree_add_7_27_groupi_n_1106 ,csa_tree_add_7_27_groupi_n_68 ,csa_tree_add_7_27_groupi_n_118);
  nor csa_tree_add_7_27_groupi_g6078(csa_tree_add_7_27_groupi_n_1105 ,csa_tree_add_7_27_groupi_n_341 ,csa_tree_add_7_27_groupi_n_146);
  nor csa_tree_add_7_27_groupi_g6079(csa_tree_add_7_27_groupi_n_1104 ,csa_tree_add_7_27_groupi_n_302 ,csa_tree_add_7_27_groupi_n_145);
  nor csa_tree_add_7_27_groupi_g6080(csa_tree_add_7_27_groupi_n_1103 ,csa_tree_add_7_27_groupi_n_353 ,csa_tree_add_7_27_groupi_n_160);
  nor csa_tree_add_7_27_groupi_g6081(csa_tree_add_7_27_groupi_n_1102 ,csa_tree_add_7_27_groupi_n_335 ,csa_tree_add_7_27_groupi_n_161);
  nor csa_tree_add_7_27_groupi_g6082(csa_tree_add_7_27_groupi_n_1101 ,csa_tree_add_7_27_groupi_n_53 ,csa_tree_add_7_27_groupi_n_161);
  nor csa_tree_add_7_27_groupi_g6083(csa_tree_add_7_27_groupi_n_1100 ,csa_tree_add_7_27_groupi_n_332 ,csa_tree_add_7_27_groupi_n_119);
  nor csa_tree_add_7_27_groupi_g6084(csa_tree_add_7_27_groupi_n_1099 ,csa_tree_add_7_27_groupi_n_369 ,csa_tree_add_7_27_groupi_n_160);
  nor csa_tree_add_7_27_groupi_g6085(csa_tree_add_7_27_groupi_n_1098 ,csa_tree_add_7_27_groupi_n_50 ,csa_tree_add_7_27_groupi_n_229);
  nor csa_tree_add_7_27_groupi_g6086(csa_tree_add_7_27_groupi_n_1097 ,csa_tree_add_7_27_groupi_n_78 ,csa_tree_add_7_27_groupi_n_229);
  nor csa_tree_add_7_27_groupi_g6087(csa_tree_add_7_27_groupi_n_1096 ,csa_tree_add_7_27_groupi_n_266 ,csa_tree_add_7_27_groupi_n_230);
  nor csa_tree_add_7_27_groupi_g6088(csa_tree_add_7_27_groupi_n_1095 ,csa_tree_add_7_27_groupi_n_257 ,csa_tree_add_7_27_groupi_n_179);
  nor csa_tree_add_7_27_groupi_g6089(csa_tree_add_7_27_groupi_n_1094 ,csa_tree_add_7_27_groupi_n_58 ,csa_tree_add_7_27_groupi_n_179);
  nor csa_tree_add_7_27_groupi_g6090(csa_tree_add_7_27_groupi_n_1093 ,csa_tree_add_7_27_groupi_n_389 ,csa_tree_add_7_27_groupi_n_131);
  nor csa_tree_add_7_27_groupi_g6091(csa_tree_add_7_27_groupi_n_1092 ,csa_tree_add_7_27_groupi_n_37 ,csa_tree_add_7_27_groupi_n_178);
  nor csa_tree_add_7_27_groupi_g6092(csa_tree_add_7_27_groupi_n_1091 ,csa_tree_add_7_27_groupi_n_44 ,csa_tree_add_7_27_groupi_n_214);
  nor csa_tree_add_7_27_groupi_g6093(csa_tree_add_7_27_groupi_n_1090 ,csa_tree_add_7_27_groupi_n_433 ,csa_tree_add_7_27_groupi_n_220);
  nor csa_tree_add_7_27_groupi_g6094(csa_tree_add_7_27_groupi_n_1089 ,csa_tree_add_7_27_groupi_n_28 ,csa_tree_add_7_27_groupi_n_221);
  nor csa_tree_add_7_27_groupi_g6095(csa_tree_add_7_27_groupi_n_1088 ,csa_tree_add_7_27_groupi_n_372 ,csa_tree_add_7_27_groupi_n_221);
  nor csa_tree_add_7_27_groupi_g6096(csa_tree_add_7_27_groupi_n_1087 ,csa_tree_add_7_27_groupi_n_421 ,csa_tree_add_7_27_groupi_n_128);
  nor csa_tree_add_7_27_groupi_g6097(csa_tree_add_7_27_groupi_n_1086 ,csa_tree_add_7_27_groupi_n_88 ,csa_tree_add_7_27_groupi_n_220);
  nor csa_tree_add_7_27_groupi_g6098(csa_tree_add_7_27_groupi_n_1085 ,csa_tree_add_7_27_groupi_n_401 ,csa_tree_add_7_27_groupi_n_181);
  nor csa_tree_add_7_27_groupi_g6099(csa_tree_add_7_27_groupi_n_1084 ,csa_tree_add_7_27_groupi_n_413 ,csa_tree_add_7_27_groupi_n_169);
  nor csa_tree_add_7_27_groupi_g6100(csa_tree_add_7_27_groupi_n_1083 ,csa_tree_add_7_27_groupi_n_31 ,csa_tree_add_7_27_groupi_n_182);
  nor csa_tree_add_7_27_groupi_g6101(csa_tree_add_7_27_groupi_n_1082 ,csa_tree_add_7_27_groupi_n_263 ,csa_tree_add_7_27_groupi_n_214);
  nor csa_tree_add_7_27_groupi_g6102(csa_tree_add_7_27_groupi_n_1081 ,csa_tree_add_7_27_groupi_n_447 ,csa_tree_add_7_27_groupi_n_182);
  nor csa_tree_add_7_27_groupi_g6103(csa_tree_add_7_27_groupi_n_1080 ,csa_tree_add_7_27_groupi_n_444 ,csa_tree_add_7_27_groupi_n_125);
  nor csa_tree_add_7_27_groupi_g6104(csa_tree_add_7_27_groupi_n_1079 ,csa_tree_add_7_27_groupi_n_320 ,csa_tree_add_7_27_groupi_n_169);
  nor csa_tree_add_7_27_groupi_g6105(csa_tree_add_7_27_groupi_n_1078 ,csa_tree_add_7_27_groupi_n_428 ,csa_tree_add_7_27_groupi_n_215);
  nor csa_tree_add_7_27_groupi_g6106(csa_tree_add_7_27_groupi_n_1077 ,csa_tree_add_7_27_groupi_n_410 ,csa_tree_add_7_27_groupi_n_181);
  nor csa_tree_add_7_27_groupi_g6107(csa_tree_add_7_27_groupi_n_1076 ,csa_tree_add_7_27_groupi_n_85 ,csa_tree_add_7_27_groupi_n_196);
  and csa_tree_add_7_27_groupi_g6108(csa_tree_add_7_27_groupi_n_1174 ,csa_tree_add_7_27_groupi_n_875 ,csa_tree_add_7_27_groupi_n_924);
  or csa_tree_add_7_27_groupi_g6109(csa_tree_add_7_27_groupi_n_1173 ,csa_tree_add_7_27_groupi_n_898 ,csa_tree_add_7_27_groupi_n_930);
  or csa_tree_add_7_27_groupi_g6110(csa_tree_add_7_27_groupi_n_1172 ,csa_tree_add_7_27_groupi_n_854 ,csa_tree_add_7_27_groupi_n_918);
  or csa_tree_add_7_27_groupi_g6111(csa_tree_add_7_27_groupi_n_1171 ,csa_tree_add_7_27_groupi_n_886 ,csa_tree_add_7_27_groupi_n_926);
  or csa_tree_add_7_27_groupi_g6112(csa_tree_add_7_27_groupi_n_1170 ,csa_tree_add_7_27_groupi_n_879 ,csa_tree_add_7_27_groupi_n_917);
  or csa_tree_add_7_27_groupi_g6113(csa_tree_add_7_27_groupi_n_1169 ,csa_tree_add_7_27_groupi_n_883 ,csa_tree_add_7_27_groupi_n_927);
  and csa_tree_add_7_27_groupi_g6114(csa_tree_add_7_27_groupi_n_1168 ,in3[15] ,csa_tree_add_7_27_groupi_n_969);
  or csa_tree_add_7_27_groupi_g6115(csa_tree_add_7_27_groupi_n_1167 ,csa_tree_add_7_27_groupi_n_857 ,csa_tree_add_7_27_groupi_n_931);
  or csa_tree_add_7_27_groupi_g6116(csa_tree_add_7_27_groupi_n_1166 ,csa_tree_add_7_27_groupi_n_855 ,csa_tree_add_7_27_groupi_n_925);
  or csa_tree_add_7_27_groupi_g6117(csa_tree_add_7_27_groupi_n_1164 ,csa_tree_add_7_27_groupi_n_876 ,csa_tree_add_7_27_groupi_n_923);
  or csa_tree_add_7_27_groupi_g6118(csa_tree_add_7_27_groupi_n_1162 ,csa_tree_add_7_27_groupi_n_882 ,csa_tree_add_7_27_groupi_n_920);
  or csa_tree_add_7_27_groupi_g6119(csa_tree_add_7_27_groupi_n_1161 ,csa_tree_add_7_27_groupi_n_874 ,csa_tree_add_7_27_groupi_n_929);
  or csa_tree_add_7_27_groupi_g6120(csa_tree_add_7_27_groupi_n_1159 ,csa_tree_add_7_27_groupi_n_853 ,csa_tree_add_7_27_groupi_n_928);
  or csa_tree_add_7_27_groupi_g6121(csa_tree_add_7_27_groupi_n_1157 ,csa_tree_add_7_27_groupi_n_849 ,csa_tree_add_7_27_groupi_n_921);
  or csa_tree_add_7_27_groupi_g6122(csa_tree_add_7_27_groupi_n_1156 ,csa_tree_add_7_27_groupi_n_860 ,csa_tree_add_7_27_groupi_n_919);
  or csa_tree_add_7_27_groupi_g6123(csa_tree_add_7_27_groupi_n_1153 ,csa_tree_add_7_27_groupi_n_848 ,csa_tree_add_7_27_groupi_n_922);
  not csa_tree_add_7_27_groupi_g6124(csa_tree_add_7_27_groupi_n_1074 ,csa_tree_add_7_27_groupi_n_1073);
  not csa_tree_add_7_27_groupi_g6125(csa_tree_add_7_27_groupi_n_1072 ,csa_tree_add_7_27_groupi_n_491);
  not csa_tree_add_7_27_groupi_g6127(csa_tree_add_7_27_groupi_n_1071 ,csa_tree_add_7_27_groupi_n_1073);
  not csa_tree_add_7_27_groupi_g6128(csa_tree_add_7_27_groupi_n_1070 ,csa_tree_add_7_27_groupi_n_1069);
  not csa_tree_add_7_27_groupi_g6129(csa_tree_add_7_27_groupi_n_1068 ,csa_tree_add_7_27_groupi_n_494);
  not csa_tree_add_7_27_groupi_g6131(csa_tree_add_7_27_groupi_n_1067 ,csa_tree_add_7_27_groupi_n_1069);
  not csa_tree_add_7_27_groupi_g6132(csa_tree_add_7_27_groupi_n_1066 ,csa_tree_add_7_27_groupi_n_1065);
  not csa_tree_add_7_27_groupi_g6133(csa_tree_add_7_27_groupi_n_1064 ,csa_tree_add_7_27_groupi_n_492);
  not csa_tree_add_7_27_groupi_g6135(csa_tree_add_7_27_groupi_n_1063 ,csa_tree_add_7_27_groupi_n_1065);
  not csa_tree_add_7_27_groupi_g6136(csa_tree_add_7_27_groupi_n_1062 ,csa_tree_add_7_27_groupi_n_1061);
  not csa_tree_add_7_27_groupi_g6137(csa_tree_add_7_27_groupi_n_1060 ,csa_tree_add_7_27_groupi_n_493);
  not csa_tree_add_7_27_groupi_g6139(csa_tree_add_7_27_groupi_n_1059 ,csa_tree_add_7_27_groupi_n_1061);
  nor csa_tree_add_7_27_groupi_g6140(csa_tree_add_7_27_groupi_n_1058 ,csa_tree_add_7_27_groupi_n_398 ,csa_tree_add_7_27_groupi_n_224);
  nor csa_tree_add_7_27_groupi_g6141(csa_tree_add_7_27_groupi_n_1057 ,csa_tree_add_7_27_groupi_n_262 ,csa_tree_add_7_27_groupi_n_170);
  nor csa_tree_add_7_27_groupi_g6142(csa_tree_add_7_27_groupi_n_1056 ,csa_tree_add_7_27_groupi_n_361 ,csa_tree_add_7_27_groupi_n_155);
  nor csa_tree_add_7_27_groupi_g6143(csa_tree_add_7_27_groupi_n_1055 ,csa_tree_add_7_27_groupi_n_361 ,csa_tree_add_7_27_groupi_n_238);
  nor csa_tree_add_7_27_groupi_g6144(csa_tree_add_7_27_groupi_n_1054 ,csa_tree_add_7_27_groupi_n_451 ,csa_tree_add_7_27_groupi_n_188);
  nor csa_tree_add_7_27_groupi_g6145(csa_tree_add_7_27_groupi_n_1053 ,csa_tree_add_7_27_groupi_n_250 ,csa_tree_add_7_27_groupi_n_241);
  nor csa_tree_add_7_27_groupi_g6146(csa_tree_add_7_27_groupi_n_1052 ,csa_tree_add_7_27_groupi_n_374 ,csa_tree_add_7_27_groupi_n_218);
  nor csa_tree_add_7_27_groupi_g6147(csa_tree_add_7_27_groupi_n_1051 ,csa_tree_add_7_27_groupi_n_337 ,csa_tree_add_7_27_groupi_n_209);
  nor csa_tree_add_7_27_groupi_g6148(csa_tree_add_7_27_groupi_n_1050 ,csa_tree_add_7_27_groupi_n_350 ,csa_tree_add_7_27_groupi_n_203);
  nor csa_tree_add_7_27_groupi_g6149(csa_tree_add_7_27_groupi_n_1049 ,csa_tree_add_7_27_groupi_n_377 ,csa_tree_add_7_27_groupi_n_244);
  nor csa_tree_add_7_27_groupi_g6150(csa_tree_add_7_27_groupi_n_1048 ,csa_tree_add_7_27_groupi_n_367 ,csa_tree_add_7_27_groupi_n_212);
  nor csa_tree_add_7_27_groupi_g6151(csa_tree_add_7_27_groupi_n_1047 ,csa_tree_add_7_27_groupi_n_251 ,csa_tree_add_7_27_groupi_n_247);
  nor csa_tree_add_7_27_groupi_g6152(csa_tree_add_7_27_groupi_n_1046 ,csa_tree_add_7_27_groupi_n_331 ,csa_tree_add_7_27_groupi_n_200);
  nor csa_tree_add_7_27_groupi_g6153(csa_tree_add_7_27_groupi_n_1045 ,csa_tree_add_7_27_groupi_n_262 ,csa_tree_add_7_27_groupi_n_167);
  nor csa_tree_add_7_27_groupi_g6154(csa_tree_add_7_27_groupi_n_1044 ,csa_tree_add_7_27_groupi_n_383 ,csa_tree_add_7_27_groupi_n_211);
  nor csa_tree_add_7_27_groupi_g6155(csa_tree_add_7_27_groupi_n_1043 ,csa_tree_add_7_27_groupi_n_56 ,csa_tree_add_7_27_groupi_n_134);
  nor csa_tree_add_7_27_groupi_g6156(csa_tree_add_7_27_groupi_n_1042 ,csa_tree_add_7_27_groupi_n_334 ,csa_tree_add_7_27_groupi_n_199);
  nor csa_tree_add_7_27_groupi_g6157(csa_tree_add_7_27_groupi_n_1041 ,csa_tree_add_7_27_groupi_n_393 ,csa_tree_add_7_27_groupi_n_227);
  nor csa_tree_add_7_27_groupi_g6158(csa_tree_add_7_27_groupi_n_1040 ,csa_tree_add_7_27_groupi_n_313 ,csa_tree_add_7_27_groupi_n_158);
  nor csa_tree_add_7_27_groupi_g6159(csa_tree_add_7_27_groupi_n_1039 ,csa_tree_add_7_27_groupi_n_265 ,csa_tree_add_7_27_groupi_n_166);
  nor csa_tree_add_7_27_groupi_g6160(csa_tree_add_7_27_groupi_n_1038 ,csa_tree_add_7_27_groupi_n_301 ,csa_tree_add_7_27_groupi_n_226);
  nor csa_tree_add_7_27_groupi_g6161(csa_tree_add_7_27_groupi_n_1037 ,csa_tree_add_7_27_groupi_n_352 ,csa_tree_add_7_27_groupi_n_187);
  nor csa_tree_add_7_27_groupi_g6162(csa_tree_add_7_27_groupi_n_1036 ,csa_tree_add_7_27_groupi_n_390 ,csa_tree_add_7_27_groupi_n_248);
  nor csa_tree_add_7_27_groupi_g6163(csa_tree_add_7_27_groupi_n_1035 ,csa_tree_add_7_27_groupi_n_280 ,csa_tree_add_7_27_groupi_n_157);
  nor csa_tree_add_7_27_groupi_g6164(csa_tree_add_7_27_groupi_n_1034 ,csa_tree_add_7_27_groupi_n_256 ,csa_tree_add_7_27_groupi_n_133);
  nor csa_tree_add_7_27_groupi_g6165(csa_tree_add_7_27_groupi_n_1033 ,csa_tree_add_7_27_groupi_n_387 ,csa_tree_add_7_27_groupi_n_122);
  nor csa_tree_add_7_27_groupi_g6166(csa_tree_add_7_27_groupi_n_1032 ,csa_tree_add_7_27_groupi_n_331 ,csa_tree_add_7_27_groupi_n_239);
  nor csa_tree_add_7_27_groupi_g6167(csa_tree_add_7_27_groupi_n_1031 ,csa_tree_add_7_27_groupi_n_256 ,csa_tree_add_7_27_groupi_n_227);
  nor csa_tree_add_7_27_groupi_g6168(csa_tree_add_7_27_groupi_n_1030 ,csa_tree_add_7_27_groupi_n_265 ,csa_tree_add_7_27_groupi_n_191);
  nor csa_tree_add_7_27_groupi_g6169(csa_tree_add_7_27_groupi_n_1029 ,csa_tree_add_7_27_groupi_n_301 ,csa_tree_add_7_27_groupi_n_121);
  nor csa_tree_add_7_27_groupi_g6170(csa_tree_add_7_27_groupi_n_1028 ,csa_tree_add_7_27_groupi_n_319 ,csa_tree_add_7_27_groupi_n_206);
  nor csa_tree_add_7_27_groupi_g6171(csa_tree_add_7_27_groupi_n_1027 ,csa_tree_add_7_27_groupi_n_385 ,csa_tree_add_7_27_groupi_n_188);
  nor csa_tree_add_7_27_groupi_g6172(csa_tree_add_7_27_groupi_n_1026 ,csa_tree_add_7_27_groupi_n_313 ,csa_tree_add_7_27_groupi_n_190);
  nor csa_tree_add_7_27_groupi_g6173(csa_tree_add_7_27_groupi_n_1025 ,csa_tree_add_7_27_groupi_n_292 ,csa_tree_add_7_27_groupi_n_158);
  nor csa_tree_add_7_27_groupi_g6174(csa_tree_add_7_27_groupi_n_1024 ,csa_tree_add_7_27_groupi_n_292 ,csa_tree_add_7_27_groupi_n_245);
  nor csa_tree_add_7_27_groupi_g6175(csa_tree_add_7_27_groupi_n_1023 ,csa_tree_add_7_27_groupi_n_397 ,csa_tree_add_7_27_groupi_n_191);
  nor csa_tree_add_7_27_groupi_g6176(csa_tree_add_7_27_groupi_n_1022 ,csa_tree_add_7_27_groupi_n_430 ,csa_tree_add_7_27_groupi_n_205);
  nor csa_tree_add_7_27_groupi_g6177(csa_tree_add_7_27_groupi_n_1021 ,csa_tree_add_7_27_groupi_n_352 ,csa_tree_add_7_27_groupi_n_247);
  nor csa_tree_add_7_27_groupi_g6178(csa_tree_add_7_27_groupi_n_1020 ,csa_tree_add_7_27_groupi_n_334 ,csa_tree_add_7_27_groupi_n_244);
  nor csa_tree_add_7_27_groupi_g6179(csa_tree_add_7_27_groupi_n_1019 ,csa_tree_add_7_27_groupi_n_403 ,csa_tree_add_7_27_groupi_n_187);
  nor csa_tree_add_7_27_groupi_g6180(csa_tree_add_7_27_groupi_n_1018 ,csa_tree_add_7_27_groupi_n_280 ,csa_tree_add_7_27_groupi_n_200);
  nor csa_tree_add_7_27_groupi_g6181(csa_tree_add_7_27_groupi_n_1017 ,csa_tree_add_7_27_groupi_n_415 ,csa_tree_add_7_27_groupi_n_238);
  nor csa_tree_add_7_27_groupi_g6182(csa_tree_add_7_27_groupi_n_1016 ,csa_tree_add_7_27_groupi_n_420 ,csa_tree_add_7_27_groupi_n_242);
  nor csa_tree_add_7_27_groupi_g6183(csa_tree_add_7_27_groupi_n_1015 ,csa_tree_add_7_27_groupi_n_432 ,csa_tree_add_7_27_groupi_n_139);
  nor csa_tree_add_7_27_groupi_g6184(csa_tree_add_7_27_groupi_n_1014 ,csa_tree_add_7_27_groupi_n_392 ,csa_tree_add_7_27_groupi_n_196);
  nor csa_tree_add_7_27_groupi_g6185(csa_tree_add_7_27_groupi_n_1013 ,csa_tree_add_7_27_groupi_n_42 ,csa_tree_add_7_27_groupi_n_212);
  nor csa_tree_add_7_27_groupi_g6186(csa_tree_add_7_27_groupi_n_1012 ,csa_tree_add_7_27_groupi_n_289 ,csa_tree_add_7_27_groupi_n_226);
  nor csa_tree_add_7_27_groupi_g6187(csa_tree_add_7_27_groupi_n_1011 ,csa_tree_add_7_27_groupi_n_435 ,csa_tree_add_7_27_groupi_n_140);
  nor csa_tree_add_7_27_groupi_g6188(csa_tree_add_7_27_groupi_n_1010 ,csa_tree_add_7_27_groupi_n_289 ,csa_tree_add_7_27_groupi_n_157);
  nor csa_tree_add_7_27_groupi_g6189(csa_tree_add_7_27_groupi_n_1009 ,csa_tree_add_7_27_groupi_n_323 ,csa_tree_add_7_27_groupi_n_134);
  nor csa_tree_add_7_27_groupi_g6190(csa_tree_add_7_27_groupi_n_1008 ,csa_tree_add_7_27_groupi_n_409 ,csa_tree_add_7_27_groupi_n_206);
  nor csa_tree_add_7_27_groupi_g6191(csa_tree_add_7_27_groupi_n_1007 ,csa_tree_add_7_27_groupi_n_260 ,csa_tree_add_7_27_groupi_n_223);
  nor csa_tree_add_7_27_groupi_g6192(csa_tree_add_7_27_groupi_n_1006 ,csa_tree_add_7_27_groupi_n_395 ,csa_tree_add_7_27_groupi_n_140);
  nor csa_tree_add_7_27_groupi_g6193(csa_tree_add_7_27_groupi_n_1005 ,csa_tree_add_7_27_groupi_n_405 ,csa_tree_add_7_27_groupi_n_122);
  nor csa_tree_add_7_27_groupi_g6194(csa_tree_add_7_27_groupi_n_1004 ,csa_tree_add_7_27_groupi_n_296 ,csa_tree_add_7_27_groupi_n_190);
  nor csa_tree_add_7_27_groupi_g6195(csa_tree_add_7_27_groupi_n_1003 ,csa_tree_add_7_27_groupi_n_254 ,csa_tree_add_7_27_groupi_n_202);
  nor csa_tree_add_7_27_groupi_g6196(csa_tree_add_7_27_groupi_n_1002 ,csa_tree_add_7_27_groupi_n_287 ,csa_tree_add_7_27_groupi_n_202);
  nor csa_tree_add_7_27_groupi_g6197(csa_tree_add_7_27_groupi_n_1001 ,csa_tree_add_7_27_groupi_n_423 ,csa_tree_add_7_27_groupi_n_139);
  nor csa_tree_add_7_27_groupi_g6198(csa_tree_add_7_27_groupi_n_1000 ,csa_tree_add_7_27_groupi_n_441 ,csa_tree_add_7_27_groupi_n_241);
  nor csa_tree_add_7_27_groupi_g6199(csa_tree_add_7_27_groupi_n_999 ,csa_tree_add_7_27_groupi_n_439 ,csa_tree_add_7_27_groupi_n_208);
  nor csa_tree_add_7_27_groupi_g6200(csa_tree_add_7_27_groupi_n_998 ,csa_tree_add_7_27_groupi_n_427 ,csa_tree_add_7_27_groupi_n_203);
  nor csa_tree_add_7_27_groupi_g6201(csa_tree_add_7_27_groupi_n_997 ,csa_tree_add_7_27_groupi_n_400 ,csa_tree_add_7_27_groupi_n_217);
  nor csa_tree_add_7_27_groupi_g6202(csa_tree_add_7_27_groupi_n_996 ,csa_tree_add_7_27_groupi_n_364 ,csa_tree_add_7_27_groupi_n_167);
  nor csa_tree_add_7_27_groupi_g6203(csa_tree_add_7_27_groupi_n_995 ,csa_tree_add_7_27_groupi_n_272 ,csa_tree_add_7_27_groupi_n_205);
  nor csa_tree_add_7_27_groupi_g6204(csa_tree_add_7_27_groupi_n_994 ,csa_tree_add_7_27_groupi_n_382 ,csa_tree_add_7_27_groupi_n_208);
  nor csa_tree_add_7_27_groupi_g6205(csa_tree_add_7_27_groupi_n_993 ,csa_tree_add_7_27_groupi_n_364 ,csa_tree_add_7_27_groupi_n_199);
  nor csa_tree_add_7_27_groupi_g6206(csa_tree_add_7_27_groupi_n_992 ,csa_tree_add_7_27_groupi_n_446 ,csa_tree_add_7_27_groupi_n_217);
  nor csa_tree_add_7_27_groupi_g6207(csa_tree_add_7_27_groupi_n_991 ,csa_tree_add_7_27_groupi_n_449 ,csa_tree_add_7_27_groupi_n_209);
  nor csa_tree_add_7_27_groupi_g6208(csa_tree_add_7_27_groupi_n_990 ,csa_tree_add_7_27_groupi_n_443 ,csa_tree_add_7_27_groupi_n_154);
  nor csa_tree_add_7_27_groupi_g6209(csa_tree_add_7_27_groupi_n_989 ,csa_tree_add_7_27_groupi_n_371 ,csa_tree_add_7_27_groupi_n_218);
  nor csa_tree_add_7_27_groupi_g6210(csa_tree_add_7_27_groupi_n_988 ,csa_tree_add_7_27_groupi_n_359 ,csa_tree_add_7_27_groupi_n_223);
  nor csa_tree_add_7_27_groupi_g6211(csa_tree_add_7_27_groupi_n_987 ,csa_tree_add_7_27_groupi_n_412 ,csa_tree_add_7_27_groupi_n_133);
  nor csa_tree_add_7_27_groupi_g6212(csa_tree_add_7_27_groupi_n_986 ,csa_tree_add_7_27_groupi_n_417 ,csa_tree_add_7_27_groupi_n_154);
  nor csa_tree_add_7_27_groupi_g6213(csa_tree_add_7_27_groupi_n_985 ,csa_tree_add_7_27_groupi_n_275 ,csa_tree_add_7_27_groupi_n_155);
  nor csa_tree_add_7_27_groupi_g6214(csa_tree_add_7_27_groupi_n_984 ,csa_tree_add_7_27_groupi_n_308 ,csa_tree_add_7_27_groupi_n_166);
  nor csa_tree_add_7_27_groupi_g6215(csa_tree_add_7_27_groupi_n_983 ,csa_tree_add_7_27_groupi_n_347 ,csa_tree_add_7_27_groupi_n_224);
  nor csa_tree_add_7_27_groupi_g6216(csa_tree_add_7_27_groupi_n_982 ,csa_tree_add_7_27_groupi_n_326 ,csa_tree_add_7_27_groupi_n_211);
  nor csa_tree_add_7_27_groupi_g6217(csa_tree_add_7_27_groupi_n_981 ,csa_tree_add_7_27_groupi_n_98 ,csa_tree_add_7_27_groupi_n_505);
  nor csa_tree_add_7_27_groupi_g6218(csa_tree_add_7_27_groupi_n_980 ,csa_tree_add_7_27_groupi_n_369 ,csa_tree_add_7_27_groupi_n_197);
  and csa_tree_add_7_27_groupi_g6219(csa_tree_add_7_27_groupi_n_979 ,csa_tree_add_7_27_groupi_n_66 ,csa_tree_add_7_27_groupi_n_130);
  and csa_tree_add_7_27_groupi_g6220(csa_tree_add_7_27_groupi_n_978 ,csa_tree_add_7_27_groupi_n_17 ,csa_tree_add_7_27_groupi_n_127);
  and csa_tree_add_7_27_groupi_g6221(csa_tree_add_7_27_groupi_n_977 ,csa_tree_add_7_27_groupi_n_48 ,csa_tree_add_7_27_groupi_n_124);
  nor csa_tree_add_7_27_groupi_g6222(csa_tree_add_7_27_groupi_n_976 ,csa_tree_add_7_27_groupi_n_106 ,csa_tree_add_7_27_groupi_n_866);
  nor csa_tree_add_7_27_groupi_g6223(csa_tree_add_7_27_groupi_n_975 ,csa_tree_add_7_27_groupi_n_100 ,csa_tree_add_7_27_groupi_n_506);
  nor csa_tree_add_7_27_groupi_g6224(csa_tree_add_7_27_groupi_n_974 ,csa_tree_add_7_27_groupi_n_104 ,csa_tree_add_7_27_groupi_n_866);
  nor csa_tree_add_7_27_groupi_g6225(csa_tree_add_7_27_groupi_n_973 ,csa_tree_add_7_27_groupi_n_102 ,csa_tree_add_7_27_groupi_n_506);
  and csa_tree_add_7_27_groupi_g6226(csa_tree_add_7_27_groupi_n_972 ,csa_tree_add_7_27_groupi_n_35 ,csa_tree_add_7_27_groupi_n_121);
  and csa_tree_add_7_27_groupi_g6227(csa_tree_add_7_27_groupi_n_971 ,csa_tree_add_7_27_groupi_n_94 ,csa_tree_add_7_27_groupi_n_118);
  xnor csa_tree_add_7_27_groupi_g6228(csa_tree_add_7_27_groupi_n_1075 ,csa_tree_add_7_27_groupi_n_790 ,csa_tree_add_7_27_groupi_n_835);
  or csa_tree_add_7_27_groupi_g6229(csa_tree_add_7_27_groupi_n_1073 ,csa_tree_add_7_27_groupi_n_947 ,csa_tree_add_7_27_groupi_n_946);
  or csa_tree_add_7_27_groupi_g6230(csa_tree_add_7_27_groupi_n_1069 ,csa_tree_add_7_27_groupi_n_934 ,csa_tree_add_7_27_groupi_n_952);
  or csa_tree_add_7_27_groupi_g6231(csa_tree_add_7_27_groupi_n_1065 ,csa_tree_add_7_27_groupi_n_944 ,csa_tree_add_7_27_groupi_n_933);
  or csa_tree_add_7_27_groupi_g6232(csa_tree_add_7_27_groupi_n_1061 ,csa_tree_add_7_27_groupi_n_962 ,csa_tree_add_7_27_groupi_n_948);
  nor csa_tree_add_7_27_groupi_g6234(csa_tree_add_7_27_groupi_n_962 ,csa_tree_add_7_27_groupi_n_743 ,csa_tree_add_7_27_groupi_n_903);
  nor csa_tree_add_7_27_groupi_g6235(csa_tree_add_7_27_groupi_n_961 ,csa_tree_add_7_27_groupi_n_290 ,csa_tree_add_7_27_groupi_n_164);
  nor csa_tree_add_7_27_groupi_g6236(csa_tree_add_7_27_groupi_n_960 ,csa_tree_add_7_27_groupi_n_302 ,csa_tree_add_7_27_groupi_n_149);
  nor csa_tree_add_7_27_groupi_g6237(csa_tree_add_7_27_groupi_n_959 ,csa_tree_add_7_27_groupi_n_335 ,csa_tree_add_7_27_groupi_n_235);
  nor csa_tree_add_7_27_groupi_g6238(csa_tree_add_7_27_groupi_n_958 ,csa_tree_add_7_27_groupi_n_332 ,csa_tree_add_7_27_groupi_n_173);
  nor csa_tree_add_7_27_groupi_g6239(csa_tree_add_7_27_groupi_n_957 ,csa_tree_add_7_27_groupi_n_337 ,csa_tree_add_7_27_groupi_n_172);
  nor csa_tree_add_7_27_groupi_g6240(csa_tree_add_7_27_groupi_n_956 ,csa_tree_add_7_27_groupi_n_362 ,csa_tree_add_7_27_groupi_n_164);
  nor csa_tree_add_7_27_groupi_g6241(csa_tree_add_7_27_groupi_n_955 ,csa_tree_add_7_27_groupi_n_257 ,csa_tree_add_7_27_groupi_n_163);
  nor csa_tree_add_7_27_groupi_g6242(csa_tree_add_7_27_groupi_n_954 ,csa_tree_add_7_27_groupi_n_293 ,csa_tree_add_7_27_groupi_n_236);
  nor csa_tree_add_7_27_groupi_g6243(csa_tree_add_7_27_groupi_n_953 ,csa_tree_add_7_27_groupi_n_236 ,csa_tree_add_7_27_groupi_n_566);
  and csa_tree_add_7_27_groupi_g6244(csa_tree_add_7_27_groupi_n_952 ,csa_tree_add_7_27_groupi_n_477 ,csa_tree_add_7_27_groupi_n_900);
  nor csa_tree_add_7_27_groupi_g6245(csa_tree_add_7_27_groupi_n_951 ,csa_tree_add_7_27_groupi_n_263 ,csa_tree_add_7_27_groupi_n_235);
  nor csa_tree_add_7_27_groupi_g6246(csa_tree_add_7_27_groupi_n_950 ,csa_tree_add_7_27_groupi_n_281 ,csa_tree_add_7_27_groupi_n_173);
  nor csa_tree_add_7_27_groupi_g6247(csa_tree_add_7_27_groupi_n_949 ,csa_tree_add_7_27_groupi_n_365 ,csa_tree_add_7_27_groupi_n_163);
  and csa_tree_add_7_27_groupi_g6248(csa_tree_add_7_27_groupi_n_948 ,csa_tree_add_7_27_groupi_n_480 ,csa_tree_add_7_27_groupi_n_904);
  nor csa_tree_add_7_27_groupi_g6249(csa_tree_add_7_27_groupi_n_947 ,csa_tree_add_7_27_groupi_n_745 ,csa_tree_add_7_27_groupi_n_901);
  and csa_tree_add_7_27_groupi_g6250(csa_tree_add_7_27_groupi_n_946 ,csa_tree_add_7_27_groupi_n_474 ,csa_tree_add_7_27_groupi_n_906);
  nor csa_tree_add_7_27_groupi_g6251(csa_tree_add_7_27_groupi_n_945 ,csa_tree_add_7_27_groupi_n_353 ,csa_tree_add_7_27_groupi_n_148);
  nor csa_tree_add_7_27_groupi_g6252(csa_tree_add_7_27_groupi_n_944 ,csa_tree_add_7_27_groupi_n_746 ,csa_tree_add_7_27_groupi_n_905);
  and csa_tree_add_7_27_groupi_g6253(csa_tree_add_7_27_groupi_n_970 ,csa_tree_add_7_27_groupi_n_780 ,csa_tree_add_7_27_groupi_n_895);
  and csa_tree_add_7_27_groupi_g6254(csa_tree_add_7_27_groupi_n_969 ,in1[0] ,csa_tree_add_7_27_groupi_n_560);
  and csa_tree_add_7_27_groupi_g6255(csa_tree_add_7_27_groupi_n_968 ,csa_tree_add_7_27_groupi_n_891 ,csa_tree_add_7_27_groupi_n_888);
  and csa_tree_add_7_27_groupi_g6256(csa_tree_add_7_27_groupi_n_967 ,csa_tree_add_7_27_groupi_n_897 ,csa_tree_add_7_27_groupi_n_889);
  or csa_tree_add_7_27_groupi_g6257(csa_tree_add_7_27_groupi_n_966 ,csa_tree_add_7_27_groupi_n_759 ,csa_tree_add_7_27_groupi_n_871);
  and csa_tree_add_7_27_groupi_g6258(csa_tree_add_7_27_groupi_n_965 ,csa_tree_add_7_27_groupi_n_892 ,csa_tree_add_7_27_groupi_n_887);
  and csa_tree_add_7_27_groupi_g6259(csa_tree_add_7_27_groupi_n_964 ,csa_tree_add_7_27_groupi_n_896 ,csa_tree_add_7_27_groupi_n_893);
  or csa_tree_add_7_27_groupi_g6260(csa_tree_add_7_27_groupi_n_963 ,csa_tree_add_7_27_groupi_n_759 ,csa_tree_add_7_27_groupi_n_872);
  nor csa_tree_add_7_27_groupi_g6261(csa_tree_add_7_27_groupi_n_935 ,csa_tree_add_7_27_groupi_n_341 ,csa_tree_add_7_27_groupi_n_148);
  nor csa_tree_add_7_27_groupi_g6262(csa_tree_add_7_27_groupi_n_934 ,csa_tree_add_7_27_groupi_n_744 ,csa_tree_add_7_27_groupi_n_902);
  and csa_tree_add_7_27_groupi_g6263(csa_tree_add_7_27_groupi_n_933 ,csa_tree_add_7_27_groupi_n_471 ,csa_tree_add_7_27_groupi_n_899);
  nor csa_tree_add_7_27_groupi_g6264(csa_tree_add_7_27_groupi_n_932 ,csa_tree_add_7_27_groupi_n_266 ,csa_tree_add_7_27_groupi_n_149);
  and csa_tree_add_7_27_groupi_g6265(csa_tree_add_7_27_groupi_n_931 ,in1[15] ,csa_tree_add_7_27_groupi_n_563);
  and csa_tree_add_7_27_groupi_g6266(csa_tree_add_7_27_groupi_n_930 ,in1[1] ,csa_tree_add_7_27_groupi_n_560);
  and csa_tree_add_7_27_groupi_g6267(csa_tree_add_7_27_groupi_n_929 ,in1[10] ,csa_tree_add_7_27_groupi_n_482);
  and csa_tree_add_7_27_groupi_g6268(csa_tree_add_7_27_groupi_n_928 ,in1[11] ,csa_tree_add_7_27_groupi_n_564);
  and csa_tree_add_7_27_groupi_g6269(csa_tree_add_7_27_groupi_n_927 ,in1[6] ,csa_tree_add_7_27_groupi_n_483);
  and csa_tree_add_7_27_groupi_g6270(csa_tree_add_7_27_groupi_n_926 ,in1[2] ,csa_tree_add_7_27_groupi_n_558);
  and csa_tree_add_7_27_groupi_g6271(csa_tree_add_7_27_groupi_n_925 ,in1[14] ,csa_tree_add_7_27_groupi_n_558);
  or csa_tree_add_7_27_groupi_g6272(csa_tree_add_7_27_groupi_n_924 ,csa_tree_add_7_27_groupi_n_32 ,csa_tree_add_7_27_groupi_n_863);
  and csa_tree_add_7_27_groupi_g6273(csa_tree_add_7_27_groupi_n_923 ,in1[7] ,csa_tree_add_7_27_groupi_n_563);
  and csa_tree_add_7_27_groupi_g6274(csa_tree_add_7_27_groupi_n_922 ,in1[13] ,csa_tree_add_7_27_groupi_n_557);
  and csa_tree_add_7_27_groupi_g6275(csa_tree_add_7_27_groupi_n_921 ,in1[4] ,csa_tree_add_7_27_groupi_n_483);
  and csa_tree_add_7_27_groupi_g6276(csa_tree_add_7_27_groupi_n_920 ,in1[8] ,csa_tree_add_7_27_groupi_n_561);
  and csa_tree_add_7_27_groupi_g6277(csa_tree_add_7_27_groupi_n_919 ,in1[5] ,csa_tree_add_7_27_groupi_n_561);
  and csa_tree_add_7_27_groupi_g6278(csa_tree_add_7_27_groupi_n_918 ,in1[9] ,csa_tree_add_7_27_groupi_n_557);
  and csa_tree_add_7_27_groupi_g6279(csa_tree_add_7_27_groupi_n_917 ,in1[12] ,csa_tree_add_7_27_groupi_n_564);
  nor csa_tree_add_7_27_groupi_g6280(csa_tree_add_7_27_groupi_n_916 ,csa_tree_add_7_27_groupi_n_314 ,csa_tree_add_7_27_groupi_n_172);
  or csa_tree_add_7_27_groupi_g6281(csa_tree_add_7_27_groupi_n_943 ,csa_tree_add_7_27_groupi_n_867 ,csa_tree_add_7_27_groupi_n_908);
  or csa_tree_add_7_27_groupi_g6282(csa_tree_add_7_27_groupi_n_942 ,csa_tree_add_7_27_groupi_n_869 ,csa_tree_add_7_27_groupi_n_910);
  or csa_tree_add_7_27_groupi_g6283(csa_tree_add_7_27_groupi_n_941 ,csa_tree_add_7_27_groupi_n_868 ,csa_tree_add_7_27_groupi_n_912);
  or csa_tree_add_7_27_groupi_g6284(csa_tree_add_7_27_groupi_n_940 ,csa_tree_add_7_27_groupi_n_870 ,csa_tree_add_7_27_groupi_n_914);
  or csa_tree_add_7_27_groupi_g6285(csa_tree_add_7_27_groupi_n_939 ,csa_tree_add_7_27_groupi_n_913 ,csa_tree_add_7_27_groupi_n_868);
  or csa_tree_add_7_27_groupi_g6286(csa_tree_add_7_27_groupi_n_938 ,csa_tree_add_7_27_groupi_n_915 ,csa_tree_add_7_27_groupi_n_870);
  or csa_tree_add_7_27_groupi_g6287(csa_tree_add_7_27_groupi_n_937 ,csa_tree_add_7_27_groupi_n_911 ,csa_tree_add_7_27_groupi_n_869);
  or csa_tree_add_7_27_groupi_g6288(csa_tree_add_7_27_groupi_n_936 ,csa_tree_add_7_27_groupi_n_909 ,csa_tree_add_7_27_groupi_n_867);
  not csa_tree_add_7_27_groupi_g6289(csa_tree_add_7_27_groupi_n_915 ,csa_tree_add_7_27_groupi_n_914);
  not csa_tree_add_7_27_groupi_g6290(csa_tree_add_7_27_groupi_n_913 ,csa_tree_add_7_27_groupi_n_912);
  not csa_tree_add_7_27_groupi_g6291(csa_tree_add_7_27_groupi_n_911 ,csa_tree_add_7_27_groupi_n_910);
  not csa_tree_add_7_27_groupi_g6292(csa_tree_add_7_27_groupi_n_909 ,csa_tree_add_7_27_groupi_n_908);
  nor csa_tree_add_7_27_groupi_g6293(csa_tree_add_7_27_groupi_n_906 ,in2[9] ,csa_tree_add_7_27_groupi_n_821);
  or csa_tree_add_7_27_groupi_g6294(csa_tree_add_7_27_groupi_n_905 ,csa_tree_add_7_27_groupi_n_739 ,csa_tree_add_7_27_groupi_n_822);
  nor csa_tree_add_7_27_groupi_g6295(csa_tree_add_7_27_groupi_n_904 ,in2[6] ,csa_tree_add_7_27_groupi_n_817);
  or csa_tree_add_7_27_groupi_g6296(csa_tree_add_7_27_groupi_n_903 ,csa_tree_add_7_27_groupi_n_755 ,csa_tree_add_7_27_groupi_n_814);
  or csa_tree_add_7_27_groupi_g6297(csa_tree_add_7_27_groupi_n_902 ,csa_tree_add_7_27_groupi_n_756 ,csa_tree_add_7_27_groupi_n_826);
  or csa_tree_add_7_27_groupi_g6298(csa_tree_add_7_27_groupi_n_901 ,csa_tree_add_7_27_groupi_n_740 ,csa_tree_add_7_27_groupi_n_818);
  nor csa_tree_add_7_27_groupi_g6299(csa_tree_add_7_27_groupi_n_900 ,in2[12] ,csa_tree_add_7_27_groupi_n_829);
  nor csa_tree_add_7_27_groupi_g6300(csa_tree_add_7_27_groupi_n_899 ,in2[3] ,csa_tree_add_7_27_groupi_n_825);
  nor csa_tree_add_7_27_groupi_g6301(csa_tree_add_7_27_groupi_n_898 ,csa_tree_add_7_27_groupi_n_116 ,csa_tree_add_7_27_groupi_n_719);
  or csa_tree_add_7_27_groupi_g6302(csa_tree_add_7_27_groupi_n_897 ,csa_tree_add_7_27_groupi_n_745 ,csa_tree_add_7_27_groupi_n_808);
  or csa_tree_add_7_27_groupi_g6303(csa_tree_add_7_27_groupi_n_896 ,csa_tree_add_7_27_groupi_n_743 ,csa_tree_add_7_27_groupi_n_800);
  nor csa_tree_add_7_27_groupi_g6305(csa_tree_add_7_27_groupi_n_894 ,csa_tree_add_7_27_groupi_n_233 ,csa_tree_add_7_27_groupi_n_567);
  or csa_tree_add_7_27_groupi_g6306(csa_tree_add_7_27_groupi_n_893 ,in2[5] ,csa_tree_add_7_27_groupi_n_802);
  or csa_tree_add_7_27_groupi_g6307(csa_tree_add_7_27_groupi_n_892 ,csa_tree_add_7_27_groupi_n_476 ,csa_tree_add_7_27_groupi_n_803);
  or csa_tree_add_7_27_groupi_g6308(csa_tree_add_7_27_groupi_n_891 ,csa_tree_add_7_27_groupi_n_746 ,csa_tree_add_7_27_groupi_n_804);
  nor csa_tree_add_7_27_groupi_g6309(csa_tree_add_7_27_groupi_n_890 ,csa_tree_add_7_27_groupi_n_72 ,csa_tree_add_7_27_groupi_n_152);
  or csa_tree_add_7_27_groupi_g6310(csa_tree_add_7_27_groupi_n_889 ,in2[8] ,csa_tree_add_7_27_groupi_n_805);
  or csa_tree_add_7_27_groupi_g6311(csa_tree_add_7_27_groupi_n_888 ,in2[2] ,csa_tree_add_7_27_groupi_n_806);
  or csa_tree_add_7_27_groupi_g6312(csa_tree_add_7_27_groupi_n_887 ,in2[11] ,csa_tree_add_7_27_groupi_n_807);
  nor csa_tree_add_7_27_groupi_g6313(csa_tree_add_7_27_groupi_n_886 ,csa_tree_add_7_27_groupi_n_20 ,csa_tree_add_7_27_groupi_n_718);
  nor csa_tree_add_7_27_groupi_g6314(csa_tree_add_7_27_groupi_n_885 ,csa_tree_add_7_27_groupi_n_96 ,csa_tree_add_7_27_groupi_n_232);
  nor csa_tree_add_7_27_groupi_g6315(csa_tree_add_7_27_groupi_n_884 ,csa_tree_add_7_27_groupi_n_13 ,csa_tree_add_7_27_groupi_n_137);
  nor csa_tree_add_7_27_groupi_g6316(csa_tree_add_7_27_groupi_n_883 ,csa_tree_add_7_27_groupi_n_51 ,csa_tree_add_7_27_groupi_n_716);
  nor csa_tree_add_7_27_groupi_g6317(csa_tree_add_7_27_groupi_n_882 ,csa_tree_add_7_27_groupi_n_86 ,csa_tree_add_7_27_groupi_n_718);
  nor csa_tree_add_7_27_groupi_g6318(csa_tree_add_7_27_groupi_n_881 ,csa_tree_add_7_27_groupi_n_32 ,csa_tree_add_7_27_groupi_n_136);
  nor csa_tree_add_7_27_groupi_g6319(csa_tree_add_7_27_groupi_n_880 ,csa_tree_add_7_27_groupi_n_319 ,csa_tree_add_7_27_groupi_n_185);
  nor csa_tree_add_7_27_groupi_g6320(csa_tree_add_7_27_groupi_n_879 ,csa_tree_add_7_27_groupi_n_29 ,csa_tree_add_7_27_groupi_n_674);
  nor csa_tree_add_7_27_groupi_g6321(csa_tree_add_7_27_groupi_n_878 ,csa_tree_add_7_27_groupi_n_45 ,csa_tree_add_7_27_groupi_n_184);
  nor csa_tree_add_7_27_groupi_g6322(csa_tree_add_7_27_groupi_n_877 ,csa_tree_add_7_27_groupi_n_22 ,csa_tree_add_7_27_groupi_n_233);
  nor csa_tree_add_7_27_groupi_g6323(csa_tree_add_7_27_groupi_n_876 ,csa_tree_add_7_27_groupi_n_59 ,csa_tree_add_7_27_groupi_n_673);
  or csa_tree_add_7_27_groupi_g6324(csa_tree_add_7_27_groupi_n_875 ,csa_tree_add_7_27_groupi_n_7 ,csa_tree_add_7_27_groupi_n_673);
  nor csa_tree_add_7_27_groupi_g6325(csa_tree_add_7_27_groupi_n_874 ,csa_tree_add_7_27_groupi_n_63 ,csa_tree_add_7_27_groupi_n_715);
  or csa_tree_add_7_27_groupi_g6326(csa_tree_add_7_27_groupi_n_914 ,csa_tree_add_7_27_groupi_n_815 ,csa_tree_add_7_27_groupi_n_816);
  or csa_tree_add_7_27_groupi_g6327(csa_tree_add_7_27_groupi_n_873 ,csa_tree_add_7_27_groupi_n_96 ,csa_tree_add_7_27_groupi_n_676);
  or csa_tree_add_7_27_groupi_g6328(csa_tree_add_7_27_groupi_n_912 ,csa_tree_add_7_27_groupi_n_819 ,csa_tree_add_7_27_groupi_n_820);
  or csa_tree_add_7_27_groupi_g6329(csa_tree_add_7_27_groupi_n_910 ,csa_tree_add_7_27_groupi_n_827 ,csa_tree_add_7_27_groupi_n_828);
  or csa_tree_add_7_27_groupi_g6330(csa_tree_add_7_27_groupi_n_908 ,csa_tree_add_7_27_groupi_n_823 ,csa_tree_add_7_27_groupi_n_824);
  or csa_tree_add_7_27_groupi_g6331(csa_tree_add_7_27_groupi_n_907 ,in2[0] ,csa_tree_add_7_27_groupi_n_791);
  not csa_tree_add_7_27_groupi_g6332(csa_tree_add_7_27_groupi_n_872 ,csa_tree_add_7_27_groupi_n_871);
  not csa_tree_add_7_27_groupi_g6333(csa_tree_add_7_27_groupi_n_865 ,csa_tree_add_7_27_groupi_n_863);
  not csa_tree_add_7_27_groupi_g6334(csa_tree_add_7_27_groupi_n_864 ,csa_tree_add_7_27_groupi_n_863);
  nor csa_tree_add_7_27_groupi_g6335(csa_tree_add_7_27_groupi_n_862 ,csa_tree_add_7_27_groupi_n_26 ,csa_tree_add_7_27_groupi_n_185);
  nor csa_tree_add_7_27_groupi_g6336(csa_tree_add_7_27_groupi_n_861 ,csa_tree_add_7_27_groupi_n_76 ,csa_tree_add_7_27_groupi_n_232);
  nor csa_tree_add_7_27_groupi_g6337(csa_tree_add_7_27_groupi_n_860 ,csa_tree_add_7_27_groupi_n_89 ,csa_tree_add_7_27_groupi_n_716);
  nor csa_tree_add_7_27_groupi_g6338(csa_tree_add_7_27_groupi_n_859 ,csa_tree_add_7_27_groupi_n_79 ,csa_tree_add_7_27_groupi_n_137);
  nor csa_tree_add_7_27_groupi_g6339(csa_tree_add_7_27_groupi_n_858 ,csa_tree_add_7_27_groupi_n_81 ,csa_tree_add_7_27_groupi_n_184);
  nor csa_tree_add_7_27_groupi_g6340(csa_tree_add_7_27_groupi_n_857 ,csa_tree_add_7_27_groupi_n_74 ,csa_tree_add_7_27_groupi_n_715);
  nor csa_tree_add_7_27_groupi_g6341(csa_tree_add_7_27_groupi_n_856 ,csa_tree_add_7_27_groupi_n_38 ,csa_tree_add_7_27_groupi_n_151);
  nor csa_tree_add_7_27_groupi_g6342(csa_tree_add_7_27_groupi_n_855 ,csa_tree_add_7_27_groupi_n_54 ,csa_tree_add_7_27_groupi_n_719);
  nor csa_tree_add_7_27_groupi_g6343(csa_tree_add_7_27_groupi_n_854 ,csa_tree_add_7_27_groupi_n_40 ,csa_tree_add_7_27_groupi_n_677);
  nor csa_tree_add_7_27_groupi_g6344(csa_tree_add_7_27_groupi_n_853 ,csa_tree_add_7_27_groupi_n_15 ,csa_tree_add_7_27_groupi_n_674);
  nor csa_tree_add_7_27_groupi_g6345(csa_tree_add_7_27_groupi_n_852 ,csa_tree_add_7_27_groupi_n_83 ,csa_tree_add_7_27_groupi_n_151);
  nor csa_tree_add_7_27_groupi_g6346(csa_tree_add_7_27_groupi_n_851 ,csa_tree_add_7_27_groupi_n_69 ,csa_tree_add_7_27_groupi_n_152);
  nor csa_tree_add_7_27_groupi_g6347(csa_tree_add_7_27_groupi_n_850 ,csa_tree_add_7_27_groupi_n_24 ,csa_tree_add_7_27_groupi_n_136);
  nor csa_tree_add_7_27_groupi_g6348(csa_tree_add_7_27_groupi_n_849 ,csa_tree_add_7_27_groupi_n_418 ,csa_tree_add_7_27_groupi_n_677);
  nor csa_tree_add_7_27_groupi_g6349(csa_tree_add_7_27_groupi_n_848 ,csa_tree_add_7_27_groupi_n_61 ,csa_tree_add_7_27_groupi_n_676);
  xnor csa_tree_add_7_27_groupi_g6350(csa_tree_add_7_27_groupi_n_847 ,in1[12] ,in1[11]);
  xnor csa_tree_add_7_27_groupi_g6351(csa_tree_add_7_27_groupi_n_846 ,in1[6] ,in1[5]);
  xnor csa_tree_add_7_27_groupi_g6352(csa_tree_add_7_27_groupi_n_871 ,csa_tree_add_7_27_groupi_n_471 ,in2[1]);
  xnor csa_tree_add_7_27_groupi_g6353(csa_tree_add_7_27_groupi_n_845 ,in2[8] ,in3[6]);
  xnor csa_tree_add_7_27_groupi_g6354(csa_tree_add_7_27_groupi_n_870 ,in2[6] ,in2[5]);
  xnor csa_tree_add_7_27_groupi_g6355(csa_tree_add_7_27_groupi_n_844 ,in2[11] ,in3[9]);
  xnor csa_tree_add_7_27_groupi_g6356(csa_tree_add_7_27_groupi_n_843 ,in2[5] ,in3[3]);
  xnor csa_tree_add_7_27_groupi_g6357(csa_tree_add_7_27_groupi_n_869 ,in2[12] ,in2[11]);
  xnor csa_tree_add_7_27_groupi_g6358(csa_tree_add_7_27_groupi_n_868 ,in2[9] ,in2[8]);
  xnor csa_tree_add_7_27_groupi_g6359(csa_tree_add_7_27_groupi_n_867 ,in2[3] ,in2[2]);
  xnor csa_tree_add_7_27_groupi_g6360(csa_tree_add_7_27_groupi_n_842 ,in2[14] ,in3[12]);
  xnor csa_tree_add_7_27_groupi_g6361(csa_tree_add_7_27_groupi_n_841 ,in1[3] ,in1[2]);
  xnor csa_tree_add_7_27_groupi_g6362(csa_tree_add_7_27_groupi_n_840 ,in1[14] ,in1[13]);
  xnor csa_tree_add_7_27_groupi_g6363(csa_tree_add_7_27_groupi_n_839 ,in1[7] ,in1[6]);
  xnor csa_tree_add_7_27_groupi_g6364(csa_tree_add_7_27_groupi_n_838 ,in1[9] ,in1[8]);
  xnor csa_tree_add_7_27_groupi_g6365(csa_tree_add_7_27_groupi_n_837 ,in1[11] ,in1[10]);
  xnor csa_tree_add_7_27_groupi_g6366(csa_tree_add_7_27_groupi_n_836 ,in1[15] ,in1[14]);
  xnor csa_tree_add_7_27_groupi_g6367(csa_tree_add_7_27_groupi_n_835 ,in1[2] ,in1[1]);
  xnor csa_tree_add_7_27_groupi_g6368(csa_tree_add_7_27_groupi_n_834 ,in1[13] ,in1[12]);
  xnor csa_tree_add_7_27_groupi_g6369(csa_tree_add_7_27_groupi_n_833 ,in1[4] ,in1[3]);
  xnor csa_tree_add_7_27_groupi_g6370(csa_tree_add_7_27_groupi_n_832 ,in1[8] ,in1[7]);
  xnor csa_tree_add_7_27_groupi_g6371(csa_tree_add_7_27_groupi_n_831 ,in1[5] ,in1[4]);
  xnor csa_tree_add_7_27_groupi_g6372(csa_tree_add_7_27_groupi_n_830 ,in1[10] ,in1[9]);
  xnor csa_tree_add_7_27_groupi_g6373(csa_tree_add_7_27_groupi_n_866 ,in1[1] ,in1[0]);
  or csa_tree_add_7_27_groupi_g6374(csa_tree_add_7_27_groupi_n_863 ,csa_tree_add_7_27_groupi_n_490 ,csa_tree_add_7_27_groupi_n_777);
  not csa_tree_add_7_27_groupi_g6375(csa_tree_add_7_27_groupi_n_829 ,csa_tree_add_7_27_groupi_n_828);
  not csa_tree_add_7_27_groupi_g6376(csa_tree_add_7_27_groupi_n_827 ,csa_tree_add_7_27_groupi_n_826);
  not csa_tree_add_7_27_groupi_g6377(csa_tree_add_7_27_groupi_n_825 ,csa_tree_add_7_27_groupi_n_824);
  not csa_tree_add_7_27_groupi_g6378(csa_tree_add_7_27_groupi_n_823 ,csa_tree_add_7_27_groupi_n_822);
  not csa_tree_add_7_27_groupi_g6379(csa_tree_add_7_27_groupi_n_821 ,csa_tree_add_7_27_groupi_n_820);
  not csa_tree_add_7_27_groupi_g6380(csa_tree_add_7_27_groupi_n_819 ,csa_tree_add_7_27_groupi_n_818);
  not csa_tree_add_7_27_groupi_g6381(csa_tree_add_7_27_groupi_n_817 ,csa_tree_add_7_27_groupi_n_816);
  not csa_tree_add_7_27_groupi_g6382(csa_tree_add_7_27_groupi_n_815 ,csa_tree_add_7_27_groupi_n_814);
  not csa_tree_add_7_27_groupi_g6383(csa_tree_add_7_27_groupi_n_812 ,csa_tree_add_7_27_groupi_n_490);
  not csa_tree_add_7_27_groupi_g6385(csa_tree_add_7_27_groupi_n_811 ,csa_tree_add_7_27_groupi_n_810);
  nor csa_tree_add_7_27_groupi_g6387(csa_tree_add_7_27_groupi_n_809 ,in1[12] ,in1[11]);
  or csa_tree_add_7_27_groupi_g6388(csa_tree_add_7_27_groupi_n_808 ,csa_tree_add_7_27_groupi_n_740 ,in2[10]);
  or csa_tree_add_7_27_groupi_g6389(csa_tree_add_7_27_groupi_n_807 ,csa_tree_add_7_27_groupi_n_758 ,in2[12]);
  or csa_tree_add_7_27_groupi_g6390(csa_tree_add_7_27_groupi_n_806 ,csa_tree_add_7_27_groupi_n_741 ,in2[3]);
  or csa_tree_add_7_27_groupi_g6391(csa_tree_add_7_27_groupi_n_805 ,csa_tree_add_7_27_groupi_n_757 ,in2[9]);
  or csa_tree_add_7_27_groupi_g6392(csa_tree_add_7_27_groupi_n_804 ,csa_tree_add_7_27_groupi_n_739 ,in2[4]);
  or csa_tree_add_7_27_groupi_g6393(csa_tree_add_7_27_groupi_n_803 ,csa_tree_add_7_27_groupi_n_756 ,in2[13]);
  or csa_tree_add_7_27_groupi_g6394(csa_tree_add_7_27_groupi_n_802 ,csa_tree_add_7_27_groupi_n_760 ,in2[6]);
  and csa_tree_add_7_27_groupi_g6395(csa_tree_add_7_27_groupi_n_801 ,in2[5] ,in3[3]);
  or csa_tree_add_7_27_groupi_g6396(csa_tree_add_7_27_groupi_n_800 ,csa_tree_add_7_27_groupi_n_755 ,in2[7]);
  nor csa_tree_add_7_27_groupi_g6397(csa_tree_add_7_27_groupi_n_799 ,in1[9] ,in1[8]);
  or csa_tree_add_7_27_groupi_g6398(csa_tree_add_7_27_groupi_n_798 ,csa_tree_add_7_27_groupi_n_29 ,csa_tree_add_7_27_groupi_n_38);
  nor csa_tree_add_7_27_groupi_g6399(csa_tree_add_7_27_groupi_n_797 ,in1[4] ,in1[3]);
  or csa_tree_add_7_27_groupi_g6400(csa_tree_add_7_27_groupi_n_796 ,csa_tree_add_7_27_groupi_n_54 ,csa_tree_add_7_27_groupi_n_69);
  nor csa_tree_add_7_27_groupi_g6401(csa_tree_add_7_27_groupi_n_795 ,in1[10] ,in1[9]);
  nor csa_tree_add_7_27_groupi_g6403(csa_tree_add_7_27_groupi_n_793 ,in1[14] ,in1[13]);
  or csa_tree_add_7_27_groupi_g6404(csa_tree_add_7_27_groupi_n_792 ,csa_tree_add_7_27_groupi_n_79 ,csa_tree_add_7_27_groupi_n_83);
  and csa_tree_add_7_27_groupi_g6405(csa_tree_add_7_27_groupi_n_828 ,in2[14] ,csa_tree_add_7_27_groupi_n_758);
  or csa_tree_add_7_27_groupi_g6406(csa_tree_add_7_27_groupi_n_826 ,csa_tree_add_7_27_groupi_n_758 ,in2[14]);
  or csa_tree_add_7_27_groupi_g6407(csa_tree_add_7_27_groupi_n_791 ,csa_tree_add_7_27_groupi_n_470 ,in2[1]);
  and csa_tree_add_7_27_groupi_g6408(csa_tree_add_7_27_groupi_n_824 ,in2[5] ,csa_tree_add_7_27_groupi_n_741);
  or csa_tree_add_7_27_groupi_g6409(csa_tree_add_7_27_groupi_n_822 ,csa_tree_add_7_27_groupi_n_741 ,in2[5]);
  and csa_tree_add_7_27_groupi_g6410(csa_tree_add_7_27_groupi_n_820 ,in2[11] ,csa_tree_add_7_27_groupi_n_757);
  or csa_tree_add_7_27_groupi_g6411(csa_tree_add_7_27_groupi_n_818 ,csa_tree_add_7_27_groupi_n_757 ,in2[11]);
  and csa_tree_add_7_27_groupi_g6412(csa_tree_add_7_27_groupi_n_816 ,in2[8] ,csa_tree_add_7_27_groupi_n_760);
  or csa_tree_add_7_27_groupi_g6413(csa_tree_add_7_27_groupi_n_814 ,csa_tree_add_7_27_groupi_n_760 ,in2[8]);
  or csa_tree_add_7_27_groupi_g6414(csa_tree_add_7_27_groupi_n_813 ,csa_tree_add_7_27_groupi_n_742 ,in2[0]);
  and csa_tree_add_7_27_groupi_g6415(csa_tree_add_7_27_groupi_n_810 ,in2[15] ,in2[14]);
  or csa_tree_add_7_27_groupi_g6416(csa_tree_add_7_27_groupi_n_789 ,in2[5] ,in3[3]);
  or csa_tree_add_7_27_groupi_g6417(csa_tree_add_7_27_groupi_n_788 ,csa_tree_add_7_27_groupi_n_42 ,csa_tree_add_7_27_groupi_n_91);
  or csa_tree_add_7_27_groupi_g6418(csa_tree_add_7_27_groupi_n_787 ,csa_tree_add_7_27_groupi_n_72 ,csa_tree_add_7_27_groupi_n_45);
  or csa_tree_add_7_27_groupi_g6419(csa_tree_add_7_27_groupi_n_786 ,in2[11] ,in3[9]);
  nor csa_tree_add_7_27_groupi_g6420(csa_tree_add_7_27_groupi_n_785 ,in1[13] ,in1[12]);
  nor csa_tree_add_7_27_groupi_g6421(csa_tree_add_7_27_groupi_n_784 ,in1[7] ,in1[6]);
  nor csa_tree_add_7_27_groupi_g6422(csa_tree_add_7_27_groupi_n_783 ,in1[11] ,in1[10]);
  nor csa_tree_add_7_27_groupi_g6423(csa_tree_add_7_27_groupi_n_782 ,in1[15] ,in1[14]);
  or csa_tree_add_7_27_groupi_g6424(csa_tree_add_7_27_groupi_n_781 ,csa_tree_add_7_27_groupi_n_89 ,csa_tree_add_7_27_groupi_n_56);
  or csa_tree_add_7_27_groupi_g6425(csa_tree_add_7_27_groupi_n_780 ,csa_tree_add_7_27_groupi_n_7 ,csa_tree_add_7_27_groupi_n_20);
  or csa_tree_add_7_27_groupi_g6426(csa_tree_add_7_27_groupi_n_779 ,csa_tree_add_7_27_groupi_n_86 ,csa_tree_add_7_27_groupi_n_59);
  or csa_tree_add_7_27_groupi_g6427(csa_tree_add_7_27_groupi_n_778 ,csa_tree_add_7_27_groupi_n_26 ,csa_tree_add_7_27_groupi_n_51);
  nor csa_tree_add_7_27_groupi_g6428(csa_tree_add_7_27_groupi_n_777 ,in2[15] ,in2[14]);
  or csa_tree_add_7_27_groupi_g6429(csa_tree_add_7_27_groupi_n_776 ,csa_tree_add_7_27_groupi_n_24 ,csa_tree_add_7_27_groupi_n_81);
  or csa_tree_add_7_27_groupi_g6430(csa_tree_add_7_27_groupi_n_775 ,in2[2] ,in3[0]);
  and csa_tree_add_7_27_groupi_g6431(csa_tree_add_7_27_groupi_n_774 ,in2[2] ,in3[0]);
  or csa_tree_add_7_27_groupi_g6432(csa_tree_add_7_27_groupi_n_773 ,csa_tree_add_7_27_groupi_n_10 ,csa_tree_add_7_27_groupi_n_74);
  or csa_tree_add_7_27_groupi_g6433(csa_tree_add_7_27_groupi_n_772 ,in2[8] ,in3[6]);
  nor csa_tree_add_7_27_groupi_g6434(csa_tree_add_7_27_groupi_n_771 ,in1[5] ,in1[4]);
  or csa_tree_add_7_27_groupi_g6435(csa_tree_add_7_27_groupi_n_770 ,csa_tree_add_7_27_groupi_n_40 ,csa_tree_add_7_27_groupi_n_76);
  nor csa_tree_add_7_27_groupi_g6436(csa_tree_add_7_27_groupi_n_769 ,in1[8] ,in1[7]);
  or csa_tree_add_7_27_groupi_g6437(csa_tree_add_7_27_groupi_n_768 ,csa_tree_add_7_27_groupi_n_15 ,csa_tree_add_7_27_groupi_n_63);
  nor csa_tree_add_7_27_groupi_g6438(csa_tree_add_7_27_groupi_n_767 ,in1[3] ,in1[2]);
  or csa_tree_add_7_27_groupi_g6439(csa_tree_add_7_27_groupi_n_766 ,csa_tree_add_7_27_groupi_n_61 ,csa_tree_add_7_27_groupi_n_22);
  and csa_tree_add_7_27_groupi_g6440(csa_tree_add_7_27_groupi_n_765 ,in2[8] ,in3[6]);
  or csa_tree_add_7_27_groupi_g6441(csa_tree_add_7_27_groupi_n_764 ,in2[14] ,in3[12]);
  and csa_tree_add_7_27_groupi_g6442(csa_tree_add_7_27_groupi_n_763 ,in2[14] ,in3[12]);
  nor csa_tree_add_7_27_groupi_g6443(csa_tree_add_7_27_groupi_n_762 ,in1[6] ,in1[5]);
  and csa_tree_add_7_27_groupi_g6444(csa_tree_add_7_27_groupi_n_761 ,in2[11] ,in3[9]);
  or csa_tree_add_7_27_groupi_g6445(csa_tree_add_7_27_groupi_n_790 ,csa_tree_add_7_27_groupi_n_13 ,csa_tree_add_7_27_groupi_n_115);
  not csa_tree_add_7_27_groupi_g6446(csa_tree_add_7_27_groupi_n_760 ,in2[7]);
  not csa_tree_add_7_27_groupi_g6447(csa_tree_add_7_27_groupi_n_759 ,in2[0]);
  not csa_tree_add_7_27_groupi_g6448(csa_tree_add_7_27_groupi_n_758 ,in2[13]);
  not csa_tree_add_7_27_groupi_g6449(csa_tree_add_7_27_groupi_n_757 ,in2[10]);
  not csa_tree_add_7_27_groupi_g6450(csa_tree_add_7_27_groupi_n_756 ,in2[12]);
  not csa_tree_add_7_27_groupi_g6451(csa_tree_add_7_27_groupi_n_755 ,in2[6]);
  not csa_tree_add_7_27_groupi_g6452(csa_tree_add_7_27_groupi_n_754 ,in1[0]);
  not csa_tree_add_7_27_groupi_g6453(csa_tree_add_7_27_groupi_n_753 ,in1[4]);
  not csa_tree_add_7_27_groupi_g6454(csa_tree_add_7_27_groupi_n_752 ,in1[12]);
  not csa_tree_add_7_27_groupi_g6455(csa_tree_add_7_27_groupi_n_751 ,in1[13]);
  not csa_tree_add_7_27_groupi_g6456(csa_tree_add_7_27_groupi_n_750 ,in1[11]);
  not csa_tree_add_7_27_groupi_g6457(csa_tree_add_7_27_groupi_n_749 ,in1[8]);
  not csa_tree_add_7_27_groupi_g6458(csa_tree_add_7_27_groupi_n_748 ,in1[3]);
  not csa_tree_add_7_27_groupi_g6459(csa_tree_add_7_27_groupi_n_747 ,in1[7]);
  not csa_tree_add_7_27_groupi_g6460(csa_tree_add_7_27_groupi_n_746 ,in2[2]);
  not csa_tree_add_7_27_groupi_g6461(csa_tree_add_7_27_groupi_n_745 ,in2[8]);
  not csa_tree_add_7_27_groupi_g6462(csa_tree_add_7_27_groupi_n_744 ,in2[11]);
  not csa_tree_add_7_27_groupi_g6463(csa_tree_add_7_27_groupi_n_743 ,in2[5]);
  not csa_tree_add_7_27_groupi_g6464(csa_tree_add_7_27_groupi_n_742 ,in2[1]);
  not csa_tree_add_7_27_groupi_g6465(csa_tree_add_7_27_groupi_n_741 ,in2[4]);
  not csa_tree_add_7_27_groupi_g6466(csa_tree_add_7_27_groupi_n_740 ,in2[9]);
  not csa_tree_add_7_27_groupi_g6467(csa_tree_add_7_27_groupi_n_739 ,in2[3]);
  not csa_tree_add_7_27_groupi_g6468(csa_tree_add_7_27_groupi_n_738 ,in1[15]);
  not csa_tree_add_7_27_groupi_g6469(csa_tree_add_7_27_groupi_n_737 ,in1[1]);
  not csa_tree_add_7_27_groupi_g6470(csa_tree_add_7_27_groupi_n_736 ,in1[10]);
  not csa_tree_add_7_27_groupi_g6471(csa_tree_add_7_27_groupi_n_735 ,in1[5]);
  not csa_tree_add_7_27_groupi_g6472(csa_tree_add_7_27_groupi_n_734 ,in1[6]);
  not csa_tree_add_7_27_groupi_g6473(csa_tree_add_7_27_groupi_n_733 ,in1[2]);
  not csa_tree_add_7_27_groupi_g6474(csa_tree_add_7_27_groupi_n_732 ,in1[9]);
  not csa_tree_add_7_27_groupi_g6475(csa_tree_add_7_27_groupi_n_731 ,in1[14]);
  not csa_tree_add_7_27_groupi_g6476(csa_tree_add_7_27_groupi_n_730 ,in2[14]);
  not csa_tree_add_7_27_groupi_drc_bufs6724(csa_tree_add_7_27_groupi_n_721 ,csa_tree_add_7_27_groupi_n_720);
  not csa_tree_add_7_27_groupi_drc_bufs6726(csa_tree_add_7_27_groupi_n_720 ,csa_tree_add_7_27_groupi_n_1154);
  not csa_tree_add_7_27_groupi_drc_bufs6832(csa_tree_add_7_27_groupi_n_719 ,csa_tree_add_7_27_groupi_n_717);
  not csa_tree_add_7_27_groupi_drc_bufs6833(csa_tree_add_7_27_groupi_n_718 ,csa_tree_add_7_27_groupi_n_717);
  not csa_tree_add_7_27_groupi_drc_bufs6834(csa_tree_add_7_27_groupi_n_717 ,csa_tree_add_7_27_groupi_n_812);
  not csa_tree_add_7_27_groupi_drc_bufs6836(csa_tree_add_7_27_groupi_n_716 ,csa_tree_add_7_27_groupi_n_714);
  not csa_tree_add_7_27_groupi_drc_bufs6837(csa_tree_add_7_27_groupi_n_715 ,csa_tree_add_7_27_groupi_n_714);
  not csa_tree_add_7_27_groupi_drc_bufs6838(csa_tree_add_7_27_groupi_n_714 ,csa_tree_add_7_27_groupi_n_811);
  not csa_tree_add_7_27_groupi_drc_bufs6840(csa_tree_add_7_27_groupi_n_713 ,csa_tree_add_7_27_groupi_n_711);
  not csa_tree_add_7_27_groupi_drc_bufs6841(csa_tree_add_7_27_groupi_n_712 ,csa_tree_add_7_27_groupi_n_711);
  not csa_tree_add_7_27_groupi_drc_bufs6842(csa_tree_add_7_27_groupi_n_711 ,csa_tree_add_7_27_groupi_n_1059);
  not csa_tree_add_7_27_groupi_drc_bufs6844(csa_tree_add_7_27_groupi_n_710 ,csa_tree_add_7_27_groupi_n_708);
  not csa_tree_add_7_27_groupi_drc_bufs6845(csa_tree_add_7_27_groupi_n_709 ,csa_tree_add_7_27_groupi_n_708);
  not csa_tree_add_7_27_groupi_drc_bufs6846(csa_tree_add_7_27_groupi_n_708 ,csa_tree_add_7_27_groupi_n_1072);
  not csa_tree_add_7_27_groupi_drc_bufs6848(csa_tree_add_7_27_groupi_n_707 ,csa_tree_add_7_27_groupi_n_705);
  not csa_tree_add_7_27_groupi_drc_bufs6849(csa_tree_add_7_27_groupi_n_706 ,csa_tree_add_7_27_groupi_n_705);
  not csa_tree_add_7_27_groupi_drc_bufs6850(csa_tree_add_7_27_groupi_n_705 ,csa_tree_add_7_27_groupi_n_726);
  not csa_tree_add_7_27_groupi_drc_bufs6852(csa_tree_add_7_27_groupi_n_704 ,csa_tree_add_7_27_groupi_n_702);
  not csa_tree_add_7_27_groupi_drc_bufs6853(csa_tree_add_7_27_groupi_n_703 ,csa_tree_add_7_27_groupi_n_702);
  not csa_tree_add_7_27_groupi_drc_bufs6854(csa_tree_add_7_27_groupi_n_702 ,csa_tree_add_7_27_groupi_n_1071);
  not csa_tree_add_7_27_groupi_drc_bufs6856(csa_tree_add_7_27_groupi_n_701 ,csa_tree_add_7_27_groupi_n_699);
  not csa_tree_add_7_27_groupi_drc_bufs6857(csa_tree_add_7_27_groupi_n_700 ,csa_tree_add_7_27_groupi_n_699);
  not csa_tree_add_7_27_groupi_drc_bufs6858(csa_tree_add_7_27_groupi_n_699 ,csa_tree_add_7_27_groupi_n_1068);
  not csa_tree_add_7_27_groupi_drc_bufs6860(csa_tree_add_7_27_groupi_n_698 ,csa_tree_add_7_27_groupi_n_696);
  not csa_tree_add_7_27_groupi_drc_bufs6861(csa_tree_add_7_27_groupi_n_697 ,csa_tree_add_7_27_groupi_n_696);
  not csa_tree_add_7_27_groupi_drc_bufs6862(csa_tree_add_7_27_groupi_n_696 ,csa_tree_add_7_27_groupi_n_725);
  not csa_tree_add_7_27_groupi_drc_bufs6864(csa_tree_add_7_27_groupi_n_695 ,csa_tree_add_7_27_groupi_n_693);
  not csa_tree_add_7_27_groupi_drc_bufs6865(csa_tree_add_7_27_groupi_n_694 ,csa_tree_add_7_27_groupi_n_693);
  not csa_tree_add_7_27_groupi_drc_bufs6866(csa_tree_add_7_27_groupi_n_693 ,csa_tree_add_7_27_groupi_n_1067);
  not csa_tree_add_7_27_groupi_drc_bufs6868(csa_tree_add_7_27_groupi_n_692 ,csa_tree_add_7_27_groupi_n_690);
  not csa_tree_add_7_27_groupi_drc_bufs6869(csa_tree_add_7_27_groupi_n_691 ,csa_tree_add_7_27_groupi_n_690);
  not csa_tree_add_7_27_groupi_drc_bufs6870(csa_tree_add_7_27_groupi_n_690 ,csa_tree_add_7_27_groupi_n_1064);
  not csa_tree_add_7_27_groupi_drc_bufs6872(csa_tree_add_7_27_groupi_n_689 ,csa_tree_add_7_27_groupi_n_687);
  not csa_tree_add_7_27_groupi_drc_bufs6873(csa_tree_add_7_27_groupi_n_688 ,csa_tree_add_7_27_groupi_n_687);
  not csa_tree_add_7_27_groupi_drc_bufs6874(csa_tree_add_7_27_groupi_n_687 ,csa_tree_add_7_27_groupi_n_724);
  not csa_tree_add_7_27_groupi_drc_bufs6876(csa_tree_add_7_27_groupi_n_686 ,csa_tree_add_7_27_groupi_n_684);
  not csa_tree_add_7_27_groupi_drc_bufs6877(csa_tree_add_7_27_groupi_n_685 ,csa_tree_add_7_27_groupi_n_684);
  not csa_tree_add_7_27_groupi_drc_bufs6878(csa_tree_add_7_27_groupi_n_684 ,csa_tree_add_7_27_groupi_n_1063);
  not csa_tree_add_7_27_groupi_drc_bufs6880(csa_tree_add_7_27_groupi_n_683 ,csa_tree_add_7_27_groupi_n_681);
  not csa_tree_add_7_27_groupi_drc_bufs6881(csa_tree_add_7_27_groupi_n_682 ,csa_tree_add_7_27_groupi_n_681);
  not csa_tree_add_7_27_groupi_drc_bufs6882(csa_tree_add_7_27_groupi_n_681 ,csa_tree_add_7_27_groupi_n_1060);
  not csa_tree_add_7_27_groupi_drc_bufs6884(csa_tree_add_7_27_groupi_n_680 ,csa_tree_add_7_27_groupi_n_678);
  not csa_tree_add_7_27_groupi_drc_bufs6885(csa_tree_add_7_27_groupi_n_679 ,csa_tree_add_7_27_groupi_n_678);
  not csa_tree_add_7_27_groupi_drc_bufs6886(csa_tree_add_7_27_groupi_n_678 ,csa_tree_add_7_27_groupi_n_723);
  not csa_tree_add_7_27_groupi_drc_bufs6888(csa_tree_add_7_27_groupi_n_677 ,csa_tree_add_7_27_groupi_n_675);
  not csa_tree_add_7_27_groupi_drc_bufs6889(csa_tree_add_7_27_groupi_n_676 ,csa_tree_add_7_27_groupi_n_675);
  not csa_tree_add_7_27_groupi_drc_bufs6890(csa_tree_add_7_27_groupi_n_675 ,csa_tree_add_7_27_groupi_n_722);
  not csa_tree_add_7_27_groupi_drc_bufs6892(csa_tree_add_7_27_groupi_n_674 ,csa_tree_add_7_27_groupi_n_672);
  not csa_tree_add_7_27_groupi_drc_bufs6893(csa_tree_add_7_27_groupi_n_673 ,csa_tree_add_7_27_groupi_n_672);
  not csa_tree_add_7_27_groupi_drc_bufs6894(csa_tree_add_7_27_groupi_n_672 ,csa_tree_add_7_27_groupi_n_811);
  not csa_tree_add_7_27_groupi_drc_bufs6897(csa_tree_add_7_27_groupi_n_671 ,csa_tree_add_7_27_groupi_n_670);
  not csa_tree_add_7_27_groupi_drc_bufs6898(csa_tree_add_7_27_groupi_n_670 ,csa_tree_add_7_27_groupi_n_1164);
  not csa_tree_add_7_27_groupi_drc_bufs6901(csa_tree_add_7_27_groupi_n_669 ,csa_tree_add_7_27_groupi_n_668);
  not csa_tree_add_7_27_groupi_drc_bufs6902(csa_tree_add_7_27_groupi_n_668 ,csa_tree_add_7_27_groupi_n_1161);
  not csa_tree_add_7_27_groupi_drc_bufs6909(csa_tree_add_7_27_groupi_n_667 ,csa_tree_add_7_27_groupi_n_666);
  not csa_tree_add_7_27_groupi_drc_bufs6911(csa_tree_add_7_27_groupi_n_666 ,csa_tree_add_7_27_groupi_n_1074);
  not csa_tree_add_7_27_groupi_drc_bufs6913(csa_tree_add_7_27_groupi_n_665 ,csa_tree_add_7_27_groupi_n_664);
  not csa_tree_add_7_27_groupi_drc_bufs6915(csa_tree_add_7_27_groupi_n_664 ,csa_tree_add_7_27_groupi_n_1070);
  not csa_tree_add_7_27_groupi_drc_bufs6917(csa_tree_add_7_27_groupi_n_663 ,csa_tree_add_7_27_groupi_n_662);
  not csa_tree_add_7_27_groupi_drc_bufs6919(csa_tree_add_7_27_groupi_n_662 ,csa_tree_add_7_27_groupi_n_1066);
  not csa_tree_add_7_27_groupi_drc_bufs6921(csa_tree_add_7_27_groupi_n_661 ,csa_tree_add_7_27_groupi_n_660);
  not csa_tree_add_7_27_groupi_drc_bufs6923(csa_tree_add_7_27_groupi_n_660 ,csa_tree_add_7_27_groupi_n_1062);
  not csa_tree_add_7_27_groupi_drc_bufs7097(csa_tree_add_7_27_groupi_n_659 ,csa_tree_add_7_27_groupi_n_658);
  not csa_tree_add_7_27_groupi_drc_bufs7098(csa_tree_add_7_27_groupi_n_658 ,csa_tree_add_7_27_groupi_n_1163);
  not csa_tree_add_7_27_groupi_drc_bufs7101(csa_tree_add_7_27_groupi_n_657 ,csa_tree_add_7_27_groupi_n_656);
  not csa_tree_add_7_27_groupi_drc_bufs7102(csa_tree_add_7_27_groupi_n_656 ,csa_tree_add_7_27_groupi_n_1160);
  buf csa_tree_add_7_27_groupi_drc_bufs7257(n_8 ,csa_tree_add_7_27_groupi_n_1783);
  buf csa_tree_add_7_27_groupi_drc_bufs7258(n_17 ,csa_tree_add_7_27_groupi_n_2308);
  buf csa_tree_add_7_27_groupi_drc_bufs7259(n_24 ,csa_tree_add_7_27_groupi_n_2329);
  buf csa_tree_add_7_27_groupi_drc_bufs7260(n_25 ,csa_tree_add_7_27_groupi_n_2332);
  buf csa_tree_add_7_27_groupi_drc_bufs7261(n_2 ,csa_tree_add_7_27_groupi_n_1511);
  buf csa_tree_add_7_27_groupi_drc_bufs7262(n_3 ,csa_tree_add_7_27_groupi_n_1536);
  not csa_tree_add_7_27_groupi_drc_bufs7293(csa_tree_add_7_27_groupi_n_649 ,csa_tree_add_7_27_groupi_n_647);
  not csa_tree_add_7_27_groupi_drc_bufs7294(csa_tree_add_7_27_groupi_n_648 ,csa_tree_add_7_27_groupi_n_647);
  not csa_tree_add_7_27_groupi_drc_bufs7295(csa_tree_add_7_27_groupi_n_647 ,csa_tree_add_7_27_groupi_n_937);
  not csa_tree_add_7_27_groupi_drc_bufs7298(csa_tree_add_7_27_groupi_n_646 ,csa_tree_add_7_27_groupi_n_644);
  not csa_tree_add_7_27_groupi_drc_bufs7299(csa_tree_add_7_27_groupi_n_645 ,csa_tree_add_7_27_groupi_n_644);
  not csa_tree_add_7_27_groupi_drc_bufs7300(csa_tree_add_7_27_groupi_n_644 ,csa_tree_add_7_27_groupi_n_936);
  not csa_tree_add_7_27_groupi_drc_bufs7303(csa_tree_add_7_27_groupi_n_643 ,csa_tree_add_7_27_groupi_n_641);
  not csa_tree_add_7_27_groupi_drc_bufs7304(csa_tree_add_7_27_groupi_n_642 ,csa_tree_add_7_27_groupi_n_641);
  not csa_tree_add_7_27_groupi_drc_bufs7305(csa_tree_add_7_27_groupi_n_641 ,csa_tree_add_7_27_groupi_n_939);
  not csa_tree_add_7_27_groupi_drc_bufs7308(csa_tree_add_7_27_groupi_n_640 ,csa_tree_add_7_27_groupi_n_638);
  not csa_tree_add_7_27_groupi_drc_bufs7309(csa_tree_add_7_27_groupi_n_639 ,csa_tree_add_7_27_groupi_n_638);
  not csa_tree_add_7_27_groupi_drc_bufs7310(csa_tree_add_7_27_groupi_n_638 ,csa_tree_add_7_27_groupi_n_963);
  not csa_tree_add_7_27_groupi_drc_bufs7313(csa_tree_add_7_27_groupi_n_637 ,csa_tree_add_7_27_groupi_n_635);
  not csa_tree_add_7_27_groupi_drc_bufs7314(csa_tree_add_7_27_groupi_n_636 ,csa_tree_add_7_27_groupi_n_635);
  not csa_tree_add_7_27_groupi_drc_bufs7315(csa_tree_add_7_27_groupi_n_635 ,csa_tree_add_7_27_groupi_n_938);
  not csa_tree_add_7_27_groupi_drc_bufs7323(csa_tree_add_7_27_groupi_n_634 ,csa_tree_add_7_27_groupi_n_632);
  not csa_tree_add_7_27_groupi_drc_bufs7324(csa_tree_add_7_27_groupi_n_633 ,csa_tree_add_7_27_groupi_n_632);
  not csa_tree_add_7_27_groupi_drc_bufs7325(csa_tree_add_7_27_groupi_n_632 ,csa_tree_add_7_27_groupi_n_752);
  not csa_tree_add_7_27_groupi_drc_bufs7333(csa_tree_add_7_27_groupi_n_631 ,csa_tree_add_7_27_groupi_n_629);
  not csa_tree_add_7_27_groupi_drc_bufs7334(csa_tree_add_7_27_groupi_n_630 ,csa_tree_add_7_27_groupi_n_629);
  not csa_tree_add_7_27_groupi_drc_bufs7335(csa_tree_add_7_27_groupi_n_629 ,csa_tree_add_7_27_groupi_n_747);
  not csa_tree_add_7_27_groupi_drc_bufs7343(csa_tree_add_7_27_groupi_n_628 ,csa_tree_add_7_27_groupi_n_626);
  not csa_tree_add_7_27_groupi_drc_bufs7344(csa_tree_add_7_27_groupi_n_627 ,csa_tree_add_7_27_groupi_n_626);
  not csa_tree_add_7_27_groupi_drc_bufs7345(csa_tree_add_7_27_groupi_n_626 ,csa_tree_add_7_27_groupi_n_737);
  not csa_tree_add_7_27_groupi_drc_bufs7353(csa_tree_add_7_27_groupi_n_625 ,csa_tree_add_7_27_groupi_n_623);
  not csa_tree_add_7_27_groupi_drc_bufs7354(csa_tree_add_7_27_groupi_n_624 ,csa_tree_add_7_27_groupi_n_623);
  not csa_tree_add_7_27_groupi_drc_bufs7355(csa_tree_add_7_27_groupi_n_623 ,csa_tree_add_7_27_groupi_n_736);
  not csa_tree_add_7_27_groupi_drc_bufs7363(csa_tree_add_7_27_groupi_n_622 ,csa_tree_add_7_27_groupi_n_620);
  not csa_tree_add_7_27_groupi_drc_bufs7364(csa_tree_add_7_27_groupi_n_621 ,csa_tree_add_7_27_groupi_n_620);
  not csa_tree_add_7_27_groupi_drc_bufs7365(csa_tree_add_7_27_groupi_n_620 ,csa_tree_add_7_27_groupi_n_735);
  not csa_tree_add_7_27_groupi_drc_bufs7373(csa_tree_add_7_27_groupi_n_619 ,csa_tree_add_7_27_groupi_n_617);
  not csa_tree_add_7_27_groupi_drc_bufs7374(csa_tree_add_7_27_groupi_n_618 ,csa_tree_add_7_27_groupi_n_617);
  not csa_tree_add_7_27_groupi_drc_bufs7375(csa_tree_add_7_27_groupi_n_617 ,csa_tree_add_7_27_groupi_n_734);
  not csa_tree_add_7_27_groupi_drc_bufs7383(csa_tree_add_7_27_groupi_n_616 ,csa_tree_add_7_27_groupi_n_614);
  not csa_tree_add_7_27_groupi_drc_bufs7384(csa_tree_add_7_27_groupi_n_615 ,csa_tree_add_7_27_groupi_n_614);
  not csa_tree_add_7_27_groupi_drc_bufs7385(csa_tree_add_7_27_groupi_n_614 ,csa_tree_add_7_27_groupi_n_732);
  not csa_tree_add_7_27_groupi_drc_bufs7393(csa_tree_add_7_27_groupi_n_613 ,csa_tree_add_7_27_groupi_n_611);
  not csa_tree_add_7_27_groupi_drc_bufs7394(csa_tree_add_7_27_groupi_n_612 ,csa_tree_add_7_27_groupi_n_611);
  not csa_tree_add_7_27_groupi_drc_bufs7395(csa_tree_add_7_27_groupi_n_611 ,csa_tree_add_7_27_groupi_n_731);
  not csa_tree_add_7_27_groupi_drc_bufs7403(csa_tree_add_7_27_groupi_n_610 ,csa_tree_add_7_27_groupi_n_608);
  not csa_tree_add_7_27_groupi_drc_bufs7404(csa_tree_add_7_27_groupi_n_609 ,csa_tree_add_7_27_groupi_n_608);
  not csa_tree_add_7_27_groupi_drc_bufs7405(csa_tree_add_7_27_groupi_n_608 ,csa_tree_add_7_27_groupi_n_753);
  not csa_tree_add_7_27_groupi_drc_bufs7423(csa_tree_add_7_27_groupi_n_607 ,csa_tree_add_7_27_groupi_n_605);
  not csa_tree_add_7_27_groupi_drc_bufs7424(csa_tree_add_7_27_groupi_n_606 ,csa_tree_add_7_27_groupi_n_605);
  not csa_tree_add_7_27_groupi_drc_bufs7425(csa_tree_add_7_27_groupi_n_605 ,csa_tree_add_7_27_groupi_n_751);
  not csa_tree_add_7_27_groupi_drc_bufs7433(csa_tree_add_7_27_groupi_n_604 ,csa_tree_add_7_27_groupi_n_602);
  not csa_tree_add_7_27_groupi_drc_bufs7434(csa_tree_add_7_27_groupi_n_603 ,csa_tree_add_7_27_groupi_n_602);
  not csa_tree_add_7_27_groupi_drc_bufs7435(csa_tree_add_7_27_groupi_n_602 ,csa_tree_add_7_27_groupi_n_750);
  not csa_tree_add_7_27_groupi_drc_bufs7438(csa_tree_add_7_27_groupi_n_601 ,csa_tree_add_7_27_groupi_n_599);
  not csa_tree_add_7_27_groupi_drc_bufs7439(csa_tree_add_7_27_groupi_n_600 ,csa_tree_add_7_27_groupi_n_599);
  not csa_tree_add_7_27_groupi_drc_bufs7440(csa_tree_add_7_27_groupi_n_599 ,csa_tree_add_7_27_groupi_n_748);
  not csa_tree_add_7_27_groupi_drc_bufs7448(csa_tree_add_7_27_groupi_n_598 ,csa_tree_add_7_27_groupi_n_596);
  not csa_tree_add_7_27_groupi_drc_bufs7449(csa_tree_add_7_27_groupi_n_597 ,csa_tree_add_7_27_groupi_n_596);
  not csa_tree_add_7_27_groupi_drc_bufs7450(csa_tree_add_7_27_groupi_n_596 ,csa_tree_add_7_27_groupi_n_749);
  not csa_tree_add_7_27_groupi_drc_bufs7453(csa_tree_add_7_27_groupi_n_595 ,csa_tree_add_7_27_groupi_n_593);
  not csa_tree_add_7_27_groupi_drc_bufs7454(csa_tree_add_7_27_groupi_n_594 ,csa_tree_add_7_27_groupi_n_593);
  not csa_tree_add_7_27_groupi_drc_bufs7455(csa_tree_add_7_27_groupi_n_593 ,csa_tree_add_7_27_groupi_n_733);
  not csa_tree_add_7_27_groupi_drc_bufs7458(csa_tree_add_7_27_groupi_n_592 ,csa_tree_add_7_27_groupi_n_590);
  not csa_tree_add_7_27_groupi_drc_bufs7459(csa_tree_add_7_27_groupi_n_591 ,csa_tree_add_7_27_groupi_n_590);
  not csa_tree_add_7_27_groupi_drc_bufs7460(csa_tree_add_7_27_groupi_n_590 ,csa_tree_add_7_27_groupi_n_738);
  not csa_tree_add_7_27_groupi_drc_bufs7498(csa_tree_add_7_27_groupi_n_589 ,csa_tree_add_7_27_groupi_n_588);
  not csa_tree_add_7_27_groupi_drc_bufs7500(csa_tree_add_7_27_groupi_n_588 ,csa_tree_add_7_27_groupi_n_907);
  not csa_tree_add_7_27_groupi_drc_bufs7503(csa_tree_add_7_27_groupi_n_587 ,csa_tree_add_7_27_groupi_n_586);
  not csa_tree_add_7_27_groupi_drc_bufs7505(csa_tree_add_7_27_groupi_n_586 ,csa_tree_add_7_27_groupi_n_813);
  not csa_tree_add_7_27_groupi_drc_bufs7528(csa_tree_add_7_27_groupi_n_585 ,csa_tree_add_7_27_groupi_n_584);
  not csa_tree_add_7_27_groupi_drc_bufs7530(csa_tree_add_7_27_groupi_n_584 ,csa_tree_add_7_27_groupi_n_967);
  not csa_tree_add_7_27_groupi_drc_bufs7533(csa_tree_add_7_27_groupi_n_583 ,csa_tree_add_7_27_groupi_n_582);
  not csa_tree_add_7_27_groupi_drc_bufs7535(csa_tree_add_7_27_groupi_n_582 ,csa_tree_add_7_27_groupi_n_965);
  not csa_tree_add_7_27_groupi_drc_bufs7538(csa_tree_add_7_27_groupi_n_581 ,csa_tree_add_7_27_groupi_n_580);
  not csa_tree_add_7_27_groupi_drc_bufs7540(csa_tree_add_7_27_groupi_n_580 ,csa_tree_add_7_27_groupi_n_964);
  not csa_tree_add_7_27_groupi_drc_bufs7543(csa_tree_add_7_27_groupi_n_579 ,csa_tree_add_7_27_groupi_n_578);
  not csa_tree_add_7_27_groupi_drc_bufs7545(csa_tree_add_7_27_groupi_n_578 ,csa_tree_add_7_27_groupi_n_968);
  not csa_tree_add_7_27_groupi_drc_bufs7548(csa_tree_add_7_27_groupi_n_577 ,csa_tree_add_7_27_groupi_n_576);
  not csa_tree_add_7_27_groupi_drc_bufs7550(csa_tree_add_7_27_groupi_n_576 ,csa_tree_add_7_27_groupi_n_942);
  not csa_tree_add_7_27_groupi_drc_bufs7553(csa_tree_add_7_27_groupi_n_575 ,csa_tree_add_7_27_groupi_n_574);
  not csa_tree_add_7_27_groupi_drc_bufs7555(csa_tree_add_7_27_groupi_n_574 ,csa_tree_add_7_27_groupi_n_966);
  not csa_tree_add_7_27_groupi_drc_bufs7558(csa_tree_add_7_27_groupi_n_573 ,csa_tree_add_7_27_groupi_n_572);
  not csa_tree_add_7_27_groupi_drc_bufs7560(csa_tree_add_7_27_groupi_n_572 ,csa_tree_add_7_27_groupi_n_940);
  not csa_tree_add_7_27_groupi_drc_bufs7563(csa_tree_add_7_27_groupi_n_571 ,csa_tree_add_7_27_groupi_n_570);
  not csa_tree_add_7_27_groupi_drc_bufs7565(csa_tree_add_7_27_groupi_n_570 ,csa_tree_add_7_27_groupi_n_943);
  not csa_tree_add_7_27_groupi_drc_bufs7568(csa_tree_add_7_27_groupi_n_569 ,csa_tree_add_7_27_groupi_n_568);
  not csa_tree_add_7_27_groupi_drc_bufs7570(csa_tree_add_7_27_groupi_n_568 ,csa_tree_add_7_27_groupi_n_941);
  not csa_tree_add_7_27_groupi_drc_bufs7577(csa_tree_add_7_27_groupi_n_567 ,csa_tree_add_7_27_groupi_n_565);
  not csa_tree_add_7_27_groupi_drc_bufs7578(csa_tree_add_7_27_groupi_n_566 ,csa_tree_add_7_27_groupi_n_565);
  not csa_tree_add_7_27_groupi_drc_bufs7579(csa_tree_add_7_27_groupi_n_565 ,csa_tree_add_7_27_groupi_n_754);
  not csa_tree_add_7_27_groupi_drc_bufs7581(csa_tree_add_7_27_groupi_n_564 ,csa_tree_add_7_27_groupi_n_562);
  not csa_tree_add_7_27_groupi_drc_bufs7582(csa_tree_add_7_27_groupi_n_563 ,csa_tree_add_7_27_groupi_n_562);
  not csa_tree_add_7_27_groupi_drc_bufs7583(csa_tree_add_7_27_groupi_n_562 ,csa_tree_add_7_27_groupi_n_865);
  not csa_tree_add_7_27_groupi_drc_bufs7585(csa_tree_add_7_27_groupi_n_561 ,csa_tree_add_7_27_groupi_n_559);
  not csa_tree_add_7_27_groupi_drc_bufs7586(csa_tree_add_7_27_groupi_n_560 ,csa_tree_add_7_27_groupi_n_559);
  not csa_tree_add_7_27_groupi_drc_bufs7587(csa_tree_add_7_27_groupi_n_559 ,csa_tree_add_7_27_groupi_n_865);
  not csa_tree_add_7_27_groupi_drc_bufs7589(csa_tree_add_7_27_groupi_n_558 ,csa_tree_add_7_27_groupi_n_556);
  not csa_tree_add_7_27_groupi_drc_bufs7590(csa_tree_add_7_27_groupi_n_557 ,csa_tree_add_7_27_groupi_n_556);
  not csa_tree_add_7_27_groupi_drc_bufs7591(csa_tree_add_7_27_groupi_n_556 ,csa_tree_add_7_27_groupi_n_864);
  not csa_tree_add_7_27_groupi_drc_bufs7593(csa_tree_add_7_27_groupi_n_555 ,csa_tree_add_7_27_groupi_n_553);
  not csa_tree_add_7_27_groupi_drc_bufs7594(csa_tree_add_7_27_groupi_n_554 ,csa_tree_add_7_27_groupi_n_553);
  not csa_tree_add_7_27_groupi_drc_bufs7595(csa_tree_add_7_27_groupi_n_553 ,csa_tree_add_7_27_groupi_n_1672);
  not csa_tree_add_7_27_groupi_drc_bufs7597(csa_tree_add_7_27_groupi_n_552 ,csa_tree_add_7_27_groupi_n_550);
  not csa_tree_add_7_27_groupi_drc_bufs7598(csa_tree_add_7_27_groupi_n_551 ,csa_tree_add_7_27_groupi_n_550);
  not csa_tree_add_7_27_groupi_drc_bufs7599(csa_tree_add_7_27_groupi_n_550 ,csa_tree_add_7_27_groupi_n_1566);
  not csa_tree_add_7_27_groupi_drc_bufs7601(csa_tree_add_7_27_groupi_n_549 ,csa_tree_add_7_27_groupi_n_547);
  not csa_tree_add_7_27_groupi_drc_bufs7602(csa_tree_add_7_27_groupi_n_548 ,csa_tree_add_7_27_groupi_n_547);
  not csa_tree_add_7_27_groupi_drc_bufs7603(csa_tree_add_7_27_groupi_n_547 ,csa_tree_add_7_27_groupi_n_1375);
  not csa_tree_add_7_27_groupi_drc_bufs7605(csa_tree_add_7_27_groupi_n_546 ,csa_tree_add_7_27_groupi_n_544);
  not csa_tree_add_7_27_groupi_drc_bufs7606(csa_tree_add_7_27_groupi_n_545 ,csa_tree_add_7_27_groupi_n_544);
  not csa_tree_add_7_27_groupi_drc_bufs7607(csa_tree_add_7_27_groupi_n_544 ,csa_tree_add_7_27_groupi_n_1512);
  not csa_tree_add_7_27_groupi_drc_bufs7609(csa_tree_add_7_27_groupi_n_543 ,csa_tree_add_7_27_groupi_n_542);
  not csa_tree_add_7_27_groupi_drc_bufs7611(csa_tree_add_7_27_groupi_n_542 ,csa_tree_add_7_27_groupi_n_2040);
  not csa_tree_add_7_27_groupi_drc_bufs7613(csa_tree_add_7_27_groupi_n_541 ,csa_tree_add_7_27_groupi_n_539);
  not csa_tree_add_7_27_groupi_drc_bufs7614(csa_tree_add_7_27_groupi_n_540 ,csa_tree_add_7_27_groupi_n_539);
  not csa_tree_add_7_27_groupi_drc_bufs7615(csa_tree_add_7_27_groupi_n_539 ,csa_tree_add_7_27_groupi_n_2040);
  not csa_tree_add_7_27_groupi_drc_bufs7617(csa_tree_add_7_27_groupi_n_538 ,csa_tree_add_7_27_groupi_n_536);
  not csa_tree_add_7_27_groupi_drc_bufs7618(csa_tree_add_7_27_groupi_n_537 ,csa_tree_add_7_27_groupi_n_536);
  not csa_tree_add_7_27_groupi_drc_bufs7619(csa_tree_add_7_27_groupi_n_536 ,csa_tree_add_7_27_groupi_n_1784);
  not csa_tree_add_7_27_groupi_drc_bufs7621(csa_tree_add_7_27_groupi_n_535 ,csa_tree_add_7_27_groupi_n_533);
  not csa_tree_add_7_27_groupi_drc_bufs7622(csa_tree_add_7_27_groupi_n_534 ,csa_tree_add_7_27_groupi_n_533);
  not csa_tree_add_7_27_groupi_drc_bufs7623(csa_tree_add_7_27_groupi_n_533 ,csa_tree_add_7_27_groupi_n_1835);
  not csa_tree_add_7_27_groupi_drc_bufs7625(csa_tree_add_7_27_groupi_n_532 ,csa_tree_add_7_27_groupi_n_530);
  not csa_tree_add_7_27_groupi_drc_bufs7626(csa_tree_add_7_27_groupi_n_531 ,csa_tree_add_7_27_groupi_n_530);
  not csa_tree_add_7_27_groupi_drc_bufs7627(csa_tree_add_7_27_groupi_n_530 ,csa_tree_add_7_27_groupi_n_1878);
  not csa_tree_add_7_27_groupi_drc_bufs7629(csa_tree_add_7_27_groupi_n_529 ,csa_tree_add_7_27_groupi_n_528);
  not csa_tree_add_7_27_groupi_drc_bufs7631(csa_tree_add_7_27_groupi_n_528 ,csa_tree_add_7_27_groupi_n_1620);
  not csa_tree_add_7_27_groupi_drc_bufs7633(csa_tree_add_7_27_groupi_n_527 ,csa_tree_add_7_27_groupi_n_525);
  not csa_tree_add_7_27_groupi_drc_bufs7634(csa_tree_add_7_27_groupi_n_526 ,csa_tree_add_7_27_groupi_n_525);
  not csa_tree_add_7_27_groupi_drc_bufs7635(csa_tree_add_7_27_groupi_n_525 ,csa_tree_add_7_27_groupi_n_1725);
  not csa_tree_add_7_27_groupi_drc_bufs7637(csa_tree_add_7_27_groupi_n_524 ,csa_tree_add_7_27_groupi_n_522);
  not csa_tree_add_7_27_groupi_drc_bufs7638(csa_tree_add_7_27_groupi_n_523 ,csa_tree_add_7_27_groupi_n_522);
  not csa_tree_add_7_27_groupi_drc_bufs7639(csa_tree_add_7_27_groupi_n_522 ,csa_tree_add_7_27_groupi_n_1438);
  not csa_tree_add_7_27_groupi_drc_bufs7641(csa_tree_add_7_27_groupi_n_521 ,csa_tree_add_7_27_groupi_n_519);
  not csa_tree_add_7_27_groupi_drc_bufs7642(csa_tree_add_7_27_groupi_n_520 ,csa_tree_add_7_27_groupi_n_519);
  not csa_tree_add_7_27_groupi_drc_bufs7643(csa_tree_add_7_27_groupi_n_519 ,csa_tree_add_7_27_groupi_n_1994);
  not csa_tree_add_7_27_groupi_drc_bufs7645(csa_tree_add_7_27_groupi_n_518 ,csa_tree_add_7_27_groupi_n_516);
  not csa_tree_add_7_27_groupi_drc_bufs7646(csa_tree_add_7_27_groupi_n_517 ,csa_tree_add_7_27_groupi_n_516);
  not csa_tree_add_7_27_groupi_drc_bufs7647(csa_tree_add_7_27_groupi_n_516 ,csa_tree_add_7_27_groupi_n_1932);
  not csa_tree_add_7_27_groupi_drc_bufs7649(csa_tree_add_7_27_groupi_n_515 ,csa_tree_add_7_27_groupi_n_513);
  not csa_tree_add_7_27_groupi_drc_bufs7650(csa_tree_add_7_27_groupi_n_514 ,csa_tree_add_7_27_groupi_n_513);
  not csa_tree_add_7_27_groupi_drc_bufs7651(csa_tree_add_7_27_groupi_n_513 ,csa_tree_add_7_27_groupi_n_1075);
  not csa_tree_add_7_27_groupi_drc_bufs7653(csa_tree_add_7_27_groupi_n_512 ,csa_tree_add_7_27_groupi_n_510);
  not csa_tree_add_7_27_groupi_drc_bufs7654(csa_tree_add_7_27_groupi_n_511 ,csa_tree_add_7_27_groupi_n_510);
  not csa_tree_add_7_27_groupi_drc_bufs7655(csa_tree_add_7_27_groupi_n_510 ,csa_tree_add_7_27_groupi_n_1236);
  not csa_tree_add_7_27_groupi_drc_bufs7657(csa_tree_add_7_27_groupi_n_509 ,csa_tree_add_7_27_groupi_n_507);
  not csa_tree_add_7_27_groupi_drc_bufs7658(csa_tree_add_7_27_groupi_n_508 ,csa_tree_add_7_27_groupi_n_507);
  not csa_tree_add_7_27_groupi_drc_bufs7659(csa_tree_add_7_27_groupi_n_507 ,csa_tree_add_7_27_groupi_n_2053);
  not csa_tree_add_7_27_groupi_drc_bufs7661(csa_tree_add_7_27_groupi_n_506 ,csa_tree_add_7_27_groupi_n_504);
  not csa_tree_add_7_27_groupi_drc_bufs7662(csa_tree_add_7_27_groupi_n_505 ,csa_tree_add_7_27_groupi_n_504);
  not csa_tree_add_7_27_groupi_drc_bufs7663(csa_tree_add_7_27_groupi_n_504 ,csa_tree_add_7_27_groupi_n_866);
  not csa_tree_add_7_27_groupi_drc_bufs7665(csa_tree_add_7_27_groupi_n_503 ,csa_tree_add_7_27_groupi_n_502);
  not csa_tree_add_7_27_groupi_drc_bufs7667(csa_tree_add_7_27_groupi_n_502 ,csa_tree_add_7_27_groupi_n_1162);
  not csa_tree_add_7_27_groupi_drc_bufs7669(csa_tree_add_7_27_groupi_n_501 ,csa_tree_add_7_27_groupi_n_499);
  not csa_tree_add_7_27_groupi_drc_bufs7670(csa_tree_add_7_27_groupi_n_500 ,csa_tree_add_7_27_groupi_n_499);
  not csa_tree_add_7_27_groupi_drc_bufs7671(csa_tree_add_7_27_groupi_n_499 ,csa_tree_add_7_27_groupi_n_1157);
  not csa_tree_add_7_27_groupi_drc_bufs7673(csa_tree_add_7_27_groupi_n_498 ,csa_tree_add_7_27_groupi_n_497);
  not csa_tree_add_7_27_groupi_drc_bufs7675(csa_tree_add_7_27_groupi_n_497 ,csa_tree_add_7_27_groupi_n_1156);
  not csa_tree_add_7_27_groupi_drc_bufs7677(csa_tree_add_7_27_groupi_n_496 ,csa_tree_add_7_27_groupi_n_495);
  not csa_tree_add_7_27_groupi_drc_bufs7679(csa_tree_add_7_27_groupi_n_495 ,csa_tree_add_7_27_groupi_n_1159);
  not csa_tree_add_7_27_groupi_drc_bufs7681(csa_tree_add_7_27_groupi_n_494 ,csa_tree_add_7_27_groupi_n_725);
  not csa_tree_add_7_27_groupi_drc_bufs7683(csa_tree_add_7_27_groupi_n_725 ,csa_tree_add_7_27_groupi_n_1069);
  not csa_tree_add_7_27_groupi_drc_bufs7685(csa_tree_add_7_27_groupi_n_493 ,csa_tree_add_7_27_groupi_n_723);
  not csa_tree_add_7_27_groupi_drc_bufs7687(csa_tree_add_7_27_groupi_n_723 ,csa_tree_add_7_27_groupi_n_1061);
  not csa_tree_add_7_27_groupi_drc_bufs7689(csa_tree_add_7_27_groupi_n_492 ,csa_tree_add_7_27_groupi_n_724);
  not csa_tree_add_7_27_groupi_drc_bufs7691(csa_tree_add_7_27_groupi_n_724 ,csa_tree_add_7_27_groupi_n_1065);
  not csa_tree_add_7_27_groupi_drc_bufs7693(csa_tree_add_7_27_groupi_n_491 ,csa_tree_add_7_27_groupi_n_726);
  not csa_tree_add_7_27_groupi_drc_bufs7695(csa_tree_add_7_27_groupi_n_726 ,csa_tree_add_7_27_groupi_n_1073);
  not csa_tree_add_7_27_groupi_drc_bufs7697(csa_tree_add_7_27_groupi_n_490 ,csa_tree_add_7_27_groupi_n_722);
  not csa_tree_add_7_27_groupi_drc_bufs7699(csa_tree_add_7_27_groupi_n_722 ,csa_tree_add_7_27_groupi_n_810);
  not csa_tree_add_7_27_groupi_drc_bufs7701(csa_tree_add_7_27_groupi_n_489 ,csa_tree_add_7_27_groupi_n_487);
  not csa_tree_add_7_27_groupi_drc_bufs7702(csa_tree_add_7_27_groupi_n_488 ,csa_tree_add_7_27_groupi_n_487);
  not csa_tree_add_7_27_groupi_drc_bufs7703(csa_tree_add_7_27_groupi_n_487 ,csa_tree_add_7_27_groupi_n_1154);
  not csa_tree_add_7_27_groupi_drc_bufs7706(csa_tree_add_7_27_groupi_n_486 ,csa_tree_add_7_27_groupi_n_728);
  not csa_tree_add_7_27_groupi_drc_bufs7707(csa_tree_add_7_27_groupi_n_728 ,csa_tree_add_7_27_groupi_n_1159);
  not csa_tree_add_7_27_groupi_drc_bufs7710(csa_tree_add_7_27_groupi_n_485 ,csa_tree_add_7_27_groupi_n_727);
  not csa_tree_add_7_27_groupi_drc_bufs7711(csa_tree_add_7_27_groupi_n_727 ,csa_tree_add_7_27_groupi_n_1156);
  not csa_tree_add_7_27_groupi_drc_bufs7714(csa_tree_add_7_27_groupi_n_484 ,csa_tree_add_7_27_groupi_n_729);
  not csa_tree_add_7_27_groupi_drc_bufs7715(csa_tree_add_7_27_groupi_n_729 ,csa_tree_add_7_27_groupi_n_1162);
  not csa_tree_add_7_27_groupi_drc_bufs7717(csa_tree_add_7_27_groupi_n_483 ,csa_tree_add_7_27_groupi_n_481);
  not csa_tree_add_7_27_groupi_drc_bufs7718(csa_tree_add_7_27_groupi_n_482 ,csa_tree_add_7_27_groupi_n_481);
  not csa_tree_add_7_27_groupi_drc_bufs7719(csa_tree_add_7_27_groupi_n_481 ,csa_tree_add_7_27_groupi_n_864);
  not csa_tree_add_7_27_groupi_drc_bufs7721(csa_tree_add_7_27_groupi_n_480 ,csa_tree_add_7_27_groupi_n_478);
  not csa_tree_add_7_27_groupi_drc_bufs7722(csa_tree_add_7_27_groupi_n_479 ,csa_tree_add_7_27_groupi_n_478);
  not csa_tree_add_7_27_groupi_drc_bufs7723(csa_tree_add_7_27_groupi_n_478 ,csa_tree_add_7_27_groupi_n_743);
  not csa_tree_add_7_27_groupi_drc_bufs7725(csa_tree_add_7_27_groupi_n_477 ,csa_tree_add_7_27_groupi_n_475);
  not csa_tree_add_7_27_groupi_drc_bufs7726(csa_tree_add_7_27_groupi_n_476 ,csa_tree_add_7_27_groupi_n_475);
  not csa_tree_add_7_27_groupi_drc_bufs7727(csa_tree_add_7_27_groupi_n_475 ,csa_tree_add_7_27_groupi_n_744);
  not csa_tree_add_7_27_groupi_drc_bufs7729(csa_tree_add_7_27_groupi_n_474 ,csa_tree_add_7_27_groupi_n_472);
  not csa_tree_add_7_27_groupi_drc_bufs7730(csa_tree_add_7_27_groupi_n_473 ,csa_tree_add_7_27_groupi_n_472);
  not csa_tree_add_7_27_groupi_drc_bufs7731(csa_tree_add_7_27_groupi_n_472 ,csa_tree_add_7_27_groupi_n_745);
  not csa_tree_add_7_27_groupi_drc_bufs7733(csa_tree_add_7_27_groupi_n_471 ,csa_tree_add_7_27_groupi_n_469);
  not csa_tree_add_7_27_groupi_drc_bufs7734(csa_tree_add_7_27_groupi_n_470 ,csa_tree_add_7_27_groupi_n_469);
  not csa_tree_add_7_27_groupi_drc_bufs7735(csa_tree_add_7_27_groupi_n_469 ,csa_tree_add_7_27_groupi_n_746);
  not csa_tree_add_7_27_groupi_drc_bufs7737(csa_tree_add_7_27_groupi_n_468 ,csa_tree_add_7_27_groupi_n_466);
  not csa_tree_add_7_27_groupi_drc_bufs7738(csa_tree_add_7_27_groupi_n_467 ,csa_tree_add_7_27_groupi_n_466);
  not csa_tree_add_7_27_groupi_drc_bufs7739(csa_tree_add_7_27_groupi_n_466 ,csa_tree_add_7_27_groupi_n_937);
  not csa_tree_add_7_27_groupi_drc_bufs7741(csa_tree_add_7_27_groupi_n_465 ,csa_tree_add_7_27_groupi_n_463);
  not csa_tree_add_7_27_groupi_drc_bufs7742(csa_tree_add_7_27_groupi_n_464 ,csa_tree_add_7_27_groupi_n_463);
  not csa_tree_add_7_27_groupi_drc_bufs7743(csa_tree_add_7_27_groupi_n_463 ,csa_tree_add_7_27_groupi_n_936);
  not csa_tree_add_7_27_groupi_drc_bufs7745(csa_tree_add_7_27_groupi_n_462 ,csa_tree_add_7_27_groupi_n_460);
  not csa_tree_add_7_27_groupi_drc_bufs7746(csa_tree_add_7_27_groupi_n_461 ,csa_tree_add_7_27_groupi_n_460);
  not csa_tree_add_7_27_groupi_drc_bufs7747(csa_tree_add_7_27_groupi_n_460 ,csa_tree_add_7_27_groupi_n_963);
  not csa_tree_add_7_27_groupi_drc_bufs7749(csa_tree_add_7_27_groupi_n_459 ,csa_tree_add_7_27_groupi_n_457);
  not csa_tree_add_7_27_groupi_drc_bufs7750(csa_tree_add_7_27_groupi_n_458 ,csa_tree_add_7_27_groupi_n_457);
  not csa_tree_add_7_27_groupi_drc_bufs7751(csa_tree_add_7_27_groupi_n_457 ,csa_tree_add_7_27_groupi_n_938);
  not csa_tree_add_7_27_groupi_drc_bufs7753(csa_tree_add_7_27_groupi_n_456 ,csa_tree_add_7_27_groupi_n_454);
  not csa_tree_add_7_27_groupi_drc_bufs7754(csa_tree_add_7_27_groupi_n_455 ,csa_tree_add_7_27_groupi_n_454);
  not csa_tree_add_7_27_groupi_drc_bufs7755(csa_tree_add_7_27_groupi_n_454 ,csa_tree_add_7_27_groupi_n_939);
  not csa_tree_add_7_27_groupi_drc_bufs7758(csa_tree_add_7_27_groupi_n_453 ,csa_tree_add_7_27_groupi_n_452);
  not csa_tree_add_7_27_groupi_drc_bufs7759(csa_tree_add_7_27_groupi_n_452 ,csa_tree_add_7_27_groupi_n_643);
  not csa_tree_add_7_27_groupi_drc_bufs7762(csa_tree_add_7_27_groupi_n_451 ,csa_tree_add_7_27_groupi_n_450);
  not csa_tree_add_7_27_groupi_drc_bufs7763(csa_tree_add_7_27_groupi_n_450 ,csa_tree_add_7_27_groupi_n_628);
  not csa_tree_add_7_27_groupi_drc_bufs7766(csa_tree_add_7_27_groupi_n_449 ,csa_tree_add_7_27_groupi_n_448);
  not csa_tree_add_7_27_groupi_drc_bufs7767(csa_tree_add_7_27_groupi_n_448 ,csa_tree_add_7_27_groupi_n_607);
  not csa_tree_add_7_27_groupi_drc_bufs7769(csa_tree_add_7_27_groupi_n_447 ,csa_tree_add_7_27_groupi_n_445);
  not csa_tree_add_7_27_groupi_drc_bufs7770(csa_tree_add_7_27_groupi_n_446 ,csa_tree_add_7_27_groupi_n_445);
  not csa_tree_add_7_27_groupi_drc_bufs7771(csa_tree_add_7_27_groupi_n_445 ,csa_tree_add_7_27_groupi_n_750);
  not csa_tree_add_7_27_groupi_drc_bufs7773(csa_tree_add_7_27_groupi_n_444 ,csa_tree_add_7_27_groupi_n_442);
  not csa_tree_add_7_27_groupi_drc_bufs7774(csa_tree_add_7_27_groupi_n_443 ,csa_tree_add_7_27_groupi_n_442);
  not csa_tree_add_7_27_groupi_drc_bufs7775(csa_tree_add_7_27_groupi_n_442 ,csa_tree_add_7_27_groupi_n_736);
  not csa_tree_add_7_27_groupi_drc_bufs7778(csa_tree_add_7_27_groupi_n_441 ,csa_tree_add_7_27_groupi_n_440);
  not csa_tree_add_7_27_groupi_drc_bufs7779(csa_tree_add_7_27_groupi_n_440 ,csa_tree_add_7_27_groupi_n_604);
  not csa_tree_add_7_27_groupi_drc_bufs7782(csa_tree_add_7_27_groupi_n_439 ,csa_tree_add_7_27_groupi_n_438);
  not csa_tree_add_7_27_groupi_drc_bufs7783(csa_tree_add_7_27_groupi_n_438 ,csa_tree_add_7_27_groupi_n_601);
  not csa_tree_add_7_27_groupi_drc_bufs7786(csa_tree_add_7_27_groupi_n_437 ,csa_tree_add_7_27_groupi_n_436);
  not csa_tree_add_7_27_groupi_drc_bufs7787(csa_tree_add_7_27_groupi_n_436 ,csa_tree_add_7_27_groupi_n_640);
  not csa_tree_add_7_27_groupi_drc_bufs7790(csa_tree_add_7_27_groupi_n_435 ,csa_tree_add_7_27_groupi_n_434);
  not csa_tree_add_7_27_groupi_drc_bufs7791(csa_tree_add_7_27_groupi_n_434 ,csa_tree_add_7_27_groupi_n_625);
  not csa_tree_add_7_27_groupi_drc_bufs7793(csa_tree_add_7_27_groupi_n_433 ,csa_tree_add_7_27_groupi_n_431);
  not csa_tree_add_7_27_groupi_drc_bufs7794(csa_tree_add_7_27_groupi_n_432 ,csa_tree_add_7_27_groupi_n_431);
  not csa_tree_add_7_27_groupi_drc_bufs7795(csa_tree_add_7_27_groupi_n_431 ,csa_tree_add_7_27_groupi_n_749);
  not csa_tree_add_7_27_groupi_drc_bufs7798(csa_tree_add_7_27_groupi_n_430 ,csa_tree_add_7_27_groupi_n_429);
  not csa_tree_add_7_27_groupi_drc_bufs7799(csa_tree_add_7_27_groupi_n_429 ,csa_tree_add_7_27_groupi_n_598);
  not csa_tree_add_7_27_groupi_drc_bufs7801(csa_tree_add_7_27_groupi_n_428 ,csa_tree_add_7_27_groupi_n_426);
  not csa_tree_add_7_27_groupi_drc_bufs7802(csa_tree_add_7_27_groupi_n_427 ,csa_tree_add_7_27_groupi_n_426);
  not csa_tree_add_7_27_groupi_drc_bufs7803(csa_tree_add_7_27_groupi_n_426 ,csa_tree_add_7_27_groupi_n_735);
  not csa_tree_add_7_27_groupi_drc_bufs7806(csa_tree_add_7_27_groupi_n_425 ,csa_tree_add_7_27_groupi_n_424);
  not csa_tree_add_7_27_groupi_drc_bufs7807(csa_tree_add_7_27_groupi_n_424 ,csa_tree_add_7_27_groupi_n_637);
  not csa_tree_add_7_27_groupi_drc_bufs7810(csa_tree_add_7_27_groupi_n_423 ,csa_tree_add_7_27_groupi_n_422);
  not csa_tree_add_7_27_groupi_drc_bufs7811(csa_tree_add_7_27_groupi_n_422 ,csa_tree_add_7_27_groupi_n_622);
  not csa_tree_add_7_27_groupi_drc_bufs7813(csa_tree_add_7_27_groupi_n_421 ,csa_tree_add_7_27_groupi_n_419);
  not csa_tree_add_7_27_groupi_drc_bufs7814(csa_tree_add_7_27_groupi_n_420 ,csa_tree_add_7_27_groupi_n_419);
  not csa_tree_add_7_27_groupi_drc_bufs7815(csa_tree_add_7_27_groupi_n_419 ,csa_tree_add_7_27_groupi_n_734);
  not csa_tree_add_7_27_groupi_drc_bufs7817(csa_tree_add_7_27_groupi_n_418 ,csa_tree_add_7_27_groupi_n_416);
  not csa_tree_add_7_27_groupi_drc_bufs7818(csa_tree_add_7_27_groupi_n_417 ,csa_tree_add_7_27_groupi_n_416);
  not csa_tree_add_7_27_groupi_drc_bufs7819(csa_tree_add_7_27_groupi_n_416 ,csa_tree_add_7_27_groupi_n_748);
  not csa_tree_add_7_27_groupi_drc_bufs7822(csa_tree_add_7_27_groupi_n_415 ,csa_tree_add_7_27_groupi_n_414);
  not csa_tree_add_7_27_groupi_drc_bufs7823(csa_tree_add_7_27_groupi_n_414 ,csa_tree_add_7_27_groupi_n_619);
  not csa_tree_add_7_27_groupi_drc_bufs7825(csa_tree_add_7_27_groupi_n_413 ,csa_tree_add_7_27_groupi_n_411);
  not csa_tree_add_7_27_groupi_drc_bufs7826(csa_tree_add_7_27_groupi_n_412 ,csa_tree_add_7_27_groupi_n_411);
  not csa_tree_add_7_27_groupi_drc_bufs7827(csa_tree_add_7_27_groupi_n_411 ,csa_tree_add_7_27_groupi_n_752);
  not csa_tree_add_7_27_groupi_drc_bufs7829(csa_tree_add_7_27_groupi_n_410 ,csa_tree_add_7_27_groupi_n_408);
  not csa_tree_add_7_27_groupi_drc_bufs7830(csa_tree_add_7_27_groupi_n_409 ,csa_tree_add_7_27_groupi_n_408);
  not csa_tree_add_7_27_groupi_drc_bufs7831(csa_tree_add_7_27_groupi_n_408 ,csa_tree_add_7_27_groupi_n_732);
  not csa_tree_add_7_27_groupi_drc_bufs7834(csa_tree_add_7_27_groupi_n_407 ,csa_tree_add_7_27_groupi_n_406);
  not csa_tree_add_7_27_groupi_drc_bufs7835(csa_tree_add_7_27_groupi_n_406 ,csa_tree_add_7_27_groupi_n_649);
  not csa_tree_add_7_27_groupi_drc_bufs7838(csa_tree_add_7_27_groupi_n_405 ,csa_tree_add_7_27_groupi_n_404);
  not csa_tree_add_7_27_groupi_drc_bufs7839(csa_tree_add_7_27_groupi_n_404 ,csa_tree_add_7_27_groupi_n_634);
  not csa_tree_add_7_27_groupi_drc_bufs7842(csa_tree_add_7_27_groupi_n_403 ,csa_tree_add_7_27_groupi_n_402);
  not csa_tree_add_7_27_groupi_drc_bufs7843(csa_tree_add_7_27_groupi_n_402 ,csa_tree_add_7_27_groupi_n_616);
  not csa_tree_add_7_27_groupi_drc_bufs7845(csa_tree_add_7_27_groupi_n_401 ,csa_tree_add_7_27_groupi_n_399);
  not csa_tree_add_7_27_groupi_drc_bufs7846(csa_tree_add_7_27_groupi_n_400 ,csa_tree_add_7_27_groupi_n_399);
  not csa_tree_add_7_27_groupi_drc_bufs7847(csa_tree_add_7_27_groupi_n_399 ,csa_tree_add_7_27_groupi_n_731);
  not csa_tree_add_7_27_groupi_drc_bufs7849(csa_tree_add_7_27_groupi_n_398 ,csa_tree_add_7_27_groupi_n_396);
  not csa_tree_add_7_27_groupi_drc_bufs7850(csa_tree_add_7_27_groupi_n_397 ,csa_tree_add_7_27_groupi_n_396);
  not csa_tree_add_7_27_groupi_drc_bufs7851(csa_tree_add_7_27_groupi_n_396 ,csa_tree_add_7_27_groupi_n_747);
  not csa_tree_add_7_27_groupi_drc_bufs7854(csa_tree_add_7_27_groupi_n_395 ,csa_tree_add_7_27_groupi_n_394);
  not csa_tree_add_7_27_groupi_drc_bufs7855(csa_tree_add_7_27_groupi_n_394 ,csa_tree_add_7_27_groupi_n_613);
  not csa_tree_add_7_27_groupi_drc_bufs7857(csa_tree_add_7_27_groupi_n_393 ,csa_tree_add_7_27_groupi_n_391);
  not csa_tree_add_7_27_groupi_drc_bufs7858(csa_tree_add_7_27_groupi_n_392 ,csa_tree_add_7_27_groupi_n_391);
  not csa_tree_add_7_27_groupi_drc_bufs7859(csa_tree_add_7_27_groupi_n_391 ,csa_tree_add_7_27_groupi_n_753);
  not csa_tree_add_7_27_groupi_drc_bufs7861(csa_tree_add_7_27_groupi_n_390 ,csa_tree_add_7_27_groupi_n_388);
  not csa_tree_add_7_27_groupi_drc_bufs7862(csa_tree_add_7_27_groupi_n_389 ,csa_tree_add_7_27_groupi_n_388);
  not csa_tree_add_7_27_groupi_drc_bufs7863(csa_tree_add_7_27_groupi_n_388 ,csa_tree_add_7_27_groupi_n_748);
  not csa_tree_add_7_27_groupi_drc_bufs7866(csa_tree_add_7_27_groupi_n_387 ,csa_tree_add_7_27_groupi_n_386);
  not csa_tree_add_7_27_groupi_drc_bufs7867(csa_tree_add_7_27_groupi_n_386 ,csa_tree_add_7_27_groupi_n_631);
  not csa_tree_add_7_27_groupi_drc_bufs7870(csa_tree_add_7_27_groupi_n_385 ,csa_tree_add_7_27_groupi_n_384);
  not csa_tree_add_7_27_groupi_drc_bufs7871(csa_tree_add_7_27_groupi_n_384 ,csa_tree_add_7_27_groupi_n_610);
  not csa_tree_add_7_27_groupi_drc_bufs7873(csa_tree_add_7_27_groupi_n_383 ,csa_tree_add_7_27_groupi_n_381);
  not csa_tree_add_7_27_groupi_drc_bufs7874(csa_tree_add_7_27_groupi_n_382 ,csa_tree_add_7_27_groupi_n_381);
  not csa_tree_add_7_27_groupi_drc_bufs7875(csa_tree_add_7_27_groupi_n_381 ,csa_tree_add_7_27_groupi_n_733);
  not csa_tree_add_7_27_groupi_drc_bufs7878(csa_tree_add_7_27_groupi_n_380 ,csa_tree_add_7_27_groupi_n_379);
  not csa_tree_add_7_27_groupi_drc_bufs7879(csa_tree_add_7_27_groupi_n_379 ,csa_tree_add_7_27_groupi_n_646);
  not csa_tree_add_7_27_groupi_drc_bufs7881(csa_tree_add_7_27_groupi_n_378 ,csa_tree_add_7_27_groupi_n_376);
  not csa_tree_add_7_27_groupi_drc_bufs7882(csa_tree_add_7_27_groupi_n_377 ,csa_tree_add_7_27_groupi_n_376);
  not csa_tree_add_7_27_groupi_drc_bufs7883(csa_tree_add_7_27_groupi_n_376 ,csa_tree_add_7_27_groupi_n_738);
  not csa_tree_add_7_27_groupi_drc_bufs7885(csa_tree_add_7_27_groupi_n_375 ,csa_tree_add_7_27_groupi_n_373);
  not csa_tree_add_7_27_groupi_drc_bufs7886(csa_tree_add_7_27_groupi_n_374 ,csa_tree_add_7_27_groupi_n_373);
  not csa_tree_add_7_27_groupi_drc_bufs7887(csa_tree_add_7_27_groupi_n_373 ,csa_tree_add_7_27_groupi_n_737);
  not csa_tree_add_7_27_groupi_drc_bufs7889(csa_tree_add_7_27_groupi_n_372 ,csa_tree_add_7_27_groupi_n_370);
  not csa_tree_add_7_27_groupi_drc_bufs7890(csa_tree_add_7_27_groupi_n_371 ,csa_tree_add_7_27_groupi_n_370);
  not csa_tree_add_7_27_groupi_drc_bufs7891(csa_tree_add_7_27_groupi_n_370 ,csa_tree_add_7_27_groupi_n_751);
  not csa_tree_add_7_27_groupi_drc_bufs7893(csa_tree_add_7_27_groupi_n_369 ,csa_tree_add_7_27_groupi_n_368);
  not csa_tree_add_7_27_groupi_drc_bufs7895(csa_tree_add_7_27_groupi_n_368 ,csa_tree_add_7_27_groupi_n_594);
  not csa_tree_add_7_27_groupi_drc_bufs7897(csa_tree_add_7_27_groupi_n_367 ,csa_tree_add_7_27_groupi_n_366);
  not csa_tree_add_7_27_groupi_drc_bufs7899(csa_tree_add_7_27_groupi_n_366 ,csa_tree_add_7_27_groupi_n_591);
  not csa_tree_add_7_27_groupi_drc_bufs7901(csa_tree_add_7_27_groupi_n_365 ,csa_tree_add_7_27_groupi_n_363);
  not csa_tree_add_7_27_groupi_drc_bufs7902(csa_tree_add_7_27_groupi_n_364 ,csa_tree_add_7_27_groupi_n_363);
  not csa_tree_add_7_27_groupi_drc_bufs7903(csa_tree_add_7_27_groupi_n_363 ,csa_tree_add_7_27_groupi_n_751);
  not csa_tree_add_7_27_groupi_drc_bufs7905(csa_tree_add_7_27_groupi_n_362 ,csa_tree_add_7_27_groupi_n_360);
  not csa_tree_add_7_27_groupi_drc_bufs7906(csa_tree_add_7_27_groupi_n_361 ,csa_tree_add_7_27_groupi_n_360);
  not csa_tree_add_7_27_groupi_drc_bufs7907(csa_tree_add_7_27_groupi_n_360 ,csa_tree_add_7_27_groupi_n_737);
  not csa_tree_add_7_27_groupi_drc_bufs7909(csa_tree_add_7_27_groupi_n_359 ,csa_tree_add_7_27_groupi_n_357);
  not csa_tree_add_7_27_groupi_drc_bufs7910(csa_tree_add_7_27_groupi_n_358 ,csa_tree_add_7_27_groupi_n_357);
  not csa_tree_add_7_27_groupi_drc_bufs7911(csa_tree_add_7_27_groupi_n_357 ,csa_tree_add_7_27_groupi_n_606);
  not csa_tree_add_7_27_groupi_drc_bufs7913(csa_tree_add_7_27_groupi_n_356 ,csa_tree_add_7_27_groupi_n_354);
  not csa_tree_add_7_27_groupi_drc_bufs7914(csa_tree_add_7_27_groupi_n_355 ,csa_tree_add_7_27_groupi_n_354);
  not csa_tree_add_7_27_groupi_drc_bufs7915(csa_tree_add_7_27_groupi_n_354 ,csa_tree_add_7_27_groupi_n_645);
  not csa_tree_add_7_27_groupi_drc_bufs7917(csa_tree_add_7_27_groupi_n_353 ,csa_tree_add_7_27_groupi_n_351);
  not csa_tree_add_7_27_groupi_drc_bufs7918(csa_tree_add_7_27_groupi_n_352 ,csa_tree_add_7_27_groupi_n_351);
  not csa_tree_add_7_27_groupi_drc_bufs7919(csa_tree_add_7_27_groupi_n_351 ,csa_tree_add_7_27_groupi_n_750);
  not csa_tree_add_7_27_groupi_drc_bufs7921(csa_tree_add_7_27_groupi_n_350 ,csa_tree_add_7_27_groupi_n_348);
  not csa_tree_add_7_27_groupi_drc_bufs7922(csa_tree_add_7_27_groupi_n_349 ,csa_tree_add_7_27_groupi_n_348);
  not csa_tree_add_7_27_groupi_drc_bufs7923(csa_tree_add_7_27_groupi_n_348 ,csa_tree_add_7_27_groupi_n_627);
  not csa_tree_add_7_27_groupi_drc_bufs7925(csa_tree_add_7_27_groupi_n_347 ,csa_tree_add_7_27_groupi_n_345);
  not csa_tree_add_7_27_groupi_drc_bufs7926(csa_tree_add_7_27_groupi_n_346 ,csa_tree_add_7_27_groupi_n_345);
  not csa_tree_add_7_27_groupi_drc_bufs7927(csa_tree_add_7_27_groupi_n_345 ,csa_tree_add_7_27_groupi_n_603);
  not csa_tree_add_7_27_groupi_drc_bufs7929(csa_tree_add_7_27_groupi_n_344 ,csa_tree_add_7_27_groupi_n_342);
  not csa_tree_add_7_27_groupi_drc_bufs7930(csa_tree_add_7_27_groupi_n_343 ,csa_tree_add_7_27_groupi_n_342);
  not csa_tree_add_7_27_groupi_drc_bufs7931(csa_tree_add_7_27_groupi_n_342 ,csa_tree_add_7_27_groupi_n_939);
  not csa_tree_add_7_27_groupi_drc_bufs7933(csa_tree_add_7_27_groupi_n_341 ,csa_tree_add_7_27_groupi_n_339);
  not csa_tree_add_7_27_groupi_drc_bufs7934(csa_tree_add_7_27_groupi_n_340 ,csa_tree_add_7_27_groupi_n_339);
  not csa_tree_add_7_27_groupi_drc_bufs7935(csa_tree_add_7_27_groupi_n_339 ,csa_tree_add_7_27_groupi_n_600);
  not csa_tree_add_7_27_groupi_drc_bufs7937(csa_tree_add_7_27_groupi_n_338 ,csa_tree_add_7_27_groupi_n_336);
  not csa_tree_add_7_27_groupi_drc_bufs7938(csa_tree_add_7_27_groupi_n_337 ,csa_tree_add_7_27_groupi_n_336);
  not csa_tree_add_7_27_groupi_drc_bufs7939(csa_tree_add_7_27_groupi_n_336 ,csa_tree_add_7_27_groupi_n_592);
  not csa_tree_add_7_27_groupi_drc_bufs7941(csa_tree_add_7_27_groupi_n_335 ,csa_tree_add_7_27_groupi_n_333);
  not csa_tree_add_7_27_groupi_drc_bufs7942(csa_tree_add_7_27_groupi_n_334 ,csa_tree_add_7_27_groupi_n_333);
  not csa_tree_add_7_27_groupi_drc_bufs7943(csa_tree_add_7_27_groupi_n_333 ,csa_tree_add_7_27_groupi_n_736);
  not csa_tree_add_7_27_groupi_drc_bufs7945(csa_tree_add_7_27_groupi_n_332 ,csa_tree_add_7_27_groupi_n_330);
  not csa_tree_add_7_27_groupi_drc_bufs7946(csa_tree_add_7_27_groupi_n_331 ,csa_tree_add_7_27_groupi_n_330);
  not csa_tree_add_7_27_groupi_drc_bufs7947(csa_tree_add_7_27_groupi_n_330 ,csa_tree_add_7_27_groupi_n_749);
  not csa_tree_add_7_27_groupi_drc_bufs7949(csa_tree_add_7_27_groupi_n_329 ,csa_tree_add_7_27_groupi_n_327);
  not csa_tree_add_7_27_groupi_drc_bufs7950(csa_tree_add_7_27_groupi_n_328 ,csa_tree_add_7_27_groupi_n_327);
  not csa_tree_add_7_27_groupi_drc_bufs7951(csa_tree_add_7_27_groupi_n_327 ,csa_tree_add_7_27_groupi_n_642);
  not csa_tree_add_7_27_groupi_drc_bufs7953(csa_tree_add_7_27_groupi_n_326 ,csa_tree_add_7_27_groupi_n_324);
  not csa_tree_add_7_27_groupi_drc_bufs7954(csa_tree_add_7_27_groupi_n_325 ,csa_tree_add_7_27_groupi_n_324);
  not csa_tree_add_7_27_groupi_drc_bufs7955(csa_tree_add_7_27_groupi_n_324 ,csa_tree_add_7_27_groupi_n_624);
  not csa_tree_add_7_27_groupi_drc_bufs7957(csa_tree_add_7_27_groupi_n_323 ,csa_tree_add_7_27_groupi_n_321);
  not csa_tree_add_7_27_groupi_drc_bufs7958(csa_tree_add_7_27_groupi_n_322 ,csa_tree_add_7_27_groupi_n_321);
  not csa_tree_add_7_27_groupi_drc_bufs7959(csa_tree_add_7_27_groupi_n_321 ,csa_tree_add_7_27_groupi_n_597);
  not csa_tree_add_7_27_groupi_drc_bufs7961(csa_tree_add_7_27_groupi_n_320 ,csa_tree_add_7_27_groupi_n_318);
  not csa_tree_add_7_27_groupi_drc_bufs7962(csa_tree_add_7_27_groupi_n_319 ,csa_tree_add_7_27_groupi_n_318);
  not csa_tree_add_7_27_groupi_drc_bufs7963(csa_tree_add_7_27_groupi_n_318 ,csa_tree_add_7_27_groupi_n_595);
  not csa_tree_add_7_27_groupi_drc_bufs7965(csa_tree_add_7_27_groupi_n_317 ,csa_tree_add_7_27_groupi_n_315);
  not csa_tree_add_7_27_groupi_drc_bufs7966(csa_tree_add_7_27_groupi_n_316 ,csa_tree_add_7_27_groupi_n_315);
  not csa_tree_add_7_27_groupi_drc_bufs7967(csa_tree_add_7_27_groupi_n_315 ,csa_tree_add_7_27_groupi_n_937);
  not csa_tree_add_7_27_groupi_drc_bufs7969(csa_tree_add_7_27_groupi_n_314 ,csa_tree_add_7_27_groupi_n_312);
  not csa_tree_add_7_27_groupi_drc_bufs7970(csa_tree_add_7_27_groupi_n_313 ,csa_tree_add_7_27_groupi_n_312);
  not csa_tree_add_7_27_groupi_drc_bufs7971(csa_tree_add_7_27_groupi_n_312 ,csa_tree_add_7_27_groupi_n_735);
  not csa_tree_add_7_27_groupi_drc_bufs7973(csa_tree_add_7_27_groupi_n_311 ,csa_tree_add_7_27_groupi_n_309);
  not csa_tree_add_7_27_groupi_drc_bufs7974(csa_tree_add_7_27_groupi_n_310 ,csa_tree_add_7_27_groupi_n_309);
  not csa_tree_add_7_27_groupi_drc_bufs7975(csa_tree_add_7_27_groupi_n_309 ,csa_tree_add_7_27_groupi_n_639);
  not csa_tree_add_7_27_groupi_drc_bufs7977(csa_tree_add_7_27_groupi_n_308 ,csa_tree_add_7_27_groupi_n_306);
  not csa_tree_add_7_27_groupi_drc_bufs7978(csa_tree_add_7_27_groupi_n_307 ,csa_tree_add_7_27_groupi_n_306);
  not csa_tree_add_7_27_groupi_drc_bufs7979(csa_tree_add_7_27_groupi_n_306 ,csa_tree_add_7_27_groupi_n_621);
  not csa_tree_add_7_27_groupi_drc_bufs7981(csa_tree_add_7_27_groupi_n_305 ,csa_tree_add_7_27_groupi_n_303);
  not csa_tree_add_7_27_groupi_drc_bufs7982(csa_tree_add_7_27_groupi_n_304 ,csa_tree_add_7_27_groupi_n_303);
  not csa_tree_add_7_27_groupi_drc_bufs7983(csa_tree_add_7_27_groupi_n_303 ,csa_tree_add_7_27_groupi_n_963);
  not csa_tree_add_7_27_groupi_drc_bufs7985(csa_tree_add_7_27_groupi_n_302 ,csa_tree_add_7_27_groupi_n_300);
  not csa_tree_add_7_27_groupi_drc_bufs7986(csa_tree_add_7_27_groupi_n_301 ,csa_tree_add_7_27_groupi_n_300);
  not csa_tree_add_7_27_groupi_drc_bufs7987(csa_tree_add_7_27_groupi_n_300 ,csa_tree_add_7_27_groupi_n_734);
  not csa_tree_add_7_27_groupi_drc_bufs7989(csa_tree_add_7_27_groupi_n_299 ,csa_tree_add_7_27_groupi_n_297);
  not csa_tree_add_7_27_groupi_drc_bufs7990(csa_tree_add_7_27_groupi_n_298 ,csa_tree_add_7_27_groupi_n_297);
  not csa_tree_add_7_27_groupi_drc_bufs7991(csa_tree_add_7_27_groupi_n_297 ,csa_tree_add_7_27_groupi_n_636);
  not csa_tree_add_7_27_groupi_drc_bufs7993(csa_tree_add_7_27_groupi_n_296 ,csa_tree_add_7_27_groupi_n_294);
  not csa_tree_add_7_27_groupi_drc_bufs7994(csa_tree_add_7_27_groupi_n_295 ,csa_tree_add_7_27_groupi_n_294);
  not csa_tree_add_7_27_groupi_drc_bufs7995(csa_tree_add_7_27_groupi_n_294 ,csa_tree_add_7_27_groupi_n_618);
  not csa_tree_add_7_27_groupi_drc_bufs7997(csa_tree_add_7_27_groupi_n_293 ,csa_tree_add_7_27_groupi_n_291);
  not csa_tree_add_7_27_groupi_drc_bufs7998(csa_tree_add_7_27_groupi_n_292 ,csa_tree_add_7_27_groupi_n_291);
  not csa_tree_add_7_27_groupi_drc_bufs7999(csa_tree_add_7_27_groupi_n_291 ,csa_tree_add_7_27_groupi_n_732);
  not csa_tree_add_7_27_groupi_drc_bufs8001(csa_tree_add_7_27_groupi_n_290 ,csa_tree_add_7_27_groupi_n_288);
  not csa_tree_add_7_27_groupi_drc_bufs8002(csa_tree_add_7_27_groupi_n_289 ,csa_tree_add_7_27_groupi_n_288);
  not csa_tree_add_7_27_groupi_drc_bufs8003(csa_tree_add_7_27_groupi_n_288 ,csa_tree_add_7_27_groupi_n_752);
  not csa_tree_add_7_27_groupi_drc_bufs8005(csa_tree_add_7_27_groupi_n_287 ,csa_tree_add_7_27_groupi_n_285);
  not csa_tree_add_7_27_groupi_drc_bufs8006(csa_tree_add_7_27_groupi_n_286 ,csa_tree_add_7_27_groupi_n_285);
  not csa_tree_add_7_27_groupi_drc_bufs8007(csa_tree_add_7_27_groupi_n_285 ,csa_tree_add_7_27_groupi_n_615);
  not csa_tree_add_7_27_groupi_drc_bufs8009(csa_tree_add_7_27_groupi_n_284 ,csa_tree_add_7_27_groupi_n_282);
  not csa_tree_add_7_27_groupi_drc_bufs8010(csa_tree_add_7_27_groupi_n_283 ,csa_tree_add_7_27_groupi_n_282);
  not csa_tree_add_7_27_groupi_drc_bufs8011(csa_tree_add_7_27_groupi_n_282 ,csa_tree_add_7_27_groupi_n_938);
  not csa_tree_add_7_27_groupi_drc_bufs8013(csa_tree_add_7_27_groupi_n_281 ,csa_tree_add_7_27_groupi_n_279);
  not csa_tree_add_7_27_groupi_drc_bufs8014(csa_tree_add_7_27_groupi_n_280 ,csa_tree_add_7_27_groupi_n_279);
  not csa_tree_add_7_27_groupi_drc_bufs8015(csa_tree_add_7_27_groupi_n_279 ,csa_tree_add_7_27_groupi_n_731);
  not csa_tree_add_7_27_groupi_drc_bufs8017(csa_tree_add_7_27_groupi_n_278 ,csa_tree_add_7_27_groupi_n_276);
  not csa_tree_add_7_27_groupi_drc_bufs8018(csa_tree_add_7_27_groupi_n_277 ,csa_tree_add_7_27_groupi_n_276);
  not csa_tree_add_7_27_groupi_drc_bufs8019(csa_tree_add_7_27_groupi_n_276 ,csa_tree_add_7_27_groupi_n_648);
  not csa_tree_add_7_27_groupi_drc_bufs8021(csa_tree_add_7_27_groupi_n_275 ,csa_tree_add_7_27_groupi_n_273);
  not csa_tree_add_7_27_groupi_drc_bufs8022(csa_tree_add_7_27_groupi_n_274 ,csa_tree_add_7_27_groupi_n_273);
  not csa_tree_add_7_27_groupi_drc_bufs8023(csa_tree_add_7_27_groupi_n_273 ,csa_tree_add_7_27_groupi_n_633);
  not csa_tree_add_7_27_groupi_drc_bufs8025(csa_tree_add_7_27_groupi_n_272 ,csa_tree_add_7_27_groupi_n_270);
  not csa_tree_add_7_27_groupi_drc_bufs8026(csa_tree_add_7_27_groupi_n_271 ,csa_tree_add_7_27_groupi_n_270);
  not csa_tree_add_7_27_groupi_drc_bufs8027(csa_tree_add_7_27_groupi_n_270 ,csa_tree_add_7_27_groupi_n_612);
  not csa_tree_add_7_27_groupi_drc_bufs8029(csa_tree_add_7_27_groupi_n_269 ,csa_tree_add_7_27_groupi_n_267);
  not csa_tree_add_7_27_groupi_drc_bufs8030(csa_tree_add_7_27_groupi_n_268 ,csa_tree_add_7_27_groupi_n_267);
  not csa_tree_add_7_27_groupi_drc_bufs8031(csa_tree_add_7_27_groupi_n_267 ,csa_tree_add_7_27_groupi_n_936);
  not csa_tree_add_7_27_groupi_drc_bufs8033(csa_tree_add_7_27_groupi_n_266 ,csa_tree_add_7_27_groupi_n_264);
  not csa_tree_add_7_27_groupi_drc_bufs8034(csa_tree_add_7_27_groupi_n_265 ,csa_tree_add_7_27_groupi_n_264);
  not csa_tree_add_7_27_groupi_drc_bufs8035(csa_tree_add_7_27_groupi_n_264 ,csa_tree_add_7_27_groupi_n_753);
  not csa_tree_add_7_27_groupi_drc_bufs8037(csa_tree_add_7_27_groupi_n_263 ,csa_tree_add_7_27_groupi_n_261);
  not csa_tree_add_7_27_groupi_drc_bufs8038(csa_tree_add_7_27_groupi_n_262 ,csa_tree_add_7_27_groupi_n_261);
  not csa_tree_add_7_27_groupi_drc_bufs8039(csa_tree_add_7_27_groupi_n_261 ,csa_tree_add_7_27_groupi_n_747);
  not csa_tree_add_7_27_groupi_drc_bufs8041(csa_tree_add_7_27_groupi_n_260 ,csa_tree_add_7_27_groupi_n_258);
  not csa_tree_add_7_27_groupi_drc_bufs8042(csa_tree_add_7_27_groupi_n_259 ,csa_tree_add_7_27_groupi_n_258);
  not csa_tree_add_7_27_groupi_drc_bufs8043(csa_tree_add_7_27_groupi_n_258 ,csa_tree_add_7_27_groupi_n_609);
  not csa_tree_add_7_27_groupi_drc_bufs8045(csa_tree_add_7_27_groupi_n_257 ,csa_tree_add_7_27_groupi_n_255);
  not csa_tree_add_7_27_groupi_drc_bufs8046(csa_tree_add_7_27_groupi_n_256 ,csa_tree_add_7_27_groupi_n_255);
  not csa_tree_add_7_27_groupi_drc_bufs8047(csa_tree_add_7_27_groupi_n_255 ,csa_tree_add_7_27_groupi_n_733);
  not csa_tree_add_7_27_groupi_drc_bufs8049(csa_tree_add_7_27_groupi_n_254 ,csa_tree_add_7_27_groupi_n_252);
  not csa_tree_add_7_27_groupi_drc_bufs8050(csa_tree_add_7_27_groupi_n_253 ,csa_tree_add_7_27_groupi_n_252);
  not csa_tree_add_7_27_groupi_drc_bufs8051(csa_tree_add_7_27_groupi_n_252 ,csa_tree_add_7_27_groupi_n_630);
  not csa_tree_add_7_27_groupi_drc_bufs8053(csa_tree_add_7_27_groupi_n_251 ,csa_tree_add_7_27_groupi_n_249);
  not csa_tree_add_7_27_groupi_drc_bufs8054(csa_tree_add_7_27_groupi_n_250 ,csa_tree_add_7_27_groupi_n_249);
  not csa_tree_add_7_27_groupi_drc_bufs8055(csa_tree_add_7_27_groupi_n_249 ,csa_tree_add_7_27_groupi_n_738);
  not csa_tree_add_7_27_groupi_drc_bufs8057(csa_tree_add_7_27_groupi_n_248 ,csa_tree_add_7_27_groupi_n_246);
  not csa_tree_add_7_27_groupi_drc_bufs8058(csa_tree_add_7_27_groupi_n_247 ,csa_tree_add_7_27_groupi_n_246);
  not csa_tree_add_7_27_groupi_drc_bufs8059(csa_tree_add_7_27_groupi_n_246 ,csa_tree_add_7_27_groupi_n_968);
  not csa_tree_add_7_27_groupi_drc_bufs8061(csa_tree_add_7_27_groupi_n_245 ,csa_tree_add_7_27_groupi_n_243);
  not csa_tree_add_7_27_groupi_drc_bufs8062(csa_tree_add_7_27_groupi_n_244 ,csa_tree_add_7_27_groupi_n_243);
  not csa_tree_add_7_27_groupi_drc_bufs8063(csa_tree_add_7_27_groupi_n_243 ,csa_tree_add_7_27_groupi_n_967);
  not csa_tree_add_7_27_groupi_drc_bufs8065(csa_tree_add_7_27_groupi_n_242 ,csa_tree_add_7_27_groupi_n_240);
  not csa_tree_add_7_27_groupi_drc_bufs8066(csa_tree_add_7_27_groupi_n_241 ,csa_tree_add_7_27_groupi_n_240);
  not csa_tree_add_7_27_groupi_drc_bufs8067(csa_tree_add_7_27_groupi_n_240 ,csa_tree_add_7_27_groupi_n_965);
  not csa_tree_add_7_27_groupi_drc_bufs8069(csa_tree_add_7_27_groupi_n_239 ,csa_tree_add_7_27_groupi_n_237);
  not csa_tree_add_7_27_groupi_drc_bufs8070(csa_tree_add_7_27_groupi_n_238 ,csa_tree_add_7_27_groupi_n_237);
  not csa_tree_add_7_27_groupi_drc_bufs8071(csa_tree_add_7_27_groupi_n_237 ,csa_tree_add_7_27_groupi_n_964);
  not csa_tree_add_7_27_groupi_drc_bufs8073(csa_tree_add_7_27_groupi_n_236 ,csa_tree_add_7_27_groupi_n_234);
  not csa_tree_add_7_27_groupi_drc_bufs8074(csa_tree_add_7_27_groupi_n_235 ,csa_tree_add_7_27_groupi_n_234);
  not csa_tree_add_7_27_groupi_drc_bufs8075(csa_tree_add_7_27_groupi_n_234 ,csa_tree_add_7_27_groupi_n_907);
  not csa_tree_add_7_27_groupi_drc_bufs8077(csa_tree_add_7_27_groupi_n_233 ,csa_tree_add_7_27_groupi_n_231);
  not csa_tree_add_7_27_groupi_drc_bufs8078(csa_tree_add_7_27_groupi_n_232 ,csa_tree_add_7_27_groupi_n_231);
  not csa_tree_add_7_27_groupi_drc_bufs8079(csa_tree_add_7_27_groupi_n_231 ,csa_tree_add_7_27_groupi_n_813);
  not csa_tree_add_7_27_groupi_drc_bufs8081(csa_tree_add_7_27_groupi_n_230 ,csa_tree_add_7_27_groupi_n_228);
  not csa_tree_add_7_27_groupi_drc_bufs8082(csa_tree_add_7_27_groupi_n_229 ,csa_tree_add_7_27_groupi_n_228);
  not csa_tree_add_7_27_groupi_drc_bufs8083(csa_tree_add_7_27_groupi_n_228 ,csa_tree_add_7_27_groupi_n_571);
  not csa_tree_add_7_27_groupi_drc_bufs8085(csa_tree_add_7_27_groupi_n_227 ,csa_tree_add_7_27_groupi_n_225);
  not csa_tree_add_7_27_groupi_drc_bufs8086(csa_tree_add_7_27_groupi_n_226 ,csa_tree_add_7_27_groupi_n_225);
  not csa_tree_add_7_27_groupi_drc_bufs8087(csa_tree_add_7_27_groupi_n_225 ,csa_tree_add_7_27_groupi_n_968);
  not csa_tree_add_7_27_groupi_drc_bufs8089(csa_tree_add_7_27_groupi_n_224 ,csa_tree_add_7_27_groupi_n_222);
  not csa_tree_add_7_27_groupi_drc_bufs8090(csa_tree_add_7_27_groupi_n_223 ,csa_tree_add_7_27_groupi_n_222);
  not csa_tree_add_7_27_groupi_drc_bufs8091(csa_tree_add_7_27_groupi_n_222 ,csa_tree_add_7_27_groupi_n_581);
  not csa_tree_add_7_27_groupi_drc_bufs8093(csa_tree_add_7_27_groupi_n_221 ,csa_tree_add_7_27_groupi_n_219);
  not csa_tree_add_7_27_groupi_drc_bufs8094(csa_tree_add_7_27_groupi_n_220 ,csa_tree_add_7_27_groupi_n_219);
  not csa_tree_add_7_27_groupi_drc_bufs8095(csa_tree_add_7_27_groupi_n_219 ,csa_tree_add_7_27_groupi_n_941);
  not csa_tree_add_7_27_groupi_drc_bufs8097(csa_tree_add_7_27_groupi_n_218 ,csa_tree_add_7_27_groupi_n_216);
  not csa_tree_add_7_27_groupi_drc_bufs8098(csa_tree_add_7_27_groupi_n_217 ,csa_tree_add_7_27_groupi_n_216);
  not csa_tree_add_7_27_groupi_drc_bufs8099(csa_tree_add_7_27_groupi_n_216 ,csa_tree_add_7_27_groupi_n_585);
  not csa_tree_add_7_27_groupi_drc_bufs8101(csa_tree_add_7_27_groupi_n_215 ,csa_tree_add_7_27_groupi_n_213);
  not csa_tree_add_7_27_groupi_drc_bufs8102(csa_tree_add_7_27_groupi_n_214 ,csa_tree_add_7_27_groupi_n_213);
  not csa_tree_add_7_27_groupi_drc_bufs8103(csa_tree_add_7_27_groupi_n_213 ,csa_tree_add_7_27_groupi_n_577);
  not csa_tree_add_7_27_groupi_drc_bufs8105(csa_tree_add_7_27_groupi_n_212 ,csa_tree_add_7_27_groupi_n_210);
  not csa_tree_add_7_27_groupi_drc_bufs8106(csa_tree_add_7_27_groupi_n_211 ,csa_tree_add_7_27_groupi_n_210);
  not csa_tree_add_7_27_groupi_drc_bufs8107(csa_tree_add_7_27_groupi_n_210 ,csa_tree_add_7_27_groupi_n_581);
  not csa_tree_add_7_27_groupi_drc_bufs8109(csa_tree_add_7_27_groupi_n_209 ,csa_tree_add_7_27_groupi_n_207);
  not csa_tree_add_7_27_groupi_drc_bufs8110(csa_tree_add_7_27_groupi_n_208 ,csa_tree_add_7_27_groupi_n_207);
  not csa_tree_add_7_27_groupi_drc_bufs8111(csa_tree_add_7_27_groupi_n_207 ,csa_tree_add_7_27_groupi_n_575);
  not csa_tree_add_7_27_groupi_drc_bufs8113(csa_tree_add_7_27_groupi_n_206 ,csa_tree_add_7_27_groupi_n_204);
  not csa_tree_add_7_27_groupi_drc_bufs8114(csa_tree_add_7_27_groupi_n_205 ,csa_tree_add_7_27_groupi_n_204);
  not csa_tree_add_7_27_groupi_drc_bufs8115(csa_tree_add_7_27_groupi_n_204 ,csa_tree_add_7_27_groupi_n_965);
  not csa_tree_add_7_27_groupi_drc_bufs8117(csa_tree_add_7_27_groupi_n_203 ,csa_tree_add_7_27_groupi_n_201);
  not csa_tree_add_7_27_groupi_drc_bufs8118(csa_tree_add_7_27_groupi_n_202 ,csa_tree_add_7_27_groupi_n_201);
  not csa_tree_add_7_27_groupi_drc_bufs8119(csa_tree_add_7_27_groupi_n_201 ,csa_tree_add_7_27_groupi_n_579);
  not csa_tree_add_7_27_groupi_drc_bufs8121(csa_tree_add_7_27_groupi_n_200 ,csa_tree_add_7_27_groupi_n_198);
  not csa_tree_add_7_27_groupi_drc_bufs8122(csa_tree_add_7_27_groupi_n_199 ,csa_tree_add_7_27_groupi_n_198);
  not csa_tree_add_7_27_groupi_drc_bufs8123(csa_tree_add_7_27_groupi_n_198 ,csa_tree_add_7_27_groupi_n_579);
  not csa_tree_add_7_27_groupi_drc_bufs8125(csa_tree_add_7_27_groupi_n_197 ,csa_tree_add_7_27_groupi_n_195);
  not csa_tree_add_7_27_groupi_drc_bufs8126(csa_tree_add_7_27_groupi_n_196 ,csa_tree_add_7_27_groupi_n_195);
  not csa_tree_add_7_27_groupi_drc_bufs8127(csa_tree_add_7_27_groupi_n_195 ,csa_tree_add_7_27_groupi_n_573);
  not csa_tree_add_7_27_groupi_drc_bufs8129(csa_tree_add_7_27_groupi_n_194 ,csa_tree_add_7_27_groupi_n_192);
  not csa_tree_add_7_27_groupi_drc_bufs8130(csa_tree_add_7_27_groupi_n_193 ,csa_tree_add_7_27_groupi_n_192);
  not csa_tree_add_7_27_groupi_drc_bufs8131(csa_tree_add_7_27_groupi_n_192 ,csa_tree_add_7_27_groupi_n_940);
  not csa_tree_add_7_27_groupi_drc_bufs8133(csa_tree_add_7_27_groupi_n_191 ,csa_tree_add_7_27_groupi_n_189);
  not csa_tree_add_7_27_groupi_drc_bufs8134(csa_tree_add_7_27_groupi_n_190 ,csa_tree_add_7_27_groupi_n_189);
  not csa_tree_add_7_27_groupi_drc_bufs8135(csa_tree_add_7_27_groupi_n_189 ,csa_tree_add_7_27_groupi_n_967);
  not csa_tree_add_7_27_groupi_drc_bufs8137(csa_tree_add_7_27_groupi_n_188 ,csa_tree_add_7_27_groupi_n_186);
  not csa_tree_add_7_27_groupi_drc_bufs8138(csa_tree_add_7_27_groupi_n_187 ,csa_tree_add_7_27_groupi_n_186);
  not csa_tree_add_7_27_groupi_drc_bufs8139(csa_tree_add_7_27_groupi_n_186 ,csa_tree_add_7_27_groupi_n_966);
  not csa_tree_add_7_27_groupi_drc_bufs8141(csa_tree_add_7_27_groupi_n_185 ,csa_tree_add_7_27_groupi_n_183);
  not csa_tree_add_7_27_groupi_drc_bufs8142(csa_tree_add_7_27_groupi_n_184 ,csa_tree_add_7_27_groupi_n_183);
  not csa_tree_add_7_27_groupi_drc_bufs8143(csa_tree_add_7_27_groupi_n_183 ,csa_tree_add_7_27_groupi_n_813);
  not csa_tree_add_7_27_groupi_drc_bufs8145(csa_tree_add_7_27_groupi_n_182 ,csa_tree_add_7_27_groupi_n_180);
  not csa_tree_add_7_27_groupi_drc_bufs8146(csa_tree_add_7_27_groupi_n_181 ,csa_tree_add_7_27_groupi_n_180);
  not csa_tree_add_7_27_groupi_drc_bufs8147(csa_tree_add_7_27_groupi_n_180 ,csa_tree_add_7_27_groupi_n_940);
  not csa_tree_add_7_27_groupi_drc_bufs8149(csa_tree_add_7_27_groupi_n_179 ,csa_tree_add_7_27_groupi_n_177);
  not csa_tree_add_7_27_groupi_drc_bufs8150(csa_tree_add_7_27_groupi_n_178 ,csa_tree_add_7_27_groupi_n_177);
  not csa_tree_add_7_27_groupi_drc_bufs8151(csa_tree_add_7_27_groupi_n_177 ,csa_tree_add_7_27_groupi_n_942);
  not csa_tree_add_7_27_groupi_drc_bufs8153(csa_tree_add_7_27_groupi_n_176 ,csa_tree_add_7_27_groupi_n_174);
  not csa_tree_add_7_27_groupi_drc_bufs8154(csa_tree_add_7_27_groupi_n_175 ,csa_tree_add_7_27_groupi_n_174);
  not csa_tree_add_7_27_groupi_drc_bufs8155(csa_tree_add_7_27_groupi_n_174 ,csa_tree_add_7_27_groupi_n_941);
  not csa_tree_add_7_27_groupi_drc_bufs8157(csa_tree_add_7_27_groupi_n_173 ,csa_tree_add_7_27_groupi_n_171);
  not csa_tree_add_7_27_groupi_drc_bufs8158(csa_tree_add_7_27_groupi_n_172 ,csa_tree_add_7_27_groupi_n_171);
  not csa_tree_add_7_27_groupi_drc_bufs8159(csa_tree_add_7_27_groupi_n_171 ,csa_tree_add_7_27_groupi_n_589);
  not csa_tree_add_7_27_groupi_drc_bufs8161(csa_tree_add_7_27_groupi_n_170 ,csa_tree_add_7_27_groupi_n_168);
  not csa_tree_add_7_27_groupi_drc_bufs8162(csa_tree_add_7_27_groupi_n_169 ,csa_tree_add_7_27_groupi_n_168);
  not csa_tree_add_7_27_groupi_drc_bufs8163(csa_tree_add_7_27_groupi_n_168 ,csa_tree_add_7_27_groupi_n_569);
  not csa_tree_add_7_27_groupi_drc_bufs8165(csa_tree_add_7_27_groupi_n_167 ,csa_tree_add_7_27_groupi_n_165);
  not csa_tree_add_7_27_groupi_drc_bufs8166(csa_tree_add_7_27_groupi_n_166 ,csa_tree_add_7_27_groupi_n_165);
  not csa_tree_add_7_27_groupi_drc_bufs8167(csa_tree_add_7_27_groupi_n_165 ,csa_tree_add_7_27_groupi_n_583);
  not csa_tree_add_7_27_groupi_drc_bufs8169(csa_tree_add_7_27_groupi_n_164 ,csa_tree_add_7_27_groupi_n_162);
  not csa_tree_add_7_27_groupi_drc_bufs8170(csa_tree_add_7_27_groupi_n_163 ,csa_tree_add_7_27_groupi_n_162);
  not csa_tree_add_7_27_groupi_drc_bufs8171(csa_tree_add_7_27_groupi_n_162 ,csa_tree_add_7_27_groupi_n_907);
  not csa_tree_add_7_27_groupi_drc_bufs8173(csa_tree_add_7_27_groupi_n_161 ,csa_tree_add_7_27_groupi_n_159);
  not csa_tree_add_7_27_groupi_drc_bufs8174(csa_tree_add_7_27_groupi_n_160 ,csa_tree_add_7_27_groupi_n_159);
  not csa_tree_add_7_27_groupi_drc_bufs8175(csa_tree_add_7_27_groupi_n_159 ,csa_tree_add_7_27_groupi_n_943);
  not csa_tree_add_7_27_groupi_drc_bufs8177(csa_tree_add_7_27_groupi_n_158 ,csa_tree_add_7_27_groupi_n_156);
  not csa_tree_add_7_27_groupi_drc_bufs8178(csa_tree_add_7_27_groupi_n_157 ,csa_tree_add_7_27_groupi_n_156);
  not csa_tree_add_7_27_groupi_drc_bufs8179(csa_tree_add_7_27_groupi_n_156 ,csa_tree_add_7_27_groupi_n_964);
  not csa_tree_add_7_27_groupi_drc_bufs8181(csa_tree_add_7_27_groupi_n_155 ,csa_tree_add_7_27_groupi_n_153);
  not csa_tree_add_7_27_groupi_drc_bufs8182(csa_tree_add_7_27_groupi_n_154 ,csa_tree_add_7_27_groupi_n_153);
  not csa_tree_add_7_27_groupi_drc_bufs8183(csa_tree_add_7_27_groupi_n_153 ,csa_tree_add_7_27_groupi_n_583);
  not csa_tree_add_7_27_groupi_drc_bufs8185(csa_tree_add_7_27_groupi_n_152 ,csa_tree_add_7_27_groupi_n_150);
  not csa_tree_add_7_27_groupi_drc_bufs8186(csa_tree_add_7_27_groupi_n_151 ,csa_tree_add_7_27_groupi_n_150);
  not csa_tree_add_7_27_groupi_drc_bufs8187(csa_tree_add_7_27_groupi_n_150 ,csa_tree_add_7_27_groupi_n_587);
  not csa_tree_add_7_27_groupi_drc_bufs8189(csa_tree_add_7_27_groupi_n_149 ,csa_tree_add_7_27_groupi_n_147);
  not csa_tree_add_7_27_groupi_drc_bufs8190(csa_tree_add_7_27_groupi_n_148 ,csa_tree_add_7_27_groupi_n_147);
  not csa_tree_add_7_27_groupi_drc_bufs8191(csa_tree_add_7_27_groupi_n_147 ,csa_tree_add_7_27_groupi_n_589);
  not csa_tree_add_7_27_groupi_drc_bufs8193(csa_tree_add_7_27_groupi_n_146 ,csa_tree_add_7_27_groupi_n_144);
  not csa_tree_add_7_27_groupi_drc_bufs8194(csa_tree_add_7_27_groupi_n_145 ,csa_tree_add_7_27_groupi_n_144);
  not csa_tree_add_7_27_groupi_drc_bufs8195(csa_tree_add_7_27_groupi_n_144 ,csa_tree_add_7_27_groupi_n_943);
  not csa_tree_add_7_27_groupi_drc_bufs8197(csa_tree_add_7_27_groupi_n_143 ,csa_tree_add_7_27_groupi_n_141);
  not csa_tree_add_7_27_groupi_drc_bufs8198(csa_tree_add_7_27_groupi_n_142 ,csa_tree_add_7_27_groupi_n_141);
  not csa_tree_add_7_27_groupi_drc_bufs8199(csa_tree_add_7_27_groupi_n_141 ,csa_tree_add_7_27_groupi_n_942);
  not csa_tree_add_7_27_groupi_drc_bufs8201(csa_tree_add_7_27_groupi_n_140 ,csa_tree_add_7_27_groupi_n_138);
  not csa_tree_add_7_27_groupi_drc_bufs8202(csa_tree_add_7_27_groupi_n_139 ,csa_tree_add_7_27_groupi_n_138);
  not csa_tree_add_7_27_groupi_drc_bufs8203(csa_tree_add_7_27_groupi_n_138 ,csa_tree_add_7_27_groupi_n_966);
  not csa_tree_add_7_27_groupi_drc_bufs8205(csa_tree_add_7_27_groupi_n_137 ,csa_tree_add_7_27_groupi_n_135);
  not csa_tree_add_7_27_groupi_drc_bufs8206(csa_tree_add_7_27_groupi_n_136 ,csa_tree_add_7_27_groupi_n_135);
  not csa_tree_add_7_27_groupi_drc_bufs8207(csa_tree_add_7_27_groupi_n_135 ,csa_tree_add_7_27_groupi_n_587);
  not csa_tree_add_7_27_groupi_drc_bufs8209(csa_tree_add_7_27_groupi_n_134 ,csa_tree_add_7_27_groupi_n_132);
  not csa_tree_add_7_27_groupi_drc_bufs8210(csa_tree_add_7_27_groupi_n_133 ,csa_tree_add_7_27_groupi_n_132);
  not csa_tree_add_7_27_groupi_drc_bufs8211(csa_tree_add_7_27_groupi_n_132 ,csa_tree_add_7_27_groupi_n_585);
  not csa_tree_add_7_27_groupi_drc_bufs8213(csa_tree_add_7_27_groupi_n_131 ,csa_tree_add_7_27_groupi_n_129);
  not csa_tree_add_7_27_groupi_drc_bufs8214(csa_tree_add_7_27_groupi_n_130 ,csa_tree_add_7_27_groupi_n_129);
  not csa_tree_add_7_27_groupi_drc_bufs8215(csa_tree_add_7_27_groupi_n_129 ,csa_tree_add_7_27_groupi_n_577);
  not csa_tree_add_7_27_groupi_drc_bufs8217(csa_tree_add_7_27_groupi_n_128 ,csa_tree_add_7_27_groupi_n_126);
  not csa_tree_add_7_27_groupi_drc_bufs8218(csa_tree_add_7_27_groupi_n_127 ,csa_tree_add_7_27_groupi_n_126);
  not csa_tree_add_7_27_groupi_drc_bufs8219(csa_tree_add_7_27_groupi_n_126 ,csa_tree_add_7_27_groupi_n_569);
  not csa_tree_add_7_27_groupi_drc_bufs8221(csa_tree_add_7_27_groupi_n_125 ,csa_tree_add_7_27_groupi_n_123);
  not csa_tree_add_7_27_groupi_drc_bufs8222(csa_tree_add_7_27_groupi_n_124 ,csa_tree_add_7_27_groupi_n_123);
  not csa_tree_add_7_27_groupi_drc_bufs8223(csa_tree_add_7_27_groupi_n_123 ,csa_tree_add_7_27_groupi_n_573);
  not csa_tree_add_7_27_groupi_drc_bufs8225(csa_tree_add_7_27_groupi_n_122 ,csa_tree_add_7_27_groupi_n_120);
  not csa_tree_add_7_27_groupi_drc_bufs8226(csa_tree_add_7_27_groupi_n_121 ,csa_tree_add_7_27_groupi_n_120);
  not csa_tree_add_7_27_groupi_drc_bufs8227(csa_tree_add_7_27_groupi_n_120 ,csa_tree_add_7_27_groupi_n_575);
  not csa_tree_add_7_27_groupi_drc_bufs8229(csa_tree_add_7_27_groupi_n_119 ,csa_tree_add_7_27_groupi_n_117);
  not csa_tree_add_7_27_groupi_drc_bufs8230(csa_tree_add_7_27_groupi_n_118 ,csa_tree_add_7_27_groupi_n_117);
  not csa_tree_add_7_27_groupi_drc_bufs8231(csa_tree_add_7_27_groupi_n_117 ,csa_tree_add_7_27_groupi_n_571);
  not csa_tree_add_7_27_groupi_drc_bufs8233(csa_tree_add_7_27_groupi_n_116 ,csa_tree_add_7_27_groupi_n_114);
  not csa_tree_add_7_27_groupi_drc_bufs8234(csa_tree_add_7_27_groupi_n_115 ,csa_tree_add_7_27_groupi_n_114);
  not csa_tree_add_7_27_groupi_drc_bufs8235(csa_tree_add_7_27_groupi_n_114 ,csa_tree_add_7_27_groupi_n_754);
  not csa_tree_add_7_27_groupi_drc_bufs8237(csa_tree_add_7_27_groupi_n_113 ,csa_tree_add_7_27_groupi_n_112);
  not csa_tree_add_7_27_groupi_drc_bufs8239(csa_tree_add_7_27_groupi_n_112 ,csa_tree_add_7_27_groupi_n_567);
  not csa_tree_add_7_27_groupi_drc_bufs8241(csa_tree_add_7_27_groupi_n_111 ,csa_tree_add_7_27_groupi_n_109);
  not csa_tree_add_7_27_groupi_drc_bufs8242(csa_tree_add_7_27_groupi_n_110 ,csa_tree_add_7_27_groupi_n_109);
  not csa_tree_add_7_27_groupi_drc_bufs8243(csa_tree_add_7_27_groupi_n_109 ,csa_tree_add_7_27_groupi_n_754);
  not csa_tree_add_7_27_groupi_drc_bufs8245(csa_tree_add_7_27_groupi_n_108 ,csa_tree_add_7_27_groupi_n_107);
  not csa_tree_add_7_27_groupi_drc_bufs8247(csa_tree_add_7_27_groupi_n_107 ,csa_tree_add_7_27_groupi_n_566);
  not csa_tree_add_7_27_groupi_drc_bufs8249(csa_tree_add_7_27_groupi_n_106 ,csa_tree_add_7_27_groupi_n_105);
  not csa_tree_add_7_27_groupi_drc_bufs8251(csa_tree_add_7_27_groupi_n_105 ,csa_tree_add_7_27_groupi_n_468);
  not csa_tree_add_7_27_groupi_drc_bufs8253(csa_tree_add_7_27_groupi_n_104 ,csa_tree_add_7_27_groupi_n_103);
  not csa_tree_add_7_27_groupi_drc_bufs8255(csa_tree_add_7_27_groupi_n_103 ,csa_tree_add_7_27_groupi_n_465);
  not csa_tree_add_7_27_groupi_drc_bufs8257(csa_tree_add_7_27_groupi_n_102 ,csa_tree_add_7_27_groupi_n_101);
  not csa_tree_add_7_27_groupi_drc_bufs8259(csa_tree_add_7_27_groupi_n_101 ,csa_tree_add_7_27_groupi_n_459);
  not csa_tree_add_7_27_groupi_drc_bufs8261(csa_tree_add_7_27_groupi_n_100 ,csa_tree_add_7_27_groupi_n_99);
  not csa_tree_add_7_27_groupi_drc_bufs8263(csa_tree_add_7_27_groupi_n_99 ,csa_tree_add_7_27_groupi_n_456);
  not csa_tree_add_7_27_groupi_drc_bufs8265(csa_tree_add_7_27_groupi_n_98 ,csa_tree_add_7_27_groupi_n_97);
  not csa_tree_add_7_27_groupi_drc_bufs8267(csa_tree_add_7_27_groupi_n_97 ,csa_tree_add_7_27_groupi_n_462);
  not csa_tree_add_7_27_groupi_drc_bufs8269(csa_tree_add_7_27_groupi_n_96 ,csa_tree_add_7_27_groupi_n_95);
  not csa_tree_add_7_27_groupi_drc_bufs8271(csa_tree_add_7_27_groupi_n_95 ,csa_tree_add_7_27_groupi_n_378);
  not csa_tree_add_7_27_groupi_drc_bufs8273(csa_tree_add_7_27_groupi_n_94 ,csa_tree_add_7_27_groupi_n_92);
  not csa_tree_add_7_27_groupi_drc_bufs8274(csa_tree_add_7_27_groupi_n_93 ,csa_tree_add_7_27_groupi_n_92);
  not csa_tree_add_7_27_groupi_drc_bufs8275(csa_tree_add_7_27_groupi_n_92 ,csa_tree_add_7_27_groupi_n_646);
  not csa_tree_add_7_27_groupi_drc_bufs8277(csa_tree_add_7_27_groupi_n_91 ,csa_tree_add_7_27_groupi_n_90);
  not csa_tree_add_7_27_groupi_drc_bufs8279(csa_tree_add_7_27_groupi_n_90 ,csa_tree_add_7_27_groupi_n_383);
  not csa_tree_add_7_27_groupi_drc_bufs8281(csa_tree_add_7_27_groupi_n_89 ,csa_tree_add_7_27_groupi_n_87);
  not csa_tree_add_7_27_groupi_drc_bufs8282(csa_tree_add_7_27_groupi_n_88 ,csa_tree_add_7_27_groupi_n_87);
  not csa_tree_add_7_27_groupi_drc_bufs8283(csa_tree_add_7_27_groupi_n_87 ,csa_tree_add_7_27_groupi_n_610);
  not csa_tree_add_7_27_groupi_drc_bufs8285(csa_tree_add_7_27_groupi_n_86 ,csa_tree_add_7_27_groupi_n_84);
  not csa_tree_add_7_27_groupi_drc_bufs8286(csa_tree_add_7_27_groupi_n_85 ,csa_tree_add_7_27_groupi_n_84);
  not csa_tree_add_7_27_groupi_drc_bufs8287(csa_tree_add_7_27_groupi_n_84 ,csa_tree_add_7_27_groupi_n_631);
  not csa_tree_add_7_27_groupi_drc_bufs8289(csa_tree_add_7_27_groupi_n_83 ,csa_tree_add_7_27_groupi_n_82);
  not csa_tree_add_7_27_groupi_drc_bufs8291(csa_tree_add_7_27_groupi_n_82 ,csa_tree_add_7_27_groupi_n_372);
  not csa_tree_add_7_27_groupi_drc_bufs8293(csa_tree_add_7_27_groupi_n_81 ,csa_tree_add_7_27_groupi_n_80);
  not csa_tree_add_7_27_groupi_drc_bufs8295(csa_tree_add_7_27_groupi_n_80 ,csa_tree_add_7_27_groupi_n_393);
  not csa_tree_add_7_27_groupi_drc_bufs8297(csa_tree_add_7_27_groupi_n_79 ,csa_tree_add_7_27_groupi_n_77);
  not csa_tree_add_7_27_groupi_drc_bufs8298(csa_tree_add_7_27_groupi_n_78 ,csa_tree_add_7_27_groupi_n_77);
  not csa_tree_add_7_27_groupi_drc_bufs8299(csa_tree_add_7_27_groupi_n_77 ,csa_tree_add_7_27_groupi_n_613);
  not csa_tree_add_7_27_groupi_drc_bufs8301(csa_tree_add_7_27_groupi_n_76 ,csa_tree_add_7_27_groupi_n_75);
  not csa_tree_add_7_27_groupi_drc_bufs8303(csa_tree_add_7_27_groupi_n_75 ,csa_tree_add_7_27_groupi_n_398);
  not csa_tree_add_7_27_groupi_drc_bufs8305(csa_tree_add_7_27_groupi_n_74 ,csa_tree_add_7_27_groupi_n_73);
  not csa_tree_add_7_27_groupi_drc_bufs8307(csa_tree_add_7_27_groupi_n_73 ,csa_tree_add_7_27_groupi_n_401);
  not csa_tree_add_7_27_groupi_drc_bufs8309(csa_tree_add_7_27_groupi_n_72 ,csa_tree_add_7_27_groupi_n_70);
  not csa_tree_add_7_27_groupi_drc_bufs8310(csa_tree_add_7_27_groupi_n_71 ,csa_tree_add_7_27_groupi_n_70);
  not csa_tree_add_7_27_groupi_drc_bufs8311(csa_tree_add_7_27_groupi_n_70 ,csa_tree_add_7_27_groupi_n_616);
  not csa_tree_add_7_27_groupi_drc_bufs8313(csa_tree_add_7_27_groupi_n_69 ,csa_tree_add_7_27_groupi_n_67);
  not csa_tree_add_7_27_groupi_drc_bufs8314(csa_tree_add_7_27_groupi_n_68 ,csa_tree_add_7_27_groupi_n_67);
  not csa_tree_add_7_27_groupi_drc_bufs8315(csa_tree_add_7_27_groupi_n_67 ,csa_tree_add_7_27_groupi_n_634);
  not csa_tree_add_7_27_groupi_drc_bufs8317(csa_tree_add_7_27_groupi_n_66 ,csa_tree_add_7_27_groupi_n_64);
  not csa_tree_add_7_27_groupi_drc_bufs8318(csa_tree_add_7_27_groupi_n_65 ,csa_tree_add_7_27_groupi_n_64);
  not csa_tree_add_7_27_groupi_drc_bufs8319(csa_tree_add_7_27_groupi_n_64 ,csa_tree_add_7_27_groupi_n_649);
  not csa_tree_add_7_27_groupi_drc_bufs8321(csa_tree_add_7_27_groupi_n_63 ,csa_tree_add_7_27_groupi_n_62);
  not csa_tree_add_7_27_groupi_drc_bufs8323(csa_tree_add_7_27_groupi_n_62 ,csa_tree_add_7_27_groupi_n_410);
  not csa_tree_add_7_27_groupi_drc_bufs8325(csa_tree_add_7_27_groupi_n_61 ,csa_tree_add_7_27_groupi_n_60);
  not csa_tree_add_7_27_groupi_drc_bufs8327(csa_tree_add_7_27_groupi_n_60 ,csa_tree_add_7_27_groupi_n_413);
  not csa_tree_add_7_27_groupi_drc_bufs8329(csa_tree_add_7_27_groupi_n_59 ,csa_tree_add_7_27_groupi_n_57);
  not csa_tree_add_7_27_groupi_drc_bufs8330(csa_tree_add_7_27_groupi_n_58 ,csa_tree_add_7_27_groupi_n_57);
  not csa_tree_add_7_27_groupi_drc_bufs8331(csa_tree_add_7_27_groupi_n_57 ,csa_tree_add_7_27_groupi_n_619);
  not csa_tree_add_7_27_groupi_drc_bufs8333(csa_tree_add_7_27_groupi_n_56 ,csa_tree_add_7_27_groupi_n_55);
  not csa_tree_add_7_27_groupi_drc_bufs8335(csa_tree_add_7_27_groupi_n_55 ,csa_tree_add_7_27_groupi_n_418);
  not csa_tree_add_7_27_groupi_drc_bufs8337(csa_tree_add_7_27_groupi_n_54 ,csa_tree_add_7_27_groupi_n_52);
  not csa_tree_add_7_27_groupi_drc_bufs8338(csa_tree_add_7_27_groupi_n_53 ,csa_tree_add_7_27_groupi_n_52);
  not csa_tree_add_7_27_groupi_drc_bufs8339(csa_tree_add_7_27_groupi_n_52 ,csa_tree_add_7_27_groupi_n_607);
  not csa_tree_add_7_27_groupi_drc_bufs8341(csa_tree_add_7_27_groupi_n_51 ,csa_tree_add_7_27_groupi_n_49);
  not csa_tree_add_7_27_groupi_drc_bufs8342(csa_tree_add_7_27_groupi_n_50 ,csa_tree_add_7_27_groupi_n_49);
  not csa_tree_add_7_27_groupi_drc_bufs8343(csa_tree_add_7_27_groupi_n_49 ,csa_tree_add_7_27_groupi_n_622);
  not csa_tree_add_7_27_groupi_drc_bufs8345(csa_tree_add_7_27_groupi_n_48 ,csa_tree_add_7_27_groupi_n_46);
  not csa_tree_add_7_27_groupi_drc_bufs8346(csa_tree_add_7_27_groupi_n_47 ,csa_tree_add_7_27_groupi_n_46);
  not csa_tree_add_7_27_groupi_drc_bufs8347(csa_tree_add_7_27_groupi_n_46 ,csa_tree_add_7_27_groupi_n_637);
  not csa_tree_add_7_27_groupi_drc_bufs8349(csa_tree_add_7_27_groupi_n_45 ,csa_tree_add_7_27_groupi_n_43);
  not csa_tree_add_7_27_groupi_drc_bufs8350(csa_tree_add_7_27_groupi_n_44 ,csa_tree_add_7_27_groupi_n_43);
  not csa_tree_add_7_27_groupi_drc_bufs8351(csa_tree_add_7_27_groupi_n_43 ,csa_tree_add_7_27_groupi_n_598);
  not csa_tree_add_7_27_groupi_drc_bufs8353(csa_tree_add_7_27_groupi_n_42 ,csa_tree_add_7_27_groupi_n_41);
  not csa_tree_add_7_27_groupi_drc_bufs8355(csa_tree_add_7_27_groupi_n_41 ,csa_tree_add_7_27_groupi_n_390);
  not csa_tree_add_7_27_groupi_drc_bufs8357(csa_tree_add_7_27_groupi_n_40 ,csa_tree_add_7_27_groupi_n_39);
  not csa_tree_add_7_27_groupi_drc_bufs8359(csa_tree_add_7_27_groupi_n_39 ,csa_tree_add_7_27_groupi_n_433);
  not csa_tree_add_7_27_groupi_drc_bufs8361(csa_tree_add_7_27_groupi_n_38 ,csa_tree_add_7_27_groupi_n_36);
  not csa_tree_add_7_27_groupi_drc_bufs8362(csa_tree_add_7_27_groupi_n_37 ,csa_tree_add_7_27_groupi_n_36);
  not csa_tree_add_7_27_groupi_drc_bufs8363(csa_tree_add_7_27_groupi_n_36 ,csa_tree_add_7_27_groupi_n_625);
  not csa_tree_add_7_27_groupi_drc_bufs8365(csa_tree_add_7_27_groupi_n_35 ,csa_tree_add_7_27_groupi_n_33);
  not csa_tree_add_7_27_groupi_drc_bufs8366(csa_tree_add_7_27_groupi_n_34 ,csa_tree_add_7_27_groupi_n_33);
  not csa_tree_add_7_27_groupi_drc_bufs8367(csa_tree_add_7_27_groupi_n_33 ,csa_tree_add_7_27_groupi_n_640);
  not csa_tree_add_7_27_groupi_drc_bufs8369(csa_tree_add_7_27_groupi_n_32 ,csa_tree_add_7_27_groupi_n_30);
  not csa_tree_add_7_27_groupi_drc_bufs8370(csa_tree_add_7_27_groupi_n_31 ,csa_tree_add_7_27_groupi_n_30);
  not csa_tree_add_7_27_groupi_drc_bufs8371(csa_tree_add_7_27_groupi_n_30 ,csa_tree_add_7_27_groupi_n_601);
  not csa_tree_add_7_27_groupi_drc_bufs8373(csa_tree_add_7_27_groupi_n_29 ,csa_tree_add_7_27_groupi_n_27);
  not csa_tree_add_7_27_groupi_drc_bufs8374(csa_tree_add_7_27_groupi_n_28 ,csa_tree_add_7_27_groupi_n_27);
  not csa_tree_add_7_27_groupi_drc_bufs8375(csa_tree_add_7_27_groupi_n_27 ,csa_tree_add_7_27_groupi_n_604);
  not csa_tree_add_7_27_groupi_drc_bufs8377(csa_tree_add_7_27_groupi_n_26 ,csa_tree_add_7_27_groupi_n_25);
  not csa_tree_add_7_27_groupi_drc_bufs8379(csa_tree_add_7_27_groupi_n_25 ,csa_tree_add_7_27_groupi_n_421);
  not csa_tree_add_7_27_groupi_drc_bufs8381(csa_tree_add_7_27_groupi_n_24 ,csa_tree_add_7_27_groupi_n_23);
  not csa_tree_add_7_27_groupi_drc_bufs8383(csa_tree_add_7_27_groupi_n_23 ,csa_tree_add_7_27_groupi_n_428);
  not csa_tree_add_7_27_groupi_drc_bufs8385(csa_tree_add_7_27_groupi_n_22 ,csa_tree_add_7_27_groupi_n_21);
  not csa_tree_add_7_27_groupi_drc_bufs8387(csa_tree_add_7_27_groupi_n_21 ,csa_tree_add_7_27_groupi_n_447);
  not csa_tree_add_7_27_groupi_drc_bufs8389(csa_tree_add_7_27_groupi_n_20 ,csa_tree_add_7_27_groupi_n_18);
  not csa_tree_add_7_27_groupi_drc_bufs8390(csa_tree_add_7_27_groupi_n_19 ,csa_tree_add_7_27_groupi_n_18);
  not csa_tree_add_7_27_groupi_drc_bufs8391(csa_tree_add_7_27_groupi_n_18 ,csa_tree_add_7_27_groupi_n_628);
  not csa_tree_add_7_27_groupi_drc_bufs8393(csa_tree_add_7_27_groupi_n_17 ,csa_tree_add_7_27_groupi_n_16);
  not csa_tree_add_7_27_groupi_drc_bufs8395(csa_tree_add_7_27_groupi_n_16 ,csa_tree_add_7_27_groupi_n_643);
  not csa_tree_add_7_27_groupi_drc_bufs8397(csa_tree_add_7_27_groupi_n_15 ,csa_tree_add_7_27_groupi_n_14);
  not csa_tree_add_7_27_groupi_drc_bufs8399(csa_tree_add_7_27_groupi_n_14 ,csa_tree_add_7_27_groupi_n_444);
  not csa_tree_add_7_27_groupi_drc_bufs8401(csa_tree_add_7_27_groupi_n_13 ,csa_tree_add_7_27_groupi_n_12);
  not csa_tree_add_7_27_groupi_drc_bufs8403(csa_tree_add_7_27_groupi_n_12 ,csa_tree_add_7_27_groupi_n_375);
  not csa_tree_add_7_27_groupi_drc_bufs8405(csa_tree_add_7_27_groupi_n_11 ,csa_tree_add_7_27_groupi_n_9);
  not csa_tree_add_7_27_groupi_drc_bufs8406(csa_tree_add_7_27_groupi_n_10 ,csa_tree_add_7_27_groupi_n_9);
  not csa_tree_add_7_27_groupi_drc_bufs8407(csa_tree_add_7_27_groupi_n_9 ,csa_tree_add_7_27_groupi_n_591);
  not csa_tree_add_7_27_groupi_drc_bufs8409(csa_tree_add_7_27_groupi_n_8 ,csa_tree_add_7_27_groupi_n_6);
  not csa_tree_add_7_27_groupi_drc_bufs8410(csa_tree_add_7_27_groupi_n_7 ,csa_tree_add_7_27_groupi_n_6);
  not csa_tree_add_7_27_groupi_drc_bufs8411(csa_tree_add_7_27_groupi_n_6 ,csa_tree_add_7_27_groupi_n_594);
  xor csa_tree_add_7_27_groupi_g2(n_29 ,csa_tree_add_7_27_groupi_n_2342 ,csa_tree_add_7_27_groupi_n_2303);
  xor csa_tree_add_7_27_groupi_g8413(n_28 ,csa_tree_add_7_27_groupi_n_2340 ,csa_tree_add_7_27_groupi_n_2302);
  xor csa_tree_add_7_27_groupi_g8414(csa_tree_add_7_27_groupi_n_3 ,csa_tree_add_7_27_groupi_n_1171 ,csa_tree_add_7_27_groupi_n_1299);
  xor csa_tree_add_7_27_groupi_g8415(csa_tree_add_7_27_groupi_n_2 ,csa_tree_add_7_27_groupi_n_1168 ,csa_tree_add_7_27_groupi_n_1173);
  xor csa_tree_add_7_27_groupi_g8416(csa_tree_add_7_27_groupi_n_1 ,csa_tree_add_7_27_groupi_n_969 ,in3[15]);
  and csa_tree_add_7_27_groupi_g8417(csa_tree_add_7_27_groupi_n_0 ,csa_tree_add_7_27_groupi_n_16 ,csa_tree_add_7_27_groupi_n_528);
  xor dec_sub_8_33_g369(out2[31] ,dec_sub_8_33_n_150 ,n_33);
  xor dec_sub_8_33_g370(out2[30] ,dec_sub_8_33_n_147 ,dec_sub_8_33_n_30);
  nor dec_sub_8_33_g371(dec_sub_8_33_n_150 ,dec_sub_8_33_n_30 ,dec_sub_8_33_n_146);
  or dec_sub_8_33_g372(out2[29] ,dec_sub_8_33_n_148 ,dec_sub_8_33_n_147);
  and dec_sub_8_33_g373(dec_sub_8_33_n_148 ,dec_sub_8_33_n_11 ,dec_sub_8_33_n_143);
  not dec_sub_8_33_g374(dec_sub_8_33_n_146 ,dec_sub_8_33_n_147);
  and dec_sub_8_33_g375(dec_sub_8_33_n_147 ,dec_sub_8_33_n_62 ,dec_sub_8_33_n_144);
  xor dec_sub_8_33_g376(out2[28] ,dec_sub_8_33_n_141 ,dec_sub_8_33_n_20);
  not dec_sub_8_33_g377(dec_sub_8_33_n_144 ,dec_sub_8_33_n_143);
  or dec_sub_8_33_g378(dec_sub_8_33_n_143 ,dec_sub_8_33_n_20 ,dec_sub_8_33_n_140);
  or dec_sub_8_33_g379(out2[27] ,dec_sub_8_33_n_6 ,dec_sub_8_33_n_141);
  not dec_sub_8_33_g381(dec_sub_8_33_n_140 ,dec_sub_8_33_n_141);
  and dec_sub_8_33_g382(dec_sub_8_33_n_141 ,dec_sub_8_33_n_60 ,dec_sub_8_33_n_138);
  xor dec_sub_8_33_g384(out2[25] ,dec_sub_8_33_n_137 ,dec_sub_8_33_n_13);
  and dec_sub_8_33_g386(dec_sub_8_33_n_138 ,dec_sub_8_33_n_58 ,dec_sub_8_33_n_136);
  nor dec_sub_8_33_g388(dec_sub_8_33_n_137 ,dec_sub_8_33_n_54 ,dec_sub_8_33_n_132);
  not dec_sub_8_33_g389(dec_sub_8_33_n_136 ,dec_sub_8_33_n_135);
  or dec_sub_8_33_g390(dec_sub_8_33_n_135 ,dec_sub_8_33_n_70 ,dec_sub_8_33_n_132);
  or dec_sub_8_33_g391(out2[23] ,dec_sub_8_33_n_131 ,dec_sub_8_33_n_133);
  not dec_sub_8_33_g392(dec_sub_8_33_n_132 ,dec_sub_8_33_n_133);
  and dec_sub_8_33_g393(dec_sub_8_33_n_133 ,dec_sub_8_33_n_65 ,dec_sub_8_33_n_128);
  nor dec_sub_8_33_g394(dec_sub_8_33_n_131 ,dec_sub_8_33_n_65 ,dec_sub_8_33_n_128);
  xor dec_sub_8_33_g396(out2[21] ,dec_sub_8_33_n_124 ,dec_sub_8_33_n_34);
  xor dec_sub_8_33_g397(out2[19] ,dec_sub_8_33_n_122 ,dec_sub_8_33_n_26);
  and dec_sub_8_33_g398(dec_sub_8_33_n_128 ,dec_sub_8_33_n_64 ,dec_sub_8_33_n_123);
  xnor dec_sub_8_33_g399(out2[20] ,dec_sub_8_33_n_118 ,dec_sub_8_33_n_46);
  xnor dec_sub_8_33_g400(out2[18] ,dec_sub_8_33_n_119 ,dec_sub_8_33_n_52);
  xor dec_sub_8_33_g401(out2[17] ,dec_sub_8_33_n_120 ,dec_sub_8_33_n_18);
  nor dec_sub_8_33_g402(dec_sub_8_33_n_124 ,dec_sub_8_33_n_45 ,dec_sub_8_33_n_118);
  and dec_sub_8_33_g404(dec_sub_8_33_n_123 ,dec_sub_8_33_n_71 ,dec_sub_8_33_n_117);
  nor dec_sub_8_33_g405(dec_sub_8_33_n_122 ,dec_sub_8_33_n_51 ,dec_sub_8_33_n_119);
  xnor dec_sub_8_33_g406(out2[16] ,dec_sub_8_33_n_36 ,dec_sub_8_33_n_114);
  nor dec_sub_8_33_g407(dec_sub_8_33_n_120 ,dec_sub_8_33_n_37 ,dec_sub_8_33_n_10);
  or dec_sub_8_33_g408(dec_sub_8_33_n_119 ,dec_sub_8_33_n_74 ,dec_sub_8_33_n_10);
  not dec_sub_8_33_g409(dec_sub_8_33_n_118 ,dec_sub_8_33_n_117);
  and dec_sub_8_33_g410(dec_sub_8_33_n_117 ,dec_sub_8_33_n_86 ,dec_sub_8_33_n_115);
  or dec_sub_8_33_g411(out2[15] ,dec_sub_8_33_n_113 ,dec_sub_8_33_n_115);
  not dec_sub_8_33_g412(dec_sub_8_33_n_114 ,dec_sub_8_33_n_115);
  and dec_sub_8_33_g413(dec_sub_8_33_n_115 ,dec_sub_8_33_n_67 ,dec_sub_8_33_n_110);
  nor dec_sub_8_33_g414(dec_sub_8_33_n_113 ,dec_sub_8_33_n_67 ,dec_sub_8_33_n_110);
  xor dec_sub_8_33_g416(out2[13] ,dec_sub_8_33_n_105 ,dec_sub_8_33_n_32);
  xor dec_sub_8_33_g417(out2[11] ,dec_sub_8_33_n_104 ,dec_sub_8_33_n_22);
  and dec_sub_8_33_g418(dec_sub_8_33_n_110 ,dec_sub_8_33_n_61 ,dec_sub_8_33_n_106);
  xnor dec_sub_8_33_g419(out2[12] ,dec_sub_8_33_n_101 ,dec_sub_8_33_n_43);
  xnor dec_sub_8_33_g420(out2[10] ,dec_sub_8_33_n_99 ,dec_sub_8_33_n_49);
  xor dec_sub_8_33_g421(out2[9] ,dec_sub_8_33_n_102 ,dec_sub_8_33_n_24);
  and dec_sub_8_33_g423(dec_sub_8_33_n_106 ,dec_sub_8_33_n_69 ,dec_sub_8_33_n_100);
  nor dec_sub_8_33_g424(dec_sub_8_33_n_105 ,dec_sub_8_33_n_42 ,dec_sub_8_33_n_101);
  nor dec_sub_8_33_g425(dec_sub_8_33_n_104 ,dec_sub_8_33_n_48 ,dec_sub_8_33_n_99);
  xnor dec_sub_8_33_g426(out2[8] ,dec_sub_8_33_n_39 ,dec_sub_8_33_n_96);
  nor dec_sub_8_33_g427(dec_sub_8_33_n_102 ,dec_sub_8_33_n_40 ,dec_sub_8_33_n_8);
  not dec_sub_8_33_g428(dec_sub_8_33_n_101 ,dec_sub_8_33_n_100);
  and dec_sub_8_33_g429(dec_sub_8_33_n_100 ,dec_sub_8_33_n_87 ,dec_sub_8_33_n_97);
  or dec_sub_8_33_g430(dec_sub_8_33_n_99 ,dec_sub_8_33_n_73 ,dec_sub_8_33_n_8);
  or dec_sub_8_33_g431(out2[7] ,dec_sub_8_33_n_3 ,dec_sub_8_33_n_97);
  not dec_sub_8_33_g433(dec_sub_8_33_n_96 ,dec_sub_8_33_n_97);
  and dec_sub_8_33_g434(dec_sub_8_33_n_97 ,dec_sub_8_33_n_59 ,dec_sub_8_33_n_93);
  xnor dec_sub_8_33_g435(out2[6] ,dec_sub_8_33_n_90 ,n_8);
  xor dec_sub_8_33_g436(out2[5] ,dec_sub_8_33_n_92 ,dec_sub_8_33_n_16);
  and dec_sub_8_33_g438(dec_sub_8_33_n_93 ,dec_sub_8_33_n_68 ,dec_sub_8_33_n_91);
  nor dec_sub_8_33_g440(dec_sub_8_33_n_92 ,dec_sub_8_33_n_56 ,dec_sub_8_33_n_84);
  not dec_sub_8_33_g441(dec_sub_8_33_n_91 ,dec_sub_8_33_n_90);
  or dec_sub_8_33_g442(dec_sub_8_33_n_90 ,dec_sub_8_33_n_72 ,dec_sub_8_33_n_84);
  or dec_sub_8_33_g443(out2[3] ,dec_sub_8_33_n_88 ,dec_sub_8_33_n_85);
  and dec_sub_8_33_g444(dec_sub_8_33_n_88 ,dec_sub_8_33_n_14 ,dec_sub_8_33_n_79);
  nor dec_sub_8_33_g445(dec_sub_8_33_n_87 ,dec_sub_8_33_n_49 ,dec_sub_8_33_n_82);
  nor dec_sub_8_33_g446(dec_sub_8_33_n_86 ,dec_sub_8_33_n_52 ,dec_sub_8_33_n_81);
  not dec_sub_8_33_g447(dec_sub_8_33_n_84 ,dec_sub_8_33_n_85);
  and dec_sub_8_33_g448(dec_sub_8_33_n_85 ,dec_sub_8_33_n_57 ,dec_sub_8_33_n_80);
  xor dec_sub_8_33_g449(out2[2] ,dec_sub_8_33_n_77 ,dec_sub_8_33_n_28);
  or dec_sub_8_33_g450(dec_sub_8_33_n_82 ,dec_sub_8_33_n_22 ,dec_sub_8_33_n_73);
  or dec_sub_8_33_g451(dec_sub_8_33_n_81 ,dec_sub_8_33_n_26 ,dec_sub_8_33_n_74);
  not dec_sub_8_33_g452(dec_sub_8_33_n_80 ,dec_sub_8_33_n_79);
  or dec_sub_8_33_g453(dec_sub_8_33_n_79 ,dec_sub_8_33_n_28 ,dec_sub_8_33_n_76);
  or dec_sub_8_33_g454(out2[1] ,dec_sub_8_33_n_75 ,dec_sub_8_33_n_77);
  not dec_sub_8_33_g455(dec_sub_8_33_n_76 ,dec_sub_8_33_n_77);
  and dec_sub_8_33_g456(dec_sub_8_33_n_77 ,dec_sub_8_33_n_63 ,dec_sub_8_33_n_66);
  nor dec_sub_8_33_g457(dec_sub_8_33_n_75 ,dec_sub_8_33_n_63 ,dec_sub_8_33_n_66);
  or dec_sub_8_33_g458(dec_sub_8_33_n_74 ,dec_sub_8_33_n_18 ,dec_sub_8_33_n_36);
  or dec_sub_8_33_g459(dec_sub_8_33_n_73 ,dec_sub_8_33_n_24 ,dec_sub_8_33_n_39);
  or dec_sub_8_33_g460(dec_sub_8_33_n_72 ,dec_sub_8_33_n_16 ,dec_sub_8_33_n_56);
  nor dec_sub_8_33_g461(dec_sub_8_33_n_71 ,dec_sub_8_33_n_34 ,dec_sub_8_33_n_46);
  or dec_sub_8_33_g462(dec_sub_8_33_n_70 ,dec_sub_8_33_n_13 ,dec_sub_8_33_n_54);
  nor dec_sub_8_33_g463(dec_sub_8_33_n_69 ,dec_sub_8_33_n_32 ,dec_sub_8_33_n_43);
  not dec_sub_8_33_g467(dec_sub_8_33_n_68 ,n_8);
  not dec_sub_8_33_g468(dec_sub_8_33_n_67 ,n_17);
  not dec_sub_8_33_g469(dec_sub_8_33_n_66 ,n_2);
  not dec_sub_8_33_g470(dec_sub_8_33_n_65 ,n_25);
  not dec_sub_8_33_g473(dec_sub_8_33_n_64 ,n_24);
  not dec_sub_8_33_g474(dec_sub_8_33_n_63 ,n_3);
  not dec_sub_8_33_drc_bufs(dec_sub_8_33_n_56 ,dec_sub_8_33_n_55);
  not dec_sub_8_33_drc_bufs477(dec_sub_8_33_n_55 ,n_6);
  not dec_sub_8_33_drc_bufs479(dec_sub_8_33_n_54 ,dec_sub_8_33_n_53);
  not dec_sub_8_33_drc_bufs481(dec_sub_8_33_n_53 ,n_26);
  not dec_sub_8_33_drc_bufs483(dec_sub_8_33_n_52 ,dec_sub_8_33_n_50);
  not dec_sub_8_33_drc_bufs484(dec_sub_8_33_n_51 ,dec_sub_8_33_n_50);
  not dec_sub_8_33_drc_bufs485(dec_sub_8_33_n_50 ,n_20);
  not dec_sub_8_33_drc_bufs487(dec_sub_8_33_n_49 ,dec_sub_8_33_n_47);
  not dec_sub_8_33_drc_bufs488(dec_sub_8_33_n_48 ,dec_sub_8_33_n_47);
  not dec_sub_8_33_drc_bufs489(dec_sub_8_33_n_47 ,n_12);
  not dec_sub_8_33_drc_bufs491(dec_sub_8_33_n_46 ,dec_sub_8_33_n_44);
  not dec_sub_8_33_drc_bufs492(dec_sub_8_33_n_45 ,dec_sub_8_33_n_44);
  not dec_sub_8_33_drc_bufs493(dec_sub_8_33_n_44 ,n_22);
  not dec_sub_8_33_drc_bufs495(dec_sub_8_33_n_43 ,dec_sub_8_33_n_41);
  not dec_sub_8_33_drc_bufs496(dec_sub_8_33_n_42 ,dec_sub_8_33_n_41);
  not dec_sub_8_33_drc_bufs497(dec_sub_8_33_n_41 ,n_14);
  not dec_sub_8_33_drc_bufs499(dec_sub_8_33_n_40 ,dec_sub_8_33_n_38);
  not dec_sub_8_33_drc_bufs500(dec_sub_8_33_n_39 ,dec_sub_8_33_n_38);
  not dec_sub_8_33_drc_bufs501(dec_sub_8_33_n_38 ,n_10);
  not dec_sub_8_33_drc_bufs503(dec_sub_8_33_n_37 ,dec_sub_8_33_n_35);
  not dec_sub_8_33_drc_bufs504(dec_sub_8_33_n_36 ,dec_sub_8_33_n_35);
  not dec_sub_8_33_drc_bufs505(dec_sub_8_33_n_35 ,n_18);
  not dec_sub_8_33_drc_bufs507(dec_sub_8_33_n_34 ,dec_sub_8_33_n_33);
  not dec_sub_8_33_drc_bufs509(dec_sub_8_33_n_33 ,n_23);
  not dec_sub_8_33_drc_bufs511(dec_sub_8_33_n_32 ,dec_sub_8_33_n_31);
  not dec_sub_8_33_drc_bufs513(dec_sub_8_33_n_31 ,n_15);
  not dec_sub_8_33_drc_bufs515(dec_sub_8_33_n_30 ,dec_sub_8_33_n_29);
  not dec_sub_8_33_drc_bufs517(dec_sub_8_33_n_29 ,n_32);
  not dec_sub_8_33_drc_bufs521(dec_sub_8_33_n_61 ,n_16);
  not dec_sub_8_33_drc_bufs523(dec_sub_8_33_n_28 ,dec_sub_8_33_n_27);
  not dec_sub_8_33_drc_bufs525(dec_sub_8_33_n_27 ,n_4);
  not dec_sub_8_33_drc_bufs527(dec_sub_8_33_n_26 ,dec_sub_8_33_n_25);
  not dec_sub_8_33_drc_bufs529(dec_sub_8_33_n_25 ,n_21);
  not dec_sub_8_33_drc_bufs531(dec_sub_8_33_n_24 ,dec_sub_8_33_n_23);
  not dec_sub_8_33_drc_bufs533(dec_sub_8_33_n_23 ,n_11);
  not dec_sub_8_33_drc_bufs535(dec_sub_8_33_n_22 ,dec_sub_8_33_n_21);
  not dec_sub_8_33_drc_bufs537(dec_sub_8_33_n_21 ,n_13);
  not dec_sub_8_33_drc_bufs539(dec_sub_8_33_n_20 ,dec_sub_8_33_n_19);
  not dec_sub_8_33_drc_bufs541(dec_sub_8_33_n_19 ,n_30);
  not dec_sub_8_33_drc_bufs543(dec_sub_8_33_n_18 ,dec_sub_8_33_n_17);
  not dec_sub_8_33_drc_bufs545(dec_sub_8_33_n_17 ,n_19);
  not dec_sub_8_33_drc_bufs549(dec_sub_8_33_n_59 ,n_9);
  not dec_sub_8_33_drc_bufs553(dec_sub_8_33_n_60 ,n_29);
  not dec_sub_8_33_drc_bufs555(dec_sub_8_33_n_16 ,dec_sub_8_33_n_15);
  not dec_sub_8_33_drc_bufs557(dec_sub_8_33_n_15 ,n_7);
  not dec_sub_8_33_drc_bufs561(dec_sub_8_33_n_58 ,n_28);
  not dec_sub_8_33_drc_bufs564(dec_sub_8_33_n_14 ,dec_sub_8_33_n_57);
  not dec_sub_8_33_drc_bufs565(dec_sub_8_33_n_57 ,n_5);
  not dec_sub_8_33_drc_bufs567(dec_sub_8_33_n_13 ,dec_sub_8_33_n_12);
  not dec_sub_8_33_drc_bufs569(dec_sub_8_33_n_12 ,n_27);
  not dec_sub_8_33_drc_bufs572(dec_sub_8_33_n_11 ,dec_sub_8_33_n_62);
  not dec_sub_8_33_drc_bufs573(dec_sub_8_33_n_62 ,n_31);
  not dec_sub_8_33_drc_bufs576(dec_sub_8_33_n_10 ,dec_sub_8_33_n_9);
  not dec_sub_8_33_drc_bufs578(dec_sub_8_33_n_9 ,dec_sub_8_33_n_114);
  not dec_sub_8_33_drc_bufs580(dec_sub_8_33_n_8 ,dec_sub_8_33_n_7);
  not dec_sub_8_33_drc_bufs582(dec_sub_8_33_n_7 ,dec_sub_8_33_n_96);
  nor dec_sub_8_33_g2(dec_sub_8_33_n_6 ,dec_sub_8_33_n_60 ,dec_sub_8_33_n_138);
  xor dec_sub_8_33_g586(out2[22] ,dec_sub_8_33_n_123 ,n_24);
  xnor dec_sub_8_33_g587(out2[14] ,dec_sub_8_33_n_106 ,dec_sub_8_33_n_61);
  nor dec_sub_8_33_g588(dec_sub_8_33_n_3 ,dec_sub_8_33_n_59 ,dec_sub_8_33_n_93);
  xnor dec_sub_8_33_g589(out2[4] ,dec_sub_8_33_n_85 ,dec_sub_8_33_n_55);
  xnor dec_sub_8_33_g590(out2[24] ,dec_sub_8_33_n_133 ,dec_sub_8_33_n_53);
  xor dec_sub_8_33_g591(out2[26] ,dec_sub_8_33_n_135 ,dec_sub_8_33_n_58);
  xnor inc_add_7_33_g381(out1[31] ,inc_add_7_33_n_147 ,n_33);
  or inc_add_7_33_g383(inc_add_7_33_n_147 ,inc_add_7_33_n_58 ,inc_add_7_33_n_146);
  or inc_add_7_33_g385(inc_add_7_33_n_146 ,inc_add_7_33_n_51 ,inc_add_7_33_n_145);
  or inc_add_7_33_g387(inc_add_7_33_n_145 ,inc_add_7_33_n_52 ,inc_add_7_33_n_144);
  or inc_add_7_33_g389(inc_add_7_33_n_144 ,inc_add_7_33_n_46 ,inc_add_7_33_n_140);
  and inc_add_7_33_g390(out1[26] ,inc_add_7_33_n_141 ,inc_add_7_33_n_140);
  xnor inc_add_7_33_g391(out1[25] ,inc_add_7_33_n_139 ,inc_add_7_33_n_22);
  or inc_add_7_33_g392(inc_add_7_33_n_141 ,inc_add_7_33_n_20 ,inc_add_7_33_n_137);
  or inc_add_7_33_g393(inc_add_7_33_n_140 ,inc_add_7_33_n_53 ,inc_add_7_33_n_138);
  or inc_add_7_33_g395(inc_add_7_33_n_139 ,inc_add_7_33_n_66 ,inc_add_7_33_n_135);
  not inc_add_7_33_g396(inc_add_7_33_n_138 ,inc_add_7_33_n_137);
  and inc_add_7_33_g397(inc_add_7_33_n_137 ,inc_add_7_33_n_76 ,inc_add_7_33_n_134);
  xnor inc_add_7_33_g398(out1[23] ,inc_add_7_33_n_131 ,n_25);
  not inc_add_7_33_g399(inc_add_7_33_n_135 ,inc_add_7_33_n_134);
  and inc_add_7_33_g400(inc_add_7_33_n_134 ,n_25 ,inc_add_7_33_n_132);
  nor inc_add_7_33_g401(inc_add_7_33_n_133 ,inc_add_7_33_n_132 ,inc_add_7_33_n_130);
  not inc_add_7_33_g404(inc_add_7_33_n_132 ,inc_add_7_33_n_131);
  or inc_add_7_33_g405(inc_add_7_33_n_131 ,inc_add_7_33_n_71 ,inc_add_7_33_n_127);
  and inc_add_7_33_g406(inc_add_7_33_n_130 ,inc_add_7_33_n_71 ,inc_add_7_33_n_127);
  xor inc_add_7_33_g407(out1[20] ,inc_add_7_33_n_119 ,inc_add_7_33_n_36);
  xor inc_add_7_33_g408(out1[18] ,inc_add_7_33_n_121 ,inc_add_7_33_n_40);
  or inc_add_7_33_g410(inc_add_7_33_n_127 ,inc_add_7_33_n_82 ,inc_add_7_33_n_120);
  or inc_add_7_33_g411(inc_add_7_33_n_126 ,inc_add_7_33_n_69 ,inc_add_7_33_n_120);
  or inc_add_7_33_g412(inc_add_7_33_n_125 ,inc_add_7_33_n_65 ,inc_add_7_33_n_122);
  xnor inc_add_7_33_g413(out1[16] ,inc_add_7_33_n_117 ,inc_add_7_33_n_30);
  or inc_add_7_33_g414(inc_add_7_33_n_123 ,inc_add_7_33_n_68 ,inc_add_7_33_n_117);
  not inc_add_7_33_g415(inc_add_7_33_n_122 ,inc_add_7_33_n_121);
  and inc_add_7_33_g416(inc_add_7_33_n_121 ,inc_add_7_33_n_78 ,inc_add_7_33_n_116);
  not inc_add_7_33_g417(inc_add_7_33_n_120 ,inc_add_7_33_n_119);
  and inc_add_7_33_g418(inc_add_7_33_n_119 ,inc_add_7_33_n_91 ,inc_add_7_33_n_116);
  xnor inc_add_7_33_g419(out1[15] ,inc_add_7_33_n_113 ,n_17);
  not inc_add_7_33_g420(inc_add_7_33_n_116 ,inc_add_7_33_n_117);
  or inc_add_7_33_g421(inc_add_7_33_n_117 ,inc_add_7_33_n_59 ,inc_add_7_33_n_114);
  xnor inc_add_7_33_g422(out1[14] ,inc_add_7_33_n_110 ,inc_add_7_33_n_26);
  or inc_add_7_33_g425(inc_add_7_33_n_114 ,inc_add_7_33_n_64 ,inc_add_7_33_n_110);
  or inc_add_7_33_g426(inc_add_7_33_n_113 ,inc_add_7_33_n_59 ,inc_add_7_33_n_110);
  xor inc_add_7_33_g427(out1[12] ,inc_add_7_33_n_104 ,inc_add_7_33_n_34);
  xor inc_add_7_33_g428(out1[10] ,inc_add_7_33_n_102 ,inc_add_7_33_n_38);
  or inc_add_7_33_g430(inc_add_7_33_n_110 ,inc_add_7_33_n_81 ,inc_add_7_33_n_105);
  or inc_add_7_33_g431(inc_add_7_33_n_109 ,inc_add_7_33_n_67 ,inc_add_7_33_n_105);
  or inc_add_7_33_g432(inc_add_7_33_n_108 ,inc_add_7_33_n_60 ,inc_add_7_33_n_103);
  xnor inc_add_7_33_g433(out1[8] ,inc_add_7_33_n_101 ,inc_add_7_33_n_32);
  or inc_add_7_33_g434(inc_add_7_33_n_106 ,inc_add_7_33_n_63 ,inc_add_7_33_n_101);
  not inc_add_7_33_g435(inc_add_7_33_n_105 ,inc_add_7_33_n_104);
  and inc_add_7_33_g436(inc_add_7_33_n_104 ,inc_add_7_33_n_92 ,inc_add_7_33_n_100);
  not inc_add_7_33_g437(inc_add_7_33_n_103 ,inc_add_7_33_n_102);
  and inc_add_7_33_g438(inc_add_7_33_n_102 ,inc_add_7_33_n_80 ,inc_add_7_33_n_100);
  not inc_add_7_33_g440(inc_add_7_33_n_100 ,inc_add_7_33_n_101);
  or inc_add_7_33_g441(inc_add_7_33_n_101 ,inc_add_7_33_n_16 ,inc_add_7_33_n_96);
  xnor inc_add_7_33_g442(out1[6] ,inc_add_7_33_n_93 ,inc_add_7_33_n_62);
  xnor inc_add_7_33_g443(out1[5] ,inc_add_7_33_n_95 ,inc_add_7_33_n_19);
  or inc_add_7_33_g444(inc_add_7_33_n_97 ,inc_add_7_33_n_16 ,inc_add_7_33_n_94);
  or inc_add_7_33_g445(inc_add_7_33_n_96 ,inc_add_7_33_n_56 ,inc_add_7_33_n_94);
  or inc_add_7_33_g447(inc_add_7_33_n_95 ,inc_add_7_33_n_70 ,inc_add_7_33_n_90);
  not inc_add_7_33_g448(inc_add_7_33_n_94 ,inc_add_7_33_n_93);
  and inc_add_7_33_g449(inc_add_7_33_n_93 ,inc_add_7_33_n_75 ,inc_add_7_33_n_89);
  nor inc_add_7_33_g451(inc_add_7_33_n_92 ,inc_add_7_33_n_60 ,inc_add_7_33_n_87);
  nor inc_add_7_33_g452(inc_add_7_33_n_91 ,inc_add_7_33_n_65 ,inc_add_7_33_n_86);
  not inc_add_7_33_g453(inc_add_7_33_n_89 ,inc_add_7_33_n_90);
  or inc_add_7_33_g454(inc_add_7_33_n_90 ,inc_add_7_33_n_48 ,inc_add_7_33_n_84);
  xnor inc_add_7_33_g455(out1[2] ,inc_add_7_33_n_28 ,inc_add_7_33_n_24);
  or inc_add_7_33_g456(inc_add_7_33_n_87 ,inc_add_7_33_n_50 ,inc_add_7_33_n_79);
  or inc_add_7_33_g457(inc_add_7_33_n_86 ,inc_add_7_33_n_45 ,inc_add_7_33_n_77);
  or inc_add_7_33_g458(inc_add_7_33_n_85 ,inc_add_7_33_n_61 ,inc_add_7_33_n_28);
  or inc_add_7_33_g459(inc_add_7_33_n_84 ,inc_add_7_33_n_61 ,inc_add_7_33_n_73);
  and inc_add_7_33_g460(out1[1] ,inc_add_7_33_n_73 ,inc_add_7_33_n_74);
  or inc_add_7_33_g461(inc_add_7_33_n_82 ,inc_add_7_33_n_47 ,inc_add_7_33_n_69);
  or inc_add_7_33_g462(inc_add_7_33_n_81 ,inc_add_7_33_n_54 ,inc_add_7_33_n_67);
  not inc_add_7_33_g463(inc_add_7_33_n_80 ,inc_add_7_33_n_79);
  or inc_add_7_33_g464(inc_add_7_33_n_79 ,inc_add_7_33_n_49 ,inc_add_7_33_n_63);
  not inc_add_7_33_g465(inc_add_7_33_n_78 ,inc_add_7_33_n_77);
  or inc_add_7_33_g466(inc_add_7_33_n_77 ,inc_add_7_33_n_55 ,inc_add_7_33_n_68);
  and inc_add_7_33_g467(inc_add_7_33_n_76 ,inc_add_7_33_n_22 ,inc_add_7_33_n_42);
  and inc_add_7_33_g468(inc_add_7_33_n_75 ,inc_add_7_33_n_19 ,inc_add_7_33_n_44);
  or inc_add_7_33_g469(inc_add_7_33_n_74 ,n_3 ,inc_add_7_33_n_17);
  or inc_add_7_33_g470(inc_add_7_33_n_73 ,inc_add_7_33_n_72 ,inc_add_7_33_n_57);
  not inc_add_7_33_g471(inc_add_7_33_n_72 ,n_3);
  not inc_add_7_33_g472(inc_add_7_33_n_71 ,n_24);
  not inc_add_7_33_g477(inc_add_7_33_n_70 ,inc_add_7_33_n_44);
  not inc_add_7_33_g478(inc_add_7_33_n_69 ,inc_add_7_33_n_36);
  not inc_add_7_33_g479(inc_add_7_33_n_68 ,inc_add_7_33_n_30);
  not inc_add_7_33_g480(inc_add_7_33_n_67 ,inc_add_7_33_n_34);
  not inc_add_7_33_g481(inc_add_7_33_n_66 ,inc_add_7_33_n_42);
  not inc_add_7_33_g482(inc_add_7_33_n_65 ,inc_add_7_33_n_40);
  not inc_add_7_33_g487(inc_add_7_33_n_64 ,n_17);
  not inc_add_7_33_g491(inc_add_7_33_n_63 ,inc_add_7_33_n_32);
  not inc_add_7_33_g492(inc_add_7_33_n_62 ,n_8);
  not inc_add_7_33_g493(inc_add_7_33_n_61 ,inc_add_7_33_n_24);
  not inc_add_7_33_g494(inc_add_7_33_n_60 ,inc_add_7_33_n_38);
  not inc_add_7_33_g496(inc_add_7_33_n_59 ,inc_add_7_33_n_26);
  not inc_add_7_33_drc_bufs(inc_add_7_33_n_44 ,inc_add_7_33_n_43);
  not inc_add_7_33_drc_bufs500(inc_add_7_33_n_43 ,n_6);
  not inc_add_7_33_drc_bufs502(inc_add_7_33_n_42 ,inc_add_7_33_n_41);
  not inc_add_7_33_drc_bufs504(inc_add_7_33_n_41 ,n_26);
  not inc_add_7_33_drc_bufs506(inc_add_7_33_n_40 ,inc_add_7_33_n_39);
  not inc_add_7_33_drc_bufs508(inc_add_7_33_n_39 ,n_20);
  not inc_add_7_33_drc_bufs510(inc_add_7_33_n_38 ,inc_add_7_33_n_37);
  not inc_add_7_33_drc_bufs512(inc_add_7_33_n_37 ,n_12);
  not inc_add_7_33_drc_bufs514(inc_add_7_33_n_36 ,inc_add_7_33_n_35);
  not inc_add_7_33_drc_bufs516(inc_add_7_33_n_35 ,n_22);
  not inc_add_7_33_drc_bufs518(inc_add_7_33_n_34 ,inc_add_7_33_n_33);
  not inc_add_7_33_drc_bufs520(inc_add_7_33_n_33 ,n_14);
  not inc_add_7_33_drc_bufs522(inc_add_7_33_n_32 ,inc_add_7_33_n_31);
  not inc_add_7_33_drc_bufs524(inc_add_7_33_n_31 ,n_10);
  not inc_add_7_33_drc_bufs526(inc_add_7_33_n_30 ,inc_add_7_33_n_29);
  not inc_add_7_33_drc_bufs528(inc_add_7_33_n_29 ,n_18);
  not inc_add_7_33_drc_bufs531(inc_add_7_33_n_28 ,inc_add_7_33_n_27);
  not inc_add_7_33_drc_bufs532(inc_add_7_33_n_27 ,inc_add_7_33_n_73);
  not inc_add_7_33_drc_bufs536(inc_add_7_33_n_47 ,n_23);
  not inc_add_7_33_drc_bufs540(inc_add_7_33_n_54 ,n_15);
  not inc_add_7_33_drc_bufs544(inc_add_7_33_n_58 ,n_32);
  not inc_add_7_33_drc_bufs546(inc_add_7_33_n_26 ,inc_add_7_33_n_25);
  not inc_add_7_33_drc_bufs548(inc_add_7_33_n_25 ,n_16);
  not inc_add_7_33_drc_bufs550(inc_add_7_33_n_24 ,inc_add_7_33_n_23);
  not inc_add_7_33_drc_bufs552(inc_add_7_33_n_23 ,n_4);
  not inc_add_7_33_drc_bufs556(inc_add_7_33_n_45 ,n_21);
  not inc_add_7_33_drc_bufs560(inc_add_7_33_n_49 ,n_11);
  not inc_add_7_33_drc_bufs564(inc_add_7_33_n_50 ,n_13);
  not inc_add_7_33_drc_bufs568(inc_add_7_33_n_52 ,n_30);
  not inc_add_7_33_drc_bufs572(inc_add_7_33_n_55 ,n_19);
  not inc_add_7_33_drc_bufs574(inc_add_7_33_n_22 ,inc_add_7_33_n_21);
  not inc_add_7_33_drc_bufs576(inc_add_7_33_n_21 ,n_27);
  not inc_add_7_33_drc_bufs580(inc_add_7_33_n_48 ,n_5);
  not inc_add_7_33_drc_bufs584(inc_add_7_33_n_56 ,n_9);
  not inc_add_7_33_drc_bufs588(inc_add_7_33_n_51 ,n_31);
  not inc_add_7_33_drc_bufs591(inc_add_7_33_n_20 ,inc_add_7_33_n_53);
  not inc_add_7_33_drc_bufs592(inc_add_7_33_n_53 ,n_28);
  not inc_add_7_33_drc_bufs596(inc_add_7_33_n_46 ,n_29);
  not inc_add_7_33_drc_bufs598(inc_add_7_33_n_19 ,inc_add_7_33_n_18);
  not inc_add_7_33_drc_bufs600(inc_add_7_33_n_18 ,n_7);
  not inc_add_7_33_drc_bufs603(inc_add_7_33_n_17 ,inc_add_7_33_n_57);
  not inc_add_7_33_drc_bufs604(inc_add_7_33_n_57 ,n_2);
  not inc_add_7_33_drc_bufs607(inc_add_7_33_n_16 ,inc_add_7_33_n_15);
  not inc_add_7_33_drc_bufs608(inc_add_7_33_n_15 ,inc_add_7_33_n_62);
  buf inc_add_7_33_drc_bufs610(out1[22] ,inc_add_7_33_n_133);
  xor inc_add_7_33_g2(out1[4] ,inc_add_7_33_n_90 ,inc_add_7_33_n_43);
  xor inc_add_7_33_g621(out1[24] ,inc_add_7_33_n_135 ,inc_add_7_33_n_41);
  xor inc_add_7_33_g622(out1[21] ,inc_add_7_33_n_126 ,inc_add_7_33_n_47);
  xor inc_add_7_33_g623(out1[13] ,inc_add_7_33_n_109 ,inc_add_7_33_n_54);
  xor inc_add_7_33_g624(out1[30] ,inc_add_7_33_n_146 ,inc_add_7_33_n_58);
  xor inc_add_7_33_g625(out1[19] ,inc_add_7_33_n_125 ,inc_add_7_33_n_45);
  xor inc_add_7_33_g626(out1[9] ,inc_add_7_33_n_106 ,inc_add_7_33_n_49);
  xor inc_add_7_33_g627(out1[11] ,inc_add_7_33_n_108 ,inc_add_7_33_n_50);
  xor inc_add_7_33_g628(out1[28] ,inc_add_7_33_n_144 ,inc_add_7_33_n_52);
  xor inc_add_7_33_g629(out1[17] ,inc_add_7_33_n_123 ,inc_add_7_33_n_55);
  xor inc_add_7_33_g630(out1[3] ,inc_add_7_33_n_85 ,inc_add_7_33_n_48);
  xor inc_add_7_33_g631(out1[7] ,inc_add_7_33_n_97 ,inc_add_7_33_n_56);
  xor inc_add_7_33_g632(out1[29] ,inc_add_7_33_n_145 ,inc_add_7_33_n_51);
  xor inc_add_7_33_g633(out1[27] ,inc_add_7_33_n_140 ,inc_add_7_33_n_46);
  buf g8418(csa_tree_add_7_27_groupi_n_895 ,csa_tree_add_7_27_groupi_n_790);
endmodule
