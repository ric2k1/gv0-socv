module top( n7 , n9 , n12 , n18 , n19 , n33 , n38 , n39 , n56 , n60 , n61 , n64 , n66 , n67 , n75 , n77 , n83 , n84 , n92 , n101 , n107 , n112 , n117 , n119 , n123 , n128 , n129 , n130 , n132 , n157 , n158 , n165 , n168 , n173 , n179 , n186 , n187 , n190 , n193 , n211 , n222 , n228 , n235 , n236 , n238 , n239 , n245 , n249 , n257 , n259 , n261 , n262 , n264 , n270 , n288 , n297 , n307 , n315 , n319 , n320 , n321 , n326 , n335 , n337 , n342 , n357 , n361 , n370 , n371 , n375 , n377 , n378 , n379 , n380 , n381 , n384 , n386 , n387 , n389 , n403 , n413 , n417 , n448 , n454 , n456 , n457 , n476 , n482 , n487 , n488 , n495 , n504 , n516 , n520 , n530 , n541 , n542 , n544 , n547 , n560 , n564 , n565 , n566 , n567 , n574 , n579 , n591 , n596 , n600 , n601 , n606 , n611 , n617 , n623 , n627 , n635 , n636 , n643 , n649 , n661 , n668 , n673 , n676 , n697 , n708 , n714 , n715 , n721 , n722 , n754 , n758 , n760 , n765 , n776 , n779 , n786 , n793 , n801 , n807 , n813 , n824 , n830 , n840 , n841 , n845 , n849 , n850 , n860 , n878 , n882 , n887 , n889 , n894 , n912 , n917 , n918 , n937 , n944 , n946 , n951 , n955 , n961 , n962 , n964 , n966 , n967 , n971 , n974 , n984 , n999 , n1016 , n1027 , n1033 , n1039 , n1043 , n1044 , n1047 , n1050 , n1058 , n1065 , n1087 , n1088 , n1095 , n1096 , n1097 , n1100 , n1110 , n1119 , n1125 , n1135 , n1140 , n1150 , n1163 , n1172 , n1175 , n1177 , n1180 , n1181 , n1182 , n1186 , n1205 , n1207 , n1219 , n1224 , n1227 , n1233 , n1238 , n1269 , n1270 , n1279 , n1281 , n1288 , n1297 , n1299 , n1314 , n1322 , n1338 , n1346 , n1353 , n1355 , n1357 , n1361 , n1362 , n1363 , n1366 , n1370 , n1377 , n1378 , n1390 , n1391 , n1396 , n1402 , n1406 , n1408 , n1409 , n1414 , n1425 , n1426 , n1427 , n1435 , n1436 , n1454 , n1462 , n1463 , n1464 , n1471 , n1485 , n1491 , n1495 , n1498 , n1503 , n1510 , n1511 , n1515 , n1518 , n1519 , n1534 , n1540 , n1543 , n1553 , n1568 , n1575 , n1584 , n1587 , n1598 , n1613 , n1631 , n1632 , n1633 , n1649 , n1654 , n1655 , n1657 , n1660 , n1663 , n1674 , n1675 , n1676 , n1682 , n1697 , n1698 , n1700 , n1707 , n1708 , n1710 , n1721 , n1729 , n1733 , n1740 , n1743 , n1753 , n1755 , n1756 , n1761 , n1768 , n1780 , n1784 , n1788 , n1790 , n1793 , n1794 );
    input n7 , n9 , n12 , n19 , n33 , n38 , n39 , n60 , n64 , n77 , n84 , n92 , n119 , n128 , n132 , n157 , n179 , n186 , n187 , n190 , n228 , n236 , n238 , n239 , n257 , n261 , n270 , n288 , n297 , n307 , n319 , n321 , n326 , n335 , n342 , n371 , n377 , n378 , n380 , n384 , n386 , n387 , n389 , n403 , n448 , n457 , n482 , n488 , n495 , n504 , n516 , n520 , n530 , n541 , n544 , n560 , n564 , n565 , n566 , n579 , n591 , n600 , n601 , n606 , n617 , n627 , n636 , n643 , n668 , n676 , n697 , n708 , n714 , n715 , n721 , n754 , n758 , n760 , n779 , n801 , n807 , n813 , n830 , n841 , n850 , n887 , n894 , n912 , n917 , n918 , n937 , n946 , n955 , n961 , n962 , n966 , n971 , n984 , n999 , n1016 , n1033 , n1039 , n1043 , n1058 , n1088 , n1095 , n1097 , n1100 , n1119 , n1125 , n1135 , n1150 , n1172 , n1175 , n1177 , n1180 , n1181 , n1182 , n1205 , n1207 , n1219 , n1227 , n1238 , n1279 , n1281 , n1288 , n1299 , n1338 , n1353 , n1357 , n1361 , n1362 , n1363 , n1366 , n1391 , n1396 , n1402 , n1406 , n1408 , n1426 , n1427 , n1435 , n1436 , n1454 , n1463 , n1471 , n1485 , n1498 , n1503 , n1515 , n1518 , n1519 , n1534 , n1540 , n1553 , n1568 , n1575 , n1598 , n1613 , n1632 , n1633 , n1649 , n1655 , n1660 , n1663 , n1674 , n1675 , n1700 , n1707 , n1729 , n1740 , n1743 , n1753 , n1755 , n1756 , n1768 , n1788 , n1790 ;
    output n18 , n56 , n61 , n66 , n67 , n75 , n83 , n101 , n107 , n112 , n117 , n123 , n129 , n130 , n158 , n165 , n168 , n173 , n193 , n211 , n222 , n235 , n245 , n249 , n259 , n262 , n264 , n315 , n320 , n337 , n357 , n361 , n370 , n375 , n379 , n381 , n413 , n417 , n454 , n456 , n476 , n487 , n542 , n547 , n567 , n574 , n596 , n611 , n623 , n635 , n649 , n661 , n673 , n722 , n765 , n776 , n786 , n793 , n824 , n840 , n845 , n849 , n860 , n878 , n882 , n889 , n944 , n951 , n964 , n967 , n974 , n1027 , n1044 , n1047 , n1050 , n1065 , n1087 , n1096 , n1110 , n1140 , n1163 , n1186 , n1224 , n1233 , n1269 , n1270 , n1297 , n1314 , n1322 , n1346 , n1355 , n1370 , n1377 , n1378 , n1390 , n1409 , n1414 , n1425 , n1462 , n1464 , n1491 , n1495 , n1510 , n1511 , n1543 , n1584 , n1587 , n1631 , n1654 , n1657 , n1676 , n1682 , n1697 , n1698 , n1708 , n1710 , n1721 , n1733 , n1761 , n1780 , n1784 , n1793 , n1794 ;
    wire n0 , n1 , n2 , n3 , n4 , n5 , n6 , n8 , n10 , n11 , n13 , n14 , n15 , n16 , n17 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n34 , n35 , n36 , n37 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n57 , n58 , n59 , n62 , n63 , n65 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n76 , n78 , n79 , n80 , n81 , n82 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n102 , n103 , n104 , n105 , n106 , n108 , n109 , n110 , n111 , n113 , n114 , n115 , n116 , n118 , n120 , n121 , n122 , n124 , n125 , n126 , n127 , n131 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n159 , n160 , n161 , n162 , n163 , n164 , n166 , n167 , n169 , n170 , n171 , n172 , n174 , n175 , n176 , n177 , n178 , n180 , n181 , n182 , n183 , n184 , n185 , n188 , n189 , n191 , n192 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n223 , n224 , n225 , n226 , n227 , n229 , n230 , n231 , n232 , n233 , n234 , n237 , n240 , n241 , n242 , n243 , n244 , n246 , n247 , n248 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n258 , n260 , n263 , n265 , n266 , n267 , n268 , n269 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n316 , n317 , n318 , n322 , n323 , n324 , n325 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n336 , n338 , n339 , n340 , n341 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n358 , n359 , n360 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n372 , n373 , n374 , n376 , n382 , n383 , n385 , n388 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n414 , n415 , n416 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n449 , n450 , n451 , n452 , n453 , n455 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n477 , n478 , n479 , n480 , n481 , n483 , n484 , n485 , n486 , n489 , n490 , n491 , n492 , n493 , n494 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n517 , n518 , n519 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n543 , n545 , n546 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n561 , n562 , n563 , n568 , n569 , n570 , n571 , n572 , n573 , n575 , n576 , n577 , n578 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n592 , n593 , n594 , n595 , n597 , n598 , n599 , n602 , n603 , n604 , n605 , n607 , n608 , n609 , n610 , n612 , n613 , n614 , n615 , n616 , n618 , n619 , n620 , n621 , n622 , n624 , n625 , n626 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n637 , n638 , n639 , n640 , n641 , n642 , n644 , n645 , n646 , n647 , n648 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n662 , n663 , n664 , n665 , n666 , n667 , n669 , n670 , n671 , n672 , n674 , n675 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n709 , n710 , n711 , n712 , n713 , n716 , n717 , n718 , n719 , n720 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n755 , n756 , n757 , n759 , n761 , n762 , n763 , n764 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n777 , n778 , n780 , n781 , n782 , n783 , n784 , n785 , n787 , n788 , n789 , n790 , n791 , n792 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n802 , n803 , n804 , n805 , n806 , n808 , n809 , n810 , n811 , n812 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n825 , n826 , n827 , n828 , n829 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n842 , n843 , n844 , n846 , n847 , n848 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n879 , n880 , n881 , n883 , n884 , n885 , n886 , n888 , n890 , n891 , n892 , n893 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n913 , n914 , n915 , n916 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n938 , n939 , n940 , n941 , n942 , n943 , n945 , n947 , n948 , n949 , n950 , n952 , n953 , n954 , n956 , n957 , n958 , n959 , n960 , n963 , n965 , n968 , n969 , n970 , n972 , n973 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1028 , n1029 , n1030 , n1031 , n1032 , n1034 , n1035 , n1036 , n1037 , n1038 , n1040 , n1041 , n1042 , n1045 , n1046 , n1048 , n1049 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1098 , n1099 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1120 , n1121 , n1122 , n1123 , n1124 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1136 , n1137 , n1138 , n1139 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1173 , n1174 , n1176 , n1178 , n1179 , n1183 , n1184 , n1185 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1206 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1220 , n1221 , n1222 , n1223 , n1225 , n1226 , n1228 , n1229 , n1230 , n1231 , n1232 , n1234 , n1235 , n1236 , n1237 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1280 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1298 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1354 , n1356 , n1358 , n1359 , n1360 , n1364 , n1365 , n1367 , n1368 , n1369 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1392 , n1393 , n1394 , n1395 , n1397 , n1398 , n1399 , n1400 , n1401 , n1403 , n1404 , n1405 , n1407 , n1410 , n1411 , n1412 , n1413 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1486 , n1487 , n1488 , n1489 , n1490 , n1492 , n1493 , n1494 , n1496 , n1497 , n1499 , n1500 , n1501 , n1502 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1512 , n1513 , n1514 , n1516 , n1517 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1535 , n1536 , n1537 , n1538 , n1539 , n1541 , n1542 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1585 , n1586 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1650 , n1651 , n1652 , n1653 , n1656 , n1658 , n1659 , n1661 , n1662 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1677 , n1678 , n1679 , n1680 , n1681 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1699 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1709 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1730 , n1731 , n1732 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1741 , n1742 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1754 , n1757 , n1758 , n1759 , n1760 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1781 , n1782 , n1783 , n1785 , n1786 , n1787 , n1789 , n1791 , n1792 , n1795 , n1796 , n1797 ;
assign n1319 = ~(n228 | n95);
assign n996 = ~n1457;
assign n337 = ~(n220 | n140);
assign n1099 = ~(n539 | n1022);
assign n464 = n24 | n465;
assign n1648 = n1081 | n1694;
assign n507 = n616 | n68;
assign n1741 = ~(n1718 ^ n1332);
assign n586 = n1103 & n81;
assign n1600 = ~(n1618 | n807);
assign n1442 = n1439 | n1316;
assign n1011 = n186 | n1027;
assign n1782 = n1690 | n1694;
assign n1306 = n723 & n1251;
assign n491 = ~n1397;
assign n1677 = ~(n525 ^ n578);
assign n1034 = n588 | n1497;
assign n1603 = n627 | n964;
assign n1090 = n1146 | n1407;
assign n237 = ~(n261 | n1028);
assign n562 = n842 & n356;
assign n840 = n452 | n421;
assign n218 = n1668 & n590;
assign n1040 = ~(n1395 | n354);
assign n24 = ~(n44 | n282);
assign n890 = n579 | n150;
assign n1171 = n99 & n1531;
assign n670 = ~(n1435 ^ n1043);
assign n1237 = ~(n1788 | n1457);
assign n551 = n579 | n1189;
assign n1469 = n186 | n75;
assign n932 = ~(n261 | n281);
assign n1221 = ~(n378 | n1268);
assign n1548 = n186 | n370;
assign n399 = n1326;
assign n674 = ~(n261 | n1746);
assign n1003 = ~n903;
assign n1720 = ~n240;
assign n48 = n669 | n77;
assign n1533 = n307 | n964;
assign n63 = n1391 & n713;
assign n1110 = n215 & n1764;
assign n1679 = ~(n473 | n1480);
assign n166 = ~(n1660 | n714);
assign n1480 = n1301 | n214;
assign n1616 = ~(n378 | n324);
assign n1597 = ~n884;
assign n436 = ~(n1765 | n219);
assign n503 = ~(n193 | n1662);
assign n1433 = ~n1039;
assign n557 = ~(n1619 ^ n1555);
assign n1048 = ~(n550 ^ n685);
assign n1035 = ~(n778 ^ n1294);
assign n1766 = ~n1545;
assign n1697 = n1414;
assign n1550 = ~n1085;
assign n1614 = ~(n1281 | n339);
assign n1023 = ~(n188 | n807);
assign n561 = ~n1506;
assign n862 = n909;
assign n1046 = n1235 & n1636;
assign n1528 = n1295 | n947;
assign n518 = n302 & n1244;
assign n1437 = n396 & n55;
assign n1179 = ~(n44 | n881);
assign n1722 = n186 | n1314;
assign n891 = n627 | n1110;
assign n428 = ~n538;
assign n1318 = n307 | n1710;
assign n134 = ~n1172;
assign n1290 = n213 | n613;
assign n1750 = ~n1437;
assign n1452 = ~(n44 | n1563);
assign n1355 = n288;
assign n700 = n307 | n905;
assign n67 = ~(n402 | n544);
assign n397 = n1106 | n1257;
assign n137 = n1205 | n964;
assign n1458 = ~(n377 | n701);
assign n175 = n764 | n1200;
assign n1060 = n462 | n1694;
assign n202 = ~(n669 | n504);
assign n1693 = n1205 | n1027;
assign n838 = n1072 | n1694;
assign n770 = ~(n862 | n355);
assign n160 = ~(n560 | n1018);
assign n242 = n139 & n436;
assign n286 = n1147 | n1749;
assign n232 = ~(n200 | n288);
assign n1761 = n1684 | n762;
assign n133 = ~(n1172 | n1519);
assign n944 = ~(n220 | n70);
assign n1460 = n1146 | n698;
assign n1667 = ~(n579 | n647);
assign n95 = n1205 | n168;
assign n1520 = ~(n1241 | n1585);
assign n1692 = n1113 | n998;
assign n1438 = n990 | n1200;
assign n1158 = ~(n704 | n144);
assign n251 = ~(n1681 | n479);
assign n805 = n1205 | n370;
assign n476 = n1613 & n1716;
assign n746 = ~(n560 | n1011);
assign n1051 = ~(n428 ^ n916);
assign n1670 = ~(n560 | n1380);
assign n1627 = ~(n94 | n1215);
assign n845 = n1613;
assign n208 = ~(n946 | n714);
assign n469 = n73 & n575;
assign n369 = n579 | n562;
assign n628 = n2 & n1204;
assign n1772 = n1744 | n229;
assign n266 = ~(n654 ^ n1741);
assign n1285 = n694 | n227;
assign n1012 = n1295 | n1793;
assign n595 = n186 | n487;
assign n950 = n1295 | n1010;
assign n1508 = n651 | n942;
assign n1785 = ~n1598;
assign n1669 = ~(n412 ^ n1108);
assign n759 = ~(n1580 | n1330);
assign n366 = ~(n853 | n1118);
assign n826 = n1280 | n394;
assign n1304 = n398 | n1694;
assign n735 = n1792 | n628;
assign n191 = n1585 & n1545;
assign n429 = ~(n378 | n1111);
assign n91 = n780 | n1440;
assign n1403 = ~(n1166 | n319);
assign n907 = ~n89;
assign n505 = n1349 | n1562;
assign n1145 = n63 | n176;
assign n1291 = ~(n1755 | n343);
assign n828 = n1660 & n1288;
assign n23 = ~n286;
assign n110 = ~(n1335 | n797);
assign n1676 = ~n1338;
assign n1297 = n203 | n349;
assign n842 = n298 | n1190;
assign n880 = ~n1226;
assign n741 = n147 & n1626;
assign n435 = n749 | n585;
assign n75 = n1453 & n241;
assign n1604 = n1235 & n252;
assign n1428 = n1374 | n1524;
assign n1546 = n1295 | n1422;
assign n1260 = n627 | n168;
assign n1410 = n206 | n879;
assign n361 = n1116 | n1692;
assign n1541 = ~(n377 | n1714);
assign n1341 = n1473 | n1211;
assign n345 = ~n1391;
assign n774 = ~n1663;
assign n215 = n1146 | n156;
assign n1369 = n703 & n243;
assign n669 = ~n617;
assign n130 = n1523 | n770;
assign n1647 = ~(n517 ^ n1445);
assign n1691 = ~(n579 | n1145);
assign n1282 = n1298 | n579;
assign n666 = ~(n526 ^ n1217);
assign n888 = n774 | n1694;
assign n856 = ~(n1032 | n1129);
assign n1244 = n777 & n185;
assign n259 = n732 & n858;
assign n1696 = ~n147;
assign n211 = n1602 | n605;
assign n1292 = n1618 | n1312;
assign n1066 = n1205 | n259;
assign n121 = n1384 | n1571;
assign n656 = n1482 | n480;
assign n1615 = ~n1097;
assign n1252 = n1054 | n268;
assign n1496 = n307 | n1346;
assign n388 = ~(n560 | n310);
assign n1524 = n348 | n283;
assign n1622 = ~(n1681 | n1363);
assign n698 = n1488 | n579;
assign n85 = n1419 | n1694;
assign n373 = n1037 & n65;
assign n223 = n982 | n1561;
assign n1287 = ~(n44 | n877);
assign n1007 = ~(n380 | n1227);
assign n784 = n271 | n1512;
assign n1412 = n857 | n809;
assign n332 = ~n758;
assign n168 = n74 & n712;
assign n347 = ~(n472 | n591);
assign n437 = ~n12;
assign n936 = ~n1171;
assign n143 = ~(n1162 | n1572);
assign n647 = ~(n353 | n1003);
assign n1681 = ~n1281;
assign n1431 = ~(n1600 | n1748);
assign n1509 = n1146 | n1282;
assign n975 = n338 | n1234;
assign n184 = n828 | n1398;
assign n1141 = ~(n545 | n1309);
assign n974 = n709 | n1290;
assign n1202 = ~(n832 | n708);
assign n1167 = n435 | n91;
assign n585 = n495 & n426;
assign n461 = n992 | n22;
assign n1744 = ~(n1162 | n908);
assign n1283 = ~(n1249 ^ n1);
assign n1185 = n344 | n695;
assign n330 = ~(n1713 | n807);
assign n57 = n1146 & n1400;
assign n519 = n1295 | n1779;
assign n1661 = ~n1047;
assign n512 = ~(n228 | n1187);
assign n443 = ~(n1281 | n254);
assign n494 = n1125 & n76;
assign n90 = ~(n1162 | n874);
assign n295 = n1135 & n407;
assign n539 = ~n560;
assign n1206 = ~(n261 | n1494);
assign n1745 = ~(n261 | n1758);
assign n317 = n1536 | n276;
assign n1731 = ~(n1591 | n1642);
assign n691 = n1295 | n960;
assign n183 = n1670 | n533;
assign n49 = n675 | n1146;
assign n230 = n1375 | n1200;
assign n1718 = n930 | n232;
assign n82 = n1417 | n579;
assign n1429 = ~n708;
assign n1711 = ~(n1755 | n592);
assign n398 = ~n606;
assign n432 = n1334 | n1694;
assign n1087 = n1460 & n292;
assign n1184 = ~(n378 | n608);
assign n1333 = n1429 | n614;
assign n1415 = ~(n438 ^ n825);
assign n1041 = ~n482;
assign n1724 = ~(n378 | n113);
assign n956 = ~n1279;
assign n277 = ~(n560 | n305);
assign n1147 = ~n1406;
assign n930 = ~(n710 | n614);
assign n903 = ~(n1093 ^ n1329);
assign n572 = ~(n966 | n1227);
assign n1257 = n396 & n1795;
assign n61 = ~n1503;
assign n511 = ~(n560 | n1424);
assign n1188 = n1105 | n1043;
assign n1642 = ~n278;
assign n1254 = ~(n378 | n1603);
assign n1153 = ~(n832 | n1043);
assign n1763 = ~(n438 | n1569);
assign n768 = n821 | n268;
assign n1082 = ~(n579 | n1672);
assign n699 = n442 | n1589;
assign n679 = n50 | n903;
assign n1026 = ~n326;
assign n744 = n1426 & n600;
assign n194 = n781 | n1312;
assign n447 = n1515 & n591;
assign n1739 = ~(n1155 | n1594);
assign n453 = ~(n748 | n1288);
assign n22 = ~(n1166 | n1238);
assign n1264 = ~n19;
assign n1261 = ~(n1388 | n438);
assign n192 = n191 | n1566;
assign n570 = n895 & n1079;
assign n417 = n972 | n997;
assign n659 = n1402 & n929;
assign n671 = n60 & n1121;
assign n250 = ~n548;
assign n1064 = n1690 | n1200;
assign n465 = ~(n378 | n1036);
assign n513 = ~(n743 | n820);
assign n1726 = n311 | n763;
assign n649 = n1613 & n915;
assign n906 = ~(n523 | n504);
assign n1209 = ~(n1553 | n721);
assign n1056 = ~(n625 | n674);
assign n526 = ~(n711 ^ n719);
assign n1160 = n909 & n280;
assign n1773 = n946 & n1118;
assign n446 = ~(n44 | n1154);
assign n532 = ~n403;
assign n485 = n996 & n1356;
assign n1246 = n1205 | n454;
assign n210 = n25 | n609;
assign n1358 = ~n1718;
assign n439 = ~n504;
assign n1747 = ~(n200 | n319);
assign n1268 = n957 | n1200;
assign n34 = n326 | n1590;
assign n176 = n1607 & n536;
assign n678 = ~(n428 ^ n467);
assign n878 = n1131 ^ n364;
assign n664 = n186 | n905;
assign n100 = n472 | n77;
assign n652 = n1466 | n359;
assign n1148 = n307 | n1087;
assign n1010 = n1446 & n317;
assign n374 = n1295 | n1002;
assign n552 = n342 & n1524;
assign n300 = n228 & n1078;
assign n1127 = n252 | n835;
assign n734 = n1295 | n1025;
assign n231 = n1089 | n667;
assign n827 = ~(n1162 | n873);
assign n707 = ~(n200 | n708);
assign n515 = ~(n228 | n289);
assign n783 = n602 | n1061;
assign n235 = n1721;
assign n400 = n1574 | n1413;
assign n802 = ~n715;
assign n1594 = ~(n261 | n796);
assign n1053 = n627 | n75;
assign n456 = n1509 & n1539;
assign n161 = ~(n1146 | n1686);
assign n109 = n1295 | n427;
assign n650 = ~(n1681 | n437);
assign n127 = n1280 | n1208;
assign n578 = ~(n1070 ^ n652);
assign n808 = n1244 & n645;
assign n1787 = n1045 & n484;
assign n925 = ~(n1435 | n714);
assign n1017 = n1464 | n1662;
assign n1143 = ~(n719 ^ n1623);
assign n340 = ~(n539 | n1671);
assign n1532 = ~(n209 | n87);
assign n661 = n72 | n102;
assign n1274 = ~(n377 | n1601);
assign n1599 = ~(n378 | n180);
assign n725 = ~(n44 | n1005);
assign n124 = n1588 & n309;
assign n909 = n154 | n1226;
assign n213 = n1146 & n1628;
assign n45 = ~(n627 | n123);
assign n1037 = n523 | n1312;
assign n1130 = ~(n1401 ^ n1391);
assign n1250 = n60 & n1070;
assign n1128 = ~n676;
assign n673 = n703 & n859;
assign n1447 = n1771 | n1184;
assign n52 = n1797 | n876;
assign n1107 = n1518 & n1662;
assign n290 = n1169 | n268;
assign n1086 = ~(n1166 | n1729);
assign n1013 = ~n1104;
assign n1571 = n825 | n548;
assign n798 = ~(n472 | n807);
assign n959 = n159 | n752;
assign n182 = n789 | n62;
assign n773 = ~(n539 | n1730);
assign n884 = ~(n624 ^ n558);
assign n214 = ~(n1395 | n308);
assign n990 = ~n830;
assign n1527 = ~n1463;
assign n933 = ~(n818 ^ n14);
assign n199 = ~(n378 | n1644);
assign n268 = ~n307;
assign n823 = n1191 | n814;
assign n1059 = ~(n820 ^ n711);
assign n1247 = n1757 | n511;
assign n1654 = ~n457;
assign n1620 = n39 & n1508;
assign n817 = n1341 | n993;
assign n150 = ~n265;
assign n1451 = ~n342;
assign n607 = n1146 | n441;
assign n1270 = ~(n220 | n80);
assign n618 = n764 | n1694;
assign n1301 = ~(n228 | n1214);
assign n249 = ~(n220 | n1371);
assign n1775 = ~n1135;
assign n1607 = n748 | n77;
assign n726 = ~(n228 | n833);
assign n1307 = ~n1180;
assign n1154 = n627 | n259;
assign n94 = n1146 & n1691;
assign n255 = n1388 & n1569;
assign n816 = n1074 | n478;
assign n499 = n1436 & n504;
assign n103 = ~(n560 | n1469);
assign n383 = n961 & n504;
assign n1619 = ~(n1226 ^ n154);
assign n555 = n450 | n579;
assign n712 = ~(n724 | n1529);
assign n1446 = n260 | n192;
assign n1047 = n92 & n457;
assign n655 = n1775 | n1086;
assign n1397 = ~(n1241 ^ n1790);
assign n2 = n956 | n1774;
assign n1634 = ~(n954 | n869);
assign n1077 = n1241 | n1160;
assign n1063 = n117 | n53;
assign n152 = n307 | n454;
assign n1716 = n1490 | n40;
assign n1161 = ~(n708 ^ n1660);
assign n421 = n1541 | n108;
assign n1473 = n851 & n1091;
assign n1474 = ~(n1238 | n1227);
assign n794 = ~(n228 | n279);
assign n165 = ~(n240 | n1389);
assign n173 = n84;
assign n574 = n1703 | n117;
assign n98 = n1146 | n1340;
assign n1539 = ~(n1258 | n164);
assign n25 = ~(n1395 | n838);
assign n42 = ~(n560 | n1478);
assign n1737 = n1383 | n1542;
assign n1690 = ~n1033;
assign n372 = n579 | n1358;
assign n1152 = ~n747;
assign n920 = ~n485;
assign n41 = ~n984;
assign n857 = ~(n481 | n151);
assign n1350 = ~(n134 | n1288);
assign n474 = n626 | n791;
assign n812 = n583 | n1552;
assign n430 = n1645;
assign n1224 = ~(n368 | n1537);
assign n227 = ~n186;
assign n588 = ~(n1395 | n1648);
assign n1157 = n388 | n376;
assign n1295 = ~n579;
assign n987 = n1146 | n1259;
assign n364 = ~(n868 ^ n1161);
assign n271 = ~(n1235 ^ n1231);
assign n1651 = ~(n1435 | n1227);
assign n31 = ~(n377 | n178);
assign n44 = ~n378;
assign n333 = n579 | n28;
assign n278 = ~(n35 ^ n1386);
assign n1343 = n445 | n1725;
assign n65 = n1105 | n319;
assign n577 = ~(n656 | n198);
assign n1529 = ~(n261 | n931);
assign n1000 = ~(n1162 | n522);
assign n693 = n864 | n815;
assign n506 = n1350 | n731;
assign n1784 = ~(n220 | n1328);
assign n1093 = ~(n1664 ^ n466);
assign n1481 = n11 | n160;
assign n958 = n847 | n1514;
assign n865 = ~n962;
assign n320 = ~(n933 ^ n26);
assign n407 = n963 | n221;
assign n1547 = ~(n1166 | n1660);
assign n993 = n265 | n1347;
assign n1717 = ~(n261 | n519);
assign n685 = n499 | n906;
assign n1440 = n495 & n552;
assign n1321 = n966 & n1662;
assign n391 = ~(n748 | n591);
assign n935 = ~(n1618 | n591);
assign n385 = n1136 | n419;
assign n824 = n5 | n1759;
assign n395 = ~n1435;
assign n811 = n1135 & n550;
assign n790 = n1250 | n174;
assign n1085 = ~(n667 ^ n273);
assign n1094 = n1476 | n1777;
assign n587 = n946 & n614;
assign n1630 = n1696 | n1571;
assign n780 = ~(n495 | n1174);
assign n1124 = n186 | n1710;
assign n1762 = ~(n1293 ^ n1051);
assign n1407 = n1210 | n579;
assign n1065 = n220 | n242;
assign n1008 = n307 | n259;
assign n785 = ~(n377 | n1533);
assign n195 = ~(n740 ^ n313);
assign n1430 = n844 | n1694;
assign n536 = ~(n1391 | n1526);
assign n943 = ~(n1700 | n1281);
assign n344 = ~(n228 | n137);
assign n810 = n1125 & n580;
assign n799 = n1477 | n655;
assign n787 = ~(n378 | n969);
assign n138 = ~(n756 | n1521);
assign n1061 = n100 & n1291;
assign n1286 = ~n1768;
assign n1401 = n589 | n425;
assign n1096 = n693 | n1410;
assign n234 = ~n711;
assign n1323 = ~(n200 | n1729);
assign n1544 = ~(n1713 | n591);
assign n701 = n307 | n1495;
assign n1190 = ~n1288;
assign n1081 = ~n335;
assign n1296 = n332 | n1694;
assign n1557 = n319 & n591;
assign n1116 = n148 | n1364;
assign n1273 = n251 | n1614;
assign n357 = ~n566;
assign n207 = ~(n325 ^ n1582);
assign n1253 = ~n9;
assign n309 = n1004 | n1302;
assign n224 = ~(n377 | n1530);
assign n902 = ~(n44 | n1277);
assign n948 = n428 | n920;
assign n1265 = n1307 | n1200;
assign n1584 = n1613 & n912;
assign n1022 = n186 | n469;
assign n481 = ~n147;
assign n1475 = n1205 | n469;
assign n722 = n1772 | n1344;
assign n1665 = ~(n377 | n365);
assign n269 = n579 | n1196;
assign n620 = n904 & n822;
assign n1200 = ~n627;
assign n1457 = n733 | n848;
assign n1543 = n1343 | n834;
assign n1164 = ~n276;
assign n1220 = n718 | n726;
assign n819 = ~(n1570 | n1283);
assign n1656 = n186 | n259;
assign n350 = ~(n380 | n721);
assign n406 = ~(n1395 | n1709);
assign n542 = n84;
assign n1348 = n1295 | n1578;
assign n710 = ~n288;
assign n632 = ~n510;
assign n229 = ~(n377 | n314);
assign n351 = n1292 & n17;
assign n875 = n111 | n227;
assign n1309 = ~(n1039 | n1223);
assign n745 = ~(n1669 | n390);
assign n1186 = ~(n220 | n1317);
assign n646 = n455 | n1567;
assign n792 = ~(n1281 | n1020);
assign n534 = ~(n580 ^ n1125);
assign n43 = n1279 & n1289;
assign n1129 = n1599 | n1062;
assign n1280 = ~n1755;
assign n1390 = n78 | n1641;
assign n325 = ~(n540 | n1711);
assign n1591 = ~n266;
assign n814 = ~(n228 | n432);
assign n533 = ~(n539 | n336);
assign n524 = n1402 | n373;
assign n1316 = n169 | n1403;
assign n1684 = n1500 | n1556;
assign n527 = ~(n261 | n890);
assign n1778 = ~(n261 | n1348);
assign n941 = n643 & n1662;
assign n263 = ~n1125;
assign n1 = ~(n940 ^ n122);
assign n1421 = ~(n1448 | n414);
assign n114 = ~(n745 | n167);
assign n1570 = ~n0;
assign n120 = n188 | n1312;
assign n1420 = ~(n472 | n1288);
assign n1491 = n1286 | n1574;
assign n929 = n1557 | n163;
assign n280 = ~n1236;
assign n873 = n307 | n1631;
assign n431 = ~(n1342 ^ n1783);
assign n20 = ~(n272 | n1763);
assign n363 = n1573 | n1031;
assign n3 = n1126 | n268;
assign n594 = n1146 | n563;
assign n1174 = n1041 | n1451;
assign n1596 = n569 | n327;
assign n205 = n1017 & n1472;
assign n1699 = ~(n669 | n1288);
assign n886 = n1019 & n1188;
assign n416 = n512 | n181;
assign n73 = n1194 | n1146;
assign n1345 = ~(n261 | n622);
assign n1552 = ~(n706 | n867);
assign n486 = ~n850;
assign n1497 = ~(n228 | n153);
assign n1337 = n395 | n1312;
assign n181 = ~(n1395 | n1073);
assign n602 = n1755 & n69;
assign n204 = n1081 | n1200;
assign n747 = n529 | n54;
assign n226 = ~(n560 | n664);
assign n56 = ~(n220 | n1399);
assign n898 = ~(n617 | n1519);
assign n1272 = n23 | n106;
assign n549 = ~n1579;
assign n675 = ~n321;
assign n716 = n1435 & n1288;
assign n1339 = ~(n1175 | n644);
assign n1794 = ~(n220 | n1723);
assign n1537 = n1596 | n1467;
assign n1611 = ~(n378 | n1064);
assign n1425 = n1534;
assign n1639 = ~(n1162 | n1148);
assign n1121 = n1549 | n1202;
assign n1131 = ~(n1284 ^ n177);
assign n592 = ~(n798 | n672);
assign n1723 = ~(n210 | n1159);
assign n1695 = n23 | n880;
assign n498 = ~(n560 | n597);
assign n1118 = ~n591;
assign n148 = n579 & n261;
assign n393 = n988 | n820;
assign n1441 = ~(n378 | n1053);
assign n1386 = ~(n1638 ^ n581);
assign n493 = n1585 | n1719;
assign n1517 = ~(n228 | n888);
assign n281 = n1295 | n870;
assign n1617 = ~(n377 | n1576);
assign n1736 = ~n1313;
assign n1637 = ~(n1162 | n290);
assign n786 = ~(n220 | n1505);
assign n1492 = ~n668;
assign n1770 = ~(n593 | n201);
assign n970 = ~(n377 | n1071);
assign n719 = ~(n901 ^ n697);
assign n426 = ~(n342 | n491);
assign n626 = n1391 & n1401;
assign n654 = ~(n1535 ^ n1423);
assign n1567 = n1423 | n1014;
assign n177 = ~(n1729 ^ n319);
assign n1248 = n952 | n268;
assign n1183 = n458 | n43;
assign n1144 = n1143 & n820;
assign n1625 = n1205 | n1346;
assign n1601 = n1178 | n268;
assign n1641 = n1305 | n692;
assign n1042 = n197 | n268;
assign n853 = ~n1043;
assign n575 = n1564 | n299;
assign n1149 = n1286 | n1222;
assign n1328 = ~(n823 | n653);
assign n1530 = n307 | n1314;
assign n475 = ~(n1125 | n27);
assign n302 = ~(n652 ^ n1575);
assign n743 = n159 & n752;
assign n1168 = n194 & n604;
assign n101 = n223 | n1030;
assign n1032 = n1404 | n1611;
assign n1234 = n1674 & n439;
assign n531 = ~n896;
assign n365 = n307 | n75;
assign n368 = n737 | n1144;
assign n831 = ~(n1498 | n1519);
assign n945 = n1046 | n1114;
assign n1029 = ~(n1160 ^ n1695);
assign n1439 = n319 & n1288;
assign n1512 = ~(n1130 ^ n945);
assign n483 = n600 & n541;
assign n301 = n1146 | n1057;
assign n623 = n1622 | n1063;
assign n672 = ~(n1553 | n714);
assign n30 = ~(n378 | n142);
assign n1735 = n900 | n227;
assign n66 = n389;
assign n899 = n490 | n227;
assign n1757 = ~(n539 | n728);
assign n651 = ~(n669 | n1118);
assign n1044 = ~n918;
assign n546 = n1204 & n884;
assign n667 = ~n88;
assign n728 = n1522 | n227;
assign n795 = n295 | n346;
assign n848 = n1515 & n1662;
assign n1468 = ~(n216 ^ n509);
assign n1728 = ~(n472 | n504);
assign n216 = ~(n686 ^ n39);
assign n1294 = ~(n288 ^ n1518);
assign n240 = n334 | n800;
assign n1376 = n48 & n727;
assign n129 = n566;
assign n537 = ~n841;
assign n1769 = n1773 | n638;
assign n1236 = n493 | n430;
assign n155 = ~n1636;
assign n360 = ~(n534 ^ n1457);
assign n1191 = ~(n1395 | n618);
assign n1389 = n415 | n855;
assign n704 = ~(n261 | n369);
assign n782 = n990 | n1694;
assign n1311 = n1295 | n1085;
assign n354 = n1205 | n456;
assign n522 = n1689 | n268;
assign n1370 = ~n92;
assign n136 = n610 | n293;
assign n1786 = n1628 | n131;
assign n753 = ~(n186 | n123);
assign n922 = n117 | n943;
assign n1228 = n503 | n444;
assign n72 = n96 | n1262;
assign n500 = n531 & n43;
assign n53 = ~(n257 | n1281);
assign n253 = ~(n1162 | n470);
assign n1036 = n1419 | n1200;
assign n468 = ~(n1672 ^ n1770);
assign n1112 = ~(n1162 | n1248);
assign n32 = ~(n748 | n807);
assign n452 = n1637 | n1459;
assign n316 = ~(n1395 | n1683);
assign n115 = n1791 | n268;
assign n571 = ~n1175;
assign n382 = ~n195;
assign n1504 = n1326;
assign n1417 = ~n813;
assign n803 = n340 | n911;
assign n418 = ~(n757 | n590);
assign n1713 = ~n1498;
assign n1793 = ~n1524;
assign n633 = n702 | n1200;
assign n285 = ~(n1395 | n4);
assign n1204 = n121 & n20;
assign n681 = n1485 & n504;
assign n291 = n1545 & n909;
assign n74 = n1146 | n1303;
assign n283 = n1256 & n1706;
assign n629 = ~(n377 | n1042);
assign n348 = ~(n1565 | n1566);
assign n1797 = ~(n560 | n1722);
assign n509 = n741 | n809;
assign n298 = ~n238;
assign n1561 = ~(n560 | n1285);
assign n144 = ~(n261 | n691);
assign n1049 = ~n663;
assign n1466 = n801 & n504;
assign n713 = n453 | n350;
assign n703 = ~n1327;
assign n750 = ~(n380 | n714);
assign n1314 = n987 & n861;
assign n724 = ~(n261 | n551);
assign n1708 = n562 & n46;
assign n267 = n1337 & n1434;
assign n1365 = ~(n560 | n968);
assign n885 = ~(n378 | n1006);
assign n401 = n209 & n1235;
assign n1235 = ~n149;
assign n254 = ~n1299;
assign n346 = n1137 & n410;
assign n872 = ~(n1175 | n546);
assign n1629 = n1054 | n227;
assign n1449 = n120 & n769;
assign n855 = n687 | n1428;
assign n331 = n669 | n614;
assign n1572 = n1128 | n268;
assign n818 = ~(n1585 ^ n1241);
assign n605 = n103 | n1525;
assign n327 = n1550 | n1506;
assign n89 = ~(n1226 ^ n1566);
assign n1521 = ~(n261 | n1193);
assign n112 = ~n448;
assign n324 = n462 | n1200;
assign n107 = n1672 & n1331;
assign n1217 = ~(n243 ^ n1623);
assign n459 = ~(n233 | n1320);
assign n68 = n946 & n1662;
assign n879 = ~(n1162 | n1318);
assign n767 = n843 | n440;
assign n1582 = ~(n1727 | n977);
assign n1315 = n411 & n475;
assign n1271 = ~(n560 | n341);
assign n1694 = ~n1205;
assign n441 = n1041 | n579;
assign n1245 = ~(n579 | n1229);
assign n1371 = ~(n1102 | n816);
assign n1646 = ~n1088;
assign n246 = ~(n539 | n1656);
assign n376 = ~(n539 | n1548);
assign n308 = n1205 | n1087;
assign n1156 = ~(n1166 | n1435);
assign n1719 = ~n258;
assign n1381 = n342 | n1358;
assign n1021 = n184 & n1098;
assign n1303 = n1492 | n579;
assign n339 = ~n371;
assign n998 = ~n1083;
assign n489 = ~n1638;
assign n40 = n792;
assign n140 = ~(n323 | n1176);
assign n1585 = n287 | n1107;
assign n409 = n579 & n195;
assign n637 = ~(n1515 ^ n643);
assign n299 = n261 | n409;
assign n1006 = n1785 | n1200;
assign n1578 = n1132 & n735;
assign n1259 = n1170 | n579;
assign n947 = ~n1512;
assign n756 = ~(n261 | n269);
assign n905 = n49 & n1786;
assign n1113 = n1146 & n1564;
assign n1795 = ~n1244;
assign n118 = n186 | n1631;
assign n910 = n627 | n1495;
assign n1558 = n1441 | n1452;
assign n1752 = n483 | n941;
assign n763 = ~n231;
assign n1070 = n358 | n1310;
assign n558 = ~(n526 ^ n949);
assign n260 = ~(n1585 | n1545);
assign n241 = ~(n1745 | n212);
assign n1499 = ~(n1162 | n141);
assign n490 = ~n1119;
assign n1501 = n147 & n1382;
assign n1765 = ~(n228 | n1266);
assign n5 = n1379 | n1617;
assign n1583 = ~(n1619 ^ n1029);
assign n1721 = n1520 & n477;
assign n871 = n1604 | n1114;
assign n4 = n1205 | n1631;
assign n508 = n887 & n504;
assign n219 = ~(n1395 | n1475);
assign n123 = n471 & n51;
assign n424 = n134 | n77;
assign n1631 = n301 & n1444;
assign n1443 = ~(n216 ^ n10);
assign n1556 = ~(n560 | n1629);
assign n414 = n238 & n1118;
assign n705 = n794 | n1040;
assign n843 = ~(n1395 | n782);
assign n1423 = n136 & n34;
assign n1216 = n398 | n1200;
assign n478 = ~(n44 | n303);
assign n225 = ~(n307 | n123);
assign n501 = n966 & n614;
assign n545 = ~(n1544 | n1324);
assign n93 = ~(n560 | n621);
assign n739 = ~(n391 | n892);
assign n599 = n1146 | n1483;
assign n1394 = n725 | n1221;
assign n1549 = n708 & n591;
assign n265 = n799 & n1487;
assign n1734 = n1112 | n1712;
assign n106 = ~n154;
assign n895 = ~(n1367 | n787);
assign n449 = ~(n377 | n700);
assign n1222 = n400 | n1593;
assign n644 = ~(n927 ^ n126);
assign n1764 = ~(n1345 | n1608);
assign n35 = ~(n1421 ^ n736);
assign n289 = n1205 | n487;
assign n1199 = ~n1645;
assign n29 = ~(n261 | n1479);
assign n375 = n84;
assign n206 = ~(n377 | n1486);
assign n653 = n8 | n285;
assign n1673 = ~n1229;
assign n126 = ~(n47 ^ n431);
assign n1104 = n896 | n216;
assign n914 = n720 | n268;
assign n1685 = ~n1089;
assign n963 = n1729 & n591;
assign n1404 = ~(n44 | n1438);
assign n1322 = n220 | n570;
assign n1069 = ~n1578;
assign n1593 = n547 | n976;
assign n158 = ~(n220 | n856);
assign n1434 = n1105 | n1435;
assign n1239 = ~(n228 | n1060);
assign n444 = ~(n395 | n600);
assign n1510 = n1732 | n1055;
assign n736 = ~(n739 | n1052);
assign n201 = ~(n1575 | n738);
assign n1680 = ~(n438 ^ n1412);
assign n470 = n307 | n370;
assign n454 = n196 & n1455;
assign n1293 = ~(n149 ^ n1668);
assign n466 = n1620 | n1373;
assign n1760 = n1791 | n227;
assign n1001 = ~(n377 | n1513);
assign n896 = ~(n747 ^ n1039);
assign n1215 = ~(n261 | n1528);
assign n79 = ~n601;
assign n942 = ~(n832 | n617);
assign n1083 = n1295 | n382;
assign n164 = ~(n261 | n374);
assign n1054 = ~n760;
assign n1379 = ~(n1162 | n914);
assign n596 = n1481 | n183;
assign n1139 = ~(n1162 | n768);
assign n167 = n1366 | n772;
assign n1650 = n1287 | n885;
assign n450 = ~n1095;
assign n1193 = n1295 | n561;
assign n1327 = ~(n1070 ^ n60);
assign n1605 = ~(n1457 ^ n1752);
assign n1302 = ~n15;
assign n169 = ~n1402;
assign n318 = ~(n767 | n37);
assign n1335 = ~(n935 | n1278);
assign n203 = n1502 | n498;
assign n1166 = ~n721;
assign n1114 = ~n1255;
assign n1385 = n1326;
assign n548 = n363 | n896;
assign n147 = ~(n1308 ^ n1402);
assign n1324 = n1433 | n641;
assign n1210 = ~n1633;
assign n1109 = ~(n904 | n15);
assign n78 = n143 | n629;
assign n314 = n995 | n268;
assign n866 = n1369 | n97;
assign n1645 = n23 & n106;
assign n125 = ~(n539 | n118);
assign n145 = ~(n408 ^ n1401);
assign n37 = n1754 | n300;
assign n217 = n307 | n1110;
assign n727 = ~(n39 | n898);
assign n1123 = n620 | n1109;
assign n1698 = n673;
assign n104 = ~(n1162 | n991);
assign n131 = n261 | n1325;
assign n6 = ~(n781 | n504);
assign n1399 = ~(n573 | n1609);
assign n256 = ~(n560 | n1760);
assign n1671 = n720 | n227;
assign n1683 = n1205 | n1710;
assign n188 = ~n1660;
assign n1212 = n821 | n227;
assign n1359 = n913 | n1728;
assign n1636 = n538 & n1507;
assign n1197 = ~(n1612 | n1206);
assign n683 = ~(n57 | n306);
assign n440 = ~(n228 | n1782);
assign n1414 = n790 | n1450;
assign n402 = ~n1471;
assign n1103 = n1336 | n1230;
assign n1075 = ~n1361;
assign n877 = n1072 | n1200;
assign n852 = n1146 | n555;
assign n968 = n186 | n1495;
assign n638 = n1147 | n1405;
assign n832 = ~n1227;
assign n978 = n1235 & n87;
assign n1310 = n708 & n439;
assign n1375 = ~n128;
assign n1240 = n1742 | n612;
assign n769 = n1105 | n1660;
assign n928 = n1678 | n443;
assign n8 = ~(n228 | n742);
assign n1308 = ~n685;
assign n535 = ~(n395 | n807);
assign n1038 = ~(n1228 ^ n580);
assign n274 = n275 | n248;
assign n995 = ~n384;
assign n1170 = ~n1740;
assign n404 = ~(n761 ^ n380);
assign n1330 = n1789 | n1651;
assign n804 = ~(n808 ^ n1470);
assign n1777 = n1726 | n1275;
assign n645 = ~n55;
assign n1453 = n1146 | n82;
assign n480 = ~(n378 | n230);
assign n392 = n428 | n854;
assign n99 = n716 | n362;
assign n1340 = n41 | n579;
assign n86 = ~(n832 | n1515);
assign n749 = ~(n495 | n1381);
assign n423 = n1610 | n227;
assign n445 = ~(n1162 | n775);
assign n1478 = n1178 | n227;
assign n689 = ~n678;
assign n1514 = ~(n1172 | n1227);
assign n523 = ~n319;
assign n233 = n1351 | n939;
assign n1419 = ~n530;
assign n292 = ~(n1781 | n1778);
assign n1476 = n88 & n500;
assign n809 = ~n10;
assign n355 = n1585 | n1004;
assign n597 = n197 | n227;
assign n752 = ~n719;
assign n1666 = n1724 | n446;
assign n367 = n1204 | n1643;
assign n1672 = n671 | n171;
assign n1057 = n1624 | n579;
assign n1162 = ~n377;
assign n1482 = ~(n44 | n965);
assign n547 = n1203 ^ n1677;
assign n1418 = n1699 | n21;
assign n1225 = n266 | n278;
assign n1618 = ~n1238;
assign n1352 = ~(n966 | n714);
assign n156 = n1253 | n579;
assign n502 = n494 | n1315;
assign n262 = ~(n220 | n665);
assign n200 = ~n714;
assign n1523 = n1241 | n1236;
assign n329 = n571 | n170;
assign n1484 = ~(n134 | n807);
assign n1424 = n1126 | n227;
assign n1489 = ~(n1293 ^ n1461);
assign n122 = n458 | n1289;
assign n608 = n658 | n1200;
assign n294 = n659 | n1787;
assign n419 = n284 | n948;
assign n718 = ~(n1395 | n598);
assign n1243 = ~(n134 | n591);
assign n1214 = n1205 | n75;
assign n980 = ~(n200 | n617);
assign n1395 = ~n228;
assign n1266 = n1205 | n905;
assign n1117 = ~(n1162 | n217);
assign n584 = n560 & n753;
assign n59 = ~n901;
assign n825 = ~n88;
assign n927 = ~(n1443 ^ n576);
assign n1488 = ~n386;
assign n858 = ~(n1198 | n1717);
assign n1115 = ~(n378 | n660);
assign n1231 = n155 & n1108;
assign n1658 = ~(n261 | n1267);
assign n1080 = n1615 | n579;
assign n634 = n825 | n1104;
assign n1076 = n957 | n1694;
assign n859 = n1437 & n1501;
assign n569 = n1368 | n663;
assign n994 = ~(n1605 ^ n1038);
assign n151 = ~n1476;
assign n797 = ~(n1100 | n1431);
assign n258 = n1026 | n434;
assign n991 = n307 | n469;
assign n658 = ~n270;
assign n1151 = n872 & n367;
assign n1122 = ~n190;
assign n1555 = ~(n1236 ^ n286);
assign n1526 = ~(n380 | n1519);
assign n1774 = ~n1501;
assign n27 = ~(n200 | n1043);
assign n988 = ~(n703 ^ n397);
assign n821 = ~n1150;
assign n185 = ~n743;
assign n1574 = ~n119;
assign n1465 = n61 | n1661;
assign n323 = n433 | n619;
assign n358 = n1408 & n504;
assign n359 = ~(n188 | n504);
assign n1071 = n1432 | n268;
assign n528 = n1139 | n970;
assign n1091 = n1100 | n351;
assign n529 = n1632 & n504;
assign n1662 = ~n600;
assign n1263 = ~(n1484 | n839);
assign n189 = n865 | n1694;
assign n972 = n1000 | n1001;
assign n517 = ~(n686 ^ n975);
assign n252 = ~n948;
assign n17 = n1105 | n1238;
assign n1098 = n1575 | n1449;
assign n212 = ~(n261 | n950);
assign n788 = ~(n1034 | n705);
assign n612 = ~(n1498 | n721);
assign n81 = n1125 | n886;
assign n379 = n1613 & n172;
assign n1262 = ~(n560 | n875);
assign n630 = ~n1575;
assign n1659 = n953 | n1696;
assign n28 = ~n1535;
assign n733 = ~(n1676 | n1662);
assign n1780 = n84 & n1058;
assign n36 = ~(n587 | n208);
assign n849 = ~n516;
assign n311 = ~n953;
assign n108 = ~(n1162 | n1496);
assign n1002 = ~n368;
assign n343 = ~(n1553 | n1519);
assign n981 = n1384 | n634;
assign n1486 = n307 | n487;
assign n154 = ~(n717 ^ n326);
assign n83 = n1247 | n505;
assign n1284 = ~(n1024 ^ n863);
assign n926 = ~(n579 | n274);
assign n1608 = ~(n261 | n1311);
assign n1689 = ~n754;
assign n1136 = ~n1788;
assign n1317 = ~(n1447 | n322);
assign n1628 = n1225 & n1581;
assign n1495 = n852 & n1627;
assign n648 = n1396 & n504;
assign n434 = ~n717;
assign n1686 = ~n33;
assign n1472 = n710 | n600;
assign n854 = n996 | n534;
assign n1643 = ~(n804 ^ n666);
assign n1313 = n1551 | n1376;
assign n1377 = n553 | n730;
assign n1102 = n554 | n199;
assign n1445 = ~(n747 ^ n1579);
assign n1531 = n1016 | n267;
assign n657 = n924 | n579;
assign n1134 = ~(n818 ^ n291);
assign n1456 = n1522 | n268;
assign n1730 = n1264 | n227;
assign n328 = ~(n642 ^ n557);
assign n1455 = ~(n29 | n71);
assign n939 = ~(n378 | n1265);
assign n415 = n979 | n784;
assign n1559 = ~(n134 | n504);
assign n883 = ~(n44 | n891);
assign n1536 = ~(n1585 ^ n291);
assign n1624 = ~n157;
assign n1073 = n1205 | n1110;
assign n793 = n544;
assign n589 = n1707 & n600;
assign n860 = n623;
assign n583 = n706 & n1597;
assign n492 = ~(n228 | n1246);
assign n863 = ~(n1238 ^ n1498);
assign n1089 = n1433 | n1152;
assign n1289 = ~n216;
assign n174 = n1106 & n703;
assign n1573 = ~n39;
assign n1479 = n579 | n1638;
assign n487 = n594 & n1158;
assign n778 = ~(n966 ^ n946);
assign n1108 = n1532 & n392;
assign n1137 = n781 | n614;
assign n1249 = ~(n1195 ^ n1415);
assign n1388 = n169 | n1308;
assign n1138 = n486 | n579;
assign n1025 = ~(n996 ^ n1788);
assign n662 = n1406 | n36;
assign n113 = n627 | n454;
assign n455 = n1171 | n1535;
assign n916 = ~(n485 | n412);
assign n1398 = n630 | n1547;
assign n102 = n226 | n1099;
assign n305 = n186 | n454;
assign n663 = ~(n896 ^ n1183);
assign n695 = ~(n1395 | n805);
assign n771 = ~(n1660 | n1227);
assign n761 = ~(n637 ^ n670);
assign n1332 = ~n1737;
assign n420 = ~(n261 | n1012);
assign n1687 = ~(n1650 | n1652);
assign n413 = n528 | n1738;
assign n47 = ~(n1777 ^ n363);
assign n1165 = n1662 | n1568;
assign n1483 = n1372 | n579;
assign n1334 = ~n1743;
assign n834 = n785 | n253;
assign n1331 = ~(n817 | n182);
assign n116 = ~(n378 | n1260);
assign n1562 = ~(n539 | n1124);
assign n1367 = ~(n44 | n521);
assign n451 = ~n1219;
assign n1467 = n496 | n1387;
assign n876 = ~(n539 | n985);
assign n1767 = ~(n1395 | n1430);
assign n901 = n681 | n1559;
assign n1507 = n1788 & n485;
assign n1727 = ~(n1243 | n958);
assign n1019 = n853 | n1312;
assign n117 = n79 | n537;
assign n1079 = ~(n1115 | n1606);
assign n1356 = ~n534;
assign n687 = n146 | n89;
assign n1187 = n1205 | n1314;
assign n940 = ~(n1626 | n1777);
assign n1586 = n186 | n1346;
assign n953 = n992 | n549;
assign n135 = ~(n1276 | n420);
assign n692 = ~(n1162 | n1008);
assign n1078 = ~(n1205 | n123);
assign n954 = n897 | n1616;
assign n1565 = ~(n1236 ^ n205);
assign n892 = n345 | n1007;
assign n1275 = ~n1571;
assign n573 = n406 | n1538;
assign n609 = ~(n228 | n304);
assign n170 = ~(n0 | n766);
assign n1374 = ~n1010;
assign n861 = ~(n237 | n1658);
assign n1256 = n205 | n1360;
assign n686 = n648 | n202;
assign n639 = n1295 | n1776;
assign n581 = ~(n1702 ^ n502);
assign n1169 = ~n179;
assign n1062 = n378 & n45;
assign n665 = ~(n1394 | n1666);
assign n772 = ~(n296 | n1489);
assign n1602 = n582 | n93;
assign n559 = ~(n1645 | n1164);
assign n1354 = ~(n1016 | n1516);
assign n1748 = ~(n1238 | n714);
assign n1626 = ~n634;
assign n422 = ~n132;
assign n1027 = n607 & n135;
assign n313 = n1151 | n1705;
assign n1111 = n627 | n882;
assign n296 = ~n1669;
assign n180 = n627 | n1027;
assign n1020 = ~n1181;
assign n1506 = ~(n481 ^ n1094);
assign n874 = n490 | n268;
assign n1733 = ~(n220 | n1634);
assign n247 = n627 | n487;
assign n1267 = n1295 | n689;
assign n1746 = n1295 | n1049;
assign n427 = ~n1680;
assign n624 = ~(n1470 ^ n1795);
assign n1701 = ~(n703 | n243);
assign n800 = n1192 & n1566;
assign n839 = ~(n1172 | n714);
assign n983 = n1689 | n227;
assign n1146 = ~n261;
assign n1461 = ~(n534 ^ n919);
assign n1732 = n688 | n42;
assign n1052 = ~(n1391 | n1009);
assign n613 = ~n639;
assign n50 = ~n353;
assign n982 = ~(n539 | n983);
assign n341 = n186 | n168;
assign n640 = n1128 | n227;
assign n273 = ~(n1342 | n500);
assign n46 = ~(n699 | n646);
assign n757 = n238 & n1165;
assign n243 = n1437 | n397;
assign n603 = n1133 | n755;
assign n1715 = ~(n261 | n109);
assign n957 = ~n1675;
assign n275 = n697 & n506;
assign n590 = n401 | n978;
assign n720 = ~n564;
assign n1444 = ~(n527 | n1715);
assign n934 = n1146 & n1082;
assign n276 = n385 & n1004;
assign n1490 = n1326 | n650;
assign n425 = ~(n748 | n600);
assign n869 = n30 | n883;
assign n567 = ~(n220 | n1687);
assign n582 = ~(n539 | n423);
assign n977 = ~(n697 | n1263);
assign n615 = ~(n377 | n1068);
assign n1230 = n263 | n1621;
assign n965 = n802 | n1200;
assign n986 = ~(n188 | n591);
assign n610 = n966 & n1118;
assign n463 = ~(n438 | n825);
assign n1346 = n1090 & n1056;
assign n1004 = n1173 & n682;
assign n738 = ~(n1023 | n166);
assign n1189 = ~n586;
assign n791 = n757 & n1668;
assign n1373 = n331 & n989;
assign n51 = ~(n934 | n932);
assign n1564 = n679 & n1667;
assign n1387 = n1069 | n1595;
assign n1610 = ~n297;
assign n730 = n1458 | n827;
assign n1595 = ~n870;
assign n677 = ~(n514 | n1204);
assign n87 = n810 & n538;
assign n1493 = ~(n1395 | n1066);
assign n867 = ~n1643;
assign n222 = ~(n220 | n577);
assign n322 = n429 | n1179;
assign n1342 = n1685 | n250;
assign n576 = ~(n88 ^ n531);
assign n69 = n1420 | n1209;
assign n411 = n853 | n614;
assign n1705 = n1175 & n812;
assign n1045 = n523 | n614;
assign n789 = n1021 | n497;
assign n462 = ~n387;
assign n172 = n1385 | n1273;
assign n1459 = ~(n377 | n1252);
assign n631 = ~(n1681 | n38);
assign n1709 = n702 | n1694;
assign n362 = n1789 | n1156;
assign n969 = n774 | n1200;
assign n1581 = ~(n579 | n1731);
assign n1704 = ~(n1498 | n714);
assign n911 = ~(n560 | n1735);
assign n1664 = ~(n1141 ^ n110);
assign n777 = n847 | n59;
assign n171 = n1333 & n1577;
assign n915 = n399 | n928;
assign n1464 = ~n389;
assign n1545 = n258 & n1199;
assign n1502 = ~(n539 | n640);
assign n951 = n631 | n922;
assign n1005 = n332 | n1200;
assign n1014 = ~n1145;
assign n837 = ~(n378 | n247);
assign n851 = n105 | n461;
assign n806 = n518 | n820;
assign n960 = ~n271;
assign n1588 = ~(n1366 | n690);
assign n0 = ~(n751 ^ n1468);
assign n352 = n1307 | n1694;
assign n1229 = n921 | n1306;
assign n1163 = n1527 | n117;
assign n844 = ~n1353;
assign n870 = n393 & n866;
assign n315 = ~(n220 | n788);
assign n964 = n1392 & n1197;
assign n729 = n186 | n1087;
assign n244 = ~n1473;
assign n1255 = n460 & n418;
assign n1142 = ~(n1127 ^ n871);
assign n822 = ~n328;
assign n1173 = n284 | n392;
assign n833 = n1375 | n1694;
assign n1566 = ~n276;
assign n196 = n1146 | n657;
assign n1360 = ~n1160;
assign n593 = ~(n986 | n1592);
assign n438 = ~(n550 ^ n1135);
assign n1372 = ~n999;
assign n1211 = ~n274;
assign n1623 = n159 | n234;
assign n467 = n1507 | n412;
assign n76 = n366 | n1153;
assign n349 = n277 | n246;
assign n563 = n1075 | n579;
assign n1050 = ~(n220 | n459);
assign n1298 = ~n779;
assign n1031 = ~n686;
assign n1276 = ~(n261 | n372);
assign n635 = n1734 | n923;
assign n709 = n148 | n161;
assign n1606 = ~(n44 | n556);
assign n1383 = n1518 & n591;
assign n938 = n124 | n543;
assign n997 = n615 | n973;
assign n1349 = ~(n560 | n595);
assign n405 = ~(n1762 ^ n16);
assign n1305 = ~(n377 | n152);
assign n1092 = n1146 | n162;
assign n622 = n579 | n244;
assign n1269 = n1411 & n1167;
assign n193 = ~n937;
assign n96 = ~(n539 | n836);
assign n625 = n1146 & n1245;
assign n88 = ~(n549 ^ n1100);
assign n1678 = ~(n1681 | n532);
assign n1178 = ~n239;
assign n1233 = n1044;
assign n1542 = ~(n832 | n1518);
assign n1792 = ~(n302 ^ n808);
assign n1771 = ~(n44 | n204);
assign n1587 = ~(n220 | n1679);
assign n1500 = ~(n539 | n58);
assign n1364 = ~(n1146 | n422);
assign n370 = n98 & n683;
assign n1392 = n1146 | n1080;
assign n1791 = ~n955;
assign n111 = ~n1756;
assign n412 = n810 | n696;
assign n1494 = n1295 | n907;
assign n1589 = n1718 | n586;
assign n711 = ~(n1359 ^ n1755);
assign n740 = ~(n1339 | n1300);
assign n989 = ~(n39 | n980);
assign n1413 = n849 | n878;
assign n1232 = n1366 & n405;
assign n62 = n1673 | n1736;
assign n641 = ~(n1498 | n1227);
assign n1644 = n1334 | n1200;
assign n1759 = n224 | n1117;
assign n1710 = n599 & n138;
assign n1378 = n84;
assign n1198 = n1146 & n1120;
assign n1635 = ~(n1618 | n504);
assign n15 = ~(n1134 ^ n1583);
assign n696 = ~n854;
assign n1776 = ~(n938 ^ n684);
assign n54 = ~(n1713 | n504);
assign n737 = n959 & n513;
assign n1140 = ~n1568;
assign n58 = n1169 | n227;
assign n334 = n1272 & n559;
assign n146 = ~n1025;
assign n1176 = n492 | n1493;
assign n766 = ~n1283;
assign n153 = n658 | n1694;
assign n751 = ~(n147 ^ n531);
assign n765 = n1044;
assign n1551 = n39 & n1418;
assign n1712 = ~(n377 | n312);
assign n904 = n419 & n1004;
assign n1278 = n992 | n1474;
assign n1067 = ~(n853 | n600);
assign n604 = n1105 | n1729;
assign n142 = n627 | n1314;
assign n1592 = n630 | n771;
assign n1590 = ~(n501 | n1352);
assign n105 = n1238 & n1288;
assign n755 = ~(n1281 | n451);
assign n1416 = n481 | n231;
assign n976 = n1511 | n320;
assign n1577 = ~(n60 | n707);
assign n1384 = n438 | n481;
assign n514 = n1327 | n1750;
assign n924 = ~n1753;
assign n471 = n1146 | n1138;
assign n284 = n149 | n1130;
assign n1084 = ~(n1395 | n189);
assign n1192 = ~(n154 ^ n1695);
assign n16 = ~(n1142 ^ n360);
assign n836 = n952 | n227;
assign n553 = n90 | n1274;
assign n10 = n1630 & n255;
assign n556 = n627 | n469;
assign n1682 = n130;
assign n1258 = n1146 & n926;
assign n1706 = n1077 & n1164;
assign n497 = n1442 & n524;
assign n1638 = n447 | n86;
assign n776 = n1613;
assign n619 = ~(n228 | n1076);
assign n732 = n1146 | n1688;
assign n1505 = ~(n1220 | n1185);
assign n882 = n1092 & n1739;
assign n221 = ~(n832 | n1729);
assign n1072 = ~n1362;
assign n949 = ~(n397 ^ n826);
assign n1068 = n307 | n1027;
assign n396 = ~n302;
assign n835 = ~n1108;
assign n1796 = n703 & n1257;
assign n1422 = ~n1059;
assign n1074 = ~(n378 | n910);
assign n408 = ~n1165;
assign n479 = ~n636;
assign n1009 = ~(n32 | n750);
assign n70 = ~(n464 | n1558);
assign n921 = n1039 & n1240;
assign n197 = ~n1207;
assign n1738 = n31 | n1499;
assign n764 = ~n236;
assign n1213 = n1504 | n603;
assign n356 = n238 | n77;
assign n264 = ~(n1465 | n1149);
assign n1196 = ~n497;
assign n1159 = n515 | n316;
assign n1563 = n627 | n1087;
assign n543 = n1366 & n1123;
assign n272 = n811 | n1261;
assign n410 = ~(n1135 | n1323);
assign n1251 = ~(n1039 | n831);
assign n442 = n1332 | n489;
assign n1312 = ~n77;
assign n477 = ~(n909 | n419);
assign n538 = n1228 ^ n1016;
assign n149 = n408 ^ n238;
assign n390 = ~n1489;
assign n985 = n186 | n1110;
assign n1325 = ~(n1295 | n1776);
assign n1703 = ~n1454;
assign n702 = ~n7;
assign n496 = n1680 | n1059;
assign n80 = ~(n568 | n416);
assign n598 = n802 | n1694;
assign n1018 = n1432 | n227;
assign n1242 = n627 | n1346;
assign n680 = n627 | n1710;
assign n568 = n1393 | n1239;
assign n1382 = n463 & n1013;
assign n796 = n1295 | n1720;
assign n682 = ~(n474 | n218);
assign n1511 = n404 ^ n1035;
assign n1462 = ~(n220 | n318);
assign n923 = n449 | n104;
assign n1277 = n627 | n370;
assign n1513 = n694 | n268;
assign n1223 = ~(n330 | n1704);
assign n304 = n1785 | n1694;
assign n1203 = ~(n1647 ^ n1048);
assign n306 = ~(n261 | n1546);
assign n694 = ~n1177;
assign n55 = n752 & n234;
assign n820 = ~n628;
assign n868 = ~(n1172 ^ n1553);
assign n18 = n1201 | n1157;
assign n139 = ~(n1084 | n1517);
assign n521 = n865 | n1200;
assign n163 = ~(n832 | n319);
assign n310 = n186 | n964;
assign n900 = ~n1655;
assign n908 = n1610 | n268;
assign n580 = n1015 | n1067;
assign n1133 = ~(n1681 | n1646);
assign n510 = ~(n534 ^ n1237);
assign n1688 = n1122 | n579;
assign n1554 = ~(n1395 | n1625);
assign n642 = ~(n818 ^ n1766);
assign n717 = n744 | n1321;
assign n484 = ~(n1402 | n1747);
assign n1326 = n117;
assign n1208 = ~(n1553 | n1227);
assign n21 = ~(n617 | n721);
assign n1024 = ~(n617 ^ n1674);
assign n621 = n995 | n227;
assign n460 = n149 | n392;
assign n381 = n803 | n52;
assign n1758 = n579 | n1737;
assign n1028 = n579 | n936;
assign n688 = ~(n539 | n899);
assign n731 = ~(n1172 | n721);
assign n1789 = ~n1016;
assign n1226 = ~(n507 ^ n1406);
assign n893 = ~(n228 | n85);
assign n1657 = n389;
assign n1653 = ~(n44 | n680);
assign n1405 = ~(n946 | n1227);
assign n1477 = n1729 & n1288;
assign n472 = ~n1553;
assign n1714 = n307 | n168;
assign n897 = ~(n44 | n1216);
assign n952 = ~n187;
assign n1105 = ~n1519;
assign n1126 = ~n1540;
assign n1015 = ~(n112 | n1662);
assign n1621 = ~(n1166 | n1043);
assign n198 = n1254 | n902;
assign n967 = n357;
assign n1120 = ~(n579 | n1313);
assign n473 = n1767 | n893;
assign n159 = ~n826;
assign n1106 = n1575 & n652;
assign n1201 = n773 | n256;
assign n1101 = ~(n539 | n1586);
assign n611 = n84;
assign n279 = n1205 | n882;
assign n1380 = n186 | n882;
assign n1579 = n383 | n1635;
assign n846 = ~n1182;
assign n1522 = ~n565;
assign n762 = n1271 | n1101;
assign n616 = n894 & n600;
assign n1450 = n1796 | n677;
assign n1132 = n1257 | n806;
assign n1195 = ~(n1342 | n1013);
assign n781 = ~n1729;
assign n1749 = ~n507;
assign n1400 = ~(n579 | n783);
assign n1640 = n579 | n1218;
assign n550 = n508 | n6;
assign n1569 = n1659 & n1416;
assign n1218 = ~n1423;
assign n1779 = ~n1368;
assign n829 = ~n1021;
assign n1725 = ~(n377 | n115);
assign n1652 = n837 | n1653;
assign n13 = ~(n697 | n133);
assign n973 = n377 & n225;
assign n97 = n1701 | n628;
assign n690 = n1004 & n328;
assign n1609 = n1319 | n1554;
assign n614 = ~n807;
assign n723 = n1713 | n77;
assign n209 = n1016 & n1228;
assign n1448 = ~(n614 | n238);
assign n312 = n111 | n268;
assign n1538 = ~(n228 | n352);
assign n992 = ~n1100;
assign n458 = ~n363;
assign n293 = n1026 | n572;
assign n554 = ~(n44 | n175);
assign n1580 = ~(n395 | n591);
assign n1393 = ~(n1395 | n1304);
assign n1194 = ~n520;
assign n14 = ~(n717 ^ n507);
assign n706 = n981 & n1204;
assign n815 = ~(n377 | n3);
assign n1329 = ~(n795 ^ n294);
assign n660 = n627 | n905;
assign n1344 = n1665 | n1639;
assign n919 = ~(n428 ^ n1255);
assign n931 = n1295 | n510;
assign n1516 = ~(n535 | n925);
assign n1055 = n1365 | n125;
assign n1525 = ~(n539 | n729);
assign n287 = n971 & n600;
assign n26 = ~(n145 ^ n994);
assign n847 = ~n697;
assign n1560 = ~(n44 | n1242);
assign n141 = n307 | n456;
assign n394 = ~n1359;
assign n11 = ~(n539 | n1212);
assign n1155 = ~(n261 | n1640);
assign n162 = n846 | n579;
assign n1668 = ~n1130;
assign n1781 = ~(n261 | n1751);
assign n245 = n1613 & n1213;
assign n338 = n504 & n64;
assign n1612 = ~(n261 | n333);
assign n1783 = ~(n438 ^ n1696);
assign n1347 = ~n783;
assign n1535 = n1769 & n662;
assign n1751 = n579 | n829;
assign n1336 = n1043 & n1288;
assign n303 = n627 | n1631;
assign n1300 = ~(n819 | n329);
assign n178 = n307 | n882;
assign n1576 = n900 | n268;
assign n282 = n844 | n1200;
assign n864 = ~(n1162 | n1456);
assign n748 = ~n380;
assign n684 = n114 | n1232;
assign n889 = ~(n1793 ^ n1397);
assign n913 = n917 & n504;
assign n540 = ~(n347 | n127);
assign n1030 = n746 | n584;
assign n775 = n1264 | n268;
assign n742 = n1205 | n1495;
assign n1742 = ~(n1713 | n1288);
assign n1351 = ~(n44 | n633);
assign n1470 = ~(n703 ^ n396);
assign n336 = n186 | n456;
assign n1432 = ~n488;
assign n1487 = n1135 | n1168;
assign n1409 = n537 | n1427;
assign n1368 = ~(n216 ^ n1279);
assign n979 = n632 | n678;
assign n1754 = ~(n228 | n1693);
assign n220 = ~n1534;
assign n881 = n627 | n456;
assign n525 = ~(n901 ^ n1359);
assign n1411 = ~(n1357 & n1649);
assign n353 = ~(n468 ^ n207);
assign n248 = n424 & n13;
assign n71 = ~(n261 | n734);
assign n1241 = ~n205;
assign n433 = ~(n1395 | n1296);
assign n1702 = ~(n759 | n1354);
assign n1320 = n116 | n1560;
endmodule
