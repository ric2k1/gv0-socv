module top( 1_n1 , 1_n4 , 1_n5 , 1_n6 , 1_n11 , 1_n16 , 1_n19 , 1_n24 , 1_n35 , 1_n36 , 1_n39 , 1_n44 , 1_n45 , 1_n46 , 1_n48 , 1_n49 );
    input 1_n1 , 1_n4 , 1_n5 , 1_n11 , 1_n19 , 1_n24 , 1_n35 , 1_n39 , 1_n45 , 1_n46 , 1_n48 , 1_n49 ;
    output 1_n6 , 1_n16 , 1_n36 , 1_n44 ;
    wire 1_n0 , 1_n2 , 1_n3 , 1_n7 , 1_n8 , 1_n9 , 1_n10 , 1_n12 , 1_n13 , 1_n14 , 1_n15 , 1_n17 , 1_n18 , 1_n20 , 1_n21 , 1_n22 , 1_n23 , 1_n25 , 1_n26 , 1_n27 , 1_n28 , 1_n29 , 1_n30 , 1_n31 , 1_n32 , 1_n33 , 1_n34 , 1_n37 , 1_n38 , 1_n40 , 1_n41 , 1_n42 , 1_n43 , 1_n47 ;
assign 1_n38 = ~1_n11;
assign 1_n43 = ~(1_n47 ^ 1_n49);
assign 1_n10 = ~1_n30;
assign 1_n6 = ~(1_n7 ^ 1_n23);
assign 1_n34 = 1_n26 | 1_n8;
assign 1_n15 = ~(1_n20 | 1_n7);
assign 1_n27 = ~(1_n35 ^ 1_n48);
assign 1_n41 = ~(1_n5 ^ 1_n4);
assign 1_n14 = ~(1_n18 ^ 1_n3);
assign 1_n23 = ~(1_n14 ^ 1_n19);
assign 1_n31 = ~(1_n24 ^ 1_n39);
assign 1_n13 = ~(1_n35 & 1_n48);
assign 1_n25 = ~(1_n0 ^ 1_n11);
assign 1_n28 = ~(1_n22 | 1_n18);
assign 1_n36 = ~(1_n31 ^ 1_n46);
assign 1_n18 = 1_n32 & 1_n13;
assign 1_n8 = ~1_n39;
assign 1_n30 = 1_n21 & 1_n46;
assign 1_n22 = ~(1_n45 | 1_n1);
assign 1_n0 = ~(1_n34 ^ 1_n27);
assign 1_n9 = ~(1_n35 | 1_n48);
assign 1_n3 = ~(1_n45 ^ 1_n1);
assign 1_n12 = 1_n38 | 1_n10;
assign 1_n7 = 1_n2 & 1_n12;
assign 1_n20 = 1_n14 & 1_n29;
assign 1_n21 = ~1_n31;
assign 1_n17 = 1_n40 | 1_n15;
assign 1_n2 = 1_n0 | 1_n37;
assign 1_n32 = 1_n9 | 1_n34;
assign 1_n42 = ~(1_n41 ^ 1_n17);
assign 1_n16 = ~(1_n43 ^ 1_n42);
assign 1_n33 = 1_n1 & 1_n45;
assign 1_n37 = ~(1_n11 | 1_n30);
assign 1_n44 = ~(1_n10 ^ 1_n25);
assign 1_n26 = ~1_n24;
assign 1_n29 = ~1_n19;
assign 1_n40 = ~(1_n29 | 1_n14);
assign 1_n47 = 1_n33 | 1_n28;
endmodule
