module top( n1 , n3 , n4 , n15 , n21 , n23 , n28 , n32 , n37 , n38 , n40 , n45 , n47 , n50 , n52 , n53 , n54 , n60 , n72 , n75 , n79 , n81 , n83 , n86 , n87 , n91 , n95 , n97 , n99 , n105 , n111 , n114 , n117 , n122 , n139 , n152 , n154 , n155 , n160 , n162 , n168 , n176 , n183 , n185 , n187 , n191 , n194 , n197 , n198 , n200 , n205 , n206 , n208 , n211 , n214 , n215 , n218 , n220 , n227 , n228 , n231 , n242 , n243 , n248 , n254 , n262 , n265 , n269 , n273 , n276 , n278 , n280 , n283 );
    input n1 , n4 , n15 , n21 , n23 , n28 , n37 , n38 , n45 , n52 , n53 , n60 , n75 , n79 , n83 , n87 , n95 , n105 , n114 , n117 , n122 , n152 , n155 , n160 , n162 , n168 , n183 , n187 , n194 , n198 , n206 , n215 , n218 , n227 , n228 , n231 , n242 , n269 , n276 , n278 , n280 ;
    output n3 , n32 , n40 , n47 , n50 , n54 , n72 , n81 , n86 , n91 , n97 , n99 , n111 , n139 , n154 , n176 , n185 , n191 , n197 , n200 , n205 , n208 , n211 , n214 , n220 , n243 , n248 , n254 , n262 , n265 , n273 , n283 ;
    wire n0 , n2 , n5 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n16 , n17 , n18 , n19 , n20 , n22 , n24 , n25 , n26 , n27 , n29 , n30 , n31 , n33 , n34 , n35 , n36 , n39 , n41 , n42 , n43 , n44 , n46 , n48 , n49 , n51 , n55 , n56 , n57 , n58 , n59 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n73 , n74 , n76 , n77 , n78 , n80 , n82 , n84 , n85 , n88 , n89 , n90 , n92 , n93 , n94 , n96 , n98 , n100 , n101 , n102 , n103 , n104 , n106 , n107 , n108 , n109 , n110 , n112 , n113 , n115 , n116 , n118 , n119 , n120 , n121 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n153 , n156 , n157 , n158 , n159 , n161 , n163 , n164 , n165 , n166 , n167 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n177 , n178 , n179 , n180 , n181 , n182 , n184 , n186 , n188 , n189 , n190 , n192 , n193 , n195 , n196 , n199 , n201 , n202 , n203 , n204 , n207 , n209 , n210 , n212 , n213 , n216 , n217 , n219 , n221 , n222 , n223 , n224 , n225 , n226 , n229 , n230 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n244 , n245 , n246 , n247 , n249 , n250 , n251 , n252 , n253 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n263 , n264 , n266 , n267 , n268 , n270 , n271 , n272 , n274 , n275 , n277 , n279 , n281 , n282 , n284 , n285 ;
assign n140 = n247 & n201;
assign n72 = ~(n126 ^ n162);
assign n244 = n173 | n230;
assign n18 = n141 | n136;
assign n43 = ~n4;
assign n177 = ~n198;
assign n16 = ~(n215 ^ n206);
assign n80 = n237 | n252;
assign n81 = ~(n216 ^ n194);
assign n261 = ~n193;
assign n55 = ~n172;
assign n148 = ~n168;
assign n136 = ~(n209 ^ n77);
assign n263 = ~(n206 ^ n183);
assign n257 = ~(n280 ^ n21);
assign n159 = ~(n285 ^ n24);
assign n254 = n0 ^ n28;
assign n33 = n115 | n256;
assign n110 = n55 | n18;
assign n68 = ~(n227 ^ n21);
assign n181 = ~(n187 ^ n45);
assign n49 = ~n26;
assign n126 = n90 | n235;
assign n225 = ~n12;
assign n202 = n103 | n235;
assign n200 = ~(n186 ^ n23);
assign n30 = n78 | n101;
assign n123 = ~n137;
assign n281 = n193 | n169;
assign n50 = ~(n179 ^ n87);
assign n164 = ~(n28 ^ n15);
assign n47 = n272 ^ n38;
assign n137 = ~n35;
assign n27 = n142 | n5;
assign n175 = ~n128;
assign n277 = n223 | n108;
assign n149 = n2 & n240;
assign n213 = ~(n89 ^ n165);
assign n66 = ~n275;
assign n103 = ~n224;
assign n190 = n226 | n281;
assign n115 = ~n224;
assign n42 = n137 | n222;
assign n56 = ~n114;
assign n283 = ~(n48 ^ n105);
assign n259 = n59 | n43;
assign n48 = n195 | n157;
assign n11 = ~n199;
assign n104 = n7 | n232;
assign n209 = ~(n170 ^ n188);
assign n78 = ~n250;
assign n174 = n55 | n150;
assign n239 = ~n2;
assign n176 = ~(n33 ^ n95);
assign n17 = n173 | n235;
assign n219 = ~(n112 ^ n16);
assign n249 = ~n60;
assign n40 = ~(n147 ^ n183);
assign n134 = n203 | n43;
assign n274 = n65 & n239;
assign n41 = n107 | n266;
assign n236 = ~(n228 ^ n95);
assign n77 = ~(n279 ^ n258);
assign n119 = n49 | n88;
assign n74 = ~(n278 ^ n52);
assign n270 = n161 & n7;
assign n163 = n78 | n19;
assign n100 = ~(n82 ^ n74);
assign n284 = ~(n271 ^ n20);
assign n241 = ~(n75 ^ n45);
assign n131 = n249 | n127;
assign n97 = ~(n27 ^ n53);
assign n94 = ~(n138 ^ n212);
assign n54 = ~(n124 ^ n160);
assign n224 = ~n104;
assign n237 = ~n149;
assign n31 = ~(n152 ^ n280);
assign n203 = ~n218;
assign n165 = ~(n152 ^ n227);
assign n129 = ~(n237 | n190);
assign n193 = ~(n71 ^ n62);
assign n166 = ~n26;
assign n256 = ~n247;
assign n107 = ~n136;
assign n144 = n166 | n163;
assign n2 = ~(n245 ^ n217);
assign n240 = ~n65;
assign n153 = ~(n276 ^ n95);
assign n111 = ~(n264 ^ n83);
assign n268 = n173 | n36;
assign n29 = ~(n28 ^ n1);
assign n125 = ~(n8 ^ n31);
assign n51 = n180 | n196;
assign n272 = ~(n182 | n190);
assign n19 = n121 | n260;
assign n141 = ~n266;
assign n118 = ~n210;
assign n5 = n252 | n275;
assign n212 = ~(n23 ^ n83);
assign n179 = n115 | n230;
assign n88 = n174 | n196;
assign n245 = ~(n9 ^ n68);
assign n91 = ~(n119 ^ n152);
assign n92 = n26 & n46;
assign n71 = ~(n8 ^ n178);
assign n26 = n6 & n35;
assign n82 = ~(n242 ^ n87);
assign n143 = n226 | n36;
assign n20 = ~(n219 ^ n134);
assign n170 = ~(n167 ^ n257);
assign n196 = n261 | n96;
assign n169 = n192 | n123;
assign n7 = ~n225;
assign n172 = ~n58;
assign n204 = ~(n135 ^ n73);
assign n246 = n169 | n19;
assign n161 = ~n41;
assign n147 = n260 | n143;
assign n69 = ~n210;
assign n138 = ~(n53 ^ n155);
assign n130 = n103 | n282;
assign n265 = n238 ^ n79;
assign n262 = n129 ^ n1;
assign n90 = ~n270;
assign n3 = ~(n130 ^ n278);
assign n22 = ~(n100 ^ n263);
assign n234 = ~(n83 ^ n52);
assign n145 = n275 | n19;
assign n208 = ~(n63 ^ n52);
assign n184 = n177 | n108;
assign n73 = n148 | n127;
assign n207 = ~(n105 ^ n194);
assign n98 = ~(n1 ^ n38);
assign n135 = ~(n153 ^ n102);
assign n217 = ~(n234 ^ n76);
assign n85 = ~(n162 ^ n183);
assign n93 = n180 | n101;
assign n112 = ~(n122 ^ n187);
assign n267 = n69 | n80;
assign n157 = n128 | n174;
assign n106 = n56 | n221;
assign n271 = ~(n23 ^ n278);
assign n199 = n92 & n149;
assign n84 = n173 | n80;
assign n142 = ~n158;
assign n61 = n222 | n123;
assign n191 = ~(n133 ^ n215);
assign n101 = ~n92;
assign n158 = ~n233;
assign n243 = ~(n202 ^ n45);
assign n222 = ~n192;
assign n235 = n182 | n128;
assign n279 = ~(n79 ^ n276);
assign n230 = n142 | n281;
assign n201 = ~n110;
assign n12 = ~(n116 ^ n151);
assign n156 = ~n231;
assign n260 = ~n274;
assign n180 = ~n66;
assign n24 = ~(n9 ^ n277);
assign n197 = ~(n44 ^ n242);
assign n39 = ~(n170 ^ n259);
assign n57 = ~(n98 ^ n39);
assign n109 = ~(n213 ^ n184);
assign n133 = n90 | n80;
assign n25 = n156 | n221;
assign n238 = n199 & n201;
assign n250 = ~n174;
assign n8 = ~(n13 ^ n29);
assign n89 = ~(n105 ^ n160);
assign n275 = n12 | n41;
assign n96 = ~n149;
assign n178 = ~(n160 ^ n37);
assign n285 = ~(n53 ^ n242);
assign n233 = n240 | n239;
assign n9 = ~(n241 ^ n85);
assign n210 = ~n104;
assign n70 = ~n233;
assign n221 = ~n4;
assign n132 = n118 | n11;
assign n226 = n58 | n232;
assign n58 = ~n12;
assign n151 = ~(n236 ^ n10);
assign n128 = n121 | n42;
assign n186 = n166 | n51;
assign n59 = ~n269;
assign n86 = ~(n244 ^ n37);
assign n171 = ~(n155 ^ n87);
assign n62 = ~(n171 ^ n204);
assign n6 = ~(n146 ^ n159);
assign n223 = ~n117;
assign n264 = n49 | n145;
assign n113 = ~(n215 ^ n162);
assign n167 = ~(n194 ^ n37);
assign n127 = ~n4;
assign n258 = ~(n213 ^ n131);
assign n13 = ~(n79 ^ n228);
assign n108 = ~n4;
assign n139 = n189 ^ n155;
assign n220 = ~(n144 ^ n227);
assign n44 = n195 | n251;
assign n65 = ~(n125 ^ n284);
assign n247 = n92 & n274;
assign n102 = ~(n15 ^ n38);
assign n252 = ~n175;
assign n255 = ~(n94 ^ n113);
assign n150 = n136 | n266;
assign n229 = ~n70;
assign n0 = n199 & n270;
assign n182 = ~n274;
assign n67 = ~(n164 ^ n109);
assign n173 = n110;
assign n214 = ~(n267 ^ n187);
assign n121 = ~n34;
assign n188 = ~(n122 ^ n75);
assign n116 = ~(n100 ^ n181);
assign n216 = n229 | n268;
assign n14 = n173 | n282;
assign n192 = ~n6;
assign n146 = ~(n219 ^ n207);
assign n36 = n261 | n61;
assign n154 = ~(n64 ^ n206);
assign n120 = n247 & n270;
assign n32 = ~(n132 ^ n228);
assign n189 = ~(n233 | n93);
assign n205 = ~(n253 ^ n21);
assign n266 = ~(n255 ^ n67);
assign n35 = ~(n22 ^ n57);
assign n185 = n140 ^ n276;
assign n211 = ~(n84 ^ n122);
assign n46 = ~n193;
assign n64 = n96 | n143;
assign n253 = n173 | n246;
assign n195 = ~n158;
assign n34 = ~n46;
assign n124 = n229 | n30;
assign n232 = n107 | n141;
assign n10 = ~(n94 ^ n106);
assign n63 = n69 | n246;
assign n273 = ~(n17 ^ n75);
assign n251 = n36 | n118;
assign n248 = n120 ^ n15;
assign n76 = ~(n135 ^ n25);
assign n282 = n169 | n196;
assign n99 = ~(n14 ^ n280);
endmodule
