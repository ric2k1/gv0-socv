module top( n5 , n13 , n17 , n20 , n27 , n36 , n37 , n53 , n62 , 
n75 , n80 , n86 , n93 , n105 , n106 , n111 , n117 , n139 , n145 , 
n147 , n157 , n161 , n175 , n176 , n182 , n190 , n198 , n204 , n208 , 
n214 , n217 , n219 , n224 , n225 , n226 , n229 , n235 , n241 , n244 , 
n249 , n256 , n281 , n287 , n289 , n294 , n300 , n303 , n319 , n345 , 
n346 , n364 , n365 , n368 , n384 , n387 , n389 , n393 , n403 , n409 , 
n410 , n417 , n430 , n439 , n442 , n457 , n465 , n473 , n477 , n489 , 
n491 , n493 , n503 , n506 , n511 , n515 , n518 , n521 , n532 , n537 , 
n587 , n588 , n593 , n594 , n595 , n606 , n618 , n630 , n642 , n648 , 
n656 , n671 , n680 , n684 , n690 , n691 , n693 , n699 , n702 , n703 , 
n704 , n706 , n716 , n741 , n742 , n743 , n746 , n753 , n756 , n765 , 
n777 , n782 , n788 );
    input n5 , n13 , n17 , n20 , n36 , n37 , n53 , n75 , n80 , 
n86 , n93 , n105 , n106 , n111 , n117 , n139 , n147 , n157 , n161 , 
n182 , n190 , n198 , n204 , n208 , n214 , n217 , n219 , n224 , n226 , 
n229 , n235 , n244 , n249 , n281 , n287 , n289 , n300 , n303 , n319 , 
n346 , n364 , n365 , n368 , n384 , n393 , n403 , n409 , n410 , n417 , 
n439 , n457 , n465 , n473 , n477 , n503 , n506 , n511 , n518 , n521 , 
n532 , n537 , n587 , n588 , n593 , n594 , n595 , n606 , n642 , n648 , 
n656 , n671 , n680 , n684 , n690 , n693 , n699 , n702 , n706 , n716 , 
n741 , n742 , n743 , n746 , n777 , n782 , n788 ;
    output n27 , n62 , n145 , n175 , n176 , n225 , n241 , n256 , n294 , 
n345 , n387 , n389 , n430 , n442 , n489 , n491 , n493 , n515 , n618 , 
n630 , n691 , n703 , n704 , n753 , n756 , n765 ;
    wire n0 , n1 , n2 , n3 , n4 , n6 , n7 , n8 , n9 , 
n10 , n11 , n12 , n14 , n15 , n16 , n18 , n19 , n21 , n22 , 
n23 , n24 , n25 , n26 , n28 , n29 , n30 , n31 , n32 , n33 , 
n34 , n35 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , 
n46 , n47 , n48 , n49 , n50 , n51 , n52 , n54 , n55 , n56 , 
n57 , n58 , n59 , n60 , n61 , n63 , n64 , n65 , n66 , n67 , 
n68 , n69 , n70 , n71 , n72 , n73 , n74 , n76 , n77 , n78 , 
n79 , n81 , n82 , n83 , n84 , n85 , n87 , n88 , n89 , n90 , 
n91 , n92 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , 
n102 , n103 , n104 , n107 , n108 , n109 , n110 , n112 , n113 , n114 , 
n115 , n116 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , 
n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , 
n136 , n137 , n138 , n140 , n141 , n142 , n143 , n144 , n146 , n148 , 
n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n158 , n159 , 
n160 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , 
n171 , n172 , n173 , n174 , n177 , n178 , n179 , n180 , n181 , n183 , 
n184 , n185 , n186 , n187 , n188 , n189 , n191 , n192 , n193 , n194 , 
n195 , n196 , n197 , n199 , n200 , n201 , n202 , n203 , n205 , n206 , 
n207 , n209 , n210 , n211 , n212 , n213 , n215 , n216 , n218 , n220 , 
n221 , n222 , n223 , n227 , n228 , n230 , n231 , n232 , n233 , n234 , 
n236 , n237 , n238 , n239 , n240 , n242 , n243 , n245 , n246 , n247 , 
n248 , n250 , n251 , n252 , n253 , n254 , n255 , n257 , n258 , n259 , 
n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , 
n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , 
n280 , n282 , n283 , n284 , n285 , n286 , n288 , n290 , n291 , n292 , 
n293 , n295 , n296 , n297 , n298 , n299 , n301 , n302 , n304 , n305 , 
n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , 
n316 , n317 , n318 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , 
n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , 
n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n347 , n348 , 
n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , 
n359 , n360 , n361 , n362 , n363 , n366 , n367 , n369 , n370 , n371 , 
n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , 
n382 , n383 , n385 , n386 , n388 , n390 , n391 , n392 , n394 , n395 , 
n396 , n397 , n398 , n399 , n400 , n401 , n402 , n404 , n405 , n406 , 
n407 , n408 , n411 , n412 , n413 , n414 , n415 , n416 , n418 , n419 , 
n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , 
n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n440 , n441 , 
n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , 
n453 , n454 , n455 , n456 , n458 , n459 , n460 , n461 , n462 , n463 , 
n464 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n474 , n475 , 
n476 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , 
n487 , n488 , n490 , n492 , n494 , n495 , n496 , n497 , n498 , n499 , 
n500 , n501 , n502 , n504 , n505 , n507 , n508 , n509 , n510 , n512 , 
n513 , n514 , n516 , n517 , n519 , n520 , n522 , n523 , n524 , n525 , 
n526 , n527 , n528 , n529 , n530 , n531 , n533 , n534 , n535 , n536 , 
n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , 
n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , 
n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , 
n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , 
n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n589 , 
n590 , n591 , n592 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , 
n603 , n604 , n605 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , 
n614 , n615 , n616 , n617 , n619 , n620 , n621 , n622 , n623 , n624 , 
n625 , n626 , n627 , n628 , n629 , n631 , n632 , n633 , n634 , n635 , 
n636 , n637 , n638 , n639 , n640 , n641 , n643 , n644 , n645 , n646 , 
n647 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n657 , n658 , 
n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , 
n669 , n670 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , 
n681 , n682 , n683 , n685 , n686 , n687 , n688 , n689 , n692 , n694 , 
n695 , n696 , n697 , n698 , n700 , n701 , n705 , n707 , n708 , n709 , 
n710 , n711 , n712 , n713 , n714 , n715 , n717 , n718 , n719 , n720 , 
n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , 
n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , 
n744 , n745 , n747 , n748 , n749 , n750 , n751 , n752 , n754 , n755 , 
n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n766 , n767 , 
n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n778 , 
n779 , n780 , n781 , n783 , n784 , n785 , n786 , n787 , n789 ;
    or g0 ( n8 , n559 , n136 );
    and g1 ( n676 , n578 , n778 );
    nor g2 ( n683 , n403 , n783 );
    or g3 ( n213 , n293 , n774 );
    nor g4 ( n273 , n300 , n250 );
    nor g5 ( n34 , n196 , n40 );
    and g6 ( n109 , n787 , n405 );
    and g7 ( n122 , n114 , n600 );
    nor g8 ( n645 , n452 , n488 );
    or g9 ( n621 , n433 , n106 );
    or g10 ( n312 , n381 , n296 );
    not g11 ( n534 , n226 );
    or g12 ( n657 , n341 , n59 );
    nor g13 ( n6 , n393 , n447 );
    not g14 ( n778 , n268 );
    or g15 ( n673 , n717 , n737 );
    and g16 ( n634 , n692 , n597 );
    nor g17 ( n719 , n452 , n655 );
    xnor g18 ( n644 , n475 , n716 );
    nor g19 ( n323 , n648 , n223 );
    not g20 ( n646 , n5 );
    and g21 ( n369 , n46 , n230 );
    not g22 ( n681 , n521 );
    and g23 ( n411 , n760 , n88 );
    nor g24 ( n600 , n656 , n155 );
    nor g25 ( n698 , n452 , n552 );
    and g26 ( n774 , n656 , n695 );
    xnor g27 ( n311 , n751 , n680 );
    or g28 ( n586 , n391 , n652 );
    or g29 ( n206 , n165 , n153 );
    not g30 ( n760 , n202 );
    not g31 ( n628 , n157 );
    and g32 ( n91 , n165 , n153 );
    or g33 ( n493 , n309 , n12 );
    or g34 ( n203 , n38 , n697 );
    or g35 ( n375 , n686 , n772 );
    or g36 ( n288 , n150 , n598 );
    and g37 ( n268 , n522 , n443 );
    or g38 ( n31 , n459 , n656 );
    nor g39 ( n415 , n98 , n363 );
    or g40 ( n685 , n546 , n276 );
    and g41 ( n63 , n131 , n627 );
    and g42 ( n764 , n656 , n135 );
    or g43 ( n707 , n452 , n761 );
    and g44 ( n450 , n666 , n257 );
    and g45 ( n52 , n391 , n767 );
    or g46 ( n772 , n452 , n270 );
    nor g47 ( n252 , n166 , n189 );
    and g48 ( n466 , n75 , n452 );
    not g49 ( n399 , n603 );
    and g50 ( n16 , n42 , n29 );
    nor g51 ( n207 , n537 , n212 );
    and g52 ( n277 , n581 , n248 );
    not g53 ( n407 , n749 );
    or g54 ( n574 , n607 , n264 );
    not g55 ( n383 , n520 );
    not g56 ( n169 , n236 );
    or g57 ( n97 , n537 , n300 );
    not g58 ( n559 , n393 );
    xnor g59 ( n14 , n440 , n19 );
    nor g60 ( n762 , n484 , n635 );
    nor g61 ( n589 , n656 , n568 );
    or g62 ( n462 , n42 , n29 );
    nor g63 ( n110 , n403 , n590 );
    or g64 ( n258 , n331 , n121 );
    and g65 ( n257 , n546 , n757 );
    or g66 ( n639 , n16 , n752 );
    not g67 ( n661 , n351 );
    not g68 ( n127 , n106 );
    xnor g69 ( n655 , n749 , n163 );
    nor g70 ( n48 , n656 , n674 );
    nor g71 ( n678 , n417 , n550 );
    not g72 ( n381 , n439 );
    xnor g73 ( n65 , n582 , n788 );
    and g74 ( n153 , n609 , n81 );
    xnor g75 ( n615 , n409 , n642 );
    not g76 ( n264 , n584 );
    not g77 ( n452 , n656 );
    xnor g78 ( n177 , n643 , n780 );
    or g79 ( n200 , n728 , n694 );
    and g80 ( n42 , n591 , n288 );
    and g81 ( n173 , n330 , n599 );
    nor g82 ( n533 , n452 , n676 );
    nor g83 ( n269 , n439 , n117 );
    or g84 ( n233 , n559 , n779 );
    not g85 ( n167 , n300 );
    xnor g86 ( n552 , n228 , n487 );
    or g87 ( n76 , n766 , n158 );
    not g88 ( n664 , n642 );
    or g89 ( n471 , n559 , n436 );
    not g90 ( n186 , n713 );
    or g91 ( n456 , n300 , n106 );
    nor g92 ( n604 , n656 , n3 );
    and g93 ( n557 , n37 , n501 );
    or g94 ( n643 , n460 , n7 );
    nor g95 ( n56 , n656 , n140 );
    not g96 ( n688 , n700 );
    not g97 ( n519 , n17 );
    and g98 ( n199 , n362 , n397 );
    not g99 ( n602 , n786 );
    or g100 ( n251 , n127 , n74 );
    and g101 ( n766 , n503 , n182 );
    not g102 ( n126 , n657 );
    and g103 ( n185 , n660 , n441 );
    or g104 ( n755 , n202 , n560 );
    nor g105 ( n154 , n384 , n129 );
    nor g106 ( n133 , n693 , n17 );
    and g107 ( n659 , n746 , n127 );
    and g108 ( n163 , n152 , n596 );
    and g109 ( n274 , n656 , n776 );
    nor g110 ( n733 , n214 , n69 );
    nor g111 ( n514 , n355 , n536 );
    and g112 ( n77 , n656 , n71 );
    nor g113 ( n336 , n228 , n372 );
    nor g114 ( n115 , n452 , n544 );
    or g115 ( n376 , n656 , n563 );
    not g116 ( n222 , n148 );
    or g117 ( n597 , n393 , n454 );
    or g118 ( n360 , n356 , n299 );
    or g119 ( n228 , n535 , n274 );
    not g120 ( n391 , n680 );
    or g121 ( n636 , n626 , n641 );
    or g122 ( n350 , n458 , n613 );
    nor g123 ( n170 , n649 , n376 );
    nor g124 ( n461 , n350 , n0 );
    and g125 ( n181 , n595 , n452 );
    xor g126 ( n526 , n767 , n453 );
    or g127 ( n316 , n393 , n508 );
    xnor g128 ( n516 , n439 , n742 );
    nor g129 ( n686 , n513 , n28 );
    and g130 ( n50 , n218 , n396 );
    and g131 ( n168 , n656 , n444 );
    not g132 ( n480 , n592 );
    nor g133 ( n70 , n656 , n631 );
    not g134 ( n441 , n19 );
    or g135 ( n549 , n628 , n340 );
    and g136 ( n490 , n228 , n372 );
    and g137 ( n497 , n656 , n408 );
    and g138 ( n267 , n403 , n311 );
    or g139 ( n174 , n23 , n520 );
    not g140 ( n581 , n159 );
    or g141 ( n30 , n519 , n423 );
    and g142 ( n143 , n366 , n369 );
    nor g143 ( n502 , n705 , n251 );
    or g144 ( n582 , n125 , n353 );
    and g145 ( n380 , n462 , n639 );
    nor g146 ( n529 , n656 , n388 );
    or g147 ( n736 , n621 , n553 );
    nor g148 ( n540 , n759 , n246 );
    and g149 ( n607 , n690 , n217 );
    or g150 ( n58 , n687 , n148 );
    xnor g151 ( n404 , n189 , n61 );
    or g152 ( n618 , n589 , n576 );
    nor g153 ( n763 , n300 , n789 );
    or g154 ( n753 , n47 , n395 );
    and g155 ( n561 , n547 , n260 );
    nor g156 ( n102 , n452 , n385 );
    not g157 ( n29 , n68 );
    nor g158 ( n39 , n452 , n33 );
    not g159 ( n292 , n287 );
    nor g160 ( n573 , n440 , n441 );
    not g161 ( n354 , n330 );
    or g162 ( n262 , n525 , n524 );
    nor g163 ( n197 , n157 , n303 );
    and g164 ( n332 , n174 , n509 );
    or g165 ( n396 , n549 , n374 );
    or g166 ( n114 , n297 , n60 );
    xnor g167 ( n520 , n574 , n690 );
    nor g168 ( n339 , n527 , n667 );
    nor g169 ( n25 , n537 , n286 );
    nor g170 ( n494 , n724 , n35 );
    and g171 ( n592 , n506 , n169 );
    nor g172 ( n155 , n495 , n556 );
    or g173 ( n241 , n731 , n698 );
    xnor g174 ( n130 , n76 , n777 );
    and g175 ( n270 , n513 , n28 );
    and g176 ( n221 , n518 , n452 );
    and g177 ( n717 , n352 , n516 );
    nor g178 ( n507 , n726 , n193 );
    or g179 ( n726 , n754 , n497 );
    and g180 ( n230 , n608 , n237 );
    xnor g181 ( n385 , n213 , n230 );
    xnor g182 ( n555 , n17 , n13 );
    not g183 ( n340 , n303 );
    or g184 ( n756 , n386 , n172 );
    and g185 ( n560 , n688 , n314 );
    nor g186 ( n98 , n78 , n470 );
    and g187 ( n322 , n656 , n344 );
    or g188 ( n697 , n403 , n537 );
    or g189 ( n565 , n73 , n446 );
    nor g190 ( n119 , n787 , n405 );
    or g191 ( n663 , n735 , n200 );
    nor g192 ( n370 , n185 , n727 );
    or g193 ( n256 , n160 , n321 );
    or g194 ( n749 , n632 , n476 );
    not g195 ( n694 , n76 );
    or g196 ( n327 , n127 , n714 );
    not g197 ( n735 , n281 );
    nor g198 ( n486 , n452 , n432 );
    not g199 ( n132 , n200 );
    not g200 ( n296 , n742 );
    not g201 ( n525 , n648 );
    nor g202 ( n499 , n300 , n485 );
    or g203 ( n227 , n15 , n668 );
    xnor g204 ( n695 , n236 , n506 );
    and g205 ( n725 , n373 , n101 );
    not g206 ( n331 , n417 );
    and g207 ( n438 , n368 , n452 );
    not g208 ( n547 , n549 );
    or g209 ( n400 , n292 , n656 );
    xnor g210 ( n246 , n355 , n141 );
    or g211 ( n701 , n660 , n19 );
    or g212 ( n189 , n32 , n658 );
    and g213 ( n476 , n656 , n770 );
    or g214 ( n583 , n44 , n380 );
    not g215 ( n566 , n636 );
    or g216 ( n131 , n412 , n787 );
    not g217 ( n530 , n299 );
    not g218 ( n687 , n672 );
    and g219 ( n789 , n137 , n327 );
    or g220 ( n239 , n608 , n636 );
    and g221 ( n348 , n20 , n57 );
    or g222 ( n669 , n666 , n685 );
    not g223 ( n46 , n213 );
    and g224 ( n341 , n161 , n452 );
    nor g225 ( n286 , n313 , n763 );
    xnor g226 ( n108 , n350 , n369 );
    and g227 ( n771 , n78 , n470 );
    or g228 ( n430 , n494 , n307 );
    or g229 ( n609 , n688 , n164 );
    or g230 ( n148 , n407 , n232 );
    xnor g231 ( n775 , n5 , n157 );
    or g232 ( n692 , n559 , n418 );
    and g233 ( n32 , n439 , n117 );
    xnor g234 ( n263 , n258 , n20 );
    nor g235 ( n454 , n358 , n482 );
    not g236 ( n479 , n606 );
    not g237 ( n255 , n490 );
    or g238 ( n62 , n604 , n87 );
    or g239 ( n489 , n56 , n102 );
    or g240 ( n142 , n559 , n722 );
    and g241 ( n193 , n687 , n392 );
    nor g242 ( n548 , n759 , n615 );
    nor g243 ( n278 , n64 , n625 );
    or g244 ( n470 , n495 , n778 );
    and g245 ( n202 , n700 , n164 );
    and g246 ( n55 , n244 , n452 );
    and g247 ( n469 , n656 , n65 );
    or g248 ( n247 , n547 , n197 );
    nor g249 ( n144 , n656 , n496 );
    or g250 ( n553 , n272 , n97 );
    and g251 ( n750 , n24 , n193 );
    and g252 ( n329 , n532 , n452 );
    and g253 ( n632 , n743 , n452 );
    and g254 ( n611 , n715 , n623 );
    and g255 ( n220 , n702 , n452 );
    xnor g256 ( n405 , n184 , n422 );
    not g257 ( n759 , n537 );
    or g258 ( n343 , n116 , n603 );
    xnor g259 ( n483 , n159 , n248 );
    or g260 ( n345 , n144 , n696 );
    and g261 ( n712 , n14 , n173 );
    or g262 ( n95 , n429 , n539 );
    not g263 ( n183 , n706 );
    and g264 ( n458 , n224 , n452 );
    nor g265 ( n783 , n577 , n207 );
    or g266 ( n603 , n24 , n58 );
    not g267 ( n758 , n384 );
    nor g268 ( n211 , n94 , n169 );
    not g269 ( n652 , n594 );
    or g270 ( n382 , n455 , n747 );
    nor g271 ( n569 , n452 , n10 );
    and g272 ( n429 , n235 , n452 );
    or g273 ( n721 , n46 , n239 );
    nor g274 ( n242 , n540 , n191 );
    and g275 ( n492 , n300 , n404 );
    xnor g276 ( n445 , n439 , n117 );
    xnor g277 ( n435 , n700 , n314 );
    and g278 ( n640 , n412 , n787 );
    or g279 ( n41 , n662 , n480 );
    and g280 ( n402 , n400 , n375 );
    nor g281 ( n201 , n377 , n647 );
    nor g282 ( n421 , n284 , n380 );
    and g283 ( n724 , n617 , n638 );
    and g284 ( n428 , n184 , n240 );
    xnor g285 ( n413 , n349 , n445 );
    or g286 ( n243 , n452 , n379 );
    not g287 ( n660 , n440 );
    or g288 ( n424 , n620 , n178 );
    not g289 ( n146 , n190 );
    or g290 ( n704 , n624 , n533 );
    or g291 ( n362 , n472 , n335 );
    nor g292 ( n158 , n720 , n28 );
    not g293 ( n614 , n582 );
    xnor g294 ( n123 , n217 , n365 );
    nor g295 ( n770 , n154 , n661 );
    not g296 ( n718 , n663 );
    and g297 ( n576 , n206 , n134 );
    not g298 ( n527 , n382 );
    nor g299 ( n45 , n298 , n718 );
    not g300 ( n24 , n726 );
    nor g301 ( n658 , n349 , n269 );
    or g302 ( n769 , n610 , n650 );
    not g303 ( n113 , n685 );
    and g304 ( n28 , n586 , n781 );
    nor g305 ( n1 , n452 , n177 );
    or g306 ( n596 , n185 , n173 );
    nor g307 ( n196 , n741 , n713 );
    or g308 ( n440 , n221 , n261 );
    nor g309 ( n408 , n323 , n390 );
    nor g310 ( n612 , n36 , n348 );
    and g311 ( n460 , n587 , n452 );
    nor g312 ( n482 , n403 , n242 );
    not g313 ( n103 , n669 );
    and g314 ( n238 , n249 , n439 );
    not g315 ( n394 , n564 );
    not g316 ( n558 , n214 );
    and g317 ( n500 , n120 , n748 );
    or g318 ( n578 , n522 , n443 );
    or g319 ( n156 , n336 , n490 );
    not g320 ( n554 , n741 );
    nor g321 ( n416 , n367 , n171 );
    not g322 ( n0 , n721 );
    or g323 ( n101 , n478 , n290 );
    not g324 ( n727 , n152 );
    and g325 ( n314 , n481 , n85 );
    and g326 ( n129 , n699 , n718 );
    and g327 ( n512 , n364 , n452 );
    nor g328 ( n508 , n267 , n110 );
    xnor g329 ( n317 , n619 , n503 );
    nor g330 ( n149 , n656 , n538 );
    not g331 ( n23 , n503 );
    nor g332 ( n682 , n700 , n314 );
    xnor g333 ( n544 , n505 , n257 );
    or g334 ( n635 , n656 , n2 );
    nor g335 ( n517 , n359 , n128 );
    and g336 ( n780 , n179 , n487 );
    or g337 ( n89 , n628 , n739 );
    or g338 ( n225 , n271 , n531 );
    or g339 ( n351 , n758 , n320 );
    not g340 ( n356 , n245 );
    nor g341 ( n309 , n461 , n670 );
    or g342 ( n218 , n646 , n107 );
    not g343 ( n231 , n402 );
    not g344 ( n412 , n184 );
    not g345 ( n324 , n69 );
    xnor g346 ( n371 , n657 , n567 );
    and g347 ( n732 , n537 , n304 );
    and g348 ( n359 , n473 , n127 );
    and g349 ( n484 , n435 , n285 );
    xnor g350 ( n54 , n495 , n268 );
    xnor g351 ( n118 , n749 , n49 );
    or g352 ( n605 , n428 , n580 );
    and g353 ( n487 , n116 , n750 );
    or g354 ( n398 , n416 , n113 );
    nor g355 ( n357 , n334 , n354 );
    and g356 ( n740 , n157 , n393 );
    and g357 ( n84 , n343 , n529 );
    nor g358 ( n307 , n452 , n26 );
    or g359 ( n786 , n558 , n324 );
    nor g360 ( n776 , n678 , n57 );
    not g361 ( n297 , n495 );
    and g362 ( n443 , n356 , n143 );
    nor g363 ( n590 , n732 , n572 );
    and g364 ( n510 , n229 , n452 );
    xor g365 ( n260 , n5 , n671 );
    nor g366 ( n531 , n452 , n679 );
    and g367 ( n501 , n53 , n602 );
    and g368 ( n74 , n30 , n729 );
    and g369 ( n620 , n503 , n611 );
    or g370 ( n389 , n72 , n543 );
    nor g371 ( n321 , n452 , n483 );
    not g372 ( n768 , n240 );
    or g373 ( n22 , n55 , n708 );
    or g374 ( n236 , n681 , n4 );
    or g375 ( n378 , n14 , n173 );
    or g376 ( n349 , n664 , n479 );
    or g377 ( n495 , n310 , n83 );
    not g378 ( n641 , n446 );
    nor g379 ( n67 , n284 , n420 );
    nor g380 ( n172 , n452 , n371 );
    xnor g381 ( n432 , n629 , n755 );
    or g382 ( n81 , n682 , n21 );
    xnor g383 ( n474 , n78 , n114 );
    nor g384 ( n747 , n452 , n247 );
    and g385 ( n290 , n51 , n504 );
    nor g386 ( n209 , n672 , n222 );
    nor g387 ( n73 , n159 , n318 );
    xnor g388 ( n406 , n663 , n699 );
    xnor g389 ( n3 , n290 , n67 );
    and g390 ( n59 , n656 , n644 );
    or g391 ( n505 , n512 , n469 );
    xnor g392 ( n308 , n672 , n392 );
    nor g393 ( n444 , n612 , n614 );
    or g394 ( n35 , n656 , n11 );
    not g395 ( n546 , n367 );
    or g396 ( n737 , n127 , n315 );
    and g397 ( n386 , n419 , n434 );
    or g398 ( n330 , n472 , n677 );
    nor g399 ( n134 , n452 , n91 );
    not g400 ( n730 , n41 );
    nor g401 ( n773 , n452 , n130 );
    nor g402 ( n467 , n657 , n563 );
    nor g403 ( n622 , n452 , n712 );
    and g404 ( n223 , n457 , n661 );
    or g405 ( n591 , n183 , n656 );
    or g406 ( n691 , n9 , n415 );
    and g407 ( n302 , n42 , n68 );
    nor g408 ( n434 , n656 , n467 );
    or g409 ( n138 , n656 , n556 );
    or g410 ( n145 , n84 , n39 );
    xnor g411 ( n675 , n505 , n113 );
    not g412 ( n433 , n319 );
    not g413 ( n472 , n283 );
    not g414 ( n563 , n333 );
    or g415 ( n51 , n42 , n68 );
    or g416 ( n187 , n220 , n99 );
    or g417 ( n668 , n347 , n266 );
    xnor g418 ( n723 , n95 , n450 );
    and g419 ( n535 , n465 , n452 );
    nor g420 ( n9 , n656 , n474 );
    nor g421 ( n191 , n537 , n431 );
    or g422 ( n387 , n170 , n637 );
    or g423 ( n475 , n554 , n186 );
    xnor g424 ( n513 , n503 , n182 );
    not g425 ( n528 , n574 );
    nor g426 ( n192 , n167 , n413 );
    or g427 ( n667 , n740 , n295 );
    and g428 ( n250 , n90 , n673 );
    or g429 ( n66 , n534 , n656 );
    and g430 ( n305 , n522 , n360 );
    and g431 ( n100 , n785 , n424 );
    and g432 ( n585 , n656 , n45 );
    nor g433 ( n254 , n187 , n566 );
    or g434 ( n333 , n275 , n669 );
    xnor g435 ( n104 , n680 , n594 );
    xnor g436 ( n551 , n786 , n53 );
    and g437 ( n754 , n588 , n452 );
    or g438 ( n152 , n660 , n441 );
    and g439 ( n69 , n208 , n730 );
    not g440 ( n784 , n111 );
    nor g441 ( n447 , n403 , n18 );
    and g442 ( n64 , n693 , n17 );
    or g443 ( n781 , n280 , n50 );
    not g444 ( n194 , n210 );
    or g445 ( n373 , n402 , n210 );
    xnor g446 ( n463 , n367 , n757 );
    or g447 ( n175 , n768 , n339 );
    nor g448 ( n377 , n17 , n782 );
    nor g449 ( n610 , n37 , n501 );
    xnor g450 ( n779 , n332 , n43 );
    xnor g451 ( n26 , n605 , n616 );
    and g452 ( n488 , n44 , n380 );
    and g453 ( n99 , n656 , n211 );
    or g454 ( n347 , n393 , n403 );
    or g455 ( n283 , n151 , n585 );
    not g456 ( n353 , n348 );
    or g457 ( n703 , n48 , n1 );
    and g458 ( n729 , n312 , n326 );
    xnor g459 ( n291 , n642 , n606 );
    xnor g460 ( n638 , n42 , n29 );
    nor g461 ( n448 , n283 , n677 );
    and g462 ( n248 , n126 , n567 );
    xnor g463 ( n679 , n245 , n143 );
    nor g464 ( n395 , n452 , n451 );
    or g465 ( n625 , n238 , n514 );
    xnor g466 ( n71 , n162 , n147 );
    nor g467 ( n731 , n656 , n156 );
    not g468 ( n38 , n93 );
    or g469 ( n363 , n452 , n771 );
    nor g470 ( n124 , n739 , n279 );
    nor g471 ( n374 , n5 , n671 );
    xnor g472 ( n538 , n188 , n446 );
    nor g473 ( n426 , n555 , n729 );
    or g474 ( n579 , n656 , n109 );
    and g475 ( n295 , n89 , n6 );
    or g476 ( n584 , n449 , n265 );
    or g477 ( n650 , n452 , n557 );
    or g478 ( n15 , n711 , n106 );
    nor g479 ( n313 , n167 , n291 );
    nor g480 ( n82 , n184 , n240 );
    nor g481 ( n536 , n249 , n439 );
    nor g482 ( n710 , n633 , n730 );
    or g483 ( n361 , n573 , n199 );
    and g484 ( n564 , n716 , n40 );
    and g485 ( n392 , n407 , n163 );
    not g486 ( n121 , n550 );
    or g487 ( n491 , n70 , n498 );
    not g488 ( n179 , n228 );
    nor g489 ( n562 , n452 , n54 );
    or g490 ( n623 , n52 , n123 );
    xnor g491 ( n33 , n22 , n750 );
    and g492 ( n180 , n147 , n523 );
    not g493 ( n285 , n725 );
    and g494 ( n68 , n112 , n316 );
    nor g495 ( n478 , n231 , n194 );
    nor g496 ( n498 , n507 , n243 );
    or g497 ( n715 , n391 , n767 );
    not g498 ( n320 , n129 );
    not g499 ( n677 , n335 );
    not g500 ( n92 , n511 );
    and g501 ( n79 , n104 , n50 );
    nor g502 ( n212 , n201 , n499 );
    xnor g503 ( n575 , n188 , n277 );
    or g504 ( n326 , n352 , n216 );
    and g505 ( n713 , n788 , n614 );
    not g506 ( n709 , n643 );
    or g507 ( n437 , n393 , n651 );
    and g508 ( n379 , n726 , n193 );
    not g509 ( n275 , n95 );
    not g510 ( n116 , n22 );
    nor g511 ( n388 , n22 , n399 );
    and g512 ( n310 , n410 , n452 );
    not g513 ( n556 , n60 );
    nor g514 ( n651 , n601 , n683 );
    and g515 ( n601 , n403 , n317 );
    and g516 ( n335 , n736 , n233 );
    not g517 ( n739 , n403 );
    or g518 ( n276 , n709 , n255 );
    or g519 ( n515 , n653 , n719 );
    or g520 ( n481 , n393 , n427 );
    and g521 ( n571 , n656 , n195 );
    not g522 ( n617 , n63 );
    and g523 ( n696 , n378 , n622 );
    nor g524 ( n464 , n452 , n575 );
    or g525 ( n245 , n466 , n571 );
    or g526 ( n672 , n438 , n322 );
    or g527 ( n504 , n302 , n63 );
    or g528 ( n176 , n762 , n486 );
    nor g529 ( n271 , n656 , n541 );
    or g530 ( n419 , n126 , n333 );
    and g531 ( n522 , n31 , n707 );
    xnor g532 ( n165 , n283 , n335 );
    or g533 ( n670 , n656 , n530 );
    nor g534 ( n11 , n617 , n638 );
    and g535 ( n261 , n656 , n406 );
    xnor g536 ( n568 , n411 , n357 );
    nor g537 ( n150 , n104 , n50 );
    xnor g538 ( n141 , n249 , n439 );
    not g539 ( n662 , n86 );
    not g540 ( n734 , n58 );
    not g541 ( n40 , n475 );
    xnor g542 ( n401 , n262 , n204 );
    or g543 ( n397 , n448 , n411 );
    or g544 ( n112 , n559 , n526 );
    and g545 ( n334 , n472 , n677 );
    and g546 ( n567 , n275 , n450 );
    nor g547 ( n572 , n537 , n328 );
    not g548 ( n171 , n276 );
    or g549 ( n294 , n342 , n115 );
    nor g550 ( n748 , n452 , n561 );
    or g551 ( n509 , n205 , n100 );
    or g552 ( n159 , n329 , n764 );
    or g553 ( n272 , n393 , n403 );
    or g554 ( n352 , n664 , n784 );
    nor g555 ( n282 , n456 , n203 );
    and g556 ( n19 , n227 , n142 );
    nor g557 ( n94 , n521 , n180 );
    nor g558 ( n580 , n82 , n422 );
    or g559 ( n279 , n23 , n619 );
    nor g560 ( n280 , n680 , n594 );
    and g561 ( n7 , n656 , n263 );
    xnor g562 ( n616 , n42 , n68 );
    not g563 ( n265 , n365 );
    not g564 ( n423 , n13 );
    or g565 ( n751 , n646 , n628 );
    not g566 ( n523 , n162 );
    nor g567 ( n425 , n452 , n463 );
    not g568 ( n125 , n36 );
    not g569 ( n372 , n343 );
    and g570 ( n253 , n346 , n452 );
    xnor g571 ( n665 , n693 , n17 );
    nor g572 ( n160 , n656 , n565 );
    nor g573 ( n633 , n86 , n592 );
    or g574 ( n627 , n640 , n634 );
    xnor g575 ( n195 , n41 , n208 );
    not g576 ( n390 , n262 );
    and g577 ( n446 , n159 , n318 );
    xnor g578 ( n631 , n726 , n734 );
    not g579 ( n542 , n239 );
    not g580 ( n711 , n139 );
    nor g581 ( n577 , n133 , n325 );
    and g582 ( n87 , n583 , n645 );
    and g583 ( n708 , n656 , n401 );
    xnor g584 ( n744 , n178 , n503 );
    or g585 ( n599 , n334 , n153 );
    or g586 ( n598 , n452 , n79 );
    or g587 ( n43 , n215 , n528 );
    or g588 ( n761 , n733 , n602 );
    not g589 ( n422 , n634 );
    and g590 ( n78 , n66 , n769 );
    not g591 ( n366 , n350 );
    and g592 ( n757 , n709 , n780 );
    xnor g593 ( n418 , n5 , n365 );
    nor g594 ( n649 , n95 , n103 );
    and g595 ( n284 , n402 , n194 );
    not g596 ( n215 , n690 );
    not g597 ( n414 , n409 );
    nor g598 ( n720 , n503 , n182 );
    xnor g599 ( n451 , n240 , n405 );
    or g600 ( n442 , n122 , n562 );
    or g601 ( n325 , n759 , n278 );
    nor g602 ( n745 , n300 , n517 );
    not g603 ( n107 , n671 );
    not g604 ( n626 , n188 );
    or g605 ( n240 , n382 , n689 );
    and g606 ( n420 , n231 , n210 );
    nor g607 ( n135 , n545 , n523 );
    or g608 ( n301 , n127 , n738 );
    xnor g609 ( n674 , n643 , n490 );
    xnor g610 ( n44 , n231 , n210 );
    nor g611 ( n96 , n306 , n100 );
    nor g612 ( n205 , n503 , n383 );
    nor g613 ( n315 , n352 , n516 );
    or g614 ( n367 , n181 , n168 );
    not g615 ( n57 , n258 );
    nor g616 ( n705 , n17 , n13 );
    xnor g617 ( n61 , n17 , n782 );
    and g618 ( n550 , n204 , n390 );
    nor g619 ( n624 , n305 , n138 );
    not g620 ( n164 , n314 );
    xnor g621 ( n714 , n642 , n111 );
    not g622 ( n468 , n289 );
    nor g623 ( n47 , n119 , n579 );
    not g624 ( n608 , n187 );
    or g625 ( n647 , n167 , n252 );
    or g626 ( n629 , n420 , n421 );
    or g627 ( n700 , n253 , n773 );
    or g628 ( n630 , n234 , n425 );
    nor g629 ( n654 , n209 , n734 );
    nor g630 ( n216 , n439 , n742 );
    and g631 ( n293 , n80 , n452 );
    or g632 ( n266 , n537 , n300 );
    not g633 ( n728 , n777 );
    nor g634 ( n128 , n426 , n301 );
    not g635 ( n449 , n217 );
    not g636 ( n689 , n667 );
    and g637 ( n337 , n593 , n452 );
    nor g638 ( n2 , n435 , n285 );
    or g639 ( n765 , n338 , n569 );
    or g640 ( n162 , n146 , n394 );
    xnor g641 ( n140 , n213 , n542 );
    and g642 ( n436 , n306 , n100 );
    nor g643 ( n338 , n656 , n570 );
    and g644 ( n237 , n626 , n277 );
    xnor g645 ( n136 , n611 , n744 );
    not g646 ( n752 , n605 );
    or g647 ( n619 , n391 , n751 );
    or g648 ( n18 , n548 , n25 );
    nor g649 ( n485 , n659 , n502 );
    nor g650 ( n543 , n452 , n308 );
    nor g651 ( n342 , n656 , n675 );
    not g652 ( n4 , n180 );
    and g653 ( n539 , n656 , n34 );
    nor g654 ( n431 , n192 , n273 );
    and g655 ( n455 , n684 , n452 );
    or g656 ( n90 , n92 , n106 );
    or g657 ( n137 , n468 , n106 );
    xnor g658 ( n304 , n625 , n665 );
    and g659 ( n232 , n701 , n361 );
    or g660 ( n85 , n96 , n471 );
    or g661 ( n785 , n503 , n611 );
    or g662 ( n27 , n149 , n464 );
    not g663 ( n666 , n505 );
    and g664 ( n210 , n437 , n8 );
    nor g665 ( n358 , n739 , n775 );
    xnor g666 ( n496 , n199 , n370 );
    not g667 ( n21 , n629 );
    or g668 ( n184 , n337 , n500 );
    xnor g669 ( n259 , n584 , n217 );
    xnor g670 ( n541 , n245 , n530 );
    nor g671 ( n298 , n281 , n132 );
    not g672 ( n49 , n232 );
    xnor g673 ( n10 , n187 , n237 );
    or g674 ( n299 , n366 , n721 );
    or g675 ( n722 , n43 , n332 );
    or g676 ( n88 , n560 , n725 );
    xnor g677 ( n344 , n351 , n457 );
    nor g678 ( n12 , n452 , n108 );
    or g679 ( n188 , n510 , n77 );
    nor g680 ( n653 , n656 , n118 );
    not g681 ( n459 , n105 );
    xnor g682 ( n178 , n259 , n690 );
    nor g683 ( n427 , n124 , n282 );
    nor g684 ( n328 , n492 , n745 );
    or g685 ( n355 , n414 , n664 );
    nor g686 ( n545 , n190 , n564 );
    or g687 ( n767 , n646 , n265 );
    and g688 ( n613 , n656 , n710 );
    or g689 ( n120 , n547 , n260 );
    or g690 ( n570 , n254 , n542 );
    not g691 ( n318 , n419 );
    and g692 ( n151 , n219 , n452 );
    nor g693 ( n637 , n452 , n723 );
    xnor g694 ( n306 , n383 , n503 );
    xnor g695 ( n453 , n123 , n680 );
    not g696 ( n524 , n223 );
    or g697 ( n787 , n527 , n689 );
    and g698 ( n72 , n452 , n654 );
    nor g699 ( n234 , n656 , n398 );
    and g700 ( n166 , n17 , n782 );
    or g701 ( n60 , n522 , n360 );
    and g702 ( n738 , n555 , n729 );
    and g703 ( n83 , n656 , n551 );
endmodule
