// Benchmark "top" written by ABC on Mon Jun 12 20:56:48 2023

module top ( 
    \1_n0 , \1_n1005 , \1_n1022 , \1_n1029 , \1_n1035 , \1_n1036 ,
    \1_n104 , \1_n1041 , \1_n1044 , \1_n1045 , \1_n1048 , \1_n1064 ,
    \1_n1067 , \1_n1069 , \1_n107 , \1_n1072 , \1_n1073 , \1_n1077 ,
    \1_n108 , \1_n1080 , \1_n1081 , \1_n1089 , \1_n1091 , \1_n1097 ,
    \1_n1098 , \1_n1120 , \1_n1131 , \1_n1132 , \1_n1140 , \1_n1141 ,
    \1_n1143 , \1_n1146 , \1_n1151 , \1_n116 , \1_n1163 , \1_n1164 ,
    \1_n1180 , \1_n1191 , \1_n1198 , \1_n1219 , \1_n122 , \1_n1226 ,
    \1_n1229 , \1_n1231 , \1_n1236 , \1_n1257 , \1_n1269 , \1_n127 ,
    \1_n1273 , \1_n1277 , \1_n1279 , \1_n128 , \1_n1298 , \1_n1308 ,
    \1_n1311 , \1_n1321 , \1_n1326 , \1_n1342 , \1_n1344 , \1_n1352 ,
    \1_n138 , \1_n153 , \1_n192 , \1_n196 , \1_n200 , \1_n208 , \1_n21 ,
    \1_n221 , \1_n231 , \1_n236 , \1_n244 , \1_n245 , \1_n246 , \1_n252 ,
    \1_n258 , \1_n260 , \1_n262 , \1_n267 , \1_n268 , \1_n281 , \1_n284 ,
    \1_n288 , \1_n301 , \1_n305 , \1_n310 , \1_n319 , \1_n323 , \1_n324 ,
    \1_n332 , \1_n336 , \1_n359 , \1_n36 , \1_n360 , \1_n364 , \1_n366 ,
    \1_n38 , \1_n381 , \1_n384 , \1_n393 , \1_n398 , \1_n421 , \1_n423 ,
    \1_n431 , \1_n433 , \1_n438 , \1_n439 , \1_n441 , \1_n444 , \1_n448 ,
    \1_n449 , \1_n45 , \1_n475 , \1_n49 , \1_n491 , \1_n500 , \1_n505 ,
    \1_n507 , \1_n510 , \1_n519 , \1_n532 , \1_n536 , \1_n540 , \1_n571 ,
    \1_n577 , \1_n589 , \1_n599 , \1_n610 , \1_n631 , \1_n635 , \1_n640 ,
    \1_n644 , \1_n650 , \1_n657 , \1_n667 , \1_n685 , \1_n688 , \1_n695 ,
    \1_n714 , \1_n716 , \1_n741 , \1_n745 , \1_n749 , \1_n766 , \1_n767 ,
    \1_n77 , \1_n771 , \1_n774 , \1_n787 , \1_n802 , \1_n804 , \1_n806 ,
    \1_n818 , \1_n819 , \1_n823 , \1_n825 , \1_n826 , \1_n833 , \1_n839 ,
    \1_n841 , \1_n845 , \1_n851 , \1_n857 , \1_n862 , \1_n863 , \1_n866 ,
    \1_n870 , \1_n879 , \1_n893 , \1_n896 , \1_n901 , \1_n928 , \1_n929 ,
    \1_n936 , \1_n944 , \1_n95 , \1_n952 , \1_n955 , \1_n961 , \1_n975 ,
    \1_n976 , \1_n98 , \1_n986 , \1_n997 , \2_n1023 , \2_n1040 , \2_n1044 ,
    \2_n1054 , \2_n1061 , \2_n107 , \2_n1071 , \2_n1095 , \2_n11 ,
    \2_n1103 , \2_n1114 , \2_n1121 , \2_n1138 , \2_n1152 , \2_n1154 ,
    \2_n1156 , \2_n1164 , \2_n117 , \2_n1172 , \2_n1175 , \2_n1187 ,
    \2_n1191 , \2_n1193 , \2_n1205 , \2_n1225 , \2_n1227 , \2_n1239 ,
    \2_n1246 , \2_n1250 , \2_n1263 , \2_n1278 , \2_n1281 , \2_n1283 ,
    \2_n1286 , \2_n1289 , \2_n1299 , \2_n1301 , \2_n1305 , \2_n1345 ,
    \2_n1346 , \2_n1350 , \2_n1361 , \2_n138 , \2_n1386 , \2_n1387 ,
    \2_n1389 , \2_n1393 , \2_n1401 , \2_n1411 , \2_n1415 , \2_n1418 ,
    \2_n1428 , \2_n143 , \2_n1435 , \2_n1438 , \2_n1443 , \2_n1446 ,
    \2_n1448 , \2_n1463 , \2_n1470 , \2_n1474 , \2_n1476 , \2_n1500 ,
    \2_n1502 , \2_n1506 , \2_n1516 , \2_n1520 , \2_n1521 , \2_n1523 ,
    \2_n153 , \2_n1536 , \2_n155 , \2_n156 , \2_n1566 , \2_n1569 ,
    \2_n1576 , \2_n1586 , \2_n159 , \2_n1592 , \2_n1609 , \2_n1613 ,
    \2_n1616 , \2_n1626 , \2_n1627 , \2_n1644 , \2_n1647 , \2_n1656 ,
    \2_n1750 , \2_n1753 , \2_n200 , \2_n21 , \2_n219 , \2_n220 , \2_n222 ,
    \2_n223 , \2_n243 , \2_n244 , \2_n246 , \2_n251 , \2_n254 , \2_n262 ,
    \2_n268 , \2_n273 , \2_n284 , \2_n288 , \2_n29 , \2_n293 , \2_n299 ,
    \2_n300 , \2_n307 , \2_n310 , \2_n312 , \2_n314 , \2_n315 , \2_n318 ,
    \2_n341 , \2_n344 , \2_n346 , \2_n374 , \2_n376 , \2_n380 , \2_n391 ,
    \2_n392 , \2_n399 , \2_n40 , \2_n408 , \2_n409 , \2_n416 , \2_n420 ,
    \2_n430 , \2_n45 , \2_n477 , \2_n478 , \2_n487 , \2_n489 , \2_n50 ,
    \2_n502 , \2_n506 , \2_n507 , \2_n510 , \2_n52 , \2_n54 , \2_n545 ,
    \2_n559 , \2_n56 , \2_n560 , \2_n561 , \2_n567 , \2_n574 , \2_n58 ,
    \2_n581 , \2_n582 , \2_n589 , \2_n593 , \2_n598 , \2_n600 , \2_n607 ,
    \2_n608 , \2_n609 , \2_n626 , \2_n641 , \2_n645 , \2_n663 , \2_n671 ,
    \2_n676 , \2_n690 , \2_n695 , \2_n701 , \2_n71 , \2_n710 , \2_n727 ,
    \2_n729 , \2_n734 , \2_n742 , \2_n743 , \2_n755 , \2_n769 , \2_n77 ,
    \2_n775 , \2_n778 , \2_n779 , \2_n787 , \2_n790 , \2_n82 , \2_n823 ,
    \2_n831 , \2_n832 , \2_n839 , \2_n849 , \2_n86 , \2_n87 , \2_n879 ,
    \2_n882 , \2_n885 , \2_n905 , \2_n920 , \2_n936 , \2_n94 , \2_n947 ,
    \2_n953 , \2_n961 , \2_n969 , \2_n980 , \2_n984 , \2_n986 , \2_n992 ,
    \2_n997 ,
    \1_n1023 , \1_n1027 , \1_n1057 , \1_n1059 , \1_n1061 , \1_n1085 ,
    \1_n1099 , \1_n112 , \1_n1150 , \1_n1153 , \1_n1178 , \1_n1184 ,
    \1_n1194 , \1_n1202 , \1_n1206 , \1_n1232 , \1_n1239 , \1_n1259 ,
    \1_n1264 , \1_n1288 , \1_n129 , \1_n130 , \1_n1301 , \1_n135 ,
    \1_n150 , \1_n159 , \1_n167 , \1_n168 , \1_n175 , \1_n185 , \1_n190 ,
    \1_n193 , \1_n204 , \1_n206 , \1_n207 , \1_n218 , \1_n223 , \1_n227 ,
    \1_n228 , \1_n229 , \1_n240 , \1_n275 , \1_n29 , \1_n299 , \1_n307 ,
    \1_n34 , \1_n342 , \1_n347 , \1_n374 , \1_n383 , \1_n389 , \1_n408 ,
    \1_n409 , \1_n410 , \1_n415 , \1_n432 , \1_n452 , \1_n456 , \1_n492 ,
    \1_n516 , \1_n554 , \1_n580 , \1_n592 , \1_n598 , \1_n60 , \1_n607 ,
    \1_n608 , \1_n613 , \1_n617 , \1_n621 , \1_n623 , \1_n627 , \1_n638 ,
    \1_n651 , \1_n653 , \1_n662 , \1_n679 , \1_n683 , \1_n707 , \1_n710 ,
    \1_n718 , \1_n723 , \1_n733 , \1_n734 , \1_n747 , \1_n779 , \1_n785 ,
    \1_n801 , \1_n807 , \1_n808 , \1_n81 , \1_n817 , \1_n82 , \1_n835 ,
    \1_n842 , \1_n853 , \1_n854 , \1_n877 , \1_n88 , \1_n90 , \1_n905 ,
    \1_n908 , \1_n91 , \1_n927 , \1_n962 , \1_n966 , \1_n973 , \1_n999 ,
    \2_n1006 , \2_n1017 , \2_n1042 , \2_n1050 , \2_n1051 , \2_n1058 ,
    \2_n1060 , \2_n1063 , \2_n1065 , \2_n112 , \2_n1177 , \2_n1186 ,
    \2_n1195 , \2_n1209 , \2_n1211 , \2_n1231 , \2_n1234 , \2_n1253 ,
    \2_n126 , \2_n1285 , \2_n1288 , \2_n1292 , \2_n1296 , \2_n130 ,
    \2_n1302 , \2_n1306 , \2_n1320 , \2_n1322 , \2_n1337 , \2_n1359 ,
    \2_n1368 , \2_n1375 , \2_n1391 , \2_n1420 , \2_n1421 , \2_n1427 ,
    \2_n1527 , \2_n1534 , \2_n1547 , \2_n1548 , \2_n1588 , \2_n1594 ,
    \2_n161 , \2_n1632 , \2_n1639 , \2_n164 , \2_n1645 , \2_n1687 ,
    \2_n1729 , \2_n173 , \2_n1738 , \2_n1752 , \2_n181 , \2_n184 ,
    \2_n216 , \2_n22 , \2_n23 , \2_n230 , \2_n233 , \2_n247 , \2_n27 ,
    \2_n275 , \2_n292 , \2_n30 , \2_n301 , \2_n304 , \2_n337 , \2_n352 ,
    \2_n362 , \2_n364 , \2_n370 , \2_n378 , \2_n396 , \2_n417 , \2_n428 ,
    \2_n453 , \2_n457 , \2_n460 , \2_n497 , \2_n498 , \2_n501 , \2_n509 ,
    \2_n516 , \2_n517 , \2_n534 , \2_n553 , \2_n585 , \2_n595 , \2_n597 ,
    \2_n625 , \2_n638 , \2_n640 , \2_n669 , \2_n693 , \2_n714 , \2_n719 ,
    \2_n726 , \2_n773 , \2_n782 , \2_n794 , \2_n821 , \2_n842 , \2_n85 ,
    \2_n894 , \2_n916 , \2_n918 , \2_n952 , \2_n990   );
  input  \1_n0 , \1_n1005 , \1_n1022 , \1_n1029 , \1_n1035 , \1_n1036 ,
    \1_n104 , \1_n1041 , \1_n1044 , \1_n1045 , \1_n1048 , \1_n1064 ,
    \1_n1067 , \1_n1069 , \1_n107 , \1_n1072 , \1_n1073 , \1_n1077 ,
    \1_n108 , \1_n1080 , \1_n1081 , \1_n1089 , \1_n1091 , \1_n1097 ,
    \1_n1098 , \1_n1120 , \1_n1131 , \1_n1132 , \1_n1140 , \1_n1141 ,
    \1_n1143 , \1_n1146 , \1_n1151 , \1_n116 , \1_n1163 , \1_n1164 ,
    \1_n1180 , \1_n1191 , \1_n1198 , \1_n1219 , \1_n122 , \1_n1226 ,
    \1_n1229 , \1_n1231 , \1_n1236 , \1_n1257 , \1_n1269 , \1_n127 ,
    \1_n1273 , \1_n1277 , \1_n1279 , \1_n128 , \1_n1298 , \1_n1308 ,
    \1_n1311 , \1_n1321 , \1_n1326 , \1_n1342 , \1_n1344 , \1_n1352 ,
    \1_n138 , \1_n153 , \1_n192 , \1_n196 , \1_n200 , \1_n208 , \1_n21 ,
    \1_n221 , \1_n231 , \1_n236 , \1_n244 , \1_n245 , \1_n246 , \1_n252 ,
    \1_n258 , \1_n260 , \1_n262 , \1_n267 , \1_n268 , \1_n281 , \1_n284 ,
    \1_n288 , \1_n301 , \1_n305 , \1_n310 , \1_n319 , \1_n323 , \1_n324 ,
    \1_n332 , \1_n336 , \1_n359 , \1_n36 , \1_n360 , \1_n364 , \1_n366 ,
    \1_n38 , \1_n381 , \1_n384 , \1_n393 , \1_n398 , \1_n421 , \1_n423 ,
    \1_n431 , \1_n433 , \1_n438 , \1_n439 , \1_n441 , \1_n444 , \1_n448 ,
    \1_n449 , \1_n45 , \1_n475 , \1_n49 , \1_n491 , \1_n500 , \1_n505 ,
    \1_n507 , \1_n510 , \1_n519 , \1_n532 , \1_n536 , \1_n540 , \1_n571 ,
    \1_n577 , \1_n589 , \1_n599 , \1_n610 , \1_n631 , \1_n635 , \1_n640 ,
    \1_n644 , \1_n650 , \1_n657 , \1_n667 , \1_n685 , \1_n688 , \1_n695 ,
    \1_n714 , \1_n716 , \1_n741 , \1_n745 , \1_n749 , \1_n766 , \1_n767 ,
    \1_n77 , \1_n771 , \1_n774 , \1_n787 , \1_n802 , \1_n804 , \1_n806 ,
    \1_n818 , \1_n819 , \1_n823 , \1_n825 , \1_n826 , \1_n833 , \1_n839 ,
    \1_n841 , \1_n845 , \1_n851 , \1_n857 , \1_n862 , \1_n863 , \1_n866 ,
    \1_n870 , \1_n879 , \1_n893 , \1_n896 , \1_n901 , \1_n928 , \1_n929 ,
    \1_n936 , \1_n944 , \1_n95 , \1_n952 , \1_n955 , \1_n961 , \1_n975 ,
    \1_n976 , \1_n98 , \1_n986 , \1_n997 , \2_n1023 , \2_n1040 , \2_n1044 ,
    \2_n1054 , \2_n1061 , \2_n107 , \2_n1071 , \2_n1095 , \2_n11 ,
    \2_n1103 , \2_n1114 , \2_n1121 , \2_n1138 , \2_n1152 , \2_n1154 ,
    \2_n1156 , \2_n1164 , \2_n117 , \2_n1172 , \2_n1175 , \2_n1187 ,
    \2_n1191 , \2_n1193 , \2_n1205 , \2_n1225 , \2_n1227 , \2_n1239 ,
    \2_n1246 , \2_n1250 , \2_n1263 , \2_n1278 , \2_n1281 , \2_n1283 ,
    \2_n1286 , \2_n1289 , \2_n1299 , \2_n1301 , \2_n1305 , \2_n1345 ,
    \2_n1346 , \2_n1350 , \2_n1361 , \2_n138 , \2_n1386 , \2_n1387 ,
    \2_n1389 , \2_n1393 , \2_n1401 , \2_n1411 , \2_n1415 , \2_n1418 ,
    \2_n1428 , \2_n143 , \2_n1435 , \2_n1438 , \2_n1443 , \2_n1446 ,
    \2_n1448 , \2_n1463 , \2_n1470 , \2_n1474 , \2_n1476 , \2_n1500 ,
    \2_n1502 , \2_n1506 , \2_n1516 , \2_n1520 , \2_n1521 , \2_n1523 ,
    \2_n153 , \2_n1536 , \2_n155 , \2_n156 , \2_n1566 , \2_n1569 ,
    \2_n1576 , \2_n1586 , \2_n159 , \2_n1592 , \2_n1609 , \2_n1613 ,
    \2_n1616 , \2_n1626 , \2_n1627 , \2_n1644 , \2_n1647 , \2_n1656 ,
    \2_n1750 , \2_n1753 , \2_n200 , \2_n21 , \2_n219 , \2_n220 , \2_n222 ,
    \2_n223 , \2_n243 , \2_n244 , \2_n246 , \2_n251 , \2_n254 , \2_n262 ,
    \2_n268 , \2_n273 , \2_n284 , \2_n288 , \2_n29 , \2_n293 , \2_n299 ,
    \2_n300 , \2_n307 , \2_n310 , \2_n312 , \2_n314 , \2_n315 , \2_n318 ,
    \2_n341 , \2_n344 , \2_n346 , \2_n374 , \2_n376 , \2_n380 , \2_n391 ,
    \2_n392 , \2_n399 , \2_n40 , \2_n408 , \2_n409 , \2_n416 , \2_n420 ,
    \2_n430 , \2_n45 , \2_n477 , \2_n478 , \2_n487 , \2_n489 , \2_n50 ,
    \2_n502 , \2_n506 , \2_n507 , \2_n510 , \2_n52 , \2_n54 , \2_n545 ,
    \2_n559 , \2_n56 , \2_n560 , \2_n561 , \2_n567 , \2_n574 , \2_n58 ,
    \2_n581 , \2_n582 , \2_n589 , \2_n593 , \2_n598 , \2_n600 , \2_n607 ,
    \2_n608 , \2_n609 , \2_n626 , \2_n641 , \2_n645 , \2_n663 , \2_n671 ,
    \2_n676 , \2_n690 , \2_n695 , \2_n701 , \2_n71 , \2_n710 , \2_n727 ,
    \2_n729 , \2_n734 , \2_n742 , \2_n743 , \2_n755 , \2_n769 , \2_n77 ,
    \2_n775 , \2_n778 , \2_n779 , \2_n787 , \2_n790 , \2_n82 , \2_n823 ,
    \2_n831 , \2_n832 , \2_n839 , \2_n849 , \2_n86 , \2_n87 , \2_n879 ,
    \2_n882 , \2_n885 , \2_n905 , \2_n920 , \2_n936 , \2_n94 , \2_n947 ,
    \2_n953 , \2_n961 , \2_n969 , \2_n980 , \2_n984 , \2_n986 , \2_n992 ,
    \2_n997 ;
  output \1_n1023 , \1_n1027 , \1_n1057 , \1_n1059 , \1_n1061 , \1_n1085 ,
    \1_n1099 , \1_n112 , \1_n1150 , \1_n1153 , \1_n1178 , \1_n1184 ,
    \1_n1194 , \1_n1202 , \1_n1206 , \1_n1232 , \1_n1239 , \1_n1259 ,
    \1_n1264 , \1_n1288 , \1_n129 , \1_n130 , \1_n1301 , \1_n135 ,
    \1_n150 , \1_n159 , \1_n167 , \1_n168 , \1_n175 , \1_n185 , \1_n190 ,
    \1_n193 , \1_n204 , \1_n206 , \1_n207 , \1_n218 , \1_n223 , \1_n227 ,
    \1_n228 , \1_n229 , \1_n240 , \1_n275 , \1_n29 , \1_n299 , \1_n307 ,
    \1_n34 , \1_n342 , \1_n347 , \1_n374 , \1_n383 , \1_n389 , \1_n408 ,
    \1_n409 , \1_n410 , \1_n415 , \1_n432 , \1_n452 , \1_n456 , \1_n492 ,
    \1_n516 , \1_n554 , \1_n580 , \1_n592 , \1_n598 , \1_n60 , \1_n607 ,
    \1_n608 , \1_n613 , \1_n617 , \1_n621 , \1_n623 , \1_n627 , \1_n638 ,
    \1_n651 , \1_n653 , \1_n662 , \1_n679 , \1_n683 , \1_n707 , \1_n710 ,
    \1_n718 , \1_n723 , \1_n733 , \1_n734 , \1_n747 , \1_n779 , \1_n785 ,
    \1_n801 , \1_n807 , \1_n808 , \1_n81 , \1_n817 , \1_n82 , \1_n835 ,
    \1_n842 , \1_n853 , \1_n854 , \1_n877 , \1_n88 , \1_n90 , \1_n905 ,
    \1_n908 , \1_n91 , \1_n927 , \1_n962 , \1_n966 , \1_n973 , \1_n999 ,
    \2_n1006 , \2_n1017 , \2_n1042 , \2_n1050 , \2_n1051 , \2_n1058 ,
    \2_n1060 , \2_n1063 , \2_n1065 , \2_n112 , \2_n1177 , \2_n1186 ,
    \2_n1195 , \2_n1209 , \2_n1211 , \2_n1231 , \2_n1234 , \2_n1253 ,
    \2_n126 , \2_n1285 , \2_n1288 , \2_n1292 , \2_n1296 , \2_n130 ,
    \2_n1302 , \2_n1306 , \2_n1320 , \2_n1322 , \2_n1337 , \2_n1359 ,
    \2_n1368 , \2_n1375 , \2_n1391 , \2_n1420 , \2_n1421 , \2_n1427 ,
    \2_n1527 , \2_n1534 , \2_n1547 , \2_n1548 , \2_n1588 , \2_n1594 ,
    \2_n161 , \2_n1632 , \2_n1639 , \2_n164 , \2_n1645 , \2_n1687 ,
    \2_n1729 , \2_n173 , \2_n1738 , \2_n1752 , \2_n181 , \2_n184 ,
    \2_n216 , \2_n22 , \2_n23 , \2_n230 , \2_n233 , \2_n247 , \2_n27 ,
    \2_n275 , \2_n292 , \2_n30 , \2_n301 , \2_n304 , \2_n337 , \2_n352 ,
    \2_n362 , \2_n364 , \2_n370 , \2_n378 , \2_n396 , \2_n417 , \2_n428 ,
    \2_n453 , \2_n457 , \2_n460 , \2_n497 , \2_n498 , \2_n501 , \2_n509 ,
    \2_n516 , \2_n517 , \2_n534 , \2_n553 , \2_n585 , \2_n595 , \2_n597 ,
    \2_n625 , \2_n638 , \2_n640 , \2_n669 , \2_n693 , \2_n714 , \2_n719 ,
    \2_n726 , \2_n773 , \2_n782 , \2_n794 , \2_n821 , \2_n842 , \2_n85 ,
    \2_n894 , \2_n916 , \2_n918 , \2_n952 , \2_n990 ;
  wire new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n932_,
    new_n933_, new_n934_, new_n935_, new_n936_, new_n937_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n964_, new_n965_, new_n966_, new_n967_, new_n968_, new_n969_,
    new_n970_, new_n971_, new_n972_, new_n973_, new_n974_, new_n975_,
    new_n976_, new_n977_, new_n978_, new_n979_, new_n980_, new_n981_,
    new_n982_, new_n983_, new_n984_, new_n985_, new_n986_, new_n987_,
    new_n988_, new_n989_, new_n990_, new_n991_, new_n992_, new_n993_,
    new_n994_, new_n995_, new_n996_, new_n997_, new_n998_, new_n999_,
    new_n1000_, new_n1001_, new_n1002_, new_n1003_, new_n1004_, new_n1005_,
    new_n1006_, new_n1007_, new_n1008_, new_n1009_, new_n1010_, new_n1011_,
    new_n1012_, new_n1013_, new_n1014_, new_n1015_, new_n1016_, new_n1017_,
    new_n1018_, new_n1019_, new_n1020_, new_n1021_, new_n1022_, new_n1023_,
    new_n1024_, new_n1025_, new_n1026_, new_n1027_, new_n1028_, new_n1029_,
    new_n1030_, new_n1031_, new_n1032_, new_n1033_, new_n1034_, new_n1035_,
    new_n1036_, new_n1037_, new_n1038_, new_n1039_, new_n1040_, new_n1041_,
    new_n1042_, new_n1043_, new_n1044_, new_n1045_, new_n1046_, new_n1047_,
    new_n1048_, new_n1049_, new_n1050_, new_n1051_, new_n1052_, new_n1053_,
    new_n1054_, new_n1055_, new_n1056_, new_n1057_, new_n1058_, new_n1059_,
    new_n1060_, new_n1061_, new_n1062_, new_n1063_, new_n1064_, new_n1065_,
    new_n1066_, new_n1067_, new_n1068_, new_n1069_, new_n1070_, new_n1071_,
    new_n1072_, new_n1073_, new_n1074_, new_n1075_, new_n1076_, new_n1077_,
    new_n1078_, new_n1079_, new_n1080_, new_n1081_, new_n1082_, new_n1083_,
    new_n1084_, new_n1085_, new_n1086_, new_n1087_, new_n1088_, new_n1089_,
    new_n1090_, new_n1091_, new_n1092_, new_n1093_, new_n1094_, new_n1095_,
    new_n1096_, new_n1098_, new_n1099_, new_n1102_, new_n1103_, new_n1104_,
    new_n1105_, new_n1106_, new_n1107_, new_n1108_, new_n1109_, new_n1110_,
    new_n1111_, new_n1112_, new_n1113_, new_n1115_, new_n1116_, new_n1118_,
    new_n1119_, new_n1120_, new_n1121_, new_n1122_, new_n1123_, new_n1124_,
    new_n1125_, new_n1126_, new_n1127_, new_n1128_, new_n1129_, new_n1130_,
    new_n1131_, new_n1132_, new_n1133_, new_n1134_, new_n1135_, new_n1136_,
    new_n1137_, new_n1138_, new_n1139_, new_n1141_, new_n1142_, new_n1143_,
    new_n1145_, new_n1146_, new_n1148_, new_n1149_, new_n1150_, new_n1151_,
    new_n1152_, new_n1153_, new_n1154_, new_n1155_, new_n1156_, new_n1157_,
    new_n1158_, new_n1159_, new_n1160_, new_n1161_, new_n1162_, new_n1163_,
    new_n1164_, new_n1165_, new_n1166_, new_n1167_, new_n1168_, new_n1169_,
    new_n1170_, new_n1171_, new_n1172_, new_n1173_, new_n1174_, new_n1175_,
    new_n1176_, new_n1177_, new_n1178_, new_n1179_, new_n1180_, new_n1181_,
    new_n1182_, new_n1183_, new_n1184_, new_n1185_, new_n1186_, new_n1187_,
    new_n1188_, new_n1189_, new_n1190_, new_n1191_, new_n1192_, new_n1193_,
    new_n1194_, new_n1195_, new_n1196_, new_n1197_, new_n1198_, new_n1199_,
    new_n1200_, new_n1201_, new_n1202_, new_n1203_, new_n1204_, new_n1205_,
    new_n1206_, new_n1207_, new_n1208_, new_n1209_, new_n1210_, new_n1211_,
    new_n1212_, new_n1213_, new_n1214_, new_n1215_, new_n1216_, new_n1217_,
    new_n1218_, new_n1219_, new_n1220_, new_n1221_, new_n1222_, new_n1223_,
    new_n1224_, new_n1225_, new_n1226_, new_n1227_, new_n1228_, new_n1229_,
    new_n1231_, new_n1232_, new_n1234_, new_n1235_, new_n1236_, new_n1237_,
    new_n1238_, new_n1239_, new_n1240_, new_n1241_, new_n1242_, new_n1243_,
    new_n1244_, new_n1245_, new_n1246_, new_n1247_, new_n1248_, new_n1249_,
    new_n1250_, new_n1252_, new_n1253_, new_n1254_, new_n1256_, new_n1260_,
    new_n1262_, new_n1263_, new_n1264_, new_n1265_, new_n1266_, new_n1267_,
    new_n1268_, new_n1269_, new_n1270_, new_n1271_, new_n1272_, new_n1273_,
    new_n1274_, new_n1275_, new_n1276_, new_n1277_, new_n1278_, new_n1279_,
    new_n1280_, new_n1281_, new_n1282_, new_n1283_, new_n1284_, new_n1285_,
    new_n1286_, new_n1287_, new_n1288_, new_n1289_, new_n1290_, new_n1291_,
    new_n1292_, new_n1293_, new_n1294_, new_n1295_, new_n1296_, new_n1297_,
    new_n1298_, new_n1299_, new_n1300_, new_n1301_, new_n1302_, new_n1303_,
    new_n1304_, new_n1305_, new_n1306_, new_n1307_, new_n1308_, new_n1309_,
    new_n1310_, new_n1311_, new_n1312_, new_n1313_, new_n1314_, new_n1315_,
    new_n1316_, new_n1317_, new_n1318_, new_n1319_, new_n1320_, new_n1321_,
    new_n1322_, new_n1323_, new_n1324_, new_n1325_, new_n1326_, new_n1327_,
    new_n1328_, new_n1329_, new_n1330_, new_n1331_, new_n1332_, new_n1333_,
    new_n1334_, new_n1335_, new_n1336_, new_n1337_, new_n1338_, new_n1339_,
    new_n1340_, new_n1341_, new_n1342_, new_n1343_, new_n1344_, new_n1345_,
    new_n1346_, new_n1347_, new_n1348_, new_n1349_, new_n1351_, new_n1353_,
    new_n1354_, new_n1355_, new_n1356_, new_n1357_, new_n1358_, new_n1359_,
    new_n1360_, new_n1361_, new_n1362_, new_n1363_, new_n1364_, new_n1365_,
    new_n1366_, new_n1367_, new_n1368_, new_n1369_, new_n1370_, new_n1371_,
    new_n1372_, new_n1373_, new_n1374_, new_n1375_, new_n1376_, new_n1377_,
    new_n1378_, new_n1379_, new_n1380_, new_n1381_, new_n1382_, new_n1383_,
    new_n1384_, new_n1385_, new_n1386_, new_n1387_, new_n1388_, new_n1389_,
    new_n1390_, new_n1391_, new_n1392_, new_n1393_, new_n1394_, new_n1395_,
    new_n1396_, new_n1397_, new_n1398_, new_n1399_, new_n1400_, new_n1401_,
    new_n1402_, new_n1403_, new_n1404_, new_n1405_, new_n1406_, new_n1407_,
    new_n1408_, new_n1409_, new_n1410_, new_n1411_, new_n1412_, new_n1413_,
    new_n1414_, new_n1415_, new_n1416_, new_n1417_, new_n1418_, new_n1419_,
    new_n1420_, new_n1421_, new_n1422_, new_n1423_, new_n1424_, new_n1425_,
    new_n1426_, new_n1427_, new_n1428_, new_n1429_, new_n1430_, new_n1431_,
    new_n1432_, new_n1433_, new_n1434_, new_n1435_, new_n1436_, new_n1437_,
    new_n1438_, new_n1439_, new_n1440_, new_n1441_, new_n1442_, new_n1443_,
    new_n1444_, new_n1445_, new_n1446_, new_n1447_, new_n1448_, new_n1449_,
    new_n1450_, new_n1451_, new_n1452_, new_n1453_, new_n1454_, new_n1455_,
    new_n1456_, new_n1457_, new_n1458_, new_n1459_, new_n1460_, new_n1462_,
    new_n1463_, new_n1464_, new_n1465_, new_n1466_, new_n1467_, new_n1468_,
    new_n1469_, new_n1470_, new_n1471_, new_n1472_, new_n1473_, new_n1474_,
    new_n1475_, new_n1476_, new_n1477_, new_n1478_, new_n1479_, new_n1480_,
    new_n1481_, new_n1485_, new_n1487_, new_n1488_, new_n1489_, new_n1490_,
    new_n1492_, new_n1493_, new_n1494_, new_n1496_, new_n1498_, new_n1499_,
    new_n1500_, new_n1501_, new_n1502_, new_n1503_, new_n1504_, new_n1505_,
    new_n1506_, new_n1507_, new_n1508_, new_n1509_, new_n1510_, new_n1511_,
    new_n1512_, new_n1513_, new_n1514_, new_n1515_, new_n1516_, new_n1517_,
    new_n1518_, new_n1519_, new_n1520_, new_n1521_, new_n1522_, new_n1523_,
    new_n1524_, new_n1525_, new_n1526_, new_n1527_, new_n1528_, new_n1529_,
    new_n1530_, new_n1531_, new_n1532_, new_n1533_, new_n1534_, new_n1535_,
    new_n1536_, new_n1537_, new_n1538_, new_n1539_, new_n1540_, new_n1541_,
    new_n1542_, new_n1543_, new_n1544_, new_n1545_, new_n1546_, new_n1547_,
    new_n1548_, new_n1549_, new_n1550_, new_n1551_, new_n1552_, new_n1553_,
    new_n1554_, new_n1555_, new_n1556_, new_n1557_, new_n1558_, new_n1559_,
    new_n1560_, new_n1561_, new_n1562_, new_n1563_, new_n1564_, new_n1565_,
    new_n1566_, new_n1567_, new_n1568_, new_n1569_, new_n1570_, new_n1571_,
    new_n1572_, new_n1573_, new_n1574_, new_n1575_, new_n1576_, new_n1577_,
    new_n1578_, new_n1579_, new_n1580_, new_n1581_, new_n1582_, new_n1583_,
    new_n1584_, new_n1585_, new_n1586_, new_n1587_, new_n1588_, new_n1589_,
    new_n1590_, new_n1591_, new_n1592_, new_n1593_, new_n1594_, new_n1595_,
    new_n1597_, new_n1598_, new_n1599_, new_n1600_, new_n1602_, new_n1604_,
    new_n1606_, new_n1608_, new_n1609_, new_n1610_, new_n1611_, new_n1612_,
    new_n1614_, new_n1616_, new_n1617_, new_n1619_, new_n1620_, new_n1621_,
    new_n1622_, new_n1623_, new_n1624_, new_n1625_, new_n1626_, new_n1627_,
    new_n1628_, new_n1629_, new_n1630_, new_n1631_, new_n1632_, new_n1633_,
    new_n1634_, new_n1635_, new_n1636_, new_n1637_, new_n1638_, new_n1639_,
    new_n1640_, new_n1641_, new_n1642_, new_n1643_, new_n1644_, new_n1645_,
    new_n1646_, new_n1647_, new_n1648_, new_n1649_, new_n1650_, new_n1651_,
    new_n1652_, new_n1653_, new_n1654_, new_n1655_, new_n1656_, new_n1657_,
    new_n1658_, new_n1659_, new_n1660_, new_n1661_, new_n1662_, new_n1663_,
    new_n1664_, new_n1665_, new_n1666_, new_n1667_, new_n1668_, new_n1669_,
    new_n1670_, new_n1671_, new_n1672_, new_n1673_, new_n1674_, new_n1675_,
    new_n1676_, new_n1677_, new_n1678_, new_n1679_, new_n1680_, new_n1681_,
    new_n1682_, new_n1683_, new_n1684_, new_n1685_, new_n1686_, new_n1687_,
    new_n1688_, new_n1689_, new_n1690_, new_n1691_, new_n1692_, new_n1693_,
    new_n1694_, new_n1695_, new_n1696_, new_n1697_, new_n1698_, new_n1699_,
    new_n1700_, new_n1701_, new_n1702_, new_n1703_, new_n1704_, new_n1705_,
    new_n1706_, new_n1707_, new_n1708_, new_n1709_, new_n1710_, new_n1711_,
    new_n1712_, new_n1713_, new_n1714_, new_n1715_, new_n1716_, new_n1717_,
    new_n1718_, new_n1719_, new_n1720_, new_n1721_, new_n1722_, new_n1723_,
    new_n1724_, new_n1726_, new_n1727_, new_n1728_, new_n1729_, new_n1730_,
    new_n1732_, new_n1733_, new_n1735_, new_n1736_, new_n1738_, new_n1739_,
    new_n1740_, new_n1741_, new_n1743_, new_n1744_, new_n1745_, new_n1746_,
    new_n1747_, new_n1750_, new_n1751_, new_n1752_, new_n1753_, new_n1755_,
    new_n1756_, new_n1757_, new_n1759_, new_n1761_, new_n1763_, new_n1765_,
    new_n1766_, new_n1767_, new_n1768_, new_n1769_, new_n1770_, new_n1771_,
    new_n1772_, new_n1773_, new_n1774_, new_n1775_, new_n1776_, new_n1777_,
    new_n1778_, new_n1779_, new_n1780_, new_n1781_, new_n1782_, new_n1783_,
    new_n1784_, new_n1785_, new_n1786_, new_n1787_, new_n1788_, new_n1789_,
    new_n1790_, new_n1791_, new_n1792_, new_n1793_, new_n1794_, new_n1795_,
    new_n1796_, new_n1797_, new_n1798_, new_n1799_, new_n1800_, new_n1801_,
    new_n1802_, new_n1803_, new_n1804_, new_n1805_, new_n1806_, new_n1807_,
    new_n1808_, new_n1809_, new_n1810_, new_n1811_, new_n1812_, new_n1813_,
    new_n1814_, new_n1815_, new_n1816_, new_n1817_, new_n1818_, new_n1819_,
    new_n1820_, new_n1821_, new_n1822_, new_n1823_, new_n1824_, new_n1825_,
    new_n1826_, new_n1827_, new_n1828_, new_n1829_, new_n1830_, new_n1831_,
    new_n1832_, new_n1833_, new_n1834_, new_n1835_, new_n1836_, new_n1837_,
    new_n1838_, new_n1839_, new_n1840_, new_n1841_, new_n1842_, new_n1843_,
    new_n1844_, new_n1845_, new_n1846_, new_n1847_, new_n1848_, new_n1849_,
    new_n1850_, new_n1851_, new_n1852_, new_n1853_, new_n1855_, new_n1856_,
    new_n1857_, new_n1859_, new_n1861_, new_n1862_, new_n1863_, new_n1864_,
    new_n1866_, new_n1867_, new_n1868_, new_n1869_, new_n1871_, new_n1872_,
    new_n1873_, new_n1874_, new_n1875_, new_n1876_, new_n1877_, new_n1878_,
    new_n1879_, new_n1880_, new_n1881_, new_n1882_, new_n1883_, new_n1884_,
    new_n1885_, new_n1886_, new_n1887_, new_n1888_, new_n1889_, new_n1890_,
    new_n1891_, new_n1892_, new_n1893_, new_n1894_, new_n1895_, new_n1896_,
    new_n1897_, new_n1898_, new_n1899_, new_n1900_, new_n1901_, new_n1902_,
    new_n1903_, new_n1904_, new_n1905_, new_n1906_, new_n1907_, new_n1908_,
    new_n1909_, new_n1910_, new_n1911_, new_n1912_, new_n1913_, new_n1914_,
    new_n1915_, new_n1916_, new_n1917_, new_n1918_, new_n1919_, new_n1920_,
    new_n1921_, new_n1922_, new_n1923_, new_n1924_, new_n1925_, new_n1926_,
    new_n1928_, new_n1930_, new_n1931_, new_n1932_, new_n1933_, new_n1934_,
    new_n1935_, new_n1936_, new_n1937_, new_n1938_, new_n1939_, new_n1940_,
    new_n1941_, new_n1942_, new_n1943_, new_n1944_, new_n1945_, new_n1946_,
    new_n1947_, new_n1948_, new_n1949_, new_n1950_, new_n1951_, new_n1952_,
    new_n1953_, new_n1954_, new_n1955_, new_n1956_, new_n1957_, new_n1958_,
    new_n1959_, new_n1960_, new_n1961_, new_n1962_, new_n1963_, new_n1964_,
    new_n1965_, new_n1966_, new_n1967_, new_n1968_, new_n1969_, new_n1970_,
    new_n1971_, new_n1972_, new_n1973_, new_n1974_, new_n1975_, new_n1976_,
    new_n1977_, new_n1978_, new_n1979_, new_n1980_, new_n1981_, new_n1982_,
    new_n1983_, new_n1984_, new_n1985_, new_n1986_, new_n1987_, new_n1988_,
    new_n1989_, new_n1990_, new_n1991_, new_n1992_, new_n1993_, new_n1994_,
    new_n1995_, new_n1996_, new_n1997_, new_n1998_, new_n1999_, new_n2000_,
    new_n2001_, new_n2002_, new_n2003_, new_n2004_, new_n2005_, new_n2006_,
    new_n2007_, new_n2008_, new_n2009_, new_n2010_, new_n2011_, new_n2012_,
    new_n2013_, new_n2014_, new_n2015_, new_n2016_, new_n2017_, new_n2018_,
    new_n2019_, new_n2020_, new_n2021_, new_n2022_, new_n2023_, new_n2024_,
    new_n2025_, new_n2026_, new_n2027_, new_n2028_, new_n2029_, new_n2030_,
    new_n2031_, new_n2032_, new_n2033_, new_n2034_, new_n2035_, new_n2036_,
    new_n2037_, new_n2038_, new_n2039_, new_n2040_, new_n2041_, new_n2042_,
    new_n2043_, new_n2044_, new_n2045_, new_n2046_, new_n2047_, new_n2048_,
    new_n2049_, new_n2050_, new_n2051_, new_n2052_, new_n2053_, new_n2054_,
    new_n2055_, new_n2056_, new_n2057_, new_n2058_, new_n2059_, new_n2060_,
    new_n2061_, new_n2062_, new_n2063_, new_n2064_, new_n2065_, new_n2066_,
    new_n2067_, new_n2069_, new_n2070_, new_n2071_, new_n2072_, new_n2073_,
    new_n2074_, new_n2075_, new_n2076_, new_n2078_, new_n2079_, new_n2080_,
    new_n2081_, new_n2082_, new_n2083_, new_n2084_, new_n2085_, new_n2086_,
    new_n2087_, new_n2088_, new_n2089_, new_n2091_, new_n2092_, new_n2094_,
    new_n2095_, new_n2096_, new_n2097_, new_n2098_, new_n2099_, new_n2100_,
    new_n2101_, new_n2102_, new_n2103_, new_n2104_, new_n2105_, new_n2106_,
    new_n2107_, new_n2108_, new_n2109_, new_n2110_, new_n2111_, new_n2112_,
    new_n2113_, new_n2114_, new_n2115_, new_n2116_, new_n2117_, new_n2118_,
    new_n2119_, new_n2120_, new_n2121_, new_n2122_, new_n2123_, new_n2124_,
    new_n2125_, new_n2126_, new_n2127_, new_n2128_, new_n2129_, new_n2130_,
    new_n2131_, new_n2132_, new_n2133_, new_n2134_, new_n2135_, new_n2136_,
    new_n2137_, new_n2138_, new_n2139_, new_n2140_, new_n2141_, new_n2142_,
    new_n2143_, new_n2144_, new_n2145_, new_n2146_, new_n2147_, new_n2148_,
    new_n2149_, new_n2150_, new_n2151_, new_n2152_, new_n2153_, new_n2154_,
    new_n2155_, new_n2156_, new_n2157_, new_n2158_, new_n2159_, new_n2160_,
    new_n2161_, new_n2162_, new_n2163_, new_n2164_, new_n2165_, new_n2166_,
    new_n2167_, new_n2168_, new_n2169_, new_n2170_, new_n2171_, new_n2172_,
    new_n2173_, new_n2174_, new_n2175_, new_n2176_, new_n2177_, new_n2178_,
    new_n2179_, new_n2180_, new_n2181_, new_n2182_, new_n2183_, new_n2184_,
    new_n2185_, new_n2186_, new_n2187_, new_n2188_, new_n2189_, new_n2190_,
    new_n2191_, new_n2192_, new_n2193_, new_n2194_, new_n2195_, new_n2196_,
    new_n2197_, new_n2198_, new_n2199_, new_n2200_, new_n2201_, new_n2202_,
    new_n2203_, new_n2204_, new_n2205_, new_n2206_, new_n2207_, new_n2208_,
    new_n2209_, new_n2210_, new_n2211_, new_n2212_, new_n2213_, new_n2214_,
    new_n2215_, new_n2216_, new_n2217_, new_n2218_, new_n2219_, new_n2220_,
    new_n2221_, new_n2222_, new_n2223_, new_n2224_, new_n2225_, new_n2226_,
    new_n2227_, new_n2228_, new_n2229_, new_n2230_, new_n2231_, new_n2232_,
    new_n2233_, new_n2234_, new_n2235_, new_n2236_, new_n2237_, new_n2238_,
    new_n2239_, new_n2240_, new_n2241_, new_n2242_, new_n2243_, new_n2244_,
    new_n2245_, new_n2246_, new_n2247_, new_n2248_, new_n2249_, new_n2250_,
    new_n2251_, new_n2252_, new_n2253_, new_n2254_, new_n2255_, new_n2257_,
    new_n2258_, new_n2260_, new_n2261_, new_n2262_, new_n2263_, new_n2264_,
    new_n2265_, new_n2266_, new_n2267_, new_n2268_, new_n2269_, new_n2270_,
    new_n2271_, new_n2272_, new_n2273_, new_n2274_, new_n2275_, new_n2276_,
    new_n2277_, new_n2278_, new_n2279_, new_n2280_, new_n2281_, new_n2282_,
    new_n2283_, new_n2284_, new_n2285_, new_n2286_, new_n2287_, new_n2288_,
    new_n2289_, new_n2290_, new_n2291_, new_n2292_, new_n2293_, new_n2294_,
    new_n2295_, new_n2296_, new_n2297_, new_n2298_, new_n2299_, new_n2300_,
    new_n2301_, new_n2302_, new_n2303_, new_n2304_, new_n2305_, new_n2306_,
    new_n2307_, new_n2308_, new_n2309_, new_n2310_, new_n2311_, new_n2312_,
    new_n2313_, new_n2314_, new_n2315_, new_n2316_, new_n2317_, new_n2318_,
    new_n2319_, new_n2320_, new_n2321_, new_n2322_, new_n2323_, new_n2324_,
    new_n2325_, new_n2326_, new_n2327_, new_n2328_, new_n2329_, new_n2330_,
    new_n2331_, new_n2332_, new_n2333_, new_n2335_, new_n2336_, new_n2337_,
    new_n2338_, new_n2339_, new_n2340_, new_n2341_, new_n2342_, new_n2343_,
    new_n2344_, new_n2346_, new_n2347_, new_n2348_, new_n2349_, new_n2350_,
    new_n2351_, new_n2352_, new_n2353_, new_n2354_, new_n2355_, new_n2356_,
    new_n2357_, new_n2358_, new_n2359_, new_n2360_, new_n2361_, new_n2362_,
    new_n2363_, new_n2364_, new_n2365_, new_n2366_, new_n2367_, new_n2368_,
    new_n2369_, new_n2370_, new_n2371_, new_n2372_, new_n2373_, new_n2374_,
    new_n2375_, new_n2376_, new_n2377_, new_n2378_, new_n2379_, new_n2380_,
    new_n2381_, new_n2382_, new_n2383_, new_n2384_, new_n2385_, new_n2386_,
    new_n2387_, new_n2388_, new_n2389_, new_n2390_, new_n2391_, new_n2392_,
    new_n2393_, new_n2394_, new_n2395_, new_n2396_, new_n2397_, new_n2398_,
    new_n2399_, new_n2400_, new_n2401_, new_n2402_, new_n2403_, new_n2404_,
    new_n2405_, new_n2406_, new_n2407_, new_n2408_, new_n2409_, new_n2410_,
    new_n2411_, new_n2412_, new_n2413_, new_n2414_, new_n2415_, new_n2416_,
    new_n2417_, new_n2418_, new_n2419_, new_n2420_, new_n2421_, new_n2422_,
    new_n2423_, new_n2424_, new_n2425_, new_n2426_, new_n2427_, new_n2428_,
    new_n2429_, new_n2430_, new_n2431_, new_n2432_, new_n2433_, new_n2434_,
    new_n2435_, new_n2436_, new_n2437_, new_n2438_, new_n2439_, new_n2440_,
    new_n2441_, new_n2442_, new_n2443_, new_n2444_, new_n2445_, new_n2446_,
    new_n2447_, new_n2448_, new_n2449_, new_n2450_, new_n2451_, new_n2452_,
    new_n2453_, new_n2454_, new_n2455_, new_n2456_, new_n2457_, new_n2458_,
    new_n2459_, new_n2460_, new_n2461_, new_n2462_, new_n2463_, new_n2464_,
    new_n2465_, new_n2466_, new_n2467_, new_n2468_, new_n2469_, new_n2470_,
    new_n2471_, new_n2472_, new_n2473_, new_n2474_, new_n2475_, new_n2476_,
    new_n2477_, new_n2478_, new_n2479_, new_n2480_, new_n2481_, new_n2482_,
    new_n2483_, new_n2484_, new_n2485_, new_n2486_, new_n2487_, new_n2488_,
    new_n2489_, new_n2490_, new_n2491_, new_n2492_, new_n2493_, new_n2494_,
    new_n2495_, new_n2496_, new_n2497_, new_n2498_, new_n2499_, new_n2500_,
    new_n2501_, new_n2502_, new_n2503_, new_n2504_, new_n2505_, new_n2506_,
    new_n2507_, new_n2508_, new_n2509_, new_n2510_, new_n2511_, new_n2512_,
    new_n2513_, new_n2514_, new_n2515_, new_n2516_, new_n2517_, new_n2518_,
    new_n2519_, new_n2520_, new_n2521_, new_n2522_, new_n2523_, new_n2524_,
    new_n2525_, new_n2526_, new_n2527_, new_n2528_, new_n2529_, new_n2530_,
    new_n2531_, new_n2532_, new_n2533_, new_n2534_, new_n2535_, new_n2536_,
    new_n2537_, new_n2538_, new_n2539_, new_n2540_, new_n2541_, new_n2542_,
    new_n2543_, new_n2544_, new_n2545_, new_n2546_, new_n2547_, new_n2548_,
    new_n2549_, new_n2550_, new_n2551_, new_n2552_, new_n2553_, new_n2554_,
    new_n2555_, new_n2556_, new_n2557_, new_n2558_, new_n2559_, new_n2560_,
    new_n2561_, new_n2562_, new_n2563_, new_n2564_, new_n2565_, new_n2566_,
    new_n2567_, new_n2568_, new_n2569_, new_n2570_, new_n2571_, new_n2572_,
    new_n2573_, new_n2574_, new_n2575_, new_n2576_, new_n2577_, new_n2578_,
    new_n2579_, new_n2580_, new_n2581_, new_n2582_, new_n2583_, new_n2584_,
    new_n2585_, new_n2586_, new_n2587_, new_n2588_, new_n2589_, new_n2590_,
    new_n2591_, new_n2592_, new_n2593_, new_n2594_, new_n2595_, new_n2596_,
    new_n2597_, new_n2598_, new_n2599_, new_n2600_, new_n2601_, new_n2602_,
    new_n2603_, new_n2604_, new_n2605_, new_n2606_, new_n2607_, new_n2608_,
    new_n2609_, new_n2610_, new_n2611_, new_n2612_, new_n2613_, new_n2614_,
    new_n2615_, new_n2616_, new_n2617_, new_n2618_, new_n2619_, new_n2620_,
    new_n2621_, new_n2622_, new_n2623_, new_n2624_, new_n2625_, new_n2626_,
    new_n2627_, new_n2628_, new_n2629_, new_n2630_, new_n2631_, new_n2632_,
    new_n2633_, new_n2634_, new_n2635_, new_n2636_, new_n2637_, new_n2638_,
    new_n2639_, new_n2640_, new_n2641_, new_n2642_, new_n2643_, new_n2644_,
    new_n2645_, new_n2646_, new_n2647_, new_n2648_, new_n2649_, new_n2650_,
    new_n2651_, new_n2652_, new_n2653_, new_n2654_, new_n2655_, new_n2656_,
    new_n2657_, new_n2658_, new_n2659_, new_n2660_, new_n2661_, new_n2662_,
    new_n2663_, new_n2664_, new_n2665_, new_n2666_, new_n2667_, new_n2668_,
    new_n2669_, new_n2670_, new_n2671_, new_n2672_, new_n2673_, new_n2674_,
    new_n2675_, new_n2676_, new_n2677_, new_n2678_, new_n2679_, new_n2680_,
    new_n2681_, new_n2682_, new_n2683_, new_n2684_, new_n2685_, new_n2686_,
    new_n2687_, new_n2688_, new_n2689_, new_n2690_, new_n2691_, new_n2692_,
    new_n2693_, new_n2694_, new_n2695_, new_n2696_, new_n2697_, new_n2698_,
    new_n2699_, new_n2700_, new_n2701_, new_n2702_, new_n2703_, new_n2704_,
    new_n2705_, new_n2706_, new_n2707_, new_n2708_, new_n2709_, new_n2710_,
    new_n2711_, new_n2712_, new_n2713_, new_n2714_, new_n2715_, new_n2716_,
    new_n2717_, new_n2718_, new_n2719_, new_n2720_, new_n2721_, new_n2722_,
    new_n2723_, new_n2724_, new_n2725_, new_n2726_, new_n2727_, new_n2728_,
    new_n2729_, new_n2730_, new_n2731_, new_n2732_, new_n2733_, new_n2734_,
    new_n2735_, new_n2736_, new_n2737_, new_n2738_, new_n2739_, new_n2740_,
    new_n2741_, new_n2742_, new_n2743_, new_n2744_, new_n2745_, new_n2746_,
    new_n2747_, new_n2748_, new_n2749_, new_n2751_, new_n2752_, new_n2754_,
    new_n2755_, new_n2756_, new_n2757_, new_n2758_, new_n2759_, new_n2760_,
    new_n2761_, new_n2762_, new_n2763_, new_n2764_, new_n2765_, new_n2766_,
    new_n2767_, new_n2768_, new_n2769_, new_n2770_, new_n2771_, new_n2772_,
    new_n2773_, new_n2774_, new_n2775_, new_n2776_, new_n2777_, new_n2778_,
    new_n2779_, new_n2780_, new_n2781_, new_n2782_, new_n2783_, new_n2784_,
    new_n2785_, new_n2786_, new_n2787_, new_n2788_, new_n2789_, new_n2790_,
    new_n2791_, new_n2792_, new_n2793_, new_n2794_, new_n2795_, new_n2796_,
    new_n2797_, new_n2798_, new_n2799_, new_n2800_, new_n2801_, new_n2802_,
    new_n2803_, new_n2804_, new_n2805_, new_n2806_, new_n2807_, new_n2808_,
    new_n2809_, new_n2810_, new_n2811_, new_n2812_, new_n2813_, new_n2814_,
    new_n2815_, new_n2816_, new_n2817_, new_n2818_, new_n2819_, new_n2820_,
    new_n2821_, new_n2822_, new_n2823_, new_n2824_, new_n2825_, new_n2826_,
    new_n2827_, new_n2828_, new_n2829_, new_n2830_, new_n2831_, new_n2832_,
    new_n2833_, new_n2834_, new_n2835_, new_n2836_, new_n2837_, new_n2838_,
    new_n2839_, new_n2840_, new_n2841_, new_n2842_, new_n2843_, new_n2844_,
    new_n2845_, new_n2846_, new_n2847_, new_n2848_, new_n2849_, new_n2850_,
    new_n2851_, new_n2852_, new_n2853_, new_n2854_, new_n2855_, new_n2856_,
    new_n2857_, new_n2858_, new_n2859_, new_n2860_, new_n2861_, new_n2862_,
    new_n2863_, new_n2864_, new_n2865_, new_n2866_, new_n2867_, new_n2868_,
    new_n2869_, new_n2870_, new_n2871_, new_n2872_, new_n2874_, new_n2875_,
    new_n2876_, new_n2877_, new_n2879_, new_n2880_, new_n2882_, new_n2883_,
    new_n2884_, new_n2885_, new_n2886_, new_n2887_, new_n2888_, new_n2889_,
    new_n2890_, new_n2891_, new_n2892_, new_n2893_, new_n2894_, new_n2895_,
    new_n2896_, new_n2897_, new_n2898_, new_n2899_, new_n2900_, new_n2901_,
    new_n2902_, new_n2903_, new_n2904_, new_n2905_, new_n2906_, new_n2907_,
    new_n2908_, new_n2909_, new_n2910_, new_n2911_, new_n2912_, new_n2913_,
    new_n2914_, new_n2915_, new_n2916_, new_n2917_, new_n2918_, new_n2919_,
    new_n2920_, new_n2921_, new_n2922_, new_n2923_, new_n2924_, new_n2925_,
    new_n2926_, new_n2927_, new_n2928_, new_n2929_, new_n2930_, new_n2931_,
    new_n2932_, new_n2933_, new_n2934_, new_n2935_, new_n2936_, new_n2937_,
    new_n2938_, new_n2939_, new_n2940_, new_n2941_, new_n2942_, new_n2943_,
    new_n2944_, new_n2945_, new_n2946_, new_n2947_, new_n2948_, new_n2949_,
    new_n2950_, new_n2951_, new_n2952_, new_n2953_, new_n2954_, new_n2955_,
    new_n2956_, new_n2957_, new_n2958_, new_n2959_, new_n2960_, new_n2961_,
    new_n2962_, new_n2963_, new_n2964_, new_n2965_, new_n2966_, new_n2967_,
    new_n2968_, new_n2969_, new_n2970_, new_n2971_, new_n2972_, new_n2973_,
    new_n2974_, new_n2975_, new_n2976_, new_n2977_, new_n2978_, new_n2979_,
    new_n2980_, new_n2981_, new_n2982_, new_n2983_, new_n2984_, new_n2985_,
    new_n2986_, new_n2987_, new_n2988_, new_n2989_, new_n2990_, new_n2991_,
    new_n2992_, new_n2993_, new_n2994_, new_n2995_, new_n2996_, new_n2997_,
    new_n2998_, new_n2999_, new_n3000_, new_n3001_, new_n3002_, new_n3003_,
    new_n3004_, new_n3005_, new_n3007_, new_n3008_, new_n3010_, new_n3011_,
    new_n3012_, new_n3013_, new_n3014_, new_n3015_, new_n3016_, new_n3017_,
    new_n3018_, new_n3019_, new_n3020_, new_n3021_, new_n3022_, new_n3023_,
    new_n3024_, new_n3025_, new_n3026_, new_n3027_, new_n3028_, new_n3029_,
    new_n3030_, new_n3031_, new_n3032_, new_n3033_, new_n3034_, new_n3035_,
    new_n3036_, new_n3037_, new_n3038_, new_n3039_, new_n3040_, new_n3041_,
    new_n3042_, new_n3043_, new_n3044_, new_n3045_, new_n3046_, new_n3047_,
    new_n3048_, new_n3049_, new_n3050_, new_n3051_, new_n3052_, new_n3053_,
    new_n3054_, new_n3055_, new_n3056_, new_n3057_, new_n3058_, new_n3059_,
    new_n3060_, new_n3061_, new_n3062_, new_n3063_, new_n3064_, new_n3065_,
    new_n3066_, new_n3067_, new_n3068_, new_n3069_, new_n3070_, new_n3071_,
    new_n3072_, new_n3073_, new_n3074_, new_n3075_, new_n3076_, new_n3077_,
    new_n3078_, new_n3079_, new_n3080_, new_n3081_, new_n3082_, new_n3083_,
    new_n3084_, new_n3085_, new_n3086_, new_n3087_, new_n3088_, new_n3089_,
    new_n3090_, new_n3091_, new_n3092_, new_n3093_, new_n3094_, new_n3095_,
    new_n3096_, new_n3097_, new_n3098_, new_n3099_, new_n3100_, new_n3101_,
    new_n3102_, new_n3103_, new_n3104_, new_n3105_, new_n3106_, new_n3107_,
    new_n3108_, new_n3109_, new_n3110_, new_n3111_, new_n3112_, new_n3113_,
    new_n3114_, new_n3115_, new_n3116_, new_n3117_, new_n3118_, new_n3119_,
    new_n3120_, new_n3121_, new_n3122_, new_n3123_, new_n3124_, new_n3125_,
    new_n3126_, new_n3127_, new_n3129_, new_n3130_, new_n3131_, new_n3132_,
    new_n3133_, new_n3134_, new_n3136_, new_n3137_, new_n3138_, new_n3140_,
    new_n3141_, new_n3142_, new_n3143_, new_n3144_, new_n3145_, new_n3146_,
    new_n3147_, new_n3149_, new_n3151_, new_n3152_, new_n3153_, new_n3154_,
    new_n3155_, new_n3156_, new_n3157_, new_n3158_, new_n3159_, new_n3161_,
    new_n3162_, new_n3164_, new_n3165_, new_n3166_, new_n3167_, new_n3168_,
    new_n3169_, new_n3170_, new_n3171_, new_n3173_, new_n3174_, new_n3175_,
    new_n3176_, new_n3177_, new_n3178_, new_n3179_, new_n3180_, new_n3182_,
    new_n3183_, new_n3184_, new_n3185_, new_n3187_, new_n3188_, new_n3189_,
    new_n3190_, new_n3191_, new_n3192_, new_n3193_, new_n3194_, new_n3195_,
    new_n3196_, new_n3198_, new_n3199_, new_n3201_, new_n3202_, new_n3203_,
    new_n3204_, new_n3206_, new_n3207_, new_n3208_, new_n3209_, new_n3211_,
    new_n3212_, new_n3213_, new_n3214_, new_n3215_, new_n3216_, new_n3217_,
    new_n3218_, new_n3220_, new_n3221_, new_n3222_, new_n3223_, new_n3224_,
    new_n3225_, new_n3226_, new_n3227_, new_n3228_, new_n3229_, new_n3230_,
    new_n3231_, new_n3232_, new_n3233_, new_n3234_, new_n3235_, new_n3236_,
    new_n3237_, new_n3238_, new_n3239_, new_n3240_, new_n3241_, new_n3242_,
    new_n3243_, new_n3244_, new_n3245_, new_n3246_, new_n3247_, new_n3248_,
    new_n3249_, new_n3250_, new_n3251_, new_n3252_, new_n3253_, new_n3254_,
    new_n3255_, new_n3256_, new_n3257_, new_n3258_, new_n3259_, new_n3260_,
    new_n3261_, new_n3262_, new_n3263_, new_n3264_, new_n3265_, new_n3266_,
    new_n3267_, new_n3268_, new_n3269_, new_n3270_, new_n3271_, new_n3272_,
    new_n3273_, new_n3274_, new_n3275_, new_n3276_, new_n3277_, new_n3278_,
    new_n3279_, new_n3280_, new_n3281_, new_n3282_, new_n3283_, new_n3284_,
    new_n3285_, new_n3286_, new_n3287_, new_n3288_, new_n3289_, new_n3290_,
    new_n3291_, new_n3292_, new_n3293_, new_n3294_, new_n3295_, new_n3296_,
    new_n3297_, new_n3298_, new_n3299_, new_n3300_, new_n3301_, new_n3302_,
    new_n3303_, new_n3304_, new_n3305_, new_n3306_, new_n3307_, new_n3308_,
    new_n3309_, new_n3310_, new_n3311_, new_n3312_, new_n3313_, new_n3314_,
    new_n3316_, new_n3317_, new_n3318_, new_n3319_, new_n3320_, new_n3321_,
    new_n3322_, new_n3326_, new_n3327_, new_n3328_, new_n3329_, new_n3330_,
    new_n3331_, new_n3332_, new_n3333_, new_n3335_, new_n3336_, new_n3337_,
    new_n3338_, new_n3339_, new_n3340_, new_n3341_, new_n3342_, new_n3344_,
    new_n3345_, new_n3346_, new_n3347_, new_n3348_, new_n3349_, new_n3350_,
    new_n3351_, new_n3352_, new_n3353_, new_n3354_, new_n3355_, new_n3356_,
    new_n3357_, new_n3358_, new_n3359_, new_n3360_, new_n3361_, new_n3362_,
    new_n3363_, new_n3364_, new_n3365_, new_n3366_, new_n3367_, new_n3368_,
    new_n3369_, new_n3370_, new_n3371_, new_n3372_, new_n3373_, new_n3374_,
    new_n3375_, new_n3376_, new_n3377_, new_n3378_, new_n3379_, new_n3380_,
    new_n3381_, new_n3382_, new_n3383_, new_n3384_, new_n3385_, new_n3386_,
    new_n3387_, new_n3388_, new_n3389_, new_n3390_, new_n3391_, new_n3392_,
    new_n3393_, new_n3394_, new_n3395_, new_n3396_, new_n3397_, new_n3398_,
    new_n3399_, new_n3400_, new_n3401_, new_n3402_, new_n3403_, new_n3404_,
    new_n3405_, new_n3406_, new_n3407_, new_n3408_, new_n3409_, new_n3410_,
    new_n3411_, new_n3412_, new_n3413_, new_n3414_, new_n3415_, new_n3416_,
    new_n3417_, new_n3419_, new_n3420_, new_n3421_, new_n3422_, new_n3423_,
    new_n3424_, new_n3425_, new_n3427_, new_n3428_, new_n3429_, new_n3430_,
    new_n3431_, new_n3432_, new_n3433_, new_n3434_, new_n3435_, new_n3436_,
    new_n3437_, new_n3439_, new_n3440_, new_n3441_, new_n3442_, new_n3444_,
    new_n3445_, new_n3446_, new_n3447_, new_n3448_, new_n3449_, new_n3450_,
    new_n3451_, new_n3453_, new_n3455_, new_n3456_, new_n3457_, new_n3458_,
    new_n3459_, new_n3460_, new_n3461_, new_n3462_, new_n3463_, new_n3464_,
    new_n3465_, new_n3466_, new_n3467_, new_n3468_, new_n3469_, new_n3470_,
    new_n3471_, new_n3472_, new_n3473_, new_n3474_, new_n3475_, new_n3476_,
    new_n3477_, new_n3478_, new_n3479_, new_n3480_, new_n3481_, new_n3482_,
    new_n3483_, new_n3484_, new_n3485_, new_n3486_, new_n3487_, new_n3488_,
    new_n3489_, new_n3490_, new_n3491_, new_n3492_, new_n3493_, new_n3494_,
    new_n3495_, new_n3496_, new_n3497_, new_n3498_, new_n3499_, new_n3500_,
    new_n3501_, new_n3502_, new_n3503_, new_n3504_, new_n3505_, new_n3506_,
    new_n3507_, new_n3508_, new_n3509_, new_n3510_, new_n3511_, new_n3512_,
    new_n3513_, new_n3514_, new_n3515_, new_n3516_, new_n3517_, new_n3518_,
    new_n3519_, new_n3520_, new_n3521_, new_n3522_, new_n3523_, new_n3524_,
    new_n3525_, new_n3526_, new_n3527_, new_n3528_, new_n3529_, new_n3530_,
    new_n3531_, new_n3532_, new_n3533_, new_n3534_, new_n3535_, new_n3536_,
    new_n3537_, new_n3538_, new_n3539_, new_n3540_, new_n3541_, new_n3542_,
    new_n3543_, new_n3544_, new_n3546_, new_n3547_, new_n3549_, new_n3550_,
    new_n3551_, new_n3553_, new_n3554_, new_n3555_, new_n3556_, new_n3557_,
    new_n3558_, new_n3559_, new_n3560_, new_n3563_, new_n3564_, new_n3565_,
    new_n3567_, new_n3568_, new_n3569_, new_n3570_, new_n3572_, new_n3574_,
    new_n3575_, new_n3576_, new_n3577_, new_n3578_, new_n3580_, new_n3581_,
    new_n3582_, new_n3584_, new_n3585_, new_n3586_, new_n3587_;
  assign new_n608_ = ~\1_n839  & ~\1_n1022 ;
  assign new_n609_ = \1_n975  & new_n608_;
  assign new_n610_ = \1_n1352  & ~new_n609_;
  assign new_n611_ = ~\1_n688  & ~\1_n866 ;
  assign new_n612_ = ~\1_n95  & ~\1_n688 ;
  assign new_n613_ = new_n611_ & new_n612_;
  assign new_n614_ = \1_n336  & \1_n384 ;
  assign new_n615_ = \1_n839  & \1_n1022 ;
  assign new_n616_ = \1_n975  & ~new_n615_;
  assign new_n617_ = ~\1_n1352  & new_n616_;
  assign new_n618_ = ~new_n614_ & ~new_n617_;
  assign new_n619_ = ~new_n613_ & new_n618_;
  assign new_n620_ = ~new_n612_ & ~new_n617_;
  assign new_n621_ = ~new_n611_ & new_n620_;
  assign new_n622_ = ~new_n618_ & ~new_n621_;
  assign new_n623_ = \1_n936  & ~new_n614_;
  assign new_n624_ = ~\1_n688  & ~new_n614_;
  assign new_n625_ = ~new_n623_ & ~new_n624_;
  assign new_n626_ = ~\1_n688  & ~\1_n804 ;
  assign new_n627_ = ~new_n625_ & ~new_n626_;
  assign new_n628_ = ~\1_n667  & ~\1_n688 ;
  assign new_n629_ = \1_n928  & ~new_n614_;
  assign new_n630_ = ~new_n624_ & ~new_n629_;
  assign new_n631_ = ~new_n628_ & ~new_n630_;
  assign new_n632_ = \1_n281  & ~new_n614_;
  assign new_n633_ = ~new_n624_ & ~new_n632_;
  assign new_n634_ = \1_n640  & ~\1_n688 ;
  assign new_n635_ = ~\1_n393  & \1_n688 ;
  assign new_n636_ = ~new_n634_ & ~new_n635_;
  assign new_n637_ = ~new_n633_ & ~new_n636_;
  assign new_n638_ = \1_n284  & ~new_n614_;
  assign new_n639_ = ~new_n624_ & ~new_n638_;
  assign new_n640_ = ~\1_n519  & ~\1_n688 ;
  assign new_n641_ = ~new_n639_ & ~new_n640_;
  assign new_n642_ = ~new_n637_ & ~new_n641_;
  assign new_n643_ = \1_n688  & \1_n1044 ;
  assign new_n644_ = ~\1_n688  & \1_n695 ;
  assign new_n645_ = ~new_n643_ & ~new_n644_;
  assign new_n646_ = ~\1_n644  & \1_n688 ;
  assign new_n647_ = ~\1_n688  & \1_n1326 ;
  assign new_n648_ = ~new_n646_ & ~new_n647_;
  assign new_n649_ = ~new_n645_ & ~new_n648_;
  assign new_n650_ = \1_n196  & ~\1_n688 ;
  assign new_n651_ = \1_n688  & \1_n806 ;
  assign new_n652_ = ~new_n650_ & ~new_n651_;
  assign new_n653_ = ~\1_n332  & \1_n688 ;
  assign new_n654_ = ~\1_n688  & \1_n1091 ;
  assign new_n655_ = ~new_n653_ & ~new_n654_;
  assign new_n656_ = ~new_n652_ & new_n655_;
  assign new_n657_ = new_n652_ & ~new_n655_;
  assign new_n658_ = ~new_n656_ & ~new_n657_;
  assign new_n659_ = \1_n246  & ~\1_n688 ;
  assign new_n660_ = ~\1_n231  & \1_n688 ;
  assign new_n661_ = ~new_n659_ & ~new_n660_;
  assign new_n662_ = \1_n771  & ~new_n614_;
  assign new_n663_ = ~new_n624_ & ~new_n662_;
  assign new_n664_ = new_n661_ & ~new_n663_;
  assign new_n665_ = ~new_n661_ & new_n663_;
  assign new_n666_ = ~new_n664_ & ~new_n665_;
  assign new_n667_ = ~new_n658_ & ~new_n666_;
  assign new_n668_ = \1_n688  & \1_n745 ;
  assign new_n669_ = ~\1_n688  & \1_n825 ;
  assign new_n670_ = ~new_n668_ & ~new_n669_;
  assign new_n671_ = \1_n688  & ~\1_n716 ;
  assign new_n672_ = \1_n245  & ~\1_n688 ;
  assign new_n673_ = ~new_n671_ & ~new_n672_;
  assign new_n674_ = new_n670_ & new_n673_;
  assign new_n675_ = ~new_n670_ & ~new_n673_;
  assign new_n676_ = ~new_n674_ & ~new_n675_;
  assign new_n677_ = new_n667_ & new_n676_;
  assign new_n678_ = new_n649_ & new_n677_;
  assign new_n679_ = new_n661_ & new_n663_;
  assign new_n680_ = ~new_n655_ & ~new_n679_;
  assign new_n681_ = ~new_n652_ & new_n680_;
  assign new_n682_ = ~new_n661_ & ~new_n663_;
  assign new_n683_ = new_n667_ & ~new_n673_;
  assign new_n684_ = ~new_n670_ & new_n683_;
  assign new_n685_ = ~new_n682_ & ~new_n684_;
  assign new_n686_ = new_n645_ & new_n648_;
  assign new_n687_ = ~new_n649_ & ~new_n686_;
  assign new_n688_ = \1_n423  & ~\1_n688 ;
  assign new_n689_ = ~\1_n449  & \1_n688 ;
  assign new_n690_ = ~new_n688_ & ~new_n689_;
  assign new_n691_ = new_n687_ & ~new_n690_;
  assign new_n692_ = new_n677_ & new_n691_;
  assign new_n693_ = \1_n610  & \1_n688 ;
  assign new_n694_ = ~\1_n688  & \1_n841 ;
  assign new_n695_ = ~new_n693_ & ~new_n694_;
  assign new_n696_ = new_n692_ & ~new_n695_;
  assign new_n697_ = new_n685_ & ~new_n696_;
  assign new_n698_ = ~new_n681_ & new_n697_;
  assign new_n699_ = ~new_n678_ & new_n698_;
  assign new_n700_ = new_n625_ & new_n626_;
  assign new_n701_ = new_n628_ & new_n630_;
  assign new_n702_ = ~new_n631_ & ~new_n701_;
  assign new_n703_ = ~new_n700_ & new_n702_;
  assign new_n704_ = ~new_n627_ & new_n703_;
  assign new_n705_ = new_n633_ & new_n636_;
  assign new_n706_ = new_n639_ & new_n640_;
  assign new_n707_ = ~new_n705_ & ~new_n706_;
  assign new_n708_ = new_n704_ & new_n707_;
  assign new_n709_ = new_n642_ & new_n708_;
  assign new_n710_ = ~new_n699_ & new_n709_;
  assign new_n711_ = new_n642_ & ~new_n710_;
  assign new_n712_ = ~new_n631_ & new_n711_;
  assign new_n713_ = ~new_n627_ & new_n712_;
  assign new_n714_ = ~new_n622_ & ~new_n713_;
  assign new_n715_ = ~new_n619_ & ~new_n714_;
  assign new_n716_ = ~new_n610_ & new_n715_;
  assign new_n717_ = \1_n500  & ~\1_n688 ;
  assign new_n718_ = \1_n688  & \1_n1073 ;
  assign new_n719_ = ~new_n717_ & ~new_n718_;
  assign new_n720_ = \1_n688  & ~\1_n1311 ;
  assign new_n721_ = \1_n258  & ~\1_n688 ;
  assign new_n722_ = ~new_n720_ & ~new_n721_;
  assign new_n723_ = \1_n688  & \1_n1097 ;
  assign new_n724_ = \1_n200  & ~\1_n688 ;
  assign new_n725_ = ~new_n723_ & ~new_n724_;
  assign new_n726_ = ~\1_n571  & \1_n688 ;
  assign new_n727_ = ~\1_n688  & \1_n1131 ;
  assign new_n728_ = ~new_n726_ & ~new_n727_;
  assign new_n729_ = new_n725_ & new_n728_;
  assign new_n730_ = ~new_n725_ & ~new_n728_;
  assign new_n731_ = ~new_n729_ & ~new_n730_;
  assign new_n732_ = \1_n366  & \1_n688 ;
  assign new_n733_ = ~\1_n688  & \1_n879 ;
  assign new_n734_ = ~new_n732_ & ~new_n733_;
  assign new_n735_ = ~\1_n301  & \1_n688 ;
  assign new_n736_ = ~\1_n688  & \1_n1005 ;
  assign new_n737_ = ~new_n735_ & ~new_n736_;
  assign new_n738_ = new_n734_ & new_n737_;
  assign new_n739_ = ~new_n734_ & ~new_n737_;
  assign new_n740_ = ~new_n738_ & ~new_n739_;
  assign new_n741_ = ~\1_n688  & \1_n1069 ;
  assign new_n742_ = \1_n650  & \1_n688 ;
  assign new_n743_ = ~new_n741_ & ~new_n742_;
  assign new_n744_ = ~\1_n688  & \1_n1279 ;
  assign new_n745_ = \1_n688  & ~\1_n1321 ;
  assign new_n746_ = ~new_n744_ & ~new_n745_;
  assign new_n747_ = new_n743_ & ~new_n746_;
  assign new_n748_ = ~new_n743_ & new_n746_;
  assign new_n749_ = ~new_n747_ & ~new_n748_;
  assign new_n750_ = new_n740_ & ~new_n749_;
  assign new_n751_ = \1_n323  & ~\1_n688 ;
  assign new_n752_ = \1_n98  & \1_n688 ;
  assign new_n753_ = ~new_n751_ & ~new_n752_;
  assign new_n754_ = \1_n688  & ~\1_n1198 ;
  assign new_n755_ = \1_n262  & ~\1_n688 ;
  assign new_n756_ = ~new_n754_ & ~new_n755_;
  assign new_n757_ = new_n753_ & new_n756_;
  assign new_n758_ = ~new_n753_ & ~new_n756_;
  assign new_n759_ = ~new_n757_ & ~new_n758_;
  assign new_n760_ = \1_n441  & ~\1_n688 ;
  assign new_n761_ = ~\1_n104  & \1_n688 ;
  assign new_n762_ = ~new_n760_ & ~new_n761_;
  assign new_n763_ = \1_n688  & \1_n1064 ;
  assign new_n764_ = \1_n536  & ~\1_n688 ;
  assign new_n765_ = ~new_n763_ & ~new_n764_;
  assign new_n766_ = ~new_n762_ & ~new_n765_;
  assign new_n767_ = new_n762_ & new_n765_;
  assign new_n768_ = \1_n688  & \1_n1098 ;
  assign new_n769_ = ~\1_n688  & \1_n1229 ;
  assign new_n770_ = ~new_n768_ & ~new_n769_;
  assign new_n771_ = ~\1_n107  & \1_n688 ;
  assign new_n772_ = \1_n208  & ~\1_n688 ;
  assign new_n773_ = ~new_n771_ & ~new_n772_;
  assign new_n774_ = new_n770_ & new_n773_;
  assign new_n775_ = ~new_n770_ & ~new_n773_;
  assign new_n776_ = ~new_n774_ & ~new_n775_;
  assign new_n777_ = \1_n688  & \1_n823 ;
  assign new_n778_ = \1_n631  & ~\1_n688 ;
  assign new_n779_ = ~new_n777_ & ~new_n778_;
  assign new_n780_ = \1_n77  & ~\1_n688 ;
  assign new_n781_ = ~\1_n589  & \1_n688 ;
  assign new_n782_ = ~new_n780_ & ~new_n781_;
  assign new_n783_ = new_n779_ & ~new_n782_;
  assign new_n784_ = ~new_n779_ & new_n782_;
  assign new_n785_ = ~new_n783_ & ~new_n784_;
  assign new_n786_ = new_n776_ & ~new_n785_;
  assign new_n787_ = \1_n657  & \1_n688 ;
  assign new_n788_ = ~\1_n688  & \1_n1132 ;
  assign new_n789_ = ~new_n787_ & ~new_n788_;
  assign new_n790_ = new_n786_ & ~new_n789_;
  assign new_n791_ = \1_n260  & ~\1_n688 ;
  assign new_n792_ = ~\1_n360  & \1_n688 ;
  assign new_n793_ = ~new_n791_ & ~new_n792_;
  assign new_n794_ = new_n786_ & ~new_n793_;
  assign new_n795_ = ~new_n790_ & ~new_n794_;
  assign new_n796_ = ~new_n767_ & ~new_n795_;
  assign new_n797_ = ~new_n766_ & new_n796_;
  assign new_n798_ = new_n759_ & new_n797_;
  assign new_n799_ = new_n750_ & new_n798_;
  assign new_n800_ = new_n731_ & new_n799_;
  assign new_n801_ = ~new_n722_ & new_n800_;
  assign new_n802_ = ~new_n719_ & new_n801_;
  assign new_n803_ = ~new_n789_ & new_n794_;
  assign new_n804_ = ~new_n779_ & ~new_n782_;
  assign new_n805_ = new_n766_ & ~new_n795_;
  assign new_n806_ = ~new_n804_ & ~new_n805_;
  assign new_n807_ = ~new_n803_ & new_n806_;
  assign new_n808_ = new_n779_ & new_n782_;
  assign new_n809_ = ~new_n773_ & ~new_n808_;
  assign new_n810_ = ~new_n770_ & new_n809_;
  assign new_n811_ = ~new_n743_ & ~new_n746_;
  assign new_n812_ = new_n743_ & new_n746_;
  assign new_n813_ = ~new_n737_ & ~new_n812_;
  assign new_n814_ = ~new_n734_ & new_n813_;
  assign new_n815_ = new_n731_ & new_n758_;
  assign new_n816_ = ~new_n730_ & ~new_n815_;
  assign new_n817_ = new_n750_ & ~new_n816_;
  assign new_n818_ = ~new_n814_ & ~new_n817_;
  assign new_n819_ = ~new_n811_ & new_n818_;
  assign new_n820_ = new_n797_ & ~new_n819_;
  assign new_n821_ = ~new_n810_ & ~new_n820_;
  assign new_n822_ = new_n807_ & new_n821_;
  assign new_n823_ = ~new_n719_ & new_n800_;
  assign new_n824_ = ~new_n801_ & ~new_n823_;
  assign new_n825_ = \1_n688  & \1_n1146 ;
  assign new_n826_ = ~\1_n688  & \1_n863 ;
  assign new_n827_ = ~new_n825_ & ~new_n826_;
  assign new_n828_ = ~\1_n688  & \1_n774 ;
  assign new_n829_ = \1_n688  & ~\1_n997 ;
  assign new_n830_ = ~new_n828_ & ~new_n829_;
  assign new_n831_ = ~new_n827_ & ~new_n830_;
  assign new_n832_ = \1_n688  & \1_n1140 ;
  assign new_n833_ = ~\1_n688  & \1_n893 ;
  assign new_n834_ = ~new_n832_ & ~new_n833_;
  assign new_n835_ = \1_n688  & ~\1_n1308 ;
  assign new_n836_ = ~\1_n688  & \1_n833 ;
  assign new_n837_ = ~new_n835_ & ~new_n836_;
  assign new_n838_ = ~new_n834_ & new_n837_;
  assign new_n839_ = new_n834_ & ~new_n837_;
  assign new_n840_ = ~new_n838_ & ~new_n839_;
  assign new_n841_ = new_n827_ & new_n830_;
  assign new_n842_ = ~new_n831_ & ~new_n841_;
  assign new_n843_ = ~new_n840_ & new_n842_;
  assign new_n844_ = \1_n688  & \1_n1080 ;
  assign new_n845_ = ~\1_n688  & \1_n1077 ;
  assign new_n846_ = ~new_n844_ & ~new_n845_;
  assign new_n847_ = ~\1_n688  & \1_n1164 ;
  assign new_n848_ = ~\1_n38  & \1_n688 ;
  assign new_n849_ = ~new_n847_ & ~new_n848_;
  assign new_n850_ = ~new_n846_ & ~new_n849_;
  assign new_n851_ = ~new_n846_ & new_n849_;
  assign new_n852_ = new_n846_ & ~new_n849_;
  assign new_n853_ = ~new_n851_ & ~new_n852_;
  assign new_n854_ = \1_n431  & \1_n688 ;
  assign new_n855_ = ~\1_n688  & \1_n741 ;
  assign new_n856_ = ~new_n854_ & ~new_n855_;
  assign new_n857_ = \1_n540  & ~\1_n688 ;
  assign new_n858_ = ~\1_n36  & \1_n688 ;
  assign new_n859_ = ~new_n857_ & ~new_n858_;
  assign new_n860_ = ~new_n856_ & ~new_n859_;
  assign new_n861_ = ~new_n853_ & new_n860_;
  assign new_n862_ = ~new_n850_ & ~new_n861_;
  assign new_n863_ = new_n843_ & ~new_n862_;
  assign new_n864_ = ~new_n831_ & ~new_n863_;
  assign new_n865_ = ~new_n837_ & ~new_n841_;
  assign new_n866_ = ~new_n834_ & new_n865_;
  assign new_n867_ = new_n864_ & ~new_n866_;
  assign new_n868_ = ~\1_n688  & \1_n1120 ;
  assign new_n869_ = ~\1_n138  & \1_n688 ;
  assign new_n870_ = ~new_n868_ & ~new_n869_;
  assign new_n871_ = \1_n305  & \1_n688 ;
  assign new_n872_ = ~\1_n688  & \1_n845 ;
  assign new_n873_ = ~new_n871_ & ~new_n872_;
  assign new_n874_ = ~new_n870_ & ~new_n873_;
  assign new_n875_ = new_n870_ & new_n873_;
  assign new_n876_ = \1_n364  & \1_n688 ;
  assign new_n877_ = \1_n221  & ~\1_n688 ;
  assign new_n878_ = ~new_n876_ & ~new_n877_;
  assign new_n879_ = ~\1_n45  & \1_n688 ;
  assign new_n880_ = \1_n510  & ~\1_n688 ;
  assign new_n881_ = ~new_n879_ & ~new_n880_;
  assign new_n882_ = new_n878_ & new_n881_;
  assign new_n883_ = ~new_n878_ & ~new_n881_;
  assign new_n884_ = ~new_n882_ & ~new_n883_;
  assign new_n885_ = \1_n688  & \1_n1219 ;
  assign new_n886_ = ~\1_n688  & \1_n1072 ;
  assign new_n887_ = ~new_n885_ & ~new_n886_;
  assign new_n888_ = ~\1_n688  & \1_n929 ;
  assign new_n889_ = \1_n688  & ~\1_n1035 ;
  assign new_n890_ = ~new_n888_ & ~new_n889_;
  assign new_n891_ = ~new_n887_ & ~new_n890_;
  assign new_n892_ = new_n887_ & new_n890_;
  assign new_n893_ = ~new_n891_ & ~new_n892_;
  assign new_n894_ = new_n884_ & new_n893_;
  assign new_n895_ = \1_n688  & \1_n714 ;
  assign new_n896_ = ~\1_n688  & \1_n1151 ;
  assign new_n897_ = ~new_n895_ & ~new_n896_;
  assign new_n898_ = new_n894_ & ~new_n897_;
  assign new_n899_ = ~\1_n688  & \1_n1141 ;
  assign new_n900_ = \1_n688  & ~\1_n1081 ;
  assign new_n901_ = ~new_n899_ & ~new_n900_;
  assign new_n902_ = new_n894_ & ~new_n901_;
  assign new_n903_ = ~new_n898_ & ~new_n902_;
  assign new_n904_ = ~new_n875_ & ~new_n903_;
  assign new_n905_ = ~new_n874_ & new_n904_;
  assign new_n906_ = ~new_n867_ & new_n905_;
  assign new_n907_ = ~new_n881_ & ~new_n892_;
  assign new_n908_ = ~new_n878_ & new_n907_;
  assign new_n909_ = ~new_n897_ & new_n902_;
  assign new_n910_ = new_n874_ & ~new_n903_;
  assign new_n911_ = ~new_n891_ & ~new_n910_;
  assign new_n912_ = ~new_n909_ & new_n911_;
  assign new_n913_ = ~new_n908_ & new_n912_;
  assign new_n914_ = ~new_n906_ & new_n913_;
  assign new_n915_ = new_n856_ & ~new_n859_;
  assign new_n916_ = ~new_n856_ & new_n859_;
  assign new_n917_ = ~new_n915_ & ~new_n916_;
  assign new_n918_ = new_n905_ & ~new_n917_;
  assign new_n919_ = new_n843_ & new_n918_;
  assign new_n920_ = ~new_n853_ & new_n919_;
  assign new_n921_ = ~\1_n685  & ~\1_n688 ;
  assign new_n922_ = ~\1_n532  & ~new_n921_;
  assign new_n923_ = \1_n685  & ~\1_n688 ;
  assign new_n924_ = \1_n532  & ~new_n923_;
  assign new_n925_ = \1_n857  & ~new_n924_;
  assign new_n926_ = ~new_n922_ & ~new_n925_;
  assign new_n927_ = new_n920_ & ~new_n926_;
  assign new_n928_ = new_n914_ & ~new_n927_;
  assign new_n929_ = ~new_n824_ & ~new_n928_;
  assign new_n930_ = new_n822_ & ~new_n929_;
  assign \1_n456  = new_n802_ | ~new_n930_;
  assign new_n932_ = new_n687_ & ~new_n695_;
  assign new_n933_ = new_n677_ & new_n932_;
  assign new_n934_ = ~new_n692_ & ~new_n933_;
  assign new_n935_ = ~new_n622_ & ~new_n934_;
  assign new_n936_ = \1_n456  & new_n935_;
  assign new_n937_ = new_n709_ & new_n936_;
  assign \1_n1259  = ~new_n716_ | new_n937_;
  assign new_n939_ = \1_n310  & \1_n688 ;
  assign new_n940_ = ~new_n669_ & ~new_n939_;
  assign new_n941_ = \1_n716  & new_n940_;
  assign new_n942_ = ~\1_n716  & ~new_n940_;
  assign new_n943_ = ~new_n941_ & ~new_n942_;
  assign new_n944_ = ~new_n644_ & ~new_n939_;
  assign new_n945_ = \1_n644  & new_n944_;
  assign new_n946_ = ~\1_n644  & ~new_n944_;
  assign new_n947_ = ~new_n945_ & ~new_n946_;
  assign new_n948_ = ~new_n694_ & ~new_n939_;
  assign new_n949_ = ~\1_n449  & ~new_n948_;
  assign new_n950_ = new_n947_ & new_n949_;
  assign new_n951_ = ~new_n946_ & ~new_n950_;
  assign new_n952_ = \1_n449  & new_n948_;
  assign new_n953_ = ~new_n949_ & ~new_n952_;
  assign new_n954_ = new_n947_ & new_n953_;
  assign new_n955_ = new_n951_ & ~new_n954_;
  assign new_n956_ = \1_n688  & \1_n1180 ;
  assign new_n957_ = ~new_n778_ & ~new_n956_;
  assign new_n958_ = ~\1_n589  & ~new_n957_;
  assign new_n959_ = \1_n589  & new_n957_;
  assign new_n960_ = ~new_n958_ & ~new_n959_;
  assign new_n961_ = ~\1_n421  & \1_n688 ;
  assign new_n962_ = ~\1_n688  & ~\1_n1229 ;
  assign new_n963_ = ~new_n961_ & ~new_n962_;
  assign new_n964_ = \1_n107  & ~new_n963_;
  assign new_n965_ = ~\1_n107  & new_n963_;
  assign new_n966_ = ~new_n964_ & ~new_n965_;
  assign new_n967_ = \1_n0  & \1_n688 ;
  assign new_n968_ = ~new_n788_ & ~new_n967_;
  assign new_n969_ = \1_n360  & new_n968_;
  assign new_n970_ = ~\1_n360  & ~new_n968_;
  assign new_n971_ = ~new_n969_ & ~new_n970_;
  assign new_n972_ = \1_n688  & \1_n1273 ;
  assign new_n973_ = ~new_n764_ & ~new_n972_;
  assign new_n974_ = ~\1_n104  & ~new_n973_;
  assign new_n975_ = new_n971_ & new_n974_;
  assign new_n976_ = ~new_n970_ & ~new_n975_;
  assign new_n977_ = new_n966_ & ~new_n976_;
  assign new_n978_ = ~new_n965_ & ~new_n977_;
  assign new_n979_ = \1_n104  & new_n973_;
  assign new_n980_ = ~new_n974_ & ~new_n979_;
  assign new_n981_ = new_n971_ & new_n980_;
  assign new_n982_ = new_n966_ & new_n981_;
  assign new_n983_ = new_n978_ & ~new_n982_;
  assign new_n984_ = \1_n688  & \1_n826 ;
  assign new_n985_ = ~new_n741_ & ~new_n984_;
  assign new_n986_ = \1_n1321  & new_n985_;
  assign new_n987_ = ~\1_n1321  & ~new_n985_;
  assign new_n988_ = ~new_n986_ & ~new_n987_;
  assign new_n989_ = \1_n688  & \1_n1045 ;
  assign new_n990_ = ~new_n733_ & ~new_n989_;
  assign new_n991_ = ~\1_n301  & ~new_n990_;
  assign new_n992_ = \1_n688  & \1_n1036 ;
  assign new_n993_ = ~new_n724_ & ~new_n992_;
  assign new_n994_ = ~\1_n571  & ~new_n993_;
  assign new_n995_ = \1_n688  & \1_n901 ;
  assign new_n996_ = ~new_n717_ & ~new_n995_;
  assign new_n997_ = ~\1_n1311  & ~new_n996_;
  assign new_n998_ = \1_n236  & \1_n688 ;
  assign new_n999_ = ~new_n751_ & ~new_n998_;
  assign new_n1000_ = \1_n1198  & new_n999_;
  assign new_n1001_ = ~\1_n1198  & ~new_n999_;
  assign new_n1002_ = ~new_n1000_ & ~new_n1001_;
  assign new_n1003_ = new_n997_ & new_n1002_;
  assign new_n1004_ = ~new_n1001_ & ~new_n1003_;
  assign new_n1005_ = \1_n571  & new_n993_;
  assign new_n1006_ = ~new_n994_ & ~new_n1005_;
  assign new_n1007_ = ~new_n1004_ & new_n1006_;
  assign new_n1008_ = ~new_n994_ & ~new_n1007_;
  assign new_n1009_ = \1_n301  & new_n990_;
  assign new_n1010_ = ~new_n991_ & ~new_n1009_;
  assign new_n1011_ = ~new_n1008_ & new_n1010_;
  assign new_n1012_ = ~new_n991_ & ~new_n1011_;
  assign new_n1013_ = \1_n688  & \1_n1089 ;
  assign new_n1014_ = ~new_n886_ & ~new_n1013_;
  assign new_n1015_ = \1_n1035  & new_n1014_;
  assign new_n1016_ = ~\1_n1035  & ~new_n1014_;
  assign new_n1017_ = ~new_n1015_ & ~new_n1016_;
  assign new_n1018_ = \1_n688  & \1_n1191 ;
  assign new_n1019_ = ~new_n877_ & ~new_n1018_;
  assign new_n1020_ = \1_n45  & new_n1019_;
  assign new_n1021_ = ~\1_n45  & ~new_n1019_;
  assign new_n1022_ = ~new_n1020_ & ~new_n1021_;
  assign new_n1023_ = \1_n688  & \1_n961 ;
  assign new_n1024_ = ~new_n896_ & ~new_n1023_;
  assign new_n1025_ = \1_n1081  & new_n1024_;
  assign new_n1026_ = ~\1_n1081  & ~new_n1024_;
  assign new_n1027_ = ~new_n1025_ & ~new_n1026_;
  assign new_n1028_ = \1_n122  & \1_n688 ;
  assign new_n1029_ = ~new_n872_ & ~new_n1028_;
  assign new_n1030_ = ~\1_n138  & ~new_n1029_;
  assign new_n1031_ = new_n1027_ & new_n1030_;
  assign new_n1032_ = ~new_n1026_ & ~new_n1031_;
  assign new_n1033_ = new_n1022_ & ~new_n1032_;
  assign new_n1034_ = ~new_n1021_ & ~new_n1033_;
  assign new_n1035_ = \1_n138  & new_n1029_;
  assign new_n1036_ = ~new_n1030_ & ~new_n1035_;
  assign new_n1037_ = new_n1027_ & new_n1036_;
  assign new_n1038_ = new_n1022_ & new_n1037_;
  assign new_n1039_ = new_n1034_ & ~new_n1038_;
  assign new_n1040_ = ~new_n826_ & ~new_n1028_;
  assign new_n1041_ = \1_n997  & new_n1040_;
  assign new_n1042_ = ~\1_n997  & ~new_n1040_;
  assign new_n1043_ = ~new_n1041_ & ~new_n1042_;
  assign new_n1044_ = ~new_n833_ & ~new_n1028_;
  assign new_n1045_ = \1_n1308  & new_n1044_;
  assign new_n1046_ = ~\1_n1308  & ~new_n1044_;
  assign new_n1047_ = ~new_n1045_ & ~new_n1046_;
  assign new_n1048_ = \1_n108  & \1_n688 ;
  assign new_n1049_ = ~new_n845_ & ~new_n1048_;
  assign new_n1050_ = \1_n38  & new_n1049_;
  assign new_n1051_ = ~\1_n38  & ~new_n1049_;
  assign new_n1052_ = ~new_n1050_ & ~new_n1051_;
  assign new_n1053_ = \1_n444  & \1_n688 ;
  assign new_n1054_ = ~new_n855_ & ~new_n1053_;
  assign new_n1055_ = \1_n36  & new_n1054_;
  assign new_n1056_ = ~\1_n36  & ~new_n1054_;
  assign new_n1057_ = ~new_n1055_ & ~new_n1056_;
  assign new_n1058_ = ~\1_n268  & new_n923_;
  assign new_n1059_ = new_n1057_ & new_n1058_;
  assign new_n1060_ = ~new_n1056_ & ~new_n1059_;
  assign new_n1061_ = new_n1052_ & ~new_n1060_;
  assign new_n1062_ = ~new_n1051_ & ~new_n1061_;
  assign new_n1063_ = new_n1047_ & ~new_n1062_;
  assign new_n1064_ = ~new_n1046_ & ~new_n1063_;
  assign new_n1065_ = \1_n268  & \1_n685 ;
  assign new_n1066_ = ~\1_n268  & ~\1_n685 ;
  assign new_n1067_ = ~new_n1065_ & ~new_n1066_;
  assign new_n1068_ = ~\1_n688  & new_n1067_;
  assign new_n1069_ = ~\1_n944  & ~new_n1068_;
  assign new_n1070_ = new_n1052_ & new_n1057_;
  assign new_n1071_ = new_n1069_ & new_n1070_;
  assign new_n1072_ = new_n1047_ & new_n1071_;
  assign new_n1073_ = new_n1064_ & ~new_n1072_;
  assign new_n1074_ = new_n1043_ & ~new_n1073_;
  assign new_n1075_ = ~new_n1042_ & ~new_n1074_;
  assign new_n1076_ = ~new_n1039_ & ~new_n1075_;
  assign new_n1077_ = new_n1034_ & ~new_n1076_;
  assign new_n1078_ = new_n1017_ & ~new_n1077_;
  assign new_n1079_ = ~new_n1016_ & ~new_n1078_;
  assign new_n1080_ = \1_n1311  & new_n996_;
  assign new_n1081_ = ~new_n997_ & ~new_n1080_;
  assign new_n1082_ = new_n1002_ & new_n1081_;
  assign new_n1083_ = new_n1006_ & new_n1082_;
  assign new_n1084_ = ~new_n1079_ & new_n1083_;
  assign new_n1085_ = new_n1010_ & new_n1084_;
  assign new_n1086_ = new_n1012_ & ~new_n1085_;
  assign new_n1087_ = new_n988_ & ~new_n1086_;
  assign new_n1088_ = ~new_n987_ & ~new_n1087_;
  assign new_n1089_ = ~new_n983_ & ~new_n1088_;
  assign new_n1090_ = new_n978_ & ~new_n1089_;
  assign new_n1091_ = new_n960_ & ~new_n1090_;
  assign new_n1092_ = ~new_n958_ & ~new_n1091_;
  assign new_n1093_ = new_n951_ & new_n1092_;
  assign new_n1094_ = ~new_n955_ & ~new_n1093_;
  assign new_n1095_ = ~new_n943_ & ~new_n1094_;
  assign new_n1096_ = new_n943_ & new_n1094_;
  assign \1_n81  = ~new_n1095_ & ~new_n1096_;
  assign new_n1098_ = new_n980_ & ~new_n1088_;
  assign new_n1099_ = ~new_n980_ & new_n1088_;
  assign \1_n90  = ~new_n1098_ & ~new_n1099_;
  assign \1_n112  = \1_n116  & \1_n1257 ;
  assign new_n1102_ = ~new_n650_ & ~new_n939_;
  assign new_n1103_ = \1_n332  & new_n1102_;
  assign new_n1104_ = ~\1_n332  & ~new_n1102_;
  assign new_n1105_ = ~new_n1103_ & ~new_n1104_;
  assign new_n1106_ = new_n943_ & ~new_n951_;
  assign new_n1107_ = ~new_n942_ & ~new_n1106_;
  assign new_n1108_ = new_n953_ & ~new_n1092_;
  assign new_n1109_ = new_n943_ & new_n947_;
  assign new_n1110_ = new_n1108_ & new_n1109_;
  assign new_n1111_ = new_n1107_ & ~new_n1110_;
  assign new_n1112_ = ~new_n1105_ & new_n1111_;
  assign new_n1113_ = new_n1105_ & ~new_n1111_;
  assign \1_n129  = ~new_n1112_ & ~new_n1113_;
  assign new_n1115_ = new_n1079_ & ~new_n1081_;
  assign new_n1116_ = ~new_n1079_ & new_n1081_;
  assign \1_n135  = ~new_n1115_ & ~new_n1116_;
  assign new_n1118_ = ~new_n614_ & new_n939_;
  assign new_n1119_ = ~new_n624_ & ~new_n1118_;
  assign new_n1120_ = \1_n599  & ~new_n614_;
  assign new_n1121_ = ~new_n624_ & ~new_n1120_;
  assign new_n1122_ = new_n1119_ & new_n1121_;
  assign new_n1123_ = ~\1_n231  & ~new_n1119_;
  assign new_n1124_ = new_n1105_ & ~new_n1107_;
  assign new_n1125_ = ~new_n1104_ & ~new_n1124_;
  assign new_n1126_ = new_n1105_ & new_n1110_;
  assign new_n1127_ = new_n1125_ & ~new_n1126_;
  assign new_n1128_ = \1_n231  & ~new_n1119_;
  assign new_n1129_ = ~\1_n231  & new_n1119_;
  assign new_n1130_ = ~new_n1128_ & ~new_n1129_;
  assign new_n1131_ = ~new_n1127_ & ~new_n1130_;
  assign new_n1132_ = ~new_n1123_ & ~new_n1131_;
  assign new_n1133_ = \1_n393  & ~new_n1119_;
  assign new_n1134_ = ~\1_n393  & new_n1119_;
  assign new_n1135_ = ~new_n1133_ & ~new_n1134_;
  assign new_n1136_ = ~new_n1132_ & ~new_n1135_;
  assign new_n1137_ = new_n1122_ & ~new_n1136_;
  assign new_n1138_ = new_n1119_ & ~new_n1136_;
  assign new_n1139_ = ~new_n1121_ & ~new_n1138_;
  assign \1_n150  = new_n1137_ | new_n1139_;
  assign new_n1141_ = ~new_n949_ & ~new_n1108_;
  assign new_n1142_ = ~new_n947_ & new_n1141_;
  assign new_n1143_ = new_n947_ & ~new_n1141_;
  assign \1_n167  = ~new_n1142_ & ~new_n1143_;
  assign new_n1145_ = \1_n802  & \1_n1344 ;
  assign new_n1146_ = \1_n288  & \1_n359 ;
  assign \1_n168  = new_n1145_ & new_n1146_;
  assign new_n1148_ = new_n1122_ & ~new_n1134_;
  assign new_n1149_ = \1_n1298  & ~new_n614_;
  assign new_n1150_ = ~new_n624_ & ~new_n1149_;
  assign new_n1151_ = ~new_n1121_ & new_n1150_;
  assign new_n1152_ = new_n1121_ & ~new_n1150_;
  assign new_n1153_ = ~new_n1151_ & ~new_n1152_;
  assign new_n1154_ = \1_n393  & ~new_n1153_;
  assign new_n1155_ = ~\1_n393  & new_n1153_;
  assign new_n1156_ = ~new_n1154_ & ~new_n1155_;
  assign new_n1157_ = ~new_n1148_ & new_n1156_;
  assign new_n1158_ = ~new_n1132_ & new_n1157_;
  assign new_n1159_ = new_n1122_ & ~new_n1156_;
  assign new_n1160_ = new_n1135_ & new_n1159_;
  assign new_n1161_ = ~new_n1132_ & new_n1160_;
  assign new_n1162_ = new_n1122_ & new_n1134_;
  assign new_n1163_ = ~new_n1122_ & ~new_n1134_;
  assign new_n1164_ = ~new_n1162_ & ~new_n1163_;
  assign new_n1165_ = ~new_n1153_ & ~new_n1164_;
  assign new_n1166_ = new_n1153_ & new_n1164_;
  assign new_n1167_ = ~new_n1165_ & ~new_n1166_;
  assign new_n1168_ = ~new_n1119_ & new_n1167_;
  assign new_n1169_ = new_n1119_ & ~new_n1167_;
  assign new_n1170_ = ~new_n1168_ & ~new_n1169_;
  assign new_n1171_ = new_n1132_ & ~new_n1170_;
  assign new_n1172_ = ~new_n1161_ & ~new_n1171_;
  assign new_n1173_ = ~new_n1158_ & new_n1172_;
  assign new_n1174_ = new_n1107_ & ~new_n1109_;
  assign new_n1175_ = new_n953_ & new_n1174_;
  assign new_n1176_ = new_n949_ & new_n1107_;
  assign new_n1177_ = ~new_n949_ & ~new_n1107_;
  assign new_n1178_ = ~new_n1176_ & ~new_n1177_;
  assign new_n1179_ = ~new_n953_ & ~new_n1178_;
  assign new_n1180_ = ~new_n1175_ & ~new_n1179_;
  assign new_n1181_ = ~new_n943_ & new_n955_;
  assign new_n1182_ = new_n943_ & ~new_n955_;
  assign new_n1183_ = ~new_n1181_ & ~new_n1182_;
  assign new_n1184_ = new_n1130_ & ~new_n1183_;
  assign new_n1185_ = ~new_n1130_ & new_n1183_;
  assign new_n1186_ = ~new_n1184_ & ~new_n1185_;
  assign new_n1187_ = ~new_n1180_ & new_n1186_;
  assign new_n1188_ = new_n1180_ & ~new_n1186_;
  assign new_n1189_ = ~new_n1187_ & ~new_n1188_;
  assign new_n1190_ = ~new_n953_ & ~new_n1125_;
  assign new_n1191_ = new_n1105_ & new_n1109_;
  assign new_n1192_ = new_n1125_ & ~new_n1191_;
  assign new_n1193_ = new_n953_ & new_n1192_;
  assign new_n1194_ = ~new_n1190_ & ~new_n1193_;
  assign new_n1195_ = ~new_n1105_ & new_n1194_;
  assign new_n1196_ = new_n1105_ & ~new_n1194_;
  assign new_n1197_ = ~new_n1195_ & ~new_n1196_;
  assign new_n1198_ = ~new_n947_ & new_n1197_;
  assign new_n1199_ = new_n947_ & ~new_n1197_;
  assign new_n1200_ = ~new_n1198_ & ~new_n1199_;
  assign new_n1201_ = ~new_n1189_ & new_n1200_;
  assign new_n1202_ = new_n1189_ & ~new_n1200_;
  assign new_n1203_ = ~new_n1201_ & ~new_n1202_;
  assign new_n1204_ = ~new_n1092_ & ~new_n1203_;
  assign new_n1205_ = new_n1105_ & new_n1130_;
  assign new_n1206_ = ~new_n1105_ & ~new_n1130_;
  assign new_n1207_ = ~new_n1205_ & ~new_n1206_;
  assign new_n1208_ = new_n951_ & ~new_n1207_;
  assign new_n1209_ = ~new_n951_ & new_n1207_;
  assign new_n1210_ = ~new_n1208_ & ~new_n1209_;
  assign new_n1211_ = new_n1178_ & new_n1210_;
  assign new_n1212_ = ~new_n1178_ & ~new_n1210_;
  assign new_n1213_ = ~new_n1211_ & ~new_n1212_;
  assign new_n1214_ = ~new_n947_ & new_n1125_;
  assign new_n1215_ = new_n947_ & ~new_n1125_;
  assign new_n1216_ = ~new_n1214_ & ~new_n1215_;
  assign new_n1217_ = new_n953_ & new_n1216_;
  assign new_n1218_ = ~new_n953_ & ~new_n1216_;
  assign new_n1219_ = ~new_n1217_ & ~new_n1218_;
  assign new_n1220_ = ~new_n943_ & ~new_n1219_;
  assign new_n1221_ = new_n943_ & new_n1219_;
  assign new_n1222_ = ~new_n1220_ & ~new_n1221_;
  assign new_n1223_ = ~new_n1213_ & new_n1222_;
  assign new_n1224_ = new_n1213_ & ~new_n1222_;
  assign new_n1225_ = ~new_n1223_ & ~new_n1224_;
  assign new_n1226_ = new_n1092_ & ~new_n1225_;
  assign new_n1227_ = ~new_n1204_ & ~new_n1226_;
  assign new_n1228_ = ~new_n1173_ & ~new_n1227_;
  assign new_n1229_ = new_n1173_ & new_n1227_;
  assign \1_n190  = ~new_n1228_ & ~new_n1229_;
  assign new_n1231_ = \1_n393  & new_n1132_;
  assign new_n1232_ = ~new_n1119_ & ~new_n1231_;
  assign \1_n204  = new_n1138_ | new_n1232_;
  assign new_n1234_ = new_n1137_ & new_n1150_;
  assign new_n1235_ = \1_n398  & ~new_n614_;
  assign new_n1236_ = ~new_n624_ & ~new_n1235_;
  assign new_n1237_ = \1_n505  & ~new_n614_;
  assign new_n1238_ = ~new_n624_ & ~new_n1237_;
  assign new_n1239_ = new_n1236_ & new_n1238_;
  assign new_n1240_ = \1_n986  & ~new_n614_;
  assign new_n1241_ = ~new_n624_ & ~new_n1240_;
  assign new_n1242_ = new_n1239_ & new_n1241_;
  assign new_n1243_ = new_n1234_ & new_n1242_;
  assign new_n1244_ = \1_n896  & ~new_n614_;
  assign new_n1245_ = ~new_n624_ & ~new_n1244_;
  assign new_n1246_ = new_n1243_ & new_n1245_;
  assign new_n1247_ = \1_n749  & ~new_n614_;
  assign new_n1248_ = ~new_n624_ & ~new_n1247_;
  assign new_n1249_ = ~new_n1246_ & ~new_n1248_;
  assign new_n1250_ = new_n1246_ & new_n1248_;
  assign \1_n206  = new_n1249_ | new_n1250_;
  assign new_n1252_ = new_n1234_ & new_n1239_;
  assign new_n1253_ = new_n1234_ & new_n1238_;
  assign new_n1254_ = ~new_n1236_ & ~new_n1253_;
  assign \1_n218  = new_n1252_ | new_n1254_;
  assign new_n1256_ = \1_n944  & new_n1068_;
  assign \1_n228  = ~new_n1069_ & ~new_n1256_;
  assign \1_n679  = \1_n1352  | ~new_n1250_;
  assign \1_n299  = \1_n679 ;
  assign new_n1260_ = ~new_n1250_ & \1_n299 ;
  assign \1_n229  = ~\1_n679  | new_n1260_;
  assign new_n1262_ = new_n1058_ & ~new_n1062_;
  assign new_n1263_ = ~new_n1058_ & new_n1062_;
  assign new_n1264_ = ~new_n1262_ & ~new_n1263_;
  assign new_n1265_ = ~new_n1047_ & new_n1060_;
  assign new_n1266_ = new_n1047_ & ~new_n1060_;
  assign new_n1267_ = ~new_n1265_ & ~new_n1266_;
  assign new_n1268_ = new_n1043_ & ~new_n1267_;
  assign new_n1269_ = ~new_n1043_ & new_n1267_;
  assign new_n1270_ = ~new_n1268_ & ~new_n1269_;
  assign new_n1271_ = ~new_n1264_ & new_n1270_;
  assign new_n1272_ = new_n1264_ & ~new_n1270_;
  assign new_n1273_ = ~new_n1271_ & ~new_n1272_;
  assign new_n1274_ = ~new_n1057_ & new_n1068_;
  assign new_n1275_ = new_n1057_ & ~new_n1068_;
  assign new_n1276_ = ~new_n1274_ & ~new_n1275_;
  assign new_n1277_ = ~new_n1052_ & new_n1276_;
  assign new_n1278_ = new_n1052_ & ~new_n1276_;
  assign new_n1279_ = ~new_n1277_ & ~new_n1278_;
  assign new_n1280_ = ~new_n1064_ & new_n1279_;
  assign new_n1281_ = new_n1064_ & ~new_n1279_;
  assign new_n1282_ = ~new_n1280_ & ~new_n1281_;
  assign new_n1283_ = ~new_n1273_ & new_n1282_;
  assign new_n1284_ = new_n1273_ & ~new_n1282_;
  assign new_n1285_ = ~new_n1283_ & ~new_n1284_;
  assign new_n1286_ = \1_n944  & new_n1285_;
  assign new_n1287_ = new_n1060_ & ~new_n1275_;
  assign new_n1288_ = new_n1043_ & new_n1287_;
  assign new_n1289_ = ~new_n1043_ & ~new_n1287_;
  assign new_n1290_ = ~new_n1288_ & ~new_n1289_;
  assign new_n1291_ = ~new_n1052_ & new_n1290_;
  assign new_n1292_ = new_n1052_ & ~new_n1290_;
  assign new_n1293_ = ~new_n1291_ & ~new_n1292_;
  assign new_n1294_ = new_n1062_ & ~new_n1070_;
  assign new_n1295_ = ~new_n1068_ & new_n1294_;
  assign new_n1296_ = new_n1068_ & new_n1264_;
  assign new_n1297_ = ~new_n1295_ & ~new_n1296_;
  assign new_n1298_ = ~new_n1064_ & new_n1068_;
  assign new_n1299_ = new_n1047_ & new_n1070_;
  assign new_n1300_ = new_n1064_ & ~new_n1299_;
  assign new_n1301_ = ~new_n1068_ & new_n1300_;
  assign new_n1302_ = ~new_n1298_ & ~new_n1301_;
  assign new_n1303_ = ~new_n1047_ & new_n1302_;
  assign new_n1304_ = new_n1047_ & ~new_n1302_;
  assign new_n1305_ = ~new_n1303_ & ~new_n1304_;
  assign new_n1306_ = ~new_n1057_ & new_n1305_;
  assign new_n1307_ = new_n1057_ & ~new_n1305_;
  assign new_n1308_ = ~new_n1306_ & ~new_n1307_;
  assign new_n1309_ = ~new_n1297_ & new_n1308_;
  assign new_n1310_ = new_n1297_ & ~new_n1308_;
  assign new_n1311_ = ~new_n1309_ & ~new_n1310_;
  assign new_n1312_ = ~new_n1293_ & new_n1311_;
  assign new_n1313_ = new_n1293_ & ~new_n1311_;
  assign new_n1314_ = ~new_n1312_ & ~new_n1313_;
  assign new_n1315_ = ~\1_n944  & ~new_n1314_;
  assign new_n1316_ = ~new_n1286_ & ~new_n1315_;
  assign new_n1317_ = ~new_n1027_ & ~new_n1036_;
  assign new_n1318_ = ~new_n1037_ & ~new_n1317_;
  assign new_n1319_ = ~new_n1034_ & ~new_n1318_;
  assign new_n1320_ = new_n1034_ & new_n1318_;
  assign new_n1321_ = ~new_n1319_ & ~new_n1320_;
  assign new_n1322_ = new_n1030_ & new_n1321_;
  assign new_n1323_ = ~new_n1030_ & ~new_n1321_;
  assign new_n1324_ = ~new_n1322_ & ~new_n1323_;
  assign new_n1325_ = new_n1032_ & new_n1324_;
  assign new_n1326_ = ~new_n1032_ & ~new_n1324_;
  assign new_n1327_ = ~new_n1325_ & ~new_n1326_;
  assign new_n1328_ = new_n1075_ & new_n1327_;
  assign new_n1329_ = new_n1032_ & ~new_n1037_;
  assign new_n1330_ = ~new_n1030_ & ~new_n1036_;
  assign new_n1331_ = new_n1039_ & new_n1318_;
  assign new_n1332_ = ~new_n1039_ & ~new_n1318_;
  assign new_n1333_ = ~new_n1331_ & ~new_n1332_;
  assign new_n1334_ = ~new_n1330_ & new_n1333_;
  assign new_n1335_ = new_n1330_ & ~new_n1333_;
  assign new_n1336_ = ~new_n1334_ & ~new_n1335_;
  assign new_n1337_ = new_n1329_ & new_n1336_;
  assign new_n1338_ = ~new_n1329_ & ~new_n1336_;
  assign new_n1339_ = ~new_n1337_ & ~new_n1338_;
  assign new_n1340_ = ~new_n1075_ & ~new_n1339_;
  assign new_n1341_ = ~new_n1328_ & ~new_n1340_;
  assign new_n1342_ = ~new_n1022_ & ~new_n1341_;
  assign new_n1343_ = new_n1022_ & new_n1341_;
  assign new_n1344_ = ~new_n1342_ & ~new_n1343_;
  assign new_n1345_ = ~new_n1017_ & new_n1344_;
  assign new_n1346_ = new_n1017_ & ~new_n1344_;
  assign new_n1347_ = ~new_n1345_ & ~new_n1346_;
  assign new_n1348_ = ~new_n1316_ & new_n1347_;
  assign new_n1349_ = new_n1316_ & ~new_n1347_;
  assign \1_n240  = ~new_n1348_ & ~new_n1349_;
  assign new_n1351_ = ~new_n1241_ & ~new_n1252_;
  assign \1_n389  = new_n1243_ | new_n1351_;
  assign new_n1353_ = ~new_n870_ & new_n901_;
  assign new_n1354_ = new_n870_ & ~new_n901_;
  assign new_n1355_ = ~new_n1353_ & ~new_n1354_;
  assign new_n1356_ = ~new_n890_ & ~new_n1355_;
  assign new_n1357_ = new_n890_ & new_n1355_;
  assign new_n1358_ = ~new_n1356_ & ~new_n1357_;
  assign new_n1359_ = ~new_n881_ & new_n1358_;
  assign new_n1360_ = new_n881_ & ~new_n1358_;
  assign new_n1361_ = ~new_n1359_ & ~new_n1360_;
  assign new_n1362_ = ~\1_n268  & \1_n688 ;
  assign new_n1363_ = ~\1_n688  & \1_n857 ;
  assign new_n1364_ = ~new_n1362_ & ~new_n1363_;
  assign new_n1365_ = ~\1_n381  & \1_n688 ;
  assign new_n1366_ = ~\1_n688  & \1_n1269 ;
  assign new_n1367_ = ~new_n1365_ & ~new_n1366_;
  assign new_n1368_ = ~new_n1364_ & ~new_n1367_;
  assign new_n1369_ = new_n1364_ & new_n1367_;
  assign new_n1370_ = ~new_n1368_ & ~new_n1369_;
  assign new_n1371_ = new_n849_ & ~new_n859_;
  assign new_n1372_ = ~new_n849_ & new_n859_;
  assign new_n1373_ = ~new_n1371_ & ~new_n1372_;
  assign new_n1374_ = ~new_n1370_ & new_n1373_;
  assign new_n1375_ = new_n1370_ & ~new_n1373_;
  assign new_n1376_ = ~new_n1374_ & ~new_n1375_;
  assign new_n1377_ = ~new_n830_ & new_n1376_;
  assign new_n1378_ = new_n830_ & ~new_n1376_;
  assign new_n1379_ = ~new_n1377_ & ~new_n1378_;
  assign new_n1380_ = ~new_n837_ & new_n1379_;
  assign new_n1381_ = new_n837_ & ~new_n1379_;
  assign new_n1382_ = ~new_n1380_ & ~new_n1381_;
  assign new_n1383_ = ~new_n1361_ & new_n1382_;
  assign new_n1384_ = new_n1361_ & ~new_n1382_;
  assign new_n1385_ = ~new_n1383_ & ~new_n1384_;
  assign new_n1386_ = ~new_n762_ & new_n782_;
  assign new_n1387_ = new_n762_ & ~new_n782_;
  assign new_n1388_ = ~new_n1386_ & ~new_n1387_;
  assign new_n1389_ = new_n793_ & new_n1388_;
  assign new_n1390_ = ~new_n793_ & ~new_n1388_;
  assign new_n1391_ = ~new_n1389_ & ~new_n1390_;
  assign new_n1392_ = ~new_n773_ & new_n1391_;
  assign new_n1393_ = new_n773_ & ~new_n1391_;
  assign new_n1394_ = ~new_n1392_ & ~new_n1393_;
  assign new_n1395_ = \1_n688  & ~\1_n1342 ;
  assign new_n1396_ = \1_n267  & ~\1_n688 ;
  assign new_n1397_ = ~new_n1395_ & ~new_n1396_;
  assign new_n1398_ = ~new_n722_ & ~new_n1397_;
  assign new_n1399_ = new_n722_ & new_n1397_;
  assign new_n1400_ = ~new_n1398_ & ~new_n1399_;
  assign new_n1401_ = ~new_n756_ & new_n1400_;
  assign new_n1402_ = new_n756_ & ~new_n1400_;
  assign new_n1403_ = ~new_n1401_ & ~new_n1402_;
  assign new_n1404_ = ~new_n728_ & new_n1403_;
  assign new_n1405_ = new_n728_ & ~new_n1403_;
  assign new_n1406_ = ~new_n1404_ & ~new_n1405_;
  assign new_n1407_ = ~new_n737_ & new_n1406_;
  assign new_n1408_ = new_n737_ & ~new_n1406_;
  assign new_n1409_ = ~new_n1407_ & ~new_n1408_;
  assign new_n1410_ = ~new_n746_ & new_n1409_;
  assign new_n1411_ = new_n746_ & ~new_n1409_;
  assign new_n1412_ = ~new_n1410_ & ~new_n1411_;
  assign new_n1413_ = ~new_n1394_ & new_n1412_;
  assign new_n1414_ = new_n1394_ & ~new_n1412_;
  assign new_n1415_ = ~new_n1413_ & ~new_n1414_;
  assign new_n1416_ = ~new_n626_ & new_n640_;
  assign new_n1417_ = new_n626_ & ~new_n640_;
  assign new_n1418_ = ~new_n1416_ & ~new_n1417_;
  assign new_n1419_ = new_n636_ & new_n1418_;
  assign new_n1420_ = ~new_n636_ & ~new_n1418_;
  assign new_n1421_ = ~new_n1419_ & ~new_n1420_;
  assign new_n1422_ = new_n655_ & new_n661_;
  assign new_n1423_ = ~new_n655_ & ~new_n661_;
  assign new_n1424_ = ~new_n1422_ & ~new_n1423_;
  assign new_n1425_ = \1_n688  & ~\1_n819 ;
  assign new_n1426_ = ~\1_n688  & \1_n818 ;
  assign new_n1427_ = ~new_n1425_ & ~new_n1426_;
  assign new_n1428_ = ~new_n690_ & ~new_n1427_;
  assign new_n1429_ = new_n690_ & new_n1427_;
  assign new_n1430_ = ~new_n1428_ & ~new_n1429_;
  assign new_n1431_ = ~new_n648_ & new_n1430_;
  assign new_n1432_ = new_n648_ & ~new_n1430_;
  assign new_n1433_ = ~new_n1431_ & ~new_n1432_;
  assign new_n1434_ = ~new_n673_ & new_n1433_;
  assign new_n1435_ = new_n673_ & ~new_n1433_;
  assign new_n1436_ = ~new_n1434_ & ~new_n1435_;
  assign new_n1437_ = new_n1424_ & new_n1436_;
  assign new_n1438_ = ~new_n1424_ & ~new_n1436_;
  assign new_n1439_ = ~new_n1437_ & ~new_n1438_;
  assign new_n1440_ = ~new_n628_ & new_n1439_;
  assign new_n1441_ = new_n628_ & ~new_n1439_;
  assign new_n1442_ = ~new_n1440_ & ~new_n1441_;
  assign new_n1443_ = ~new_n1421_ & new_n1442_;
  assign new_n1444_ = new_n1421_ & ~new_n1442_;
  assign new_n1445_ = ~new_n1443_ & ~new_n1444_;
  assign new_n1446_ = ~new_n1415_ & ~new_n1445_;
  assign new_n1447_ = ~new_n1385_ & new_n1446_;
  assign new_n1448_ = \1_n839  & ~\1_n1022 ;
  assign new_n1449_ = ~\1_n839  & \1_n1022 ;
  assign new_n1450_ = ~new_n1448_ & ~new_n1449_;
  assign new_n1451_ = ~\1_n688  & ~new_n1450_;
  assign new_n1452_ = ~\1_n475  & \1_n688 ;
  assign new_n1453_ = ~\1_n688  & \1_n1231 ;
  assign new_n1454_ = ~new_n1452_ & ~new_n1453_;
  assign new_n1455_ = ~new_n611_ & new_n1454_;
  assign new_n1456_ = new_n611_ & ~new_n1454_;
  assign new_n1457_ = ~new_n1455_ & ~new_n1456_;
  assign new_n1458_ = ~new_n1451_ & new_n1457_;
  assign new_n1459_ = new_n1451_ & ~new_n1457_;
  assign new_n1460_ = ~new_n1458_ & ~new_n1459_;
  assign \1_n408  = new_n1447_ & new_n1460_;
  assign new_n1462_ = ~new_n1245_ & new_n1248_;
  assign new_n1463_ = new_n1245_ & ~new_n1248_;
  assign new_n1464_ = ~new_n1462_ & ~new_n1463_;
  assign new_n1465_ = ~new_n1236_ & ~new_n1241_;
  assign new_n1466_ = new_n1236_ & new_n1241_;
  assign new_n1467_ = ~new_n1465_ & ~new_n1466_;
  assign new_n1468_ = new_n1238_ & ~new_n1467_;
  assign new_n1469_ = ~new_n1238_ & new_n1467_;
  assign new_n1470_ = ~new_n1468_ & ~new_n1469_;
  assign new_n1471_ = new_n1238_ & ~new_n1239_;
  assign new_n1472_ = ~new_n1242_ & ~new_n1471_;
  assign new_n1473_ = new_n1234_ & new_n1472_;
  assign new_n1474_ = new_n1470_ & ~new_n1473_;
  assign new_n1475_ = ~new_n1470_ & new_n1473_;
  assign new_n1476_ = ~new_n1474_ & ~new_n1475_;
  assign new_n1477_ = ~new_n1246_ & new_n1476_;
  assign new_n1478_ = ~new_n1464_ & new_n1477_;
  assign new_n1479_ = new_n1464_ & ~new_n1477_;
  assign new_n1480_ = ~new_n1478_ & ~new_n1479_;
  assign new_n1481_ = \1_n1352  & new_n1250_;
  assign \1_n409  = ~new_n1480_ & ~new_n1481_;
  assign \1_n432  = \1_n127  | \1_n976 ;
  assign \1_n592  = \1_n432 ;
  assign new_n1485_ = \1_n491  & \1_n787 ;
  assign \1_n598  = \1_n432 ;
  assign new_n1487_ = new_n981_ & ~new_n1088_;
  assign new_n1488_ = new_n976_ & ~new_n1487_;
  assign new_n1489_ = ~new_n966_ & new_n1488_;
  assign new_n1490_ = new_n966_ & ~new_n1488_;
  assign \1_n607  = ~new_n1489_ & ~new_n1490_;
  assign new_n1492_ = new_n1062_ & ~new_n1071_;
  assign new_n1493_ = ~new_n1047_ & new_n1492_;
  assign new_n1494_ = new_n1047_ & ~new_n1492_;
  assign \1_n621  = ~new_n1493_ & ~new_n1494_;
  assign new_n1496_ = ~new_n953_ & new_n1092_;
  assign \1_n627  = ~new_n1108_ & ~new_n1496_;
  assign new_n1498_ = ~new_n968_ & new_n973_;
  assign new_n1499_ = new_n968_ & ~new_n973_;
  assign new_n1500_ = ~new_n1498_ & ~new_n1499_;
  assign new_n1501_ = new_n957_ & new_n1500_;
  assign new_n1502_ = ~new_n957_ & ~new_n1500_;
  assign new_n1503_ = ~new_n1501_ & ~new_n1502_;
  assign new_n1504_ = ~new_n963_ & new_n1503_;
  assign new_n1505_ = new_n963_ & ~new_n1503_;
  assign new_n1506_ = ~new_n1504_ & ~new_n1505_;
  assign new_n1507_ = \1_n688  & \1_n767 ;
  assign new_n1508_ = \1_n192  & ~\1_n688 ;
  assign new_n1509_ = ~new_n1507_ & ~new_n1508_;
  assign new_n1510_ = new_n996_ & ~new_n1509_;
  assign new_n1511_ = ~new_n996_ & new_n1509_;
  assign new_n1512_ = ~new_n1510_ & ~new_n1511_;
  assign new_n1513_ = ~new_n993_ & new_n999_;
  assign new_n1514_ = new_n993_ & ~new_n999_;
  assign new_n1515_ = ~new_n1513_ & ~new_n1514_;
  assign new_n1516_ = ~new_n1512_ & new_n1515_;
  assign new_n1517_ = new_n1512_ & ~new_n1515_;
  assign new_n1518_ = ~new_n1516_ & ~new_n1517_;
  assign new_n1519_ = new_n985_ & new_n1518_;
  assign new_n1520_ = ~new_n985_ & ~new_n1518_;
  assign new_n1521_ = ~new_n1519_ & ~new_n1520_;
  assign new_n1522_ = new_n990_ & new_n1521_;
  assign new_n1523_ = ~new_n990_ & ~new_n1521_;
  assign new_n1524_ = ~new_n1522_ & ~new_n1523_;
  assign new_n1525_ = ~new_n1506_ & new_n1524_;
  assign new_n1526_ = new_n1506_ & ~new_n1524_;
  assign new_n1527_ = ~new_n1525_ & ~new_n1526_;
  assign new_n1528_ = \1_n688  & \1_n1163 ;
  assign new_n1529_ = ~\1_n688  & \1_n1143 ;
  assign new_n1530_ = ~new_n1528_ & ~new_n1529_;
  assign new_n1531_ = new_n948_ & ~new_n1530_;
  assign new_n1532_ = ~new_n948_ & new_n1530_;
  assign new_n1533_ = ~new_n1531_ & ~new_n1532_;
  assign new_n1534_ = new_n1102_ & new_n1533_;
  assign new_n1535_ = ~new_n1102_ & ~new_n1533_;
  assign new_n1536_ = ~new_n1534_ & ~new_n1535_;
  assign new_n1537_ = ~new_n1119_ & new_n1536_;
  assign new_n1538_ = new_n1119_ & ~new_n1536_;
  assign new_n1539_ = ~new_n1537_ & ~new_n1538_;
  assign new_n1540_ = ~new_n1153_ & ~new_n1539_;
  assign new_n1541_ = new_n1153_ & new_n1539_;
  assign new_n1542_ = ~new_n1540_ & ~new_n1541_;
  assign new_n1543_ = new_n944_ & new_n1542_;
  assign new_n1544_ = ~new_n944_ & ~new_n1542_;
  assign new_n1545_ = ~new_n1543_ & ~new_n1544_;
  assign new_n1546_ = new_n940_ & new_n1545_;
  assign new_n1547_ = ~new_n940_ & ~new_n1545_;
  assign new_n1548_ = ~new_n1546_ & ~new_n1547_;
  assign new_n1549_ = \1_n507  & ~new_n614_;
  assign new_n1550_ = ~new_n624_ & ~new_n1549_;
  assign new_n1551_ = ~new_n614_ & ~new_n624_;
  assign new_n1552_ = ~\1_n439  & new_n1551_;
  assign new_n1553_ = ~new_n1470_ & ~new_n1552_;
  assign new_n1554_ = new_n1470_ & new_n1552_;
  assign new_n1555_ = ~new_n1553_ & ~new_n1554_;
  assign new_n1556_ = ~new_n1464_ & ~new_n1555_;
  assign new_n1557_ = new_n1464_ & new_n1555_;
  assign new_n1558_ = ~new_n1556_ & ~new_n1557_;
  assign new_n1559_ = new_n1550_ & new_n1558_;
  assign new_n1560_ = ~new_n1550_ & ~new_n1558_;
  assign new_n1561_ = ~new_n1559_ & ~new_n1560_;
  assign new_n1562_ = ~new_n1548_ & ~new_n1561_;
  assign new_n1563_ = ~new_n1527_ & new_n1562_;
  assign new_n1564_ = ~new_n1024_ & new_n1029_;
  assign new_n1565_ = new_n1024_ & ~new_n1029_;
  assign new_n1566_ = ~new_n1564_ & ~new_n1565_;
  assign new_n1567_ = new_n1019_ & new_n1566_;
  assign new_n1568_ = ~new_n1019_ & ~new_n1566_;
  assign new_n1569_ = ~new_n1567_ & ~new_n1568_;
  assign new_n1570_ = new_n1014_ & new_n1569_;
  assign new_n1571_ = ~new_n1014_ & ~new_n1569_;
  assign new_n1572_ = ~new_n1570_ & ~new_n1571_;
  assign new_n1573_ = ~new_n1049_ & new_n1054_;
  assign new_n1574_ = new_n1049_ & ~new_n1054_;
  assign new_n1575_ = ~new_n1573_ & ~new_n1574_;
  assign new_n1576_ = \1_n128  & \1_n688 ;
  assign new_n1577_ = \1_n153  & ~\1_n688 ;
  assign new_n1578_ = ~new_n1576_ & ~new_n1577_;
  assign new_n1579_ = \1_n252  & \1_n688 ;
  assign new_n1580_ = ~new_n923_ & ~new_n1579_;
  assign new_n1581_ = new_n1578_ & ~new_n1580_;
  assign new_n1582_ = ~new_n1578_ & new_n1580_;
  assign new_n1583_ = ~new_n1581_ & ~new_n1582_;
  assign new_n1584_ = ~new_n1575_ & new_n1583_;
  assign new_n1585_ = new_n1575_ & ~new_n1583_;
  assign new_n1586_ = ~new_n1584_ & ~new_n1585_;
  assign new_n1587_ = new_n1040_ & new_n1586_;
  assign new_n1588_ = ~new_n1040_ & ~new_n1586_;
  assign new_n1589_ = ~new_n1587_ & ~new_n1588_;
  assign new_n1590_ = new_n1044_ & new_n1589_;
  assign new_n1591_ = ~new_n1044_ & ~new_n1589_;
  assign new_n1592_ = ~new_n1590_ & ~new_n1591_;
  assign new_n1593_ = ~new_n1572_ & new_n1592_;
  assign new_n1594_ = new_n1572_ & ~new_n1592_;
  assign new_n1595_ = ~new_n1593_ & ~new_n1594_;
  assign \1_n653  = new_n1563_ & ~new_n1595_;
  assign new_n1597_ = new_n1037_ & ~new_n1075_;
  assign new_n1598_ = new_n1032_ & ~new_n1597_;
  assign new_n1599_ = ~new_n1022_ & new_n1598_;
  assign new_n1600_ = new_n1022_ & ~new_n1598_;
  assign \1_n662  = ~new_n1599_ & ~new_n1600_;
  assign new_n1602_ = new_n1127_ & new_n1130_;
  assign \1_n707  = ~new_n1131_ & ~new_n1602_;
  assign new_n1604_ = ~new_n1017_ & new_n1077_;
  assign \1_n723  = ~new_n1078_ & ~new_n1604_;
  assign new_n1606_ = new_n1132_ & new_n1135_;
  assign \1_n733  = ~new_n1136_ & ~new_n1606_;
  assign new_n1608_ = ~new_n974_ & ~new_n980_;
  assign new_n1609_ = ~new_n974_ & new_n1088_;
  assign new_n1610_ = ~new_n1608_ & ~new_n1609_;
  assign new_n1611_ = new_n971_ & new_n1610_;
  assign new_n1612_ = ~new_n971_ & ~new_n1610_;
  assign \1_n747  = ~new_n1611_ & ~new_n1612_;
  assign new_n1614_ = ~new_n1137_ & ~new_n1150_;
  assign \1_n779  = new_n1234_ | new_n1614_;
  assign new_n1616_ = new_n1036_ & ~new_n1075_;
  assign new_n1617_ = ~new_n1036_ & new_n1075_;
  assign \1_n808  = ~new_n1616_ & ~new_n1617_;
  assign new_n1619_ = new_n873_ & ~new_n897_;
  assign new_n1620_ = ~new_n873_ & new_n897_;
  assign new_n1621_ = ~new_n1619_ & ~new_n1620_;
  assign new_n1622_ = new_n878_ & new_n1621_;
  assign new_n1623_ = ~new_n878_ & ~new_n1621_;
  assign new_n1624_ = ~new_n1622_ & ~new_n1623_;
  assign new_n1625_ = new_n887_ & new_n1624_;
  assign new_n1626_ = ~new_n887_ & ~new_n1624_;
  assign new_n1627_ = ~new_n1625_ & ~new_n1626_;
  assign new_n1628_ = ~\1_n153  & ~\1_n688 ;
  assign new_n1629_ = ~new_n921_ & new_n1628_;
  assign new_n1630_ = new_n921_ & ~new_n1628_;
  assign new_n1631_ = ~new_n1629_ & ~new_n1630_;
  assign new_n1632_ = ~new_n846_ & new_n856_;
  assign new_n1633_ = new_n846_ & ~new_n856_;
  assign new_n1634_ = ~new_n1632_ & ~new_n1633_;
  assign new_n1635_ = ~new_n1631_ & new_n1634_;
  assign new_n1636_ = new_n1631_ & ~new_n1634_;
  assign new_n1637_ = ~new_n1635_ & ~new_n1636_;
  assign new_n1638_ = new_n827_ & new_n1637_;
  assign new_n1639_ = ~new_n827_ & ~new_n1637_;
  assign new_n1640_ = ~new_n1638_ & ~new_n1639_;
  assign new_n1641_ = new_n834_ & new_n1640_;
  assign new_n1642_ = ~new_n834_ & ~new_n1640_;
  assign new_n1643_ = ~new_n1641_ & ~new_n1642_;
  assign new_n1644_ = ~new_n1627_ & new_n1643_;
  assign new_n1645_ = new_n1627_ & ~new_n1643_;
  assign new_n1646_ = ~new_n1644_ & ~new_n1645_;
  assign new_n1647_ = \1_n851  & ~\1_n955 ;
  assign new_n1648_ = ~\1_n851  & \1_n955 ;
  assign new_n1649_ = ~new_n1647_ & ~new_n1648_;
  assign new_n1650_ = new_n1551_ & ~new_n1649_;
  assign new_n1651_ = ~\1_n49  & \1_n244 ;
  assign new_n1652_ = \1_n49  & ~\1_n244 ;
  assign new_n1653_ = ~new_n1651_ & ~new_n1652_;
  assign new_n1654_ = new_n1551_ & new_n1653_;
  assign new_n1655_ = ~\1_n438  & \1_n1048 ;
  assign new_n1656_ = \1_n438  & ~\1_n1048 ;
  assign new_n1657_ = ~new_n1655_ & ~new_n1656_;
  assign new_n1658_ = new_n1551_ & ~new_n1657_;
  assign new_n1659_ = ~new_n1654_ & new_n1658_;
  assign new_n1660_ = new_n1654_ & ~new_n1658_;
  assign new_n1661_ = ~new_n1659_ & ~new_n1660_;
  assign new_n1662_ = ~new_n1650_ & new_n1661_;
  assign new_n1663_ = new_n1650_ & ~new_n1661_;
  assign new_n1664_ = ~new_n1662_ & ~new_n1663_;
  assign new_n1665_ = ~\1_n433  & \1_n688 ;
  assign new_n1666_ = ~new_n1529_ & ~new_n1665_;
  assign new_n1667_ = new_n695_ & ~new_n1666_;
  assign new_n1668_ = ~new_n695_ & new_n1666_;
  assign new_n1669_ = ~new_n1667_ & ~new_n1668_;
  assign new_n1670_ = ~new_n645_ & new_n670_;
  assign new_n1671_ = new_n645_ & ~new_n670_;
  assign new_n1672_ = ~new_n1670_ & ~new_n1671_;
  assign new_n1673_ = ~new_n1669_ & new_n1672_;
  assign new_n1674_ = new_n1669_ & ~new_n1672_;
  assign new_n1675_ = ~new_n1673_ & ~new_n1674_;
  assign new_n1676_ = ~new_n652_ & new_n663_;
  assign new_n1677_ = new_n652_ & ~new_n663_;
  assign new_n1678_ = ~new_n1676_ & ~new_n1677_;
  assign new_n1679_ = ~new_n1675_ & new_n1678_;
  assign new_n1680_ = new_n1675_ & ~new_n1678_;
  assign new_n1681_ = ~new_n1679_ & ~new_n1680_;
  assign new_n1682_ = ~new_n625_ & new_n639_;
  assign new_n1683_ = new_n625_ & ~new_n639_;
  assign new_n1684_ = ~new_n1682_ & ~new_n1683_;
  assign new_n1685_ = new_n630_ & new_n1684_;
  assign new_n1686_ = ~new_n630_ & ~new_n1684_;
  assign new_n1687_ = ~new_n1685_ & ~new_n1686_;
  assign new_n1688_ = new_n633_ & new_n1687_;
  assign new_n1689_ = ~new_n633_ & ~new_n1687_;
  assign new_n1690_ = ~new_n1688_ & ~new_n1689_;
  assign new_n1691_ = ~new_n1681_ & new_n1690_;
  assign new_n1692_ = new_n1681_ & ~new_n1690_;
  assign new_n1693_ = ~new_n1691_ & ~new_n1692_;
  assign new_n1694_ = ~new_n1664_ & ~new_n1693_;
  assign new_n1695_ = ~new_n1646_ & new_n1694_;
  assign new_n1696_ = new_n765_ & ~new_n789_;
  assign new_n1697_ = ~new_n765_ & new_n789_;
  assign new_n1698_ = ~new_n1696_ & ~new_n1697_;
  assign new_n1699_ = new_n779_ & new_n1698_;
  assign new_n1700_ = ~new_n779_ & ~new_n1698_;
  assign new_n1701_ = ~new_n1699_ & ~new_n1700_;
  assign new_n1702_ = new_n770_ & new_n1701_;
  assign new_n1703_ = ~new_n770_ & ~new_n1701_;
  assign new_n1704_ = ~new_n1702_ & ~new_n1703_;
  assign new_n1705_ = new_n734_ & new_n743_;
  assign new_n1706_ = ~new_n734_ & ~new_n743_;
  assign new_n1707_ = ~new_n1705_ & ~new_n1706_;
  assign new_n1708_ = \1_n688  & ~\1_n1067 ;
  assign new_n1709_ = ~new_n1508_ & ~new_n1708_;
  assign new_n1710_ = ~new_n719_ & ~new_n1709_;
  assign new_n1711_ = new_n719_ & new_n1709_;
  assign new_n1712_ = ~new_n1710_ & ~new_n1711_;
  assign new_n1713_ = new_n753_ & new_n1712_;
  assign new_n1714_ = ~new_n753_ & ~new_n1712_;
  assign new_n1715_ = ~new_n1713_ & ~new_n1714_;
  assign new_n1716_ = new_n725_ & new_n1715_;
  assign new_n1717_ = ~new_n725_ & ~new_n1715_;
  assign new_n1718_ = ~new_n1716_ & ~new_n1717_;
  assign new_n1719_ = new_n1707_ & new_n1718_;
  assign new_n1720_ = ~new_n1707_ & ~new_n1718_;
  assign new_n1721_ = ~new_n1719_ & ~new_n1720_;
  assign new_n1722_ = ~new_n1704_ & new_n1721_;
  assign new_n1723_ = new_n1704_ & ~new_n1721_;
  assign new_n1724_ = ~new_n1722_ & ~new_n1723_;
  assign \1_n817  = new_n1695_ & new_n1724_;
  assign new_n1726_ = new_n1004_ & ~new_n1082_;
  assign new_n1727_ = new_n1004_ & new_n1079_;
  assign new_n1728_ = ~new_n1726_ & ~new_n1727_;
  assign new_n1729_ = ~new_n1006_ & ~new_n1728_;
  assign new_n1730_ = new_n1006_ & new_n1728_;
  assign \1_n835  = ~new_n1729_ & ~new_n1730_;
  assign new_n1732_ = \1_n448  & \1_n870 ;
  assign new_n1733_ = \1_n324  & \1_n577 ;
  assign \1_n854  = new_n1732_ & new_n1733_;
  assign new_n1735_ = ~new_n1234_ & new_n1238_;
  assign new_n1736_ = new_n1234_ & ~new_n1238_;
  assign \1_n905  = ~new_n1735_ & ~new_n1736_;
  assign new_n1738_ = \1_n408  & \1_n817 ;
  assign new_n1739_ = \1_n653  & new_n1738_;
  assign new_n1740_ = \1_n21  & \1_n1226 ;
  assign new_n1741_ = \1_n635  & \1_n766 ;
  assign \1_n999  = new_n1740_ & new_n1741_;
  assign new_n1743_ = new_n1739_ & \1_n999 ;
  assign new_n1744_ = \1_n168  & new_n1743_;
  assign new_n1745_ = \1_n854  & new_n1744_;
  assign new_n1746_ = \1_n319  & \1_n1236 ;
  assign new_n1747_ = \1_n952  & \1_n1029 ;
  assign \1_n1027  = new_n1746_ & new_n1747_;
  assign \1_n927  = new_n1745_ & \1_n1027 ;
  assign new_n1750_ = ~new_n1030_ & new_n1075_;
  assign new_n1751_ = ~new_n1330_ & ~new_n1750_;
  assign new_n1752_ = new_n1027_ & new_n1751_;
  assign new_n1753_ = ~new_n1027_ & ~new_n1751_;
  assign \1_n962  = ~new_n1752_ & ~new_n1753_;
  assign new_n1755_ = new_n1008_ & ~new_n1084_;
  assign new_n1756_ = new_n1010_ & ~new_n1755_;
  assign new_n1757_ = ~new_n1010_ & new_n1755_;
  assign \1_n1059  = ~new_n1756_ & ~new_n1757_;
  assign new_n1759_ = ~new_n988_ & new_n1086_;
  assign \1_n1061  = ~new_n1087_ & ~new_n1759_;
  assign new_n1761_ = ~new_n1043_ & new_n1073_;
  assign \1_n1085  = ~new_n1074_ & ~new_n1761_;
  assign new_n1763_ = ~new_n1243_ & ~new_n1245_;
  assign \1_n1099  = new_n1246_ | new_n1763_;
  assign new_n1765_ = new_n1004_ & new_n1010_;
  assign new_n1766_ = ~new_n1004_ & ~new_n1010_;
  assign new_n1767_ = ~new_n1765_ & ~new_n1766_;
  assign new_n1768_ = new_n988_ & ~new_n1767_;
  assign new_n1769_ = ~new_n988_ & new_n1767_;
  assign new_n1770_ = ~new_n1768_ & ~new_n1769_;
  assign new_n1771_ = ~new_n997_ & new_n1770_;
  assign new_n1772_ = new_n997_ & ~new_n1770_;
  assign new_n1773_ = ~new_n1771_ & ~new_n1772_;
  assign new_n1774_ = new_n1008_ & new_n1773_;
  assign new_n1775_ = ~new_n1008_ & ~new_n1773_;
  assign new_n1776_ = ~new_n1774_ & ~new_n1775_;
  assign new_n1777_ = ~new_n1012_ & ~new_n1081_;
  assign new_n1778_ = new_n1012_ & new_n1081_;
  assign new_n1779_ = ~new_n1777_ & ~new_n1778_;
  assign new_n1780_ = ~new_n1006_ & new_n1779_;
  assign new_n1781_ = new_n1006_ & ~new_n1779_;
  assign new_n1782_ = ~new_n1780_ & ~new_n1781_;
  assign new_n1783_ = new_n1002_ & new_n1782_;
  assign new_n1784_ = ~new_n1002_ & ~new_n1782_;
  assign new_n1785_ = ~new_n1783_ & ~new_n1784_;
  assign new_n1786_ = ~new_n1776_ & new_n1785_;
  assign new_n1787_ = new_n1776_ & ~new_n1785_;
  assign new_n1788_ = ~new_n1786_ & ~new_n1787_;
  assign new_n1789_ = new_n1079_ & ~new_n1788_;
  assign new_n1790_ = ~new_n988_ & new_n1006_;
  assign new_n1791_ = new_n988_ & ~new_n1006_;
  assign new_n1792_ = ~new_n1790_ & ~new_n1791_;
  assign new_n1793_ = ~new_n1726_ & ~new_n1792_;
  assign new_n1794_ = new_n1726_ & new_n1792_;
  assign new_n1795_ = ~new_n1793_ & ~new_n1794_;
  assign new_n1796_ = ~new_n997_ & ~new_n1081_;
  assign new_n1797_ = new_n1008_ & ~new_n1083_;
  assign new_n1798_ = ~new_n1796_ & new_n1797_;
  assign new_n1799_ = new_n1796_ & ~new_n1797_;
  assign new_n1800_ = ~new_n1798_ & ~new_n1799_;
  assign new_n1801_ = ~new_n1795_ & new_n1800_;
  assign new_n1802_ = new_n1795_ & ~new_n1800_;
  assign new_n1803_ = ~new_n1801_ & ~new_n1802_;
  assign new_n1804_ = new_n1010_ & new_n1083_;
  assign new_n1805_ = new_n1012_ & ~new_n1804_;
  assign new_n1806_ = new_n1081_ & new_n1805_;
  assign new_n1807_ = ~new_n1777_ & ~new_n1806_;
  assign new_n1808_ = new_n1002_ & ~new_n1010_;
  assign new_n1809_ = ~new_n1002_ & new_n1010_;
  assign new_n1810_ = ~new_n1808_ & ~new_n1809_;
  assign new_n1811_ = ~new_n1807_ & new_n1810_;
  assign new_n1812_ = new_n1807_ & ~new_n1810_;
  assign new_n1813_ = ~new_n1811_ & ~new_n1812_;
  assign new_n1814_ = ~new_n1803_ & new_n1813_;
  assign new_n1815_ = new_n1803_ & ~new_n1813_;
  assign new_n1816_ = ~new_n1814_ & ~new_n1815_;
  assign new_n1817_ = ~new_n1079_ & ~new_n1816_;
  assign new_n1818_ = ~new_n1789_ & ~new_n1817_;
  assign new_n1819_ = new_n960_ & ~new_n966_;
  assign new_n1820_ = ~new_n960_ & new_n966_;
  assign new_n1821_ = ~new_n1819_ & ~new_n1820_;
  assign new_n1822_ = new_n976_ & new_n1821_;
  assign new_n1823_ = ~new_n976_ & ~new_n1821_;
  assign new_n1824_ = ~new_n1822_ & ~new_n1823_;
  assign new_n1825_ = ~new_n971_ & ~new_n980_;
  assign new_n1826_ = ~new_n981_ & ~new_n1825_;
  assign new_n1827_ = ~new_n978_ & ~new_n1826_;
  assign new_n1828_ = new_n978_ & new_n1826_;
  assign new_n1829_ = ~new_n1827_ & ~new_n1828_;
  assign new_n1830_ = new_n974_ & ~new_n1829_;
  assign new_n1831_ = ~new_n974_ & new_n1829_;
  assign new_n1832_ = ~new_n1830_ & ~new_n1831_;
  assign new_n1833_ = new_n1824_ & new_n1832_;
  assign new_n1834_ = ~new_n1824_ & ~new_n1832_;
  assign new_n1835_ = ~new_n1833_ & ~new_n1834_;
  assign new_n1836_ = new_n1088_ & new_n1835_;
  assign new_n1837_ = new_n976_ & ~new_n981_;
  assign new_n1838_ = ~new_n1821_ & ~new_n1837_;
  assign new_n1839_ = new_n1821_ & new_n1837_;
  assign new_n1840_ = ~new_n1838_ & ~new_n1839_;
  assign new_n1841_ = new_n983_ & new_n1826_;
  assign new_n1842_ = ~new_n983_ & ~new_n1826_;
  assign new_n1843_ = ~new_n1841_ & ~new_n1842_;
  assign new_n1844_ = ~new_n1608_ & new_n1843_;
  assign new_n1845_ = new_n1608_ & ~new_n1843_;
  assign new_n1846_ = ~new_n1844_ & ~new_n1845_;
  assign new_n1847_ = ~new_n1840_ & new_n1846_;
  assign new_n1848_ = new_n1840_ & ~new_n1846_;
  assign new_n1849_ = ~new_n1847_ & ~new_n1848_;
  assign new_n1850_ = ~new_n1088_ & ~new_n1849_;
  assign new_n1851_ = ~new_n1836_ & ~new_n1850_;
  assign new_n1852_ = ~new_n1818_ & ~new_n1851_;
  assign new_n1853_ = new_n1818_ & new_n1851_;
  assign \1_n1150  = ~new_n1852_ & ~new_n1853_;
  assign new_n1855_ = ~new_n1058_ & ~new_n1069_;
  assign new_n1856_ = ~new_n1057_ & new_n1855_;
  assign new_n1857_ = new_n1057_ & ~new_n1855_;
  assign \1_n1178  = ~new_n1856_ & ~new_n1857_;
  assign new_n1859_ = ~new_n960_ & new_n1090_;
  assign \1_n1202  = ~new_n1091_ & ~new_n1859_;
  assign new_n1861_ = ~new_n997_ & new_n1079_;
  assign new_n1862_ = ~new_n1796_ & ~new_n1861_;
  assign new_n1863_ = new_n1002_ & new_n1862_;
  assign new_n1864_ = ~new_n1002_ & ~new_n1862_;
  assign \1_n1239  = ~new_n1863_ & ~new_n1864_;
  assign new_n1866_ = new_n1057_ & new_n1069_;
  assign new_n1867_ = new_n1060_ & ~new_n1866_;
  assign new_n1868_ = ~new_n1052_ & ~new_n1867_;
  assign new_n1869_ = new_n1052_ & new_n1867_;
  assign \1_n1301  = new_n1868_ | new_n1869_;
  assign new_n1871_ = \2_n1239  & \2_n312 ;
  assign new_n1872_ = ~\2_n1239  & \2_n307 ;
  assign new_n1873_ = ~new_n1871_ & ~new_n1872_;
  assign new_n1874_ = \2_n222  & new_n1873_;
  assign new_n1875_ = ~\2_n222  & ~new_n1873_;
  assign new_n1876_ = ~new_n1874_ & ~new_n1875_;
  assign new_n1877_ = \2_n1239  & \2_n1609 ;
  assign new_n1878_ = ~\2_n1239  & \2_n54 ;
  assign new_n1879_ = ~new_n1877_ & ~new_n1878_;
  assign new_n1880_ = \2_n608  & new_n1879_;
  assign new_n1881_ = ~\2_n608  & ~new_n1879_;
  assign new_n1882_ = ~new_n1880_ & ~new_n1881_;
  assign new_n1883_ = \2_n1239  & \2_n310 ;
  assign new_n1884_ = \2_n1175  & ~\2_n1239 ;
  assign new_n1885_ = ~new_n1883_ & ~new_n1884_;
  assign new_n1886_ = \2_n1071  & new_n1885_;
  assign new_n1887_ = ~\2_n1071  & ~new_n1885_;
  assign new_n1888_ = ~new_n1886_ & ~new_n1887_;
  assign new_n1889_ = new_n1882_ & new_n1888_;
  assign new_n1890_ = \2_n1239  & \2_n219 ;
  assign new_n1891_ = ~\2_n1239  & \2_n409 ;
  assign new_n1892_ = ~new_n1890_ & ~new_n1891_;
  assign new_n1893_ = \2_n45  & new_n1892_;
  assign new_n1894_ = ~\2_n45  & ~new_n1892_;
  assign new_n1895_ = ~new_n1893_ & ~new_n1894_;
  assign new_n1896_ = ~\2_n1239  & \2_n510 ;
  assign new_n1897_ = \2_n1205  & ~\2_n1239 ;
  assign new_n1898_ = new_n1896_ & ~new_n1897_;
  assign new_n1899_ = ~new_n1896_ & new_n1897_;
  assign new_n1900_ = ~new_n1898_ & ~new_n1899_;
  assign new_n1901_ = \2_n1239  & \2_n1569 ;
  assign new_n1902_ = ~\2_n1239  & \2_n1250 ;
  assign new_n1903_ = ~new_n1901_ & ~new_n1902_;
  assign new_n1904_ = \2_n695  & ~new_n1903_;
  assign new_n1905_ = ~\2_n695  & new_n1903_;
  assign new_n1906_ = ~new_n1904_ & ~new_n1905_;
  assign new_n1907_ = new_n1900_ & ~new_n1906_;
  assign new_n1908_ = new_n1895_ & new_n1907_;
  assign new_n1909_ = new_n1889_ & new_n1908_;
  assign new_n1910_ = \2_n545  & new_n1909_;
  assign new_n1911_ = new_n1888_ & new_n1894_;
  assign new_n1912_ = new_n1882_ & new_n1911_;
  assign new_n1913_ = ~\2_n695  & ~new_n1903_;
  assign new_n1914_ = new_n1895_ & new_n1913_;
  assign new_n1915_ = new_n1889_ & new_n1914_;
  assign new_n1916_ = ~new_n1912_ & ~new_n1915_;
  assign new_n1917_ = new_n1882_ & new_n1887_;
  assign new_n1918_ = ~new_n1881_ & ~new_n1917_;
  assign new_n1919_ = new_n1898_ & ~new_n1906_;
  assign new_n1920_ = new_n1895_ & new_n1919_;
  assign new_n1921_ = new_n1889_ & new_n1920_;
  assign new_n1922_ = new_n1918_ & ~new_n1921_;
  assign new_n1923_ = new_n1916_ & new_n1922_;
  assign new_n1924_ = ~new_n1910_ & new_n1923_;
  assign new_n1925_ = ~new_n1876_ & new_n1924_;
  assign new_n1926_ = new_n1876_ & ~new_n1924_;
  assign \2_n1006  = ~new_n1925_ & ~new_n1926_;
  assign new_n1928_ = \2_n380  & \2_n701 ;
  assign \2_n1050  = \2_n1361  | ~new_n1928_;
  assign new_n1930_ = \2_n1239  & \2_n598 ;
  assign new_n1931_ = ~\2_n1239  & \2_n1647 ;
  assign new_n1932_ = ~new_n1930_ & ~new_n1931_;
  assign new_n1933_ = \2_n1446  & new_n1932_;
  assign new_n1934_ = ~\2_n1446  & ~new_n1932_;
  assign new_n1935_ = ~new_n1933_ & ~new_n1934_;
  assign new_n1936_ = \2_n1239  & \2_n1415 ;
  assign new_n1937_ = ~\2_n1239  & \2_n1246 ;
  assign new_n1938_ = ~new_n1936_ & ~new_n1937_;
  assign new_n1939_ = ~\2_n1345  & ~new_n1938_;
  assign new_n1940_ = \2_n1345  & new_n1938_;
  assign new_n1941_ = ~new_n1939_ & ~new_n1940_;
  assign new_n1942_ = \2_n1239  & \2_n1350 ;
  assign new_n1943_ = ~\2_n1239  & \2_n262 ;
  assign new_n1944_ = ~new_n1942_ & ~new_n1943_;
  assign new_n1945_ = ~\2_n1301  & ~new_n1944_;
  assign new_n1946_ = \2_n1239  & \2_n676 ;
  assign new_n1947_ = \2_n1154  & ~\2_n1239 ;
  assign new_n1948_ = ~new_n1946_ & ~new_n1947_;
  assign new_n1949_ = ~\2_n1566  & ~new_n1948_;
  assign new_n1950_ = \2_n1301  & new_n1944_;
  assign new_n1951_ = ~new_n1945_ & ~new_n1950_;
  assign new_n1952_ = new_n1949_ & new_n1951_;
  assign new_n1953_ = ~new_n1945_ & ~new_n1952_;
  assign new_n1954_ = \2_n1239  & \2_n1289 ;
  assign new_n1955_ = \2_n1193  & ~\2_n1239 ;
  assign new_n1956_ = ~new_n1954_ & ~new_n1955_;
  assign new_n1957_ = ~\2_n920  & ~new_n1956_;
  assign new_n1958_ = \2_n1566  & new_n1948_;
  assign new_n1959_ = ~new_n1949_ & ~new_n1958_;
  assign new_n1960_ = new_n1957_ & new_n1959_;
  assign new_n1961_ = new_n1951_ & new_n1960_;
  assign new_n1962_ = \2_n1239  & \2_n244 ;
  assign new_n1963_ = ~\2_n1239  & \2_n641 ;
  assign new_n1964_ = ~new_n1962_ & ~new_n1963_;
  assign new_n1965_ = ~\2_n293  & ~new_n1964_;
  assign new_n1966_ = \2_n920  & new_n1956_;
  assign new_n1967_ = ~new_n1957_ & ~new_n1966_;
  assign new_n1968_ = new_n1965_ & new_n1967_;
  assign new_n1969_ = new_n1959_ & new_n1968_;
  assign new_n1970_ = new_n1951_ & new_n1969_;
  assign new_n1971_ = ~new_n1961_ & ~new_n1970_;
  assign new_n1972_ = new_n1953_ & new_n1971_;
  assign new_n1973_ = \2_n293  & new_n1964_;
  assign new_n1974_ = ~new_n1965_ & ~new_n1973_;
  assign new_n1975_ = new_n1967_ & new_n1974_;
  assign new_n1976_ = new_n1959_ & new_n1975_;
  assign new_n1977_ = new_n1951_ & new_n1976_;
  assign new_n1978_ = \2_n1239  & \2_n251 ;
  assign new_n1979_ = \2_n1172  & ~\2_n1239 ;
  assign new_n1980_ = ~new_n1978_ & ~new_n1979_;
  assign new_n1981_ = \2_n408  & new_n1980_;
  assign new_n1982_ = ~\2_n408  & ~new_n1980_;
  assign new_n1983_ = ~new_n1981_ & ~new_n1982_;
  assign new_n1984_ = \2_n1239  & \2_n790 ;
  assign new_n1985_ = ~\2_n1239  & \2_n1521 ;
  assign new_n1986_ = ~new_n1984_ & ~new_n1985_;
  assign new_n1987_ = ~\2_n823  & ~new_n1986_;
  assign new_n1988_ = \2_n1239  & \2_n1516 ;
  assign new_n1989_ = ~\2_n1239  & \2_n710 ;
  assign new_n1990_ = ~new_n1988_ & ~new_n1989_;
  assign new_n1991_ = \2_n1476  & new_n1990_;
  assign new_n1992_ = ~\2_n1476  & ~new_n1990_;
  assign new_n1993_ = ~new_n1991_ & ~new_n1992_;
  assign new_n1994_ = new_n1987_ & new_n1993_;
  assign new_n1995_ = new_n1983_ & new_n1994_;
  assign new_n1996_ = \2_n1239  & \2_n1576 ;
  assign new_n1997_ = ~\2_n1239  & \2_n1283 ;
  assign new_n1998_ = ~new_n1996_ & ~new_n1997_;
  assign new_n1999_ = ~\2_n153  & ~new_n1998_;
  assign new_n2000_ = \2_n823  & new_n1986_;
  assign new_n2001_ = ~new_n1987_ & ~new_n2000_;
  assign new_n2002_ = new_n1999_ & new_n2001_;
  assign new_n2003_ = new_n1983_ & new_n1993_;
  assign new_n2004_ = new_n2002_ & new_n2003_;
  assign new_n2005_ = ~new_n1995_ & ~new_n2004_;
  assign new_n2006_ = new_n1983_ & new_n1992_;
  assign new_n2007_ = ~new_n1982_ & ~new_n2006_;
  assign new_n2008_ = \2_n1239  & \2_n82 ;
  assign new_n2009_ = \2_n1061  & ~\2_n1239 ;
  assign new_n2010_ = ~new_n2008_ & ~new_n2009_;
  assign new_n2011_ = ~\2_n1401  & ~new_n2010_;
  assign new_n2012_ = \2_n153  & new_n1998_;
  assign new_n2013_ = ~new_n1999_ & ~new_n2012_;
  assign new_n2014_ = new_n2011_ & new_n2013_;
  assign new_n2015_ = new_n2001_ & new_n2014_;
  assign new_n2016_ = new_n2003_ & new_n2015_;
  assign new_n2017_ = new_n2007_ & ~new_n2016_;
  assign new_n2018_ = new_n2005_ & new_n2017_;
  assign new_n2019_ = new_n1977_ & ~new_n2018_;
  assign new_n2020_ = new_n1972_ & ~new_n2019_;
  assign new_n2021_ = \2_n1401  & new_n2010_;
  assign new_n2022_ = ~new_n2011_ & ~new_n2021_;
  assign new_n2023_ = new_n2013_ & new_n2022_;
  assign new_n2024_ = new_n2001_ & new_n2023_;
  assign new_n2025_ = new_n2003_ & new_n2024_;
  assign new_n2026_ = new_n1977_ & new_n2025_;
  assign new_n2027_ = \2_n1239  & \2_n645 ;
  assign new_n2028_ = ~\2_n1239  & \2_n87 ;
  assign new_n2029_ = ~new_n2027_ & ~new_n2028_;
  assign new_n2030_ = \2_n374  & new_n2029_;
  assign new_n2031_ = ~\2_n374  & ~new_n2029_;
  assign new_n2032_ = ~new_n2030_ & ~new_n2031_;
  assign new_n2033_ = \2_n1239  & \2_n268 ;
  assign new_n2034_ = ~\2_n1239  & \2_n600 ;
  assign new_n2035_ = ~new_n2033_ & ~new_n2034_;
  assign new_n2036_ = \2_n567  & ~new_n2035_;
  assign new_n2037_ = ~\2_n567  & new_n2035_;
  assign new_n2038_ = ~new_n2036_ & ~new_n2037_;
  assign new_n2039_ = new_n2032_ & ~new_n2038_;
  assign new_n2040_ = \2_n1239  & \2_n1393 ;
  assign new_n2041_ = ~\2_n1239  & \2_n254 ;
  assign new_n2042_ = ~new_n2040_ & ~new_n2041_;
  assign new_n2043_ = \2_n1463  & new_n2042_;
  assign new_n2044_ = ~\2_n1463  & ~new_n2042_;
  assign new_n2045_ = ~new_n2043_ & ~new_n2044_;
  assign new_n2046_ = new_n1876_ & new_n2045_;
  assign new_n2047_ = new_n2039_ & new_n2046_;
  assign new_n2048_ = new_n1910_ & new_n2047_;
  assign new_n2049_ = ~\2_n567  & ~new_n2035_;
  assign new_n2050_ = new_n2032_ & new_n2049_;
  assign new_n2051_ = ~new_n2031_ & ~new_n2050_;
  assign new_n2052_ = ~new_n2038_ & new_n2044_;
  assign new_n2053_ = new_n2032_ & new_n2052_;
  assign new_n2054_ = new_n1875_ & new_n2045_;
  assign new_n2055_ = ~new_n2038_ & new_n2054_;
  assign new_n2056_ = new_n2032_ & new_n2055_;
  assign new_n2057_ = ~new_n2053_ & ~new_n2056_;
  assign new_n2058_ = new_n2051_ & new_n2057_;
  assign new_n2059_ = ~new_n1923_ & new_n2047_;
  assign new_n2060_ = new_n2058_ & ~new_n2059_;
  assign new_n2061_ = ~new_n2048_ & new_n2060_;
  assign new_n2062_ = new_n2026_ & ~new_n2061_;
  assign new_n2063_ = new_n2020_ & ~new_n2062_;
  assign new_n2064_ = new_n1941_ & ~new_n2063_;
  assign new_n2065_ = ~new_n1939_ & ~new_n2064_;
  assign new_n2066_ = ~new_n1935_ & new_n2065_;
  assign new_n2067_ = new_n1935_ & ~new_n2065_;
  assign \2_n1051  = ~new_n2066_ & ~new_n2067_;
  assign new_n2069_ = \2_n545  & new_n1900_;
  assign new_n2070_ = ~new_n1906_ & new_n2069_;
  assign new_n2071_ = new_n1895_ & new_n2070_;
  assign new_n2072_ = ~new_n1914_ & ~new_n1920_;
  assign new_n2073_ = ~new_n1894_ & new_n2072_;
  assign new_n2074_ = ~new_n2071_ & new_n2073_;
  assign new_n2075_ = new_n1888_ & ~new_n2074_;
  assign new_n2076_ = ~new_n1888_ & new_n2074_;
  assign \2_n1058  = ~new_n2075_ & ~new_n2076_;
  assign new_n2078_ = ~new_n1965_ & ~new_n1967_;
  assign new_n2079_ = ~new_n1924_ & new_n2047_;
  assign new_n2080_ = new_n2058_ & ~new_n2079_;
  assign new_n2081_ = new_n2025_ & ~new_n2080_;
  assign new_n2082_ = new_n2018_ & ~new_n2081_;
  assign new_n2083_ = ~new_n1968_ & new_n2082_;
  assign new_n2084_ = ~new_n2078_ & new_n2083_;
  assign new_n2085_ = ~new_n1965_ & ~new_n1974_;
  assign new_n2086_ = new_n1967_ & new_n2085_;
  assign new_n2087_ = ~new_n1967_ & ~new_n2085_;
  assign new_n2088_ = ~new_n2086_ & ~new_n2087_;
  assign new_n2089_ = ~new_n2082_ & ~new_n2088_;
  assign \2_n1060  = new_n2084_ | new_n2089_;
  assign new_n2091_ = ~new_n2022_ & new_n2080_;
  assign new_n2092_ = new_n2022_ & ~new_n2080_;
  assign \2_n1063  = ~new_n2091_ & ~new_n2092_;
  assign new_n2094_ = \2_n11  & \2_n984 ;
  assign new_n2095_ = \2_n1239  & ~\2_n1435 ;
  assign new_n2096_ = ~new_n2094_ & ~new_n2095_;
  assign new_n2097_ = \2_n318  & ~new_n2096_;
  assign new_n2098_ = ~\2_n318  & new_n2096_;
  assign new_n2099_ = ~new_n2097_ & ~new_n2098_;
  assign new_n2100_ = \2_n1239  & \2_n58 ;
  assign new_n2101_ = ~\2_n1239  & \2_n1443 ;
  assign new_n2102_ = ~new_n2100_ & ~new_n2101_;
  assign new_n2103_ = ~\2_n1616  & ~new_n2102_;
  assign new_n2104_ = \2_n1239  & \2_n1474 ;
  assign new_n2105_ = ~\2_n1239  & \2_n1506 ;
  assign new_n2106_ = ~new_n2104_ & ~new_n2105_;
  assign new_n2107_ = \2_n1592  & new_n2106_;
  assign new_n2108_ = ~\2_n1592  & ~new_n2106_;
  assign new_n2109_ = ~new_n2107_ & ~new_n2108_;
  assign new_n2110_ = new_n2103_ & new_n2109_;
  assign new_n2111_ = new_n2099_ & new_n2110_;
  assign new_n2112_ = \2_n1616  & new_n2102_;
  assign new_n2113_ = ~new_n2103_ & ~new_n2112_;
  assign new_n2114_ = new_n1934_ & new_n2113_;
  assign new_n2115_ = new_n2099_ & new_n2109_;
  assign new_n2116_ = new_n2114_ & new_n2115_;
  assign new_n2117_ = ~new_n2111_ & ~new_n2116_;
  assign new_n2118_ = new_n2099_ & new_n2108_;
  assign new_n2119_ = ~new_n2098_ & ~new_n2118_;
  assign new_n2120_ = new_n1935_ & new_n1939_;
  assign new_n2121_ = new_n2113_ & new_n2120_;
  assign new_n2122_ = new_n2115_ & new_n2121_;
  assign new_n2123_ = new_n2119_ & ~new_n2122_;
  assign new_n2124_ = new_n2117_ & new_n2123_;
  assign new_n2125_ = \2_n1239  & ~\2_n905 ;
  assign new_n2126_ = ~new_n2094_ & ~new_n2125_;
  assign new_n2127_ = ~\2_n399  & new_n2126_;
  assign new_n2128_ = \2_n1239  & ~\2_n1278 ;
  assign new_n2129_ = ~new_n2094_ & ~new_n2128_;
  assign new_n2130_ = ~\2_n980  & new_n2129_;
  assign new_n2131_ = \2_n399  & ~new_n2126_;
  assign new_n2132_ = ~new_n2127_ & ~new_n2131_;
  assign new_n2133_ = new_n2130_ & new_n2132_;
  assign new_n2134_ = ~new_n2127_ & ~new_n2133_;
  assign new_n2135_ = \2_n1239  & ~\2_n220 ;
  assign new_n2136_ = ~new_n2094_ & ~new_n2135_;
  assign new_n2137_ = \2_n1263  & new_n2136_;
  assign new_n2138_ = ~\2_n1263  & ~new_n2136_;
  assign new_n2139_ = ~new_n2137_ & ~new_n2138_;
  assign new_n2140_ = \2_n1239  & ~\2_n391 ;
  assign new_n2141_ = ~new_n2094_ & ~new_n2140_;
  assign new_n2142_ = \2_n346  & new_n2141_;
  assign new_n2143_ = ~\2_n346  & ~new_n2141_;
  assign new_n2144_ = ~new_n2142_ & ~new_n2143_;
  assign new_n2145_ = new_n2139_ & ~new_n2144_;
  assign new_n2146_ = ~new_n2139_ & new_n2144_;
  assign new_n2147_ = ~new_n2145_ & ~new_n2146_;
  assign new_n2148_ = new_n2134_ & new_n2147_;
  assign new_n2149_ = ~new_n2134_ & ~new_n2147_;
  assign new_n2150_ = ~new_n2148_ & ~new_n2149_;
  assign new_n2151_ = \2_n980  & ~new_n2129_;
  assign new_n2152_ = ~new_n2130_ & ~new_n2151_;
  assign new_n2153_ = new_n2132_ & new_n2152_;
  assign new_n2154_ = ~new_n2132_ & ~new_n2152_;
  assign new_n2155_ = ~new_n2153_ & ~new_n2154_;
  assign new_n2156_ = ~\2_n346  & new_n2141_;
  assign new_n2157_ = new_n2127_ & ~new_n2144_;
  assign new_n2158_ = ~new_n2156_ & ~new_n2157_;
  assign new_n2159_ = new_n2133_ & ~new_n2144_;
  assign new_n2160_ = new_n2158_ & ~new_n2159_;
  assign new_n2161_ = ~new_n2130_ & new_n2160_;
  assign new_n2162_ = new_n2130_ & ~new_n2160_;
  assign new_n2163_ = ~new_n2161_ & ~new_n2162_;
  assign new_n2164_ = new_n2155_ & new_n2163_;
  assign new_n2165_ = ~new_n2155_ & ~new_n2163_;
  assign new_n2166_ = ~new_n2164_ & ~new_n2165_;
  assign new_n2167_ = ~new_n2150_ & new_n2166_;
  assign new_n2168_ = new_n2150_ & ~new_n2166_;
  assign new_n2169_ = ~new_n2167_ & ~new_n2168_;
  assign new_n2170_ = new_n2124_ & ~new_n2169_;
  assign new_n2171_ = new_n2134_ & ~new_n2153_;
  assign new_n2172_ = new_n2147_ & new_n2171_;
  assign new_n2173_ = ~new_n2147_ & ~new_n2171_;
  assign new_n2174_ = ~new_n2172_ & ~new_n2173_;
  assign new_n2175_ = ~new_n2130_ & ~new_n2152_;
  assign new_n2176_ = ~new_n2144_ & new_n2153_;
  assign new_n2177_ = new_n2160_ & ~new_n2176_;
  assign new_n2178_ = ~new_n2175_ & ~new_n2177_;
  assign new_n2179_ = new_n2175_ & new_n2177_;
  assign new_n2180_ = ~new_n2178_ & ~new_n2179_;
  assign new_n2181_ = new_n2155_ & new_n2180_;
  assign new_n2182_ = ~new_n2155_ & ~new_n2180_;
  assign new_n2183_ = ~new_n2181_ & ~new_n2182_;
  assign new_n2184_ = ~new_n2174_ & new_n2183_;
  assign new_n2185_ = new_n2174_ & ~new_n2183_;
  assign new_n2186_ = ~new_n2184_ & ~new_n2185_;
  assign new_n2187_ = ~new_n2124_ & new_n2186_;
  assign new_n2188_ = ~new_n2170_ & ~new_n2187_;
  assign new_n2189_ = new_n2063_ & ~new_n2188_;
  assign new_n2190_ = new_n1935_ & new_n1941_;
  assign new_n2191_ = new_n2113_ & new_n2190_;
  assign new_n2192_ = new_n2115_ & new_n2191_;
  assign new_n2193_ = new_n2124_ & ~new_n2192_;
  assign new_n2194_ = ~new_n2186_ & ~new_n2193_;
  assign new_n2195_ = new_n2169_ & new_n2193_;
  assign new_n2196_ = ~new_n2063_ & ~new_n2195_;
  assign new_n2197_ = ~new_n2194_ & new_n2196_;
  assign new_n2198_ = ~new_n2189_ & ~new_n2197_;
  assign new_n2199_ = ~new_n1935_ & ~new_n2113_;
  assign new_n2200_ = new_n1935_ & new_n2113_;
  assign new_n2201_ = ~new_n2199_ & ~new_n2200_;
  assign new_n2202_ = ~new_n2108_ & ~new_n2110_;
  assign new_n2203_ = ~new_n2114_ & ~new_n2121_;
  assign new_n2204_ = new_n2109_ & ~new_n2203_;
  assign new_n2205_ = new_n2202_ & ~new_n2204_;
  assign new_n2206_ = ~new_n1941_ & ~new_n2205_;
  assign new_n2207_ = new_n1941_ & new_n2205_;
  assign new_n2208_ = ~new_n2206_ & ~new_n2207_;
  assign new_n2209_ = new_n2201_ & new_n2208_;
  assign new_n2210_ = ~new_n2201_ & ~new_n2208_;
  assign new_n2211_ = ~new_n2209_ & ~new_n2210_;
  assign new_n2212_ = ~new_n2103_ & new_n2203_;
  assign new_n2213_ = ~new_n1939_ & ~new_n2212_;
  assign new_n2214_ = new_n1939_ & new_n2212_;
  assign new_n2215_ = ~new_n2213_ & ~new_n2214_;
  assign new_n2216_ = ~new_n1934_ & ~new_n2120_;
  assign new_n2217_ = ~new_n2099_ & ~new_n2109_;
  assign new_n2218_ = ~new_n2115_ & ~new_n2217_;
  assign new_n2219_ = new_n2216_ & new_n2218_;
  assign new_n2220_ = ~new_n2216_ & ~new_n2218_;
  assign new_n2221_ = ~new_n2219_ & ~new_n2220_;
  assign new_n2222_ = new_n2215_ & new_n2221_;
  assign new_n2223_ = ~new_n2215_ & ~new_n2221_;
  assign new_n2224_ = ~new_n2222_ & ~new_n2223_;
  assign new_n2225_ = ~new_n2211_ & new_n2224_;
  assign new_n2226_ = new_n2211_ & ~new_n2224_;
  assign new_n2227_ = ~new_n2225_ & ~new_n2226_;
  assign new_n2228_ = new_n2063_ & new_n2227_;
  assign new_n2229_ = ~new_n1939_ & ~new_n1941_;
  assign new_n2230_ = ~new_n2191_ & new_n2212_;
  assign new_n2231_ = ~new_n2229_ & ~new_n2230_;
  assign new_n2232_ = new_n2229_ & new_n2230_;
  assign new_n2233_ = ~new_n2231_ & ~new_n2232_;
  assign new_n2234_ = ~new_n1941_ & ~new_n2218_;
  assign new_n2235_ = new_n1941_ & new_n2218_;
  assign new_n2236_ = ~new_n2234_ & ~new_n2235_;
  assign new_n2237_ = ~new_n2190_ & new_n2216_;
  assign new_n2238_ = new_n2109_ & new_n2191_;
  assign new_n2239_ = new_n2205_ & ~new_n2238_;
  assign new_n2240_ = new_n2237_ & new_n2239_;
  assign new_n2241_ = ~new_n2237_ & ~new_n2239_;
  assign new_n2242_ = ~new_n2240_ & ~new_n2241_;
  assign new_n2243_ = ~new_n2236_ & new_n2242_;
  assign new_n2244_ = new_n2236_ & ~new_n2242_;
  assign new_n2245_ = ~new_n2243_ & ~new_n2244_;
  assign new_n2246_ = ~new_n2233_ & new_n2245_;
  assign new_n2247_ = new_n2233_ & ~new_n2245_;
  assign new_n2248_ = ~new_n2246_ & ~new_n2247_;
  assign new_n2249_ = ~new_n2201_ & new_n2248_;
  assign new_n2250_ = new_n2201_ & ~new_n2248_;
  assign new_n2251_ = ~new_n2063_ & ~new_n2250_;
  assign new_n2252_ = ~new_n2249_ & new_n2251_;
  assign new_n2253_ = ~new_n2228_ & ~new_n2252_;
  assign new_n2254_ = new_n2198_ & ~new_n2253_;
  assign new_n2255_ = ~new_n2198_ & new_n2253_;
  assign \2_n1065  = ~new_n2254_ & ~new_n2255_;
  assign new_n2257_ = new_n1974_ & ~new_n2082_;
  assign new_n2258_ = ~new_n1974_ & new_n2082_;
  assign \2_n112  = ~new_n2257_ & ~new_n2258_;
  assign new_n2260_ = \2_n156  & \2_n487 ;
  assign new_n2261_ = \2_n986  & ~new_n2260_;
  assign new_n2262_ = \2_n156  & \2_n200 ;
  assign new_n2263_ = \2_n986  & ~new_n2262_;
  assign new_n2264_ = ~new_n2261_ & ~new_n2263_;
  assign new_n2265_ = \2_n986  & new_n2260_;
  assign new_n2266_ = ~\2_n986  & ~new_n2260_;
  assign new_n2267_ = ~new_n2265_ & ~new_n2266_;
  assign new_n2268_ = \2_n986  & new_n2262_;
  assign new_n2269_ = ~\2_n986  & ~new_n2262_;
  assign new_n2270_ = ~new_n2268_ & ~new_n2269_;
  assign new_n2271_ = ~new_n2267_ & ~new_n2270_;
  assign new_n2272_ = \2_n1239  & ~\2_n582 ;
  assign new_n2273_ = ~new_n2094_ & ~new_n2272_;
  assign new_n2274_ = ~\2_n1470  & new_n2273_;
  assign new_n2275_ = \2_n1239  & ~\2_n1500 ;
  assign new_n2276_ = ~new_n2094_ & ~new_n2275_;
  assign new_n2277_ = ~\2_n138  & new_n2276_;
  assign new_n2278_ = \2_n1470  & ~new_n2273_;
  assign new_n2279_ = ~new_n2274_ & ~new_n2278_;
  assign new_n2280_ = new_n2277_ & new_n2279_;
  assign new_n2281_ = ~new_n2274_ & ~new_n2280_;
  assign new_n2282_ = \2_n138  & ~new_n2276_;
  assign new_n2283_ = ~new_n2277_ & ~new_n2282_;
  assign new_n2284_ = \2_n1239  & ~\2_n477 ;
  assign new_n2285_ = ~new_n2094_ & ~new_n2284_;
  assign new_n2286_ = ~\2_n769  & new_n2285_;
  assign new_n2287_ = ~\2_n1191  & \2_n1239 ;
  assign new_n2288_ = ~new_n2094_ & ~new_n2287_;
  assign new_n2289_ = ~\2_n626  & new_n2288_;
  assign new_n2290_ = \2_n769  & ~new_n2285_;
  assign new_n2291_ = ~new_n2286_ & ~new_n2290_;
  assign new_n2292_ = new_n2289_ & new_n2291_;
  assign new_n2293_ = ~new_n2286_ & ~new_n2292_;
  assign new_n2294_ = new_n2283_ & ~new_n2293_;
  assign new_n2295_ = new_n2279_ & new_n2294_;
  assign new_n2296_ = new_n2279_ & new_n2283_;
  assign new_n2297_ = \2_n1239  & ~\2_n430 ;
  assign new_n2298_ = ~new_n2094_ & ~new_n2297_;
  assign new_n2299_ = ~\2_n1656  & new_n2298_;
  assign new_n2300_ = \2_n626  & ~new_n2288_;
  assign new_n2301_ = ~new_n2289_ & ~new_n2300_;
  assign new_n2302_ = new_n2299_ & new_n2301_;
  assign new_n2303_ = new_n2291_ & new_n2302_;
  assign new_n2304_ = new_n2296_ & new_n2303_;
  assign new_n2305_ = ~new_n2295_ & ~new_n2304_;
  assign new_n2306_ = new_n2281_ & new_n2305_;
  assign new_n2307_ = \2_n1656  & ~new_n2298_;
  assign new_n2308_ = ~new_n2299_ & ~new_n2307_;
  assign new_n2309_ = new_n2301_ & new_n2308_;
  assign new_n2310_ = new_n2291_ & new_n2309_;
  assign new_n2311_ = new_n2296_ & new_n2310_;
  assign new_n2312_ = ~new_n2139_ & new_n2176_;
  assign new_n2313_ = new_n2192_ & new_n2312_;
  assign new_n2314_ = new_n2026_ & new_n2313_;
  assign new_n2315_ = ~new_n2060_ & new_n2314_;
  assign new_n2316_ = new_n2048_ & new_n2313_;
  assign new_n2317_ = new_n2026_ & new_n2316_;
  assign new_n2318_ = ~\2_n1263  & new_n2136_;
  assign new_n2319_ = ~new_n2139_ & new_n2156_;
  assign new_n2320_ = ~new_n2318_ & ~new_n2319_;
  assign new_n2321_ = ~new_n2139_ & new_n2157_;
  assign new_n2322_ = ~new_n2139_ & new_n2159_;
  assign new_n2323_ = ~new_n2321_ & ~new_n2322_;
  assign new_n2324_ = new_n2320_ & new_n2323_;
  assign new_n2325_ = ~new_n2124_ & new_n2312_;
  assign new_n2326_ = new_n2324_ & ~new_n2325_;
  assign new_n2327_ = ~new_n2020_ & new_n2313_;
  assign new_n2328_ = new_n2326_ & ~new_n2327_;
  assign new_n2329_ = ~new_n2317_ & new_n2328_;
  assign new_n2330_ = ~new_n2315_ & new_n2329_;
  assign new_n2331_ = new_n2311_ & ~new_n2330_;
  assign new_n2332_ = new_n2306_ & ~new_n2331_;
  assign new_n2333_ = new_n2271_ & ~new_n2332_;
  assign \2_n1186  = ~new_n2264_ | new_n2333_;
  assign new_n2335_ = ~new_n2044_ & ~new_n2054_;
  assign new_n2336_ = new_n2038_ & new_n2335_;
  assign new_n2337_ = ~new_n2038_ & ~new_n2335_;
  assign new_n2338_ = ~new_n2336_ & ~new_n2337_;
  assign new_n2339_ = new_n1924_ & new_n2338_;
  assign new_n2340_ = ~new_n2046_ & new_n2335_;
  assign new_n2341_ = ~new_n2038_ & ~new_n2340_;
  assign new_n2342_ = new_n2038_ & new_n2340_;
  assign new_n2343_ = ~new_n1924_ & ~new_n2342_;
  assign new_n2344_ = ~new_n2341_ & new_n2343_;
  assign \2_n1195  = new_n2339_ | new_n2344_;
  assign new_n2346_ = \2_n156  & ~\2_n559 ;
  assign new_n2347_ = \2_n156  & ~\2_n589 ;
  assign new_n2348_ = new_n2346_ & new_n2347_;
  assign new_n2349_ = \2_n986  & ~new_n2348_;
  assign new_n2350_ = ~\2_n986  & new_n2347_;
  assign new_n2351_ = \2_n986  & new_n2346_;
  assign new_n2352_ = ~\2_n986  & ~new_n2346_;
  assign new_n2353_ = ~new_n2351_ & ~new_n2352_;
  assign new_n2354_ = ~new_n2350_ & ~new_n2353_;
  assign new_n2355_ = \2_n1239  & ~\2_n223 ;
  assign new_n2356_ = ~new_n2094_ & ~new_n2355_;
  assign new_n2357_ = \2_n1239  & ~\2_n1470 ;
  assign new_n2358_ = ~\2_n1239  & \2_n300 ;
  assign new_n2359_ = ~new_n2357_ & ~new_n2358_;
  assign new_n2360_ = new_n2356_ & ~new_n2359_;
  assign new_n2361_ = \2_n1239  & ~\2_n138 ;
  assign new_n2362_ = ~\2_n1239  & \2_n561 ;
  assign new_n2363_ = ~new_n2361_ & ~new_n2362_;
  assign new_n2364_ = \2_n1239  & ~\2_n86 ;
  assign new_n2365_ = ~new_n2094_ & ~new_n2364_;
  assign new_n2366_ = ~new_n2356_ & ~new_n2359_;
  assign new_n2367_ = new_n2356_ & new_n2359_;
  assign new_n2368_ = ~new_n2366_ & ~new_n2367_;
  assign new_n2369_ = new_n2365_ & ~new_n2368_;
  assign new_n2370_ = ~new_n2363_ & new_n2369_;
  assign new_n2371_ = ~new_n2360_ & ~new_n2370_;
  assign new_n2372_ = \2_n1239  & ~\2_n1299 ;
  assign new_n2373_ = ~new_n2094_ & ~new_n2372_;
  assign new_n2374_ = \2_n1239  & ~\2_n769 ;
  assign new_n2375_ = ~\2_n1239  & \2_n879 ;
  assign new_n2376_ = ~new_n2374_ & ~new_n2375_;
  assign new_n2377_ = new_n2373_ & ~new_n2376_;
  assign new_n2378_ = ~new_n2363_ & ~new_n2365_;
  assign new_n2379_ = new_n2363_ & new_n2365_;
  assign new_n2380_ = ~new_n2378_ & ~new_n2379_;
  assign new_n2381_ = ~new_n2368_ & ~new_n2380_;
  assign new_n2382_ = new_n2377_ & new_n2381_;
  assign new_n2383_ = new_n2371_ & ~new_n2382_;
  assign new_n2384_ = \2_n1239  & ~\2_n1502 ;
  assign new_n2385_ = ~new_n2094_ & ~new_n2384_;
  assign new_n2386_ = ~new_n2368_ & new_n2385_;
  assign new_n2387_ = \2_n1239  & ~\2_n626 ;
  assign new_n2388_ = ~\2_n1239  & \2_n143 ;
  assign new_n2389_ = ~new_n2387_ & ~new_n2388_;
  assign new_n2390_ = new_n2373_ & new_n2376_;
  assign new_n2391_ = ~new_n2373_ & ~new_n2376_;
  assign new_n2392_ = ~new_n2390_ & ~new_n2391_;
  assign new_n2393_ = ~new_n2380_ & ~new_n2392_;
  assign new_n2394_ = ~new_n2389_ & new_n2393_;
  assign new_n2395_ = new_n2386_ & new_n2394_;
  assign new_n2396_ = ~new_n2368_ & ~new_n2392_;
  assign new_n2397_ = ~new_n2385_ & ~new_n2389_;
  assign new_n2398_ = new_n2385_ & new_n2389_;
  assign new_n2399_ = ~new_n2397_ & ~new_n2398_;
  assign new_n2400_ = \2_n1239  & ~\2_n1656 ;
  assign new_n2401_ = ~\2_n1239  & \2_n663 ;
  assign new_n2402_ = ~new_n2400_ & ~new_n2401_;
  assign new_n2403_ = ~new_n2094_ & ~new_n2402_;
  assign new_n2404_ = ~new_n2380_ & new_n2403_;
  assign new_n2405_ = ~new_n2399_ & new_n2404_;
  assign new_n2406_ = new_n2396_ & new_n2405_;
  assign new_n2407_ = ~new_n2395_ & ~new_n2406_;
  assign new_n2408_ = new_n2383_ & new_n2407_;
  assign new_n2409_ = new_n2094_ & new_n2402_;
  assign new_n2410_ = ~new_n2399_ & ~new_n2403_;
  assign new_n2411_ = ~new_n2409_ & new_n2410_;
  assign new_n2412_ = ~new_n2380_ & new_n2411_;
  assign new_n2413_ = new_n2396_ & new_n2412_;
  assign new_n2414_ = \2_n1239  & ~\2_n787 ;
  assign new_n2415_ = ~new_n2094_ & ~new_n2414_;
  assign new_n2416_ = \2_n1239  & ~\2_n399 ;
  assign new_n2417_ = \2_n1164  & ~\2_n1239 ;
  assign new_n2418_ = ~new_n2416_ & ~new_n2417_;
  assign new_n2419_ = new_n2415_ & ~new_n2418_;
  assign new_n2420_ = \2_n1239  & ~\2_n727 ;
  assign new_n2421_ = ~new_n2094_ & ~new_n2420_;
  assign new_n2422_ = \2_n1239  & ~\2_n1263 ;
  assign new_n2423_ = ~\2_n1239  & \2_n40 ;
  assign new_n2424_ = ~new_n2422_ & ~new_n2423_;
  assign new_n2425_ = ~new_n2421_ & ~new_n2424_;
  assign new_n2426_ = new_n2421_ & new_n2424_;
  assign new_n2427_ = ~new_n2425_ & ~new_n2426_;
  assign new_n2428_ = \2_n1239  & ~\2_n346 ;
  assign new_n2429_ = ~\2_n1239  & \2_n489 ;
  assign new_n2430_ = ~new_n2428_ & ~new_n2429_;
  assign new_n2431_ = \2_n1239  & ~\2_n94 ;
  assign new_n2432_ = ~new_n2094_ & ~new_n2431_;
  assign new_n2433_ = ~new_n2430_ & ~new_n2432_;
  assign new_n2434_ = new_n2430_ & new_n2432_;
  assign new_n2435_ = ~new_n2433_ & ~new_n2434_;
  assign new_n2436_ = ~new_n2427_ & ~new_n2435_;
  assign new_n2437_ = new_n2419_ & new_n2436_;
  assign new_n2438_ = \2_n1239  & ~\2_n609 ;
  assign new_n2439_ = ~new_n2094_ & ~new_n2438_;
  assign new_n2440_ = new_n2415_ & new_n2418_;
  assign new_n2441_ = ~new_n2415_ & ~new_n2418_;
  assign new_n2442_ = ~new_n2440_ & ~new_n2441_;
  assign new_n2443_ = new_n2439_ & ~new_n2442_;
  assign new_n2444_ = \2_n1239  & ~\2_n980 ;
  assign new_n2445_ = ~\2_n1239  & \2_n71 ;
  assign new_n2446_ = ~new_n2444_ & ~new_n2445_;
  assign new_n2447_ = new_n2436_ & ~new_n2446_;
  assign new_n2448_ = new_n2443_ & new_n2447_;
  assign new_n2449_ = ~new_n2437_ & ~new_n2448_;
  assign new_n2450_ = new_n2421_ & ~new_n2424_;
  assign new_n2451_ = ~new_n2427_ & new_n2432_;
  assign new_n2452_ = ~new_n2430_ & new_n2451_;
  assign new_n2453_ = ~new_n2439_ & ~new_n2446_;
  assign new_n2454_ = new_n2439_ & new_n2446_;
  assign new_n2455_ = ~new_n2453_ & ~new_n2454_;
  assign new_n2456_ = ~new_n2442_ & ~new_n2455_;
  assign new_n2457_ = new_n2436_ & new_n2456_;
  assign new_n2458_ = \2_n1239  & \2_n52 ;
  assign new_n2459_ = ~new_n2101_ & ~new_n2458_;
  assign new_n2460_ = \2_n1239  & ~\2_n1616 ;
  assign new_n2461_ = ~\2_n1239  & \2_n1418 ;
  assign new_n2462_ = ~new_n2460_ & ~new_n2461_;
  assign new_n2463_ = ~new_n2459_ & ~new_n2462_;
  assign new_n2464_ = \2_n1239  & ~\2_n1592 ;
  assign new_n2465_ = ~\2_n1239  & \2_n1305 ;
  assign new_n2466_ = ~new_n2464_ & ~new_n2465_;
  assign new_n2467_ = \2_n1239  & \2_n953 ;
  assign new_n2468_ = ~new_n2105_ & ~new_n2467_;
  assign new_n2469_ = ~new_n2466_ & new_n2468_;
  assign new_n2470_ = new_n2466_ & ~new_n2468_;
  assign new_n2471_ = ~new_n2469_ & ~new_n2470_;
  assign new_n2472_ = \2_n1239  & ~\2_n839 ;
  assign new_n2473_ = ~new_n2094_ & ~new_n2472_;
  assign new_n2474_ = \2_n1239  & ~\2_n318 ;
  assign new_n2475_ = ~\2_n1239  & \2_n1523 ;
  assign new_n2476_ = ~new_n2474_ & ~new_n2475_;
  assign new_n2477_ = ~new_n2473_ & ~new_n2476_;
  assign new_n2478_ = new_n2473_ & new_n2476_;
  assign new_n2479_ = ~new_n2477_ & ~new_n2478_;
  assign new_n2480_ = ~new_n2471_ & ~new_n2479_;
  assign new_n2481_ = new_n2463_ & new_n2480_;
  assign new_n2482_ = \2_n1239  & ~\2_n1446 ;
  assign new_n2483_ = \2_n1156  & ~\2_n1239 ;
  assign new_n2484_ = ~new_n2482_ & ~new_n2483_;
  assign new_n2485_ = new_n2459_ & ~new_n2462_;
  assign new_n2486_ = ~new_n2459_ & new_n2462_;
  assign new_n2487_ = ~new_n2485_ & ~new_n2486_;
  assign new_n2488_ = ~new_n2484_ & ~new_n2487_;
  assign new_n2489_ = \2_n1239  & \2_n1428 ;
  assign new_n2490_ = ~new_n1931_ & ~new_n2489_;
  assign new_n2491_ = new_n2480_ & ~new_n2490_;
  assign new_n2492_ = new_n2488_ & new_n2491_;
  assign new_n2493_ = ~new_n2481_ & ~new_n2492_;
  assign new_n2494_ = new_n2473_ & ~new_n2476_;
  assign new_n2495_ = ~new_n2468_ & ~new_n2479_;
  assign new_n2496_ = ~new_n2466_ & new_n2495_;
  assign new_n2497_ = ~new_n2494_ & ~new_n2496_;
  assign new_n2498_ = ~new_n2471_ & ~new_n2487_;
  assign new_n2499_ = ~new_n2484_ & new_n2490_;
  assign new_n2500_ = new_n2484_ & ~new_n2490_;
  assign new_n2501_ = ~new_n2499_ & ~new_n2500_;
  assign new_n2502_ = \2_n1239  & \2_n607 ;
  assign new_n2503_ = ~new_n1937_ & ~new_n2502_;
  assign new_n2504_ = \2_n1239  & ~\2_n1345 ;
  assign new_n2505_ = ~\2_n1239  & \2_n969 ;
  assign new_n2506_ = ~new_n2504_ & ~new_n2505_;
  assign new_n2507_ = ~new_n2503_ & ~new_n2506_;
  assign new_n2508_ = ~new_n2479_ & new_n2507_;
  assign new_n2509_ = ~new_n2501_ & new_n2508_;
  assign new_n2510_ = new_n2498_ & new_n2509_;
  assign new_n2511_ = new_n2497_ & ~new_n2510_;
  assign new_n2512_ = new_n2493_ & new_n2511_;
  assign new_n2513_ = new_n2457_ & ~new_n2512_;
  assign new_n2514_ = ~new_n2452_ & ~new_n2513_;
  assign new_n2515_ = ~new_n2450_ & new_n2514_;
  assign new_n2516_ = new_n2449_ & new_n2515_;
  assign new_n2517_ = new_n2503_ & new_n2506_;
  assign new_n2518_ = ~new_n2501_ & ~new_n2507_;
  assign new_n2519_ = ~new_n2517_ & new_n2518_;
  assign new_n2520_ = new_n2457_ & new_n2519_;
  assign new_n2521_ = ~new_n2487_ & new_n2520_;
  assign new_n2522_ = new_n2480_ & new_n2521_;
  assign new_n2523_ = \2_n1239  & \2_n885 ;
  assign new_n2524_ = ~new_n1955_ & ~new_n2523_;
  assign new_n2525_ = \2_n1239  & ~\2_n920 ;
  assign new_n2526_ = \2_n107  & ~\2_n1239 ;
  assign new_n2527_ = ~new_n2525_ & ~new_n2526_;
  assign new_n2528_ = ~new_n2524_ & ~new_n2527_;
  assign new_n2529_ = \2_n1239  & \2_n376 ;
  assign new_n2530_ = ~new_n1943_ & ~new_n2529_;
  assign new_n2531_ = \2_n1239  & ~\2_n1301 ;
  assign new_n2532_ = ~\2_n1239  & \2_n779 ;
  assign new_n2533_ = ~new_n2531_ & ~new_n2532_;
  assign new_n2534_ = new_n2530_ & ~new_n2533_;
  assign new_n2535_ = ~new_n2530_ & new_n2533_;
  assign new_n2536_ = ~new_n2534_ & ~new_n2535_;
  assign new_n2537_ = \2_n1239  & ~\2_n1566 ;
  assign new_n2538_ = ~\2_n1239  & \2_n507 ;
  assign new_n2539_ = ~new_n2537_ & ~new_n2538_;
  assign new_n2540_ = \2_n1239  & \2_n273 ;
  assign new_n2541_ = ~new_n1947_ & ~new_n2540_;
  assign new_n2542_ = ~new_n2539_ & new_n2541_;
  assign new_n2543_ = new_n2539_ & ~new_n2541_;
  assign new_n2544_ = ~new_n2542_ & ~new_n2543_;
  assign new_n2545_ = ~new_n2536_ & ~new_n2544_;
  assign new_n2546_ = new_n2528_ & new_n2545_;
  assign new_n2547_ = \2_n1239  & ~\2_n293 ;
  assign new_n2548_ = ~\2_n1239  & \2_n1448 ;
  assign new_n2549_ = ~new_n2547_ & ~new_n2548_;
  assign new_n2550_ = new_n2524_ & ~new_n2527_;
  assign new_n2551_ = ~new_n2524_ & new_n2527_;
  assign new_n2552_ = ~new_n2550_ & ~new_n2551_;
  assign new_n2553_ = ~new_n2549_ & ~new_n2552_;
  assign new_n2554_ = \2_n1239  & \2_n50 ;
  assign new_n2555_ = ~new_n1963_ & ~new_n2554_;
  assign new_n2556_ = new_n2545_ & ~new_n2555_;
  assign new_n2557_ = new_n2553_ & new_n2556_;
  assign new_n2558_ = ~new_n2546_ & ~new_n2557_;
  assign new_n2559_ = ~new_n2530_ & ~new_n2533_;
  assign new_n2560_ = ~new_n2536_ & ~new_n2539_;
  assign new_n2561_ = ~new_n2541_ & new_n2560_;
  assign new_n2562_ = ~new_n2549_ & new_n2555_;
  assign new_n2563_ = new_n2549_ & ~new_n2555_;
  assign new_n2564_ = ~new_n2562_ & ~new_n2563_;
  assign new_n2565_ = ~new_n2552_ & ~new_n2564_;
  assign new_n2566_ = new_n2545_ & new_n2565_;
  assign new_n2567_ = \2_n1239  & \2_n734 ;
  assign new_n2568_ = ~new_n1979_ & ~new_n2567_;
  assign new_n2569_ = \2_n1239  & ~\2_n408 ;
  assign new_n2570_ = \2_n1152  & ~\2_n1239 ;
  assign new_n2571_ = ~new_n2569_ & ~new_n2570_;
  assign new_n2572_ = ~new_n2568_ & ~new_n2571_;
  assign new_n2573_ = \2_n1239  & ~\2_n1476 ;
  assign new_n2574_ = ~\2_n1239  & \2_n1386 ;
  assign new_n2575_ = ~new_n2573_ & ~new_n2574_;
  assign new_n2576_ = \2_n1239  & \2_n1586 ;
  assign new_n2577_ = ~new_n1989_ & ~new_n2576_;
  assign new_n2578_ = new_n2568_ & ~new_n2571_;
  assign new_n2579_ = ~new_n2568_ & new_n2571_;
  assign new_n2580_ = ~new_n2578_ & ~new_n2579_;
  assign new_n2581_ = ~new_n2577_ & ~new_n2580_;
  assign new_n2582_ = ~new_n2575_ & new_n2581_;
  assign new_n2583_ = ~new_n2572_ & ~new_n2582_;
  assign new_n2584_ = \2_n1239  & ~\2_n153 ;
  assign new_n2585_ = ~\2_n1239  & \2_n1627 ;
  assign new_n2586_ = ~new_n2584_ & ~new_n2585_;
  assign new_n2587_ = \2_n1239  & \2_n77 ;
  assign new_n2588_ = ~new_n1985_ & ~new_n2587_;
  assign new_n2589_ = \2_n1239  & ~\2_n823 ;
  assign new_n2590_ = ~\2_n1239  & \2_n882 ;
  assign new_n2591_ = ~new_n2589_ & ~new_n2590_;
  assign new_n2592_ = new_n2588_ & ~new_n2591_;
  assign new_n2593_ = ~new_n2588_ & new_n2591_;
  assign new_n2594_ = ~new_n2592_ & ~new_n2593_;
  assign new_n2595_ = ~new_n2586_ & ~new_n2594_;
  assign new_n2596_ = \2_n1114  & \2_n1239 ;
  assign new_n2597_ = ~new_n1997_ & ~new_n2596_;
  assign new_n2598_ = ~new_n2575_ & new_n2577_;
  assign new_n2599_ = new_n2575_ & ~new_n2577_;
  assign new_n2600_ = ~new_n2598_ & ~new_n2599_;
  assign new_n2601_ = ~new_n2580_ & ~new_n2600_;
  assign new_n2602_ = ~new_n2597_ & new_n2601_;
  assign new_n2603_ = new_n2595_ & new_n2602_;
  assign new_n2604_ = new_n2583_ & ~new_n2603_;
  assign new_n2605_ = ~new_n2588_ & ~new_n2591_;
  assign new_n2606_ = new_n2601_ & new_n2605_;
  assign new_n2607_ = ~new_n2594_ & ~new_n2600_;
  assign new_n2608_ = ~new_n2586_ & new_n2597_;
  assign new_n2609_ = new_n2586_ & ~new_n2597_;
  assign new_n2610_ = ~new_n2608_ & ~new_n2609_;
  assign new_n2611_ = \2_n1239  & \2_n344 ;
  assign new_n2612_ = ~new_n2009_ & ~new_n2611_;
  assign new_n2613_ = \2_n1239  & ~\2_n1401 ;
  assign new_n2614_ = \2_n1227  & ~\2_n1239 ;
  assign new_n2615_ = ~new_n2613_ & ~new_n2614_;
  assign new_n2616_ = ~new_n2612_ & ~new_n2615_;
  assign new_n2617_ = ~new_n2580_ & new_n2616_;
  assign new_n2618_ = ~new_n2610_ & new_n2617_;
  assign new_n2619_ = new_n2607_ & new_n2618_;
  assign new_n2620_ = ~new_n2606_ & ~new_n2619_;
  assign new_n2621_ = new_n2604_ & new_n2620_;
  assign new_n2622_ = new_n2566_ & ~new_n2621_;
  assign new_n2623_ = ~new_n2561_ & ~new_n2622_;
  assign new_n2624_ = ~new_n2559_ & new_n2623_;
  assign new_n2625_ = new_n2558_ & new_n2624_;
  assign new_n2626_ = new_n2522_ & ~new_n2625_;
  assign new_n2627_ = new_n2516_ & ~new_n2626_;
  assign new_n2628_ = ~new_n2580_ & ~new_n2594_;
  assign new_n2629_ = new_n2612_ & new_n2615_;
  assign new_n2630_ = ~new_n2610_ & ~new_n2616_;
  assign new_n2631_ = ~new_n2629_ & new_n2630_;
  assign new_n2632_ = new_n2566_ & new_n2631_;
  assign new_n2633_ = ~new_n2600_ & new_n2632_;
  assign new_n2634_ = new_n2628_ & new_n2633_;
  assign new_n2635_ = \2_n1239  & \2_n392 ;
  assign new_n2636_ = ~new_n1878_ & ~new_n2635_;
  assign new_n2637_ = \2_n1239  & ~\2_n608 ;
  assign new_n2638_ = ~\2_n1239  & \2_n742 ;
  assign new_n2639_ = ~new_n2637_ & ~new_n2638_;
  assign new_n2640_ = new_n2636_ & new_n2639_;
  assign new_n2641_ = ~new_n2636_ & ~new_n2639_;
  assign new_n2642_ = ~new_n2640_ & ~new_n2641_;
  assign new_n2643_ = \2_n690  & new_n2642_;
  assign new_n2644_ = ~\2_n1071  & \2_n1239 ;
  assign new_n2645_ = ~\2_n1239  & \2_n341 ;
  assign new_n2646_ = ~new_n2644_ & ~new_n2645_;
  assign new_n2647_ = \2_n1239  & \2_n671 ;
  assign new_n2648_ = ~new_n1884_ & ~new_n2647_;
  assign new_n2649_ = ~new_n2646_ & new_n2648_;
  assign new_n2650_ = new_n2646_ & ~new_n2648_;
  assign new_n2651_ = ~new_n2649_ & ~new_n2650_;
  assign new_n2652_ = \2_n1239  & \2_n29 ;
  assign new_n2653_ = ~new_n1891_ & ~new_n2652_;
  assign new_n2654_ = \2_n1239  & ~\2_n45 ;
  assign new_n2655_ = ~\2_n1239  & \2_n849 ;
  assign new_n2656_ = ~new_n2654_ & ~new_n2655_;
  assign new_n2657_ = new_n2653_ & ~new_n2656_;
  assign new_n2658_ = ~new_n2653_ & new_n2656_;
  assign new_n2659_ = ~new_n2657_ & ~new_n2658_;
  assign new_n2660_ = ~new_n2651_ & ~new_n2659_;
  assign new_n2661_ = ~\2_n1239  & \2_n729 ;
  assign new_n2662_ = ~\2_n1239  & ~new_n2661_;
  assign new_n2663_ = ~new_n1896_ & new_n2662_;
  assign new_n2664_ = new_n1896_ & ~new_n2662_;
  assign new_n2665_ = \2_n1239  & ~\2_n695 ;
  assign new_n2666_ = ~\2_n1239  & \2_n502 ;
  assign new_n2667_ = ~new_n2665_ & ~new_n2666_;
  assign new_n2668_ = \2_n1239  & \2_n778 ;
  assign new_n2669_ = ~new_n1902_ & ~new_n2668_;
  assign new_n2670_ = ~new_n2667_ & new_n2669_;
  assign new_n2671_ = new_n2667_ & ~new_n2669_;
  assign new_n2672_ = ~new_n2670_ & ~new_n2671_;
  assign new_n2673_ = ~new_n2664_ & ~new_n2672_;
  assign new_n2674_ = ~new_n2663_ & new_n2673_;
  assign new_n2675_ = \2_n1239  & \2_n1753 ;
  assign new_n2676_ = ~new_n2028_ & ~new_n2675_;
  assign new_n2677_ = \2_n1239  & ~\2_n374 ;
  assign new_n2678_ = ~\2_n1239  & \2_n755 ;
  assign new_n2679_ = ~new_n2677_ & ~new_n2678_;
  assign new_n2680_ = new_n2676_ & ~new_n2679_;
  assign new_n2681_ = ~new_n2676_ & new_n2679_;
  assign new_n2682_ = ~new_n2680_ & ~new_n2681_;
  assign new_n2683_ = \2_n1239  & ~\2_n567 ;
  assign new_n2684_ = ~\2_n1239  & \2_n936 ;
  assign new_n2685_ = ~new_n2683_ & ~new_n2684_;
  assign new_n2686_ = \2_n1239  & \2_n288 ;
  assign new_n2687_ = ~new_n2034_ & ~new_n2686_;
  assign new_n2688_ = ~new_n2685_ & new_n2687_;
  assign new_n2689_ = new_n2685_ & ~new_n2687_;
  assign new_n2690_ = ~new_n2688_ & ~new_n2689_;
  assign new_n2691_ = ~new_n2682_ & ~new_n2690_;
  assign new_n2692_ = \2_n1239  & \2_n416 ;
  assign new_n2693_ = ~new_n2041_ & ~new_n2692_;
  assign new_n2694_ = \2_n1239  & ~\2_n1463 ;
  assign new_n2695_ = ~\2_n1239  & \2_n159 ;
  assign new_n2696_ = ~new_n2694_ & ~new_n2695_;
  assign new_n2697_ = new_n2693_ & ~new_n2696_;
  assign new_n2698_ = ~new_n2693_ & new_n2696_;
  assign new_n2699_ = ~new_n2697_ & ~new_n2698_;
  assign new_n2700_ = \2_n1239  & ~\2_n222 ;
  assign new_n2701_ = ~\2_n1239  & \2_n243 ;
  assign new_n2702_ = ~new_n2700_ & ~new_n2701_;
  assign new_n2703_ = \2_n1239  & \2_n506 ;
  assign new_n2704_ = ~new_n1872_ & ~new_n2703_;
  assign new_n2705_ = ~new_n2702_ & new_n2704_;
  assign new_n2706_ = new_n2702_ & ~new_n2704_;
  assign new_n2707_ = ~new_n2705_ & ~new_n2706_;
  assign new_n2708_ = ~new_n2699_ & ~new_n2707_;
  assign new_n2709_ = new_n2691_ & new_n2708_;
  assign new_n2710_ = new_n2674_ & new_n2709_;
  assign new_n2711_ = new_n2660_ & new_n2710_;
  assign new_n2712_ = new_n2643_ & new_n2711_;
  assign new_n2713_ = new_n2522_ & new_n2712_;
  assign new_n2714_ = new_n2634_ & new_n2713_;
  assign new_n2715_ = ~new_n2693_ & ~new_n2696_;
  assign new_n2716_ = new_n2691_ & new_n2715_;
  assign new_n2717_ = ~new_n2699_ & ~new_n2702_;
  assign new_n2718_ = new_n2691_ & ~new_n2704_;
  assign new_n2719_ = new_n2717_ & new_n2718_;
  assign new_n2720_ = ~new_n2716_ & ~new_n2719_;
  assign new_n2721_ = ~new_n2676_ & ~new_n2679_;
  assign new_n2722_ = ~new_n2682_ & ~new_n2685_;
  assign new_n2723_ = ~new_n2687_ & new_n2722_;
  assign new_n2724_ = new_n2642_ & ~new_n2648_;
  assign new_n2725_ = ~new_n2646_ & new_n2724_;
  assign new_n2726_ = ~new_n2641_ & ~new_n2725_;
  assign new_n2727_ = ~new_n2659_ & ~new_n2667_;
  assign new_n2728_ = new_n2642_ & ~new_n2651_;
  assign new_n2729_ = ~new_n2669_ & new_n2728_;
  assign new_n2730_ = new_n2727_ & new_n2729_;
  assign new_n2731_ = new_n2726_ & ~new_n2730_;
  assign new_n2732_ = ~new_n2653_ & ~new_n2656_;
  assign new_n2733_ = new_n2728_ & new_n2732_;
  assign new_n2734_ = new_n2664_ & ~new_n2672_;
  assign new_n2735_ = new_n2642_ & new_n2734_;
  assign new_n2736_ = new_n2660_ & new_n2735_;
  assign new_n2737_ = ~new_n2733_ & ~new_n2736_;
  assign new_n2738_ = new_n2731_ & new_n2737_;
  assign new_n2739_ = new_n2709_ & ~new_n2738_;
  assign new_n2740_ = ~new_n2723_ & ~new_n2739_;
  assign new_n2741_ = ~new_n2721_ & new_n2740_;
  assign new_n2742_ = new_n2720_ & new_n2741_;
  assign new_n2743_ = new_n2522_ & ~new_n2742_;
  assign new_n2744_ = new_n2634_ & new_n2743_;
  assign new_n2745_ = ~new_n2714_ & ~new_n2744_;
  assign new_n2746_ = new_n2627_ & new_n2745_;
  assign new_n2747_ = new_n2413_ & ~new_n2746_;
  assign new_n2748_ = new_n2408_ & ~new_n2747_;
  assign new_n2749_ = new_n2354_ & ~new_n2748_;
  assign \2_n1211  = new_n2349_ | new_n2749_;
  assign new_n2751_ = \2_n284  & \2_n574 ;
  assign new_n2752_ = \2_n1520  & \2_n1613 ;
  assign \2_n126  = ~new_n2751_ | ~new_n2752_;
  assign new_n2754_ = new_n2285_ & ~new_n2288_;
  assign new_n2755_ = ~new_n2285_ & new_n2288_;
  assign new_n2756_ = ~new_n2754_ & ~new_n2755_;
  assign new_n2757_ = new_n2273_ & ~new_n2276_;
  assign new_n2758_ = ~new_n2273_ & new_n2276_;
  assign new_n2759_ = ~new_n2757_ & ~new_n2758_;
  assign new_n2760_ = ~new_n2756_ & new_n2759_;
  assign new_n2761_ = new_n2756_ & ~new_n2759_;
  assign new_n2762_ = ~new_n2760_ & ~new_n2761_;
  assign new_n2763_ = \2_n1239  & ~\2_n1626 ;
  assign new_n2764_ = ~new_n2094_ & ~new_n2763_;
  assign new_n2765_ = new_n2298_ & ~new_n2764_;
  assign new_n2766_ = ~new_n2298_ & new_n2764_;
  assign new_n2767_ = ~new_n2765_ & ~new_n2766_;
  assign new_n2768_ = \2_n1239  & ~\2_n775 ;
  assign new_n2769_ = ~new_n2094_ & ~new_n2768_;
  assign new_n2770_ = ~new_n2094_ & new_n2769_;
  assign new_n2771_ = new_n2094_ & ~new_n2769_;
  assign new_n2772_ = ~new_n2770_ & ~new_n2771_;
  assign new_n2773_ = ~new_n2767_ & new_n2772_;
  assign new_n2774_ = new_n2767_ & ~new_n2772_;
  assign new_n2775_ = ~new_n2773_ & ~new_n2774_;
  assign new_n2776_ = ~new_n2762_ & new_n2775_;
  assign new_n2777_ = new_n2762_ & ~new_n2775_;
  assign new_n2778_ = ~new_n2776_ & ~new_n2777_;
  assign new_n2779_ = \2_n117  & \2_n1239 ;
  assign new_n2780_ = \2_n1103  & ~\2_n1239 ;
  assign new_n2781_ = ~new_n2779_ & ~new_n2780_;
  assign new_n2782_ = new_n1938_ & ~new_n2781_;
  assign new_n2783_ = ~new_n1938_ & new_n2781_;
  assign new_n2784_ = ~new_n2782_ & ~new_n2783_;
  assign new_n2785_ = ~new_n1932_ & new_n2102_;
  assign new_n2786_ = new_n1932_ & ~new_n2102_;
  assign new_n2787_ = ~new_n2785_ & ~new_n2786_;
  assign new_n2788_ = ~new_n2784_ & new_n2787_;
  assign new_n2789_ = new_n2784_ & ~new_n2787_;
  assign new_n2790_ = ~new_n2788_ & ~new_n2789_;
  assign new_n2791_ = ~new_n2096_ & ~new_n2106_;
  assign new_n2792_ = new_n2096_ & new_n2106_;
  assign new_n2793_ = ~new_n2791_ & ~new_n2792_;
  assign new_n2794_ = ~new_n2790_ & new_n2793_;
  assign new_n2795_ = new_n2790_ & ~new_n2793_;
  assign new_n2796_ = ~new_n2794_ & ~new_n2795_;
  assign new_n2797_ = new_n2126_ & ~new_n2129_;
  assign new_n2798_ = ~new_n2126_ & new_n2129_;
  assign new_n2799_ = ~new_n2797_ & ~new_n2798_;
  assign new_n2800_ = new_n2136_ & ~new_n2141_;
  assign new_n2801_ = ~new_n2136_ & new_n2141_;
  assign new_n2802_ = ~new_n2800_ & ~new_n2801_;
  assign new_n2803_ = ~new_n2799_ & new_n2802_;
  assign new_n2804_ = new_n2799_ & ~new_n2802_;
  assign new_n2805_ = ~new_n2803_ & ~new_n2804_;
  assign new_n2806_ = ~new_n2796_ & new_n2805_;
  assign new_n2807_ = new_n2796_ & ~new_n2805_;
  assign new_n2808_ = ~new_n2806_ & ~new_n2807_;
  assign new_n2809_ = ~new_n2778_ & ~new_n2808_;
  assign new_n2810_ = \2_n1239  & \2_n314 ;
  assign new_n2811_ = \2_n1121  & ~\2_n1239 ;
  assign new_n2812_ = ~new_n2810_ & ~new_n2811_;
  assign new_n2813_ = new_n2010_ & ~new_n2812_;
  assign new_n2814_ = ~new_n2010_ & new_n2812_;
  assign new_n2815_ = ~new_n2813_ & ~new_n2814_;
  assign new_n2816_ = new_n1986_ & ~new_n1998_;
  assign new_n2817_ = ~new_n1986_ & new_n1998_;
  assign new_n2818_ = ~new_n2816_ & ~new_n2817_;
  assign new_n2819_ = ~new_n2815_ & new_n2818_;
  assign new_n2820_ = new_n2815_ & ~new_n2818_;
  assign new_n2821_ = ~new_n2819_ & ~new_n2820_;
  assign new_n2822_ = new_n1980_ & ~new_n1990_;
  assign new_n2823_ = ~new_n1980_ & new_n1990_;
  assign new_n2824_ = ~new_n2822_ & ~new_n2823_;
  assign new_n2825_ = ~new_n2821_ & new_n2824_;
  assign new_n2826_ = new_n2821_ & ~new_n2824_;
  assign new_n2827_ = ~new_n2825_ & ~new_n2826_;
  assign new_n2828_ = new_n1956_ & ~new_n1964_;
  assign new_n2829_ = ~new_n1956_ & new_n1964_;
  assign new_n2830_ = ~new_n2828_ & ~new_n2829_;
  assign new_n2831_ = new_n1944_ & ~new_n1948_;
  assign new_n2832_ = ~new_n1944_ & new_n1948_;
  assign new_n2833_ = ~new_n2831_ & ~new_n2832_;
  assign new_n2834_ = ~new_n2830_ & new_n2833_;
  assign new_n2835_ = new_n2830_ & ~new_n2833_;
  assign new_n2836_ = ~new_n2834_ & ~new_n2835_;
  assign new_n2837_ = ~new_n2827_ & new_n2836_;
  assign new_n2838_ = new_n2827_ & ~new_n2836_;
  assign new_n2839_ = ~new_n2837_ & ~new_n2838_;
  assign new_n2840_ = \2_n1239  & \2_n961 ;
  assign new_n2841_ = ~new_n1896_ & ~new_n2840_;
  assign new_n2842_ = \2_n1239  & \2_n1281 ;
  assign new_n2843_ = ~\2_n1239  & \2_n299 ;
  assign new_n2844_ = ~new_n2842_ & ~new_n2843_;
  assign new_n2845_ = new_n2841_ & ~new_n2844_;
  assign new_n2846_ = ~new_n2841_ & new_n2844_;
  assign new_n2847_ = ~new_n2845_ & ~new_n2846_;
  assign new_n2848_ = ~new_n1892_ & ~new_n1903_;
  assign new_n2849_ = new_n1892_ & new_n1903_;
  assign new_n2850_ = ~new_n2848_ & ~new_n2849_;
  assign new_n2851_ = ~new_n2847_ & ~new_n2850_;
  assign new_n2852_ = new_n2847_ & new_n2850_;
  assign new_n2853_ = ~new_n2851_ & ~new_n2852_;
  assign new_n2854_ = new_n1879_ & ~new_n1885_;
  assign new_n2855_ = ~new_n1879_ & new_n1885_;
  assign new_n2856_ = ~new_n2854_ & ~new_n2855_;
  assign new_n2857_ = ~new_n2853_ & new_n2856_;
  assign new_n2858_ = new_n2853_ & ~new_n2856_;
  assign new_n2859_ = ~new_n2857_ & ~new_n2858_;
  assign new_n2860_ = ~new_n1873_ & new_n2042_;
  assign new_n2861_ = new_n1873_ & ~new_n2042_;
  assign new_n2862_ = ~new_n2860_ & ~new_n2861_;
  assign new_n2863_ = ~new_n2029_ & ~new_n2035_;
  assign new_n2864_ = new_n2029_ & new_n2035_;
  assign new_n2865_ = ~new_n2863_ & ~new_n2864_;
  assign new_n2866_ = ~new_n2862_ & ~new_n2865_;
  assign new_n2867_ = new_n2862_ & new_n2865_;
  assign new_n2868_ = ~new_n2866_ & ~new_n2867_;
  assign new_n2869_ = ~new_n2859_ & new_n2868_;
  assign new_n2870_ = new_n2859_ & ~new_n2868_;
  assign new_n2871_ = ~new_n2869_ & ~new_n2870_;
  assign new_n2872_ = ~new_n2839_ & ~new_n2871_;
  assign \2_n1288  = ~new_n2809_ | ~new_n2872_;
  assign new_n2874_ = new_n2308_ & ~new_n2330_;
  assign new_n2875_ = ~new_n2299_ & ~new_n2874_;
  assign new_n2876_ = ~new_n2301_ & new_n2875_;
  assign new_n2877_ = new_n2301_ & ~new_n2875_;
  assign \2_n1302  = ~new_n2876_ & ~new_n2877_;
  assign new_n2879_ = ~new_n2712_ & new_n2742_;
  assign new_n2880_ = new_n2634_ & ~new_n2879_;
  assign \2_n1306  = ~new_n2625_ | new_n2880_;
  assign new_n2882_ = ~new_n2359_ & ~new_n2363_;
  assign new_n2883_ = new_n2359_ & new_n2363_;
  assign new_n2884_ = ~new_n2882_ & ~new_n2883_;
  assign new_n2885_ = ~new_n2376_ & ~new_n2389_;
  assign new_n2886_ = new_n2376_ & new_n2389_;
  assign new_n2887_ = ~new_n2885_ & ~new_n2886_;
  assign new_n2888_ = new_n2884_ & new_n2887_;
  assign new_n2889_ = ~new_n2884_ & ~new_n2887_;
  assign new_n2890_ = ~new_n2888_ & ~new_n2889_;
  assign new_n2891_ = ~\2_n1239  & \2_n1346 ;
  assign new_n2892_ = \2_n1239  & ~\2_n831 ;
  assign new_n2893_ = ~new_n2891_ & ~new_n2892_;
  assign new_n2894_ = new_n2402_ & ~new_n2893_;
  assign new_n2895_ = ~new_n2402_ & new_n2893_;
  assign new_n2896_ = ~new_n2894_ & ~new_n2895_;
  assign new_n2897_ = ~\2_n1239  & \2_n559 ;
  assign new_n2898_ = \2_n1239  & ~\2_n487 ;
  assign new_n2899_ = ~new_n2897_ & ~new_n2898_;
  assign new_n2900_ = ~\2_n1239  & \2_n589 ;
  assign new_n2901_ = \2_n1239  & ~\2_n200 ;
  assign new_n2902_ = ~new_n2900_ & ~new_n2901_;
  assign new_n2903_ = ~new_n2899_ & ~new_n2902_;
  assign new_n2904_ = new_n2899_ & new_n2902_;
  assign new_n2905_ = ~new_n2903_ & ~new_n2904_;
  assign new_n2906_ = ~new_n2896_ & new_n2905_;
  assign new_n2907_ = new_n2896_ & ~new_n2905_;
  assign new_n2908_ = ~new_n2906_ & ~new_n2907_;
  assign new_n2909_ = ~new_n2890_ & new_n2908_;
  assign new_n2910_ = new_n2890_ & ~new_n2908_;
  assign new_n2911_ = ~new_n2909_ & ~new_n2910_;
  assign new_n2912_ = new_n2424_ & ~new_n2430_;
  assign new_n2913_ = ~new_n2424_ & new_n2430_;
  assign new_n2914_ = ~new_n2912_ & ~new_n2913_;
  assign new_n2915_ = ~new_n2418_ & ~new_n2446_;
  assign new_n2916_ = new_n2418_ & new_n2446_;
  assign new_n2917_ = ~new_n2915_ & ~new_n2916_;
  assign new_n2918_ = ~new_n2914_ & new_n2917_;
  assign new_n2919_ = new_n2914_ & ~new_n2917_;
  assign new_n2920_ = ~new_n2918_ & ~new_n2919_;
  assign new_n2921_ = ~new_n2466_ & new_n2476_;
  assign new_n2922_ = new_n2466_ & ~new_n2476_;
  assign new_n2923_ = ~new_n2921_ & ~new_n2922_;
  assign new_n2924_ = new_n2462_ & ~new_n2484_;
  assign new_n2925_ = ~new_n2462_ & new_n2484_;
  assign new_n2926_ = ~new_n2924_ & ~new_n2925_;
  assign new_n2927_ = ~\2_n1239  & \2_n1644 ;
  assign new_n2928_ = \2_n1239  & ~\2_n21 ;
  assign new_n2929_ = ~new_n2927_ & ~new_n2928_;
  assign new_n2930_ = ~new_n2506_ & ~new_n2929_;
  assign new_n2931_ = new_n2506_ & new_n2929_;
  assign new_n2932_ = ~new_n2930_ & ~new_n2931_;
  assign new_n2933_ = ~new_n2926_ & new_n2932_;
  assign new_n2934_ = new_n2926_ & ~new_n2932_;
  assign new_n2935_ = ~new_n2933_ & ~new_n2934_;
  assign new_n2936_ = ~new_n2923_ & new_n2935_;
  assign new_n2937_ = new_n2923_ & ~new_n2935_;
  assign new_n2938_ = ~new_n2936_ & ~new_n2937_;
  assign new_n2939_ = ~new_n2920_ & new_n2938_;
  assign new_n2940_ = new_n2920_ & ~new_n2938_;
  assign new_n2941_ = ~new_n2939_ & ~new_n2940_;
  assign new_n2942_ = ~new_n2911_ & ~new_n2941_;
  assign new_n2943_ = new_n2533_ & ~new_n2539_;
  assign new_n2944_ = ~new_n2533_ & new_n2539_;
  assign new_n2945_ = ~new_n2943_ & ~new_n2944_;
  assign new_n2946_ = ~new_n2527_ & ~new_n2549_;
  assign new_n2947_ = new_n2527_ & new_n2549_;
  assign new_n2948_ = ~new_n2946_ & ~new_n2947_;
  assign new_n2949_ = ~new_n2945_ & new_n2948_;
  assign new_n2950_ = new_n2945_ & ~new_n2948_;
  assign new_n2951_ = ~new_n2949_ & ~new_n2950_;
  assign new_n2952_ = new_n2571_ & ~new_n2575_;
  assign new_n2953_ = ~new_n2571_ & new_n2575_;
  assign new_n2954_ = ~new_n2952_ & ~new_n2953_;
  assign new_n2955_ = ~new_n2586_ & new_n2591_;
  assign new_n2956_ = new_n2586_ & ~new_n2591_;
  assign new_n2957_ = ~new_n2955_ & ~new_n2956_;
  assign new_n2958_ = ~\2_n1239  & \2_n1750 ;
  assign new_n2959_ = \2_n1239  & ~\2_n947 ;
  assign new_n2960_ = ~new_n2958_ & ~new_n2959_;
  assign new_n2961_ = ~new_n2615_ & ~new_n2960_;
  assign new_n2962_ = new_n2615_ & new_n2960_;
  assign new_n2963_ = ~new_n2961_ & ~new_n2962_;
  assign new_n2964_ = ~new_n2957_ & new_n2963_;
  assign new_n2965_ = new_n2957_ & ~new_n2963_;
  assign new_n2966_ = ~new_n2964_ & ~new_n2965_;
  assign new_n2967_ = ~new_n2954_ & new_n2966_;
  assign new_n2968_ = new_n2954_ & ~new_n2966_;
  assign new_n2969_ = ~new_n2967_ & ~new_n2968_;
  assign new_n2970_ = ~new_n2951_ & new_n2969_;
  assign new_n2971_ = new_n2951_ & ~new_n2969_;
  assign new_n2972_ = ~new_n2970_ & ~new_n2971_;
  assign new_n2973_ = ~new_n2679_ & ~new_n2685_;
  assign new_n2974_ = new_n2679_ & new_n2685_;
  assign new_n2975_ = ~new_n2973_ & ~new_n2974_;
  assign new_n2976_ = ~new_n2696_ & ~new_n2702_;
  assign new_n2977_ = new_n2696_ & new_n2702_;
  assign new_n2978_ = ~new_n2976_ & ~new_n2977_;
  assign new_n2979_ = new_n2975_ & new_n2978_;
  assign new_n2980_ = ~new_n2975_ & ~new_n2978_;
  assign new_n2981_ = ~new_n2979_ & ~new_n2980_;
  assign new_n2982_ = new_n2639_ & ~new_n2646_;
  assign new_n2983_ = ~new_n2639_ & new_n2646_;
  assign new_n2984_ = ~new_n2982_ & ~new_n2983_;
  assign new_n2985_ = new_n2656_ & ~new_n2667_;
  assign new_n2986_ = ~new_n2656_ & new_n2667_;
  assign new_n2987_ = ~new_n2985_ & ~new_n2986_;
  assign new_n2988_ = ~\2_n1205  & \2_n1239 ;
  assign new_n2989_ = ~new_n2661_ & ~new_n2988_;
  assign new_n2990_ = ~\2_n1239  & \2_n155 ;
  assign new_n2991_ = ~\2_n1138  & \2_n1239 ;
  assign new_n2992_ = ~new_n2990_ & ~new_n2991_;
  assign new_n2993_ = ~new_n2989_ & ~new_n2992_;
  assign new_n2994_ = new_n2989_ & new_n2992_;
  assign new_n2995_ = ~new_n2993_ & ~new_n2994_;
  assign new_n2996_ = ~new_n2987_ & new_n2995_;
  assign new_n2997_ = new_n2987_ & ~new_n2995_;
  assign new_n2998_ = ~new_n2996_ & ~new_n2997_;
  assign new_n2999_ = ~new_n2984_ & new_n2998_;
  assign new_n3000_ = new_n2984_ & ~new_n2998_;
  assign new_n3001_ = ~new_n2999_ & ~new_n3000_;
  assign new_n3002_ = ~new_n2981_ & new_n3001_;
  assign new_n3003_ = new_n2981_ & ~new_n3001_;
  assign new_n3004_ = ~new_n3002_ & ~new_n3003_;
  assign new_n3005_ = ~new_n2972_ & ~new_n3004_;
  assign \2_n1322  = ~new_n2942_ | ~new_n3005_;
  assign new_n3007_ = ~new_n2270_ & ~new_n2332_;
  assign new_n3008_ = new_n2270_ & new_n2332_;
  assign \2_n1359  = ~new_n3007_ & ~new_n3008_;
  assign new_n3010_ = ~new_n2373_ & new_n2385_;
  assign new_n3011_ = new_n2373_ & ~new_n2385_;
  assign new_n3012_ = ~new_n3010_ & ~new_n3011_;
  assign new_n3013_ = ~new_n2356_ & ~new_n2365_;
  assign new_n3014_ = new_n2356_ & new_n2365_;
  assign new_n3015_ = ~new_n3013_ & ~new_n3014_;
  assign new_n3016_ = ~new_n3012_ & ~new_n3015_;
  assign new_n3017_ = new_n3012_ & new_n3015_;
  assign new_n3018_ = ~new_n3016_ & ~new_n3017_;
  assign new_n3019_ = \2_n1239  & ~\2_n56 ;
  assign new_n3020_ = ~new_n2094_ & ~new_n3019_;
  assign new_n3021_ = ~new_n2094_ & new_n3020_;
  assign new_n3022_ = new_n2094_ & ~new_n3020_;
  assign new_n3023_ = ~new_n3021_ & ~new_n3022_;
  assign new_n3024_ = \2_n1239  & ~\2_n1389 ;
  assign new_n3025_ = ~new_n2094_ & ~new_n3024_;
  assign new_n3026_ = \2_n1239  & ~\2_n246 ;
  assign new_n3027_ = ~new_n2094_ & ~new_n3026_;
  assign new_n3028_ = ~new_n3025_ & new_n3027_;
  assign new_n3029_ = new_n3025_ & ~new_n3027_;
  assign new_n3030_ = ~new_n3028_ & ~new_n3029_;
  assign new_n3031_ = ~new_n3023_ & new_n3030_;
  assign new_n3032_ = new_n3023_ & ~new_n3030_;
  assign new_n3033_ = ~new_n3031_ & ~new_n3032_;
  assign new_n3034_ = ~new_n3018_ & new_n3033_;
  assign new_n3035_ = new_n3018_ & ~new_n3033_;
  assign new_n3036_ = ~new_n3034_ & ~new_n3035_;
  assign new_n3037_ = \2_n1023  & \2_n1239 ;
  assign new_n3038_ = ~new_n2780_ & ~new_n3037_;
  assign new_n3039_ = new_n2503_ & ~new_n3038_;
  assign new_n3040_ = ~new_n2503_ & new_n3038_;
  assign new_n3041_ = ~new_n3039_ & ~new_n3040_;
  assign new_n3042_ = ~new_n2459_ & ~new_n2490_;
  assign new_n3043_ = new_n2459_ & new_n2490_;
  assign new_n3044_ = ~new_n3042_ & ~new_n3043_;
  assign new_n3045_ = ~new_n3041_ & ~new_n3044_;
  assign new_n3046_ = new_n3041_ & new_n3044_;
  assign new_n3047_ = ~new_n3045_ & ~new_n3046_;
  assign new_n3048_ = ~new_n2468_ & ~new_n2473_;
  assign new_n3049_ = new_n2468_ & new_n2473_;
  assign new_n3050_ = ~new_n3048_ & ~new_n3049_;
  assign new_n3051_ = ~new_n3047_ & new_n3050_;
  assign new_n3052_ = new_n3047_ & ~new_n3050_;
  assign new_n3053_ = ~new_n3051_ & ~new_n3052_;
  assign new_n3054_ = new_n2415_ & ~new_n2439_;
  assign new_n3055_ = ~new_n2415_ & new_n2439_;
  assign new_n3056_ = ~new_n3054_ & ~new_n3055_;
  assign new_n3057_ = ~new_n2421_ & new_n2432_;
  assign new_n3058_ = new_n2421_ & ~new_n2432_;
  assign new_n3059_ = ~new_n3057_ & ~new_n3058_;
  assign new_n3060_ = ~new_n3056_ & new_n3059_;
  assign new_n3061_ = new_n3056_ & ~new_n3059_;
  assign new_n3062_ = ~new_n3060_ & ~new_n3061_;
  assign new_n3063_ = ~new_n3053_ & new_n3062_;
  assign new_n3064_ = new_n3053_ & ~new_n3062_;
  assign new_n3065_ = ~new_n3063_ & ~new_n3064_;
  assign new_n3066_ = ~new_n3036_ & ~new_n3065_;
  assign new_n3067_ = \2_n1239  & \2_n560 ;
  assign new_n3068_ = ~new_n2811_ & ~new_n3067_;
  assign new_n3069_ = new_n2612_ & ~new_n3068_;
  assign new_n3070_ = ~new_n2612_ & new_n3068_;
  assign new_n3071_ = ~new_n3069_ & ~new_n3070_;
  assign new_n3072_ = ~new_n2588_ & ~new_n2597_;
  assign new_n3073_ = new_n2588_ & new_n2597_;
  assign new_n3074_ = ~new_n3072_ & ~new_n3073_;
  assign new_n3075_ = ~new_n3071_ & ~new_n3074_;
  assign new_n3076_ = new_n3071_ & new_n3074_;
  assign new_n3077_ = ~new_n3075_ & ~new_n3076_;
  assign new_n3078_ = ~new_n2568_ & ~new_n2577_;
  assign new_n3079_ = new_n2568_ & new_n2577_;
  assign new_n3080_ = ~new_n3078_ & ~new_n3079_;
  assign new_n3081_ = ~new_n3077_ & ~new_n3080_;
  assign new_n3082_ = new_n3077_ & new_n3080_;
  assign new_n3083_ = ~new_n3081_ & ~new_n3082_;
  assign new_n3084_ = ~new_n2524_ & ~new_n2555_;
  assign new_n3085_ = new_n2524_ & new_n2555_;
  assign new_n3086_ = ~new_n3084_ & ~new_n3085_;
  assign new_n3087_ = ~new_n2530_ & ~new_n2541_;
  assign new_n3088_ = new_n2530_ & new_n2541_;
  assign new_n3089_ = ~new_n3087_ & ~new_n3088_;
  assign new_n3090_ = new_n3086_ & ~new_n3089_;
  assign new_n3091_ = ~new_n3086_ & new_n3089_;
  assign new_n3092_ = ~new_n3090_ & ~new_n3091_;
  assign new_n3093_ = ~new_n3083_ & new_n3092_;
  assign new_n3094_ = new_n3083_ & ~new_n3092_;
  assign new_n3095_ = ~new_n3093_ & ~new_n3094_;
  assign new_n3096_ = \2_n1239  & \2_n1411 ;
  assign new_n3097_ = ~new_n1896_ & ~new_n3096_;
  assign new_n3098_ = \2_n1044  & \2_n1239 ;
  assign new_n3099_ = ~new_n2843_ & ~new_n3098_;
  assign new_n3100_ = new_n3097_ & ~new_n3099_;
  assign new_n3101_ = ~new_n3097_ & new_n3099_;
  assign new_n3102_ = ~new_n3100_ & ~new_n3101_;
  assign new_n3103_ = ~new_n2653_ & ~new_n2669_;
  assign new_n3104_ = new_n2653_ & new_n2669_;
  assign new_n3105_ = ~new_n3103_ & ~new_n3104_;
  assign new_n3106_ = ~new_n3102_ & ~new_n3105_;
  assign new_n3107_ = new_n3102_ & new_n3105_;
  assign new_n3108_ = ~new_n3106_ & ~new_n3107_;
  assign new_n3109_ = ~new_n2636_ & ~new_n2648_;
  assign new_n3110_ = new_n2636_ & new_n2648_;
  assign new_n3111_ = ~new_n3109_ & ~new_n3110_;
  assign new_n3112_ = ~new_n3108_ & ~new_n3111_;
  assign new_n3113_ = new_n3108_ & new_n3111_;
  assign new_n3114_ = ~new_n3112_ & ~new_n3113_;
  assign new_n3115_ = ~new_n2693_ & ~new_n2704_;
  assign new_n3116_ = new_n2693_ & new_n2704_;
  assign new_n3117_ = ~new_n3115_ & ~new_n3116_;
  assign new_n3118_ = ~new_n2676_ & ~new_n2687_;
  assign new_n3119_ = new_n2676_ & new_n2687_;
  assign new_n3120_ = ~new_n3118_ & ~new_n3119_;
  assign new_n3121_ = new_n3117_ & ~new_n3120_;
  assign new_n3122_ = ~new_n3117_ & new_n3120_;
  assign new_n3123_ = ~new_n3121_ & ~new_n3122_;
  assign new_n3124_ = ~new_n3114_ & new_n3123_;
  assign new_n3125_ = new_n3114_ & ~new_n3123_;
  assign new_n3126_ = ~new_n3124_ & ~new_n3125_;
  assign new_n3127_ = ~new_n3095_ & ~new_n3126_;
  assign \2_n1375  = ~new_n3066_ | ~new_n3127_;
  assign new_n3129_ = new_n2293_ & ~new_n2303_;
  assign new_n3130_ = new_n2301_ & new_n2874_;
  assign new_n3131_ = new_n2291_ & new_n3130_;
  assign new_n3132_ = new_n3129_ & ~new_n3131_;
  assign new_n3133_ = new_n2283_ & ~new_n3132_;
  assign new_n3134_ = ~new_n2283_ & new_n3132_;
  assign \2_n1391  = ~new_n3133_ & ~new_n3134_;
  assign new_n3136_ = ~new_n1898_ & ~new_n2069_;
  assign new_n3137_ = ~new_n1906_ & ~new_n3136_;
  assign new_n3138_ = new_n1906_ & new_n3136_;
  assign \2_n1420  = ~new_n3137_ & ~new_n3138_;
  assign new_n3140_ = ~new_n1875_ & ~new_n2045_;
  assign new_n3141_ = ~new_n2054_ & ~new_n3140_;
  assign new_n3142_ = new_n1924_ & new_n3141_;
  assign new_n3143_ = ~new_n1875_ & ~new_n1876_;
  assign new_n3144_ = new_n2045_ & ~new_n3143_;
  assign new_n3145_ = ~new_n2045_ & new_n3143_;
  assign new_n3146_ = ~new_n1924_ & ~new_n3145_;
  assign new_n3147_ = ~new_n3144_ & new_n3146_;
  assign \2_n1427  = new_n3142_ | new_n3147_;
  assign new_n3149_ = ~new_n1941_ & new_n2063_;
  assign \2_n1527  = ~new_n2064_ & ~new_n3149_;
  assign new_n3151_ = ~new_n2263_ & ~new_n2267_;
  assign new_n3152_ = new_n2263_ & new_n2267_;
  assign new_n3153_ = ~new_n3151_ & ~new_n3152_;
  assign new_n3154_ = new_n2332_ & ~new_n3153_;
  assign new_n3155_ = ~new_n2263_ & new_n2270_;
  assign new_n3156_ = ~new_n2267_ & ~new_n3155_;
  assign new_n3157_ = new_n2267_ & new_n3155_;
  assign new_n3158_ = ~new_n3156_ & ~new_n3157_;
  assign new_n3159_ = ~new_n2332_ & new_n3158_;
  assign \2_n1588  = new_n3154_ | new_n3159_;
  assign new_n3161_ = \2_n1040  & \2_n1054 ;
  assign new_n3162_ = \2_n1286  & \2_n593 ;
  assign \2_n1594  = ~new_n3161_ | ~new_n3162_;
  assign new_n3164_ = new_n2354_ & ~new_n2408_;
  assign new_n3165_ = new_n2354_ & new_n2413_;
  assign new_n3166_ = ~new_n2627_ & new_n3165_;
  assign new_n3167_ = ~new_n2349_ & ~new_n3166_;
  assign new_n3168_ = ~new_n3164_ & new_n3167_;
  assign new_n3169_ = new_n2714_ & new_n3165_;
  assign new_n3170_ = new_n2744_ & new_n3165_;
  assign new_n3171_ = ~new_n3169_ & ~new_n3170_;
  assign \2_n161  = ~new_n3168_ | ~new_n3171_;
  assign new_n3173_ = new_n1888_ & new_n1908_;
  assign new_n3174_ = \2_n545  & new_n3173_;
  assign new_n3175_ = ~new_n1887_ & ~new_n1911_;
  assign new_n3176_ = new_n1888_ & ~new_n2072_;
  assign new_n3177_ = new_n3175_ & ~new_n3176_;
  assign new_n3178_ = ~new_n3174_ & new_n3177_;
  assign new_n3179_ = ~new_n1882_ & new_n3178_;
  assign new_n3180_ = new_n1882_ & ~new_n3178_;
  assign \2_n1639  = ~new_n3179_ & ~new_n3180_;
  assign new_n3182_ = ~new_n2063_ & new_n2238_;
  assign new_n3183_ = new_n2205_ & ~new_n3182_;
  assign new_n3184_ = ~new_n2099_ & new_n3183_;
  assign new_n3185_ = new_n2099_ & ~new_n3183_;
  assign \2_n164  = ~new_n3184_ & ~new_n3185_;
  assign new_n3187_ = ~new_n1957_ & ~new_n1968_;
  assign new_n3188_ = new_n1959_ & ~new_n3187_;
  assign new_n3189_ = ~new_n1959_ & new_n3187_;
  assign new_n3190_ = new_n2082_ & ~new_n3189_;
  assign new_n3191_ = ~new_n3188_ & new_n3190_;
  assign new_n3192_ = ~new_n1975_ & new_n3187_;
  assign new_n3193_ = ~new_n1959_ & ~new_n3192_;
  assign new_n3194_ = new_n1959_ & new_n3192_;
  assign new_n3195_ = ~new_n3193_ & ~new_n3194_;
  assign new_n3196_ = ~new_n2082_ & ~new_n3195_;
  assign \2_n1687  = new_n3191_ | new_n3196_;
  assign new_n3198_ = \2_n581  & \2_n743 ;
  assign new_n3199_ = \2_n1095  & \2_n478 ;
  assign \2_n1752  = ~new_n3198_ | ~new_n3199_;
  assign new_n3201_ = ~new_n2063_ & new_n2192_;
  assign new_n3202_ = new_n2124_ & ~new_n3201_;
  assign new_n3203_ = ~new_n2152_ & new_n3202_;
  assign new_n3204_ = new_n2152_ & ~new_n3202_;
  assign \2_n181  = ~new_n3203_ & ~new_n3204_;
  assign new_n3206_ = ~new_n2289_ & ~new_n2302_;
  assign new_n3207_ = ~new_n3130_ & new_n3206_;
  assign new_n3208_ = ~new_n2291_ & new_n3207_;
  assign new_n3209_ = new_n2291_ & ~new_n3207_;
  assign \2_n216  = ~new_n3208_ & ~new_n3209_;
  assign new_n3211_ = ~new_n2139_ & ~new_n2160_;
  assign new_n3212_ = new_n2139_ & new_n2160_;
  assign new_n3213_ = new_n3202_ & ~new_n3212_;
  assign new_n3214_ = ~new_n3211_ & new_n3213_;
  assign new_n3215_ = new_n2139_ & ~new_n2177_;
  assign new_n3216_ = ~new_n2139_ & new_n2177_;
  assign new_n3217_ = ~new_n3215_ & ~new_n3216_;
  assign new_n3218_ = ~new_n3202_ & ~new_n3217_;
  assign \2_n22  = new_n3214_ | new_n3218_;
  assign new_n3220_ = ~new_n2032_ & ~new_n2038_;
  assign new_n3221_ = new_n2032_ & new_n2038_;
  assign new_n3222_ = ~new_n3220_ & ~new_n3221_;
  assign new_n3223_ = new_n2335_ & new_n3222_;
  assign new_n3224_ = ~new_n2335_ & ~new_n3222_;
  assign new_n3225_ = ~new_n3223_ & ~new_n3224_;
  assign new_n3226_ = ~new_n1876_ & ~new_n2045_;
  assign new_n3227_ = ~new_n2046_ & ~new_n3226_;
  assign new_n3228_ = ~new_n2049_ & ~new_n2052_;
  assign new_n3229_ = ~new_n2055_ & new_n3228_;
  assign new_n3230_ = new_n1875_ & ~new_n3229_;
  assign new_n3231_ = ~new_n1875_ & new_n3229_;
  assign new_n3232_ = ~new_n3230_ & ~new_n3231_;
  assign new_n3233_ = new_n3227_ & new_n3232_;
  assign new_n3234_ = ~new_n3227_ & ~new_n3232_;
  assign new_n3235_ = ~new_n3233_ & ~new_n3234_;
  assign new_n3236_ = ~new_n3225_ & new_n3235_;
  assign new_n3237_ = new_n3225_ & ~new_n3235_;
  assign new_n3238_ = ~new_n3236_ & ~new_n3237_;
  assign new_n3239_ = new_n1923_ & ~new_n3238_;
  assign new_n3240_ = new_n2340_ & new_n3222_;
  assign new_n3241_ = ~new_n2340_ & ~new_n3222_;
  assign new_n3242_ = ~new_n3240_ & ~new_n3241_;
  assign new_n3243_ = ~new_n2038_ & new_n2046_;
  assign new_n3244_ = new_n3229_ & ~new_n3243_;
  assign new_n3245_ = ~new_n3143_ & ~new_n3244_;
  assign new_n3246_ = new_n3143_ & new_n3244_;
  assign new_n3247_ = ~new_n3245_ & ~new_n3246_;
  assign new_n3248_ = new_n3227_ & new_n3247_;
  assign new_n3249_ = ~new_n3227_ & ~new_n3247_;
  assign new_n3250_ = ~new_n3248_ & ~new_n3249_;
  assign new_n3251_ = ~new_n3242_ & new_n3250_;
  assign new_n3252_ = new_n3242_ & ~new_n3250_;
  assign new_n3253_ = ~new_n3251_ & ~new_n3252_;
  assign new_n3254_ = ~new_n1923_ & new_n3253_;
  assign new_n3255_ = ~new_n3239_ & ~new_n3254_;
  assign new_n3256_ = ~\2_n545  & ~new_n3255_;
  assign new_n3257_ = ~new_n1909_ & new_n1923_;
  assign new_n3258_ = new_n3238_ & new_n3257_;
  assign new_n3259_ = \2_n545  & ~new_n3258_;
  assign new_n3260_ = ~new_n3253_ & ~new_n3257_;
  assign new_n3261_ = new_n3259_ & ~new_n3260_;
  assign new_n3262_ = ~new_n3256_ & ~new_n3261_;
  assign new_n3263_ = ~new_n1913_ & ~new_n1919_;
  assign new_n3264_ = ~new_n1882_ & new_n1888_;
  assign new_n3265_ = new_n1882_ & ~new_n1888_;
  assign new_n3266_ = ~new_n3264_ & ~new_n3265_;
  assign new_n3267_ = ~new_n3263_ & new_n3266_;
  assign new_n3268_ = new_n3263_ & ~new_n3266_;
  assign new_n3269_ = ~new_n3267_ & ~new_n3268_;
  assign new_n3270_ = new_n1898_ & new_n2073_;
  assign new_n3271_ = ~new_n1898_ & ~new_n2073_;
  assign new_n3272_ = ~new_n3270_ & ~new_n3271_;
  assign new_n3273_ = ~new_n3269_ & new_n3272_;
  assign new_n3274_ = new_n3269_ & ~new_n3272_;
  assign new_n3275_ = ~new_n3273_ & ~new_n3274_;
  assign new_n3276_ = new_n1895_ & ~new_n1906_;
  assign new_n3277_ = ~new_n1895_ & new_n1906_;
  assign new_n3278_ = ~new_n3276_ & ~new_n3277_;
  assign new_n3279_ = ~new_n1900_ & ~new_n3177_;
  assign new_n3280_ = new_n1900_ & new_n3177_;
  assign new_n3281_ = ~new_n3279_ & ~new_n3280_;
  assign new_n3282_ = new_n3278_ & new_n3281_;
  assign new_n3283_ = ~new_n3278_ & ~new_n3281_;
  assign new_n3284_ = ~new_n3282_ & ~new_n3283_;
  assign new_n3285_ = ~new_n3275_ & new_n3284_;
  assign new_n3286_ = new_n3275_ & ~new_n3284_;
  assign new_n3287_ = ~new_n3285_ & ~new_n3286_;
  assign new_n3288_ = ~\2_n545  & ~new_n3287_;
  assign new_n3289_ = ~new_n1900_ & new_n3266_;
  assign new_n3290_ = new_n1900_ & ~new_n3266_;
  assign new_n3291_ = ~new_n3289_ & ~new_n3290_;
  assign new_n3292_ = ~new_n3173_ & new_n3177_;
  assign new_n3293_ = ~new_n1907_ & new_n3263_;
  assign new_n3294_ = ~new_n3292_ & ~new_n3293_;
  assign new_n3295_ = new_n3292_ & new_n3293_;
  assign new_n3296_ = ~new_n3294_ & ~new_n3295_;
  assign new_n3297_ = ~new_n3291_ & new_n3296_;
  assign new_n3298_ = new_n3291_ & ~new_n3296_;
  assign new_n3299_ = ~new_n3297_ & ~new_n3298_;
  assign new_n3300_ = ~new_n1898_ & ~new_n1900_;
  assign new_n3301_ = ~new_n1908_ & new_n2073_;
  assign new_n3302_ = new_n3300_ & ~new_n3301_;
  assign new_n3303_ = ~new_n3300_ & new_n3301_;
  assign new_n3304_ = ~new_n3302_ & ~new_n3303_;
  assign new_n3305_ = ~new_n3299_ & new_n3304_;
  assign new_n3306_ = new_n3299_ & ~new_n3304_;
  assign new_n3307_ = ~new_n3305_ & ~new_n3306_;
  assign new_n3308_ = ~new_n3278_ & ~new_n3307_;
  assign new_n3309_ = new_n3278_ & new_n3307_;
  assign new_n3310_ = \2_n545  & ~new_n3309_;
  assign new_n3311_ = ~new_n3308_ & new_n3310_;
  assign new_n3312_ = ~new_n3288_ & ~new_n3311_;
  assign new_n3313_ = ~new_n3262_ & new_n3312_;
  assign new_n3314_ = new_n3262_ & ~new_n3312_;
  assign \2_n233  = ~new_n3313_ & ~new_n3314_;
  assign new_n3316_ = ~new_n2002_ & ~new_n2015_;
  assign new_n3317_ = ~new_n1987_ & new_n3316_;
  assign new_n3318_ = new_n2013_ & new_n2092_;
  assign new_n3319_ = new_n2001_ & new_n3318_;
  assign new_n3320_ = new_n3317_ & ~new_n3319_;
  assign new_n3321_ = new_n1993_ & ~new_n3320_;
  assign new_n3322_ = ~new_n1993_ & new_n3320_;
  assign \2_n247  = ~new_n3321_ & ~new_n3322_;
  assign \2_n30  = \2_n1050 ;
  assign \2_n304  = \2_n420  & \2_n832 ;
  assign new_n3326_ = new_n2134_ & new_n2144_;
  assign new_n3327_ = ~new_n2134_ & ~new_n2144_;
  assign new_n3328_ = ~new_n3326_ & ~new_n3327_;
  assign new_n3329_ = new_n3202_ & new_n3328_;
  assign new_n3330_ = ~new_n2144_ & ~new_n2171_;
  assign new_n3331_ = new_n2144_ & new_n2171_;
  assign new_n3332_ = ~new_n3202_ & ~new_n3331_;
  assign new_n3333_ = ~new_n3330_ & new_n3332_;
  assign \2_n364  = new_n3329_ | new_n3333_;
  assign new_n3335_ = ~new_n1992_ & ~new_n1994_;
  assign new_n3336_ = new_n1993_ & ~new_n3316_;
  assign new_n3337_ = new_n3335_ & ~new_n3336_;
  assign new_n3338_ = new_n1993_ & new_n2024_;
  assign new_n3339_ = ~new_n2080_ & new_n3338_;
  assign new_n3340_ = new_n3337_ & ~new_n3339_;
  assign new_n3341_ = ~new_n1983_ & new_n3340_;
  assign new_n3342_ = new_n1983_ & ~new_n3340_;
  assign \2_n370  = ~new_n3341_ & ~new_n3342_;
  assign new_n3344_ = ~new_n2270_ & new_n3158_;
  assign new_n3345_ = new_n2270_ & ~new_n3158_;
  assign new_n3346_ = ~new_n3344_ & ~new_n3345_;
  assign new_n3347_ = ~new_n2306_ & new_n3346_;
  assign new_n3348_ = ~new_n2263_ & ~new_n2270_;
  assign new_n3349_ = new_n2263_ & new_n2270_;
  assign new_n3350_ = ~new_n3348_ & ~new_n3349_;
  assign new_n3351_ = ~new_n2267_ & new_n3350_;
  assign new_n3352_ = new_n2267_ & ~new_n3350_;
  assign new_n3353_ = ~new_n3351_ & ~new_n3352_;
  assign new_n3354_ = new_n2306_ & new_n3353_;
  assign new_n3355_ = new_n2330_ & ~new_n3354_;
  assign new_n3356_ = ~new_n3347_ & new_n3355_;
  assign new_n3357_ = new_n2306_ & ~new_n2311_;
  assign new_n3358_ = ~new_n3353_ & new_n3357_;
  assign new_n3359_ = ~new_n3346_ & ~new_n3357_;
  assign new_n3360_ = ~new_n3358_ & ~new_n3359_;
  assign new_n3361_ = ~new_n2330_ & ~new_n3360_;
  assign new_n3362_ = ~new_n3356_ & ~new_n3361_;
  assign new_n3363_ = new_n2299_ & new_n3129_;
  assign new_n3364_ = ~new_n2299_ & ~new_n3129_;
  assign new_n3365_ = ~new_n3363_ & ~new_n3364_;
  assign new_n3366_ = ~new_n2279_ & new_n2283_;
  assign new_n3367_ = new_n2279_ & ~new_n2283_;
  assign new_n3368_ = ~new_n3366_ & ~new_n3367_;
  assign new_n3369_ = new_n3206_ & new_n3368_;
  assign new_n3370_ = ~new_n3206_ & ~new_n3368_;
  assign new_n3371_ = ~new_n3369_ & ~new_n3370_;
  assign new_n3372_ = new_n3365_ & new_n3371_;
  assign new_n3373_ = ~new_n3365_ & ~new_n3371_;
  assign new_n3374_ = ~new_n3372_ & ~new_n3373_;
  assign new_n3375_ = new_n2291_ & new_n2301_;
  assign new_n3376_ = ~new_n2291_ & ~new_n2301_;
  assign new_n3377_ = ~new_n3375_ & ~new_n3376_;
  assign new_n3378_ = new_n2283_ & new_n2303_;
  assign new_n3379_ = ~new_n2277_ & ~new_n2294_;
  assign new_n3380_ = ~new_n3378_ & new_n3379_;
  assign new_n3381_ = ~new_n2308_ & ~new_n3380_;
  assign new_n3382_ = new_n2308_ & new_n3380_;
  assign new_n3383_ = ~new_n3381_ & ~new_n3382_;
  assign new_n3384_ = new_n3377_ & new_n3383_;
  assign new_n3385_ = ~new_n3377_ & ~new_n3383_;
  assign new_n3386_ = ~new_n3384_ & ~new_n3385_;
  assign new_n3387_ = ~new_n3374_ & new_n3386_;
  assign new_n3388_ = new_n3374_ & ~new_n3386_;
  assign new_n3389_ = ~new_n3387_ & ~new_n3388_;
  assign new_n3390_ = new_n2330_ & ~new_n3389_;
  assign new_n3391_ = ~new_n2299_ & ~new_n2308_;
  assign new_n3392_ = ~new_n2310_ & new_n3129_;
  assign new_n3393_ = ~new_n3391_ & ~new_n3392_;
  assign new_n3394_ = new_n3391_ & new_n3392_;
  assign new_n3395_ = ~new_n3393_ & ~new_n3394_;
  assign new_n3396_ = ~new_n2308_ & new_n3368_;
  assign new_n3397_ = new_n2308_ & ~new_n3368_;
  assign new_n3398_ = ~new_n3396_ & ~new_n3397_;
  assign new_n3399_ = ~new_n2309_ & new_n3206_;
  assign new_n3400_ = new_n2283_ & new_n2310_;
  assign new_n3401_ = new_n3380_ & ~new_n3400_;
  assign new_n3402_ = new_n3399_ & new_n3401_;
  assign new_n3403_ = ~new_n3399_ & ~new_n3401_;
  assign new_n3404_ = ~new_n3402_ & ~new_n3403_;
  assign new_n3405_ = ~new_n3398_ & new_n3404_;
  assign new_n3406_ = new_n3398_ & ~new_n3404_;
  assign new_n3407_ = ~new_n3405_ & ~new_n3406_;
  assign new_n3408_ = ~new_n3395_ & new_n3407_;
  assign new_n3409_ = new_n3395_ & ~new_n3407_;
  assign new_n3410_ = ~new_n3408_ & ~new_n3409_;
  assign new_n3411_ = ~new_n3377_ & new_n3410_;
  assign new_n3412_ = new_n3377_ & ~new_n3410_;
  assign new_n3413_ = ~new_n2330_ & ~new_n3412_;
  assign new_n3414_ = ~new_n3411_ & new_n3413_;
  assign new_n3415_ = ~new_n3390_ & ~new_n3414_;
  assign new_n3416_ = new_n3362_ & ~new_n3415_;
  assign new_n3417_ = ~new_n3362_ & new_n3415_;
  assign \2_n378  = ~new_n3416_ & ~new_n3417_;
  assign new_n3419_ = ~new_n2130_ & ~new_n2132_;
  assign new_n3420_ = new_n3202_ & ~new_n3419_;
  assign new_n3421_ = ~new_n2133_ & new_n3420_;
  assign new_n3422_ = new_n2132_ & new_n2175_;
  assign new_n3423_ = ~new_n2132_ & ~new_n2175_;
  assign new_n3424_ = ~new_n3422_ & ~new_n3423_;
  assign new_n3425_ = ~new_n3202_ & ~new_n3424_;
  assign \2_n396  = new_n3421_ | new_n3425_;
  assign new_n3427_ = ~new_n1949_ & ~new_n1960_;
  assign new_n3428_ = ~new_n1969_ & new_n3427_;
  assign new_n3429_ = new_n1951_ & ~new_n3428_;
  assign new_n3430_ = ~new_n1951_ & new_n3428_;
  assign new_n3431_ = new_n2082_ & ~new_n3430_;
  assign new_n3432_ = ~new_n3429_ & new_n3431_;
  assign new_n3433_ = ~new_n1976_ & new_n3428_;
  assign new_n3434_ = ~new_n1951_ & ~new_n3433_;
  assign new_n3435_ = new_n1951_ & new_n3433_;
  assign new_n3436_ = ~new_n3434_ & ~new_n3435_;
  assign new_n3437_ = ~new_n2082_ & ~new_n3436_;
  assign \2_n517  = new_n3432_ | new_n3437_;
  assign new_n3439_ = new_n1935_ & new_n2064_;
  assign new_n3440_ = new_n2216_ & ~new_n3439_;
  assign new_n3441_ = ~new_n2113_ & new_n3440_;
  assign new_n3442_ = new_n2113_ & ~new_n3440_;
  assign \2_n534  = ~new_n3441_ & ~new_n3442_;
  assign new_n3444_ = new_n2271_ & new_n2311_;
  assign new_n3445_ = ~new_n2328_ & new_n3444_;
  assign new_n3446_ = new_n2264_ & ~new_n3445_;
  assign new_n3447_ = new_n2271_ & ~new_n2306_;
  assign new_n3448_ = new_n2317_ & new_n3444_;
  assign new_n3449_ = new_n2315_ & new_n3444_;
  assign new_n3450_ = ~new_n3448_ & ~new_n3449_;
  assign new_n3451_ = ~new_n3447_ & new_n3450_;
  assign \2_n553  = ~new_n3446_ | ~new_n3451_;
  assign new_n3453_ = ~\2_n545  & ~new_n1900_;
  assign \2_n597  = ~new_n2069_ & ~new_n3453_;
  assign new_n3455_ = ~new_n1951_ & new_n1959_;
  assign new_n3456_ = new_n1951_ & ~new_n1959_;
  assign new_n3457_ = ~new_n3455_ & ~new_n3456_;
  assign new_n3458_ = new_n3187_ & ~new_n3457_;
  assign new_n3459_ = ~new_n3187_ & new_n3457_;
  assign new_n3460_ = ~new_n3458_ & ~new_n3459_;
  assign new_n3461_ = ~new_n1967_ & ~new_n1974_;
  assign new_n3462_ = ~new_n1975_ & ~new_n3461_;
  assign new_n3463_ = ~new_n1965_ & new_n3428_;
  assign new_n3464_ = new_n1965_ & ~new_n3428_;
  assign new_n3465_ = ~new_n3463_ & ~new_n3464_;
  assign new_n3466_ = new_n3462_ & new_n3465_;
  assign new_n3467_ = ~new_n3462_ & ~new_n3465_;
  assign new_n3468_ = ~new_n3466_ & ~new_n3467_;
  assign new_n3469_ = ~new_n3460_ & new_n3468_;
  assign new_n3470_ = new_n3460_ & ~new_n3468_;
  assign new_n3471_ = ~new_n3469_ & ~new_n3470_;
  assign new_n3472_ = new_n2018_ & ~new_n3471_;
  assign new_n3473_ = new_n2080_ & ~new_n3472_;
  assign new_n3474_ = ~new_n2085_ & new_n3433_;
  assign new_n3475_ = new_n2085_ & ~new_n3433_;
  assign new_n3476_ = ~new_n3474_ & ~new_n3475_;
  assign new_n3477_ = new_n3462_ & new_n3476_;
  assign new_n3478_ = ~new_n3462_ & ~new_n3476_;
  assign new_n3479_ = ~new_n3477_ & ~new_n3478_;
  assign new_n3480_ = ~new_n3192_ & ~new_n3457_;
  assign new_n3481_ = new_n3192_ & new_n3457_;
  assign new_n3482_ = ~new_n3480_ & ~new_n3481_;
  assign new_n3483_ = ~new_n3479_ & new_n3482_;
  assign new_n3484_ = new_n3479_ & ~new_n3482_;
  assign new_n3485_ = ~new_n3483_ & ~new_n3484_;
  assign new_n3486_ = ~new_n2018_ & new_n3485_;
  assign new_n3487_ = new_n3473_ & ~new_n3486_;
  assign new_n3488_ = new_n2018_ & ~new_n2025_;
  assign new_n3489_ = new_n3471_ & new_n3488_;
  assign new_n3490_ = ~new_n3485_ & ~new_n3488_;
  assign new_n3491_ = ~new_n3489_ & ~new_n3490_;
  assign new_n3492_ = ~new_n2080_ & ~new_n3491_;
  assign new_n3493_ = ~new_n3487_ & ~new_n3492_;
  assign new_n3494_ = new_n2001_ & new_n2013_;
  assign new_n3495_ = ~new_n2001_ & ~new_n2013_;
  assign new_n3496_ = ~new_n3494_ & ~new_n3495_;
  assign new_n3497_ = ~new_n2022_ & ~new_n3337_;
  assign new_n3498_ = new_n2022_ & new_n3337_;
  assign new_n3499_ = ~new_n3497_ & ~new_n3498_;
  assign new_n3500_ = new_n3496_ & new_n3499_;
  assign new_n3501_ = ~new_n3496_ & ~new_n3499_;
  assign new_n3502_ = ~new_n3500_ & ~new_n3501_;
  assign new_n3503_ = new_n2011_ & new_n3317_;
  assign new_n3504_ = ~new_n2011_ & ~new_n3317_;
  assign new_n3505_ = ~new_n3503_ & ~new_n3504_;
  assign new_n3506_ = ~new_n1999_ & ~new_n2014_;
  assign new_n3507_ = ~new_n1983_ & ~new_n1993_;
  assign new_n3508_ = ~new_n2003_ & ~new_n3507_;
  assign new_n3509_ = new_n3506_ & new_n3508_;
  assign new_n3510_ = ~new_n3506_ & ~new_n3508_;
  assign new_n3511_ = ~new_n3509_ & ~new_n3510_;
  assign new_n3512_ = new_n3505_ & new_n3511_;
  assign new_n3513_ = ~new_n3505_ & ~new_n3511_;
  assign new_n3514_ = ~new_n3512_ & ~new_n3513_;
  assign new_n3515_ = ~new_n3502_ & new_n3514_;
  assign new_n3516_ = new_n3502_ & ~new_n3514_;
  assign new_n3517_ = ~new_n3515_ & ~new_n3516_;
  assign new_n3518_ = new_n2080_ & new_n3517_;
  assign new_n3519_ = ~new_n2011_ & ~new_n2022_;
  assign new_n3520_ = ~new_n2024_ & new_n3317_;
  assign new_n3521_ = ~new_n3519_ & ~new_n3520_;
  assign new_n3522_ = new_n3519_ & new_n3520_;
  assign new_n3523_ = ~new_n3521_ & ~new_n3522_;
  assign new_n3524_ = ~new_n2022_ & ~new_n3508_;
  assign new_n3525_ = new_n2022_ & new_n3508_;
  assign new_n3526_ = ~new_n3524_ & ~new_n3525_;
  assign new_n3527_ = ~new_n2023_ & new_n3506_;
  assign new_n3528_ = new_n3337_ & ~new_n3338_;
  assign new_n3529_ = new_n3527_ & new_n3528_;
  assign new_n3530_ = ~new_n3527_ & ~new_n3528_;
  assign new_n3531_ = ~new_n3529_ & ~new_n3530_;
  assign new_n3532_ = ~new_n3526_ & new_n3531_;
  assign new_n3533_ = new_n3526_ & ~new_n3531_;
  assign new_n3534_ = ~new_n3532_ & ~new_n3533_;
  assign new_n3535_ = ~new_n3523_ & new_n3534_;
  assign new_n3536_ = new_n3523_ & ~new_n3534_;
  assign new_n3537_ = ~new_n3535_ & ~new_n3536_;
  assign new_n3538_ = ~new_n3496_ & new_n3537_;
  assign new_n3539_ = new_n3496_ & ~new_n3537_;
  assign new_n3540_ = ~new_n2080_ & ~new_n3539_;
  assign new_n3541_ = ~new_n3538_ & new_n3540_;
  assign new_n3542_ = ~new_n3518_ & ~new_n3541_;
  assign new_n3543_ = new_n3493_ & ~new_n3542_;
  assign new_n3544_ = ~new_n3493_ & new_n3542_;
  assign \2_n625  = ~new_n3543_ & ~new_n3544_;
  assign new_n3546_ = \2_n1438  & \2_n1536 ;
  assign new_n3547_ = \2_n315  & \2_n997 ;
  assign \2_n669  = ~new_n3546_ | ~new_n3547_;
  assign new_n3549_ = ~new_n2011_ & ~new_n2092_;
  assign new_n3550_ = ~new_n2013_ & new_n3549_;
  assign new_n3551_ = new_n2013_ & ~new_n3549_;
  assign \2_n693  = ~new_n3550_ & ~
