module top( n0 , n21 , n29 , n34 , n36 , n38 , n45 , n49 , n60 , n77 , n81 , n82 , n88 , n90 , n91 , n95 , n98 , n104 , n107 , n108 , n112 , n116 , n122 , n127 , n128 , n129 , n130 , n135 , n138 , n150 , n153 , n159 , n167 , n168 , n175 , n185 , n190 , n192 , n193 , n196 , n200 , n204 , n206 , n207 , n208 , n218 , n221 , n223 , n227 , n228 , n229 , n231 , n236 , n240 , n244 , n245 , n246 , n252 , n258 , n260 , n262 , n267 , n268 , n275 , n281 , n284 , n288 , n299 , n301 , n305 , n307 , n310 , n319 , n323 , n324 , n332 , n336 , n342 , n347 , n359 , n360 , n364 , n366 , n374 , n381 , n383 , n384 , n389 , n393 , n398 , n408 , n409 , n410 , n415 , n421 , n423 , n431 , n432 , n433 , n438 , n439 , n441 , n444 , n448 , n449 , n452 , n456 , n475 , n491 , n492 , n500 , n505 , n507 , n510 , n516 , n519 , n532 , n536 , n540 , n554 , n571 , n577 , n580 , n589 , n592 , n598 , n599 , n607 , n608 , n610 , n613 , n617 , n621 , n623 , n627 , n631 , n635 , n638 , n640 , n644 , n650 , n651 , n653 , n657 , n662 , n667 , n679 , n683 , n685 , n688 , n695 , n707 , n710 , n714 , n716 , n718 , n723 , n733 , n734 , n741 , n745 , n747 , n749 , n766 , n767 , n771 , n774 , n779 , n785 , n787 , n801 , n802 , n804 , n806 , n807 , n808 , n817 , n818 , n819 , n823 , n825 , n826 , n833 , n835 , n839 , n841 , n842 , n845 , n851 , n853 , n854 , n857 , n862 , n863 , n866 , n870 , n877 , n879 , n893 , n896 , n901 , n905 , n908 , n927 , n928 , n929 , n936 , n944 , n952 , n955 , n961 , n962 , n966 , n973 , n975 , n976 , n986 , n997 , n999 , n1005 , n1022 , n1023 , n1027 , n1029 , n1035 , n1036 , n1041 , n1044 , n1045 , n1048 , n1057 , n1059 , n1061 , n1064 , n1067 , n1069 , n1072 , n1073 , n1077 , n1080 , n1081 , n1085 , n1089 , n1091 , n1097 , n1098 , n1099 , n1120 , n1131 , n1132 , n1140 , n1141 , n1143 , n1146 , n1150 , n1151 , n1153 , n1163 , n1164 , n1178 , n1180 , n1184 , n1191 , n1194 , n1198 , n1202 , n1206 , n1219 , n1226 , n1229 , n1231 , n1232 , n1236 , n1239 , n1257 , n1259 , n1264 , n1269 , n1273 , n1277 , n1279 , n1288 , n1298 , n1301 , n1308 , n1311 , n1321 , n1326 , n1342 , n1344 , n1352 );
    input n0 , n21 , n36 , n38 , n45 , n49 , n77 , n95 , n98 , n104 , n107 , n108 , n116 , n122 , n127 , n128 , n138 , n153 , n192 , n196 , n200 , n208 , n221 , n231 , n236 , n244 , n245 , n246 , n252 , n258 , n260 , n262 , n267 , n268 , n281 , n284 , n288 , n301 , n305 , n310 , n319 , n323 , n324 , n332 , n336 , n359 , n360 , n364 , n366 , n381 , n384 , n393 , n398 , n421 , n423 , n431 , n433 , n438 , n439 , n441 , n444 , n448 , n449 , n475 , n491 , n500 , n505 , n507 , n510 , n519 , n532 , n536 , n540 , n571 , n577 , n589 , n599 , n610 , n631 , n635 , n640 , n644 , n650 , n657 , n667 , n685 , n688 , n695 , n714 , n716 , n741 , n745 , n749 , n766 , n767 , n771 , n774 , n787 , n802 , n804 , n806 , n818 , n819 , n823 , n825 , n826 , n833 , n839 , n841 , n845 , n851 , n857 , n862 , n863 , n866 , n870 , n879 , n893 , n896 , n901 , n928 , n929 , n936 , n944 , n952 , n955 , n961 , n975 , n976 , n986 , n997 , n1005 , n1022 , n1029 , n1035 , n1036 , n1041 , n1044 , n1045 , n1048 , n1064 , n1067 , n1069 , n1072 , n1073 , n1077 , n1080 , n1081 , n1089 , n1091 , n1097 , n1098 , n1120 , n1131 , n1132 , n1140 , n1141 , n1143 , n1146 , n1151 , n1163 , n1164 , n1180 , n1191 , n1198 , n1219 , n1226 , n1229 , n1231 , n1236 , n1257 , n1269 , n1273 , n1277 , n1279 , n1298 , n1308 , n1311 , n1321 , n1326 , n1342 , n1344 , n1352 ;
    output n29 , n34 , n60 , n81 , n82 , n88 , n90 , n91 , n112 , n129 , n130 , n135 , n150 , n159 , n167 , n168 , n175 , n185 , n190 , n193 , n204 , n206 , n207 , n218 , n223 , n227 , n228 , n229 , n240 , n275 , n299 , n307 , n342 , n347 , n374 , n383 , n389 , n408 , n409 , n410 , n415 , n432 , n452 , n456 , n492 , n516 , n554 , n580 , n592 , n598 , n607 , n608 , n613 , n617 , n621 , n623 , n627 , n638 , n651 , n653 , n662 , n679 , n683 , n707 , n710 , n718 , n723 , n733 , n734 , n747 , n779 , n785 , n801 , n807 , n808 , n817 , n835 , n842 , n853 , n854 , n877 , n905 , n908 , n927 , n962 , n966 , n973 , n999 , n1023 , n1027 , n1057 , n1059 , n1061 , n1085 , n1099 , n1150 , n1153 , n1178 , n1184 , n1194 , n1202 , n1206 , n1232 , n1239 , n1259 , n1264 , n1288 , n1301 ;
    wire n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n30 , n31 , n32 , n33 , n35 , n37 , n39 , n40 , n41 , n42 , n43 , n44 , n46 , n47 , n48 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n78 , n79 , n80 , n83 , n84 , n85 , n86 , n87 , n89 , n92 , n93 , n94 , n96 , n97 , n99 , n100 , n101 , n102 , n103 , n105 , n106 , n109 , n110 , n111 , n113 , n114 , n115 , n117 , n118 , n119 , n120 , n121 , n123 , n124 , n125 , n126 , n131 , n132 , n133 , n134 , n136 , n137 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n151 , n152 , n154 , n155 , n156 , n157 , n158 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n169 , n170 , n171 , n172 , n173 , n174 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n186 , n187 , n188 , n189 , n191 , n194 , n195 , n197 , n198 , n199 , n201 , n202 , n203 , n205 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n219 , n220 , n222 , n224 , n225 , n226 , n230 , n232 , n233 , n234 , n235 , n237 , n238 , n239 , n241 , n242 , n243 , n247 , n248 , n249 , n250 , n251 , n253 , n254 , n255 , n256 , n257 , n259 , n261 , n263 , n264 , n265 , n266 , n269 , n270 , n271 , n272 , n273 , n274 , n276 , n277 , n278 , n279 , n280 , n282 , n283 , n285 , n286 , n287 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n300 , n302 , n303 , n304 , n306 , n308 , n309 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n320 , n321 , n322 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n333 , n334 , n335 , n337 , n338 , n339 , n340 , n341 , n343 , n344 , n345 , n346 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n361 , n362 , n363 , n365 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n375 , n376 , n377 , n378 , n379 , n380 , n382 , n385 , n386 , n387 , n388 , n390 , n391 , n392 , n394 , n395 , n396 , n397 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n411 , n412 , n413 , n414 , n416 , n417 , n418 , n419 , n420 , n422 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n434 , n435 , n436 , n437 , n440 , n442 , n443 , n445 , n446 , n447 , n450 , n451 , n453 , n454 , n455 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n501 , n502 , n503 , n504 , n506 , n508 , n509 , n511 , n512 , n513 , n514 , n515 , n517 , n518 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n533 , n534 , n535 , n537 , n538 , n539 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n572 , n573 , n574 , n575 , n576 , n578 , n579 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n590 , n591 , n593 , n594 , n595 , n596 , n597 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n609 , n611 , n612 , n614 , n615 , n616 , n618 , n619 , n620 , n622 , n624 , n625 , n626 , n628 , n629 , n630 , n632 , n633 , n634 , n636 , n637 , n639 , n641 , n642 , n643 , n645 , n646 , n647 , n648 , n649 , n652 , n654 , n655 , n656 , n658 , n659 , n660 , n661 , n663 , n664 , n665 , n666 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n680 , n681 , n682 , n684 , n686 , n687 , n689 , n690 , n691 , n692 , n693 , n694 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n708 , n709 , n711 , n712 , n713 , n715 , n717 , n719 , n720 , n721 , n722 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n735 , n736 , n737 , n738 , n739 , n740 , n742 , n743 , n744 , n746 , n748 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n768 , n769 , n770 , n772 , n773 , n775 , n776 , n777 , n778 , n780 , n781 , n782 , n783 , n784 , n786 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n803 , n805 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n820 , n821 , n822 , n824 , n827 , n828 , n829 , n830 , n831 , n832 , n834 , n836 , n837 , n838 , n840 , n843 , n844 , n846 , n847 , n848 , n849 , n850 , n852 , n855 , n856 , n858 , n859 , n860 , n861 , n864 , n865 , n867 , n868 , n869 , n871 , n872 , n873 , n874 , n875 , n876 , n878 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n894 , n895 , n897 , n898 , n899 , n900 , n902 , n903 , n904 , n906 , n907 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n930 , n931 , n932 , n933 , n934 , n935 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n953 , n954 , n956 , n957 , n958 , n959 , n960 , n963 , n964 , n965 , n967 , n968 , n969 , n970 , n971 , n972 , n974 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n998 , n1000 , n1001 , n1002 , n1003 , n1004 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1024 , n1025 , n1026 , n1028 , n1030 , n1031 , n1032 , n1033 , n1034 , n1037 , n1038 , n1039 , n1040 , n1042 , n1043 , n1046 , n1047 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1058 , n1060 , n1062 , n1063 , n1065 , n1066 , n1068 , n1070 , n1071 , n1074 , n1075 , n1076 , n1078 , n1079 , n1082 , n1083 , n1084 , n1086 , n1087 , n1088 , n1090 , n1092 , n1093 , n1094 , n1095 , n1096 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1142 , n1144 , n1145 , n1147 , n1148 , n1149 , n1152 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1179 , n1181 , n1182 , n1183 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1192 , n1193 , n1195 , n1196 , n1197 , n1199 , n1200 , n1201 , n1203 , n1204 , n1205 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1227 , n1228 , n1230 , n1233 , n1234 , n1235 , n1237 , n1238 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1258 , n1260 , n1261 , n1262 , n1263 , n1265 , n1266 , n1267 , n1268 , n1270 , n1271 , n1272 , n1274 , n1275 , n1276 , n1278 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1299 , n1300 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1309 , n1310 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1322 , n1323 , n1324 , n1325 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1343 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1353 ;
assign n55 = n1004 | n1113;
assign n1107 = n1214 | n636;
assign n487 = ~n942;
assign n682 = n1332 & n147;
assign n1004 = n1158 ^ n974;
assign n744 = ~(n89 ^ n393);
assign n502 = ~n375;
assign n471 = ~(n643 | n52);
assign n1240 = ~(n152 ^ n499);
assign n1303 = n846 & n153;
assign n1168 = ~(n78 ^ n1156);
assign n894 = n449 | n497;
assign n472 = ~(n838 | n727);
assign n638 = n1311;
assign n313 = ~n634;
assign n216 = n579 | n1320;
assign n854 = n243 & n647;
assign n1052 = ~n505;
assign n584 = n525 & n1324;
assign n721 = ~(n920 ^ n501);
assign n356 = n1093 | n435;
assign n683 = n381;
assign n756 = ~n514;
assign n217 = ~n951;
assign n827 = ~(n440 | n522);
assign n42 = ~(n301 | n1312);
assign n652 = n1198 | n403;
assign n1100 = ~(n1224 | n317);
assign n563 = n987 & n269;
assign n1253 = ~(n1225 | n697);
assign n996 = n205 | n541;
assign n732 = n985 & n528;
assign n1109 = n1076 & n687;
assign n478 = ~(n703 | n189);
assign n509 = n1300 | n981;
assign n840 = n692 & n238;
assign n60 = n1081;
assign n184 = n1216 | n1275;
assign n254 = ~(n955 ^ n851);
assign n932 = n456 & n574;
assign n1315 = ~(n571 | n1047);
assign n836 = ~n796;
assign n490 = ~n631;
assign n1245 = ~(n1081 | n1205);
assign n1082 = n496 | n670;
assign n1332 = n1038 ^ n1311;
assign n227 = 1'b0;
assign n469 = ~n601;
assign n220 = ~n1091;
assign n415 = n997;
assign n964 = ~(n805 | n550);
assign n1150 = ~(n1015 ^ n1350);
assign n765 = ~(n1130 ^ n957);
assign n27 = ~n239;
assign n956 = ~(n1290 ^ n889);
assign n671 = n1236 & n319;
assign n871 = ~n656;
assign n941 = n1213 ^ n1081;
assign n1290 = ~(n254 | n815);
assign n377 = n1198 | n520;
assign n719 = ~(n1126 | n1313);
assign n1139 = n36 | n1317;
assign n459 = n1273 & n688;
assign n1006 = ~(n472 ^ n765);
assign n152 = n502 & n591;
assign n51 = ~n52;
assign n690 = n1351 | n214;
assign n161 = n941 | n416;
assign n969 = ~(n188 ^ n1095);
assign n279 = n871 & n1345;
assign n1280 = ~n330;
assign n443 = ~n177;
assign n1086 = n53 | n602;
assign n1026 = n584 | n1248;
assign n29 = n1259;
assign n733 = ~(n1108 ^ n744);
assign n211 = ~(n777 | n1313);
assign n698 = n471 & n995;
assign n382 = n1116 & n1307;
assign n653 = n717 & n939;
assign n890 = ~(n524 | n261);
assign n145 = n332 | n970;
assign n1250 = ~n688;
assign n614 = n1062 & n831;
assign n429 = ~(n1123 ^ n535);
assign n183 = n1222 ^ n47;
assign n927 = n824 & n1027;
assign n80 = n688 | n759;
assign n552 = n371 | n405;
assign n229 = n785;
assign n1104 = ~n3;
assign n991 = ~(n1349 ^ n138);
assign n1042 = ~n630;
assign n253 = n485 & n264;
assign n1057 = n332;
assign n177 = ~n257;
assign n1106 = ~(n821 ^ n440);
assign n568 = n716 | n891;
assign n762 = ~(n885 | n143);
assign n1203 = n40 | n660;
assign n125 = n663 | n1049;
assign n461 = n272 | n583;
assign n753 = n403 & n695;
assign n1142 = ~(n508 ^ n1034);
assign n895 = n219 | n1157;
assign n701 = ~n585;
assign n861 = n269 & n446;
assign n998 = ~(n1011 ^ n641);
assign n659 = ~(n1248 ^ n20);
assign n1058 = n198 & n131;
assign n24 = ~(n799 ^ n1200);
assign n1049 = n680;
assign n792 = ~(n559 | n457);
assign n249 = ~(n775 ^ n259);
assign n62 = n1337 & n9;
assign n570 = ~(n292 ^ n1142);
assign n830 = ~(n757 | n813);
assign n118 = ~n418;
assign n704 = ~(n1262 ^ n1211);
assign n1338 = n1020 | n1299;
assign n66 = n438 ^ n1048;
assign n1305 = n1098 & n688;
assign n643 = n1109 & n474;
assign n1285 = n688 | n100;
assign n1216 = n947 & n928;
assign n1007 = ~n991;
assign n1254 = n1018 & n585;
assign n198 = n688 | n1092;
assign n696 = n811 | n16;
assign n1155 = n350 | n743;
assign n921 = ~(n1321 | n1205);
assign n75 = n1316 & n958;
assign n731 = n1050 & n1056;
assign n357 = n1049 & n863;
assign n117 = ~n1332;
assign n847 = ~(n604 ^ n1238);
assign n700 = ~(n341 ^ n396);
assign n210 = ~n297;
assign n1255 = ~(n296 ^ n96);
assign n348 = ~(n1189 ^ n1030);
assign n1260 = ~(n1186 | n725);
assign n176 = ~n208;
assign n1137 = ~(n909 | n75);
assign n224 = n846 & n1164;
assign n865 = ~(n1323 ^ n270);
assign n634 = ~(n1190 ^ n36);
assign n492 = 1'b0;
assign n286 = ~(n25 ^ n1340);
assign n561 = n427 | n968;
assign n978 = ~(n1319 | n1192);
assign n971 = n1171 & n1207;
assign n590 = ~(n788 | n14);
assign n1293 = ~(n1349 ^ n1213);
assign n770 = ~n330;
assign n626 = n1271 | n798;
assign n1186 = ~(n609 ^ n573);
assign n764 = ~(n1123 | n457);
assign n121 = ~n1326;
assign n628 = n814 & n281;
assign n680 = ~n688;
assign n1208 = n1171 & n552;
assign n602 = n1205 & n1269;
assign n306 = ~(n247 ^ n948);
assign n946 = n1315 | n387;
assign n1178 = ~(n634 ^ n840);
assign n9 = n690 & n28;
assign n1112 = ~(n900 | n392);
assign n1284 = ~n1325;
assign n593 = n688 | n19;
assign n1084 = n706 | n357;
assign n609 = ~(n466 ^ n1117);
assign n195 = n1049 & n818;
assign n973 = n819;
assign n565 = ~(n982 | n195);
assign n178 = ~n310;
assign n604 = ~n586;
assign n776 = ~n796;
assign n1015 = ~(n792 | n912);
assign n206 = n732 | n118;
assign n1018 = ~n47;
assign n19 = ~n245;
assign n815 = ~n1330;
assign n670 = n1254 & n1222;
assign n167 = ~(n1280 ^ n394);
assign n1259 = n691 | n1183;
assign n1145 = n31 | n646;
assign n684 = ~n528;
assign n518 = n766 & n635;
assign n608 = 1'b0;
assign n307 = n1308;
assign n158 = ~n1069;
assign n1258 = ~(n953 ^ n1155);
assign n1094 = ~n744;
assign n529 = n688 | n1212;
assign n703 = ~(n241 | n907);
assign n1317 = ~n1190;
assign n967 = n1270 | n253;
assign n859 = n688 | n1229;
assign n344 = ~n75;
assign n1016 = ~(n974 ^ n659);
assign n951 = n178 | n403;
assign n1287 = n1176 & n975;
assign n465 = n772 | n693;
assign n648 = n888 | n614;
assign n112 = n116 & n1257;
assign n1021 = ~n1313;
assign n881 = ~n1058;
assign n988 = n1282 | n742;
assign n736 = ~(n291 ^ n79);
assign n915 = ~(n770 ^ n261);
assign n385 = n118 & n1147;
assign n910 = ~n75;
assign n715 = n417 & n139;
assign n511 = ~(n566 ^ n589);
assign n523 = ~(n443 ^ n231);
assign n460 = n45 | n846;
assign n506 = ~(n153 | n688);
assign n738 = n661 | n812;
assign n1012 = ~n965;
assign n812 = ~(n997 | n1049);
assign n1159 = ~(n1094 | n367);
assign n1099 = n1325 ^ n515;
assign n168 = n597 & n453;
assign n397 = n52 & n1332;
assign n32 = n419 | n1166;
assign n583 = ~n214;
assign n30 = n1246 | n295;
assign n1087 = n688 & n1163;
assign n64 = ~n1073;
assign n383 = n1321;
assign n783 = ~(n1055 ^ n216);
assign n282 = n293 & n1139;
assign n450 = n447 | n636;
assign n878 = n300 & n1207;
assign n22 = n1140 & n688;
assign n191 = ~n0;
assign n1172 = n846 & n233;
assign n1271 = ~n1249;
assign n189 = n139 | n979;
assign n706 = ~n125;
assign n109 = n217 | n102;
assign n256 = n421 | n1205;
assign n520 = ~n354;
assign n1302 = ~(n458 ^ n820);
assign n404 = n403 & n221;
assign n566 = ~n165;
assign n201 = n618 | n977;
assign n180 = ~(n576 ^ n461);
assign n661 = n846 & n774;
assign n1050 = n945 | n464;
assign n654 = ~(n84 ^ n564);
assign n613 = n592;
assign n1301 = n71 ^ n133;
assign n513 = n846 & n267;
assign n185 = n571;
assign n788 = ~n393;
assign n624 = ~n1110;
assign n902 = ~(n1011 | n1079);
assign n615 = n17 | n935;
assign n334 = n850 | n1275;
assign n123 = n436 | n187;
assign n1068 = ~(n757 | n1278);
assign n501 = n65 | n911;
assign n737 = n901 & n688;
assign n361 = n1136 | n789;
assign n585 = n965 & n7;
assign n1312 = ~n895;
assign n203 = ~(n455 | n3);
assign n1328 = ~n833;
assign n557 = n109 ^ n332;
assign n480 = n1347 | n182;
assign n413 = ~(n923 ^ n763);
assign n687 = ~(n56 ^ n571);
assign n50 = ~(n738 | n44);
assign n464 = n550 & n1101;
assign n126 = ~n67;
assign n1292 = n688 | n220;
assign n219 = n1045 & n688;
assign n1165 = n521 | n878;
assign n691 = n1002 | n1032;
assign n147 = n1311 | n83;
assign n270 = ~(n174 ^ n678);
assign n1274 = ~(n995 ^ n31);
assign n1218 = ~(n41 ^ n735);
assign n63 = ~(n1019 | n696);
assign n170 = ~(n938 ^ n1293);
assign n67 = ~n1031;
assign n1060 = ~(n1022 | n839);
assign n129 = ~(n378 ^ n352);
assign n209 = ~n1084;
assign n549 = ~n761;
assign n498 = ~n117;
assign n1333 = ~n731;
assign n402 = n274 | n1245;
assign n131 = n191 | n1049;
assign n238 = ~n600;
assign n297 = n688 | n1179;
assign n897 = ~(n1035 | n846);
assign n347 = n1342;
assign n805 = ~n1201;
assign n595 = ~(n1310 ^ n1152);
assign n272 = ~n212;
assign n406 = ~(n138 | n1049);
assign n371 = n1205 & n423;
assign n171 = n271 | n921;
assign n855 = ~(n682 | n764);
assign n1116 = ~(n57 | n772);
assign n1000 = n1286 | n1275;
assign n1296 = n1051 & n1205;
assign n427 = ~n532;
assign n1028 = n571 | n403;
assign n1322 = n173 | n76;
assign n632 = n688 | n278;
assign n495 = ~n1270;
assign n100 = ~n893;
assign n1222 = n708 & n70;
assign n748 = ~(n1004 | n1026);
assign n130 = n716;
assign n239 = ~n731;
assign n1353 = n431 & n688;
assign n391 = ~(n114 ^ n860);
assign n533 = n263 & n339;
assign n37 = ~n445;
assign n809 = n1108 & n1159;
assign n587 = ~n1270;
assign n686 = n786 | n340;
assign n1329 = ~n1330;
assign n139 = n837 & n1055;
assign n554 = n360;
assign n1154 = ~(n433 | n403);
assign n816 = ~(n589 | n165);
assign n586 = n125 & n1285;
assign n1133 = n553 ^ n1335;
assign n1061 = ~(n712 ^ n1145);
assign n1010 = ~(n890 | n382);
assign n1243 = ~(n517 ^ n1261);
assign n999 = n484 & n518;
assign n477 = ~(n39 ^ n1274);
assign n82 = n104;
assign n87 = n1105 | n276;
assign n417 = n729 | n110;
assign n993 = n364 & n688;
assign n938 = n232 | n404;
assign n1 = ~(n467 | n315);
assign n666 = ~n686;
assign n115 = n1322 | n395;
assign n837 = n222 | n588;
assign n1030 = ~(n1158 ^ n1065);
assign n1055 = n539 | n512;
assign n1235 = ~(n575 ^ n1122);
assign n909 = ~(n180 ^ n1240);
assign n1252 = ~n849;
assign n26 = ~(n152 | n1054);
assign n1090 = ~(n876 ^ n420);
assign n673 = ~n694;
assign n205 = ~n645;
assign n810 = n610 & n688;
assign n1126 = ~(n622 ^ n298);
assign n390 = ~n317;
assign n775 = ~(n37 ^ n287);
assign n25 = n746 | n210;
assign n134 = n213 & n1294;
assign n1281 = ~(n601 ^ n881);
assign n1105 = n1204 & n501;
assign n488 = n454 | n282;
assign n900 = n1172 & n1020;
assign n1083 = n45 | n829;
assign n1276 = n836 & n749;
assign n47 = n358 | n285;
assign n90 = ~(n442 ^ n375);
assign n889 = ~(n343 ^ n639);
assign n422 = ~(n439 | n1329);
assign n1350 = n1187 | n1137;
assign n1319 = ~(n1134 ^ n637);
assign n149 = ~(n895 ^ n793);
assign n1175 = n988 & n953;
assign n326 = ~n71;
assign n280 = n1311 | n846;
assign n1211 = ~(n294 ^ n904);
assign n70 = n567 | n796;
assign n1066 = n800 | n403;
assign n761 = ~n313;
assign n790 = ~n95;
assign n1283 = n280 & n632;
assign n755 = n1228 | n6;
assign n556 = n336 & n384;
assign n17 = ~(n339 | n263);
assign n462 = ~n612;
assign n1334 = ~(n37 | n141);
assign n1223 = n583 ^ n576;
assign n697 = ~(n212 | n345);
assign n1088 = n688 & n252;
assign n954 = n124 & n168;
assign n317 = n1195 | n437;
assign n234 = n944 | n596;
assign n907 = n867 | n762;
assign n752 = n444 & n688;
assign n187 = ~n1242;
assign n213 = ~n304;
assign n821 = n993 | n404;
assign n309 = ~n685;
assign n7 = n1052 | n796;
assign n822 = ~n944;
assign n940 = ~n268;
assign n656 = ~n946;
assign n15 = ~(n136 | n1071);
assign n779 = n494 | n33;
assign n18 = ~n511;
assign n832 = ~n416;
assign n1185 = ~n482;
assign n980 = ~(n1109 | n946);
assign n784 = ~n761;
assign n906 = ~(n376 ^ n120);
assign n481 = ~n1158;
assign n1201 = n1205 & n328;
assign n645 = n22 | n1268;
assign n1286 = n776 & n217;
assign n1074 = n403 & n741;
assign n674 = n289 | n30;
assign n367 = n1166 | n144;
assign n1056 = n997 | n209;
assign n54 = n58 | n414;
assign n709 = ~(n589 | n846);
assign n926 = n688 | n616;
assign n1196 = n688 | n176;
assign n257 = ~n1000;
assign n1247 = n587 ^ n1040;
assign n1336 = ~n196;
assign n965 = ~n1148;
assign n850 = n814 & n507;
assign n639 = n1330 & n66;
assign n750 = n132 | n514;
assign n232 = n1191 & n688;
assign n199 = n557 | n473;
assign n350 = n403 & n540;
assign n672 = ~(n682 ^ n980);
assign n186 = n688 | n1336;
assign n785 = n385 | n99;
assign n1267 = ~n620;
assign n658 = ~(n291 ^ n619);
assign n970 = ~n109;
assign n1031 = ~n724;
assign n1129 = n701 | n711;
assign n1187 = n1121 & n2;
assign n76 = n873 | n478;
assign n207 = n1198;
assign n913 = ~n3;
assign n1349 = ~n412;
assign n295 = n542 | n1181;
assign n580 = n449;
assign n739 = n476 & n996;
assign n1059 = ~(n553 ^ n302);
assign n223 = 1'b0;
assign n607 = ~(n1039 ^ n1253);
assign n375 = ~(n601 ^ n104);
assign n553 = ~n875;
assign n1054 = n1121 & n591;
assign n503 = ~n510;
assign n303 = ~(n626 ^ n780);
assign n1266 = n234 | n751;
assign n89 = ~n527;
assign n525 = n688 | n1125;
assign n91 = n1259;
assign n948 = ~(n1144 ^ n998);
assign n1209 = ~(n475 | n846);
assign n271 = n1205 & n1279;
assign n942 = n356 ^ n1321;
assign n1130 = ~n313;
assign n846 = n680;
assign n853 = n589;
assign n84 = ~(n688 | n726);
assign n56 = n963 | n843;
assign n780 = ~(n1124 ^ n794);
assign n793 = ~(n356 ^ n105);
assign n1037 = ~n562;
assign n315 = ~n157;
assign n485 = n514 | n894;
assign n1239 = ~(n1043 ^ n855);
assign n120 = ~(n831 ^ n339);
assign n803 = ~(n1118 ^ n837);
assign n136 = n1017 | n11;
assign n197 = ~n451;
assign n1121 = ~n344;
assign n1202 = ~(n511 ^ n62);
assign n179 = ~n480;
assign n538 = n1129 & n47;
assign n1108 = ~n913;
assign n1246 = n1001 & n920;
assign n53 = ~(n381 | n846);
assign n947 = ~n796;
assign n340 = n1185 | n582;
assign n372 = ~(n720 ^ n321);
assign n572 = n629 & n501;
assign n798 = ~n630;
assign n799 = ~(n79 ^ n426);
assign n174 = n166 | n1303;
assign n175 = n138;
assign n773 = n1205 & n77;
assign n354 = n119 | n430;
assign n97 = n655 ^ n915;
assign n515 = n1267 & n670;
assign n867 = n369 & n1167;
assign n582 = n142 & n1094;
assign n1002 = ~(n1233 | n250);
assign n578 = n1008 | n13;
assign n437 = ~n322;
assign n751 = n454 | n784;
assign n882 = ~(n72 ^ n795);
assign n106 = ~n1333;
assign n418 = ~n730;
assign n1278 = n611 | n164;
assign n1085 = ~(n694 ^ n464);
assign n689 = n142 & n1114;
assign n374 = 1'b0;
assign n786 = n581 | n285;
assign n534 = ~n720;
assign n1189 = n1167 ^ n1309;
assign n376 = n43 | n984;
assign n3 = n917 | n887;
assign n1212 = ~n1077;
assign n442 = ~n910;
assign n600 = ~n234;
assign n717 = ~(n308 | n54);
assign n1340 = n983 | n753;
assign n1169 = n881 ^ n360;
assign n222 = n846 & n441;
assign n304 = ~n834;
assign n497 = ~n361;
assign n71 = ~(n462 ^ n38);
assign n33 = ~n711;
assign n226 = n1081 | n73;
assign n265 = ~n365;
assign n923 = ~(n391 ^ n722);
assign n241 = n101 & n171;
assign n290 = ~n796;
assign n1162 = ~(n946 ^ n429);
assign n992 = n644 | n1205;
assign n172 = n544 & n1217;
assign n758 = ~(n1100 | n79);
assign n1033 = ~n796;
assign n486 = n1205 & n857;
assign n1310 = ~n326;
assign n289 = ~(n94 ^ n1155);
assign n1153 = n231;
assign n1251 = ~n557;
assign n1177 = n1087 | n316;
assign n454 = ~n71;
assign n1020 = n1205 & n790;
assign n1264 = n116;
assign n702 = ~(n265 ^ n1010);
assign n655 = ~n1014;
assign n1265 = ~(n360 | n1049);
assign n746 = n745 & n688;
assign n1197 = n943 | n1205;
assign n52 = n42 | n279;
assign n165 = n322 & n728;
assign n1316 = n942 | n1348;
assign n740 = n1078 | n630;
assign n58 = ~(n407 ^ n700);
assign n248 = n1263 & n1309;
assign n934 = n950 | n897;
assign n242 = ~(n303 | n731);
assign n1123 = ~n147;
assign n341 = n1136 | n753;
assign n188 = ~n255;
assign n829 = ~n938;
assign n1327 = n1097 & n688;
assign n924 = n315 & n1109;
assign n983 = n1044 & n688;
assign n85 = n408 & n817;
assign n591 = n104 | n469;
assign n849 = ~n1169;
assign n218 = n545 | n538;
assign n368 = ~n67;
assign n1345 = ~(n895 ^ n301);
assign n163 = ~(n268 | n403);
assign n235 = ~(n1209 | n160);
assign n1192 = n24 | n1295;
assign n1092 = ~n1132;
assign n111 = n151 ^ n1248;
assign n445 = n1025 | n1275;
assign n6 = n830 & n333;
assign n1125 = ~n323;
assign n164 = ~n1155;
assign n151 = ~n584;
assign n318 = ~(n1147 | n349);
assign n575 = ~(n504 ^ n672);
assign n1188 = n1351 | n212;
assign n842 = n1184;
assign n243 = n448 & n870;
assign n74 = ~n1079;
assign n333 = n338 | n1256;
assign n483 = n754 ^ n991;
assign n337 = ~(n919 | n590);
assign n269 = n740 & n1083;
assign n1103 = ~(n154 ^ n834);
assign n824 = n954 & n854;
assign n1119 = n1110 & n1307;
assign n4 = n827 & n821;
assign n576 = ~(n1039 ^ n511);
assign n1233 = ~n1352;
assign n642 = ~n340;
assign n1330 = n708 & n947;
assign n325 = ~(n380 ^ n400);
assign n5 = ~(n1019 ^ n304);
assign n388 = ~(n132 | n509);
assign n931 = ~(n777 ^ n194);
assign n20 = ~(n1283 ^ n903);
assign n995 = ~n498;
assign n1289 = n543 & n971;
assign n293 = n549 | n692;
assign n352 = ~(n1215 | n428);
assign n1176 = ~(n1022 & n839);
assign n1306 = n290 & n936;
assign n99 = n299 & n349;
assign n1299 = n1287 & n1233;
assign n496 = ~(n701 | n1254);
assign n943 = ~n650;
assign n266 = ~(n874 | n876);
assign n1268 = ~n1285;
assign n1323 = ~(n1190 ^ n462);
assign n251 = ~(n922 ^ n286);
assign n754 = ~n782;
assign n1275 = n1148;
assign n162 = ~n582;
assign n772 = ~n261;
assign n396 = ~(n775 ^ n933);
assign n403 = n1250;
assign n1001 = n1314 | n406;
assign n778 = ~(n689 | n531);
assign n1224 = n773 | n709;
assign n1166 = n1000 | n445;
assign n114 = ~n187;
assign n1076 = n669 & n255;
assign n541 = n664 | n50;
assign n31 = ~n51;
assign n757 = ~(n953 ^ n988);
assign n463 = ~(n1115 | n113);
assign n1205 = n1250;
assign n14 = ~n1104;
assign n409 = ~(n633 | n318);
assign n1237 = n110 & n216;
assign n1337 = n994 | n442;
assign n562 = n361 ^ n449;
assign n782 = ~n941;
assign n641 = ~(n660 ^ n1046);
assign n72 = ~n832;
assign n569 = ~n172;
assign n629 = n1106 & n555;
assign n299 = n1352 | n730;
assign n194 = n557 ^ n523;
assign n1034 = n1272 | n242;
assign n379 = ~(n1289 | n300);
assign n601 = n459 | n512;
assign n887 = n465 & n468;
assign n618 = n436 & n368;
assign n1291 = ~n390;
assign n1213 = ~n73;
assign n559 = ~(n1162 ^ n1173);
assign n228 = n238 & n883;
assign n308 = ~(n372 ^ n149);
assign n1173 = ~(n188 ^ n477);
assign n1307 = ~n655;
assign n573 = ~(n645 ^ n181);
assign n581 = n776 & n1298;
assign n1038 = n737 | n675;
assign n1256 = n561 & n857;
assign n1039 = ~(n720 ^ n107);
assign n1117 = ~(n821 ^ n721);
assign n342 = n299;
assign n10 = n424 & n86;
assign n596 = n1201;
assign n953 = n224 | n46;
assign n864 = n846 & n246;
assign n886 = ~n648;
assign n292 = ~(n480 ^ n1035);
assign n296 = ~(n425 ^ n546);
assign n504 = ~(n1009 ^ n353);
assign n1160 = n1161 & n677;
assign n922 = ~(n1207 ^ n949);
assign n230 = n688 | n121;
assign n918 = n1242 & n1266;
assign n694 = ~(n1084 ^ n997);
assign n888 = n294 & n376;
assign n985 = ~n1241;
assign n516 = n301;
assign n405 = ~(n449 | n403);
assign n322 = n688 | n490;
assign n373 = ~(n1124 | n8);
assign n791 = n305 & n688;
assign n1078 = ~n508;
assign n456 = n215 | n115;
assign n789 = n846 & n841;
assign n977 = ~n681;
assign n369 = ~(n603 | n248);
assign n435 = ~n146;
assign n1228 = n1341 | n1127;
assign n489 = n1219 & n688;
assign n1217 = n1035 | n179;
assign n225 = n63 | n1165;
assign n950 = n846 & n929;
assign n378 = ~n365;
assign n436 = ~n751;
assign n1171 = ~(n1340 ^ n660);
assign n1325 = n848 | n285;
assign n1127 = n4 | n87;
assign n214 = n872 & n61;
assign n419 = n937 & n788;
assign n1314 = n1049 & n1120;
assign n844 = n403 & n1229;
assign n676 = n346 | n715;
assign n1204 = n629 & n402;
assign n544 = n1331 | n563;
assign n440 = n460 & n363;
assign n302 = n871 | n924;
assign n560 = n1013 & n392;
assign n588 = ~(n104 | n403);
assign n904 = ~(n184 ^ n1135);
assign n1046 = ~(n565 ^ n552);
assign n669 = ~n498;
assign n820 = n402 ^ n1001;
assign n335 = n107 | n1049;
assign n1149 = ~n1076;
assign n291 = n1305 | n844;
assign n276 = n35 | n769;
assign n446 = n1078 | n1249;
assign n1215 = ~n473;
assign n416 = n138 | n412;
assign n617 = n598;
assign n1309 = n146 & n1197;
assign n637 = ~(n664 ^ n1090);
assign n528 = n1276 | n1275;
assign n781 = n1308 | n1049;
assign n817 = n1260 & n493;
assign n215 = ~(n1160 | n451);
assign n1027 = n671 & n1221;
assign n974 = n1028 & n926;
assign n742 = ~n529;
assign n712 = ~n487;
assign n660 = n992 & n230;
assign n370 = ~(n1249 | n27);
assign n699 = ~n1345;
assign n1148 = ~n237;
assign n858 = n126 ^ n282;
assign n545 = n1267 & n1254;
assign n868 = n38 | n612;
assign n59 = ~n1041;
assign n412 = n125 & n80;
assign n1110 = ~n1021;
assign n524 = ~n1346;
assign n81 = ~(n495 ^ n351);
assign n994 = n9 & n1188;
assign n451 = n1283 | n55;
assign n883 = n822 | n805;
assign n801 = ~n385;
assign n1241 = n515 & n1284;
assign n159 = 1'b0;
assign n558 = ~n687;
assign n508 = ~(n938 ^ n45);
assign n182 = n403 & n1072;
assign n726 = ~(n1022 ^ n839);
assign n287 = ~n786;
assign n298 = ~(n587 ^ n97);
assign n808 = ~(n106 ^ n991);
assign n285 = n1296;
assign n979 = n140 | n914;
assign n877 = n679;
assign n1263 = ~n171;
assign n166 = n688 & n128;
assign n1156 = n422 ^ n41;
assign n1071 = ~(n1175 | n1068);
assign n1221 = n1029 & n952;
assign n551 = ~n239;
assign n875 = ~n1095;
assign n410 = 1'b0;
assign n1318 = ~(n234 | n549);
assign n627 = ~(n524 ^ n624);
assign n144 = ~(n775 ^ n393);
assign n1096 = ~(n1130 ^ n596);
assign n872 = n1252 | n380;
assign n720 = n256 & n859;
assign n96 = ~(n770 ^ n702);
assign n1242 = n488 & n868;
assign n574 = ~(n560 | n379);
assign n1324 = n537 | n1049;
assign n358 = n836 & n398;
assign n311 = ~(n960 ^ n1086);
assign n813 = n136 | n674;
assign n620 = ~n33;
assign n722 = ~(n673 ^ n858);
assign n860 = n968 & n940;
assign n960 = ~(n163 | n486);
assign n92 = ~(n481 | n974);
assign n1282 = n1080 & n688;
assign n1348 = ~n1145;
assign n110 = n12 & n797;
assign n259 = n1185 ^ n419;
assign n1008 = ~(n247 | n137);
assign n1261 = ~(n94 ^ n988);
assign n420 = ~(n311 ^ n1258);
assign n79 = n335 & n1196;
assign n1070 = n985 & n1218;
assign n1009 = n1335 & n1149;
assign n962 = ~(n941 ^ n373);
assign n1195 = n823 & n688;
assign n1032 = n1112 | n605;
assign n707 = ~(n523 ^ n465);
assign n1075 = ~n591;
assign n729 = n12 & n216;
assign n48 = ~(n434 | n273);
assign n939 = n1174 ^ n847;
assign n1304 = n1252 ^ n375;
assign n61 = n360 | n1058;
assign n531 = n809 | n203;
assign n78 = ~(n528 ^ n1325);
assign n193 = n644;
assign n647 = n324 & n577;
assign n597 = n1344 & n802;
assign n912 = ~(n1235 | n172);
assign n351 = n1040 | n211;
assign n425 = ~(n388 | n1343);
assign n432 = n976 | n127;
assign n69 = ~n1005;
assign n233 = ~n866;
assign n1313 = n816 | n1210;
assign n903 = n169 | n513;
assign n914 = ~n417;
assign n386 = ~(n376 | n294);
assign n795 = ~(n269 ^ n483);
assign n835 = ~(n687 ^ n990);
assign n711 = ~n666;
assign n1065 = ~(n151 ^ n1297);
assign n1346 = ~n1014;
assign n616 = ~n1131;
assign n981 = ~n473;
assign n86 = ~(n386 | n760);
assign n675 = ~n1161;
assign n1230 = ~(n1019 ^ n811);
assign n2 = ~(n1223 ^ n325);
assign n493 = ~(n658 ^ n348);
assign n1014 = ~n562;
assign n530 = ~(n603 ^ n1016);
assign n1093 = n826 & n688;
assign n362 = ~(n101 ^ n171);
assign n880 = n846 & n309;
assign n395 = n705 & n755;
assign n892 = ~(n1160 | n55);
assign n327 = n1308 | n586;
assign n1181 = ~n713;
assign n1351 = ~n1039;
assign n294 = n628 | n1275;
assign n1019 = n186 & n470;
assign n394 = ~(n989 | n1119);
assign n314 = n301 | n1049;
assign n103 = ~n262;
assign n499 = ~(n1304 ^ n994);
assign n154 = ~n869;
assign n1157 = n1049 & n879;
assign n278 = ~n258;
assign n1184 = ~n862;
assign n623 = 1'b0;
assign n919 = ~n177;
assign n664 = n781 & n1102;
assign n621 = ~(n126 ^ n918);
assign n989 = ~n894;
assign n1170 = n724 | n114;
assign n625 = ~n80;
assign n41 = n1227 ^ n183;
assign n665 = ~n1224;
assign n567 = ~n986;
assign n1238 = ~(n1084 ^ n865);
assign n622 = ~(n899 ^ n931);
assign n283 = ~n108;
assign n564 = ~(n1172 ^ n235);
assign n796 = n556;
assign n1190 = n752 | n1074;
assign n157 = ~n569;
assign n1193 = n1111 | n719;
assign n546 = ~(n468 ^ n1247);
assign n339 = n688 | n804;
assign n807 = n45;
assign n1270 = n407 ^ n716;
assign n273 = ~(n944 | n93);
assign n1335 = n649 & n377;
assign n13 = n648 | n925;
assign n1102 = n688 | n1328;
assign n550 = ~n977;
assign n710 = n36;
assign n713 = n572 | n1204;
assign n937 = ~n527;
assign n39 = ~n558;
assign n1183 = n932 & n155;
assign n401 = n688 | n69;
assign n916 = ~(n533 | n578);
assign n677 = n64 | n1049;
assign n155 = n10 & n886;
assign n547 = ~n1180;
assign n105 = ~(n23 ^ n856);
assign n681 = n1170 & n327;
assign n428 = n1119 & n1300;
assign n1011 = n331 & n593;
assign n1115 = ~(n596 | n784);
assign n1232 = n268;
assign n312 = ~n341;
assign n760 = ~(n831 | n1062);
assign n470 = n972 | n846;
assign n473 = n967 & n568;
assign n843 = n1205 & n200;
assign n204 = n337 | n141;
assign n728 = n547 | n1049;
assign n458 = ~n934;
assign n646 = n924 & n474;
assign n414 = ~(n334 ^ n1168);
assign n543 = n74 & n479;
assign n930 = n85 & n653;
assign n1300 = n1280 & n495;
assign n831 = n688 | n519;
assign n1138 = n846 & n260;
assign n963 = n1036 & n688;
assign n202 = n111 | n189;
assign n263 = n1306 | n1275;
assign n619 = ~(n1291 ^ n783);
assign n40 = ~n1340;
assign n982 = ~(n819 | n846);
assign n848 = n1033 & n896;
assign n542 = ~(n920 | n1001);
assign n1167 = n668 | n1157;
assign n1297 = ~(n1160 ^ n1107);
assign n876 = ~n738;
assign n141 = n162 & n937;
assign n1194 = n116;
assign n349 = ~n730;
assign n814 = ~n796;
assign n662 = ~(n508 ^ n277);
assign n73 = n548 & n1066;
assign n1161 = n688 | n1024;
assign n453 = n288 & n359;
assign n1025 = n290 & n599;
assign n1295 = ~(n906 ^ n306);
assign n611 = ~n94;
assign n11 = n874 ^ n738;
assign n468 = ~n523;
assign n150 = n642 | n1334;
assign n579 = n657 & n688;
assign n747 = ~(n1169 ^ n26);
assign n972 = ~n806;
assign n1062 = n329 | n285;
assign n331 = n716 | n403;
assign n1210 = ~(n18 | n62);
assign n320 = ~(n798 ^ n882);
assign n759 = ~n845;
assign n455 = ~(n89 ^ n249);
assign n958 = n1321 | n594;
assign n16 = ~(n1294 | n213);
assign n261 = n199 & n145;
assign n1320 = ~n198;
assign n363 = n688 | n503;
assign n539 = n1064 & n688;
assign n763 = ~(n681 ^ n1199);
assign n181 = ~(n44 ^ n1243);
assign n1128 = n1167 ^ n603;
assign n12 = n736 & n1234;
assign n1047 = ~n56;
assign n838 = ~(n596 | n123);
assign n355 = ~n1151;
assign n484 = n21 & n1226;
assign n1220 = ~(n397 | n698);
assign n1343 = n899 & n562;
assign n83 = ~n1038;
assign n400 = n9 ^ n1304;
assign n668 = n366 & n688;
assign n408 = n978 & n654;
assign n743 = ~(n36 | n1205);
assign n316 = n1049 & n1143;
assign n1294 = n864 | n884;
assign n237 = ~n1296;
assign n537 = ~n98;
assign n274 = n403 & n1141;
assign n346 = n1291 & n1224;
assign n1003 = n332 | n846;
assign n735 = n1082 | n686;
assign n160 = n1205 & n1231;
assign n389 = n515 | n68;
assign n693 = n428 & n265;
assign n1053 = n1033 & n771;
assign n447 = n688 & n767;
assign n692 = ~n860;
assign n135 = ~(n669 ^ n172);
assign n28 = n107 | n534;
assign n94 = n1353 | n1074;
assign n411 = ~(n1203 | n1063);
assign n1199 = ~(n1310 ^ n1096);
assign n908 = n801;
assign n527 = ~n257;
assign n1234 = n317 ^ n1118;
assign n1200 = ~(n1263 ^ n530);
assign n68 = ~(n1222 | n545);
assign n512 = n1205 & n536;
assign n1051 = ~n796;
assign n8 = n106 & n416;
assign n1134 = ~(n440 ^ n1302);
assign n212 = n502 | n1169;
assign n1063 = ~n543;
assign n885 = ~(n92 | n748);
assign n1017 = ~(n205 ^ n664);
assign n343 = ~(n768 | n815);
assign n1174 = ~(n480 ^ n170);
assign n365 = ~n1251;
assign n594 = ~n356;
assign n35 = ~(n399 | n458);
assign n1111 = ~(n1255 | n624);
assign n457 = ~n157;
assign n452 = n393;
assign n1182 = n902 & n25;
assign n338 = ~(n532 | n880);
assign n173 = n1237 | n676;
assign n476 = ~(n266 | n15);
assign n143 = n1128 | n362;
assign n156 = n1146 & n688;
assign n1179 = ~n825;
assign n633 = ~(n78 ^ n1070);
assign n1288 = n1035;
assign n727 = n391 & n596;
assign n137 = ~n184;
assign n869 = ~n1294;
assign n113 = ~n282;
assign n102 = ~n186;
assign n917 = ~(n231 | n443);
assign n725 = n956 | n704;
assign n935 = n247 ^ n184;
assign n598 = n127 | n606;
assign n140 = ~(n1055 | n837);
assign n957 = ~(n368 ^ n526);
assign n142 = ~n1104;
assign n329 = n1051 & n284;
assign n353 = n558 ^ n942;
assign n65 = n714 & n688;
assign n43 = n403 & n640;
assign n1101 = n724 | n1266;
assign n603 = n314 & n401;
assign n1206 = 1'b0;
assign n1124 = n72 & n1007;
assign n240 = ~(n48 ^ n570);
assign n1207 = n810 | n789;
assign n535 = ~(n712 ^ n1133);
assign n46 = ~(n38 | n1049);
assign n1147 = ~n1352;
assign n1214 = ~(n1067 | n403);
assign n514 = n341 ^ n644;
assign n1152 = ~(n673 ^ n463);
assign n777 = ~n253;
assign n1244 = ~(n596 | n201);
assign n856 = ~(n354 ^ n56);
assign n1095 = ~n1345;
assign n606 = ~(n787 & n491);
assign n34 = n116;
assign n555 = ~(n399 ^ n934);
assign n968 = n1049 & n685;
assign n399 = ~n466;
assign n920 = n791 | n625;
assign n275 = n1277;
assign n387 = n467 & n39;
assign n769 = n713 & n1246;
assign n649 = n147 | n1043;
assign n1331 = ~n292;
assign n88 = 1'b0;
assign n1227 = ~n585;
assign n874 = ~n44;
assign n1339 = ~n667;
assign n23 = ~(n1038 ^ n450);
assign n987 = n861 | n551;
assign n899 = n981 ^ n989;
assign n612 = n529 & n148;
assign n905 = ~(n1227 ^ n686);
assign n424 = ~(n533 | n615);
assign n321 = ~(n566 ^ n1281);
assign n605 = ~(n560 | n916);
assign n124 = n930 & n999;
assign n891 = n951 & n297;
assign n526 = ~(n964 | n1244);
assign n146 = n688 | n158;
assign n1158 = n1327 | n843;
assign n1023 = n38;
assign n250 = n1060 & n975;
assign n630 = n161 & n226;
assign n548 = n688 | n355;
assign n1122 = ~(n1220 ^ n969);
assign n828 = ~(n361 ^ n1177);
assign n898 = ~(n109 ^ n828);
assign n479 = ~(n25 ^ n1011);
assign n1136 = ~n951;
assign n169 = ~(n1342 | n1205);
assign n945 = ~n694;
assign n1013 = n1172 | n1338;
assign n517 = ~(n880 ^ n506);
assign n800 = ~n961;
assign n1249 = n754 | n1007;
assign n380 = ~n1075;
assign n679 = ~n385;
assign n730 = n1241 & n684;
assign n873 = n758 & n291;
assign n1118 = ~n665;
assign n724 = n604 ^ n1308;
assign n794 = ~(n483 ^ n861);
assign n723 = ~(n292 ^ n563);
assign n133 = n1318 | n113;
assign n101 = ~n1309;
assign n521 = n134 | n1182;
assign n430 = ~n525;
assign n190 = ~(n778 ^ n1193);
assign n330 = ~n756;
assign n990 = n1009 | n1;
assign n663 = ~n122;
assign n1144 = n154 ^ n811;
assign n119 = n236 & n688;
assign n1079 = n1230 | n1103;
assign n247 = n1205 & n1339;
assign n132 = ~n1037;
assign n705 = n892 | n197;
assign n797 = n1138 | n1265;
assign n651 = n1184;
assign n148 = n283 | n1049;
assign n1135 = ~(n1062 ^ n263);
assign n300 = n543 & n1208;
assign n1272 = n551 & n320;
assign n434 = n413 & n944;
assign n392 = n796 | n1299;
assign n911 = ~n548;
assign n345 = ~n344;
assign n93 = ~(n595 ^ n1006);
assign n1040 = n253 & n750;
assign n768 = n49 ^ n244;
assign n884 = ~(n231 | n1205);
assign n426 = ~(n797 ^ n803);
assign n592 = n127 | n59;
assign n255 = ~(n354 ^ n1198);
assign n1225 = ~n214;
assign n949 = n1154 | n316;
assign n933 = n919 ^ n898;
assign n328 = ~(n940 ^ n685);
assign n984 = ~(n393 | n1049);
assign n718 = n116;
assign n734 = n475;
assign n834 = n1053 | n1275;
assign n1113 = n143 | n202;
assign n1262 = ~(n251 ^ n5);
assign n466 = n489 | n182;
assign n482 = ~n1166;
assign n1347 = n1089 & n688;
assign n708 = ~n1012;
assign n44 = n156 | n357;
assign n1024 = ~n500;
assign n474 = ~n699;
assign n1114 = n32 & n144;
assign n277 = ~(n1042 | n370);
assign n407 = ~n891;
assign n494 = ~(n287 | n642);
assign n636 = n403 & n192;
assign n264 = n644 | n312;
assign n678 = n1088 | n968;
assign n1043 = ~n255;
assign n522 = ~(n934 | n466);
assign n1341 = ~(n739 | n30);
assign n852 = n688 | n103;
assign n1248 = n652 & n852;
assign n959 = n411 | n225;
assign n57 = n1300 & n378;
assign n925 = n959 & n155;
assign n966 = n107;
assign n467 = ~n1335;
assign n811 = n1003 & n1292;
endmodule
