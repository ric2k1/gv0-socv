module a;
integer [31:0]w;
endmodule

