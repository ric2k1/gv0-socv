module top(in1, in2, in3, out1, out2);
  input [7:0] in1, in2, in3;
  output [23:0] out1;
  output [15:0] out2;
  wire [7:0] in1, in2, in3;
  wire [23:0] out1;
  wire [15:0] out2;
  wire mul_7_27_n_0, mul_7_27_n_1, mul_7_27_n_2, mul_7_27_n_3, mul_7_27_n_4, mul_7_27_n_5, mul_7_27_n_9, mul_7_27_n_10;
  wire mul_7_27_n_11, mul_7_27_n_12, mul_7_27_n_13, mul_7_27_n_14, mul_7_27_n_15, mul_7_27_n_16, mul_7_27_n_17, mul_7_27_n_18;
  wire mul_7_27_n_19, mul_7_27_n_20, mul_7_27_n_21, mul_7_27_n_22, mul_7_27_n_23, mul_7_27_n_24, mul_7_27_n_25, mul_7_27_n_26;
  wire mul_7_27_n_27, mul_7_27_n_28, mul_7_27_n_29, mul_7_27_n_30, mul_7_27_n_31, mul_7_27_n_32, mul_7_27_n_33, mul_7_27_n_34;
  wire mul_7_27_n_35, mul_7_27_n_36, mul_7_27_n_37, mul_7_27_n_38, mul_7_27_n_39, mul_7_27_n_40, mul_7_27_n_41, mul_7_27_n_42;
  wire mul_7_27_n_43, mul_7_27_n_44, mul_7_27_n_45, mul_7_27_n_46, mul_7_27_n_47, mul_7_27_n_48, mul_7_27_n_49, mul_7_27_n_50;
  wire mul_7_27_n_51, mul_7_27_n_52, mul_7_27_n_53, mul_7_27_n_54, mul_7_27_n_55, mul_7_27_n_56, mul_7_27_n_57, mul_7_27_n_58;
  wire mul_7_27_n_59, mul_7_27_n_60, mul_7_27_n_61, mul_7_27_n_62, mul_7_27_n_63, mul_7_27_n_64, mul_7_27_n_65, mul_7_27_n_66;
  wire mul_7_27_n_67, mul_7_27_n_68, mul_7_27_n_69, mul_7_27_n_70, mul_7_27_n_71, mul_7_27_n_72, mul_7_27_n_73, mul_7_27_n_74;
  wire mul_7_27_n_75, mul_7_27_n_76, mul_7_27_n_77, mul_7_27_n_78, mul_7_27_n_79, mul_7_27_n_80, mul_7_27_n_81, mul_7_27_n_82;
  wire mul_7_27_n_83, mul_7_27_n_84, mul_7_27_n_85, mul_7_27_n_86, mul_7_27_n_87, mul_7_27_n_88, mul_7_27_n_89, mul_7_27_n_90;
  wire mul_7_27_n_91, mul_7_27_n_92, mul_7_27_n_93, mul_7_27_n_94, mul_7_27_n_95, mul_7_27_n_96, mul_7_27_n_97, mul_7_27_n_98;
  wire mul_7_27_n_99, mul_7_27_n_100, mul_7_27_n_101, mul_7_27_n_102, mul_7_27_n_103, mul_7_27_n_104, mul_7_27_n_105, mul_7_27_n_106;
  wire mul_7_27_n_107, mul_7_27_n_108, mul_7_27_n_109, mul_7_27_n_110, mul_7_27_n_111, mul_7_27_n_112, mul_7_27_n_113, mul_7_27_n_114;
  wire mul_7_27_n_115, mul_7_27_n_116, mul_7_27_n_117, mul_7_27_n_118, mul_7_27_n_119, mul_7_27_n_120, mul_7_27_n_121, mul_7_27_n_122;
  wire mul_7_27_n_123, mul_7_27_n_124, mul_7_27_n_125, mul_7_27_n_126, mul_7_27_n_127, mul_7_27_n_128, mul_7_27_n_129, mul_7_27_n_130;
  wire mul_7_27_n_131, mul_7_27_n_132, mul_7_27_n_133, mul_7_27_n_134, mul_7_27_n_135, mul_7_27_n_136, mul_7_27_n_137, mul_7_27_n_138;
  wire mul_7_27_n_139, mul_7_27_n_140, mul_7_27_n_141, mul_7_27_n_142, mul_7_27_n_143, mul_7_27_n_144, mul_7_27_n_145, mul_7_27_n_146;
  wire mul_7_27_n_147, mul_7_27_n_148, mul_7_27_n_149, mul_7_27_n_150, mul_7_27_n_151, mul_7_27_n_152, mul_7_27_n_153, mul_7_27_n_154;
  wire mul_7_27_n_155, mul_7_27_n_156, mul_7_27_n_157, mul_7_27_n_158, mul_7_27_n_159, mul_7_27_n_160, mul_7_27_n_161, mul_7_27_n_162;
  wire mul_7_27_n_163, mul_7_27_n_164, mul_7_27_n_165, mul_7_27_n_166, mul_7_27_n_167, mul_7_27_n_168, mul_7_27_n_169, mul_7_27_n_170;
  wire mul_7_27_n_171, mul_7_27_n_172, mul_7_27_n_173, mul_7_27_n_174, mul_7_27_n_175, mul_7_27_n_176, mul_7_27_n_177, mul_7_27_n_178;
  wire mul_7_27_n_179, mul_7_27_n_180, mul_7_27_n_181, mul_7_27_n_182, mul_7_27_n_183, mul_7_27_n_184, mul_7_27_n_185, mul_7_27_n_186;
  wire mul_7_27_n_187, mul_7_27_n_188, mul_7_27_n_189, mul_7_27_n_190, mul_7_27_n_191, mul_7_27_n_192, mul_7_27_n_193, mul_7_27_n_194;
  wire mul_7_27_n_195, mul_7_27_n_196, mul_7_27_n_197, mul_7_27_n_198, mul_7_27_n_199, mul_7_27_n_200, mul_7_27_n_201, mul_7_27_n_202;
  wire mul_7_27_n_203, mul_7_27_n_204, mul_7_27_n_205, mul_7_27_n_206, mul_7_27_n_207, mul_7_27_n_208, mul_7_27_n_209, mul_7_27_n_210;
  wire mul_7_27_n_211, mul_7_27_n_212, mul_7_27_n_213, mul_7_27_n_214, mul_7_27_n_215, mul_7_27_n_216, mul_7_27_n_217, mul_7_27_n_218;
  wire mul_7_27_n_219, mul_7_27_n_220, mul_7_27_n_221, mul_7_27_n_222, mul_7_27_n_223, mul_7_27_n_224, mul_7_27_n_225, mul_7_27_n_226;
  wire mul_7_27_n_227, mul_7_27_n_228, mul_7_27_n_229, mul_7_27_n_230, mul_7_27_n_231, mul_7_27_n_232, mul_7_27_n_233, mul_7_27_n_234;
  wire mul_7_27_n_235, mul_7_27_n_236, mul_7_27_n_237, mul_7_27_n_238, mul_7_27_n_239, mul_7_27_n_240, mul_7_27_n_241, mul_7_27_n_242;
  wire mul_7_27_n_243, mul_7_27_n_244, mul_7_27_n_245, mul_7_27_n_246, mul_7_27_n_247, mul_7_27_n_248, mul_7_27_n_249, mul_7_27_n_250;
  wire mul_7_27_n_251, mul_7_27_n_252, mul_7_27_n_253, mul_7_27_n_254, mul_7_27_n_255, mul_7_27_n_256, mul_7_27_n_257, mul_7_27_n_258;
  wire mul_7_27_n_259, mul_7_27_n_260, mul_7_27_n_261, mul_7_27_n_262, mul_7_27_n_263, mul_7_27_n_264, mul_7_27_n_265, mul_7_27_n_266;
  wire mul_7_27_n_267, mul_7_27_n_268, mul_7_27_n_269, mul_7_27_n_270, mul_7_27_n_271, mul_7_27_n_272, mul_7_27_n_273, mul_7_27_n_274;
  wire mul_7_27_n_275, mul_7_27_n_276, mul_7_27_n_277, mul_7_27_n_279, mul_7_27_n_280, mul_7_27_n_281, mul_7_27_n_282, mul_7_27_n_283;
  wire mul_7_27_n_284, mul_7_27_n_285, mul_7_27_n_286, mul_7_27_n_287, mul_7_27_n_288, mul_7_27_n_289, mul_7_27_n_290, mul_7_27_n_291;
  wire mul_7_27_n_292, mul_7_27_n_293, mul_7_27_n_294, mul_7_27_n_295, mul_7_27_n_296, mul_7_27_n_297, mul_7_27_n_298, mul_7_27_n_299;
  wire mul_7_27_n_300, mul_7_27_n_301, mul_7_27_n_302, mul_7_27_n_303, mul_7_27_n_304, mul_7_27_n_305, mul_7_27_n_306, mul_7_27_n_307;
  wire mul_7_27_n_308, mul_7_27_n_309, mul_7_27_n_310, mul_7_27_n_311, mul_7_27_n_312, mul_7_27_n_313, mul_7_27_n_314, mul_7_27_n_315;
  wire mul_7_27_n_316, mul_7_27_n_317, mul_7_27_n_318, mul_7_27_n_319, mul_7_27_n_320, mul_7_27_n_321, mul_7_27_n_322, mul_7_27_n_323;
  wire mul_7_27_n_324, mul_7_27_n_325, mul_7_27_n_326, mul_7_27_n_327, mul_7_27_n_328, mul_7_27_n_329, mul_7_27_n_330, mul_7_27_n_331;
  wire mul_7_27_n_332, mul_7_27_n_333, mul_7_27_n_334, mul_7_27_n_335, mul_7_27_n_336, mul_7_27_n_337, mul_7_27_n_338, mul_7_27_n_339;
  wire mul_7_27_n_340, mul_7_27_n_341, mul_7_27_n_342, mul_7_27_n_343, mul_7_27_n_344, mul_7_27_n_345, mul_7_27_n_346, mul_7_27_n_347;
  wire mul_7_27_n_348, mul_7_27_n_349, mul_7_27_n_350, mul_7_27_n_351, mul_7_27_n_352, mul_7_27_n_353, mul_7_27_n_354, mul_7_27_n_355;
  wire mul_7_27_n_356, mul_7_27_n_357, mul_7_27_n_358, mul_7_27_n_359, mul_7_27_n_360, mul_7_27_n_361, mul_7_27_n_362, mul_7_27_n_363;
  wire mul_7_27_n_364, mul_7_27_n_365, mul_7_27_n_366, mul_7_27_n_367, mul_7_27_n_368, mul_7_27_n_369, mul_7_27_n_370, mul_7_27_n_371;
  wire mul_7_27_n_372, mul_7_27_n_373, mul_7_27_n_374, mul_7_27_n_375, mul_7_27_n_376, mul_7_27_n_377, mul_7_27_n_378, mul_7_27_n_379;
  wire mul_7_27_n_381, mul_7_27_n_382, mul_7_27_n_383, mul_7_27_n_384, mul_7_27_n_385, mul_7_27_n_386, mul_7_27_n_387, mul_7_27_n_388;
  wire mul_7_27_n_389, mul_7_27_n_390, mul_7_27_n_391, mul_7_27_n_392, mul_7_27_n_393, mul_7_27_n_394, mul_7_27_n_395, mul_7_27_n_396;
  wire mul_7_27_n_397, mul_7_27_n_398, mul_7_27_n_399, mul_7_27_n_400, mul_7_27_n_401, mul_7_27_n_402, mul_7_27_n_403, mul_7_27_n_404;
  wire mul_7_27_n_405, mul_7_27_n_406, mul_7_27_n_407, mul_7_27_n_408, mul_7_27_n_409, mul_7_27_n_410, mul_7_27_n_411, mul_7_27_n_412;
  wire mul_7_27_n_413, mul_7_27_n_414, mul_7_27_n_415, mul_7_27_n_416, mul_7_27_n_417, mul_7_27_n_418, mul_7_27_n_419, mul_7_27_n_420;
  wire mul_7_27_n_421, mul_7_27_n_422, mul_7_27_n_423, mul_7_27_n_424, mul_7_27_n_425, mul_7_27_n_426, mul_7_27_n_427, mul_7_27_n_428;
  wire mul_7_27_n_429, mul_7_27_n_430, mul_7_27_n_431, mul_7_27_n_432, mul_7_27_n_433, mul_7_27_n_434, mul_7_27_n_435, mul_7_27_n_436;
  wire mul_7_27_n_437, mul_7_27_n_438, mul_7_27_n_439, mul_7_27_n_440, mul_7_27_n_441, mul_7_27_n_442, mul_7_27_n_443, mul_7_27_n_444;
  wire mul_7_27_n_445, mul_7_27_n_446, mul_7_27_n_447, mul_7_27_n_448, mul_7_27_n_449, mul_7_27_n_450, mul_7_27_n_451, mul_7_27_n_452;
  wire mul_7_27_n_453, mul_7_27_n_454, mul_7_27_n_455, mul_7_27_n_456, mul_7_27_n_457, mul_7_27_n_458, mul_7_27_n_459, mul_7_27_n_460;
  wire mul_7_27_n_461, mul_7_27_n_462, mul_7_27_n_463, mul_7_27_n_464, mul_7_27_n_465, mul_7_27_n_466, mul_7_27_n_467, mul_7_27_n_468;
  wire mul_7_27_n_469, mul_7_27_n_470, mul_7_27_n_471, mul_7_27_n_472, mul_7_27_n_473, mul_7_27_n_474, mul_7_27_n_475, mul_7_27_n_476;
  wire mul_7_27_n_477, mul_7_27_n_478, mul_7_27_n_479, mul_7_27_n_480, mul_7_27_n_481, mul_7_27_n_482, mul_7_27_n_483, mul_7_27_n_484;
  wire mul_7_27_n_485, mul_7_27_n_486, mul_7_27_n_487, mul_7_27_n_488, mul_7_27_n_489, mul_7_27_n_490, mul_7_27_n_491, mul_7_27_n_492;
  wire mul_7_27_n_493, mul_7_27_n_494, mul_7_27_n_495, mul_7_27_n_496, mul_7_27_n_497, mul_7_27_n_498, mul_7_27_n_499, mul_7_27_n_500;
  wire mul_7_27_n_501, mul_7_27_n_502, mul_7_27_n_503, mul_7_27_n_504, mul_7_27_n_505, mul_7_27_n_506, mul_7_27_n_507, mul_7_27_n_508;
  wire mul_7_27_n_509, mul_7_27_n_510, mul_7_27_n_511, mul_7_27_n_512, mul_7_27_n_513, mul_7_27_n_514, mul_7_27_n_515, mul_7_27_n_516;
  wire mul_7_27_n_517, mul_7_27_n_518, mul_7_27_n_519, mul_7_27_n_520, mul_7_27_n_521, mul_7_27_n_522, mul_7_27_n_523, mul_7_27_n_524;
  wire mul_7_27_n_525, mul_7_27_n_526, mul_7_27_n_527, mul_7_27_n_528, mul_7_27_n_529, mul_7_27_n_530, mul_7_27_n_531, mul_7_27_n_532;
  wire mul_7_27_n_533, mul_7_27_n_534, mul_7_27_n_535, mul_7_27_n_536, mul_7_27_n_537, mul_7_27_n_538, mul_7_27_n_539, mul_7_27_n_540;
  wire mul_7_27_n_541, mul_7_27_n_542, mul_7_27_n_543, mul_7_27_n_544, mul_7_27_n_545, mul_7_27_n_546, mul_7_27_n_547, mul_7_27_n_548;
  wire mul_7_27_n_549, mul_7_27_n_550, mul_7_27_n_551, mul_7_27_n_552, mul_7_27_n_553, mul_7_27_n_554, mul_7_27_n_555, mul_7_27_n_556;
  wire mul_7_27_n_557, mul_7_27_n_558, mul_7_27_n_559, mul_7_27_n_560, mul_7_27_n_561, mul_7_27_n_562, mul_7_27_n_563, mul_7_27_n_564;
  wire mul_7_27_n_565, mul_7_27_n_566, mul_7_27_n_567, mul_7_27_n_568, mul_7_27_n_569, mul_7_27_n_570, mul_7_27_n_571, mul_7_27_n_572;
  wire mul_7_27_n_573, mul_7_27_n_574, mul_7_27_n_575, mul_7_27_n_576, mul_7_27_n_577, mul_7_27_n_578, mul_7_27_n_579, mul_7_27_n_580;
  wire mul_7_27_n_581, mul_7_27_n_582, mul_7_27_n_583, mul_7_27_n_584, mul_7_27_n_585, mul_7_27_n_586, mul_7_27_n_587, mul_7_27_n_588;
  wire mul_7_27_n_589, mul_7_27_n_590, mul_7_27_n_591, mul_7_27_n_592, mul_7_27_n_593, mul_7_27_n_594, mul_7_27_n_595, mul_7_27_n_596;
  wire mul_7_27_n_597, mul_7_27_n_598, mul_7_27_n_599, mul_7_27_n_600, mul_7_27_n_601, mul_7_27_n_602, mul_7_27_n_603, mul_7_27_n_604;
  wire mul_7_27_n_605, mul_7_27_n_606, mul_7_27_n_607, mul_7_27_n_608, mul_7_27_n_609, mul_7_27_n_610, mul_7_27_n_611, mul_7_27_n_612;
  wire mul_7_27_n_613, mul_7_27_n_614, mul_7_27_n_615, mul_7_27_n_616, mul_7_27_n_617, mul_7_27_n_618, mul_7_27_n_619, mul_7_27_n_620;
  wire mul_7_27_n_621, mul_7_27_n_622, mul_7_27_n_623, mul_7_27_n_624, mul_7_27_n_625, mul_7_27_n_626, mul_7_27_n_627, mul_7_27_n_628;
  wire mul_7_27_n_629, mul_7_27_n_630, mul_7_27_n_631, mul_7_27_n_632, mul_7_27_n_633, mul_7_27_n_634, mul_7_27_n_635, mul_7_27_n_636;
  wire mul_7_27_n_637, mul_7_27_n_638, mul_7_27_n_639, mul_7_27_n_640, mul_7_27_n_641, mul_7_27_n_642, mul_7_27_n_643, mul_7_27_n_644;
  wire mul_7_27_n_645, mul_7_27_n_646, mul_7_27_n_647, mul_7_27_n_648, mul_7_27_n_649, mul_7_27_n_650, mul_7_27_n_651, mul_7_27_n_652;
  wire mul_7_27_n_653, mul_7_27_n_654, mul_7_27_n_655, mul_7_27_n_656, mul_7_27_n_657, mul_7_27_n_658, mul_7_27_n_659, mul_7_27_n_660;
  wire mul_7_27_n_661, mul_7_27_n_662, mul_7_27_n_663, mul_7_27_n_664, mul_7_27_n_665, mul_7_27_n_666, mul_7_27_n_667, mul_7_27_n_668;
  wire mul_7_27_n_669, mul_7_27_n_670, mul_7_27_n_671, mul_7_27_n_672, mul_7_27_n_673, mul_7_27_n_674, mul_7_27_n_675, mul_7_27_n_676;
  wire mul_7_27_n_677, mul_7_27_n_678, mul_7_27_n_679, mul_7_27_n_680, mul_7_27_n_681, mul_7_27_n_682, mul_7_27_n_683, mul_7_27_n_684;
  wire mul_7_27_n_685, mul_7_27_n_686, mul_7_27_n_687, mul_7_27_n_688, mul_7_27_n_689, mul_7_27_n_690, mul_7_27_n_691, mul_7_27_n_692;
  wire mul_7_27_n_693, mul_7_27_n_694, mul_7_27_n_695, mul_7_27_n_696, mul_7_27_n_697, mul_7_27_n_698, mul_7_27_n_699, mul_7_27_n_700;
  wire mul_7_27_n_701, mul_7_27_n_702, mul_7_27_n_703, mul_7_27_n_704, mul_7_27_n_705, mul_7_27_n_706, mul_7_27_n_707, mul_7_27_n_708;
  wire mul_7_27_n_709, mul_7_27_n_710, mul_7_27_n_711, mul_7_27_n_712, mul_7_27_n_713, mul_7_27_n_714, mul_7_27_n_715, mul_7_27_n_716;
  wire mul_7_27_n_717, mul_7_27_n_718, mul_7_27_n_719, mul_7_27_n_720, mul_7_27_n_721, mul_7_27_n_722, mul_7_27_n_723, mul_7_27_n_724;
  wire mul_7_27_n_725, mul_7_27_n_726, mul_7_27_n_727, mul_7_27_n_728, mul_7_27_n_729, mul_7_27_n_730, mul_7_27_n_731, mul_7_27_n_732;
  wire mul_7_27_n_733, mul_7_27_n_734, mul_7_27_n_735, mul_7_27_n_736, mul_7_27_n_737, mul_7_27_n_738, mul_7_27_n_739, mul_7_27_n_740;
  wire mul_7_27_n_741, mul_7_27_n_742, mul_7_27_n_743, mul_7_27_n_744, mul_7_27_n_745, mul_7_27_n_746, mul_7_27_n_747, mul_7_27_n_748;
  wire mul_7_27_n_749, mul_7_27_n_750, mul_7_27_n_751, mul_7_27_n_752, mul_7_27_n_753, mul_7_27_n_754, mul_7_27_n_755, mul_7_27_n_756;
  wire mul_7_27_n_757, mul_7_27_n_758, mul_7_27_n_759, mul_7_27_n_760, mul_7_27_n_761, mul_7_27_n_762, mul_7_27_n_763, mul_7_27_n_764;
  wire mul_7_27_n_765, mul_7_27_n_766, mul_7_27_n_767, mul_7_27_n_768, mul_7_27_n_769, mul_7_27_n_770, mul_7_27_n_771, mul_7_27_n_772;
  wire mul_7_27_n_773, mul_7_27_n_774, mul_7_27_n_775, mul_7_27_n_776, mul_7_27_n_777, mul_7_27_n_778, mul_7_27_n_779, mul_7_27_n_780;
  wire mul_7_27_n_781, mul_7_27_n_782, mul_7_27_n_783, mul_7_27_n_784, mul_7_27_n_786, mul_7_27_n_787, mul_7_27_n_788, mul_7_27_n_789;
  wire mul_7_27_n_790, mul_7_27_n_791, mul_7_27_n_792, mul_7_27_n_793, mul_7_27_n_794, mul_7_27_n_795, mul_7_27_n_796, mul_7_27_n_797;
  wire mul_7_27_n_798, mul_7_27_n_799, mul_7_27_n_800, mul_7_27_n_801, mul_7_27_n_802, mul_7_27_n_803, mul_7_27_n_804, mul_7_27_n_805;
  wire mul_7_27_n_806, mul_7_27_n_807, mul_7_27_n_808, mul_7_27_n_809, mul_7_27_n_810, mul_7_27_n_811, mul_7_27_n_812, mul_7_27_n_813;
  wire mul_7_27_n_814, mul_7_27_n_815, mul_7_27_n_816, mul_7_27_n_817, mul_7_27_n_818, mul_7_27_n_819, mul_7_27_n_820, mul_7_27_n_821;
  wire mul_7_27_n_822, mul_7_27_n_823, mul_7_27_n_824, mul_7_27_n_825, mul_7_27_n_826, mul_7_27_n_827, mul_7_27_n_828, mul_7_27_n_829;
  wire mul_7_27_n_830, mul_7_27_n_831, mul_7_27_n_832, mul_7_27_n_833, mul_7_27_n_834, mul_7_27_n_835, mul_7_27_n_836, mul_7_27_n_837;
  wire mul_7_27_n_838, mul_7_27_n_839, mul_7_27_n_840, mul_7_27_n_842, mul_7_27_n_843, mul_7_27_n_844, mul_7_27_n_845, mul_7_27_n_846;
  wire mul_7_27_n_847, mul_7_27_n_848, mul_7_27_n_849, mul_7_27_n_850, mul_7_27_n_851, mul_7_27_n_852, mul_7_27_n_853, mul_7_27_n_854;
  wire mul_7_27_n_855, mul_7_27_n_856, mul_7_27_n_857, mul_7_27_n_858, mul_7_27_n_859, mul_7_27_n_860, mul_7_27_n_861, mul_7_27_n_862;
  wire mul_7_27_n_863, mul_7_27_n_864, mul_7_27_n_865, mul_7_27_n_866, mul_7_27_n_867, mul_7_27_n_868, mul_7_27_n_869, mul_7_27_n_870;
  wire mul_7_27_n_871, mul_7_27_n_872, mul_7_27_n_873, mul_7_27_n_874, mul_7_27_n_875, mul_7_27_n_876, mul_7_27_n_877, mul_7_27_n_878;
  wire mul_7_27_n_879, mul_7_27_n_880, mul_7_27_n_881, mul_7_27_n_882, mul_7_27_n_883, mul_7_27_n_884, mul_7_27_n_885, mul_7_27_n_886;
  wire mul_7_27_n_887, mul_7_27_n_888, mul_7_27_n_889, mul_7_27_n_890, mul_7_27_n_891, mul_7_27_n_892, mul_7_27_n_893, mul_7_27_n_894;
  wire mul_7_27_n_895, mul_7_27_n_896, mul_7_27_n_897, mul_7_27_n_898, mul_7_27_n_899, mul_7_27_n_900, mul_7_27_n_901, mul_7_27_n_902;
  wire mul_7_27_n_903, mul_7_27_n_904, mul_7_27_n_905, mul_7_27_n_906, mul_7_27_n_907, mul_7_27_n_908, mul_7_27_n_909, mul_7_27_n_910;
  wire mul_7_27_n_911, mul_7_27_n_913, mul_7_27_n_914, mul_7_27_n_915, mul_7_27_n_916, mul_7_27_n_917, mul_7_27_n_918, mul_7_27_n_919;
  wire mul_7_27_n_920, mul_7_27_n_921, mul_7_27_n_922, mul_7_27_n_923, mul_7_27_n_924, mul_7_27_n_925, mul_7_27_n_926, mul_7_27_n_927;
  wire mul_7_27_n_928, mul_7_27_n_929, mul_7_27_n_930, mul_7_27_n_931, mul_7_27_n_932, mul_7_27_n_933, mul_7_27_n_934, mul_7_27_n_935;
  wire mul_7_27_n_936, mul_7_27_n_937, mul_7_27_n_938, mul_7_27_n_939, mul_7_27_n_940, mul_7_27_n_941, mul_7_27_n_942, mul_7_27_n_943;
  wire mul_7_27_n_944, mul_7_27_n_945, mul_7_27_n_946, mul_7_27_n_947, mul_7_27_n_948, mul_7_27_n_949, mul_7_27_n_950, mul_7_27_n_951;
  wire mul_7_27_n_952, mul_7_27_n_953, mul_7_27_n_954, mul_7_27_n_955, mul_7_27_n_956, mul_7_27_n_957, mul_7_27_n_958, mul_7_27_n_959;
  wire mul_7_27_n_960, mul_7_27_n_961, mul_7_27_n_962, mul_7_27_n_963, mul_7_27_n_964, mul_7_27_n_965, mul_7_27_n_966, mul_7_27_n_967;
  wire mul_7_27_n_968, mul_7_27_n_969, mul_7_27_n_970, mul_7_27_n_972, mul_7_27_n_973, mul_7_27_n_974, mul_7_27_n_975, mul_7_27_n_976;
  wire mul_7_27_n_977, mul_7_27_n_978, mul_7_27_n_979, mul_7_27_n_980, mul_7_27_n_981, mul_7_27_n_982, mul_7_27_n_983, mul_7_27_n_984;
  wire mul_7_27_n_985, mul_7_27_n_986, mul_7_27_n_987, mul_7_27_n_988, mul_7_27_n_989, mul_7_27_n_990, mul_7_27_n_991, mul_7_27_n_992;
  wire mul_7_27_n_993, mul_7_27_n_994, mul_7_27_n_995, mul_7_27_n_996, mul_7_27_n_997, mul_7_27_n_998, mul_7_27_n_999, mul_7_27_n_1001;
  wire mul_7_27_n_1002, mul_7_27_n_1004, mul_7_27_n_1005, mul_7_27_n_1007, mul_7_27_n_1008, mul_7_27_n_1010, mul_7_27_n_1011, mul_7_27_n_1013;
  wire mul_7_27_n_1014, mul_7_27_n_1016, mul_7_27_n_1017, mul_7_27_n_1019, mul_7_27_n_1020, mul_7_27_n_1021, mul_7_27_n_1022, mul_7_27_n_1023;
  wire mul_7_27_n_1024, mul_7_27_n_1025, mul_7_27_n_1026, mul_7_27_n_1028, mul_7_27_n_1029, mul_7_27_n_1031, mul_7_27_n_1032, mul_7_27_n_1034;
  wire mul_7_27_n_1035, mul_7_27_n_1037, mul_7_27_n_1038, mul_7_27_n_1040, mul_7_27_n_1041, mul_7_27_n_1043, mul_7_27_n_1044, mul_7_27_n_1046;
  wire mul_8_23_n_0, mul_8_23_n_1, mul_8_23_n_2, mul_8_23_n_3, mul_8_23_n_4, mul_8_23_n_5, mul_8_23_n_6, mul_8_23_n_7;
  wire mul_8_23_n_8, mul_8_23_n_9, mul_8_23_n_10, mul_8_23_n_11, mul_8_23_n_12, mul_8_23_n_13, mul_8_23_n_14, mul_8_23_n_15;
  wire mul_8_23_n_16, mul_8_23_n_17, mul_8_23_n_18, mul_8_23_n_19, mul_8_23_n_20, mul_8_23_n_21, mul_8_23_n_22, mul_8_23_n_23;
  wire mul_8_23_n_24, mul_8_23_n_25, mul_8_23_n_26, mul_8_23_n_27, mul_8_23_n_28, mul_8_23_n_29, mul_8_23_n_30, mul_8_23_n_31;
  wire mul_8_23_n_32, mul_8_23_n_33, mul_8_23_n_34, mul_8_23_n_35, mul_8_23_n_36, mul_8_23_n_37, mul_8_23_n_38, mul_8_23_n_39;
  wire mul_8_23_n_40, mul_8_23_n_41, mul_8_23_n_42, mul_8_23_n_43, mul_8_23_n_44, mul_8_23_n_45, mul_8_23_n_46, mul_8_23_n_47;
  wire mul_8_23_n_48, mul_8_23_n_49, mul_8_23_n_50, mul_8_23_n_51, mul_8_23_n_52, mul_8_23_n_53, mul_8_23_n_54, mul_8_23_n_55;
  wire mul_8_23_n_56, mul_8_23_n_57, mul_8_23_n_58, mul_8_23_n_59, mul_8_23_n_60, mul_8_23_n_61, mul_8_23_n_62, mul_8_23_n_63;
  wire mul_8_23_n_64, mul_8_23_n_65, mul_8_23_n_66, mul_8_23_n_67, mul_8_23_n_68, mul_8_23_n_69, mul_8_23_n_70, mul_8_23_n_71;
  wire mul_8_23_n_72, mul_8_23_n_73, mul_8_23_n_74, mul_8_23_n_75, mul_8_23_n_76, mul_8_23_n_77, mul_8_23_n_78, mul_8_23_n_79;
  wire mul_8_23_n_80, mul_8_23_n_81, mul_8_23_n_82, mul_8_23_n_83, mul_8_23_n_84, mul_8_23_n_85, mul_8_23_n_87, mul_8_23_n_88;
  wire mul_8_23_n_89, mul_8_23_n_90, mul_8_23_n_91, mul_8_23_n_92, mul_8_23_n_93, mul_8_23_n_94, mul_8_23_n_95, mul_8_23_n_96;
  wire mul_8_23_n_97, mul_8_23_n_98, mul_8_23_n_99, mul_8_23_n_100, mul_8_23_n_101, mul_8_23_n_102, mul_8_23_n_103, mul_8_23_n_104;
  wire mul_8_23_n_105, mul_8_23_n_106, mul_8_23_n_107, mul_8_23_n_108, mul_8_23_n_109, mul_8_23_n_110, mul_8_23_n_111, mul_8_23_n_112;
  wire mul_8_23_n_113, mul_8_23_n_114, mul_8_23_n_115, mul_8_23_n_116, mul_8_23_n_117, mul_8_23_n_118, mul_8_23_n_119, mul_8_23_n_120;
  wire mul_8_23_n_121, mul_8_23_n_122, mul_8_23_n_123, mul_8_23_n_124, mul_8_23_n_125, mul_8_23_n_126, mul_8_23_n_127, mul_8_23_n_128;
  wire mul_8_23_n_129, mul_8_23_n_130, mul_8_23_n_131, mul_8_23_n_132, mul_8_23_n_133, mul_8_23_n_134, mul_8_23_n_135, mul_8_23_n_136;
  wire mul_8_23_n_137, mul_8_23_n_138, mul_8_23_n_139, mul_8_23_n_140, mul_8_23_n_141, mul_8_23_n_142, mul_8_23_n_143, mul_8_23_n_144;
  wire mul_8_23_n_145, mul_8_23_n_146, mul_8_23_n_147, mul_8_23_n_148, mul_8_23_n_149, mul_8_23_n_150, mul_8_23_n_151, mul_8_23_n_152;
  wire mul_8_23_n_153, mul_8_23_n_154, mul_8_23_n_155, mul_8_23_n_156, mul_8_23_n_157, mul_8_23_n_158, mul_8_23_n_159, mul_8_23_n_160;
  wire mul_8_23_n_161, mul_8_23_n_162, mul_8_23_n_163, mul_8_23_n_164, mul_8_23_n_165, mul_8_23_n_166, mul_8_23_n_167, mul_8_23_n_168;
  wire mul_8_23_n_169, mul_8_23_n_170, mul_8_23_n_171, mul_8_23_n_172, mul_8_23_n_173, mul_8_23_n_174, mul_8_23_n_175, mul_8_23_n_176;
  wire mul_8_23_n_177, mul_8_23_n_178, mul_8_23_n_179, mul_8_23_n_180, mul_8_23_n_181, mul_8_23_n_182, mul_8_23_n_183, mul_8_23_n_184;
  wire mul_8_23_n_185, mul_8_23_n_186, mul_8_23_n_187, mul_8_23_n_188, mul_8_23_n_189, mul_8_23_n_190, mul_8_23_n_191, mul_8_23_n_192;
  wire mul_8_23_n_193, mul_8_23_n_194, mul_8_23_n_195, mul_8_23_n_196, mul_8_23_n_197, mul_8_23_n_198, mul_8_23_n_199, mul_8_23_n_200;
  wire mul_8_23_n_201, mul_8_23_n_202, mul_8_23_n_203, mul_8_23_n_204, mul_8_23_n_205, mul_8_23_n_206, mul_8_23_n_207, mul_8_23_n_208;
  wire mul_8_23_n_209, mul_8_23_n_210, mul_8_23_n_211, mul_8_23_n_212, mul_8_23_n_213, mul_8_23_n_214, mul_8_23_n_215, mul_8_23_n_216;
  wire mul_8_23_n_217, mul_8_23_n_218, mul_8_23_n_219, mul_8_23_n_220, mul_8_23_n_221, mul_8_23_n_222, mul_8_23_n_223, mul_8_23_n_224;
  wire mul_8_23_n_225, mul_8_23_n_226, mul_8_23_n_227, mul_8_23_n_228, mul_8_23_n_229, mul_8_23_n_230, mul_8_23_n_231, mul_8_23_n_232;
  wire mul_8_23_n_233, mul_8_23_n_234, mul_8_23_n_235, mul_8_23_n_236, mul_8_23_n_237, mul_8_23_n_238, mul_8_23_n_239, mul_8_23_n_240;
  wire mul_8_23_n_241, mul_8_23_n_242, mul_8_23_n_243, mul_8_23_n_244, mul_8_23_n_245, mul_8_23_n_246, mul_8_23_n_247, mul_8_23_n_248;
  wire mul_8_23_n_250, mul_8_23_n_251, mul_8_23_n_252, mul_8_23_n_253, mul_8_23_n_254, mul_8_23_n_255, mul_8_23_n_256, mul_8_23_n_257;
  wire mul_8_23_n_258, mul_8_23_n_259, mul_8_23_n_260, mul_8_23_n_261, mul_8_23_n_262, mul_8_23_n_263, mul_8_23_n_264, mul_8_23_n_265;
  wire mul_8_23_n_266, mul_8_23_n_267, mul_8_23_n_269, mul_8_23_n_270, mul_8_23_n_271, mul_8_23_n_272, mul_8_23_n_273, mul_8_23_n_274;
  wire mul_8_23_n_275, mul_8_23_n_276, mul_8_23_n_277, mul_8_23_n_278, mul_8_23_n_279, mul_8_23_n_280, mul_8_23_n_281, mul_8_23_n_282;
  wire mul_8_23_n_283, mul_8_23_n_284, mul_8_23_n_285, mul_8_23_n_286, mul_8_23_n_287, mul_8_23_n_288, mul_8_23_n_289, mul_8_23_n_290;
  wire mul_8_23_n_291, mul_8_23_n_292, mul_8_23_n_293, mul_8_23_n_294, mul_8_23_n_295, mul_8_23_n_296, mul_8_23_n_297, mul_8_23_n_298;
  wire mul_8_23_n_299, mul_8_23_n_300, mul_8_23_n_301, mul_8_23_n_302, mul_8_23_n_303, mul_8_23_n_304, mul_8_23_n_305, mul_8_23_n_306;
  wire mul_8_23_n_307, mul_8_23_n_308, mul_8_23_n_309, mul_8_23_n_310, mul_8_23_n_311, mul_8_23_n_312, mul_8_23_n_313, mul_8_23_n_314;
  wire mul_8_23_n_315, mul_8_23_n_316, mul_8_23_n_317, mul_8_23_n_318, mul_8_23_n_319, mul_8_23_n_320, mul_8_23_n_321, mul_8_23_n_322;
  wire mul_8_23_n_323, mul_8_23_n_324, mul_8_23_n_325, mul_8_23_n_326, mul_8_23_n_327, mul_8_23_n_328, mul_8_23_n_329, mul_8_23_n_330;
  wire mul_8_23_n_331, mul_8_23_n_332, mul_8_23_n_333, mul_8_23_n_334, mul_8_23_n_335, mul_8_23_n_336, mul_8_23_n_337, mul_8_23_n_338;
  wire mul_8_23_n_339, mul_8_23_n_340, mul_8_23_n_341, mul_8_23_n_342, mul_8_23_n_343, mul_8_23_n_344, mul_8_23_n_345, mul_8_23_n_346;
  wire mul_8_23_n_347, mul_8_23_n_348, mul_8_23_n_349, mul_8_23_n_350, mul_8_23_n_351, mul_8_23_n_352, mul_8_23_n_353, mul_8_23_n_354;
  wire mul_8_23_n_355, mul_8_23_n_356, mul_8_23_n_358, mul_8_23_n_359, mul_8_23_n_360, mul_8_23_n_361, mul_8_23_n_362, mul_8_23_n_363;
  wire mul_8_23_n_364, mul_8_23_n_365, mul_8_23_n_366, mul_8_23_n_367, mul_8_23_n_368, mul_8_23_n_369, mul_8_23_n_370, mul_8_23_n_371;
  wire mul_8_23_n_372, mul_8_23_n_373, mul_8_23_n_374, mul_8_23_n_375, mul_8_23_n_376, mul_8_23_n_377, mul_8_23_n_378, mul_8_23_n_379;
  wire mul_8_23_n_380, mul_8_23_n_381, mul_8_23_n_382, mul_8_23_n_383, mul_8_23_n_384, mul_8_23_n_385, mul_8_23_n_386, mul_8_23_n_387;
  wire mul_8_23_n_388, mul_8_23_n_389, mul_8_23_n_390, mul_8_23_n_391, mul_8_23_n_392, mul_8_23_n_393, mul_8_23_n_395, mul_8_23_n_396;
  wire mul_8_23_n_397, mul_8_23_n_398, mul_8_23_n_399, mul_8_23_n_400, mul_8_23_n_401, mul_8_23_n_402, mul_8_23_n_403, mul_8_23_n_404;
  wire mul_8_23_n_405, mul_8_23_n_406, mul_8_23_n_407, mul_8_23_n_408, mul_8_23_n_409, mul_8_23_n_410, mul_8_23_n_411, mul_8_23_n_412;
  wire mul_8_23_n_413, mul_8_23_n_414, mul_8_23_n_415, mul_8_23_n_416, mul_8_23_n_417, mul_8_23_n_418, mul_8_23_n_419, mul_8_23_n_420;
  wire mul_8_23_n_421, mul_8_23_n_422, mul_8_23_n_423, mul_8_23_n_424, mul_8_23_n_425, mul_8_23_n_426, mul_8_23_n_427, mul_8_23_n_428;
  wire mul_8_23_n_429, mul_8_23_n_430, mul_8_23_n_431, mul_8_23_n_432, mul_8_23_n_433, mul_8_23_n_434, mul_8_23_n_435, mul_8_23_n_436;
  wire mul_8_23_n_437, mul_8_23_n_439, mul_8_23_n_440, mul_8_23_n_441, mul_8_23_n_442, mul_8_23_n_443, mul_8_23_n_444, mul_8_23_n_445;
  wire mul_8_23_n_446, mul_8_23_n_447, mul_8_23_n_448, mul_8_23_n_449, mul_8_23_n_450, mul_8_23_n_451, mul_8_23_n_452, mul_8_23_n_453;
  wire mul_8_23_n_454, mul_8_23_n_455, mul_8_23_n_456, mul_8_23_n_457, mul_8_23_n_458, mul_8_23_n_459, mul_8_23_n_460, mul_8_23_n_461;
  wire mul_8_23_n_462, mul_8_23_n_463, mul_8_23_n_465, mul_8_23_n_466, mul_8_23_n_467, mul_8_23_n_468, mul_8_23_n_469, mul_8_23_n_470;
  wire mul_8_23_n_471, mul_8_23_n_472, mul_8_23_n_473, mul_8_23_n_474, mul_8_23_n_475, mul_8_23_n_477, mul_8_23_n_478, mul_8_23_n_479;
  wire mul_8_23_n_480, mul_8_23_n_481, mul_8_23_n_482, mul_8_23_n_483, mul_8_23_n_484, mul_8_23_n_485, mul_8_23_n_486, mul_8_23_n_488;
  wire mul_8_23_n_489, mul_8_23_n_491, mul_8_23_n_492, mul_8_23_n_494, mul_8_23_n_495, mul_8_23_n_497, mul_8_23_n_498, mul_8_23_n_500;
  wire mul_8_23_n_501, mul_8_23_n_503, mul_8_23_n_504, mul_8_23_n_506, mul_8_23_n_507, n_1, n_2, n_3;
  wire n_4, n_5, n_6, n_7, n_8, n_9, n_10, n_11;
  wire n_12, n_13, n_14, square_mul_7_21_n_0, square_mul_7_21_n_1, square_mul_7_21_n_2, square_mul_7_21_n_3, square_mul_7_21_n_4;
  wire square_mul_7_21_n_5, square_mul_7_21_n_6, square_mul_7_21_n_7, square_mul_7_21_n_8, square_mul_7_21_n_9, square_mul_7_21_n_10, square_mul_7_21_n_11, square_mul_7_21_n_12;
  wire square_mul_7_21_n_13, square_mul_7_21_n_14, square_mul_7_21_n_15, square_mul_7_21_n_16, square_mul_7_21_n_17, square_mul_7_21_n_18, square_mul_7_21_n_19, square_mul_7_21_n_20;
  wire square_mul_7_21_n_21, square_mul_7_21_n_22, square_mul_7_21_n_23, square_mul_7_21_n_24, square_mul_7_21_n_25, square_mul_7_21_n_26, square_mul_7_21_n_27, square_mul_7_21_n_28;
  wire square_mul_7_21_n_29, square_mul_7_21_n_30, square_mul_7_21_n_31, square_mul_7_21_n_32, square_mul_7_21_n_33, square_mul_7_21_n_34, square_mul_7_21_n_35, square_mul_7_21_n_36;
  wire square_mul_7_21_n_37, square_mul_7_21_n_38, square_mul_7_21_n_39, square_mul_7_21_n_40, square_mul_7_21_n_41, square_mul_7_21_n_42, square_mul_7_21_n_44, square_mul_7_21_n_45;
  wire square_mul_7_21_n_46, square_mul_7_21_n_47, square_mul_7_21_n_48, square_mul_7_21_n_49, square_mul_7_21_n_50, square_mul_7_21_n_51, square_mul_7_21_n_52, square_mul_7_21_n_53;
  wire square_mul_7_21_n_54, square_mul_7_21_n_55, square_mul_7_21_n_56, square_mul_7_21_n_57, square_mul_7_21_n_58, square_mul_7_21_n_59, square_mul_7_21_n_60, square_mul_7_21_n_61;
  wire square_mul_7_21_n_62, square_mul_7_21_n_63, square_mul_7_21_n_64, square_mul_7_21_n_65, square_mul_7_21_n_66, square_mul_7_21_n_67, square_mul_7_21_n_68, square_mul_7_21_n_69;
  wire square_mul_7_21_n_70, square_mul_7_21_n_71, square_mul_7_21_n_72, square_mul_7_21_n_73, square_mul_7_21_n_74, square_mul_7_21_n_75, square_mul_7_21_n_76, square_mul_7_21_n_77;
  wire square_mul_7_21_n_78, square_mul_7_21_n_79, square_mul_7_21_n_80, square_mul_7_21_n_81, square_mul_7_21_n_82, square_mul_7_21_n_83, square_mul_7_21_n_84, square_mul_7_21_n_85;
  wire square_mul_7_21_n_86, square_mul_7_21_n_87, square_mul_7_21_n_88, square_mul_7_21_n_89, square_mul_7_21_n_90, square_mul_7_21_n_91, square_mul_7_21_n_92, square_mul_7_21_n_93;
  wire square_mul_7_21_n_94, square_mul_7_21_n_95, square_mul_7_21_n_96, square_mul_7_21_n_97, square_mul_7_21_n_98, square_mul_7_21_n_99, square_mul_7_21_n_100, square_mul_7_21_n_101;
  wire square_mul_7_21_n_102, square_mul_7_21_n_103, square_mul_7_21_n_104, square_mul_7_21_n_105, square_mul_7_21_n_106, square_mul_7_21_n_107, square_mul_7_21_n_108, square_mul_7_21_n_109;
  wire square_mul_7_21_n_110, square_mul_7_21_n_111, square_mul_7_21_n_112, square_mul_7_21_n_113, square_mul_7_21_n_114, square_mul_7_21_n_115, square_mul_7_21_n_116, square_mul_7_21_n_117;
  wire square_mul_7_21_n_118, square_mul_7_21_n_119, square_mul_7_21_n_120, square_mul_7_21_n_121, square_mul_7_21_n_122, square_mul_7_21_n_123, square_mul_7_21_n_125, square_mul_7_21_n_126;
  wire square_mul_7_21_n_127, square_mul_7_21_n_128, square_mul_7_21_n_129, square_mul_7_21_n_130, square_mul_7_21_n_131, square_mul_7_21_n_132, square_mul_7_21_n_133, square_mul_7_21_n_134;
  wire square_mul_7_21_n_137, square_mul_7_21_n_138, square_mul_7_21_n_139, square_mul_7_21_n_140, square_mul_7_21_n_141, square_mul_7_21_n_142, square_mul_7_21_n_143, square_mul_7_21_n_144;
  wire square_mul_7_21_n_145, square_mul_7_21_n_146, square_mul_7_21_n_147, square_mul_7_21_n_148, square_mul_7_21_n_149, square_mul_7_21_n_150, square_mul_7_21_n_151, square_mul_7_21_n_152;
  wire square_mul_7_21_n_153, square_mul_7_21_n_154, square_mul_7_21_n_155, square_mul_7_21_n_156, square_mul_7_21_n_157, square_mul_7_21_n_158, square_mul_7_21_n_159, square_mul_7_21_n_160;
  wire square_mul_7_21_n_161, square_mul_7_21_n_162, square_mul_7_21_n_163, square_mul_7_21_n_164, square_mul_7_21_n_165, square_mul_7_21_n_166, square_mul_7_21_n_167, square_mul_7_21_n_168;
  wire square_mul_7_21_n_169, square_mul_7_21_n_170, square_mul_7_21_n_171, square_mul_7_21_n_172, square_mul_7_21_n_173, square_mul_7_21_n_174, square_mul_7_21_n_175, square_mul_7_21_n_176;
  wire square_mul_7_21_n_178, square_mul_7_21_n_179, square_mul_7_21_n_180, square_mul_7_21_n_181, square_mul_7_21_n_182, square_mul_7_21_n_183, square_mul_7_21_n_184, square_mul_7_21_n_185;
  wire square_mul_7_21_n_186, square_mul_7_21_n_187, square_mul_7_21_n_189, square_mul_7_21_n_190, square_mul_7_21_n_191, square_mul_7_21_n_192, square_mul_7_21_n_193, square_mul_7_21_n_194;
  wire square_mul_7_21_n_195, square_mul_7_21_n_196, square_mul_7_21_n_197, square_mul_7_21_n_198, square_mul_7_21_n_199, square_mul_7_21_n_200, square_mul_7_21_n_201, square_mul_7_21_n_202;
  wire square_mul_7_21_n_203, square_mul_7_21_n_204, square_mul_7_21_n_205, square_mul_7_21_n_206, square_mul_7_21_n_207, square_mul_7_21_n_208, square_mul_7_21_n_210, square_mul_7_21_n_211;
  wire square_mul_7_21_n_212, square_mul_7_21_n_213, square_mul_7_21_n_215, square_mul_7_21_n_216, square_mul_7_21_n_218, square_mul_7_21_n_219, square_mul_7_21_n_220, square_mul_7_21_n_222;
  wire square_mul_7_21_n_223, square_mul_7_21_n_225, square_mul_7_21_n_226, square_mul_7_21_n_227, square_mul_7_21_n_229, square_mul_7_21_n_230, square_mul_7_21_n_232, square_mul_7_21_n_233;
  wire square_mul_7_21_n_234, square_mul_7_21_n_236, square_mul_7_21_n_237;
  buf constbuf_n1(out1[0], in1[0]);
  xnor mul_7_27_g2715__2398(out1[23] ,mul_7_27_n_876 ,mul_7_27_n_1046);
  nor mul_7_27_g2716__5107(mul_7_27_n_1046 ,mul_7_27_n_1044 ,mul_7_27_n_894);
  xnor mul_7_27_g2717__6260(out1[22] ,mul_7_27_n_1043 ,mul_7_27_n_910);
  nor mul_7_27_g2718__4319(mul_7_27_n_1044 ,mul_7_27_n_900 ,mul_7_27_n_1043);
  and mul_7_27_g2719__8428(mul_7_27_n_1043 ,mul_7_27_n_959 ,mul_7_27_n_1041);
  xnor mul_7_27_g2720__5526(out1[21] ,mul_7_27_n_1040 ,mul_7_27_n_967);
  or mul_7_27_g2721__6783(mul_7_27_n_1041 ,mul_7_27_n_960 ,mul_7_27_n_1040);
  and mul_7_27_g2722__3680(mul_7_27_n_1040 ,mul_7_27_n_962 ,mul_7_27_n_1038);
  xnor mul_7_27_g2723__1617(out1[20] ,mul_7_27_n_1037 ,mul_7_27_n_966);
  or mul_7_27_g2724__2802(mul_7_27_n_1038 ,mul_7_27_n_961 ,mul_7_27_n_1037);
  and mul_7_27_g2725__1705(mul_7_27_n_1037 ,mul_7_27_n_939 ,mul_7_27_n_1035);
  xnor mul_7_27_g2726__5122(out1[19] ,mul_7_27_n_1034 ,mul_7_27_n_968);
  or mul_7_27_g2727__8246(mul_7_27_n_1035 ,mul_7_27_n_958 ,mul_7_27_n_1034);
  and mul_7_27_g2728__7098(mul_7_27_n_1034 ,mul_7_27_n_975 ,mul_7_27_n_1032);
  xnor mul_7_27_g2729__6131(out1[18] ,mul_7_27_n_1031 ,mul_7_27_n_996);
  or mul_7_27_g2730__1881(mul_7_27_n_1032 ,mul_7_27_n_974 ,mul_7_27_n_1031);
  and mul_7_27_g2731__5115(mul_7_27_n_1031 ,mul_7_27_n_973 ,mul_7_27_n_1029);
  xnor mul_7_27_g2732__7482(out1[17] ,mul_7_27_n_1028 ,mul_7_27_n_995);
  or mul_7_27_g2733__4733(mul_7_27_n_1029 ,mul_7_27_n_972 ,mul_7_27_n_1028);
  and mul_7_27_g2734__6161(mul_7_27_n_1028 ,mul_7_27_n_985 ,mul_7_27_n_1026);
  xnor mul_7_27_g2735__9315(out1[16] ,mul_7_27_n_1025 ,mul_7_27_n_998);
  or mul_7_27_g2736__9945(mul_7_27_n_1026 ,mul_7_27_n_984 ,mul_7_27_n_1025);
  and mul_7_27_g2737__2883(mul_7_27_n_1025 ,mul_7_27_n_989 ,mul_7_27_n_1024);
  or mul_7_27_g2739__2346(mul_7_27_n_1024 ,mul_7_27_n_982 ,mul_7_27_n_1023);
  and mul_7_27_g2741__1666(mul_7_27_n_1023 ,mul_7_27_n_983 ,mul_7_27_n_1022);
  or mul_7_27_g2743__7410(mul_7_27_n_1022 ,mul_7_27_n_988 ,mul_7_27_n_1021);
  and mul_7_27_g2745__6417(mul_7_27_n_1021 ,mul_7_27_n_987 ,mul_7_27_n_1020);
  or mul_7_27_g2747__5477(mul_7_27_n_1020 ,mul_7_27_n_986 ,mul_7_27_n_1019);
  and mul_7_27_g2749__2398(mul_7_27_n_1019 ,mul_7_27_n_981 ,mul_7_27_n_1017);
  xnor mul_7_27_g2750__5107(out1[12] ,mul_7_27_n_1016 ,mul_7_27_n_994);
  or mul_7_27_g2751__6260(mul_7_27_n_1017 ,mul_7_27_n_980 ,mul_7_27_n_1016);
  and mul_7_27_g2752__4319(mul_7_27_n_1016 ,mul_7_27_n_955 ,mul_7_27_n_1014);
  xnor mul_7_27_g2753__8428(out1[11] ,mul_7_27_n_1013 ,mul_7_27_n_969);
  or mul_7_27_g2754__5526(mul_7_27_n_1014 ,mul_7_27_n_954 ,mul_7_27_n_1013);
  and mul_7_27_g2755__6783(mul_7_27_n_1013 ,mul_7_27_n_977 ,mul_7_27_n_1011);
  xnor mul_7_27_g2756__3680(out1[10] ,mul_7_27_n_1010 ,mul_7_27_n_997);
  or mul_7_27_g2757__1617(mul_7_27_n_1011 ,mul_7_27_n_976 ,mul_7_27_n_1010);
  and mul_7_27_g2758__2802(mul_7_27_n_1010 ,mul_7_27_n_979 ,mul_7_27_n_1008);
  xnor mul_7_27_g2759__1705(out1[9] ,mul_7_27_n_1007 ,mul_7_27_n_5);
  or mul_7_27_g2760__5122(mul_7_27_n_1008 ,mul_7_27_n_978 ,mul_7_27_n_1007);
  and mul_7_27_g2761__8246(mul_7_27_n_1007 ,mul_7_27_n_963 ,mul_7_27_n_1005);
  xnor mul_7_27_g2762__7098(out1[8] ,mul_7_27_n_1004 ,mul_7_27_n_970);
  or mul_7_27_g2763__6131(mul_7_27_n_1005 ,mul_7_27_n_957 ,mul_7_27_n_1004);
  and mul_7_27_g2764__1881(mul_7_27_n_1004 ,mul_7_27_n_924 ,mul_7_27_n_1002);
  xnor mul_7_27_g2765__5115(out1[7] ,mul_7_27_n_1001 ,mul_7_27_n_938);
  or mul_7_27_g2766__7482(mul_7_27_n_1002 ,mul_7_27_n_913 ,mul_7_27_n_1001);
  and mul_7_27_g2767__4733(mul_7_27_n_1001 ,mul_7_27_n_891 ,mul_7_27_n_999);
  xnor mul_7_27_g2768__6161(out1[6] ,mul_7_27_n_990 ,mul_7_27_n_911);
  or mul_7_27_g2769__9315(mul_7_27_n_999 ,mul_7_27_n_883 ,mul_7_27_n_990);
  xnor mul_7_27_g2770__9945(mul_7_27_n_998 ,mul_7_27_n_933 ,mul_7_27_n_947);
  xnor mul_7_27_g2771__2883(mul_7_27_n_997 ,mul_7_27_n_965 ,mul_7_27_n_951);
  xnor mul_7_27_g2772__2346(mul_7_27_n_996 ,mul_7_27_n_930 ,mul_7_27_n_949);
  xnor mul_7_27_g2773__1666(mul_7_27_n_995 ,mul_7_27_n_936 ,mul_7_27_n_953);
  xnor mul_7_27_g2774__7410(mul_7_27_n_994 ,mul_7_27_n_927 ,mul_7_27_n_942);
  xnor mul_7_27_g2776__6417(mul_7_27_n_993 ,mul_7_27_n_940 ,mul_7_27_n_931);
  xnor mul_7_27_g2777__5477(mul_7_27_n_992 ,mul_7_27_n_944 ,mul_7_27_n_934);
  xnor mul_7_27_g2778__2398(mul_7_27_n_991 ,mul_7_27_n_943 ,mul_7_27_n_928);
  or mul_7_27_g2779__5107(mul_7_27_n_989 ,mul_7_27_n_931 ,mul_7_27_n_940);
  and mul_7_27_g2780__6260(mul_7_27_n_988 ,mul_7_27_n_934 ,mul_7_27_n_944);
  or mul_7_27_g2781__4319(mul_7_27_n_987 ,mul_7_27_n_928 ,mul_7_27_n_943);
  and mul_7_27_g2782__8428(mul_7_27_n_986 ,mul_7_27_n_928 ,mul_7_27_n_943);
  or mul_7_27_g2783__5526(mul_7_27_n_985 ,mul_7_27_n_933 ,mul_7_27_n_946);
  nor mul_7_27_g2784__6783(mul_7_27_n_984 ,mul_7_27_n_932 ,mul_7_27_n_947);
  or mul_7_27_g2785__3680(mul_7_27_n_983 ,mul_7_27_n_934 ,mul_7_27_n_944);
  and mul_7_27_g2786__1617(mul_7_27_n_982 ,mul_7_27_n_931 ,mul_7_27_n_940);
  or mul_7_27_g2787__2802(mul_7_27_n_981 ,mul_7_27_n_926 ,mul_7_27_n_942);
  nor mul_7_27_g2788__1705(mul_7_27_n_980 ,mul_7_27_n_927 ,mul_7_27_n_941);
  or mul_7_27_g2789__5122(mul_7_27_n_979 ,mul_7_27_n_886 ,mul_7_27_n_945);
  and mul_7_27_g2790__8246(mul_7_27_n_990 ,mul_7_27_n_882 ,mul_7_27_n_956);
  and mul_7_27_g2791__7098(mul_7_27_n_978 ,mul_7_27_n_886 ,mul_7_27_n_945);
  or mul_7_27_g2792__6131(mul_7_27_n_977 ,mul_7_27_n_965 ,mul_7_27_n_950);
  nor mul_7_27_g2793__1881(mul_7_27_n_976 ,mul_7_27_n_964 ,mul_7_27_n_951);
  or mul_7_27_g2794__5115(mul_7_27_n_975 ,mul_7_27_n_930 ,mul_7_27_n_948);
  nor mul_7_27_g2795__7482(mul_7_27_n_974 ,mul_7_27_n_929 ,mul_7_27_n_949);
  or mul_7_27_g2796__4733(mul_7_27_n_973 ,mul_7_27_n_936 ,mul_7_27_n_952);
  nor mul_7_27_g2797__6161(mul_7_27_n_972 ,mul_7_27_n_935 ,mul_7_27_n_953);
  xnor mul_7_27_g2798__9315(out1[5] ,mul_7_27_n_937 ,mul_7_27_n_909);
  xnor mul_7_27_g2799__9945(mul_7_27_n_970 ,mul_7_27_n_904 ,mul_7_27_n_921);
  xnor mul_7_27_g2800__2883(mul_7_27_n_969 ,mul_7_27_n_885 ,mul_7_27_n_923);
  xnor mul_7_27_g2801__2346(mul_7_27_n_968 ,mul_7_27_n_906 ,mul_7_27_n_919);
  xnor mul_7_27_g2802__1666(mul_7_27_n_967 ,mul_7_27_n_908 ,mul_7_27_n_917);
  xnor mul_7_27_g2803__7410(mul_7_27_n_966 ,mul_7_27_n_902 ,mul_7_27_n_915);
  not mul_7_27_g2804(mul_7_27_n_964 ,mul_7_27_n_965);
  or mul_7_27_g2805__6417(mul_7_27_n_963 ,mul_7_27_n_904 ,mul_7_27_n_920);
  or mul_7_27_g2806__5477(mul_7_27_n_962 ,mul_7_27_n_902 ,mul_7_27_n_914);
  nor mul_7_27_g2807__2398(mul_7_27_n_961 ,mul_7_27_n_901 ,mul_7_27_n_915);
  nor mul_7_27_g2808__5107(mul_7_27_n_960 ,mul_7_27_n_907 ,mul_7_27_n_917);
  or mul_7_27_g2809__6260(mul_7_27_n_959 ,mul_7_27_n_908 ,mul_7_27_n_916);
  nor mul_7_27_g2810__4319(mul_7_27_n_958 ,mul_7_27_n_905 ,mul_7_27_n_919);
  nor mul_7_27_g2811__8428(mul_7_27_n_957 ,mul_7_27_n_903 ,mul_7_27_n_921);
  or mul_7_27_g2812__5526(mul_7_27_n_956 ,mul_7_27_n_881 ,mul_7_27_n_937);
  or mul_7_27_g2813__6783(mul_7_27_n_955 ,mul_7_27_n_885 ,mul_7_27_n_922);
  nor mul_7_27_g2814__3680(mul_7_27_n_954 ,mul_7_27_n_884 ,mul_7_27_n_923);
  and mul_7_27_g2815__1617(mul_7_27_n_965 ,mul_7_27_n_782 ,mul_7_27_n_925);
  not mul_7_27_g2816(mul_7_27_n_953 ,mul_7_27_n_952);
  not mul_7_27_g2817(mul_7_27_n_950 ,mul_7_27_n_951);
  not mul_7_27_g2818(mul_7_27_n_949 ,mul_7_27_n_948);
  not mul_7_27_g2819(mul_7_27_n_946 ,mul_7_27_n_947);
  not mul_7_27_g2821(mul_7_27_n_941 ,mul_7_27_n_942);
  or mul_7_27_g2822__2802(mul_7_27_n_939 ,mul_7_27_n_906 ,mul_7_27_n_918);
  xnor mul_7_27_g2823__1705(mul_7_27_n_938 ,mul_7_27_n_849 ,mul_7_27_n_887);
  xnor mul_7_27_g2824__5122(mul_7_27_n_952 ,mul_7_27_n_872 ,mul_7_27_n_877);
  xnor mul_7_27_g2825__8246(mul_7_27_n_951 ,mul_7_27_n_794 ,mul_7_27_n_874);
  xnor mul_7_27_g2826__7098(mul_7_27_n_948 ,mul_7_27_n_791 ,mul_7_27_n_4);
  xnor mul_7_27_g2827__6131(mul_7_27_n_947 ,mul_7_27_n_852 ,mul_7_27_n_875);
  xnor mul_7_27_g2828__1881(mul_7_27_n_945 ,mul_7_27_n_889 ,mul_7_27_n_799);
  xnor mul_7_27_g2829__5115(mul_7_27_n_944 ,mul_7_27_n_851 ,mul_7_27_n_879);
  xnor mul_7_27_g2830__7482(mul_7_27_n_943 ,mul_7_27_n_871 ,mul_7_27_n_873);
  xnor mul_7_27_g2831__4733(mul_7_27_n_942 ,mul_7_27_n_850 ,mul_7_27_n_880);
  xnor mul_7_27_g2832__6161(mul_7_27_n_940 ,mul_7_27_n_870 ,mul_7_27_n_878);
  not mul_7_27_g2833(mul_7_27_n_936 ,mul_7_27_n_935);
  not mul_7_27_g2834(mul_7_27_n_932 ,mul_7_27_n_933);
  not mul_7_27_g2835(mul_7_27_n_930 ,mul_7_27_n_929);
  not mul_7_27_g2836(mul_7_27_n_927 ,mul_7_27_n_926);
  or mul_7_27_g2837__9315(mul_7_27_n_925 ,mul_7_27_n_780 ,mul_7_27_n_889);
  or mul_7_27_g2838__9945(mul_7_27_n_924 ,mul_7_27_n_849 ,mul_7_27_n_888);
  and mul_7_27_g2839__2883(mul_7_27_n_937 ,mul_7_27_n_840 ,mul_7_27_n_890);
  or mul_7_27_g2840__2346(mul_7_27_n_935 ,mul_7_27_n_863 ,mul_7_27_n_897);
  and mul_7_27_g2841__1666(mul_7_27_n_934 ,mul_7_27_n_867 ,mul_7_27_n_893);
  and mul_7_27_g2842__7410(mul_7_27_n_933 ,mul_7_27_n_859 ,mul_7_27_n_896);
  and mul_7_27_g2843__6417(mul_7_27_n_931 ,mul_7_27_n_856 ,mul_7_27_n_895);
  or mul_7_27_g2844__5477(mul_7_27_n_929 ,mul_7_27_n_853 ,mul_7_27_n_892);
  and mul_7_27_g2845__2398(mul_7_27_n_928 ,mul_7_27_n_866 ,mul_7_27_n_899);
  and mul_7_27_g2846__5107(mul_7_27_n_926 ,mul_7_27_n_864 ,mul_7_27_n_898);
  not mul_7_27_g2847(mul_7_27_n_923 ,mul_7_27_n_922);
  not mul_7_27_g2848(mul_7_27_n_921 ,mul_7_27_n_920);
  not mul_7_27_g2849(mul_7_27_n_919 ,mul_7_27_n_918);
  not mul_7_27_g2850(mul_7_27_n_917 ,mul_7_27_n_916);
  not mul_7_27_g2851(mul_7_27_n_914 ,mul_7_27_n_915);
  and mul_7_27_g2852__6260(mul_7_27_n_913 ,mul_7_27_n_849 ,mul_7_27_n_888);
  xnor mul_7_27_g2853__4319(out1[4] ,mul_7_27_n_807 ,mul_7_27_n_836);
  xnor mul_7_27_g2854__8428(mul_7_27_n_911 ,mul_7_27_n_792 ,mul_7_27_n_845);
  xnor mul_7_27_g2855__5526(mul_7_27_n_910 ,mul_7_27_n_813 ,mul_7_27_n_869);
  xnor mul_7_27_g2856__6783(mul_7_27_n_909 ,mul_7_27_n_738 ,mul_7_27_n_848);
  xnor mul_7_27_g2857__3680(mul_7_27_n_922 ,mul_7_27_n_809 ,mul_7_27_n_833);
  xnor mul_7_27_g2858__1617(mul_7_27_n_920 ,mul_7_27_n_814 ,mul_7_27_n_832);
  xnor mul_7_27_g2859__2802(mul_7_27_n_918 ,mul_7_27_n_789 ,mul_7_27_n_834);
  xnor mul_7_27_g2860__1705(mul_7_27_n_916 ,mul_7_27_n_745 ,mul_7_27_n_1);
  xnor mul_7_27_g2861__5122(mul_7_27_n_915 ,mul_7_27_n_796 ,mul_7_27_n_835);
  not mul_7_27_g2862(mul_7_27_n_907 ,mul_7_27_n_908);
  not mul_7_27_g2863(mul_7_27_n_905 ,mul_7_27_n_906);
  not mul_7_27_g2864(mul_7_27_n_903 ,mul_7_27_n_904);
  not mul_7_27_g2865(mul_7_27_n_901 ,mul_7_27_n_902);
  and mul_7_27_g2866__8246(mul_7_27_n_900 ,mul_7_27_n_812 ,mul_7_27_n_869);
  or mul_7_27_g2867__7098(mul_7_27_n_899 ,mul_7_27_n_865 ,mul_7_27_n_850);
  or mul_7_27_g2868__6131(mul_7_27_n_898 ,mul_7_27_n_752 ,mul_7_27_n_862);
  and mul_7_27_g2869__1881(mul_7_27_n_897 ,mul_7_27_n_861 ,mul_7_27_n_852);
  or mul_7_27_g2870__5115(mul_7_27_n_896 ,mul_7_27_n_870 ,mul_7_27_n_858);
  or mul_7_27_g2871__7482(mul_7_27_n_895 ,mul_7_27_n_855 ,mul_7_27_n_851);
  and mul_7_27_g2872__4733(mul_7_27_n_894 ,mul_7_27_n_813 ,mul_7_27_n_868);
  or mul_7_27_g2873__6161(mul_7_27_n_893 ,mul_7_27_n_871 ,mul_7_27_n_857);
  and mul_7_27_g2874__9315(mul_7_27_n_892 ,mul_7_27_n_872 ,mul_7_27_n_854);
  or mul_7_27_g2875__9945(mul_7_27_n_891 ,mul_7_27_n_792 ,mul_7_27_n_846);
  or mul_7_27_g2876__2883(mul_7_27_n_890 ,mul_7_27_n_771 ,mul_7_27_n_839);
  and mul_7_27_g2877__2346(mul_7_27_n_908 ,mul_7_27_n_817 ,mul_7_27_n_844);
  and mul_7_27_g2878__1666(mul_7_27_n_906 ,mul_7_27_n_816 ,mul_7_27_n_842);
  and mul_7_27_g2879__7410(mul_7_27_n_904 ,mul_7_27_n_806 ,mul_7_27_n_843);
  and mul_7_27_g2880__6417(mul_7_27_n_902 ,mul_7_27_n_803 ,mul_7_27_n_860);
  not mul_7_27_g2881(mul_7_27_n_888 ,mul_7_27_n_887);
  not mul_7_27_g2882(mul_7_27_n_884 ,mul_7_27_n_885);
  and mul_7_27_g2883__5477(mul_7_27_n_883 ,mul_7_27_n_792 ,mul_7_27_n_846);
  or mul_7_27_g2884__2398(mul_7_27_n_882 ,mul_7_27_n_738 ,mul_7_27_n_847);
  nor mul_7_27_g2885__5107(mul_7_27_n_881 ,mul_7_27_n_737 ,mul_7_27_n_848);
  xnor mul_7_27_g2886__6260(mul_7_27_n_880 ,mul_7_27_n_829 ,mul_7_27_n_746);
  xnor mul_7_27_g2887__4319(mul_7_27_n_879 ,mul_7_27_n_828 ,mul_7_27_n_736);
  xnor mul_7_27_g2888__8428(mul_7_27_n_878 ,mul_7_27_n_808 ,mul_7_27_n_765);
  xnor mul_7_27_g2890__5526(mul_7_27_n_877 ,mul_7_27_n_719 ,mul_7_27_n_811);
  xnor mul_7_27_g2891__6783(mul_7_27_n_876 ,mul_7_27_n_756 ,mul_7_27_n_815);
  xnor mul_7_27_g2892__3680(mul_7_27_n_875 ,mul_7_27_n_827 ,mul_7_27_n_751);
  xnor mul_7_27_g2893__1617(mul_7_27_n_874 ,mul_7_27_n_830 ,mul_7_27_n_764);
  xnor mul_7_27_g2894__2802(mul_7_27_n_873 ,mul_7_27_n_810 ,mul_7_27_n_767);
  xnor mul_7_27_g2895__1705(mul_7_27_n_889 ,mul_7_27_n_543 ,mul_7_27_n_797);
  xnor mul_7_27_g2896__5122(mul_7_27_n_887 ,mul_7_27_n_762 ,mul_7_27_n_798);
  and mul_7_27_g2897__8246(mul_7_27_n_886 ,mul_7_27_n_800 ,mul_7_27_n_837);
  and mul_7_27_g2898__7098(mul_7_27_n_885 ,mul_7_27_n_821 ,mul_7_27_n_838);
  not mul_7_27_g2899(mul_7_27_n_868 ,mul_7_27_n_869);
  or mul_7_27_g2900__6131(mul_7_27_n_867 ,mul_7_27_n_767 ,mul_7_27_n_810);
  or mul_7_27_g2901__1881(mul_7_27_n_866 ,mul_7_27_n_746 ,mul_7_27_n_829);
  and mul_7_27_g2902__5115(mul_7_27_n_865 ,mul_7_27_n_746 ,mul_7_27_n_829);
  or mul_7_27_g2903__7482(mul_7_27_n_864 ,mul_7_27_n_769 ,mul_7_27_n_809);
  nor mul_7_27_g2904__4733(mul_7_27_n_863 ,mul_7_27_n_751 ,mul_7_27_n_827);
  and mul_7_27_g2905__6161(mul_7_27_n_862 ,mul_7_27_n_769 ,mul_7_27_n_809);
  or mul_7_27_g2906__9315(mul_7_27_n_861 ,mul_7_27_n_750 ,mul_7_27_n_826);
  or mul_7_27_g2907__9945(mul_7_27_n_860 ,mul_7_27_n_772 ,mul_7_27_n_802);
  or mul_7_27_g2908__2883(mul_7_27_n_859 ,mul_7_27_n_765 ,mul_7_27_n_808);
  and mul_7_27_g2909__2346(mul_7_27_n_858 ,mul_7_27_n_765 ,mul_7_27_n_808);
  and mul_7_27_g2910__1666(mul_7_27_n_857 ,mul_7_27_n_767 ,mul_7_27_n_810);
  or mul_7_27_g2911__7410(mul_7_27_n_856 ,mul_7_27_n_736 ,mul_7_27_n_828);
  and mul_7_27_g2912__6417(mul_7_27_n_855 ,mul_7_27_n_736 ,mul_7_27_n_828);
  or mul_7_27_g2913__5477(mul_7_27_n_854 ,mul_7_27_n_719 ,mul_7_27_n_3);
  nor mul_7_27_g2914__2398(mul_7_27_n_853 ,mul_7_27_n_718 ,mul_7_27_n_811);
  or mul_7_27_g2915__5107(mul_7_27_n_872 ,mul_7_27_n_660 ,mul_7_27_n_823);
  and mul_7_27_g2916__6260(mul_7_27_n_871 ,mul_7_27_n_666 ,mul_7_27_n_825);
  and mul_7_27_g2917__4319(mul_7_27_n_870 ,mul_7_27_n_626 ,mul_7_27_n_818);
  and mul_7_27_g2918__8428(mul_7_27_n_869 ,mul_7_27_n_787 ,mul_7_27_n_822);
  not mul_7_27_g2919(mul_7_27_n_847 ,mul_7_27_n_848);
  not mul_7_27_g2920(mul_7_27_n_846 ,mul_7_27_n_845);
  or mul_7_27_g2921__5526(mul_7_27_n_844 ,mul_7_27_n_796 ,mul_7_27_n_824);
  or mul_7_27_g2922__6783(mul_7_27_n_843 ,mul_7_27_n_740 ,mul_7_27_n_805);
  or mul_7_27_g2923__3680(mul_7_27_n_842 ,mul_7_27_n_831 ,mul_7_27_n_820);
  xnor mul_7_27_g2924__1617(out1[3] ,mul_7_27_n_722 ,mul_7_27_n_758);
  or mul_7_27_g2925__2802(mul_7_27_n_840 ,mul_7_27_n_639 ,mul_7_27_n_807);
  and mul_7_27_g2926__1705(mul_7_27_n_839 ,mul_7_27_n_639 ,mul_7_27_n_807);
  or mul_7_27_g2927__5122(mul_7_27_n_838 ,mul_7_27_n_830 ,mul_7_27_n_819);
  or mul_7_27_g2928__8246(mul_7_27_n_837 ,mul_7_27_n_814 ,mul_7_27_n_804);
  xnor mul_7_27_g2930__7098(mul_7_27_n_836 ,mul_7_27_n_638 ,mul_7_27_n_771);
  xnor mul_7_27_g2931__6131(mul_7_27_n_835 ,mul_7_27_n_748 ,mul_7_27_n_760);
  xnor mul_7_27_g2932__1881(mul_7_27_n_834 ,mul_7_27_n_768 ,mul_7_27_n_772);
  xnor mul_7_27_g2933__5115(mul_7_27_n_833 ,mul_7_27_n_769 ,mul_7_27_n_752);
  xnor mul_7_27_g2934__7482(mul_7_27_n_832 ,mul_7_27_n_795 ,mul_7_27_n_766);
  xnor mul_7_27_g2935__4733(mul_7_27_n_852 ,mul_7_27_n_770 ,mul_7_27_n_676);
  xnor mul_7_27_g2936__6161(mul_7_27_n_851 ,mul_7_27_n_776 ,mul_7_27_n_683);
  xnor mul_7_27_g2937__9315(mul_7_27_n_850 ,mul_7_27_n_775 ,mul_7_27_n_682);
  and mul_7_27_g2938__9945(mul_7_27_n_849 ,mul_7_27_n_699 ,mul_7_27_n_801);
  xnor mul_7_27_g2939__2883(mul_7_27_n_848 ,mul_7_27_n_536 ,mul_7_27_n_757);
  xnor mul_7_27_g2940__2346(mul_7_27_n_845 ,mul_7_27_n_773 ,mul_7_27_n_731);
  not mul_7_27_g2942(mul_7_27_n_826 ,mul_7_27_n_827);
  or mul_7_27_g2943__1666(mul_7_27_n_825 ,mul_7_27_n_654 ,mul_7_27_n_775);
  nor mul_7_27_g2944__7410(mul_7_27_n_824 ,mul_7_27_n_747 ,mul_7_27_n_760);
  and mul_7_27_g2945__6417(mul_7_27_n_823 ,mul_7_27_n_656 ,mul_7_27_n_770);
  or mul_7_27_g2946__5477(mul_7_27_n_822 ,mul_7_27_n_781 ,mul_7_27_n_774);
  or mul_7_27_g2947__2398(mul_7_27_n_821 ,mul_7_27_n_764 ,mul_7_27_n_793);
  nor mul_7_27_g2948__5107(mul_7_27_n_820 ,mul_7_27_n_716 ,mul_7_27_n_791);
  nor mul_7_27_g2949__6260(mul_7_27_n_819 ,mul_7_27_n_763 ,mul_7_27_n_794);
  or mul_7_27_g2950__4319(mul_7_27_n_818 ,mul_7_27_n_625 ,mul_7_27_n_776);
  or mul_7_27_g2951__8428(mul_7_27_n_817 ,mul_7_27_n_748 ,mul_7_27_n_759);
  or mul_7_27_g2952__5526(mul_7_27_n_816 ,mul_7_27_n_717 ,mul_7_27_n_790);
  nor mul_7_27_g2953__6783(mul_7_27_n_815 ,mul_7_27_n_608 ,mul_7_27_n_788);
  and mul_7_27_g2954__3680(mul_7_27_n_831 ,mul_7_27_n_617 ,mul_7_27_n_778);
  and mul_7_27_g2955__1617(mul_7_27_n_830 ,mul_7_27_n_643 ,mul_7_27_n_784);
  and mul_7_27_g2956__2802(mul_7_27_n_829 ,mul_7_27_n_661 ,mul_7_27_n_786);
  and mul_7_27_g2957__1705(mul_7_27_n_828 ,mul_7_27_n_670 ,mul_7_27_n_777);
  and mul_7_27_g2958__5122(mul_7_27_n_827 ,mul_7_27_n_644 ,mul_7_27_n_783);
  not mul_7_27_g2959(mul_7_27_n_812 ,mul_7_27_n_813);
  not mul_7_27_g2960(mul_7_27_n_811 ,mul_7_27_n_3);
  or mul_7_27_g2961__8246(mul_7_27_n_806 ,mul_7_27_n_539 ,mul_7_27_n_761);
  nor mul_7_27_g2962__7098(mul_7_27_n_805 ,mul_7_27_n_538 ,mul_7_27_n_762);
  and mul_7_27_g2963__6131(mul_7_27_n_804 ,mul_7_27_n_766 ,mul_7_27_n_795);
  or mul_7_27_g2964__1881(mul_7_27_n_803 ,mul_7_27_n_789 ,mul_7_27_n_768);
  and mul_7_27_g2965__5115(mul_7_27_n_802 ,mul_7_27_n_789 ,mul_7_27_n_768);
  or mul_7_27_g2966__7482(mul_7_27_n_801 ,mul_7_27_n_705 ,mul_7_27_n_773);
  or mul_7_27_g2967__4733(mul_7_27_n_800 ,mul_7_27_n_766 ,mul_7_27_n_795);
  xnor mul_7_27_g2968__6161(mul_7_27_n_799 ,mul_7_27_n_749 ,mul_7_27_n_697);
  xnor mul_7_27_g2969__9315(mul_7_27_n_798 ,mul_7_27_n_740 ,mul_7_27_n_539);
  xnor mul_7_27_g2970__9945(mul_7_27_n_797 ,mul_7_27_n_753 ,mul_7_27_n_582);
  xnor mul_7_27_g2971__2883(mul_7_27_n_814 ,mul_7_27_n_546 ,mul_7_27_n_730);
  xnor mul_7_27_g2972__2346(mul_7_27_n_813 ,mul_7_27_n_742 ,mul_7_27_n_0);
  xnor mul_7_27_g2974__1666(mul_7_27_n_810 ,mul_7_27_n_739 ,mul_7_27_n_684);
  xnor mul_7_27_g2975__7410(mul_7_27_n_809 ,mul_7_27_n_755 ,mul_7_27_n_681);
  xnor mul_7_27_g2976__6417(mul_7_27_n_808 ,mul_7_27_n_754 ,mul_7_27_n_675);
  and mul_7_27_g2977__5477(mul_7_27_n_807 ,mul_7_27_n_735 ,mul_7_27_n_779);
  not mul_7_27_g2978(mul_7_27_n_793 ,mul_7_27_n_794);
  not mul_7_27_g2979(mul_7_27_n_790 ,mul_7_27_n_791);
  nor mul_7_27_g2980__2398(mul_7_27_n_788 ,mul_7_27_n_609 ,mul_7_27_n_742);
  or mul_7_27_g2981__5107(mul_7_27_n_787 ,mul_7_27_n_87 ,mul_7_27_n_745);
  or mul_7_27_g2982__6260(mul_7_27_n_786 ,mul_7_27_n_659 ,mul_7_27_n_755);
  xnor mul_7_27_g2983__4319(out1[2] ,mul_7_27_n_698 ,mul_7_27_n_351);
  or mul_7_27_g2984__8428(mul_7_27_n_784 ,mul_7_27_n_641 ,mul_7_27_n_753);
  or mul_7_27_g2985__5526(mul_7_27_n_783 ,mul_7_27_n_646 ,mul_7_27_n_754);
  or mul_7_27_g2986__6783(mul_7_27_n_782 ,mul_7_27_n_697 ,mul_7_27_n_749);
  and mul_7_27_g2987__3680(mul_7_27_n_781 ,mul_7_27_n_89 ,mul_7_27_n_745);
  and mul_7_27_g2988__1617(mul_7_27_n_780 ,mul_7_27_n_697 ,mul_7_27_n_749);
  or mul_7_27_g2989__2802(mul_7_27_n_779 ,mul_7_27_n_722 ,mul_7_27_n_732);
  or mul_7_27_g2990__1705(mul_7_27_n_778 ,mul_7_27_n_665 ,mul_7_27_n_741);
  or mul_7_27_g2991__5122(mul_7_27_n_777 ,mul_7_27_n_651 ,mul_7_27_n_739);
  and mul_7_27_g2992__8246(mul_7_27_n_796 ,mul_7_27_n_667 ,mul_7_27_n_734);
  and mul_7_27_g2993__7098(mul_7_27_n_795 ,mul_7_27_n_633 ,mul_7_27_n_743);
  xnor mul_7_27_g2994__6131(mul_7_27_n_794 ,mul_7_27_n_671 ,mul_7_27_n_680);
  and mul_7_27_g2995__1881(mul_7_27_n_792 ,mul_7_27_n_635 ,mul_7_27_n_733);
  xnor mul_7_27_g2996__5115(mul_7_27_n_791 ,mul_7_27_n_727 ,mul_7_27_n_677);
  and mul_7_27_g2997__7482(mul_7_27_n_789 ,mul_7_27_n_649 ,mul_7_27_n_744);
  not mul_7_27_g2998(mul_7_27_n_763 ,mul_7_27_n_764);
  not mul_7_27_g2999(mul_7_27_n_761 ,mul_7_27_n_762);
  not mul_7_27_g3000(mul_7_27_n_759 ,mul_7_27_n_760);
  xnor mul_7_27_g3001__4733(mul_7_27_n_758 ,mul_7_27_n_549 ,mul_7_27_n_721);
  xnor mul_7_27_g3002__6161(mul_7_27_n_757 ,mul_7_27_n_552 ,mul_7_27_n_725);
  xnor mul_7_27_g3003__9315(mul_7_27_n_756 ,mul_7_27_n_674 ,mul_7_27_n_531);
  xnor mul_7_27_g3004__9945(mul_7_27_n_776 ,mul_7_27_n_599 ,mul_7_27_n_689);
  xnor mul_7_27_g3005__2883(mul_7_27_n_775 ,mul_7_27_n_555 ,mul_7_27_n_695);
  xnor mul_7_27_g3006__2346(mul_7_27_n_774 ,mul_7_27_n_678 ,mul_7_27_n_289);
  xnor mul_7_27_g3007__1666(mul_7_27_n_773 ,mul_7_27_n_571 ,mul_7_27_n_685);
  xnor mul_7_27_g3008__7410(mul_7_27_n_772 ,mul_7_27_n_532 ,mul_7_27_n_687);
  xnor mul_7_27_g3009__6417(mul_7_27_n_771 ,mul_7_27_n_534 ,mul_7_27_n_686);
  xnor mul_7_27_g3010__5477(mul_7_27_n_770 ,mul_7_27_n_597 ,mul_7_27_n_694);
  xnor mul_7_27_g3011__2398(mul_7_27_n_769 ,mul_7_27_n_604 ,mul_7_27_n_693);
  xnor mul_7_27_g3012__5107(mul_7_27_n_768 ,mul_7_27_n_729 ,mul_7_27_n_691);
  xnor mul_7_27_g3013__6260(mul_7_27_n_767 ,mul_7_27_n_554 ,mul_7_27_n_696);
  xnor mul_7_27_g3014__4319(mul_7_27_n_766 ,mul_7_27_n_589 ,mul_7_27_n_2);
  xnor mul_7_27_g3015__8428(mul_7_27_n_765 ,mul_7_27_n_563 ,mul_7_27_n_690);
  xnor mul_7_27_g3016__5526(mul_7_27_n_764 ,mul_7_27_n_606 ,mul_7_27_n_692);
  xnor mul_7_27_g3017__6783(mul_7_27_n_762 ,mul_7_27_n_723 ,mul_7_27_n_673);
  xnor mul_7_27_g3018__3680(mul_7_27_n_760 ,mul_7_27_n_688 ,mul_7_27_n_529);
  not mul_7_27_g3019(mul_7_27_n_750 ,mul_7_27_n_751);
  not mul_7_27_g3020(mul_7_27_n_747 ,mul_7_27_n_748);
  or mul_7_27_g3021__1617(mul_7_27_n_744 ,mul_7_27_n_642 ,mul_7_27_n_728);
  or mul_7_27_g3022__2802(mul_7_27_n_743 ,mul_7_27_n_627 ,mul_7_27_n_724);
  and mul_7_27_g3023__1705(mul_7_27_n_755 ,mul_7_27_n_658 ,mul_7_27_n_713);
  and mul_7_27_g3024__5122(mul_7_27_n_754 ,mul_7_27_n_619 ,mul_7_27_n_707);
  and mul_7_27_g3025__8246(mul_7_27_n_753 ,mul_7_27_n_664 ,mul_7_27_n_708);
  and mul_7_27_g3026__7098(mul_7_27_n_752 ,mul_7_27_n_650 ,mul_7_27_n_711);
  and mul_7_27_g3027__6131(mul_7_27_n_751 ,mul_7_27_n_648 ,mul_7_27_n_710);
  and mul_7_27_g3028__1881(mul_7_27_n_749 ,mul_7_27_n_632 ,mul_7_27_n_706);
  and mul_7_27_g3029__5115(mul_7_27_n_748 ,mul_7_27_n_629 ,mul_7_27_n_703);
  and mul_7_27_g3030__7482(mul_7_27_n_746 ,mul_7_27_n_663 ,mul_7_27_n_714);
  and mul_7_27_g3031__4733(mul_7_27_n_745 ,mul_7_27_n_610 ,mul_7_27_n_709);
  not mul_7_27_g3033(mul_7_27_n_737 ,mul_7_27_n_738);
  or mul_7_27_g3034__6161(mul_7_27_n_735 ,mul_7_27_n_549 ,mul_7_27_n_720);
  or mul_7_27_g3035__9315(mul_7_27_n_734 ,mul_7_27_n_669 ,mul_7_27_n_729);
  or mul_7_27_g3036__9945(mul_7_27_n_733 ,mul_7_27_n_652 ,mul_7_27_n_726);
  nor mul_7_27_g3037__2883(mul_7_27_n_732 ,mul_7_27_n_548 ,mul_7_27_n_721);
  xnor mul_7_27_g3038__2346(mul_7_27_n_731 ,mul_7_27_n_542 ,mul_7_27_n_637);
  xnor mul_7_27_g3039__1666(mul_7_27_n_730 ,mul_7_27_n_579 ,mul_7_27_n_640);
  and mul_7_27_g3040__7410(mul_7_27_n_742 ,mul_7_27_n_655 ,mul_7_27_n_712);
  and mul_7_27_g3041__6417(mul_7_27_n_741 ,mul_7_27_n_613 ,mul_7_27_n_702);
  and mul_7_27_g3042__5477(mul_7_27_n_740 ,mul_7_27_n_624 ,mul_7_27_n_704);
  and mul_7_27_g3043__2398(mul_7_27_n_739 ,mul_7_27_n_653 ,mul_7_27_n_700);
  and mul_7_27_g3044__5107(mul_7_27_n_738 ,mul_7_27_n_616 ,mul_7_27_n_701);
  and mul_7_27_g3045__6260(mul_7_27_n_736 ,mul_7_27_n_620 ,mul_7_27_n_715);
  not mul_7_27_g3046(mul_7_27_n_728 ,mul_7_27_n_727);
  not mul_7_27_g3047(mul_7_27_n_726 ,mul_7_27_n_725);
  not mul_7_27_g3048(mul_7_27_n_724 ,mul_7_27_n_723);
  not mul_7_27_g3049(mul_7_27_n_720 ,mul_7_27_n_721);
  not mul_7_27_g3050(mul_7_27_n_718 ,mul_7_27_n_719);
  not mul_7_27_g3051(mul_7_27_n_716 ,mul_7_27_n_717);
  or mul_7_27_g3052__4319(mul_7_27_n_715 ,mul_7_27_n_554 ,mul_7_27_n_618);
  or mul_7_27_g3053__8428(mul_7_27_n_714 ,mul_7_27_n_604 ,mul_7_27_n_662);
  or mul_7_27_g3054__5526(mul_7_27_n_713 ,mul_7_27_n_606 ,mul_7_27_n_657);
  or mul_7_27_g3055__6783(mul_7_27_n_712 ,mul_7_27_n_605 ,mul_7_27_n_628);
  or mul_7_27_g3056__3680(mul_7_27_n_711 ,mul_7_27_n_647 ,mul_7_27_n_672);
  or mul_7_27_g3057__1617(mul_7_27_n_710 ,mul_7_27_n_563 ,mul_7_27_n_645);
  or mul_7_27_g3058__2802(mul_7_27_n_709 ,mul_7_27_n_607 ,mul_7_27_n_603);
  or mul_7_27_g3059__1705(mul_7_27_n_708 ,mul_7_27_n_569 ,mul_7_27_n_634);
  or mul_7_27_g3060__5122(mul_7_27_n_707 ,mul_7_27_n_599 ,mul_7_27_n_631);
  or mul_7_27_g3061__8246(mul_7_27_n_706 ,mul_7_27_n_640 ,mul_7_27_n_630);
  nor mul_7_27_g3062__7098(mul_7_27_n_705 ,mul_7_27_n_541 ,mul_7_27_n_637);
  or mul_7_27_g3063__6131(mul_7_27_n_704 ,mul_7_27_n_600 ,mul_7_27_n_622);
  or mul_7_27_g3064__1881(mul_7_27_n_703 ,mul_7_27_n_596 ,mul_7_27_n_614);
  or mul_7_27_g3065__5115(mul_7_27_n_702 ,mul_7_27_n_598 ,mul_7_27_n_668);
  or mul_7_27_g3066__7482(mul_7_27_n_701 ,mul_7_27_n_561 ,mul_7_27_n_615);
  or mul_7_27_g3067__4733(mul_7_27_n_700 ,mul_7_27_n_555 ,mul_7_27_n_611);
  or mul_7_27_g3068__6161(mul_7_27_n_699 ,mul_7_27_n_542 ,mul_7_27_n_636);
  xnor mul_7_27_g3069__9315(mul_7_27_n_698 ,mul_7_27_n_408 ,mul_7_27_n_566);
  and mul_7_27_g3070__9945(mul_7_27_n_729 ,mul_7_27_n_346 ,mul_7_27_n_621);
  xnor mul_7_27_g3071__2883(mul_7_27_n_727 ,mul_7_27_n_556 ,mul_7_27_n_378);
  xnor mul_7_27_g3072__2346(mul_7_27_n_725 ,mul_7_27_n_487 ,mul_7_27_n_564);
  xnor mul_7_27_g3073__1666(mul_7_27_n_723 ,mul_7_27_n_485 ,mul_7_27_n_568);
  and mul_7_27_g3074__7410(mul_7_27_n_722 ,mul_7_27_n_497 ,mul_7_27_n_612);
  xnor mul_7_27_g3075__6417(mul_7_27_n_721 ,mul_7_27_n_488 ,mul_7_27_n_557);
  xnor mul_7_27_g3076__5477(mul_7_27_n_719 ,mul_7_27_n_562 ,mul_7_27_n_379);
  and mul_7_27_g3077__2398(mul_7_27_n_717 ,mul_7_27_n_345 ,mul_7_27_n_623);
  xnor mul_7_27_g3079__5107(mul_7_27_n_696 ,mul_7_27_n_550 ,mul_7_27_n_293);
  xnor mul_7_27_g3080__6260(mul_7_27_n_695 ,mul_7_27_n_551 ,mul_7_27_n_288);
  xnor mul_7_27_g3081__4319(mul_7_27_n_694 ,mul_7_27_n_584 ,mul_7_27_n_287);
  xnor mul_7_27_g3082__8428(mul_7_27_n_693 ,mul_7_27_n_592 ,mul_7_27_n_291);
  xnor mul_7_27_g3083__5526(mul_7_27_n_692 ,mul_7_27_n_580 ,mul_7_27_n_295);
  xnor mul_7_27_g3084__6783(mul_7_27_n_691 ,mul_7_27_n_576 ,mul_7_27_n_276);
  xnor mul_7_27_g3085__3680(mul_7_27_n_690 ,mul_7_27_n_553 ,mul_7_27_n_290);
  xnor mul_7_27_g3086__1617(mul_7_27_n_689 ,mul_7_27_n_533 ,mul_7_27_n_292);
  xnor mul_7_27_g3087__2802(mul_7_27_n_688 ,mul_7_27_n_603 ,mul_7_27_n_274);
  xnor mul_7_27_g3089__1705(mul_7_27_n_687 ,mul_7_27_n_596 ,in1[1]);
  xnor mul_7_27_g3090__5122(mul_7_27_n_686 ,mul_7_27_n_561 ,mul_7_27_n_410);
  xnor mul_7_27_g3091__8246(mul_7_27_n_685 ,mul_7_27_n_600 ,mul_7_27_n_409);
  xnor mul_7_27_g3092__7098(mul_7_27_n_684 ,mul_7_27_n_573 ,mul_7_27_n_535);
  xnor mul_7_27_g3093__6131(mul_7_27_n_683 ,mul_7_27_n_572 ,mul_7_27_n_540);
  xnor mul_7_27_g3094__1881(mul_7_27_n_682 ,mul_7_27_n_581 ,mul_7_27_n_537);
  xnor mul_7_27_g3095__5115(mul_7_27_n_681 ,mul_7_27_n_585 ,mul_7_27_n_547);
  xnor mul_7_27_g3096__7482(mul_7_27_n_680 ,mul_7_27_n_591 ,mul_7_27_n_545);
  xnor mul_7_27_g3097__4733(mul_7_27_n_679 ,mul_7_27_n_544 ,mul_7_27_n_594);
  xnor mul_7_27_g3098__6161(mul_7_27_n_678 ,mul_7_27_n_595 ,mul_7_27_n_605);
  xnor mul_7_27_g3099__9315(mul_7_27_n_677 ,mul_7_27_n_586 ,mul_7_27_n_590);
  xnor mul_7_27_g3100__9945(mul_7_27_n_676 ,mul_7_27_n_578 ,mul_7_27_n_588);
  xnor mul_7_27_g3101__2883(mul_7_27_n_675 ,mul_7_27_n_583 ,mul_7_27_n_575);
  xnor mul_7_27_g3102__2346(mul_7_27_n_674 ,mul_7_27_n_258 ,mul_7_27_n_570);
  xnor mul_7_27_g3103__1666(mul_7_27_n_673 ,mul_7_27_n_574 ,mul_7_27_n_593);
  xnor mul_7_27_g3104__7410(mul_7_27_n_697 ,mul_7_27_n_601 ,mul_7_27_n_559);
  not mul_7_27_g3105(mul_7_27_n_672 ,mul_7_27_n_671);
  or mul_7_27_g3106__6417(mul_7_27_n_670 ,mul_7_27_n_535 ,mul_7_27_n_573);
  and mul_7_27_g3107__5477(mul_7_27_n_669 ,mul_7_27_n_174 ,mul_7_27_n_576);
  and mul_7_27_g3108__2398(mul_7_27_n_668 ,mul_7_27_n_175 ,mul_7_27_n_584);
  or mul_7_27_g3109__5107(mul_7_27_n_667 ,mul_7_27_n_276 ,mul_7_27_n_576);
  or mul_7_27_g3110__6260(mul_7_27_n_666 ,mul_7_27_n_537 ,mul_7_27_n_581);
  and mul_7_27_g3111__4319(mul_7_27_n_665 ,mul_7_27_n_594 ,mul_7_27_n_544);
  or mul_7_27_g3112__8428(mul_7_27_n_664 ,mul_7_27_n_162 ,mul_7_27_n_589);
  or mul_7_27_g3113__5526(mul_7_27_n_663 ,mul_7_27_n_168 ,mul_7_27_n_592);
  and mul_7_27_g3114__6783(mul_7_27_n_662 ,mul_7_27_n_291 ,mul_7_27_n_592);
  or mul_7_27_g3115__3680(mul_7_27_n_661 ,mul_7_27_n_547 ,mul_7_27_n_585);
  nor mul_7_27_g3116__1617(mul_7_27_n_660 ,mul_7_27_n_588 ,mul_7_27_n_578);
  and mul_7_27_g3117__2802(mul_7_27_n_659 ,mul_7_27_n_547 ,mul_7_27_n_585);
  or mul_7_27_g3118__1705(mul_7_27_n_658 ,mul_7_27_n_173 ,mul_7_27_n_580);
  and mul_7_27_g3119__5122(mul_7_27_n_657 ,mul_7_27_n_295 ,mul_7_27_n_580);
  or mul_7_27_g3120__8246(mul_7_27_n_656 ,mul_7_27_n_587 ,mul_7_27_n_577);
  or mul_7_27_g3121__7098(mul_7_27_n_655 ,mul_7_27_n_167 ,mul_7_27_n_595);
  and mul_7_27_g3122__6131(mul_7_27_n_654 ,mul_7_27_n_537 ,mul_7_27_n_581);
  or mul_7_27_g3123__1881(mul_7_27_n_653 ,mul_7_27_n_169 ,mul_7_27_n_551);
  and mul_7_27_g3124__5115(mul_7_27_n_652 ,mul_7_27_n_536 ,mul_7_27_n_552);
  and mul_7_27_g3125__7482(mul_7_27_n_651 ,mul_7_27_n_535 ,mul_7_27_n_573);
  or mul_7_27_g3126__4733(mul_7_27_n_650 ,mul_7_27_n_545 ,mul_7_27_n_591);
  or mul_7_27_g3127__6161(mul_7_27_n_649 ,mul_7_27_n_590 ,mul_7_27_n_586);
  or mul_7_27_g3128__9315(mul_7_27_n_648 ,mul_7_27_n_171 ,mul_7_27_n_553);
  and mul_7_27_g3129__9945(mul_7_27_n_647 ,mul_7_27_n_545 ,mul_7_27_n_591);
  and mul_7_27_g3130__2883(mul_7_27_n_646 ,mul_7_27_n_575 ,mul_7_27_n_583);
  and mul_7_27_g3131__2346(mul_7_27_n_645 ,mul_7_27_n_290 ,mul_7_27_n_553);
  or mul_7_27_g3132__1666(mul_7_27_n_644 ,mul_7_27_n_575 ,mul_7_27_n_583);
  or mul_7_27_g3133__7410(mul_7_27_n_643 ,mul_7_27_n_543 ,mul_7_27_n_582);
  and mul_7_27_g3134__6417(mul_7_27_n_642 ,mul_7_27_n_590 ,mul_7_27_n_586);
  and mul_7_27_g3135__5477(mul_7_27_n_641 ,mul_7_27_n_543 ,mul_7_27_n_582);
  and mul_7_27_g3136__2398(mul_7_27_n_671 ,mul_7_27_n_560 ,mul_7_27_n_602);
  not mul_7_27_g3137(mul_7_27_n_639 ,mul_7_27_n_638);
  not mul_7_27_g3138(mul_7_27_n_636 ,mul_7_27_n_637);
  or mul_7_27_g3139__5107(mul_7_27_n_635 ,mul_7_27_n_536 ,mul_7_27_n_552);
  and mul_7_27_g3140__6260(mul_7_27_n_634 ,mul_7_27_n_162 ,mul_7_27_n_589);
  or mul_7_27_g3141__4319(mul_7_27_n_633 ,mul_7_27_n_593 ,mul_7_27_n_574);
  or mul_7_27_g3142__8428(mul_7_27_n_632 ,mul_7_27_n_546 ,mul_7_27_n_579);
  and mul_7_27_g3143__5526(mul_7_27_n_631 ,mul_7_27_n_172 ,mul_7_27_n_533);
  and mul_7_27_g3144__6783(mul_7_27_n_630 ,mul_7_27_n_546 ,mul_7_27_n_579);
  or mul_7_27_g3145__3680(mul_7_27_n_629 ,in1[1] ,mul_7_27_n_532);
  and mul_7_27_g3146__1617(mul_7_27_n_628 ,mul_7_27_n_289 ,mul_7_27_n_595);
  and mul_7_27_g3147__2802(mul_7_27_n_627 ,mul_7_27_n_593 ,mul_7_27_n_574);
  or mul_7_27_g3148__1705(mul_7_27_n_626 ,mul_7_27_n_540 ,mul_7_27_n_572);
  and mul_7_27_g3149__5122(mul_7_27_n_625 ,mul_7_27_n_540 ,mul_7_27_n_572);
  or mul_7_27_g3150__8246(mul_7_27_n_624 ,mul_7_27_n_409 ,mul_7_27_n_571);
  or mul_7_27_g3151__7098(mul_7_27_n_623 ,mul_7_27_n_343 ,mul_7_27_n_562);
  and mul_7_27_g3152__6131(mul_7_27_n_622 ,mul_7_27_n_409 ,mul_7_27_n_571);
  or mul_7_27_g3153__1881(mul_7_27_n_621 ,mul_7_27_n_344 ,mul_7_27_n_556);
  or mul_7_27_g3154__5115(mul_7_27_n_620 ,mul_7_27_n_170 ,mul_7_27_n_550);
  or mul_7_27_g3155__7482(mul_7_27_n_619 ,mul_7_27_n_292 ,mul_7_27_n_533);
  and mul_7_27_g3156__4733(mul_7_27_n_618 ,mul_7_27_n_293 ,mul_7_27_n_550);
  or mul_7_27_g3157__6161(mul_7_27_n_617 ,mul_7_27_n_594 ,mul_7_27_n_544);
  or mul_7_27_g3158__9315(mul_7_27_n_616 ,mul_7_27_n_410 ,mul_7_27_n_534);
  and mul_7_27_g3159__9945(mul_7_27_n_615 ,mul_7_27_n_410 ,mul_7_27_n_534);
  and mul_7_27_g3160__2883(mul_7_27_n_614 ,in1[1] ,mul_7_27_n_532);
  or mul_7_27_g3161__2346(mul_7_27_n_613 ,mul_7_27_n_287 ,mul_7_27_n_584);
  or mul_7_27_g3162__1666(mul_7_27_n_612 ,mul_7_27_n_498 ,mul_7_27_n_567);
  and mul_7_27_g3163__7410(mul_7_27_n_611 ,mul_7_27_n_288 ,mul_7_27_n_551);
  or mul_7_27_g3164__6417(mul_7_27_n_610 ,mul_7_27_n_274 ,mul_7_27_n_530);
  and mul_7_27_g3165__5477(mul_7_27_n_609 ,mul_7_27_n_294 ,mul_7_27_n_177);
  nor mul_7_27_g3166__2398(mul_7_27_n_608 ,mul_7_27_n_294 ,mul_7_27_n_177);
  nor mul_7_27_g3167__5107(mul_7_27_n_607 ,mul_7_27_n_273 ,mul_7_27_n_89);
  or mul_7_27_g3168__6260(mul_7_27_n_640 ,mul_7_27_n_486 ,mul_7_27_n_568);
  and mul_7_27_g3169__4319(mul_7_27_n_638 ,mul_7_27_n_488 ,mul_7_27_n_558);
  and mul_7_27_g3170__8428(mul_7_27_n_637 ,mul_7_27_n_487 ,mul_7_27_n_565);
  not mul_7_27_g3171(mul_7_27_n_602 ,mul_7_27_n_601);
  not mul_7_27_g3172(mul_7_27_n_598 ,mul_7_27_n_597);
  not mul_7_27_g3173(mul_7_27_n_587 ,mul_7_27_n_588);
  not mul_7_27_g3174(mul_7_27_n_577 ,mul_7_27_n_578);
  or mul_7_27_g3175__5526(mul_7_27_n_570 ,mul_7_27_n_416 ,mul_7_27_n_490);
  and mul_7_27_g3176__6783(mul_7_27_n_606 ,mul_7_27_n_431 ,mul_7_27_n_518);
  or mul_7_27_g3177__3680(mul_7_27_n_605 ,mul_7_27_n_413 ,mul_7_27_n_493);
  and mul_7_27_g3178__1617(mul_7_27_n_604 ,mul_7_27_n_445 ,mul_7_27_n_524);
  and mul_7_27_g3179__2802(mul_7_27_n_603 ,mul_7_27_n_388 ,mul_7_27_n_462);
  and mul_7_27_g3180__1705(mul_7_27_n_601 ,mul_7_27_n_385 ,mul_7_27_n_467);
  and mul_7_27_g3181__5122(mul_7_27_n_600 ,mul_7_27_n_432 ,mul_7_27_n_494);
  and mul_7_27_g3182__8246(mul_7_27_n_599 ,mul_7_27_n_434 ,mul_7_27_n_516);
  or mul_7_27_g3183__7098(mul_7_27_n_597 ,mul_7_27_n_282 ,mul_7_27_n_479);
  or mul_7_27_g3184__6131(mul_7_27_n_596 ,mul_7_27_n_411 ,mul_7_27_n_491);
  and mul_7_27_g3185__1881(mul_7_27_n_595 ,mul_7_27_n_407 ,mul_7_27_n_463);
  and mul_7_27_g3186__5115(mul_7_27_n_594 ,mul_7_27_n_426 ,mul_7_27_n_502);
  and mul_7_27_g3187__7482(mul_7_27_n_593 ,mul_7_27_n_430 ,mul_7_27_n_507);
  and mul_7_27_g3188__4733(mul_7_27_n_592 ,mul_7_27_n_391 ,mul_7_27_n_461);
  and mul_7_27_g3189__6161(mul_7_27_n_591 ,mul_7_27_n_419 ,mul_7_27_n_515);
  and mul_7_27_g3190__9315(mul_7_27_n_590 ,mul_7_27_n_438 ,mul_7_27_n_513);
  and mul_7_27_g3191__9945(mul_7_27_n_589 ,mul_7_27_n_420 ,mul_7_27_n_509);
  and mul_7_27_g3192__2883(mul_7_27_n_588 ,mul_7_27_n_447 ,mul_7_27_n_520);
  and mul_7_27_g3193__2346(mul_7_27_n_586 ,mul_7_27_n_390 ,mul_7_27_n_458);
  and mul_7_27_g3194__1666(mul_7_27_n_585 ,mul_7_27_n_446 ,mul_7_27_n_521);
  and mul_7_27_g3195__7410(mul_7_27_n_584 ,mul_7_27_n_387 ,mul_7_27_n_472);
  and mul_7_27_g3196__6417(mul_7_27_n_583 ,mul_7_27_n_437 ,mul_7_27_n_511);
  and mul_7_27_g3197__5477(mul_7_27_n_582 ,mul_7_27_n_429 ,mul_7_27_n_510);
  and mul_7_27_g3198__2398(mul_7_27_n_581 ,mul_7_27_n_443 ,mul_7_27_n_526);
  and mul_7_27_g3199__5107(mul_7_27_n_580 ,mul_7_27_n_392 ,mul_7_27_n_459);
  and mul_7_27_g3200__6260(mul_7_27_n_579 ,mul_7_27_n_428 ,mul_7_27_n_527);
  and mul_7_27_g3201__4319(mul_7_27_n_578 ,mul_7_27_n_440 ,mul_7_27_n_519);
  and mul_7_27_g3202__8428(mul_7_27_n_576 ,mul_7_27_n_393 ,mul_7_27_n_460);
  and mul_7_27_g3203__5526(mul_7_27_n_575 ,mul_7_27_n_435 ,mul_7_27_n_512);
  and mul_7_27_g3204__6783(mul_7_27_n_574 ,mul_7_27_n_439 ,mul_7_27_n_517);
  and mul_7_27_g3205__3680(mul_7_27_n_573 ,mul_7_27_n_418 ,mul_7_27_n_500);
  and mul_7_27_g3206__1617(mul_7_27_n_572 ,mul_7_27_n_436 ,mul_7_27_n_499);
  and mul_7_27_g3207__2802(mul_7_27_n_571 ,mul_7_27_n_448 ,mul_7_27_n_501);
  not mul_7_27_g3208(mul_7_27_n_567 ,mul_7_27_n_566);
  not mul_7_27_g3209(mul_7_27_n_565 ,mul_7_27_n_564);
  not mul_7_27_g3210(mul_7_27_n_560 ,mul_7_27_n_559);
  not mul_7_27_g3211(mul_7_27_n_558 ,mul_7_27_n_557);
  not mul_7_27_g3212(mul_7_27_n_548 ,mul_7_27_n_549);
  not mul_7_27_g3213(mul_7_27_n_541 ,mul_7_27_n_542);
  not mul_7_27_g3214(mul_7_27_n_538 ,mul_7_27_n_539);
  not mul_7_27_g3215(mul_7_27_n_530 ,mul_7_27_n_87);
  and mul_7_27_g3216__1705(mul_7_27_n_569 ,mul_7_27_n_386 ,mul_7_27_n_489);
  and mul_7_27_g3217__5122(mul_7_27_n_568 ,mul_7_27_n_415 ,mul_7_27_n_465);
  or mul_7_27_g3218__8246(mul_7_27_n_566 ,mul_7_27_n_395 ,mul_7_27_n_466);
  and mul_7_27_g3219__7098(mul_7_27_n_564 ,mul_7_27_n_441 ,mul_7_27_n_504);
  and mul_7_27_g3220__6131(mul_7_27_n_563 ,mul_7_27_n_402 ,mul_7_27_n_482);
  and mul_7_27_g3221__1881(mul_7_27_n_562 ,mul_7_27_n_422 ,mul_7_27_n_505);
  and mul_7_27_g3222__5115(mul_7_27_n_561 ,mul_7_27_n_423 ,mul_7_27_n_492);
  and mul_7_27_g3223__7482(mul_7_27_n_559 ,mul_7_27_n_424 ,mul_7_27_n_514);
  and mul_7_27_g3224__4733(mul_7_27_n_557 ,mul_7_27_n_412 ,mul_7_27_n_528);
  and mul_7_27_g3225__6161(mul_7_27_n_556 ,mul_7_27_n_412 ,mul_7_27_n_522);
  and mul_7_27_g3226__9315(mul_7_27_n_555 ,mul_7_27_n_421 ,mul_7_27_n_525);
  and mul_7_27_g3227__9945(mul_7_27_n_554 ,mul_7_27_n_442 ,mul_7_27_n_506);
  and mul_7_27_g3228__2883(mul_7_27_n_553 ,mul_7_27_n_383 ,mul_7_27_n_457);
  and mul_7_27_g3229__2346(mul_7_27_n_552 ,mul_7_27_n_414 ,mul_7_27_n_503);
  and mul_7_27_g3230__1666(mul_7_27_n_551 ,mul_7_27_n_381 ,mul_7_27_n_470);
  and mul_7_27_g3231__7410(mul_7_27_n_550 ,mul_7_27_n_394 ,mul_7_27_n_471);
  and mul_7_27_g3232__6417(mul_7_27_n_549 ,mul_7_27_n_401 ,mul_7_27_n_474);
  and mul_7_27_g3233__5477(mul_7_27_n_547 ,mul_7_27_n_404 ,mul_7_27_n_484);
  and mul_7_27_g3234__2398(mul_7_27_n_546 ,mul_7_27_n_389 ,mul_7_27_n_480);
  and mul_7_27_g3235__5107(mul_7_27_n_545 ,mul_7_27_n_403 ,mul_7_27_n_483);
  and mul_7_27_g3236__6260(mul_7_27_n_544 ,mul_7_27_n_382 ,mul_7_27_n_468);
  and mul_7_27_g3237__4319(mul_7_27_n_543 ,mul_7_27_n_444 ,mul_7_27_n_481);
  and mul_7_27_g3238__8428(mul_7_27_n_542 ,mul_7_27_n_405 ,mul_7_27_n_475);
  and mul_7_27_g3239__5526(mul_7_27_n_540 ,mul_7_27_n_400 ,mul_7_27_n_477);
  and mul_7_27_g3240__6783(mul_7_27_n_539 ,mul_7_27_n_399 ,mul_7_27_n_476);
  and mul_7_27_g3241__3680(mul_7_27_n_537 ,mul_7_27_n_397 ,mul_7_27_n_496);
  and mul_7_27_g3242__1617(mul_7_27_n_536 ,mul_7_27_n_396 ,mul_7_27_n_495);
  and mul_7_27_g3243__2802(mul_7_27_n_535 ,mul_7_27_n_398 ,mul_7_27_n_478);
  and mul_7_27_g3244__1705(mul_7_27_n_534 ,mul_7_27_n_406 ,mul_7_27_n_473);
  and mul_7_27_g3245__5122(mul_7_27_n_533 ,mul_7_27_n_384 ,mul_7_27_n_469);
  and mul_7_27_g3246__8246(mul_7_27_n_532 ,mul_7_27_n_425 ,mul_7_27_n_508);
  or mul_7_27_g3247__7098(mul_7_27_n_531 ,mul_7_27_n_416 ,mul_7_27_n_464);
  and mul_7_27_g3248__6131(mul_7_27_n_529 ,mul_7_27_n_414 ,mul_7_27_n_523);
  or mul_7_27_g3249__1881(mul_7_27_n_528 ,mul_7_27_n_297 ,mul_7_27_n_117);
  or mul_7_27_g3250__5115(mul_7_27_n_527 ,mul_7_27_n_340 ,mul_7_27_n_117);
  or mul_7_27_g3251__7482(mul_7_27_n_526 ,mul_7_27_n_322 ,mul_7_27_n_68);
  or mul_7_27_g3252__4733(mul_7_27_n_525 ,mul_7_27_n_324 ,mul_7_27_n_99);
  or mul_7_27_g3253__6161(mul_7_27_n_524 ,mul_7_27_n_338 ,mul_7_27_n_99);
  or mul_7_27_g3254__9315(mul_7_27_n_523 ,mul_7_27_n_328 ,mul_7_27_n_71);
  or mul_7_27_g3255__9945(mul_7_27_n_522 ,mul_7_27_n_332 ,mul_7_27_n_97);
  or mul_7_27_g3256__2883(mul_7_27_n_521 ,mul_7_27_n_318 ,mul_7_27_n_69);
  or mul_7_27_g3257__2346(mul_7_27_n_520 ,mul_7_27_n_320 ,mul_7_27_n_103);
  or mul_7_27_g3258__1666(mul_7_27_n_519 ,mul_7_27_n_321 ,mul_7_27_n_142);
  or mul_7_27_g3259__7410(mul_7_27_n_518 ,mul_7_27_n_335 ,mul_7_27_n_72);
  or mul_7_27_g3260__6417(mul_7_27_n_517 ,mul_7_27_n_313 ,mul_7_27_n_142);
  or mul_7_27_g3261__5477(mul_7_27_n_516 ,mul_7_27_n_325 ,mul_7_27_n_121);
  or mul_7_27_g3262__2398(mul_7_27_n_515 ,mul_7_27_n_312 ,mul_7_27_n_96);
  or mul_7_27_g3263__5107(mul_7_27_n_514 ,mul_7_27_n_319 ,mul_7_27_n_121);
  or mul_7_27_g3264__6260(mul_7_27_n_513 ,mul_7_27_n_330 ,mul_7_27_n_102);
  or mul_7_27_g3265__4319(mul_7_27_n_512 ,mul_7_27_n_316 ,mul_7_27_n_120);
  or mul_7_27_g3266__8428(mul_7_27_n_511 ,mul_7_27_n_334 ,mul_7_27_n_141);
  or mul_7_27_g3267__5526(mul_7_27_n_510 ,mul_7_27_n_336 ,mul_7_27_n_69);
  or mul_7_27_g3268__6783(mul_7_27_n_509 ,mul_7_27_n_329 ,mul_7_27_n_72);
  or mul_7_27_g3269__3680(mul_7_27_n_508 ,mul_7_27_n_317 ,mul_7_27_n_100);
  or mul_7_27_g3270__1617(mul_7_27_n_507 ,mul_7_27_n_315 ,mul_7_27_n_102);
  or mul_7_27_g3271__2802(mul_7_27_n_506 ,mul_7_27_n_326 ,mul_7_27_n_120);
  or mul_7_27_g3272__1705(mul_7_27_n_505 ,mul_7_27_n_323 ,mul_7_27_n_118);
  or mul_7_27_g3273__5122(mul_7_27_n_504 ,mul_7_27_n_314 ,mul_7_27_n_96);
  or mul_7_27_g3274__8246(mul_7_27_n_503 ,mul_7_27_n_301 ,mul_7_27_n_100);
  or mul_7_27_g3275__7098(mul_7_27_n_502 ,mul_7_27_n_337 ,mul_7_27_n_103);
  or mul_7_27_g3276__6131(mul_7_27_n_501 ,mul_7_27_n_331 ,mul_7_27_n_141);
  or mul_7_27_g3277__1881(mul_7_27_n_500 ,mul_7_27_n_311 ,mul_7_27_n_118);
  or mul_7_27_g3278__5115(mul_7_27_n_499 ,mul_7_27_n_327 ,mul_7_27_n_97);
  and mul_7_27_g3279__7482(mul_7_27_n_498 ,mul_7_27_n_164 ,mul_7_27_n_408);
  or mul_7_27_g3280__4733(mul_7_27_n_497 ,mul_7_27_n_351 ,mul_7_27_n_408);
  or mul_7_27_g3281__6161(mul_7_27_n_496 ,mul_7_27_n_360 ,mul_7_27_n_36);
  or mul_7_27_g3282__9315(mul_7_27_n_495 ,mul_7_27_n_354 ,mul_7_27_n_55);
  not mul_7_27_g3283(mul_7_27_n_494 ,mul_7_27_n_493);
  not mul_7_27_g3284(mul_7_27_n_492 ,mul_7_27_n_491);
  not mul_7_27_g3285(mul_7_27_n_490 ,mul_7_27_n_489);
  not mul_7_27_g3286(mul_7_27_n_486 ,mul_7_27_n_485);
  or mul_7_27_g3287__9945(mul_7_27_n_484 ,mul_7_27_n_356 ,mul_7_27_n_60);
  or mul_7_27_g3288__2883(mul_7_27_n_483 ,mul_7_27_n_339 ,mul_7_27_n_37);
  or mul_7_27_g3289__2346(mul_7_27_n_482 ,mul_7_27_n_357 ,mul_7_27_n_55);
  or mul_7_27_g3290__1666(mul_7_27_n_481 ,mul_7_27_n_362 ,mul_7_27_n_54);
  or mul_7_27_g3291__7410(mul_7_27_n_480 ,mul_7_27_n_355 ,mul_7_27_n_31);
  nor mul_7_27_g3292__6417(mul_7_27_n_479 ,mul_7_27_n_157 ,mul_7_27_n_353);
  or mul_7_27_g3293__5477(mul_7_27_n_478 ,mul_7_27_n_358 ,mul_7_27_n_31);
  or mul_7_27_g3294__2398(mul_7_27_n_477 ,mul_7_27_n_367 ,mul_7_27_n_61);
  or mul_7_27_g3295__5107(mul_7_27_n_476 ,mul_7_27_n_333 ,mul_7_27_n_36);
  or mul_7_27_g3296__6260(mul_7_27_n_475 ,mul_7_27_n_359 ,mul_7_27_n_54);
  or mul_7_27_g3297__4319(mul_7_27_n_474 ,mul_7_27_n_361 ,mul_7_27_n_60);
  or mul_7_27_g3298__8428(mul_7_27_n_473 ,mul_7_27_n_352 ,mul_7_27_n_37);
  or mul_7_27_g3299__5526(mul_7_27_n_472 ,mul_7_27_n_374 ,mul_7_27_n_63);
  or mul_7_27_g3300__6783(mul_7_27_n_471 ,mul_7_27_n_363 ,mul_7_27_n_58);
  or mul_7_27_g3301__3680(mul_7_27_n_470 ,mul_7_27_n_364 ,mul_7_27_n_45);
  or mul_7_27_g3302__1617(mul_7_27_n_469 ,mul_7_27_n_365 ,mul_7_27_n_45);
  or mul_7_27_g3303__2802(mul_7_27_n_468 ,mul_7_27_n_370 ,mul_7_27_n_63);
  or mul_7_27_g3304__1705(mul_7_27_n_467 ,mul_7_27_n_369 ,mul_7_27_n_46);
  or mul_7_27_g3306__5122(mul_7_27_n_465 ,mul_7_27_n_342 ,mul_7_27_n_64);
  nor mul_7_27_g3307__8246(mul_7_27_n_464 ,mul_7_27_n_64 ,mul_7_27_n_373);
  or mul_7_27_g3308__7098(mul_7_27_n_463 ,mul_7_27_n_372 ,mul_7_27_n_39);
  or mul_7_27_g3309__6131(mul_7_27_n_462 ,mul_7_27_n_368 ,mul_7_27_n_57);
  or mul_7_27_g3310__1881(mul_7_27_n_461 ,mul_7_27_n_376 ,mul_7_27_n_40);
  or mul_7_27_g3311__5115(mul_7_27_n_460 ,mul_7_27_n_377 ,mul_7_27_n_40);
  or mul_7_27_g3312__7482(mul_7_27_n_459 ,mul_7_27_n_371 ,mul_7_27_n_57);
  or mul_7_27_g3313__4733(mul_7_27_n_458 ,mul_7_27_n_375 ,mul_7_27_n_58);
  or mul_7_27_g3314__6161(mul_7_27_n_457 ,mul_7_27_n_366 ,mul_7_27_n_39);
  and mul_7_27_g3315__9315(mul_7_27_n_493 ,in1[5] ,mul_7_27_n_453);
  and mul_7_27_g3316__9945(mul_7_27_n_491 ,in1[3] ,mul_7_27_n_450);
  or mul_7_27_g3317__2883(mul_7_27_n_489 ,mul_7_27_n_51 ,mul_7_27_n_46);
  and mul_7_27_g3318__2346(mul_7_27_n_488 ,in1[3] ,mul_7_27_n_417);
  and mul_7_27_g3319__1666(mul_7_27_n_487 ,in1[5] ,mul_7_27_n_427);
  and mul_7_27_g3320__7410(mul_7_27_n_485 ,in1[7] ,mul_7_27_n_433);
  not mul_7_27_g3321(mul_7_27_n_455 ,mul_7_27_n_453);
  not mul_7_27_g3322(mul_7_27_n_454 ,mul_7_27_n_453);
  not mul_7_27_g3323(mul_7_27_n_452 ,mul_7_27_n_450);
  not mul_7_27_g3324(mul_7_27_n_451 ,mul_7_27_n_450);
  or mul_7_27_g3325__6417(mul_7_27_n_448 ,mul_7_27_n_313 ,mul_7_27_n_138);
  or mul_7_27_g3326__5477(mul_7_27_n_447 ,mul_7_27_n_337 ,mul_7_27_n_126);
  or mul_7_27_g3327__2398(mul_7_27_n_446 ,mul_7_27_n_322 ,mul_7_27_n_93);
  or mul_7_27_g3328__5107(mul_7_27_n_445 ,mul_7_27_n_324 ,mul_7_27_n_132);
  or mul_7_27_g3329__6260(mul_7_27_n_444 ,mul_7_27_n_17 ,mul_7_27_n_339);
  or mul_7_27_g3330__4319(mul_7_27_n_443 ,mul_7_27_n_311 ,mul_7_27_n_135);
  or mul_7_27_g3331__8428(mul_7_27_n_442 ,mul_7_27_n_325 ,mul_7_27_n_123);
  or mul_7_27_g3332__5526(mul_7_27_n_441 ,mul_7_27_n_331 ,mul_7_27_n_139);
  or mul_7_27_g3333__6783(mul_7_27_n_440 ,mul_7_27_n_323 ,mul_7_27_n_139);
  or mul_7_27_g3334__3680(mul_7_27_n_439 ,mul_7_27_n_340 ,mul_7_27_n_144);
  or mul_7_27_g3335__1617(mul_7_27_n_438 ,mul_7_27_n_317 ,mul_7_27_n_127);
  or mul_7_27_g3336__2802(mul_7_27_n_437 ,mul_7_27_n_321 ,mul_7_27_n_94);
  or mul_7_27_g3337__1705(mul_7_27_n_436 ,mul_7_27_n_334 ,mul_7_27_n_93);
  or mul_7_27_g3338__5122(mul_7_27_n_435 ,mul_7_27_n_320 ,mul_7_27_n_127);
  or mul_7_27_g3339__8246(mul_7_27_n_434 ,mul_7_27_n_316 ,mul_7_27_n_129);
  or mul_7_27_g3340__7098(mul_7_27_n_433 ,mul_7_27_n_262 ,mul_7_27_n_350);
  or mul_7_27_g3341__6131(mul_7_27_n_432 ,mul_7_27_n_315 ,mul_7_27_n_133);
  or mul_7_27_g3342__1881(mul_7_27_n_431 ,mul_7_27_n_338 ,mul_7_27_n_132);
  or mul_7_27_g3343__5115(mul_7_27_n_430 ,mul_7_27_n_329 ,mul_7_27_n_124);
  or mul_7_27_g3344__7482(mul_7_27_n_429 ,mul_7_27_n_312 ,mul_7_27_n_136);
  or mul_7_27_g3345__4733(mul_7_27_n_428 ,mul_7_27_n_336 ,mul_7_27_n_145);
  or mul_7_27_g3346__6161(mul_7_27_n_427 ,mul_7_27_n_283 ,mul_7_27_n_347);
  or mul_7_27_g3347__9315(mul_7_27_n_426 ,mul_7_27_n_330 ,mul_7_27_n_130);
  or mul_7_27_g3348__9945(mul_7_27_n_425 ,mul_7_27_n_328 ,mul_7_27_n_126);
  or mul_7_27_g3349__2883(mul_7_27_n_424 ,mul_7_27_n_335 ,mul_7_27_n_123);
  or mul_7_27_g3350__2346(mul_7_27_n_423 ,mul_7_27_n_314 ,mul_7_27_n_138);
  or mul_7_27_g3351__1666(mul_7_27_n_422 ,mul_7_27_n_332 ,mul_7_27_n_135);
  or mul_7_27_g3352__7410(mul_7_27_n_421 ,mul_7_27_n_326 ,mul_7_27_n_124);
  or mul_7_27_g3353__6417(mul_7_27_n_420 ,mul_7_27_n_319 ,mul_7_27_n_133);
  or mul_7_27_g3354__5477(mul_7_27_n_419 ,mul_7_27_n_318 ,mul_7_27_n_136);
  or mul_7_27_g3355__2398(mul_7_27_n_418 ,mul_7_27_n_327 ,mul_7_27_n_94);
  or mul_7_27_g3356__5107(mul_7_27_n_417 ,mul_7_27_n_264 ,mul_7_27_n_349);
  or mul_7_27_g3357__6260(mul_7_27_n_456 ,in1[0] ,mul_7_27_n_341);
  and mul_7_27_g3358__4319(mul_7_27_n_453 ,mul_7_27_n_300 ,mul_7_27_n_130);
  and mul_7_27_g3359__8428(mul_7_27_n_450 ,mul_7_27_n_298 ,mul_7_27_n_145);
  or mul_7_27_g3360__5526(mul_7_27_n_449 ,mul_7_27_n_299 ,mul_7_27_n_308);
  not mul_7_27_g3361(mul_7_27_n_416 ,mul_7_27_n_415);
  not mul_7_27_g3362(mul_7_27_n_414 ,mul_7_27_n_413);
  not mul_7_27_g3363(mul_7_27_n_412 ,mul_7_27_n_411);
  or mul_7_27_g3364__6783(mul_7_27_n_407 ,mul_7_27_n_108 ,mul_7_27_n_373);
  or mul_7_27_g3365__3680(mul_7_27_n_406 ,mul_7_27_n_26 ,mul_7_27_n_354);
  or mul_7_27_g3366__1617(mul_7_27_n_405 ,mul_7_27_n_29 ,mul_7_27_n_333);
  or mul_7_27_g3367__2802(mul_7_27_n_404 ,mul_7_27_n_23 ,mul_7_27_n_360);
  or mul_7_27_g3368__1705(mul_7_27_n_403 ,mul_7_27_n_20 ,mul_7_27_n_356);
  or mul_7_27_g3369__5122(mul_7_27_n_402 ,mul_7_27_n_14 ,mul_7_27_n_353);
  or mul_7_27_g3370__8246(mul_7_27_n_401 ,mul_7_27_n_152 ,mul_7_27_n_352);
  or mul_7_27_g3371__7098(mul_7_27_n_400 ,mul_7_27_n_154 ,mul_7_27_n_357);
  or mul_7_27_g3372__6131(mul_7_27_n_399 ,mul_7_27_n_25 ,mul_7_27_n_355);
  or mul_7_27_g3373__1881(mul_7_27_n_398 ,mul_7_27_n_16 ,mul_7_27_n_367);
  or mul_7_27_g3374__5115(mul_7_27_n_397 ,mul_7_27_n_19 ,mul_7_27_n_358);
  or mul_7_27_g3375__7482(mul_7_27_n_396 ,mul_7_27_n_22 ,mul_7_27_n_359);
  or mul_7_27_g3377__4733(mul_7_27_n_394 ,mul_7_27_n_114 ,mul_7_27_n_365);
  or mul_7_27_g3378__6161(mul_7_27_n_393 ,mul_7_27_n_105 ,mul_7_27_n_368);
  or mul_7_27_g3379__9315(mul_7_27_n_392 ,mul_7_27_n_109 ,mul_7_27_n_376);
  or mul_7_27_g3380__9945(mul_7_27_n_391 ,mul_7_27_n_109 ,mul_7_27_n_364);
  or mul_7_27_g3381__2883(mul_7_27_n_390 ,mul_7_27_n_111 ,mul_7_27_n_377);
  or mul_7_27_g3382__2346(mul_7_27_n_389 ,mul_7_27_n_13 ,mul_7_27_n_362);
  or mul_7_27_g3383__1666(mul_7_27_n_388 ,mul_7_27_n_115 ,mul_7_27_n_372);
  or mul_7_27_g3384__7410(mul_7_27_n_387 ,mul_7_27_n_114 ,mul_7_27_n_370);
  or mul_7_27_g3385__6417(mul_7_27_n_386 ,mul_7_27_n_106 ,mul_7_27_n_369);
  or mul_7_27_g3386__5477(mul_7_27_n_385 ,mul_7_27_n_112 ,mul_7_27_n_371);
  or mul_7_27_g3387__2398(mul_7_27_n_384 ,mul_7_27_n_108 ,mul_7_27_n_366);
  or mul_7_27_g3388__5107(mul_7_27_n_383 ,mul_7_27_n_105 ,mul_7_27_n_374);
  or mul_7_27_g3389__6260(mul_7_27_n_382 ,mul_7_27_n_106 ,mul_7_27_n_375);
  or mul_7_27_g3390__4319(mul_7_27_n_381 ,mul_7_27_n_115 ,mul_7_27_n_363);
  and mul_7_27_g3391__8428(out1[1] ,mul_7_27_n_348 ,mul_7_27_n_164);
  xnor mul_7_27_g3392__5526(mul_7_27_n_379 ,mul_7_27_n_166 ,in1[1]);
  xnor mul_7_27_g3393__6783(mul_7_27_n_378 ,mul_7_27_n_165 ,in1[1]);
  or mul_7_27_g3394__3680(mul_7_27_n_415 ,mul_7_27_n_34 ,mul_7_27_n_112);
  and mul_7_27_g3395__1617(mul_7_27_n_413 ,in1[5] ,mul_7_27_n_305);
  and mul_7_27_g3396__2802(mul_7_27_n_411 ,in1[3] ,mul_7_27_n_302);
  or mul_7_27_g3397__1705(mul_7_27_n_410 ,mul_7_27_n_29 ,mul_7_27_n_129);
  or mul_7_27_g3398__5122(mul_7_27_n_409 ,mul_7_27_n_23 ,mul_7_27_n_111);
  or mul_7_27_g3399__8246(mul_7_27_n_408 ,mul_7_27_n_26 ,mul_7_27_n_144);
  and mul_7_27_g3400__7098(mul_7_27_n_350 ,mul_7_27_n_17 ,mul_7_27_n_284);
  and mul_7_27_g3401__6131(mul_7_27_n_349 ,mul_7_27_n_20 ,mul_7_27_n_285);
  and mul_7_27_g3403__1881(mul_7_27_n_347 ,mul_7_27_n_14 ,mul_7_27_n_268);
  or mul_7_27_g3404__5115(mul_7_27_n_346 ,mul_7_27_n_148 ,mul_7_27_n_296);
  or mul_7_27_g3405__7482(mul_7_27_n_345 ,mul_7_27_n_150 ,mul_7_27_n_275);
  and mul_7_27_g3406__4733(mul_7_27_n_344 ,mul_7_27_n_147 ,mul_7_27_n_165);
  and mul_7_27_g3407__6161(mul_7_27_n_343 ,mul_7_27_n_10 ,mul_7_27_n_166);
  or mul_7_27_g3408__9315(mul_7_27_n_342 ,mul_7_27_n_272 ,mul_7_27_n_267);
  or mul_7_27_g3410__9945(mul_7_27_n_377 ,mul_7_27_n_273 ,mul_7_27_n_279);
  or mul_7_27_g3411__2883(mul_7_27_n_376 ,mul_7_27_n_240 ,mul_7_27_n_261);
  or mul_7_27_g3412__2346(mul_7_27_n_375 ,mul_7_27_n_238 ,mul_7_27_n_280);
  or mul_7_27_g3413__1666(mul_7_27_n_374 ,mul_7_27_n_237 ,mul_7_27_n_263);
  xnor mul_7_27_g3414__7410(mul_7_27_n_373 ,mul_7_27_n_179 ,in1[7]);
  or mul_7_27_g3415__6417(mul_7_27_n_372 ,mul_7_27_n_246 ,mul_7_27_n_259);
  or mul_7_27_g3416__5477(mul_7_27_n_371 ,mul_7_27_n_243 ,mul_7_27_n_260);
  or mul_7_27_g3417__2398(mul_7_27_n_370 ,mul_7_27_n_248 ,mul_7_27_n_281);
  or mul_7_27_g3418__5107(mul_7_27_n_369 ,mul_7_27_n_247 ,mul_7_27_n_269);
  or mul_7_27_g3419__6260(mul_7_27_n_368 ,mul_7_27_n_241 ,mul_7_27_n_270);
  xnor mul_7_27_g3420__4319(mul_7_27_n_367 ,mul_7_27_n_76 ,in1[1]);
  or mul_7_27_g3421__8428(mul_7_27_n_366 ,mul_7_27_n_239 ,mul_7_27_n_286);
  or mul_7_27_g3422__5526(mul_7_27_n_365 ,mul_7_27_n_242 ,mul_7_27_n_271);
  or mul_7_27_g3423__6783(mul_7_27_n_364 ,mul_7_27_n_245 ,mul_7_27_n_266);
  or mul_7_27_g3424__3680(mul_7_27_n_363 ,mul_7_27_n_244 ,mul_7_27_n_265);
  xnor mul_7_27_g3425__1617(mul_7_27_n_362 ,mul_7_27_n_78 ,in1[1]);
  xnor mul_7_27_g3426__2802(mul_7_27_n_361 ,mul_7_27_n_73 ,in1[1]);
  xnor mul_7_27_g3427__1705(mul_7_27_n_360 ,mul_7_27_n_74 ,in1[1]);
  xnor mul_7_27_g3428__5122(mul_7_27_n_359 ,mul_7_27_n_82 ,in1[1]);
  xnor mul_7_27_g3429__8246(mul_7_27_n_358 ,mul_7_27_n_79 ,in1[1]);
  xnor mul_7_27_g3430__7098(mul_7_27_n_357 ,mul_7_27_n_83 ,in1[1]);
  xnor mul_7_27_g3431__6131(mul_7_27_n_356 ,mul_7_27_n_81 ,in1[1]);
  xnor mul_7_27_g3432__1881(mul_7_27_n_355 ,mul_7_27_n_80 ,in1[1]);
  xnor mul_7_27_g3433__5115(mul_7_27_n_354 ,mul_7_27_n_84 ,in1[1]);
  xnor mul_7_27_g3434__7482(mul_7_27_n_353 ,mul_7_27_n_66 ,in1[1]);
  xnor mul_7_27_g3435__4733(mul_7_27_n_352 ,mul_7_27_n_85 ,in1[1]);
  not mul_7_27_g3437(mul_7_27_n_310 ,mul_7_27_n_308);
  not mul_7_27_g3438(mul_7_27_n_309 ,mul_7_27_n_308);
  not mul_7_27_g3439(mul_7_27_n_307 ,mul_7_27_n_305);
  not mul_7_27_g3440(mul_7_27_n_306 ,mul_7_27_n_305);
  not mul_7_27_g3441(mul_7_27_n_304 ,mul_7_27_n_302);
  not mul_7_27_g3442(mul_7_27_n_303 ,mul_7_27_n_302);
  xnor mul_7_27_g3443__6161(mul_7_27_n_301 ,in1[5] ,in1[0]);
  xor mul_7_27_g3444__9315(mul_7_27_n_300 ,in1[5] ,in1[4]);
  xnor mul_7_27_g3445__9945(mul_7_27_n_299 ,in1[7] ,in1[6]);
  xor mul_7_27_g3446__2883(mul_7_27_n_298 ,in1[3] ,in1[2]);
  xnor mul_7_27_g3447__2346(mul_7_27_n_297 ,in1[3] ,in1[0]);
  xnor mul_7_27_g3448__1666(mul_7_27_n_340 ,mul_7_27_n_82 ,in1[3]);
  xnor mul_7_27_g3449__7410(mul_7_27_n_339 ,mul_7_27_n_75 ,in1[1]);
  xnor mul_7_27_g3450__6417(mul_7_27_n_338 ,mul_7_27_n_77 ,in1[5]);
  xnor mul_7_27_g3451__5477(mul_7_27_n_337 ,mul_7_27_n_79 ,in1[5]);
  xnor mul_7_27_g3452__2398(mul_7_27_n_336 ,mul_7_27_n_77 ,in1[3]);
  xnor mul_7_27_g3453__5107(mul_7_27_n_335 ,mul_7_27_n_212 ,in1[5]);
  xnor mul_7_27_g3454__6260(mul_7_27_n_334 ,mul_7_27_n_200 ,in1[3]);
  xnor mul_7_27_g3455__4319(mul_7_27_n_333 ,mul_7_27_n_197 ,in1[1]);
  xnor mul_7_27_g3456__8428(mul_7_27_n_332 ,mul_7_27_n_180 ,in1[3]);
  xnor mul_7_27_g3457__5526(mul_7_27_n_331 ,mul_7_27_n_85 ,in1[3]);
  xnor mul_7_27_g3458__6783(mul_7_27_n_330 ,mul_7_27_n_76 ,in1[5]);
  xnor mul_7_27_g3459__3680(mul_7_27_n_329 ,mul_7_27_n_218 ,in1[5]);
  xnor mul_7_27_g3460__1617(mul_7_27_n_328 ,mul_7_27_n_66 ,in1[5]);
  xnor mul_7_27_g3461__2802(mul_7_27_n_327 ,mul_7_27_n_74 ,in1[3]);
  xnor mul_7_27_g3462__1705(mul_7_27_n_326 ,mul_7_27_n_78 ,in1[5]);
  xnor mul_7_27_g3463__5122(mul_7_27_n_325 ,mul_7_27_n_75 ,in1[5]);
  xnor mul_7_27_g3464__8246(mul_7_27_n_324 ,mul_7_27_n_80 ,in1[5]);
  xnor mul_7_27_g3465__7098(mul_7_27_n_323 ,mul_7_27_n_83 ,in1[3]);
  xnor mul_7_27_g3466__6131(mul_7_27_n_322 ,mul_7_27_n_209 ,in1[3]);
  xnor mul_7_27_g3467__1881(mul_7_27_n_321 ,mul_7_27_n_194 ,in1[3]);
  xnor mul_7_27_g3468__5115(mul_7_27_n_320 ,mul_7_27_n_203 ,in1[5]);
  xnor mul_7_27_g3469__7482(mul_7_27_n_319 ,mul_7_27_n_84 ,in1[5]);
  xnor mul_7_27_g3470__4733(mul_7_27_n_318 ,mul_7_27_n_185 ,in1[3]);
  xnor mul_7_27_g3471__6161(mul_7_27_n_317 ,mul_7_27_n_188 ,in1[5]);
  xnor mul_7_27_g3472__9315(mul_7_27_n_316 ,mul_7_27_n_81 ,in1[5]);
  xnor mul_7_27_g3473__9945(mul_7_27_n_315 ,mul_7_27_n_73 ,in1[5]);
  xnor mul_7_27_g3474__2883(mul_7_27_n_314 ,mul_7_27_n_182 ,in1[3]);
  xnor mul_7_27_g3475__2346(mul_7_27_n_313 ,mul_7_27_n_215 ,in1[3]);
  xnor mul_7_27_g3476__1666(mul_7_27_n_312 ,mul_7_27_n_191 ,in1[3]);
  xnor mul_7_27_g3477__7410(mul_7_27_n_311 ,mul_7_27_n_206 ,in1[3]);
  xor mul_7_27_g3478__6417(mul_7_27_n_308 ,in1[6] ,in1[5]);
  xor mul_7_27_g3479__5477(mul_7_27_n_305 ,in1[4] ,in1[3]);
  xnor mul_7_27_g3480__2398(mul_7_27_n_302 ,mul_7_27_n_11 ,in1[2]);
  nor mul_7_27_g3491__5107(mul_7_27_n_286 ,mul_7_27_n_185 ,in1[7]);
  or mul_7_27_g3492__6260(mul_7_27_n_285 ,mul_7_27_n_257 ,mul_7_27_n_11);
  or mul_7_27_g3493__4319(mul_7_27_n_284 ,mul_7_27_n_256 ,mul_7_27_n_250);
  nor mul_7_27_g3494__8428(mul_7_27_n_283 ,in1[4] ,in1[3]);
  nor mul_7_27_g3495__5526(mul_7_27_n_282 ,mul_7_27_n_154 ,mul_7_27_n_148);
  nor mul_7_27_g3496__6783(mul_7_27_n_281 ,mul_7_27_n_206 ,in1[7]);
  nor mul_7_27_g3497__3680(mul_7_27_n_280 ,mul_7_27_n_203 ,in1[7]);
  nor mul_7_27_g3498__1617(mul_7_27_n_279 ,mul_7_27_n_200 ,in1[7]);
  or mul_7_27_g3499__2802(mul_7_27_n_296 ,mul_7_27_n_233 ,mul_7_27_n_48);
  or mul_7_27_g3500__1705(mul_7_27_n_295 ,mul_7_27_n_230 ,mul_7_27_n_33);
  or mul_7_27_g3501__5122(mul_7_27_n_294 ,mul_7_27_n_225 ,mul_7_27_n_43);
  or mul_7_27_g3502__8246(mul_7_27_n_293 ,mul_7_27_n_234 ,mul_7_27_n_52);
  or mul_7_27_g3503__7098(mul_7_27_n_292 ,mul_7_27_n_228 ,mul_7_27_n_49);
  or mul_7_27_g3504__6131(mul_7_27_n_291 ,mul_7_27_n_235 ,mul_7_27_n_34);
  or mul_7_27_g3505__1881(mul_7_27_n_290 ,mul_7_27_n_229 ,mul_7_27_n_42);
  or mul_7_27_g3506__5115(mul_7_27_n_289 ,mul_7_27_n_236 ,mul_7_27_n_51);
  or mul_7_27_g3507__7482(mul_7_27_n_288 ,mul_7_27_n_226 ,mul_7_27_n_48);
  or mul_7_27_g3508__4733(mul_7_27_n_287 ,mul_7_27_n_232 ,mul_7_27_n_33);
  not mul_7_27_g3512(mul_7_27_n_273 ,mul_7_27_n_274);
  nor mul_7_27_g3514__6161(mul_7_27_n_271 ,mul_7_27_n_191 ,in1[7]);
  nor mul_7_27_g3515__9315(mul_7_27_n_270 ,mul_7_27_n_194 ,in1[7]);
  nor mul_7_27_g3516__9945(mul_7_27_n_269 ,mul_7_27_n_182 ,in1[7]);
  or mul_7_27_g3517__2883(mul_7_27_n_268 ,mul_7_27_n_252 ,mul_7_27_n_253);
  nor mul_7_27_g3518__2346(mul_7_27_n_267 ,in1[7] ,in1[0]);
  nor mul_7_27_g3519__1666(mul_7_27_n_266 ,mul_7_27_n_212 ,in1[7]);
  nor mul_7_27_g3520__7410(mul_7_27_n_265 ,mul_7_27_n_197 ,in1[7]);
  nor mul_7_27_g3521__6417(mul_7_27_n_264 ,in1[2] ,in1[1]);
  nor mul_7_27_g3522__5477(mul_7_27_n_263 ,mul_7_27_n_209 ,in1[7]);
  nor mul_7_27_g3523__2398(mul_7_27_n_262 ,in1[6] ,in1[5]);
  nor mul_7_27_g3524__5107(mul_7_27_n_261 ,mul_7_27_n_215 ,in1[7]);
  nor mul_7_27_g3525__6260(mul_7_27_n_260 ,mul_7_27_n_218 ,in1[7]);
  nor mul_7_27_g3526__4319(mul_7_27_n_259 ,mul_7_27_n_188 ,in1[7]);
  or mul_7_27_g3527__8428(mul_7_27_n_258 ,mul_7_27_n_251 ,mul_7_27_n_43);
  and mul_7_27_g3528__5526(mul_7_27_n_277 ,in1[1] ,mul_7_27_n_28);
  or mul_7_27_g3529__6783(mul_7_27_n_276 ,mul_7_27_n_231 ,mul_7_27_n_52);
  or mul_7_27_g3530__3680(mul_7_27_n_275 ,mul_7_27_n_224 ,mul_7_27_n_49);
  or mul_7_27_g3531__1617(mul_7_27_n_274 ,mul_7_27_n_227 ,mul_7_27_n_42);
  and mul_7_27_g3532__2802(mul_7_27_n_272 ,in1[7] ,in1[0]);
  not mul_7_27_g3533(mul_7_27_n_257 ,in1[2]);
  not mul_7_27_g3534(mul_7_27_n_256 ,in1[6]);
  not mul_7_27_g3541(mul_7_27_n_255 ,in1[0]);
  not mul_7_27_g3542(mul_7_27_n_254 ,in1[7]);
  not mul_7_27_g3543(mul_7_27_n_253 ,in1[3]);
  not mul_7_27_g3544(mul_7_27_n_252 ,in1[4]);
  not mul_7_27_g3546(mul_7_27_n_251 ,mul_7_27_n_180);
  not mul_7_27_g3553(mul_7_27_n_250 ,in1[5]);
  not mul_7_27_g3554(mul_7_27_n_249 ,in1[1]);
  not mul_7_27_drc_bufs(mul_7_27_n_223 ,mul_7_27_n_90);
  not mul_7_27_drc_bufs3555(mul_7_27_n_222 ,mul_7_27_n_91);
  not mul_7_27_drc_bufs3556(mul_7_27_n_221 ,mul_7_27_n_90);
  not mul_7_27_drc_bufs3557(mul_7_27_n_220 ,mul_7_27_n_91);
  not mul_7_27_drc_bufs3639(mul_7_27_n_219 ,mul_7_27_n_217);
  not mul_7_27_drc_bufs3640(mul_7_27_n_218 ,mul_7_27_n_217);
  not mul_7_27_drc_bufs3641(mul_7_27_n_217 ,n_2);
  not mul_7_27_drc_bufs3643(mul_7_27_n_216 ,mul_7_27_n_214);
  not mul_7_27_drc_bufs3644(mul_7_27_n_215 ,mul_7_27_n_214);
  not mul_7_27_drc_bufs3645(mul_7_27_n_214 ,n_3);
  not mul_7_27_drc_bufs3647(mul_7_27_n_213 ,mul_7_27_n_211);
  not mul_7_27_drc_bufs3648(mul_7_27_n_212 ,mul_7_27_n_211);
  not mul_7_27_drc_bufs3649(mul_7_27_n_211 ,n_4);
  not mul_7_27_drc_bufs3651(mul_7_27_n_210 ,mul_7_27_n_208);
  not mul_7_27_drc_bufs3652(mul_7_27_n_209 ,mul_7_27_n_208);
  not mul_7_27_drc_bufs3653(mul_7_27_n_208 ,n_8);
  not mul_7_27_drc_bufs3655(mul_7_27_n_207 ,mul_7_27_n_205);
  not mul_7_27_drc_bufs3656(mul_7_27_n_206 ,mul_7_27_n_205);
  not mul_7_27_drc_bufs3657(mul_7_27_n_205 ,n_9);
  not mul_7_27_drc_bufs3659(mul_7_27_n_204 ,mul_7_27_n_202);
  not mul_7_27_drc_bufs3660(mul_7_27_n_203 ,mul_7_27_n_202);
  not mul_7_27_drc_bufs3661(mul_7_27_n_202 ,n_10);
  not mul_7_27_drc_bufs3663(mul_7_27_n_201 ,mul_7_27_n_199);
  not mul_7_27_drc_bufs3664(mul_7_27_n_200 ,mul_7_27_n_199);
  not mul_7_27_drc_bufs3665(mul_7_27_n_199 ,n_11);
  not mul_7_27_drc_bufs3667(mul_7_27_n_198 ,mul_7_27_n_196);
  not mul_7_27_drc_bufs3668(mul_7_27_n_197 ,mul_7_27_n_196);
  not mul_7_27_drc_bufs3669(mul_7_27_n_196 ,n_5);
  not mul_7_27_drc_bufs3671(mul_7_27_n_195 ,mul_7_27_n_193);
  not mul_7_27_drc_bufs3672(mul_7_27_n_194 ,mul_7_27_n_193);
  not mul_7_27_drc_bufs3673(mul_7_27_n_193 ,n_12);
  not mul_7_27_drc_bufs3675(mul_7_27_n_192 ,mul_7_27_n_190);
  not mul_7_27_drc_bufs3676(mul_7_27_n_191 ,mul_7_27_n_190);
  not mul_7_27_drc_bufs3677(mul_7_27_n_190 ,n_6);
  not mul_7_27_drc_bufs3679(mul_7_27_n_189 ,mul_7_27_n_187);
  not mul_7_27_drc_bufs3680(mul_7_27_n_188 ,mul_7_27_n_187);
  not mul_7_27_drc_bufs3681(mul_7_27_n_187 ,n_13);
  not mul_7_27_drc_bufs3683(mul_7_27_n_186 ,mul_7_27_n_184);
  not mul_7_27_drc_bufs3684(mul_7_27_n_185 ,mul_7_27_n_184);
  not mul_7_27_drc_bufs3685(mul_7_27_n_184 ,n_7);
  not mul_7_27_drc_bufs3687(mul_7_27_n_183 ,mul_7_27_n_181);
  not mul_7_27_drc_bufs3688(mul_7_27_n_182 ,mul_7_27_n_181);
  not mul_7_27_drc_bufs3689(mul_7_27_n_181 ,n_1);
  not mul_7_27_drc_bufs3691(mul_7_27_n_180 ,mul_7_27_n_178);
  not mul_7_27_drc_bufs3692(mul_7_27_n_179 ,mul_7_27_n_178);
  not mul_7_27_drc_bufs3693(mul_7_27_n_178 ,n_14);
  not mul_7_27_drc_bufs3696(mul_7_27_n_177 ,mul_7_27_n_176);
  not mul_7_27_drc_bufs3697(mul_7_27_n_176 ,mul_7_27_n_531);
  not mul_7_27_drc_bufs3700(mul_7_27_n_175 ,mul_7_27_n_239);
  not mul_7_27_drc_bufs3701(mul_7_27_n_239 ,mul_7_27_n_287);
  not mul_7_27_drc_bufs3704(mul_7_27_n_174 ,mul_7_27_n_238);
  not mul_7_27_drc_bufs3705(mul_7_27_n_238 ,mul_7_27_n_276);
  not mul_7_27_drc_bufs3708(mul_7_27_n_173 ,mul_7_27_n_247);
  not mul_7_27_drc_bufs3709(mul_7_27_n_247 ,mul_7_27_n_295);
  not mul_7_27_drc_bufs3713(mul_7_27_n_246 ,mul_7_27_n_294);
  not mul_7_27_drc_bufs3716(mul_7_27_n_172 ,mul_7_27_n_244);
  not mul_7_27_drc_bufs3717(mul_7_27_n_244 ,mul_7_27_n_292);
  not mul_7_27_drc_bufs3720(mul_7_27_n_171 ,mul_7_27_n_242);
  not mul_7_27_drc_bufs3721(mul_7_27_n_242 ,mul_7_27_n_290);
  not mul_7_27_drc_bufs3724(mul_7_27_n_170 ,mul_7_27_n_245);
  not mul_7_27_drc_bufs3725(mul_7_27_n_245 ,mul_7_27_n_293);
  not mul_7_27_drc_bufs3728(mul_7_27_n_169 ,mul_7_27_n_240);
  not mul_7_27_drc_bufs3729(mul_7_27_n_240 ,mul_7_27_n_288);
  not mul_7_27_drc_bufs3732(mul_7_27_n_168 ,mul_7_27_n_243);
  not mul_7_27_drc_bufs3733(mul_7_27_n_243 ,mul_7_27_n_291);
  not mul_7_27_drc_bufs3736(mul_7_27_n_167 ,mul_7_27_n_241);
  not mul_7_27_drc_bufs3737(mul_7_27_n_241 ,mul_7_27_n_289);
  not mul_7_27_drc_bufs3740(mul_7_27_n_166 ,mul_7_27_n_237);
  not mul_7_27_drc_bufs3741(mul_7_27_n_237 ,mul_7_27_n_275);
  not mul_7_27_drc_bufs3744(mul_7_27_n_165 ,mul_7_27_n_248);
  not mul_7_27_drc_bufs3745(mul_7_27_n_248 ,mul_7_27_n_296);
  not mul_7_27_drc_bufs3748(mul_7_27_n_164 ,mul_7_27_n_163);
  not mul_7_27_drc_bufs3749(mul_7_27_n_163 ,mul_7_27_n_351);
  not mul_7_27_drc_bufs3756(mul_7_27_n_162 ,mul_7_27_n_272);
  not mul_7_27_drc_bufs3769(mul_7_27_n_161 ,mul_7_27_n_160);
  not mul_7_27_drc_bufs3771(mul_7_27_n_160 ,mul_7_27_n_449);
  not mul_7_27_drc_bufs3779(mul_7_27_n_159 ,mul_7_27_n_158);
  not mul_7_27_drc_bufs3781(mul_7_27_n_158 ,mul_7_27_n_254);
  not mul_7_27_drc_bufs3784(mul_7_27_n_157 ,mul_7_27_n_155);
  not mul_7_27_drc_bufs3785(mul_7_27_n_156 ,mul_7_27_n_155);
  not mul_7_27_drc_bufs3786(mul_7_27_n_155 ,mul_7_27_n_456);
  not mul_7_27_drc_bufs3796(mul_7_27_n_154 ,mul_7_27_n_153);
  not mul_7_27_drc_bufs3798(mul_7_27_n_153 ,mul_7_27_n_223);
  not mul_7_27_drc_bufs3800(mul_7_27_n_152 ,mul_7_27_n_151);
  not mul_7_27_drc_bufs3802(mul_7_27_n_151 ,mul_7_27_n_222);
  not mul_7_27_drc_bufs3804(mul_7_27_n_150 ,mul_7_27_n_149);
  not mul_7_27_drc_bufs3806(mul_7_27_n_149 ,mul_7_27_n_249);
  not mul_7_27_drc_bufs3808(mul_7_27_n_148 ,mul_7_27_n_146);
  not mul_7_27_drc_bufs3809(mul_7_27_n_147 ,mul_7_27_n_146);
  not mul_7_27_drc_bufs3810(mul_7_27_n_146 ,mul_7_27_n_249);
  not mul_7_27_drc_bufs3812(mul_7_27_n_145 ,mul_7_27_n_143);
  not mul_7_27_drc_bufs3813(mul_7_27_n_144 ,mul_7_27_n_143);
  not mul_7_27_drc_bufs3814(mul_7_27_n_143 ,mul_7_27_n_304);
  not mul_7_27_drc_bufs3816(mul_7_27_n_142 ,mul_7_27_n_140);
  not mul_7_27_drc_bufs3817(mul_7_27_n_141 ,mul_7_27_n_140);
  not mul_7_27_drc_bufs3818(mul_7_27_n_140 ,mul_7_27_n_451);
  not mul_7_27_drc_bufs3820(mul_7_27_n_139 ,mul_7_27_n_137);
  not mul_7_27_drc_bufs3821(mul_7_27_n_138 ,mul_7_27_n_137);
  not mul_7_27_drc_bufs3822(mul_7_27_n_137 ,mul_7_27_n_303);
  not mul_7_27_drc_bufs3824(mul_7_27_n_136 ,mul_7_27_n_134);
  not mul_7_27_drc_bufs3825(mul_7_27_n_135 ,mul_7_27_n_134);
  not mul_7_27_drc_bufs3826(mul_7_27_n_134 ,mul_7_27_n_303);
  not mul_7_27_drc_bufs3828(mul_7_27_n_133 ,mul_7_27_n_131);
  not mul_7_27_drc_bufs3829(mul_7_27_n_132 ,mul_7_27_n_131);
  not mul_7_27_drc_bufs3830(mul_7_27_n_131 ,mul_7_27_n_307);
  not mul_7_27_drc_bufs3832(mul_7_27_n_130 ,mul_7_27_n_128);
  not mul_7_27_drc_bufs3833(mul_7_27_n_129 ,mul_7_27_n_128);
  not mul_7_27_drc_bufs3834(mul_7_27_n_128 ,mul_7_27_n_307);
  not mul_7_27_drc_bufs3836(mul_7_27_n_127 ,mul_7_27_n_125);
  not mul_7_27_drc_bufs3837(mul_7_27_n_126 ,mul_7_27_n_125);
  not mul_7_27_drc_bufs3838(mul_7_27_n_125 ,mul_7_27_n_306);
  not mul_7_27_drc_bufs3840(mul_7_27_n_124 ,mul_7_27_n_122);
  not mul_7_27_drc_bufs3841(mul_7_27_n_123 ,mul_7_27_n_122);
  not mul_7_27_drc_bufs3842(mul_7_27_n_122 ,mul_7_27_n_306);
  not mul_7_27_drc_bufs3844(mul_7_27_n_121 ,mul_7_27_n_119);
  not mul_7_27_drc_bufs3845(mul_7_27_n_120 ,mul_7_27_n_119);
  not mul_7_27_drc_bufs3846(mul_7_27_n_119 ,mul_7_27_n_454);
  not mul_7_27_drc_bufs3848(mul_7_27_n_118 ,mul_7_27_n_116);
  not mul_7_27_drc_bufs3849(mul_7_27_n_117 ,mul_7_27_n_116);
  not mul_7_27_drc_bufs3850(mul_7_27_n_116 ,mul_7_27_n_452);
  not mul_7_27_drc_bufs3852(mul_7_27_n_115 ,mul_7_27_n_113);
  not mul_7_27_drc_bufs3853(mul_7_27_n_114 ,mul_7_27_n_113);
  not mul_7_27_drc_bufs3854(mul_7_27_n_113 ,mul_7_27_n_310);
  not mul_7_27_drc_bufs3856(mul_7_27_n_112 ,mul_7_27_n_110);
  not mul_7_27_drc_bufs3857(mul_7_27_n_111 ,mul_7_27_n_110);
  not mul_7_27_drc_bufs3858(mul_7_27_n_110 ,mul_7_27_n_310);
  not mul_7_27_drc_bufs3860(mul_7_27_n_109 ,mul_7_27_n_107);
  not mul_7_27_drc_bufs3861(mul_7_27_n_108 ,mul_7_27_n_107);
  not mul_7_27_drc_bufs3862(mul_7_27_n_107 ,mul_7_27_n_309);
  not mul_7_27_drc_bufs3864(mul_7_27_n_106 ,mul_7_27_n_104);
  not mul_7_27_drc_bufs3865(mul_7_27_n_105 ,mul_7_27_n_104);
  not mul_7_27_drc_bufs3866(mul_7_27_n_104 ,mul_7_27_n_309);
  not mul_7_27_drc_bufs3868(mul_7_27_n_103 ,mul_7_27_n_101);
  not mul_7_27_drc_bufs3869(mul_7_27_n_102 ,mul_7_27_n_101);
  not mul_7_27_drc_bufs3870(mul_7_27_n_101 ,mul_7_27_n_455);
  not mul_7_27_drc_bufs3872(mul_7_27_n_100 ,mul_7_27_n_98);
  not mul_7_27_drc_bufs3873(mul_7_27_n_99 ,mul_7_27_n_98);
  not mul_7_27_drc_bufs3874(mul_7_27_n_98 ,mul_7_27_n_455);
  not mul_7_27_drc_bufs3876(mul_7_27_n_97 ,mul_7_27_n_95);
  not mul_7_27_drc_bufs3877(mul_7_27_n_96 ,mul_7_27_n_95);
  not mul_7_27_drc_bufs3878(mul_7_27_n_95 ,mul_7_27_n_452);
  not mul_7_27_drc_bufs3880(mul_7_27_n_94 ,mul_7_27_n_92);
  not mul_7_27_drc_bufs3881(mul_7_27_n_93 ,mul_7_27_n_92);
  not mul_7_27_drc_bufs3882(mul_7_27_n_92 ,mul_7_27_n_304);
  not mul_7_27_drc_bufs3884(mul_7_27_n_91 ,mul_7_27_n_255);
  not mul_7_27_drc_bufs3885(mul_7_27_n_90 ,mul_7_27_n_255);
  not mul_7_27_drc_bufs3888(mul_7_27_n_89 ,mul_7_27_n_88);
  not mul_7_27_drc_bufs3890(mul_7_27_n_88 ,mul_7_27_n_529);
  not mul_7_27_drc_bufs3892(mul_7_27_n_87 ,mul_7_27_n_86);
  not mul_7_27_drc_bufs3894(mul_7_27_n_86 ,mul_7_27_n_529);
  not mul_7_27_drc_bufs3897(mul_7_27_n_85 ,mul_7_27_n_235);
  not mul_7_27_drc_bufs3898(mul_7_27_n_235 ,mul_7_27_n_219);
  not mul_7_27_drc_bufs3901(mul_7_27_n_84 ,mul_7_27_n_226);
  not mul_7_27_drc_bufs3902(mul_7_27_n_226 ,mul_7_27_n_216);
  not mul_7_27_drc_bufs3905(mul_7_27_n_83 ,mul_7_27_n_225);
  not mul_7_27_drc_bufs3906(mul_7_27_n_225 ,mul_7_27_n_189);
  not mul_7_27_drc_bufs3909(mul_7_27_n_82 ,mul_7_27_n_234);
  not mul_7_27_drc_bufs3910(mul_7_27_n_234 ,mul_7_27_n_213);
  not mul_7_27_drc_bufs3913(mul_7_27_n_81 ,mul_7_27_n_233);
  not mul_7_27_drc_bufs3914(mul_7_27_n_233 ,mul_7_27_n_207);
  not mul_7_27_drc_bufs3917(mul_7_27_n_80 ,mul_7_27_n_229);
  not mul_7_27_drc_bufs3918(mul_7_27_n_229 ,mul_7_27_n_192);
  not mul_7_27_drc_bufs3921(mul_7_27_n_79 ,mul_7_27_n_227);
  not mul_7_27_drc_bufs3922(mul_7_27_n_227 ,mul_7_27_n_201);
  not mul_7_27_drc_bufs3925(mul_7_27_n_78 ,mul_7_27_n_232);
  not mul_7_27_drc_bufs3926(mul_7_27_n_232 ,mul_7_27_n_186);
  not mul_7_27_drc_bufs3929(mul_7_27_n_77 ,mul_7_27_n_228);
  not mul_7_27_drc_bufs3930(mul_7_27_n_228 ,mul_7_27_n_198);
  not mul_7_27_drc_bufs3933(mul_7_27_n_76 ,mul_7_27_n_236);
  not mul_7_27_drc_bufs3934(mul_7_27_n_236 ,mul_7_27_n_195);
  not mul_7_27_drc_bufs3937(mul_7_27_n_75 ,mul_7_27_n_224);
  not mul_7_27_drc_bufs3938(mul_7_27_n_224 ,mul_7_27_n_210);
  not mul_7_27_drc_bufs3941(mul_7_27_n_74 ,mul_7_27_n_231);
  not mul_7_27_drc_bufs3942(mul_7_27_n_231 ,mul_7_27_n_204);
  not mul_7_27_drc_bufs3945(mul_7_27_n_73 ,mul_7_27_n_230);
  not mul_7_27_drc_bufs3946(mul_7_27_n_230 ,mul_7_27_n_183);
  not mul_7_27_drc_bufs3948(mul_7_27_n_72 ,mul_7_27_n_70);
  not mul_7_27_drc_bufs3949(mul_7_27_n_71 ,mul_7_27_n_70);
  not mul_7_27_drc_bufs3950(mul_7_27_n_70 ,mul_7_27_n_454);
  not mul_7_27_drc_bufs3952(mul_7_27_n_69 ,mul_7_27_n_67);
  not mul_7_27_drc_bufs3953(mul_7_27_n_68 ,mul_7_27_n_67);
  not mul_7_27_drc_bufs3954(mul_7_27_n_67 ,mul_7_27_n_451);
  not mul_7_27_drc_bufs3956(mul_7_27_n_66 ,mul_7_27_n_65);
  not mul_7_27_drc_bufs3958(mul_7_27_n_65 ,mul_7_27_n_179);
  not mul_7_27_drc_bufs3960(mul_7_27_n_64 ,mul_7_27_n_62);
  not mul_7_27_drc_bufs3961(mul_7_27_n_63 ,mul_7_27_n_62);
  not mul_7_27_drc_bufs3962(mul_7_27_n_62 ,mul_7_27_n_449);
  not mul_7_27_drc_bufs3964(mul_7_27_n_61 ,mul_7_27_n_59);
  not mul_7_27_drc_bufs3965(mul_7_27_n_60 ,mul_7_27_n_59);
  not mul_7_27_drc_bufs3966(mul_7_27_n_59 ,mul_7_27_n_456);
  not mul_7_27_drc_bufs3968(mul_7_27_n_58 ,mul_7_27_n_56);
  not mul_7_27_drc_bufs3969(mul_7_27_n_57 ,mul_7_27_n_56);
  not mul_7_27_drc_bufs3970(mul_7_27_n_56 ,mul_7_27_n_449);
  not mul_7_27_drc_bufs3972(mul_7_27_n_55 ,mul_7_27_n_53);
  not mul_7_27_drc_bufs3973(mul_7_27_n_54 ,mul_7_27_n_53);
  not mul_7_27_drc_bufs3974(mul_7_27_n_53 ,mul_7_27_n_456);
  not mul_7_27_drc_bufs3976(mul_7_27_n_52 ,mul_7_27_n_50);
  not mul_7_27_drc_bufs3977(mul_7_27_n_51 ,mul_7_27_n_50);
  not mul_7_27_drc_bufs3978(mul_7_27_n_50 ,mul_7_27_n_254);
  not mul_7_27_drc_bufs3980(mul_7_27_n_49 ,mul_7_27_n_47);
  not mul_7_27_drc_bufs3981(mul_7_27_n_48 ,mul_7_27_n_47);
  not mul_7_27_drc_bufs3982(mul_7_27_n_47 ,mul_7_27_n_159);
  not mul_7_27_drc_bufs3984(mul_7_27_n_46 ,mul_7_27_n_44);
  not mul_7_27_drc_bufs3985(mul_7_27_n_45 ,mul_7_27_n_44);
  not mul_7_27_drc_bufs3986(mul_7_27_n_44 ,mul_7_27_n_161);
  not mul_7_27_drc_bufs3988(mul_7_27_n_43 ,mul_7_27_n_41);
  not mul_7_27_drc_bufs3989(mul_7_27_n_42 ,mul_7_27_n_41);
  not mul_7_27_drc_bufs3990(mul_7_27_n_41 ,mul_7_27_n_159);
  not mul_7_27_drc_bufs3992(mul_7_27_n_40 ,mul_7_27_n_38);
  not mul_7_27_drc_bufs3993(mul_7_27_n_39 ,mul_7_27_n_38);
  not mul_7_27_drc_bufs3994(mul_7_27_n_38 ,mul_7_27_n_161);
  not mul_7_27_drc_bufs3996(mul_7_27_n_37 ,mul_7_27_n_35);
  not mul_7_27_drc_bufs3997(mul_7_27_n_36 ,mul_7_27_n_35);
  not mul_7_27_drc_bufs3998(mul_7_27_n_35 ,mul_7_27_n_156);
  not mul_7_27_drc_bufs4000(mul_7_27_n_34 ,mul_7_27_n_32);
  not mul_7_27_drc_bufs4001(mul_7_27_n_33 ,mul_7_27_n_32);
  not mul_7_27_drc_bufs4002(mul_7_27_n_32 ,mul_7_27_n_254);
  not mul_7_27_drc_bufs4005(mul_7_27_n_31 ,mul_7_27_n_30);
  not mul_7_27_drc_bufs4006(mul_7_27_n_30 ,mul_7_27_n_157);
  not mul_7_27_drc_bufs4008(mul_7_27_n_29 ,mul_7_27_n_27);
  not mul_7_27_drc_bufs4009(mul_7_27_n_28 ,mul_7_27_n_27);
  not mul_7_27_drc_bufs4010(mul_7_27_n_27 ,mul_7_27_n_222);
  not mul_7_27_drc_bufs4012(mul_7_27_n_26 ,mul_7_27_n_24);
  not mul_7_27_drc_bufs4013(mul_7_27_n_25 ,mul_7_27_n_24);
  not mul_7_27_drc_bufs4014(mul_7_27_n_24 ,mul_7_27_n_220);
  not mul_7_27_drc_bufs4016(mul_7_27_n_23 ,mul_7_27_n_21);
  not mul_7_27_drc_bufs4017(mul_7_27_n_22 ,mul_7_27_n_21);
  not mul_7_27_drc_bufs4018(mul_7_27_n_21 ,mul_7_27_n_223);
  not mul_7_27_drc_bufs4020(mul_7_27_n_20 ,mul_7_27_n_18);
  not mul_7_27_drc_bufs4021(mul_7_27_n_19 ,mul_7_27_n_18);
  not mul_7_27_drc_bufs4022(mul_7_27_n_18 ,mul_7_27_n_220);
  not mul_7_27_drc_bufs4024(mul_7_27_n_17 ,mul_7_27_n_15);
  not mul_7_27_drc_bufs4025(mul_7_27_n_16 ,mul_7_27_n_15);
  not mul_7_27_drc_bufs4026(mul_7_27_n_15 ,mul_7_27_n_221);
  not mul_7_27_drc_bufs4028(mul_7_27_n_14 ,mul_7_27_n_12);
  not mul_7_27_drc_bufs4029(mul_7_27_n_13 ,mul_7_27_n_12);
  not mul_7_27_drc_bufs4030(mul_7_27_n_12 ,mul_7_27_n_221);
  not mul_7_27_drc_bufs4032(mul_7_27_n_11 ,mul_7_27_n_9);
  not mul_7_27_drc_bufs4033(mul_7_27_n_10 ,mul_7_27_n_9);
  not mul_7_27_drc_bufs4034(mul_7_27_n_9 ,mul_7_27_n_249);
  xor mul_7_27_g2__1705(out1[15] ,mul_7_27_n_1023 ,mul_7_27_n_993);
  xor mul_7_27_g4036__5122(out1[14] ,mul_7_27_n_1021 ,mul_7_27_n_992);
  xor mul_7_27_g4037__8246(out1[13] ,mul_7_27_n_1019 ,mul_7_27_n_991);
  xor mul_7_27_g4038__7098(mul_7_27_n_5 ,mul_7_27_n_886 ,mul_7_27_n_945);
  xor mul_7_27_g4039__6131(mul_7_27_n_4 ,mul_7_27_n_717 ,mul_7_27_n_831);
  xor mul_7_27_g4040__1881(mul_7_27_n_3 ,mul_7_27_n_741 ,mul_7_27_n_679);
  xor mul_7_27_g4041__5115(mul_7_27_n_2 ,mul_7_27_n_569 ,mul_7_27_n_272);
  xor mul_7_27_g4042__7482(mul_7_27_n_1 ,mul_7_27_n_774 ,mul_7_27_n_86);
  xnor mul_7_27_g4043__4733(mul_7_27_n_0 ,mul_7_27_n_246 ,mul_7_27_n_531);
  or mul_8_23_g1307__6161(out2[15] ,mul_8_23_n_367 ,mul_8_23_n_507);
  xnor mul_8_23_g1308__9315(out2[14] ,mul_8_23_n_506 ,mul_8_23_n_375);
  and mul_8_23_g1309__9945(mul_8_23_n_507 ,mul_8_23_n_370 ,mul_8_23_n_506);
  or mul_8_23_g1310__2883(mul_8_23_n_506 ,mul_8_23_n_419 ,mul_8_23_n_504);
  xnor mul_8_23_g1311__2346(out2[13] ,mul_8_23_n_503 ,mul_8_23_n_434);
  and mul_8_23_g1312__1666(mul_8_23_n_504 ,mul_8_23_n_429 ,mul_8_23_n_503);
  or mul_8_23_g1313__7410(mul_8_23_n_503 ,mul_8_23_n_457 ,mul_8_23_n_501);
  xnor mul_8_23_g1314__6417(out2[12] ,mul_8_23_n_500 ,mul_8_23_n_463);
  and mul_8_23_g1315__5477(mul_8_23_n_501 ,mul_8_23_n_456 ,mul_8_23_n_500);
  or mul_8_23_g1316__2398(mul_8_23_n_500 ,mul_8_23_n_472 ,mul_8_23_n_498);
  xnor mul_8_23_g1317__5107(out2[11] ,mul_8_23_n_497 ,mul_8_23_n_475);
  and mul_8_23_g1318__6260(mul_8_23_n_498 ,mul_8_23_n_471 ,mul_8_23_n_497);
  or mul_8_23_g1319__4319(mul_8_23_n_497 ,mul_8_23_n_479 ,mul_8_23_n_495);
  xnor mul_8_23_g1320__8428(out2[10] ,mul_8_23_n_494 ,mul_8_23_n_484);
  and mul_8_23_g1321__5526(mul_8_23_n_495 ,mul_8_23_n_483 ,mul_8_23_n_494);
  or mul_8_23_g1322__6783(mul_8_23_n_494 ,mul_8_23_n_482 ,mul_8_23_n_492);
  xnor mul_8_23_g1323__3680(out2[9] ,mul_8_23_n_491 ,mul_8_23_n_485);
  and mul_8_23_g1324__1617(mul_8_23_n_492 ,mul_8_23_n_481 ,mul_8_23_n_491);
  or mul_8_23_g1325__2802(mul_8_23_n_491 ,mul_8_23_n_466 ,mul_8_23_n_489);
  xnor mul_8_23_g1326__1705(out2[8] ,mul_8_23_n_488 ,mul_8_23_n_478);
  and mul_8_23_g1327__5122(mul_8_23_n_489 ,mul_8_23_n_465 ,mul_8_23_n_488);
  or mul_8_23_g1328__8246(mul_8_23_n_488 ,mul_8_23_n_473 ,mul_8_23_n_486);
  xnor mul_8_23_g1329__7098(out2[7] ,mul_8_23_n_480 ,mul_8_23_n_477);
  nor mul_8_23_g1330__6131(mul_8_23_n_486 ,mul_8_23_n_474 ,mul_8_23_n_480);
  xnor mul_8_23_g1331__1881(mul_8_23_n_485 ,mul_8_23_n_454 ,mul_8_23_n_469);
  xnor mul_8_23_g1332__5115(mul_8_23_n_484 ,mul_8_23_n_468 ,mul_8_23_n_461);
  or mul_8_23_g1333__7482(mul_8_23_n_483 ,mul_8_23_n_460 ,mul_8_23_n_467);
  and mul_8_23_g1334__4733(mul_8_23_n_482 ,mul_8_23_n_454 ,mul_8_23_n_469);
  or mul_8_23_g1335__6161(mul_8_23_n_481 ,mul_8_23_n_454 ,mul_8_23_n_469);
  and mul_8_23_g1336__9315(mul_8_23_n_480 ,mul_8_23_n_440 ,mul_8_23_n_470);
  nor mul_8_23_g1337__9945(mul_8_23_n_479 ,mul_8_23_n_461 ,mul_8_23_n_468);
  xnor mul_8_23_g1338__2883(mul_8_23_n_478 ,mul_8_23_n_462 ,mul_8_23_n_453);
  xnor mul_8_23_g1339__2346(mul_8_23_n_477 ,mul_8_23_n_445 ,mul_8_23_n_451);
  xnor mul_8_23_g1340__1666(out2[6] ,mul_8_23_n_455 ,mul_8_23_n_448);
  xnor mul_8_23_g1341__7410(mul_8_23_n_475 ,mul_8_23_n_450 ,mul_8_23_n_459);
  and mul_8_23_g1342__6417(mul_8_23_n_474 ,mul_8_23_n_445 ,mul_8_23_n_452);
  nor mul_8_23_g1343__5477(mul_8_23_n_473 ,mul_8_23_n_445 ,mul_8_23_n_452);
  nor mul_8_23_g1344__2398(mul_8_23_n_472 ,mul_8_23_n_459 ,mul_8_23_n_450);
  or mul_8_23_g1345__5107(mul_8_23_n_471 ,mul_8_23_n_458 ,mul_8_23_n_449);
  or mul_8_23_g1346__6260(mul_8_23_n_470 ,mul_8_23_n_441 ,mul_8_23_n_455);
  not mul_8_23_g1347(mul_8_23_n_467 ,mul_8_23_n_468);
  and mul_8_23_g1348__4319(mul_8_23_n_466 ,mul_8_23_n_462 ,mul_8_23_n_453);
  or mul_8_23_g1349__8428(mul_8_23_n_465 ,mul_8_23_n_462 ,mul_8_23_n_453);
  xnor mul_8_23_g1350__5526(out2[5] ,mul_8_23_n_423 ,mul_8_23_n_436);
  xnor mul_8_23_g1351__6783(mul_8_23_n_463 ,mul_8_23_n_447 ,mul_8_23_n_399);
  xnor mul_8_23_g1352__3680(mul_8_23_n_469 ,mul_8_23_n_391 ,mul_8_23_n_433);
  xnor mul_8_23_g1353__1617(mul_8_23_n_468 ,mul_8_23_n_411 ,mul_8_23_n_435);
  not mul_8_23_g1354(mul_8_23_n_460 ,mul_8_23_n_461);
  not mul_8_23_g1355(mul_8_23_n_458 ,mul_8_23_n_459);
  nor mul_8_23_g1356__2802(mul_8_23_n_457 ,mul_8_23_n_84 ,mul_8_23_n_447);
  or mul_8_23_g1357__1705(mul_8_23_n_456 ,mul_8_23_n_93 ,mul_8_23_n_446);
  or mul_8_23_g1358__5122(mul_8_23_n_462 ,mul_8_23_n_427 ,mul_8_23_n_442);
  and mul_8_23_g1359__8246(mul_8_23_n_461 ,mul_8_23_n_418 ,mul_8_23_n_444);
  and mul_8_23_g1360__7098(mul_8_23_n_459 ,mul_8_23_n_430 ,mul_8_23_n_443);
  not mul_8_23_g1361(mul_8_23_n_452 ,mul_8_23_n_451);
  not mul_8_23_g1362(mul_8_23_n_449 ,mul_8_23_n_450);
  xnor mul_8_23_g1363__6131(mul_8_23_n_448 ,mul_8_23_n_410 ,mul_8_23_n_422);
  and mul_8_23_g1364__1881(mul_8_23_n_455 ,mul_8_23_n_417 ,mul_8_23_n_439);
  or mul_8_23_g1365__5115(mul_8_23_n_454 ,mul_8_23_n_431 ,mul_8_23_n_437);
  xnor mul_8_23_g1366__7482(mul_8_23_n_453 ,mul_8_23_n_397 ,mul_8_23_n_415);
  xnor mul_8_23_g1367__4733(mul_8_23_n_451 ,mul_8_23_n_400 ,mul_8_23_n_413);
  xnor mul_8_23_g1368__6161(mul_8_23_n_450 ,mul_8_23_n_412 ,mul_8_23_n_414);
  not mul_8_23_g1369(mul_8_23_n_446 ,mul_8_23_n_447);
  or mul_8_23_g1370__9315(mul_8_23_n_444 ,mul_8_23_n_391 ,mul_8_23_n_424);
  or mul_8_23_g1371__9945(mul_8_23_n_443 ,mul_8_23_n_411 ,mul_8_23_n_432);
  nor mul_8_23_g1372__2883(mul_8_23_n_442 ,mul_8_23_n_390 ,mul_8_23_n_426);
  nor mul_8_23_g1373__2346(mul_8_23_n_441 ,mul_8_23_n_409 ,mul_8_23_n_422);
  or mul_8_23_g1374__1666(mul_8_23_n_440 ,mul_8_23_n_410 ,mul_8_23_n_421);
  and mul_8_23_g1375__7410(mul_8_23_n_447 ,mul_8_23_n_405 ,mul_8_23_n_420);
  and mul_8_23_g1376__6417(mul_8_23_n_445 ,mul_8_23_n_403 ,mul_8_23_n_425);
  or mul_8_23_g1377__5477(mul_8_23_n_439 ,mul_8_23_n_416 ,mul_8_23_n_423);
  xnor mul_8_23_g1378__2398(out2[4] ,mul_8_23_n_383 ,mul_8_23_n_392);
  nor mul_8_23_g1379__5107(mul_8_23_n_437 ,mul_8_23_n_389 ,mul_8_23_n_428);
  xnor mul_8_23_g1380__6260(mul_8_23_n_436 ,mul_8_23_n_372 ,mul_8_23_n_396);
  xnor mul_8_23_g1381__4319(mul_8_23_n_435 ,mul_8_23_n_398 ,mul_8_23_n_388);
  xnor mul_8_23_g1382__8428(mul_8_23_n_434 ,mul_8_23_n_408 ,mul_8_23_n_330);
  xnor mul_8_23_g1383__5526(mul_8_23_n_433 ,mul_8_23_n_382 ,mul_8_23_n_402);
  and mul_8_23_g1384__6783(mul_8_23_n_432 ,mul_8_23_n_388 ,mul_8_23_n_398);
  nor mul_8_23_g1385__3680(mul_8_23_n_431 ,mul_8_23_n_380 ,mul_8_23_n_397);
  or mul_8_23_g1386__1617(mul_8_23_n_430 ,mul_8_23_n_388 ,mul_8_23_n_398);
  or mul_8_23_g1387__2802(mul_8_23_n_429 ,mul_8_23_n_92 ,mul_8_23_n_407);
  and mul_8_23_g1388__1705(mul_8_23_n_428 ,mul_8_23_n_380 ,mul_8_23_n_397);
  nor mul_8_23_g1389__5122(mul_8_23_n_427 ,mul_8_23_n_358 ,mul_8_23_n_400);
  and mul_8_23_g1390__8246(mul_8_23_n_426 ,mul_8_23_n_358 ,mul_8_23_n_400);
  or mul_8_23_g1391__7098(mul_8_23_n_425 ,mul_8_23_n_318 ,mul_8_23_n_406);
  nor mul_8_23_g1392__6131(mul_8_23_n_424 ,mul_8_23_n_382 ,mul_8_23_n_401);
  not mul_8_23_g1393(mul_8_23_n_421 ,mul_8_23_n_422);
  or mul_8_23_g1394__1881(mul_8_23_n_420 ,mul_8_23_n_404 ,mul_8_23_n_412);
  nor mul_8_23_g1395__5115(mul_8_23_n_419 ,mul_8_23_n_85 ,mul_8_23_n_408);
  or mul_8_23_g1396__7482(mul_8_23_n_418 ,mul_8_23_n_381 ,mul_8_23_n_402);
  or mul_8_23_g1397__4733(mul_8_23_n_417 ,mul_8_23_n_372 ,mul_8_23_n_395);
  nor mul_8_23_g1398__6161(mul_8_23_n_416 ,mul_8_23_n_371 ,mul_8_23_n_396);
  xor mul_8_23_g1399__9315(mul_8_23_n_415 ,mul_8_23_n_389 ,mul_8_23_n_380);
  xnor mul_8_23_g1400__9945(mul_8_23_n_414 ,mul_8_23_n_378 ,mul_8_23_n_348);
  xor mul_8_23_g1401__2883(mul_8_23_n_413 ,mul_8_23_n_358 ,mul_8_23_n_390);
  and mul_8_23_g1402__2346(mul_8_23_n_423 ,mul_8_23_n_377 ,mul_8_23_n_393);
  xnor mul_8_23_g1403__1666(mul_8_23_n_422 ,mul_8_23_n_379 ,mul_8_23_n_353);
  not mul_8_23_g1404(mul_8_23_n_410 ,mul_8_23_n_409);
  not mul_8_23_g1405(mul_8_23_n_407 ,mul_8_23_n_408);
  and mul_8_23_g1406__7410(mul_8_23_n_406 ,mul_8_23_n_314 ,mul_8_23_n_379);
  or mul_8_23_g1407__6417(mul_8_23_n_405 ,mul_8_23_n_348 ,mul_8_23_n_378);
  and mul_8_23_g1408__5477(mul_8_23_n_404 ,mul_8_23_n_348 ,mul_8_23_n_378);
  or mul_8_23_g1409__2398(mul_8_23_n_403 ,mul_8_23_n_314 ,mul_8_23_n_379);
  and mul_8_23_g1410__5107(mul_8_23_n_412 ,mul_8_23_n_362 ,mul_8_23_n_386);
  and mul_8_23_g1411__6260(mul_8_23_n_411 ,mul_8_23_n_345 ,mul_8_23_n_384);
  or mul_8_23_g1412__4319(mul_8_23_n_409 ,mul_8_23_n_329 ,mul_8_23_n_385);
  and mul_8_23_g1413__8428(mul_8_23_n_408 ,mul_8_23_n_339 ,mul_8_23_n_387);
  not mul_8_23_g1414(mul_8_23_n_401 ,mul_8_23_n_402);
  not mul_8_23_g1416(mul_8_23_n_395 ,mul_8_23_n_396);
  xnor mul_8_23_g1417__5526(out2[3] ,mul_8_23_n_333 ,mul_8_23_n_351);
  or mul_8_23_g1418__6783(mul_8_23_n_393 ,mul_8_23_n_383 ,mul_8_23_n_376);
  xnor mul_8_23_g1419__3680(mul_8_23_n_392 ,mul_8_23_n_317 ,mul_8_23_n_360);
  xnor mul_8_23_g1420__1617(mul_8_23_n_402 ,mul_8_23_n_373 ,mul_8_23_n_354);
  xnor mul_8_23_g1421__2802(mul_8_23_n_400 ,mul_8_23_n_284 ,mul_8_23_n_349);
  xnor mul_8_23_g1422__1705(mul_8_23_n_399 ,mul_8_23_n_374 ,mul_8_23_n_356);
  xnor mul_8_23_g1423__5122(mul_8_23_n_398 ,mul_8_23_n_331 ,mul_8_23_n_350);
  xnor mul_8_23_g1424__8246(mul_8_23_n_397 ,mul_8_23_n_332 ,mul_8_23_n_352);
  xnor mul_8_23_g1425__7098(mul_8_23_n_396 ,mul_8_23_n_361 ,mul_8_23_n_355);
  or mul_8_23_g1426__6131(mul_8_23_n_387 ,mul_8_23_n_324 ,mul_8_23_n_374);
  or mul_8_23_g1427__1881(mul_8_23_n_386 ,mul_8_23_n_283 ,mul_8_23_n_364);
  and mul_8_23_g1428__5115(mul_8_23_n_385 ,mul_8_23_n_328 ,mul_8_23_n_361);
  or mul_8_23_g1429__7482(mul_8_23_n_384 ,mul_8_23_n_337 ,mul_8_23_n_373);
  and mul_8_23_g1430__4733(mul_8_23_n_391 ,mul_8_23_n_340 ,mul_8_23_n_363);
  and mul_8_23_g1431__6161(mul_8_23_n_390 ,mul_8_23_n_338 ,mul_8_23_n_366);
  and mul_8_23_g1432__9315(mul_8_23_n_389 ,mul_8_23_n_343 ,mul_8_23_n_368);
  and mul_8_23_g1433__9945(mul_8_23_n_388 ,mul_8_23_n_344 ,mul_8_23_n_369);
  not mul_8_23_g1434(mul_8_23_n_381 ,mul_8_23_n_382);
  or mul_8_23_g1435__2883(mul_8_23_n_377 ,mul_8_23_n_317 ,mul_8_23_n_359);
  nor mul_8_23_g1436__2346(mul_8_23_n_376 ,mul_8_23_n_316 ,mul_8_23_n_360);
  xnor mul_8_23_g1437__1666(mul_8_23_n_375 ,mul_8_23_n_116 ,mul_8_23_n_347);
  and mul_8_23_g1438__7410(mul_8_23_n_383 ,mul_8_23_n_326 ,mul_8_23_n_365);
  xnor mul_8_23_g1439__6417(mul_8_23_n_382 ,mul_8_23_n_298 ,mul_8_23_n_320);
  xor mul_8_23_g1440__5477(mul_8_23_n_380 ,mul_8_23_n_272 ,mul_8_23_n_319);
  xnor mul_8_23_g1441__2398(mul_8_23_n_379 ,mul_8_23_n_299 ,mul_8_23_n_321);
  xnor mul_8_23_g1442__5107(mul_8_23_n_378 ,mul_8_23_n_303 ,mul_8_23_n_322);
  not mul_8_23_g1443(mul_8_23_n_371 ,mul_8_23_n_372);
  or mul_8_23_g1444__6260(mul_8_23_n_370 ,mul_8_23_n_115 ,mul_8_23_n_346);
  or mul_8_23_g1445__4319(mul_8_23_n_369 ,mul_8_23_n_285 ,mul_8_23_n_342);
  or mul_8_23_g1446__8428(mul_8_23_n_368 ,mul_8_23_n_284 ,mul_8_23_n_341);
  nor mul_8_23_g1447__5526(mul_8_23_n_367 ,mul_8_23_n_116 ,mul_8_23_n_347);
  or mul_8_23_g1448__6783(mul_8_23_n_366 ,mul_8_23_n_286 ,mul_8_23_n_336);
  or mul_8_23_g1449__3680(mul_8_23_n_365 ,mul_8_23_n_333 ,mul_8_23_n_323);
  and mul_8_23_g1450__1617(mul_8_23_n_364 ,mul_8_23_n_292 ,mul_8_23_n_331);
  or mul_8_23_g1451__2802(mul_8_23_n_363 ,mul_8_23_n_332 ,mul_8_23_n_334);
  or mul_8_23_g1452__1705(mul_8_23_n_362 ,mul_8_23_n_292 ,mul_8_23_n_331);
  and mul_8_23_g1453__5122(mul_8_23_n_374 ,mul_8_23_n_307 ,mul_8_23_n_325);
  and mul_8_23_g1454__8246(mul_8_23_n_373 ,mul_8_23_n_313 ,mul_8_23_n_335);
  and mul_8_23_g1455__7098(mul_8_23_n_372 ,mul_8_23_n_276 ,mul_8_23_n_327);
  not mul_8_23_g1456(mul_8_23_n_359 ,mul_8_23_n_360);
  xnor mul_8_23_g1457__6131(out2[2] ,mul_8_23_n_222 ,mul_8_23_n_288);
  xnor mul_8_23_g1458__1881(mul_8_23_n_356 ,mul_8_23_n_297 ,mul_8_23_n_279);
  xnor mul_8_23_g1459__5115(mul_8_23_n_355 ,mul_8_23_n_295 ,mul_8_23_n_281);
  xnor mul_8_23_g1460__7482(mul_8_23_n_354 ,mul_8_23_n_301 ,mul_8_23_n_315);
  xor mul_8_23_g1461__4733(mul_8_23_n_353 ,mul_8_23_n_314 ,mul_8_23_n_318);
  xnor mul_8_23_g1462__6161(mul_8_23_n_352 ,mul_8_23_n_291 ,mul_8_23_n_300);
  xnor mul_8_23_g1463__9315(mul_8_23_n_351 ,mul_8_23_n_203 ,mul_8_23_n_290);
  xnor mul_8_23_g1464__9945(mul_8_23_n_350 ,mul_8_23_n_292 ,mul_8_23_n_283);
  xnor mul_8_23_g1465__2883(mul_8_23_n_349 ,mul_8_23_n_293 ,mul_8_23_n_296);
  xnor mul_8_23_g1466__2346(mul_8_23_n_361 ,mul_8_23_n_205 ,mul_8_23_n_287);
  xnor mul_8_23_g1467__1666(mul_8_23_n_360 ,mul_8_23_n_302 ,mul_8_23_n_304);
  xor mul_8_23_g1468__7410(mul_8_23_n_358 ,mul_8_23_n_282 ,mul_8_23_n_305);
  not mul_8_23_g1469(mul_8_23_n_346 ,mul_8_23_n_347);
  or mul_8_23_g1470__6417(mul_8_23_n_345 ,mul_8_23_n_315 ,mul_8_23_n_301);
  or mul_8_23_g1471__5477(mul_8_23_n_344 ,mul_8_23_n_221 ,mul_8_23_n_298);
  or mul_8_23_g1472__2398(mul_8_23_n_343 ,mul_8_23_n_296 ,mul_8_23_n_293);
  and mul_8_23_g1473__5107(mul_8_23_n_342 ,mul_8_23_n_221 ,mul_8_23_n_298);
  and mul_8_23_g1474__6260(mul_8_23_n_341 ,mul_8_23_n_296 ,mul_8_23_n_293);
  or mul_8_23_g1475__4319(mul_8_23_n_340 ,mul_8_23_n_300 ,mul_8_23_n_291);
  or mul_8_23_g1476__8428(mul_8_23_n_339 ,mul_8_23_n_279 ,mul_8_23_n_297);
  or mul_8_23_g1477__5526(mul_8_23_n_338 ,mul_8_23_n_5 ,mul_8_23_n_299);
  and mul_8_23_g1478__6783(mul_8_23_n_337 ,mul_8_23_n_315 ,mul_8_23_n_301);
  and mul_8_23_g1479__3680(mul_8_23_n_336 ,mul_8_23_n_5 ,mul_8_23_n_299);
  or mul_8_23_g1480__1617(mul_8_23_n_335 ,mul_8_23_n_275 ,mul_8_23_n_312);
  and mul_8_23_g1481__2802(mul_8_23_n_334 ,mul_8_23_n_300 ,mul_8_23_n_291);
  and mul_8_23_g1482__1705(mul_8_23_n_348 ,mul_8_23_n_198 ,mul_8_23_n_310);
  and mul_8_23_g1483__5122(mul_8_23_n_347 ,mul_8_23_n_184 ,mul_8_23_n_308);
  nor mul_8_23_g1485__8246(mul_8_23_n_329 ,mul_8_23_n_281 ,mul_8_23_n_295);
  or mul_8_23_g1486__7098(mul_8_23_n_328 ,mul_8_23_n_280 ,mul_8_23_n_294);
  or mul_8_23_g1487__6131(mul_8_23_n_327 ,mul_8_23_n_269 ,mul_8_23_n_302);
  or mul_8_23_g1488__1881(mul_8_23_n_326 ,mul_8_23_n_202 ,mul_8_23_n_290);
  or mul_8_23_g1489__5115(mul_8_23_n_325 ,mul_8_23_n_309 ,mul_8_23_n_303);
  and mul_8_23_g1490__7482(mul_8_23_n_324 ,mul_8_23_n_279 ,mul_8_23_n_297);
  nor mul_8_23_g1491__4733(mul_8_23_n_323 ,mul_8_23_n_203 ,mul_8_23_n_289);
  xnor mul_8_23_g1492__6161(mul_8_23_n_322 ,mul_8_23_n_158 ,mul_8_23_n_270);
  xnor mul_8_23_g1493__9315(mul_8_23_n_321 ,mul_8_23_n_286 ,mul_8_23_n_5);
  xor mul_8_23_g1494__9945(mul_8_23_n_320 ,mul_8_23_n_221 ,mul_8_23_n_285);
  xnor mul_8_23_g1495__2883(mul_8_23_n_319 ,mul_8_23_n_201 ,mul_8_23_n_275);
  and mul_8_23_g1496__2346(mul_8_23_n_333 ,mul_8_23_n_264 ,mul_8_23_n_306);
  and mul_8_23_g1497__1666(mul_8_23_n_332 ,mul_8_23_n_267 ,mul_8_23_n_311);
  xnor mul_8_23_g1498__7410(mul_8_23_n_331 ,mul_8_23_n_274 ,mul_8_23_n_235);
  xnor mul_8_23_g1499__6417(mul_8_23_n_330 ,mul_8_23_n_273 ,mul_8_23_n_241);
  not mul_8_23_g1500(mul_8_23_n_316 ,mul_8_23_n_317);
  or mul_8_23_g1501__5477(mul_8_23_n_313 ,mul_8_23_n_200 ,mul_8_23_n_272);
  nor mul_8_23_g1502__2398(mul_8_23_n_312 ,mul_8_23_n_201 ,mul_8_23_n_271);
  or mul_8_23_g1503__5107(mul_8_23_n_311 ,mul_8_23_n_282 ,mul_8_23_n_277);
  or mul_8_23_g1504__6260(mul_8_23_n_310 ,mul_8_23_n_195 ,mul_8_23_n_274);
  and mul_8_23_g1505__4319(mul_8_23_n_309 ,mul_8_23_n_158 ,mul_8_23_n_270);
  or mul_8_23_g1506__8428(mul_8_23_n_308 ,mul_8_23_n_209 ,mul_8_23_n_273);
  or mul_8_23_g1507__5526(mul_8_23_n_307 ,mul_8_23_n_158 ,mul_8_23_n_270);
  xnor mul_8_23_g1509__6783(mul_8_23_n_305 ,mul_8_23_n_227 ,mul_8_23_n_7);
  xnor mul_8_23_g1510__3680(mul_8_23_n_304 ,mul_8_23_n_224 ,mul_8_23_n_3);
  and mul_8_23_g1511__1617(mul_8_23_n_318 ,mul_8_23_n_263 ,mul_8_23_n_266);
  and mul_8_23_g1512__2802(mul_8_23_n_317 ,mul_8_23_n_193 ,mul_8_23_n_265);
  and mul_8_23_g1513__1705(mul_8_23_n_315 ,mul_8_23_n_196 ,mul_8_23_n_278);
  xor mul_8_23_g1514__5122(mul_8_23_n_314 ,mul_8_23_n_228 ,mul_8_23_n_232);
  not mul_8_23_g1515(mul_8_23_n_294 ,mul_8_23_n_295);
  not mul_8_23_g1516(mul_8_23_n_289 ,mul_8_23_n_290);
  xnor mul_8_23_g1517__8246(mul_8_23_n_288 ,mul_8_23_n_122 ,mul_8_23_n_244);
  xnor mul_8_23_g1518__7098(mul_8_23_n_287 ,mul_8_23_n_148 ,mul_8_23_n_4);
  xnor mul_8_23_g1519__6131(mul_8_23_n_303 ,mul_8_23_n_130 ,mul_8_23_n_247);
  xnor mul_8_23_g1520__1881(mul_8_23_n_302 ,mul_8_23_n_150 ,mul_8_23_n_236);
  xnor mul_8_23_g1521__5115(mul_8_23_n_301 ,mul_8_23_n_173 ,mul_8_23_n_242);
  xnor mul_8_23_g1522__7482(mul_8_23_n_300 ,mul_8_23_n_118 ,mul_8_23_n_233);
  xnor mul_8_23_g1523__4733(mul_8_23_n_299 ,mul_8_23_n_159 ,mul_8_23_n_234);
  xnor mul_8_23_g1524__6161(mul_8_23_n_298 ,mul_8_23_n_141 ,mul_8_23_n_240);
  xnor mul_8_23_g1525__9315(mul_8_23_n_297 ,mul_8_23_n_142 ,mul_8_23_n_231);
  xnor mul_8_23_g1526__9945(mul_8_23_n_296 ,mul_8_23_n_117 ,mul_8_23_n_239);
  xnor mul_8_23_g1527__2883(mul_8_23_n_295 ,mul_8_23_n_155 ,mul_8_23_n_230);
  xnor mul_8_23_g1528__2346(mul_8_23_n_293 ,mul_8_23_n_162 ,mul_8_23_n_238);
  xnor mul_8_23_g1529__1666(mul_8_23_n_292 ,mul_8_23_n_140 ,mul_8_23_n_237);
  xnor mul_8_23_g1530__7410(mul_8_23_n_291 ,mul_8_23_n_245 ,mul_8_23_n_248);
  xnor mul_8_23_g1531__6417(mul_8_23_n_290 ,mul_8_23_n_6 ,mul_8_23_n_246);
  not mul_8_23_g1532(mul_8_23_n_280 ,mul_8_23_n_281);
  or mul_8_23_g1533__5477(mul_8_23_n_278 ,mul_8_23_n_211 ,mul_8_23_n_245);
  nor mul_8_23_g1534__2398(mul_8_23_n_277 ,mul_8_23_n_227 ,mul_8_23_n_243);
  or mul_8_23_g1535__5107(mul_8_23_n_276 ,mul_8_23_n_225 ,mul_8_23_n_3);
  and mul_8_23_g1536__6260(mul_8_23_n_286 ,mul_8_23_n_218 ,mul_8_23_n_258);
  and mul_8_23_g1537__4319(mul_8_23_n_285 ,mul_8_23_n_194 ,mul_8_23_n_261);
  and mul_8_23_g1538__8428(mul_8_23_n_284 ,mul_8_23_n_212 ,mul_8_23_n_260);
  and mul_8_23_g1539__5526(mul_8_23_n_283 ,mul_8_23_n_197 ,mul_8_23_n_250);
  and mul_8_23_g1540__6783(mul_8_23_n_282 ,mul_8_23_n_219 ,mul_8_23_n_254);
  and mul_8_23_g1541__3680(mul_8_23_n_281 ,mul_8_23_n_190 ,mul_8_23_n_251);
  and mul_8_23_g1542__1617(mul_8_23_n_279 ,mul_8_23_n_183 ,mul_8_23_n_259);
  not mul_8_23_g1543(mul_8_23_n_271 ,mul_8_23_n_272);
  and mul_8_23_g1544__2802(mul_8_23_n_269 ,mul_8_23_n_225 ,mul_8_23_n_3);
  or mul_8_23_g1546__1705(mul_8_23_n_267 ,mul_8_23_n_226 ,mul_8_23_n_7);
  or mul_8_23_g1547__5122(mul_8_23_n_266 ,mul_8_23_n_253 ,mul_8_23_n_4);
  or mul_8_23_g1548__8246(mul_8_23_n_265 ,mul_8_23_n_220 ,mul_8_23_n_6);
  or mul_8_23_g1549__7098(mul_8_23_n_264 ,mul_8_23_n_122 ,mul_8_23_n_244);
  and mul_8_23_g1550__6131(mul_8_23_n_275 ,mul_8_23_n_188 ,mul_8_23_n_252);
  and mul_8_23_g1551__1881(mul_8_23_n_274 ,mul_8_23_n_207 ,mul_8_23_n_257);
  and mul_8_23_g1552__5115(mul_8_23_n_273 ,mul_8_23_n_186 ,mul_8_23_n_262);
  and mul_8_23_g1553__7482(mul_8_23_n_272 ,mul_8_23_n_214 ,mul_8_23_n_255);
  and mul_8_23_g1554__4733(mul_8_23_n_270 ,mul_8_23_n_187 ,mul_8_23_n_256);
  or mul_8_23_g1555__6161(mul_8_23_n_263 ,mul_8_23_n_148 ,mul_8_23_n_204);
  or mul_8_23_g1556__9315(mul_8_23_n_262 ,mul_8_23_n_142 ,mul_8_23_n_217);
  or mul_8_23_g1557__9945(mul_8_23_n_261 ,mul_8_23_n_175 ,mul_8_23_n_213);
  or mul_8_23_g1558__2883(mul_8_23_n_260 ,mul_8_23_n_206 ,mul_8_23_n_229);
  or mul_8_23_g1559__2346(mul_8_23_n_259 ,mul_8_23_n_130 ,mul_8_23_n_182);
  or mul_8_23_g1560__1666(mul_8_23_n_258 ,mul_8_23_n_138 ,mul_8_23_n_191);
  or mul_8_23_g1561__7410(mul_8_23_n_257 ,mul_8_23_n_141 ,mul_8_23_n_192);
  or mul_8_23_g1562__6417(mul_8_23_n_256 ,mul_8_23_n_140 ,mul_8_23_n_185);
  or mul_8_23_g1563__5477(mul_8_23_n_255 ,mul_8_23_n_162 ,mul_8_23_n_189);
  or mul_8_23_g1564__2398(mul_8_23_n_254 ,mul_8_23_n_174 ,mul_8_23_n_208);
  nor mul_8_23_g1565__5107(mul_8_23_n_253 ,mul_8_23_n_147 ,mul_8_23_n_205);
  or mul_8_23_g1566__6260(mul_8_23_n_252 ,mul_8_23_n_163 ,mul_8_23_n_199);
  or mul_8_23_g1567__4319(mul_8_23_n_251 ,mul_8_23_n_136 ,mul_8_23_n_215);
  or mul_8_23_g1568__8428(mul_8_23_n_250 ,mul_8_23_n_173 ,mul_8_23_n_210);
  and mul_8_23_g1569__5526(out2[1] ,mul_8_23_n_216 ,mul_8_23_n_223);
  xnor mul_8_23_g1570__6783(mul_8_23_n_248 ,mul_8_23_n_125 ,mul_8_23_n_114);
  xnor mul_8_23_g1571__3680(mul_8_23_n_247 ,mul_8_23_n_120 ,mul_8_23_n_143);
  xnor mul_8_23_g1572__1617(mul_8_23_n_246 ,mul_8_23_n_152 ,mul_8_23_n_113);
  not mul_8_23_g1574(mul_8_23_n_243 ,mul_8_23_n_7);
  xnor mul_8_23_g1575__2802(mul_8_23_n_242 ,mul_8_23_n_154 ,mul_8_23_n_153);
  xnor mul_8_23_g1576__1705(mul_8_23_n_241 ,mul_8_23_n_145 ,mul_8_23_n_124);
  xnor mul_8_23_g1577__5122(mul_8_23_n_240 ,mul_8_23_n_157 ,mul_8_23_n_128);
  xnor mul_8_23_g1578__8246(mul_8_23_n_239 ,mul_8_23_n_163 ,mul_8_23_n_127);
  xnor mul_8_23_g1579__7098(mul_8_23_n_238 ,mul_8_23_n_149 ,mul_8_23_n_126);
  xnor mul_8_23_g1580__6131(mul_8_23_n_237 ,mul_8_23_n_161 ,mul_8_23_n_111);
  xnor mul_8_23_g1581__1881(mul_8_23_n_236 ,mul_8_23_n_136 ,mul_8_23_n_123);
  xnor mul_8_23_g1582__5115(mul_8_23_n_235 ,mul_8_23_n_121 ,mul_8_23_n_146);
  xnor mul_8_23_g1583__7482(mul_8_23_n_234 ,mul_8_23_n_174 ,mul_8_23_n_160);
  xnor mul_8_23_g1584__4733(mul_8_23_n_233 ,mul_8_23_n_175 ,mul_8_23_n_119);
  xnor mul_8_23_g1585__6161(mul_8_23_n_232 ,mul_8_23_n_156 ,mul_8_23_n_112);
  xnor mul_8_23_g1586__9315(mul_8_23_n_231 ,mul_8_23_n_151 ,mul_8_23_n_129);
  xnor mul_8_23_g1587__9945(mul_8_23_n_230 ,mul_8_23_n_138 ,mul_8_23_n_144);
  xnor mul_8_23_g1588__2883(mul_8_23_n_245 ,mul_8_23_n_137 ,mul_8_23_n_166);
  xnor mul_8_23_g1592__2346(mul_8_23_n_244 ,mul_8_23_n_178 ,mul_8_23_n_164);
  not mul_8_23_g1594(mul_8_23_n_229 ,mul_8_23_n_228);
  not mul_8_23_g1595(mul_8_23_n_226 ,mul_8_23_n_227);
  not mul_8_23_g1596(mul_8_23_n_225 ,mul_8_23_n_224);
  not mul_8_23_g1597(mul_8_23_n_223 ,mul_8_23_n_222);
  and mul_8_23_g1598__1666(mul_8_23_n_220 ,mul_8_23_n_152 ,mul_8_23_n_113);
  or mul_8_23_g1599__7410(mul_8_23_n_219 ,mul_8_23_n_160 ,mul_8_23_n_159);
  or mul_8_23_g1600__6417(mul_8_23_n_218 ,mul_8_23_n_144 ,mul_8_23_n_155);
  and mul_8_23_g1601__5477(mul_8_23_n_217 ,mul_8_23_n_151 ,mul_8_23_n_129);
  or mul_8_23_g1602__2398(mul_8_23_n_216 ,mul_8_23_n_181 ,mul_8_23_n_180);
  and mul_8_23_g1603__5107(mul_8_23_n_215 ,mul_8_23_n_123 ,mul_8_23_n_150);
  or mul_8_23_g1604__6260(mul_8_23_n_214 ,mul_8_23_n_149 ,mul_8_23_n_126);
  and mul_8_23_g1605__4319(mul_8_23_n_213 ,mul_8_23_n_119 ,mul_8_23_n_118);
  or mul_8_23_g1606__8428(mul_8_23_n_212 ,mul_8_23_n_156 ,mul_8_23_n_112);
  and mul_8_23_g1607__5526(mul_8_23_n_211 ,mul_8_23_n_125 ,mul_8_23_n_114);
  and mul_8_23_g1608__6783(mul_8_23_n_210 ,mul_8_23_n_154 ,mul_8_23_n_153);
  and mul_8_23_g1609__3680(mul_8_23_n_209 ,mul_8_23_n_145 ,mul_8_23_n_124);
  and mul_8_23_g1610__1617(mul_8_23_n_208 ,mul_8_23_n_160 ,mul_8_23_n_159);
  or mul_8_23_g1611__2802(mul_8_23_n_207 ,mul_8_23_n_157 ,mul_8_23_n_128);
  and mul_8_23_g1612__1705(mul_8_23_n_206 ,mul_8_23_n_156 ,mul_8_23_n_112);
  and mul_8_23_g1613__5122(mul_8_23_n_228 ,mul_8_23_n_132 ,mul_8_23_n_170);
  and mul_8_23_g1614__8246(mul_8_23_n_227 ,mul_8_23_n_172 ,mul_8_23_n_133);
  and mul_8_23_g1615__7098(mul_8_23_n_224 ,mul_8_23_n_168 ,mul_8_23_n_134);
  and mul_8_23_g1616__6131(mul_8_23_n_222 ,mul_8_23_n_181 ,mul_8_23_n_180);
  or mul_8_23_g1617__1881(mul_8_23_n_221 ,mul_8_23_n_137 ,mul_8_23_n_166);
  not mul_8_23_g1618(mul_8_23_n_204 ,mul_8_23_n_205);
  not mul_8_23_g1619(mul_8_23_n_202 ,mul_8_23_n_203);
  not mul_8_23_g1620(mul_8_23_n_200 ,mul_8_23_n_201);
  and mul_8_23_g1621__5115(mul_8_23_n_199 ,mul_8_23_n_117 ,mul_8_23_n_127);
  or mul_8_23_g1622__7482(mul_8_23_n_198 ,mul_8_23_n_121 ,mul_8_23_n_146);
  or mul_8_23_g1623__4733(mul_8_23_n_197 ,mul_8_23_n_154 ,mul_8_23_n_153);
  or mul_8_23_g1624__6161(mul_8_23_n_196 ,mul_8_23_n_125 ,mul_8_23_n_114);
  and mul_8_23_g1625(mul_8_23_n_195 ,mul_8_23_n_121 ,mul_8_23_n_146);
  or mul_8_23_g1626(mul_8_23_n_194 ,mul_8_23_n_119 ,mul_8_23_n_118);
  or mul_8_23_g1627(mul_8_23_n_193 ,mul_8_23_n_152 ,mul_8_23_n_113);
  and mul_8_23_g1628(mul_8_23_n_192 ,mul_8_23_n_157 ,mul_8_23_n_128);
  and mul_8_23_g1629(mul_8_23_n_191 ,mul_8_23_n_144 ,mul_8_23_n_155);
  or mul_8_23_g1630(mul_8_23_n_190 ,mul_8_23_n_123 ,mul_8_23_n_150);
  and mul_8_23_g1631(mul_8_23_n_189 ,mul_8_23_n_149 ,mul_8_23_n_126);
  or mul_8_23_g1632(mul_8_23_n_188 ,mul_8_23_n_117 ,mul_8_23_n_127);
  or mul_8_23_g1633(mul_8_23_n_187 ,mul_8_23_n_161 ,mul_8_23_n_111);
  or mul_8_23_g1634(mul_8_23_n_186 ,mul_8_23_n_151 ,mul_8_23_n_129);
  and mul_8_23_g1635(mul_8_23_n_185 ,mul_8_23_n_161 ,mul_8_23_n_111);
  or mul_8_23_g1636(mul_8_23_n_184 ,mul_8_23_n_145 ,mul_8_23_n_124);
  or mul_8_23_g1637(mul_8_23_n_183 ,mul_8_23_n_120 ,mul_8_23_n_143);
  and mul_8_23_g1638(mul_8_23_n_182 ,mul_8_23_n_120 ,mul_8_23_n_143);
  and mul_8_23_g1639(mul_8_23_n_205 ,mul_8_23_n_131 ,mul_8_23_n_177);
  and mul_8_23_g1640(mul_8_23_n_203 ,mul_8_23_n_179 ,mul_8_23_n_165);
  and mul_8_23_g1641(mul_8_23_n_201 ,mul_8_23_n_139 ,mul_8_23_n_135);
  not mul_8_23_g1642(mul_8_23_n_179 ,mul_8_23_n_178);
  not mul_8_23_g1643(mul_8_23_n_177 ,mul_8_23_n_176);
  not mul_8_23_g1644(mul_8_23_n_172 ,mul_8_23_n_171);
  not mul_8_23_g1645(mul_8_23_n_170 ,mul_8_23_n_169);
  not mul_8_23_g1646(mul_8_23_n_168 ,mul_8_23_n_167);
  not mul_8_23_g1647(mul_8_23_n_165 ,mul_8_23_n_164);
  not mul_8_23_g1648(mul_8_23_n_147 ,mul_8_23_n_148);
  and mul_8_23_g1649(mul_8_23_n_181 ,in1[0] ,in3[1]);
  and mul_8_23_g1650(mul_8_23_n_180 ,in1[1] ,in3[0]);
  or mul_8_23_g1651(mul_8_23_n_178 ,mul_8_23_n_29 ,mul_8_23_n_46);
  or mul_8_23_g1652(mul_8_23_n_176 ,mul_8_23_n_19 ,mul_8_23_n_90);
  or mul_8_23_g1653(mul_8_23_n_175 ,mul_8_23_n_22 ,mul_8_23_n_31);
  or mul_8_23_g1654(mul_8_23_n_174 ,mul_8_23_n_79 ,mul_8_23_n_76);
  or mul_8_23_g1655(mul_8_23_n_173 ,mul_8_23_n_68 ,mul_8_23_n_37);
  or mul_8_23_g1656(mul_8_23_n_171 ,mul_8_23_n_43 ,mul_8_23_n_98);
  or mul_8_23_g1657(mul_8_23_n_169 ,mul_8_23_n_40 ,mul_8_23_n_100);
  or mul_8_23_g1658(mul_8_23_n_167 ,mul_8_23_n_64 ,mul_8_23_n_88);
  or mul_8_23_g1659(mul_8_23_n_166 ,mul_8_23_n_26 ,mul_8_23_n_88);
  or mul_8_23_g1660(mul_8_23_n_164 ,mul_8_23_n_65 ,mul_8_23_n_90);
  or mul_8_23_g1661(mul_8_23_n_163 ,mul_8_23_n_74 ,mul_8_23_n_15);
  or mul_8_23_g1662(mul_8_23_n_162 ,mul_8_23_n_28 ,mul_8_23_n_61);
  or mul_8_23_g1663(mul_8_23_n_161 ,mul_8_23_n_10 ,mul_8_23_n_70);
  or mul_8_23_g1664(mul_8_23_n_160 ,mul_8_23_n_24 ,mul_8_23_n_82);
  or mul_8_23_g1665(mul_8_23_n_159 ,mul_8_23_n_68 ,mul_8_23_n_34);
  or mul_8_23_g1666(mul_8_23_n_158 ,mul_8_23_n_41 ,mul_8_23_n_55);
  or mul_8_23_g1667(mul_8_23_n_157 ,mul_8_23_n_105 ,mul_8_23_n_56);
  or mul_8_23_g1668(mul_8_23_n_156 ,mul_8_23_n_74 ,mul_8_23_n_62);
  or mul_8_23_g1669(mul_8_23_n_155 ,mul_8_23_n_21 ,mul_8_23_n_35);
  or mul_8_23_g1670(mul_8_23_n_154 ,mul_8_23_n_17 ,mul_8_23_n_49);
  or mul_8_23_g1671(mul_8_23_n_153 ,mul_8_23_n_13 ,mul_8_23_n_47);
  or mul_8_23_g1672(mul_8_23_n_152 ,mul_8_23_n_29 ,mul_8_23_n_50);
  or mul_8_23_g1673(mul_8_23_n_151 ,mul_8_23_n_99 ,mul_8_23_n_55);
  or mul_8_23_g1674(mul_8_23_n_150 ,mul_8_23_n_80 ,mul_8_23_n_34);
  or mul_8_23_g1675(mul_8_23_n_149 ,mul_8_23_n_64 ,mul_8_23_n_38);
  or mul_8_23_g1676(mul_8_23_n_148 ,mul_8_23_n_73 ,mul_8_23_n_32);
  or mul_8_23_g1677(mul_8_23_n_146 ,mul_8_23_n_44 ,mul_8_23_n_37);
  or mul_8_23_g1678(mul_8_23_n_145 ,mul_8_23_n_9 ,mul_8_23_n_59);
  or mul_8_23_g1679(mul_8_23_n_144 ,mul_8_23_n_79 ,mul_8_23_n_83);
  or mul_8_23_g1680(mul_8_23_n_143 ,mul_8_23_n_12 ,mul_8_23_n_71);
  not mul_8_23_g1687(mul_8_23_n_116 ,mul_8_23_n_115);
  nor mul_8_23_g1688(mul_8_23_n_110 ,mul_8_23_n_100 ,mul_8_23_n_1);
  or mul_8_23_g1689(mul_8_23_n_142 ,mul_8_23_n_40 ,mul_8_23_n_59);
  or mul_8_23_g1690(mul_8_23_n_141 ,mul_8_23_n_65 ,mul_8_23_n_95);
  or mul_8_23_g1691(mul_8_23_n_140 ,mul_8_23_n_94 ,mul_8_23_n_61);
  and mul_8_23_g1692(mul_8_23_n_139 ,in1[6] ,in3[1]);
  or mul_8_23_g1693(mul_8_23_n_138 ,mul_8_23_n_53 ,mul_8_23_n_77);
  or mul_8_23_g1694(mul_8_23_n_137 ,mul_8_23_n_17 ,mul_8_23_n_46);
  or mul_8_23_g1695(mul_8_23_n_136 ,mul_8_23_n_73 ,mul_8_23_n_70);
  and mul_8_23_g1696(mul_8_23_n_135 ,in1[7] ,in3[0]);
  and mul_8_23_g1697(mul_8_23_n_134 ,in1[3] ,in3[0]);
  and mul_8_23_g1698(mul_8_23_n_133 ,in1[6] ,in3[0]);
  and mul_8_23_g1699(mul_8_23_n_132 ,in1[4] ,in3[1]);
  and mul_8_23_g1700(mul_8_23_n_131 ,in1[3] ,in3[1]);
  or mul_8_23_g1701(mul_8_23_n_130 ,mul_8_23_n_67 ,mul_8_23_n_58);
  or mul_8_23_g1702(mul_8_23_n_129 ,mul_8_23_n_102 ,mul_8_23_n_31);
  or mul_8_23_g1703(mul_8_23_n_128 ,mul_8_23_n_43 ,mul_8_23_n_76);
  or mul_8_23_g1704(mul_8_23_n_127 ,mul_8_23_n_19 ,mul_8_23_n_49);
  or mul_8_23_g1705(mul_8_23_n_126 ,mul_8_23_n_41 ,mul_8_23_n_35);
  or mul_8_23_g1706(mul_8_23_n_125 ,mul_8_23_n_53 ,mul_8_23_n_15);
  or mul_8_23_g1707(mul_8_23_n_124 ,mul_8_23_n_13 ,mul_8_23_n_56);
  or mul_8_23_g1708(mul_8_23_n_123 ,mul_8_23_n_101 ,mul_8_23_n_82);
  or mul_8_23_g1709(mul_8_23_n_122 ,mul_8_23_n_52 ,mul_8_23_n_98);
  or mul_8_23_g1710(mul_8_23_n_121 ,mul_8_23_n_24 ,mul_8_23_n_58);
  or mul_8_23_g1711(mul_8_23_n_120 ,mul_8_23_n_10 ,mul_8_23_n_38);
  or mul_8_23_g1712(mul_8_23_n_119 ,mul_8_23_n_67 ,mul_8_23_n_71);
  or mul_8_23_g1713(mul_8_23_n_118 ,mul_8_23_n_44 ,mul_8_23_n_50);
  or mul_8_23_g1714(mul_8_23_n_117 ,mul_8_23_n_22 ,mul_8_23_n_77);
  and mul_8_23_g1715(mul_8_23_n_115 ,in1[7] ,in3[7]);
  or mul_8_23_g1716(mul_8_23_n_114 ,mul_8_23_n_80 ,mul_8_23_n_62);
  or mul_8_23_g1717(mul_8_23_n_113 ,mul_8_23_n_28 ,mul_8_23_n_47);
  or mul_8_23_g1718(mul_8_23_n_112 ,mul_8_23_n_52 ,mul_8_23_n_32);
  or mul_8_23_g1719(mul_8_23_n_111 ,mul_8_23_n_26 ,mul_8_23_n_83);
  not mul_8_23_g1720(mul_8_23_n_109 ,in1[0]);
  not mul_8_23_g1721(mul_8_23_n_108 ,in3[3]);
  not mul_8_23_g1722(mul_8_23_n_107 ,in1[5]);
  not mul_8_23_g1723(mul_8_23_n_106 ,in3[5]);
  not mul_8_23_g1724(mul_8_23_n_105 ,in1[3]);
  not mul_8_23_g1725(mul_8_23_n_104 ,in1[2]);
  not mul_8_23_g1726(mul_8_23_n_103 ,in3[6]);
  not mul_8_23_g1727(mul_8_23_n_102 ,in1[7]);
  not mul_8_23_g1728(mul_8_23_n_101 ,in1[1]);
  not mul_8_23_g1729(mul_8_23_n_100 ,in3[0]);
  not mul_8_23_g1730(mul_8_23_n_99 ,in1[6]);
  not mul_8_23_g1731(mul_8_23_n_98 ,in3[1]);
  not mul_8_23_g1732(mul_8_23_n_97 ,in3[2]);
  not mul_8_23_g1733(mul_8_23_n_96 ,in3[4]);
  not mul_8_23_g1734(mul_8_23_n_95 ,in3[7]);
  not mul_8_23_g1735(mul_8_23_n_94 ,in1[4]);
  not mul_8_23_drc_bufs1770(mul_8_23_n_2 ,mul_8_23_n_91);
  not mul_8_23_drc_bufs1772(mul_8_23_n_91 ,mul_8_23_n_109);
  not mul_8_23_drc_bufs1799(mul_8_23_n_90 ,mul_8_23_n_89);
  not mul_8_23_drc_bufs1800(mul_8_23_n_89 ,mul_8_23_n_100);
  not mul_8_23_drc_bufs1803(mul_8_23_n_88 ,mul_8_23_n_87);
  not mul_8_23_drc_bufs1804(mul_8_23_n_87 ,mul_8_23_n_98);
  buf mul_8_23_drc_bufs1806(out2[0] ,mul_8_23_n_110);
  not mul_8_23_drc_bufs1808(mul_8_23_n_85 ,mul_8_23_n_92);
  not mul_8_23_drc_bufs1809(mul_8_23_n_92 ,mul_8_23_n_330);
  not mul_8_23_drc_bufs1812(mul_8_23_n_84 ,mul_8_23_n_93);
  not mul_8_23_drc_bufs1813(mul_8_23_n_93 ,mul_8_23_n_399);
  not mul_8_23_drc_bufs1815(mul_8_23_n_83 ,mul_8_23_n_81);
  not mul_8_23_drc_bufs1816(mul_8_23_n_82 ,mul_8_23_n_81);
  not mul_8_23_drc_bufs1817(mul_8_23_n_81 ,mul_8_23_n_108);
  not mul_8_23_drc_bufs1819(mul_8_23_n_80 ,mul_8_23_n_78);
  not mul_8_23_drc_bufs1820(mul_8_23_n_79 ,mul_8_23_n_78);
  not mul_8_23_drc_bufs1821(mul_8_23_n_78 ,mul_8_23_n_104);
  not mul_8_23_drc_bufs1823(mul_8_23_n_77 ,mul_8_23_n_75);
  not mul_8_23_drc_bufs1824(mul_8_23_n_76 ,mul_8_23_n_75);
  not mul_8_23_drc_bufs1825(mul_8_23_n_75 ,mul_8_23_n_96);
  not mul_8_23_drc_bufs1827(mul_8_23_n_74 ,mul_8_23_n_72);
  not mul_8_23_drc_bufs1828(mul_8_23_n_73 ,mul_8_23_n_72);
  not mul_8_23_drc_bufs1829(mul_8_23_n_72 ,mul_8_23_n_109);
  not mul_8_23_drc_bufs1831(mul_8_23_n_71 ,mul_8_23_n_69);
  not mul_8_23_drc_bufs1832(mul_8_23_n_70 ,mul_8_23_n_69);
  not mul_8_23_drc_bufs1833(mul_8_23_n_69 ,mul_8_23_n_96);
  not mul_8_23_drc_bufs1835(mul_8_23_n_68 ,mul_8_23_n_66);
  not mul_8_23_drc_bufs1836(mul_8_23_n_67 ,mul_8_23_n_66);
  not mul_8_23_drc_bufs1837(mul_8_23_n_66 ,mul_8_23_n_94);
  not mul_8_23_drc_bufs1839(mul_8_23_n_65 ,mul_8_23_n_63);
  not mul_8_23_drc_bufs1840(mul_8_23_n_64 ,mul_8_23_n_63);
  not mul_8_23_drc_bufs1841(mul_8_23_n_63 ,mul_8_23_n_104);
  not mul_8_23_drc_bufs1843(mul_8_23_n_62 ,mul_8_23_n_60);
  not mul_8_23_drc_bufs1844(mul_8_23_n_61 ,mul_8_23_n_60);
  not mul_8_23_drc_bufs1845(mul_8_23_n_60 ,mul_8_23_n_103);
  not mul_8_23_drc_bufs1847(mul_8_23_n_59 ,mul_8_23_n_57);
  not mul_8_23_drc_bufs1848(mul_8_23_n_58 ,mul_8_23_n_57);
  not mul_8_23_drc_bufs1849(mul_8_23_n_57 ,mul_8_23_n_95);
  not mul_8_23_drc_bufs1851(mul_8_23_n_56 ,mul_8_23_n_54);
  not mul_8_23_drc_bufs1852(mul_8_23_n_55 ,mul_8_23_n_54);
  not mul_8_23_drc_bufs1853(mul_8_23_n_54 ,mul_8_23_n_103);
  not mul_8_23_drc_bufs1855(mul_8_23_n_53 ,mul_8_23_n_51);
  not mul_8_23_drc_bufs1856(mul_8_23_n_52 ,mul_8_23_n_51);
  not mul_8_23_drc_bufs1857(mul_8_23_n_51 ,mul_8_23_n_101);
  not mul_8_23_drc_bufs1859(mul_8_23_n_50 ,mul_8_23_n_48);
  not mul_8_23_drc_bufs1860(mul_8_23_n_49 ,mul_8_23_n_48);
  not mul_8_23_drc_bufs1861(mul_8_23_n_48 ,mul_8_23_n_108);
  not mul_8_23_drc_bufs1863(mul_8_23_n_47 ,mul_8_23_n_45);
  not mul_8_23_drc_bufs1864(mul_8_23_n_46 ,mul_8_23_n_45);
  not mul_8_23_drc_bufs1865(mul_8_23_n_45 ,mul_8_23_n_97);
  not mul_8_23_drc_bufs1867(mul_8_23_n_44 ,mul_8_23_n_42);
  not mul_8_23_drc_bufs1868(mul_8_23_n_43 ,mul_8_23_n_42);
  not mul_8_23_drc_bufs1869(mul_8_23_n_42 ,mul_8_23_n_107);
  not mul_8_23_drc_bufs1871(mul_8_23_n_41 ,mul_8_23_n_39);
  not mul_8_23_drc_bufs1872(mul_8_23_n_40 ,mul_8_23_n_39);
  not mul_8_23_drc_bufs1873(mul_8_23_n_39 ,mul_8_23_n_107);
  not mul_8_23_drc_bufs1875(mul_8_23_n_38 ,mul_8_23_n_36);
  not mul_8_23_drc_bufs1876(mul_8_23_n_37 ,mul_8_23_n_36);
  not mul_8_23_drc_bufs1877(mul_8_23_n_36 ,mul_8_23_n_106);
  not mul_8_23_drc_bufs1879(mul_8_23_n_35 ,mul_8_23_n_33);
  not mul_8_23_drc_bufs1880(mul_8_23_n_34 ,mul_8_23_n_33);
  not mul_8_23_drc_bufs1881(mul_8_23_n_33 ,mul_8_23_n_97);
  not mul_8_23_drc_bufs1883(mul_8_23_n_32 ,mul_8_23_n_30);
  not mul_8_23_drc_bufs1884(mul_8_23_n_31 ,mul_8_23_n_30);
  not mul_8_23_drc_bufs1885(mul_8_23_n_30 ,mul_8_23_n_106);
  not mul_8_23_drc_bufs1887(mul_8_23_n_1 ,mul_8_23_n_0);
  not mul_8_23_drc_bufs1888(mul_8_23_n_29 ,mul_8_23_n_0);
  not mul_8_23_drc_bufs1889(mul_8_23_n_0 ,mul_8_23_n_2);
  not mul_8_23_drc_bufs1891(mul_8_23_n_28 ,mul_8_23_n_27);
  not mul_8_23_drc_bufs1893(mul_8_23_n_27 ,mul_8_23_n_101);
  not mul_8_23_drc_bufs1895(mul_8_23_n_26 ,mul_8_23_n_25);
  not mul_8_23_drc_bufs1897(mul_8_23_n_25 ,mul_8_23_n_102);
  not mul_8_23_drc_bufs1899(mul_8_23_n_24 ,mul_8_23_n_23);
  not mul_8_23_drc_bufs1901(mul_8_23_n_23 ,mul_8_23_n_105);
  not mul_8_23_drc_bufs1903(mul_8_23_n_22 ,mul_8_23_n_20);
  not mul_8_23_drc_bufs1904(mul_8_23_n_21 ,mul_8_23_n_20);
  not mul_8_23_drc_bufs1905(mul_8_23_n_20 ,mul_8_23_n_105);
  not mul_8_23_drc_bufs1907(mul_8_23_n_19 ,mul_8_23_n_18);
  not mul_8_23_drc_bufs1909(mul_8_23_n_18 ,mul_8_23_n_94);
  not mul_8_23_drc_bufs1911(mul_8_23_n_17 ,mul_8_23_n_16);
  not mul_8_23_drc_bufs1913(mul_8_23_n_16 ,mul_8_23_n_99);
  not mul_8_23_drc_bufs1915(mul_8_23_n_15 ,mul_8_23_n_14);
  not mul_8_23_drc_bufs1917(mul_8_23_n_14 ,mul_8_23_n_95);
  not mul_8_23_drc_bufs1919(mul_8_23_n_13 ,mul_8_23_n_11);
  not mul_8_23_drc_bufs1920(mul_8_23_n_12 ,mul_8_23_n_11);
  not mul_8_23_drc_bufs1921(mul_8_23_n_11 ,mul_8_23_n_102);
  not mul_8_23_drc_bufs1923(mul_8_23_n_10 ,mul_8_23_n_8);
  not mul_8_23_drc_bufs1924(mul_8_23_n_9 ,mul_8_23_n_8);
  not mul_8_23_drc_bufs1925(mul_8_23_n_8 ,mul_8_23_n_99);
  xnor mul_8_23_g2(mul_8_23_n_7 ,mul_8_23_n_139 ,mul_8_23_n_135);
  xor mul_8_23_g1929(mul_8_23_n_6 ,mul_8_23_n_167 ,mul_8_23_n_134);
  xor mul_8_23_g1930(mul_8_23_n_5 ,mul_8_23_n_171 ,mul_8_23_n_133);
  xor mul_8_23_g1931(mul_8_23_n_4 ,mul_8_23_n_132 ,mul_8_23_n_169);
  xor mul_8_23_g1932(mul_8_23_n_3 ,mul_8_23_n_131 ,mul_8_23_n_176);
  or square_mul_7_21_g599(n_14 ,square_mul_7_21_n_100 ,square_mul_7_21_n_237);
  xnor square_mul_7_21_g600(n_13 ,square_mul_7_21_n_236 ,square_mul_7_21_n_113);
  nor square_mul_7_21_g601(square_mul_7_21_n_237 ,square_mul_7_21_n_102 ,square_mul_7_21_n_236);
  and square_mul_7_21_g602(square_mul_7_21_n_236 ,square_mul_7_21_n_157 ,square_mul_7_21_n_234);
  xnor square_mul_7_21_g603(n_12 ,square_mul_7_21_n_232 ,square_mul_7_21_n_164);
  or square_mul_7_21_g604(square_mul_7_21_n_234 ,square_mul_7_21_n_159 ,square_mul_7_21_n_233);
  not square_mul_7_21_g605(square_mul_7_21_n_233 ,square_mul_7_21_n_232);
  or square_mul_7_21_g606(square_mul_7_21_n_232 ,square_mul_7_21_n_184 ,square_mul_7_21_n_230);
  xnor square_mul_7_21_g607(n_11 ,square_mul_7_21_n_229 ,square_mul_7_21_n_187);
  nor square_mul_7_21_g608(square_mul_7_21_n_230 ,square_mul_7_21_n_185 ,square_mul_7_21_n_229);
  and square_mul_7_21_g609(square_mul_7_21_n_229 ,square_mul_7_21_n_204 ,square_mul_7_21_n_227);
  xnor square_mul_7_21_g610(n_10 ,square_mul_7_21_n_225 ,square_mul_7_21_n_208);
  or square_mul_7_21_g611(square_mul_7_21_n_227 ,square_mul_7_21_n_207 ,square_mul_7_21_n_226);
  not square_mul_7_21_g612(square_mul_7_21_n_226 ,square_mul_7_21_n_225);
  or square_mul_7_21_g613(square_mul_7_21_n_225 ,square_mul_7_21_n_206 ,square_mul_7_21_n_223);
  xnor square_mul_7_21_g614(n_9 ,square_mul_7_21_n_222 ,square_mul_7_21_n_211);
  nor square_mul_7_21_g615(square_mul_7_21_n_223 ,square_mul_7_21_n_203 ,square_mul_7_21_n_222);
  and square_mul_7_21_g616(square_mul_7_21_n_222 ,square_mul_7_21_n_201 ,square_mul_7_21_n_220);
  xnor square_mul_7_21_g617(n_8 ,square_mul_7_21_n_218 ,square_mul_7_21_n_210);
  or square_mul_7_21_g618(square_mul_7_21_n_220 ,square_mul_7_21_n_202 ,square_mul_7_21_n_219);
  not square_mul_7_21_g619(square_mul_7_21_n_219 ,square_mul_7_21_n_218);
  or square_mul_7_21_g620(square_mul_7_21_n_218 ,square_mul_7_21_n_194 ,square_mul_7_21_n_216);
  xnor square_mul_7_21_g621(n_7 ,square_mul_7_21_n_215 ,square_mul_7_21_n_200);
  and square_mul_7_21_g622(square_mul_7_21_n_216 ,square_mul_7_21_n_195 ,square_mul_7_21_n_215);
  or square_mul_7_21_g623(square_mul_7_21_n_215 ,square_mul_7_21_n_190 ,square_mul_7_21_n_213);
  xnor square_mul_7_21_g624(n_6 ,square_mul_7_21_n_212 ,square_mul_7_21_n_3);
  nor square_mul_7_21_g625(square_mul_7_21_n_213 ,square_mul_7_21_n_189 ,square_mul_7_21_n_212);
  and square_mul_7_21_g626(square_mul_7_21_n_212 ,square_mul_7_21_n_172 ,square_mul_7_21_n_205);
  xnor square_mul_7_21_g627(square_mul_7_21_n_211 ,square_mul_7_21_n_197 ,square_mul_7_21_n_192);
  xnor square_mul_7_21_g628(square_mul_7_21_n_210 ,square_mul_7_21_n_191 ,square_mul_7_21_n_182);
  xnor square_mul_7_21_g629(n_5 ,square_mul_7_21_n_198 ,square_mul_7_21_n_176);
  xnor square_mul_7_21_g630(square_mul_7_21_n_208 ,square_mul_7_21_n_196 ,square_mul_7_21_n_168);
  and square_mul_7_21_g631(square_mul_7_21_n_207 ,square_mul_7_21_n_168 ,square_mul_7_21_n_196);
  nor square_mul_7_21_g632(square_mul_7_21_n_206 ,square_mul_7_21_n_197 ,square_mul_7_21_n_193);
  or square_mul_7_21_g633(square_mul_7_21_n_205 ,square_mul_7_21_n_171 ,square_mul_7_21_n_199);
  or square_mul_7_21_g634(square_mul_7_21_n_204 ,square_mul_7_21_n_168 ,square_mul_7_21_n_196);
  and square_mul_7_21_g635(square_mul_7_21_n_203 ,square_mul_7_21_n_197 ,square_mul_7_21_n_193);
  and square_mul_7_21_g636(square_mul_7_21_n_202 ,square_mul_7_21_n_182 ,square_mul_7_21_n_191);
  or square_mul_7_21_g637(square_mul_7_21_n_201 ,square_mul_7_21_n_182 ,square_mul_7_21_n_191);
  xnor square_mul_7_21_g639(square_mul_7_21_n_200 ,square_mul_7_21_n_179 ,square_mul_7_21_n_162);
  not square_mul_7_21_g640(square_mul_7_21_n_199 ,square_mul_7_21_n_198);
  or square_mul_7_21_g641(square_mul_7_21_n_195 ,square_mul_7_21_n_161 ,square_mul_7_21_n_178);
  nor square_mul_7_21_g642(square_mul_7_21_n_194 ,square_mul_7_21_n_162 ,square_mul_7_21_n_179);
  or square_mul_7_21_g643(square_mul_7_21_n_198 ,square_mul_7_21_n_138 ,square_mul_7_21_n_183);
  and square_mul_7_21_g644(square_mul_7_21_n_197 ,square_mul_7_21_n_174 ,square_mul_7_21_n_186);
  and square_mul_7_21_g645(square_mul_7_21_n_196 ,square_mul_7_21_n_167 ,square_mul_7_21_n_181);
  not square_mul_7_21_g646(square_mul_7_21_n_193 ,square_mul_7_21_n_192);
  nor square_mul_7_21_g647(square_mul_7_21_n_190 ,square_mul_7_21_n_160 ,square_mul_7_21_n_180);
  and square_mul_7_21_g648(square_mul_7_21_n_189 ,square_mul_7_21_n_160 ,square_mul_7_21_n_180);
  xnor square_mul_7_21_g649(n_4 ,square_mul_7_21_n_169 ,square_mul_7_21_n_144);
  xnor square_mul_7_21_g650(square_mul_7_21_n_187 ,square_mul_7_21_n_175 ,square_mul_7_21_n_151);
  xnor square_mul_7_21_g651(square_mul_7_21_n_192 ,square_mul_7_21_n_150 ,square_mul_7_21_n_165);
  xnor square_mul_7_21_g652(square_mul_7_21_n_191 ,square_mul_7_21_n_153 ,square_mul_7_21_n_163);
  or square_mul_7_21_g653(square_mul_7_21_n_186 ,square_mul_7_21_n_142 ,square_mul_7_21_n_170);
  and square_mul_7_21_g654(square_mul_7_21_n_185 ,square_mul_7_21_n_175 ,square_mul_7_21_n_152);
  nor square_mul_7_21_g655(square_mul_7_21_n_184 ,square_mul_7_21_n_175 ,square_mul_7_21_n_152);
  and square_mul_7_21_g656(square_mul_7_21_n_183 ,square_mul_7_21_n_132 ,square_mul_7_21_n_169);
  and square_mul_7_21_g657(square_mul_7_21_n_182 ,square_mul_7_21_n_134 ,square_mul_7_21_n_166);
  or square_mul_7_21_g658(square_mul_7_21_n_181 ,square_mul_7_21_n_143 ,square_mul_7_21_n_173);
  xnor square_mul_7_21_g659(square_mul_7_21_n_180 ,square_mul_7_21_n_107 ,square_mul_7_21_n_145);
  not square_mul_7_21_g660(square_mul_7_21_n_178 ,square_mul_7_21_n_179);
  xnor square_mul_7_21_g661(square_mul_7_21_n_179 ,square_mul_7_21_n_154 ,square_mul_7_21_n_146);
  xor square_mul_7_21_g662(n_3 ,square_mul_7_21_n_130 ,square_mul_7_21_n_155);
  xnor square_mul_7_21_g663(square_mul_7_21_n_176 ,square_mul_7_21_n_95 ,square_mul_7_21_n_148);
  or square_mul_7_21_g664(square_mul_7_21_n_174 ,square_mul_7_21_n_104 ,square_mul_7_21_n_153);
  nor square_mul_7_21_g665(square_mul_7_21_n_173 ,square_mul_7_21_n_56 ,square_mul_7_21_n_150);
  or square_mul_7_21_g666(square_mul_7_21_n_172 ,square_mul_7_21_n_94 ,square_mul_7_21_n_147);
  nor square_mul_7_21_g667(square_mul_7_21_n_171 ,square_mul_7_21_n_95 ,square_mul_7_21_n_148);
  and square_mul_7_21_g668(square_mul_7_21_n_170 ,square_mul_7_21_n_104 ,square_mul_7_21_n_153);
  and square_mul_7_21_g669(square_mul_7_21_n_175 ,square_mul_7_21_n_90 ,square_mul_7_21_n_158);
  or square_mul_7_21_g670(square_mul_7_21_n_167 ,square_mul_7_21_n_55 ,square_mul_7_21_n_149);
  or square_mul_7_21_g671(square_mul_7_21_n_166 ,square_mul_7_21_n_131 ,square_mul_7_21_n_154);
  xor square_mul_7_21_g672(square_mul_7_21_n_165 ,square_mul_7_21_n_56 ,square_mul_7_21_n_143);
  xnor square_mul_7_21_g673(square_mul_7_21_n_164 ,square_mul_7_21_n_62 ,square_mul_7_21_n_141);
  xnor square_mul_7_21_g674(square_mul_7_21_n_163 ,square_mul_7_21_n_104 ,square_mul_7_21_n_142);
  or square_mul_7_21_g675(square_mul_7_21_n_169 ,square_mul_7_21_n_133 ,square_mul_7_21_n_156);
  xnor square_mul_7_21_g676(square_mul_7_21_n_168 ,square_mul_7_21_n_137 ,square_mul_7_21_n_110);
  not square_mul_7_21_g677(square_mul_7_21_n_161 ,square_mul_7_21_n_162);
  and square_mul_7_21_g679(square_mul_7_21_n_159 ,square_mul_7_21_n_62 ,square_mul_7_21_n_141);
  or square_mul_7_21_g680(square_mul_7_21_n_158 ,square_mul_7_21_n_89 ,square_mul_7_21_n_137);
  or square_mul_7_21_g681(square_mul_7_21_n_157 ,square_mul_7_21_n_62 ,square_mul_7_21_n_141);
  xnor square_mul_7_21_g683(square_mul_7_21_n_155 ,square_mul_7_21_n_60 ,square_mul_7_21_n_0);
  and square_mul_7_21_g684(square_mul_7_21_n_162 ,square_mul_7_21_n_123 ,square_mul_7_21_n_140);
  and square_mul_7_21_g685(square_mul_7_21_n_160 ,square_mul_7_21_n_93 ,square_mul_7_21_n_139);
  not square_mul_7_21_g686(square_mul_7_21_n_152 ,square_mul_7_21_n_151);
  not square_mul_7_21_g687(square_mul_7_21_n_149 ,square_mul_7_21_n_150);
  not square_mul_7_21_g688(square_mul_7_21_n_147 ,square_mul_7_21_n_148);
  xnor square_mul_7_21_g689(square_mul_7_21_n_146 ,square_mul_7_21_n_97 ,square_mul_7_21_n_117);
  xnor square_mul_7_21_g690(square_mul_7_21_n_145 ,square_mul_7_21_n_57 ,square_mul_7_21_n_1);
  xnor square_mul_7_21_g691(square_mul_7_21_n_144 ,square_mul_7_21_n_106 ,square_mul_7_21_n_2);
  xnor square_mul_7_21_g692(square_mul_7_21_n_154 ,square_mul_7_21_n_71 ,square_mul_7_21_n_112);
  xnor square_mul_7_21_g693(square_mul_7_21_n_153 ,square_mul_7_21_n_76 ,square_mul_7_21_n_111);
  xnor square_mul_7_21_g694(square_mul_7_21_n_151 ,square_mul_7_21_n_79 ,square_mul_7_21_n_121);
  xnor square_mul_7_21_g695(square_mul_7_21_n_150 ,square_mul_7_21_n_75 ,square_mul_7_21_n_122);
  xnor square_mul_7_21_g696(square_mul_7_21_n_148 ,square_mul_7_21_n_119 ,square_mul_7_21_n_114);
  or square_mul_7_21_g697(square_mul_7_21_n_140 ,square_mul_7_21_n_126 ,square_mul_7_21_n_1);
  or square_mul_7_21_g698(square_mul_7_21_n_139 ,square_mul_7_21_n_92 ,square_mul_7_21_n_120);
  nor square_mul_7_21_g699(square_mul_7_21_n_138 ,square_mul_7_21_n_106 ,square_mul_7_21_n_2);
  and square_mul_7_21_g700(square_mul_7_21_n_143 ,square_mul_7_21_n_85 ,square_mul_7_21_n_128);
  and square_mul_7_21_g701(square_mul_7_21_n_142 ,square_mul_7_21_n_86 ,square_mul_7_21_n_125);
  and square_mul_7_21_g702(square_mul_7_21_n_141 ,square_mul_7_21_n_88 ,square_mul_7_21_n_129);
  xor square_mul_7_21_g703(n_2 ,square_mul_7_21_n_109 ,square_mul_7_21_n_83);
  or square_mul_7_21_g705(square_mul_7_21_n_134 ,square_mul_7_21_n_96 ,square_mul_7_21_n_116);
  nor square_mul_7_21_g706(square_mul_7_21_n_133 ,square_mul_7_21_n_60 ,square_mul_7_21_n_115);
  or square_mul_7_21_g707(square_mul_7_21_n_132 ,square_mul_7_21_n_105 ,square_mul_7_21_n_118);
  nor square_mul_7_21_g708(square_mul_7_21_n_131 ,square_mul_7_21_n_97 ,square_mul_7_21_n_117);
  and square_mul_7_21_g709(square_mul_7_21_n_137 ,square_mul_7_21_n_101 ,square_mul_7_21_n_127);
  or square_mul_7_21_g710(square_mul_7_21_n_129 ,square_mul_7_21_n_79 ,square_mul_7_21_n_99);
  or square_mul_7_21_g711(square_mul_7_21_n_128 ,square_mul_7_21_n_76 ,square_mul_7_21_n_91);
  or square_mul_7_21_g712(square_mul_7_21_n_127 ,square_mul_7_21_n_75 ,square_mul_7_21_n_98);
  and square_mul_7_21_g713(square_mul_7_21_n_126 ,square_mul_7_21_n_57 ,square_mul_7_21_n_107);
  or square_mul_7_21_g714(square_mul_7_21_n_125 ,square_mul_7_21_n_63 ,square_mul_7_21_n_87);
  and square_mul_7_21_g715(n_1 ,square_mul_7_21_n_103 ,square_mul_7_21_n_109);
  or square_mul_7_21_g716(square_mul_7_21_n_123 ,square_mul_7_21_n_57 ,square_mul_7_21_n_107);
  xnor square_mul_7_21_g717(square_mul_7_21_n_122 ,square_mul_7_21_n_58 ,in1[5]);
  xnor square_mul_7_21_g718(square_mul_7_21_n_121 ,square_mul_7_21_n_52 ,in1[6]);
  and square_mul_7_21_g719(square_mul_7_21_n_130 ,square_mul_7_21_n_84 ,square_mul_7_21_n_108);
  not square_mul_7_21_g720(square_mul_7_21_n_120 ,square_mul_7_21_n_119);
  not square_mul_7_21_g721(square_mul_7_21_n_118 ,square_mul_7_21_n_2);
  not square_mul_7_21_g722(square_mul_7_21_n_116 ,square_mul_7_21_n_117);
  not square_mul_7_21_g723(square_mul_7_21_n_115 ,square_mul_7_21_n_0);
  xnor square_mul_7_21_g724(square_mul_7_21_n_114 ,square_mul_7_21_n_53 ,square_mul_7_21_n_68);
  xnor square_mul_7_21_g725(square_mul_7_21_n_113 ,square_mul_7_21_n_61 ,in1[7]);
  xnor square_mul_7_21_g726(square_mul_7_21_n_112 ,square_mul_7_21_n_70 ,square_mul_7_21_n_63);
  xnor square_mul_7_21_g727(square_mul_7_21_n_111 ,square_mul_7_21_n_73 ,square_mul_7_21_n_54);
  xnor square_mul_7_21_g728(square_mul_7_21_n_110 ,square_mul_7_21_n_69 ,square_mul_7_21_n_72);
  xnor square_mul_7_21_g730(square_mul_7_21_n_119 ,square_mul_7_21_n_64 ,in1[3]);
  xnor square_mul_7_21_g732(square_mul_7_21_n_117 ,square_mul_7_21_n_65 ,in1[4]);
  not square_mul_7_21_g734(square_mul_7_21_n_108 ,square_mul_7_21_n_109);
  not square_mul_7_21_g735(square_mul_7_21_n_106 ,square_mul_7_21_n_105);
  or square_mul_7_21_g736(square_mul_7_21_n_103 ,in1[1] ,square_mul_7_21_n_82);
  and square_mul_7_21_g744(square_mul_7_21_n_105 ,in1[2] ,square_mul_7_21_n_67);
  not square_mul_7_21_g746(square_mul_7_21_n_96 ,square_mul_7_21_n_97);
  not square_mul_7_21_g747(square_mul_7_21_n_94 ,square_mul_7_21_n_95);
  or square_mul_7_21_g748(square_mul_7_21_n_93 ,square_mul_7_21_n_53 ,square_mul_7_21_n_68);
  and square_mul_7_21_g749(square_mul_7_21_n_92 ,square_mul_7_21_n_53 ,square_mul_7_21_n_68);
  and square_mul_7_21_g750(square_mul_7_21_n_91 ,square_mul_7_21_n_73 ,square_mul_7_21_n_54);
  or square_mul_7_21_g751(square_mul_7_21_n_90 ,square_mul_7_21_n_69 ,square_mul_7_21_n_72);
  and square_mul_7_21_g752(square_mul_7_21_n_89 ,square_mul_7_21_n_69 ,square_mul_7_21_n_72);
  or square_mul_7_21_g753(square_mul_7_21_n_88 ,square_mul_7_21_n_27 ,square_mul_7_21_n_52);
  and square_mul_7_21_g754(square_mul_7_21_n_87 ,square_mul_7_21_n_71 ,square_mul_7_21_n_70);
  or square_mul_7_21_g755(square_mul_7_21_n_86 ,square_mul_7_21_n_71 ,square_mul_7_21_n_70);
  or square_mul_7_21_g756(square_mul_7_21_n_85 ,square_mul_7_21_n_73 ,square_mul_7_21_n_54);
  and square_mul_7_21_g757(square_mul_7_21_n_97 ,square_mul_7_21_n_78 ,square_mul_7_21_n_74);
  and square_mul_7_21_g758(square_mul_7_21_n_95 ,square_mul_7_21_n_80 ,square_mul_7_21_n_66);
  not square_mul_7_21_g759(square_mul_7_21_n_84 ,square_mul_7_21_n_83);
  not square_mul_7_21_g760(square_mul_7_21_n_82 ,square_mul_7_21_n_81);
  not square_mul_7_21_g762(square_mul_7_21_n_78 ,square_mul_7_21_n_77);
  or square_mul_7_21_g764(square_mul_7_21_n_83 ,square_mul_7_21_n_22 ,square_mul_7_21_n_50);
  or square_mul_7_21_g765(square_mul_7_21_n_81 ,square_mul_7_21_n_14 ,square_mul_7_21_n_9);
  and square_mul_7_21_g766(square_mul_7_21_n_80 ,in1[3] ,in1[1]);
  or square_mul_7_21_g767(square_mul_7_21_n_79 ,square_mul_7_21_n_5 ,square_mul_7_21_n_25);
  or square_mul_7_21_g768(square_mul_7_21_n_77 ,square_mul_7_21_n_25 ,square_mul_7_21_n_20);
  or square_mul_7_21_g769(square_mul_7_21_n_76 ,square_mul_7_21_n_6 ,square_mul_7_21_n_14);
  or square_mul_7_21_g770(square_mul_7_21_n_75 ,square_mul_7_21_n_39 ,square_mul_7_21_n_19);
  and square_mul_7_21_g771(square_mul_7_21_n_74 ,in1[5] ,in1[1]);
  or square_mul_7_21_g772(square_mul_7_21_n_73 ,square_mul_7_21_n_37 ,square_mul_7_21_n_17);
  or square_mul_7_21_g773(square_mul_7_21_n_72 ,square_mul_7_21_n_42 ,square_mul_7_21_n_17);
  or square_mul_7_21_g774(square_mul_7_21_n_71 ,square_mul_7_21_n_31 ,square_mul_7_21_n_49);
  or square_mul_7_21_g775(square_mul_7_21_n_70 ,square_mul_7_21_n_28 ,square_mul_7_21_n_46);
  or square_mul_7_21_g776(square_mul_7_21_n_69 ,square_mul_7_21_n_34 ,square_mul_7_21_n_51);
  or square_mul_7_21_g777(square_mul_7_21_n_68 ,square_mul_7_21_n_36 ,square_mul_7_21_n_9);
  not square_mul_7_21_g780(square_mul_7_21_n_60 ,square_mul_7_21_n_59);
  not square_mul_7_21_g781(square_mul_7_21_n_55 ,square_mul_7_21_n_56);
  and square_mul_7_21_g782(square_mul_7_21_n_67 ,in1[3] ,in1[0]);
  and square_mul_7_21_g783(square_mul_7_21_n_66 ,in1[4] ,in1[0]);
  or square_mul_7_21_g784(square_mul_7_21_n_65 ,square_mul_7_21_n_24 ,square_mul_7_21_n_45);
  or square_mul_7_21_g785(square_mul_7_21_n_64 ,square_mul_7_21_n_16 ,square_mul_7_21_n_20);
  or square_mul_7_21_g786(square_mul_7_21_n_63 ,square_mul_7_21_n_39 ,square_mul_7_21_n_50);
  or square_mul_7_21_g787(square_mul_7_21_n_62 ,square_mul_7_21_n_6 ,square_mul_7_21_n_30);
  or square_mul_7_21_g788(square_mul_7_21_n_61 ,square_mul_7_21_n_40 ,square_mul_7_21_n_27);
  and square_mul_7_21_g789(square_mul_7_21_n_59 ,in1[2] ,in1[1]);
  or square_mul_7_21_g790(square_mul_7_21_n_58 ,square_mul_7_21_n_37 ,square_mul_7_21_n_11);
  or square_mul_7_21_g791(square_mul_7_21_n_57 ,square_mul_7_21_n_33 ,square_mul_7_21_n_8);
  and square_mul_7_21_g792(square_mul_7_21_n_56 ,in1[6] ,in1[3]);
  or square_mul_7_21_g793(square_mul_7_21_n_54 ,square_mul_7_21_n_28 ,square_mul_7_21_n_22);
  or square_mul_7_21_g794(square_mul_7_21_n_53 ,square_mul_7_21_n_24 ,square_mul_7_21_n_13);
  or square_mul_7_21_g795(square_mul_7_21_n_52 ,square_mul_7_21_n_34 ,square_mul_7_21_n_31);
  not square_mul_7_21_g796(square_mul_7_21_n_51 ,in1[4]);
  not square_mul_7_21_g797(square_mul_7_21_n_50 ,in1[0]);
  not square_mul_7_21_g798(square_mul_7_21_n_49 ,in1[2]);
  not square_mul_7_21_g799(square_mul_7_21_n_48 ,in1[5]);
  not square_mul_7_21_g800(square_mul_7_21_n_47 ,in1[7]);
  not square_mul_7_21_g801(square_mul_7_21_n_46 ,in1[1]);
  not square_mul_7_21_g802(square_mul_7_21_n_45 ,in1[3]);
  not square_mul_7_21_g803(square_mul_7_21_n_44 ,in1[6]);
  not square_mul_7_21_drc_bufs839(square_mul_7_21_n_42 ,square_mul_7_21_n_41);
  not square_mul_7_21_drc_bufs840(square_mul_7_21_n_41 ,square_mul_7_21_n_47);
  not square_mul_7_21_drc_bufs842(square_mul_7_21_n_40 ,square_mul_7_21_n_38);
  not square_mul_7_21_drc_bufs843(square_mul_7_21_n_39 ,square_mul_7_21_n_38);
  not square_mul_7_21_drc_bufs844(square_mul_7_21_n_38 ,square_mul_7_21_n_47);
  not square_mul_7_21_drc_bufs846(square_mul_7_21_n_37 ,square_mul_7_21_n_35);
  not square_mul_7_21_drc_bufs847(square_mul_7_21_n_36 ,square_mul_7_21_n_35);
  not square_mul_7_21_drc_bufs848(square_mul_7_21_n_35 ,square_mul_7_21_n_48);
  not square_mul_7_21_drc_bufs850(square_mul_7_21_n_34 ,square_mul_7_21_n_32);
  not square_mul_7_21_drc_bufs851(square_mul_7_21_n_33 ,square_mul_7_21_n_32);
  not square_mul_7_21_drc_bufs852(square_mul_7_21_n_32 ,square_mul_7_21_n_44);
  not square_mul_7_21_drc_bufs854(square_mul_7_21_n_31 ,square_mul_7_21_n_29);
  not square_mul_7_21_drc_bufs855(square_mul_7_21_n_30 ,square_mul_7_21_n_29);
  not square_mul_7_21_drc_bufs856(square_mul_7_21_n_29 ,square_mul_7_21_n_48);
  not square_mul_7_21_drc_bufs858(square_mul_7_21_n_28 ,square_mul_7_21_n_26);
  not square_mul_7_21_drc_bufs859(square_mul_7_21_n_27 ,square_mul_7_21_n_26);
  not square_mul_7_21_drc_bufs860(square_mul_7_21_n_26 ,square_mul_7_21_n_44);
  not square_mul_7_21_drc_bufs862(square_mul_7_21_n_25 ,square_mul_7_21_n_23);
  not square_mul_7_21_drc_bufs863(square_mul_7_21_n_24 ,square_mul_7_21_n_23);
  not square_mul_7_21_drc_bufs864(square_mul_7_21_n_23 ,square_mul_7_21_n_51);
  not square_mul_7_21_drc_bufs866(square_mul_7_21_n_22 ,square_mul_7_21_n_21);
  not square_mul_7_21_drc_bufs868(square_mul_7_21_n_21 ,square_mul_7_21_n_49);
  not square_mul_7_21_drc_bufs870(square_mul_7_21_n_20 ,square_mul_7_21_n_18);
  not square_mul_7_21_drc_bufs871(square_mul_7_21_n_19 ,square_mul_7_21_n_18);
  not square_mul_7_21_drc_bufs872(square_mul_7_21_n_18 ,square_mul_7_21_n_49);
  not square_mul_7_21_drc_bufs874(square_mul_7_21_n_17 ,square_mul_7_21_n_15);
  not square_mul_7_21_drc_bufs875(square_mul_7_21_n_16 ,square_mul_7_21_n_15);
  not square_mul_7_21_drc_bufs876(square_mul_7_21_n_15 ,square_mul_7_21_n_45);
  not square_mul_7_21_drc_bufs878(square_mul_7_21_n_14 ,square_mul_7_21_n_12);
  not square_mul_7_21_drc_bufs879(square_mul_7_21_n_13 ,square_mul_7_21_n_12);
  not square_mul_7_21_drc_bufs880(square_mul_7_21_n_12 ,square_mul_7_21_n_46);
  not square_mul_7_21_drc_bufs882(square_mul_7_21_n_11 ,square_mul_7_21_n_10);
  not square_mul_7_21_drc_bufs884(square_mul_7_21_n_10 ,square_mul_7_21_n_51);
  not square_mul_7_21_drc_bufs886(square_mul_7_21_n_9 ,square_mul_7_21_n_7);
  not square_mul_7_21_drc_bufs887(square_mul_7_21_n_8 ,square_mul_7_21_n_7);
  not square_mul_7_21_drc_bufs888(square_mul_7_21_n_7 ,square_mul_7_21_n_50);
  not square_mul_7_21_drc_bufs890(square_mul_7_21_n_6 ,square_mul_7_21_n_4);
  not square_mul_7_21_drc_bufs891(square_mul_7_21_n_5 ,square_mul_7_21_n_4);
  not square_mul_7_21_drc_bufs892(square_mul_7_21_n_4 ,square_mul_7_21_n_47);
  xor square_mul_7_21_g2(square_mul_7_21_n_3 ,square_mul_7_21_n_160 ,square_mul_7_21_n_180);
  xnor square_mul_7_21_g894(square_mul_7_21_n_2 ,square_mul_7_21_n_80 ,square_mul_7_21_n_66);
  xor square_mul_7_21_g895(square_mul_7_21_n_1 ,square_mul_7_21_n_77 ,square_mul_7_21_n_74);
  xor square_mul_7_21_g896(square_mul_7_21_n_0 ,square_mul_7_21_n_67 ,in1[2]);
  not g4044(mul_7_27_n_341 ,in1[1]);
  buf g4045(mul_7_27_n_348 ,in1[1]);
  not g4046(square_mul_7_21_n_102 ,square_mul_7_21_n_41);
  not g4047(square_mul_7_21_n_99 ,square_mul_7_21_n_32);
  not g4048(square_mul_7_21_n_98 ,square_mul_7_21_n_35);
  not g4049(mul_8_23_n_306 ,mul_8_23_n_222);
  not g4050(square_mul_7_21_n_100 ,square_mul_7_21_n_61);
  buf g4051(square_mul_7_21_n_101 ,square_mul_7_21_n_58);
  buf g4052(square_mul_7_21_n_104 ,square_mul_7_21_n_65);
  buf g4053(square_mul_7_21_n_107 ,square_mul_7_21_n_64);
  buf g4054(square_mul_7_21_n_109 ,square_mul_7_21_n_81);
  buf g4055(mul_7_27_n_466 ,mul_7_27_n_59);
  buf g4056(square_mul_7_21_n_156 ,square_mul_7_21_n_130);
  not g4057(mul_7_27_n_351 ,mul_7_27_n_277);
  not g4058(mul_7_27_n_395 ,mul_7_27_n_361);
endmodule
