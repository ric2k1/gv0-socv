module top( 2_n2 , 2_n4 , 2_n6 , 2_n9 , 2_n12 , 2_n18 , 2_n22 , 2_n34 , 2_n35 , 2_n42 , 2_n48 , 2_n51 , 2_n56 , 2_n57 , 2_n65 , 2_n67 , 2_n68 , 2_n72 , 2_n75 , 2_n77 , 2_n78 , 2_n80 );
    input 2_n2 , 2_n4 , 2_n12 , 2_n18 , 2_n22 , 2_n34 , 2_n35 , 2_n51 , 2_n57 , 2_n67 , 2_n72 , 2_n75 , 2_n78 , 2_n80 ;
    output 2_n6 , 2_n9 , 2_n42 , 2_n48 , 2_n56 , 2_n65 , 2_n68 , 2_n77 ;
    wire 2_n0 , 2_n1 , 2_n3 , 2_n5 , 2_n7 , 2_n8 , 2_n10 , 2_n11 , 2_n13 , 2_n14 , 2_n15 , 2_n16 , 2_n17 , 2_n19 , 2_n20 , 2_n21 , 2_n23 , 2_n24 , 2_n25 , 2_n26 , 2_n27 , 2_n28 , 2_n29 , 2_n30 , 2_n31 , 2_n32 , 2_n33 , 2_n36 , 2_n37 , 2_n38 , 2_n39 , 2_n40 , 2_n41 , 2_n43 , 2_n44 , 2_n45 , 2_n46 , 2_n47 , 2_n49 , 2_n50 , 2_n52 , 2_n53 , 2_n54 , 2_n55 , 2_n58 , 2_n59 , 2_n60 , 2_n61 , 2_n62 , 2_n63 , 2_n64 , 2_n66 , 2_n69 , 2_n70 , 2_n71 , 2_n73 , 2_n74 , 2_n76 , 2_n79 , 2_n81 , 2_n82 , 2_n83 , 2_n84 , 2_n85 , 2_n86 , 2_n87 , 2_n88 , 2_n89 , 2_n90 ;
assign 2_n77 = 2_n86 | 2_n73;
assign 2_n5 = ~(2_n45 ^ 2_n53);
assign 2_n9 = 2_n61 ^ 2_n30;
assign 2_n40 = ~(2_n12 | 2_n27);
assign 2_n16 = ~2_n10;
assign 2_n81 = ~2_n84;
assign 2_n31 = 2_n34 & 2_n44;
assign 2_n26 = 2_n80 | 2_n2;
assign 2_n58 = 2_n72 & 2_n67;
assign 2_n24 = ~2_n2;
assign 2_n14 = 2_n21 | 2_n78;
assign 2_n79 = 2_n39 & 2_n1;
assign 2_n20 = 2_n80 | 2_n67;
assign 2_n7 = ~(2_n84 | 2_n76);
assign 2_n52 = 2_n72 & 2_n57;
assign 2_n50 = 2_n28 & 2_n36;
assign 2_n15 = ~2_n45;
assign 2_n69 = ~(2_n0 ^ 2_n50);
assign 2_n3 = ~(2_n72 & 2_n4);
assign 2_n43 = 2_n22 & 2_n20;
assign 2_n27 = 2_n53 & 2_n16;
assign 2_n21 = ~2_n4;
assign 2_n60 = 2_n37 | 2_n12;
assign 2_n1 = 2_n55 & 2_n70;
assign 2_n88 = ~2_n67;
assign 2_n87 = 2_n18 & 2_n26;
assign 2_n48 = ~2_n63;
assign 2_n71 = ~2_n57;
assign 2_n6 = ~(2_n60 ^ 2_n5);
assign 2_n33 = ~(2_n37 | 2_n77);
assign 2_n59 = 2_n35 & 2_n25;
assign 2_n45 = 2_n54 & 2_n43;
assign 2_n55 = 2_n52 | 2_n64;
assign 2_n29 = ~2_n75;
assign 2_n74 = ~(2_n29 | 2_n4);
assign 2_n86 = 2_n90 | 2_n11;
assign 2_n73 = 2_n66 | 2_n45;
assign 2_n42 = 2_n40 ^ 2_n69;
assign 2_n65 = 2_n19 ^ 2_n82;
assign 2_n89 = 2_n9 & 2_n65;
assign 2_n37 = ~2_n51;
assign 2_n90 = 2_n14 & 2_n59;
assign 2_n25 = 2_n80 | 2_n4;
assign 2_n49 = 2_n3 & 2_n38;
assign 2_n10 = 2_n51 & 2_n15;
assign 2_n61 = ~(2_n12 | 2_n7);
assign 2_n68 = 2_n33 | 2_n63;
assign 2_n70 = 2_n11 | 2_n47;
assign 2_n36 = ~(2_n18 | 2_n23);
assign 2_n46 = 2_n71 | 2_n78;
assign 2_n32 = ~(2_n90 | 2_n1);
assign 2_n39 = 2_n11 | 2_n81;
assign 2_n13 = ~(2_n29 | 2_n57);
assign 2_n82 = 2_n90 ^ 2_n49;
assign 2_n56 = 2_n8 & 2_n89;
assign 2_n30 = ~(2_n11 ^ 2_n55);
assign 2_n41 = 2_n22 | 2_n83;
assign 2_n54 = 2_n88 | 2_n78;
assign 2_n17 = ~2_n72;
assign 2_n19 = ~(2_n12 | 2_n79);
assign 2_n38 = ~(2_n35 | 2_n74);
assign 2_n11 = 2_n46 & 2_n31;
assign 2_n23 = ~(2_n29 | 2_n2);
assign 2_n44 = 2_n80 | 2_n57;
assign 2_n76 = 2_n50 | 2_n62;
assign 2_n66 = 2_n85 & 2_n87;
assign 2_n53 = 2_n58 | 2_n41;
assign 2_n85 = 2_n24 | 2_n78;
assign 2_n83 = ~(2_n29 | 2_n67);
assign 2_n0 = ~2_n66;
assign 2_n47 = ~2_n76;
assign 2_n63 = 2_n49 | 2_n32;
assign 2_n62 = ~(2_n53 | 2_n66);
assign 2_n8 = 2_n6 & 2_n42;
assign 2_n84 = 2_n0 & 2_n10;
assign 2_n64 = 2_n34 | 2_n13;
assign 2_n28 = 2_n17 | 2_n24;
endmodule
