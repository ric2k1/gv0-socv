module top( 1_n9 , 1_n22 , 1_n103 , 1_n124 , 1_n134 , 1_n201 , 1_n211 , 1_n287 , 1_n353 , 1_n358 , 1_n370 , 1_n389 , 1_n396 , 1_n401 , 1_n411 , 1_n443 , 1_n460 , 1_n469 , 1_n497 , 1_n499 , 1_n510 , 1_n537 , 1_n573 , 1_n603 , 1_n728 , 1_n758 , 1_n761 , 1_n762 , 1_n767 , 1_n772 , 1_n777 , 1_n800 , 1_n817 , 1_n831 , 1_n834 , 1_n846 , 1_n854 , 1_n922 , 1_n927 , 1_n937 , 1_n951 , 1_n985 , 1_n1007 , 1_n1084 , 1_n1097 , 1_n1112 , 1_n1165 , 1_n1181 , 1_n1198 , 1_n1231 , 1_n1302 , 1_n1307 , 1_n1364 , 1_n1392 , 1_n1401 , 1_n1487 , 1_n1561 , 1_n1636 , 1_n1650 , 1_n1709 , 1_n1724 , 1_n1757 , 1_n1806 , 1_n1860 , 1_n1912 , 1_n1916 , 1_n1937 , 1_n1982 , 1_n2057 , 1_n2061 , 1_n2068 , 1_n2174 , 1_n2190 , 1_n2235 , 1_n2252 , 1_n2295 , 1_n2339 , 1_n2341 , 1_n2458 , 1_n2482 , 1_n2498 , 1_n2549 , 1_n2590 , 1_n2592 , 1_n2666 , 1_n2709 , 1_n2737 , 1_n2758 , 1_n2771 , 1_n2777 , 1_n2805 , 1_n2882 , 1_n2904 , 1_n2934 , 1_n3006 , 1_n3076 , 1_n3085 , 1_n3112 , 1_n3130 , 1_n3178 , 1_n3262 , 1_n3311 , 1_n3323 , 1_n3362 , 1_n3409 , 1_n3591 , 1_n3641 , 1_n3669 , 1_n3677 , 1_n3748 , 1_n3769 , 1_n3790 , 1_n3815 , 1_n3832 , 1_n3946 , 1_n4006 , 1_n4059 , 1_n4075 , 1_n4114 , 1_n4122 , 1_n4141 , 1_n4202 , 1_n4330 , 1_n4335 , 1_n4357 , 1_n4382 , 1_n4419 , 1_n4452 , 1_n4470 , 1_n4553 , 1_n4743 , 1_n4748 , 1_n4777 , 1_n4824 , 1_n4862 , 1_n4864 , 1_n4964 , 1_n4998 , 1_n5003 , 1_n5031 , 1_n5060 , 1_n5065 , 1_n5167 , 1_n5189 , 1_n5214 , 1_n5320 , 1_n5356 , 1_n5364 , 1_n5427 , 1_n5470 , 1_n5536 , 1_n5548 , 1_n5549 , 1_n5557 , 1_n5568 , 1_n5586 , 1_n5609 , 1_n5671 , 1_n5684 , 1_n5715 , 1_n5729 , 1_n5758 , 1_n5801 , 1_n5882 , 1_n5884 , 1_n5920 , 1_n5962 , 1_n5969 , 1_n6019 , 1_n6023 , 1_n6085 , 1_n6103 , 1_n6109 , 1_n6149 , 1_n6168 , 1_n6297 , 1_n6301 , 1_n6333 , 1_n6392 , 1_n6409 , 1_n6434 , 1_n6586 , 1_n6655 , 1_n6668 , 1_n6683 , 1_n6818 , 1_n6826 , 1_n6843 , 1_n6862 , 1_n6937 , 1_n7034 , 1_n7061 , 1_n7111 , 1_n7113 , 1_n7132 , 1_n7161 , 1_n7241 , 1_n7374 , 1_n7411 , 1_n7529 , 1_n7553 , 1_n7582 , 1_n7659 , 1_n7687 , 1_n7715 , 1_n7720 , 1_n7729 , 1_n7755 , 1_n7772 , 1_n7790 , 1_n7812 , 1_n7858 , 1_n7860 , 1_n7968 , 1_n7974 , 1_n8139 , 1_n8163 , 1_n8172 , 1_n8183 , 1_n8219 , 1_n8228 , 1_n8230 , 1_n8233 , 1_n8265 , 1_n8290 , 1_n8308 , 1_n8332 , 1_n8336 , 1_n8466 , 1_n8468 , 1_n8506 , 1_n8516 , 1_n8522 , 1_n8701 , 1_n8716 , 1_n8768 , 1_n8820 , 1_n8859 , 1_n8860 , 1_n8940 , 1_n9041 , 1_n9093 , 1_n9100 , 1_n9187 , 1_n9216 , 1_n9300 , 1_n9329 , 1_n9353 , 1_n9475 , 1_n9528 , 1_n9531 , 1_n9570 , 1_n9591 , 1_n9620 , 1_n9669 , 1_n9732 , 1_n9747 , 1_n9846 , 1_n9866 , 1_n9872 , 1_n9887 , 1_n9906 , 1_n9915 , 1_n10063 , 1_n10101 , 1_n10113 , 1_n10122 , 1_n10142 , 1_n10162 , 1_n10168 , 1_n10243 , 1_n10408 , 1_n10416 , 1_n10451 , 1_n10453 , 1_n10522 , 1_n10524 , 1_n10560 , 1_n10594 , 1_n10606 , 1_n10628 , 1_n10642 , 1_n10657 , 1_n10736 , 1_n10770 , 1_n10797 , 1_n10805 , 1_n10866 , 1_n10874 , 1_n10908 , 1_n11030 , 1_n11057 , 1_n11058 , 1_n11061 , 1_n11077 , 1_n11109 , 1_n11111 , 1_n11140 , 1_n11147 , 1_n11180 , 1_n11222 , 1_n11236 , 1_n11252 , 1_n11264 , 1_n11324 , 1_n11350 , 1_n11396 , 1_n11411 , 1_n11429 , 1_n11484 , 1_n11488 , 1_n11537 , 1_n11574 , 1_n11634 , 1_n11665 , 1_n11667 , 1_n11732 , 1_n11734 , 1_n11778 , 1_n11792 , 1_n11835 , 1_n11879 , 1_n11882 , 1_n11891 , 1_n11895 , 1_n12003 , 1_n12059 , 1_n12065 , 1_n12067 , 1_n12187 , 1_n12263 , 1_n12284 , 1_n12289 , 1_n12306 , 1_n12334 , 1_n12348 , 1_n12352 , 1_n12372 , 1_n12406 , 1_n12408 , 1_n12463 , 1_n12482 , 1_n12503 , 1_n12515 , 1_n12579 , 1_n12592 , 1_n12605 , 1_n12616 , 1_n12651 , 1_n12693 , 1_n12750 , 1_n12839 , 1_n12853 , 1_n12912 , 1_n12965 , 1_n12968 , 1_n13002 , 1_n13035 , 1_n13058 , 1_n13060 , 1_n13201 );
    input 1_n9 , 1_n22 , 1_n103 , 1_n124 , 1_n287 , 1_n353 , 1_n389 , 1_n401 , 1_n411 , 1_n443 , 1_n469 , 1_n497 , 1_n499 , 1_n510 , 1_n603 , 1_n761 , 1_n767 , 1_n772 , 1_n817 , 1_n834 , 1_n854 , 1_n937 , 1_n951 , 1_n1007 , 1_n1084 , 1_n1165 , 1_n1198 , 1_n1231 , 1_n1302 , 1_n1307 , 1_n1364 , 1_n1392 , 1_n1636 , 1_n1650 , 1_n1709 , 1_n1724 , 1_n1757 , 1_n1912 , 1_n1916 , 1_n1982 , 1_n2057 , 1_n2068 , 1_n2174 , 1_n2252 , 1_n2295 , 1_n2339 , 1_n2341 , 1_n2458 , 1_n2482 , 1_n2498 , 1_n2590 , 1_n2592 , 1_n2666 , 1_n2737 , 1_n2758 , 1_n2771 , 1_n2777 , 1_n2882 , 1_n3006 , 1_n3076 , 1_n3085 , 1_n3112 , 1_n3130 , 1_n3178 , 1_n3311 , 1_n3409 , 1_n3591 , 1_n3641 , 1_n3669 , 1_n3677 , 1_n3769 , 1_n3815 , 1_n3832 , 1_n4006 , 1_n4075 , 1_n4114 , 1_n4122 , 1_n4141 , 1_n4330 , 1_n4335 , 1_n4357 , 1_n4382 , 1_n4419 , 1_n4452 , 1_n4470 , 1_n4743 , 1_n4748 , 1_n4862 , 1_n4964 , 1_n4998 , 1_n5031 , 1_n5065 , 1_n5167 , 1_n5189 , 1_n5214 , 1_n5320 , 1_n5356 , 1_n5427 , 1_n5470 , 1_n5536 , 1_n5548 , 1_n5568 , 1_n5586 , 1_n5671 , 1_n5684 , 1_n5715 , 1_n5729 , 1_n5758 , 1_n5801 , 1_n5884 , 1_n5920 , 1_n5962 , 1_n5969 , 1_n6023 , 1_n6085 , 1_n6149 , 1_n6168 , 1_n6333 , 1_n6392 , 1_n6409 , 1_n6655 , 1_n6668 , 1_n6818 , 1_n6826 , 1_n6843 , 1_n6937 , 1_n7061 , 1_n7113 , 1_n7161 , 1_n7374 , 1_n7411 , 1_n7529 , 1_n7659 , 1_n7715 , 1_n7720 , 1_n7729 , 1_n7772 , 1_n7812 , 1_n7974 , 1_n8139 , 1_n8163 , 1_n8183 , 1_n8228 , 1_n8230 , 1_n8233 , 1_n8290 , 1_n8308 , 1_n8332 , 1_n8466 , 1_n8468 , 1_n8506 , 1_n8522 , 1_n8716 , 1_n8768 , 1_n8820 , 1_n8859 , 1_n8860 , 1_n8940 , 1_n9041 , 1_n9093 , 1_n9187 , 1_n9216 , 1_n9300 , 1_n9353 , 1_n9475 , 1_n9528 , 1_n9531 , 1_n9570 , 1_n9591 , 1_n9620 , 1_n9669 , 1_n9732 , 1_n9747 , 1_n9846 , 1_n9887 , 1_n9906 , 1_n9915 , 1_n10063 , 1_n10113 , 1_n10122 , 1_n10142 , 1_n10162 , 1_n10168 , 1_n10408 , 1_n10416 , 1_n10451 , 1_n10522 , 1_n10560 , 1_n10594 , 1_n10606 , 1_n10642 , 1_n10657 , 1_n10770 , 1_n10805 , 1_n10866 , 1_n10874 , 1_n10908 , 1_n11030 , 1_n11058 , 1_n11061 , 1_n11109 , 1_n11111 , 1_n11180 , 1_n11222 , 1_n11236 , 1_n11324 , 1_n11350 , 1_n11396 , 1_n11411 , 1_n11429 , 1_n11488 , 1_n11537 , 1_n11574 , 1_n11634 , 1_n11665 , 1_n11734 , 1_n11835 , 1_n11891 , 1_n12003 , 1_n12065 , 1_n12263 , 1_n12284 , 1_n12289 , 1_n12306 , 1_n12348 , 1_n12352 , 1_n12372 , 1_n12408 , 1_n12482 , 1_n12579 , 1_n12592 , 1_n12605 , 1_n12651 , 1_n12693 , 1_n12750 , 1_n12853 , 1_n12912 , 1_n12965 , 1_n13058 , 1_n13060 , 1_n13201 ;
    output 1_n134 , 1_n201 , 1_n211 , 1_n358 , 1_n370 , 1_n396 , 1_n460 , 1_n537 , 1_n573 , 1_n728 , 1_n758 , 1_n762 , 1_n777 , 1_n800 , 1_n831 , 1_n846 , 1_n922 , 1_n927 , 1_n985 , 1_n1097 , 1_n1112 , 1_n1181 , 1_n1401 , 1_n1487 , 1_n1561 , 1_n1806 , 1_n1860 , 1_n1937 , 1_n2061 , 1_n2190 , 1_n2235 , 1_n2549 , 1_n2709 , 1_n2805 , 1_n2904 , 1_n2934 , 1_n3262 , 1_n3323 , 1_n3362 , 1_n3748 , 1_n3790 , 1_n3946 , 1_n4059 , 1_n4202 , 1_n4553 , 1_n4777 , 1_n4824 , 1_n4864 , 1_n5003 , 1_n5060 , 1_n5364 , 1_n5549 , 1_n5557 , 1_n5609 , 1_n5882 , 1_n6019 , 1_n6103 , 1_n6109 , 1_n6297 , 1_n6301 , 1_n6434 , 1_n6586 , 1_n6683 , 1_n6862 , 1_n7034 , 1_n7111 , 1_n7132 , 1_n7241 , 1_n7553 , 1_n7582 , 1_n7687 , 1_n7755 , 1_n7790 , 1_n7858 , 1_n7860 , 1_n7968 , 1_n8172 , 1_n8219 , 1_n8265 , 1_n8336 , 1_n8516 , 1_n8701 , 1_n9100 , 1_n9329 , 1_n9866 , 1_n9872 , 1_n10101 , 1_n10243 , 1_n10453 , 1_n10524 , 1_n10628 , 1_n10736 , 1_n10797 , 1_n11057 , 1_n11077 , 1_n11140 , 1_n11147 , 1_n11252 , 1_n11264 , 1_n11484 , 1_n11667 , 1_n11732 , 1_n11778 , 1_n11792 , 1_n11879 , 1_n11882 , 1_n11895 , 1_n12059 , 1_n12067 , 1_n12187 , 1_n12334 , 1_n12406 , 1_n12463 , 1_n12503 , 1_n12515 , 1_n12616 , 1_n12839 , 1_n12968 , 1_n13002 , 1_n13035 ;
    wire 1_n0 , 1_n1 , 1_n2 , 1_n3 , 1_n4 , 1_n5 , 1_n6 , 1_n7 , 1_n8 , 1_n10 , 1_n11 , 1_n12 , 1_n13 , 1_n14 , 1_n15 , 1_n16 , 1_n17 , 1_n18 , 1_n19 , 1_n20 , 1_n21 , 1_n23 , 1_n24 , 1_n25 , 1_n26 , 1_n27 , 1_n28 , 1_n29 , 1_n30 , 1_n31 , 1_n32 , 1_n33 , 1_n34 , 1_n35 , 1_n36 , 1_n37 , 1_n38 , 1_n39 , 1_n40 , 1_n41 , 1_n42 , 1_n43 , 1_n44 , 1_n45 , 1_n46 , 1_n47 , 1_n48 , 1_n49 , 1_n50 , 1_n51 , 1_n52 , 1_n53 , 1_n54 , 1_n55 , 1_n56 , 1_n57 , 1_n58 , 1_n59 , 1_n60 , 1_n61 , 1_n62 , 1_n63 , 1_n64 , 1_n65 , 1_n66 , 1_n67 , 1_n68 , 1_n69 , 1_n70 , 1_n71 , 1_n72 , 1_n73 , 1_n74 , 1_n75 , 1_n76 , 1_n77 , 1_n78 , 1_n79 , 1_n80 , 1_n81 , 1_n82 , 1_n83 , 1_n84 , 1_n85 , 1_n86 , 1_n87 , 1_n88 , 1_n89 , 1_n90 , 1_n91 , 1_n92 , 1_n93 , 1_n94 , 1_n95 , 1_n96 , 1_n97 , 1_n98 , 1_n99 , 1_n100 , 1_n101 , 1_n102 , 1_n104 , 1_n105 , 1_n106 , 1_n107 , 1_n108 , 1_n109 , 1_n110 , 1_n111 , 1_n112 , 1_n113 , 1_n114 , 1_n115 , 1_n116 , 1_n117 , 1_n118 , 1_n119 , 1_n120 , 1_n121 , 1_n122 , 1_n123 , 1_n125 , 1_n126 , 1_n127 , 1_n128 , 1_n129 , 1_n130 , 1_n131 , 1_n132 , 1_n133 , 1_n135 , 1_n136 , 1_n137 , 1_n138 , 1_n139 , 1_n140 , 1_n141 , 1_n142 , 1_n143 , 1_n144 , 1_n145 , 1_n146 , 1_n147 , 1_n148 , 1_n149 , 1_n150 , 1_n151 , 1_n152 , 1_n153 , 1_n154 , 1_n155 , 1_n156 , 1_n157 , 1_n158 , 1_n159 , 1_n160 , 1_n161 , 1_n162 , 1_n163 , 1_n164 , 1_n165 , 1_n166 , 1_n167 , 1_n168 , 1_n169 , 1_n170 , 1_n171 , 1_n172 , 1_n173 , 1_n174 , 1_n175 , 1_n176 , 1_n177 , 1_n178 , 1_n179 , 1_n180 , 1_n181 , 1_n182 , 1_n183 , 1_n184 , 1_n185 , 1_n186 , 1_n187 , 1_n188 , 1_n189 , 1_n190 , 1_n191 , 1_n192 , 1_n193 , 1_n194 , 1_n195 , 1_n196 , 1_n197 , 1_n198 , 1_n199 , 1_n200 , 1_n202 , 1_n203 , 1_n204 , 1_n205 , 1_n206 , 1_n207 , 1_n208 , 1_n209 , 1_n210 , 1_n212 , 1_n213 , 1_n214 , 1_n215 , 1_n216 , 1_n217 , 1_n218 , 1_n219 , 1_n220 , 1_n221 , 1_n222 , 1_n223 , 1_n224 , 1_n225 , 1_n226 , 1_n227 , 1_n228 , 1_n229 , 1_n230 , 1_n231 , 1_n232 , 1_n233 , 1_n234 , 1_n235 , 1_n236 , 1_n237 , 1_n238 , 1_n239 , 1_n240 , 1_n241 , 1_n242 , 1_n243 , 1_n244 , 1_n245 , 1_n246 , 1_n247 , 1_n248 , 1_n249 , 1_n250 , 1_n251 , 1_n252 , 1_n253 , 1_n254 , 1_n255 , 1_n256 , 1_n257 , 1_n258 , 1_n259 , 1_n260 , 1_n261 , 1_n262 , 1_n263 , 1_n264 , 1_n265 , 1_n266 , 1_n267 , 1_n268 , 1_n269 , 1_n270 , 1_n271 , 1_n272 , 1_n273 , 1_n274 , 1_n275 , 1_n276 , 1_n277 , 1_n278 , 1_n279 , 1_n280 , 1_n281 , 1_n282 , 1_n283 , 1_n284 , 1_n285 , 1_n286 , 1_n288 , 1_n289 , 1_n290 , 1_n291 , 1_n292 , 1_n293 , 1_n294 , 1_n295 , 1_n296 , 1_n297 , 1_n298 , 1_n299 , 1_n300 , 1_n301 , 1_n302 , 1_n303 , 1_n304 , 1_n305 , 1_n306 , 1_n307 , 1_n308 , 1_n309 , 1_n310 , 1_n311 , 1_n312 , 1_n313 , 1_n314 , 1_n315 , 1_n316 , 1_n317 , 1_n318 , 1_n319 , 1_n320 , 1_n321 , 1_n322 , 1_n323 , 1_n324 , 1_n325 , 1_n326 , 1_n327 , 1_n328 , 1_n329 , 1_n330 , 1_n331 , 1_n332 , 1_n333 , 1_n334 , 1_n335 , 1_n336 , 1_n337 , 1_n338 , 1_n339 , 1_n340 , 1_n341 , 1_n342 , 1_n343 , 1_n344 , 1_n345 , 1_n346 , 1_n347 , 1_n348 , 1_n349 , 1_n350 , 1_n351 , 1_n352 , 1_n354 , 1_n355 , 1_n356 , 1_n357 , 1_n359 , 1_n360 , 1_n361 , 1_n362 , 1_n363 , 1_n364 , 1_n365 , 1_n366 , 1_n367 , 1_n368 , 1_n369 , 1_n371 , 1_n372 , 1_n373 , 1_n374 , 1_n375 , 1_n376 , 1_n377 , 1_n378 , 1_n379 , 1_n380 , 1_n381 , 1_n382 , 1_n383 , 1_n384 , 1_n385 , 1_n386 , 1_n387 , 1_n388 , 1_n390 , 1_n391 , 1_n392 , 1_n393 , 1_n394 , 1_n395 , 1_n397 , 1_n398 , 1_n399 , 1_n400 , 1_n402 , 1_n403 , 1_n404 , 1_n405 , 1_n406 , 1_n407 , 1_n408 , 1_n409 , 1_n410 , 1_n412 , 1_n413 , 1_n414 , 1_n415 , 1_n416 , 1_n417 , 1_n418 , 1_n419 , 1_n420 , 1_n421 , 1_n422 , 1_n423 , 1_n424 , 1_n425 , 1_n426 , 1_n427 , 1_n428 , 1_n429 , 1_n430 , 1_n431 , 1_n432 , 1_n433 , 1_n434 , 1_n435 , 1_n436 , 1_n437 , 1_n438 , 1_n439 , 1_n440 , 1_n441 , 1_n442 , 1_n444 , 1_n445 , 1_n446 , 1_n447 , 1_n448 , 1_n449 , 1_n450 , 1_n451 , 1_n452 , 1_n453 , 1_n454 , 1_n455 , 1_n456 , 1_n457 , 1_n458 , 1_n459 , 1_n461 , 1_n462 , 1_n463 , 1_n464 , 1_n465 , 1_n466 , 1_n467 , 1_n468 , 1_n470 , 1_n471 , 1_n472 , 1_n473 , 1_n474 , 1_n475 , 1_n476 , 1_n477 , 1_n478 , 1_n479 , 1_n480 , 1_n481 , 1_n482 , 1_n483 , 1_n484 , 1_n485 , 1_n486 , 1_n487 , 1_n488 , 1_n489 , 1_n490 , 1_n491 , 1_n492 , 1_n493 , 1_n494 , 1_n495 , 1_n496 , 1_n498 , 1_n500 , 1_n501 , 1_n502 , 1_n503 , 1_n504 , 1_n505 , 1_n506 , 1_n507 , 1_n508 , 1_n509 , 1_n511 , 1_n512 , 1_n513 , 1_n514 , 1_n515 , 1_n516 , 1_n517 , 1_n518 , 1_n519 , 1_n520 , 1_n521 , 1_n522 , 1_n523 , 1_n524 , 1_n525 , 1_n526 , 1_n527 , 1_n528 , 1_n529 , 1_n530 , 1_n531 , 1_n532 , 1_n533 , 1_n534 , 1_n535 , 1_n536 , 1_n538 , 1_n539 , 1_n540 , 1_n541 , 1_n542 , 1_n543 , 1_n544 , 1_n545 , 1_n546 , 1_n547 , 1_n548 , 1_n549 , 1_n550 , 1_n551 , 1_n552 , 1_n553 , 1_n554 , 1_n555 , 1_n556 , 1_n557 , 1_n558 , 1_n559 , 1_n560 , 1_n561 , 1_n562 , 1_n563 , 1_n564 , 1_n565 , 1_n566 , 1_n567 , 1_n568 , 1_n569 , 1_n570 , 1_n571 , 1_n572 , 1_n574 , 1_n575 , 1_n576 , 1_n577 , 1_n578 , 1_n579 , 1_n580 , 1_n581 , 1_n582 , 1_n583 , 1_n584 , 1_n585 , 1_n586 , 1_n587 , 1_n588 , 1_n589 , 1_n590 , 1_n591 , 1_n592 , 1_n593 , 1_n594 , 1_n595 , 1_n596 , 1_n597 , 1_n598 , 1_n599 , 1_n600 , 1_n601 , 1_n602 , 1_n604 , 1_n605 , 1_n606 , 1_n607 , 1_n608 , 1_n609 , 1_n610 , 1_n611 , 1_n612 , 1_n613 , 1_n614 , 1_n615 , 1_n616 , 1_n617 , 1_n618 , 1_n619 , 1_n620 , 1_n621 , 1_n622 , 1_n623 , 1_n624 , 1_n625 , 1_n626 , 1_n627 , 1_n628 , 1_n629 , 1_n630 , 1_n631 , 1_n632 , 1_n633 , 1_n634 , 1_n635 , 1_n636 , 1_n637 , 1_n638 , 1_n639 , 1_n640 , 1_n641 , 1_n642 , 1_n643 , 1_n644 , 1_n645 , 1_n646 , 1_n647 , 1_n648 , 1_n649 , 1_n650 , 1_n651 , 1_n652 , 1_n653 , 1_n654 , 1_n655 , 1_n656 , 1_n657 , 1_n658 , 1_n659 , 1_n660 , 1_n661 , 1_n662 , 1_n663 , 1_n664 , 1_n665 , 1_n666 , 1_n667 , 1_n668 , 1_n669 , 1_n670 , 1_n671 , 1_n672 , 1_n673 , 1_n674 , 1_n675 , 1_n676 , 1_n677 , 1_n678 , 1_n679 , 1_n680 , 1_n681 , 1_n682 , 1_n683 , 1_n684 , 1_n685 , 1_n686 , 1_n687 , 1_n688 , 1_n689 , 1_n690 , 1_n691 , 1_n692 , 1_n693 , 1_n694 , 1_n695 , 1_n696 , 1_n697 , 1_n698 , 1_n699 , 1_n700 , 1_n701 , 1_n702 , 1_n703 , 1_n704 , 1_n705 , 1_n706 , 1_n707 , 1_n708 , 1_n709 , 1_n710 , 1_n711 , 1_n712 , 1_n713 , 1_n714 , 1_n715 , 1_n716 , 1_n717 , 1_n718 , 1_n719 , 1_n720 , 1_n721 , 1_n722 , 1_n723 , 1_n724 , 1_n725 , 1_n726 , 1_n727 , 1_n729 , 1_n730 , 1_n731 , 1_n732 , 1_n733 , 1_n734 , 1_n735 , 1_n736 , 1_n737 , 1_n738 , 1_n739 , 1_n740 , 1_n741 , 1_n742 , 1_n743 , 1_n744 , 1_n745 , 1_n746 , 1_n747 , 1_n748 , 1_n749 , 1_n750 , 1_n751 , 1_n752 , 1_n753 , 1_n754 , 1_n755 , 1_n756 , 1_n757 , 1_n759 , 1_n760 , 1_n763 , 1_n764 , 1_n765 , 1_n766 , 1_n768 , 1_n769 , 1_n770 , 1_n771 , 1_n773 , 1_n774 , 1_n775 , 1_n776 , 1_n778 , 1_n779 , 1_n780 , 1_n781 , 1_n782 , 1_n783 , 1_n784 , 1_n785 , 1_n786 , 1_n787 , 1_n788 , 1_n789 , 1_n790 , 1_n791 , 1_n792 , 1_n793 , 1_n794 , 1_n795 , 1_n796 , 1_n797 , 1_n798 , 1_n799 , 1_n801 , 1_n802 , 1_n803 , 1_n804 , 1_n805 , 1_n806 , 1_n807 , 1_n808 , 1_n809 , 1_n810 , 1_n811 , 1_n812 , 1_n813 , 1_n814 , 1_n815 , 1_n816 , 1_n818 , 1_n819 , 1_n820 , 1_n821 , 1_n822 , 1_n823 , 1_n824 , 1_n825 , 1_n826 , 1_n827 , 1_n828 , 1_n829 , 1_n830 , 1_n832 , 1_n833 , 1_n835 , 1_n836 , 1_n837 , 1_n838 , 1_n839 , 1_n840 , 1_n841 , 1_n842 , 1_n843 , 1_n844 , 1_n845 , 1_n847 , 1_n848 , 1_n849 , 1_n850 , 1_n851 , 1_n852 , 1_n853 , 1_n855 , 1_n856 , 1_n857 , 1_n858 , 1_n859 , 1_n860 , 1_n861 , 1_n862 , 1_n863 , 1_n864 , 1_n865 , 1_n866 , 1_n867 , 1_n868 , 1_n869 , 1_n870 , 1_n871 , 1_n872 , 1_n873 , 1_n874 , 1_n875 , 1_n876 , 1_n877 , 1_n878 , 1_n879 , 1_n880 , 1_n881 , 1_n882 , 1_n883 , 1_n884 , 1_n885 , 1_n886 , 1_n887 , 1_n888 , 1_n889 , 1_n890 , 1_n891 , 1_n892 , 1_n893 , 1_n894 , 1_n895 , 1_n896 , 1_n897 , 1_n898 , 1_n899 , 1_n900 , 1_n901 , 1_n902 , 1_n903 , 1_n904 , 1_n905 , 1_n906 , 1_n907 , 1_n908 , 1_n909 , 1_n910 , 1_n911 , 1_n912 , 1_n913 , 1_n914 , 1_n915 , 1_n916 , 1_n917 , 1_n918 , 1_n919 , 1_n920 , 1_n921 , 1_n923 , 1_n924 , 1_n925 , 1_n926 , 1_n928 , 1_n929 , 1_n930 , 1_n931 , 1_n932 , 1_n933 , 1_n934 , 1_n935 , 1_n936 , 1_n938 , 1_n939 , 1_n940 , 1_n941 , 1_n942 , 1_n943 , 1_n944 , 1_n945 , 1_n946 , 1_n947 , 1_n948 , 1_n949 , 1_n950 , 1_n952 , 1_n953 , 1_n954 , 1_n955 , 1_n956 , 1_n957 , 1_n958 , 1_n959 , 1_n960 , 1_n961 , 1_n962 , 1_n963 , 1_n964 , 1_n965 , 1_n966 , 1_n967 , 1_n968 , 1_n969 , 1_n970 , 1_n971 , 1_n972 , 1_n973 , 1_n974 , 1_n975 , 1_n976 , 1_n977 , 1_n978 , 1_n979 , 1_n980 , 1_n981 , 1_n982 , 1_n983 , 1_n984 , 1_n986 , 1_n987 , 1_n988 , 1_n989 , 1_n990 , 1_n991 , 1_n992 , 1_n993 , 1_n994 , 1_n995 , 1_n996 , 1_n997 , 1_n998 , 1_n999 , 1_n1000 , 1_n1001 , 1_n1002 , 1_n1003 , 1_n1004 , 1_n1005 , 1_n1006 , 1_n1008 , 1_n1009 , 1_n1010 , 1_n1011 , 1_n1012 , 1_n1013 , 1_n1014 , 1_n1015 , 1_n1016 , 1_n1017 , 1_n1018 , 1_n1019 , 1_n1020 , 1_n1021 , 1_n1022 , 1_n1023 , 1_n1024 , 1_n1025 , 1_n1026 , 1_n1027 , 1_n1028 , 1_n1029 , 1_n1030 , 1_n1031 , 1_n1032 , 1_n1033 , 1_n1034 , 1_n1035 , 1_n1036 , 1_n1037 , 1_n1038 , 1_n1039 , 1_n1040 , 1_n1041 , 1_n1042 , 1_n1043 , 1_n1044 , 1_n1045 , 1_n1046 , 1_n1047 , 1_n1048 , 1_n1049 , 1_n1050 , 1_n1051 , 1_n1052 , 1_n1053 , 1_n1054 , 1_n1055 , 1_n1056 , 1_n1057 , 1_n1058 , 1_n1059 , 1_n1060 , 1_n1061 , 1_n1062 , 1_n1063 , 1_n1064 , 1_n1065 , 1_n1066 , 1_n1067 , 1_n1068 , 1_n1069 , 1_n1070 , 1_n1071 , 1_n1072 , 1_n1073 , 1_n1074 , 1_n1075 , 1_n1076 , 1_n1077 , 1_n1078 , 1_n1079 , 1_n1080 , 1_n1081 , 1_n1082 , 1_n1083 , 1_n1085 , 1_n1086 , 1_n1087 , 1_n1088 , 1_n1089 , 1_n1090 , 1_n1091 , 1_n1092 , 1_n1093 , 1_n1094 , 1_n1095 , 1_n1096 , 1_n1098 , 1_n1099 , 1_n1100 , 1_n1101 , 1_n1102 , 1_n1103 , 1_n1104 , 1_n1105 , 1_n1106 , 1_n1107 , 1_n1108 , 1_n1109 , 1_n1110 , 1_n1111 , 1_n1113 , 1_n1114 , 1_n1115 , 1_n1116 , 1_n1117 , 1_n1118 , 1_n1119 , 1_n1120 , 1_n1121 , 1_n1122 , 1_n1123 , 1_n1124 , 1_n1125 , 1_n1126 , 1_n1127 , 1_n1128 , 1_n1129 , 1_n1130 , 1_n1131 , 1_n1132 , 1_n1133 , 1_n1134 , 1_n1135 , 1_n1136 , 1_n1137 , 1_n1138 , 1_n1139 , 1_n1140 , 1_n1141 , 1_n1142 , 1_n1143 , 1_n1144 , 1_n1145 , 1_n1146 , 1_n1147 , 1_n1148 , 1_n1149 , 1_n1150 , 1_n1151 , 1_n1152 , 1_n1153 , 1_n1154 , 1_n1155 , 1_n1156 , 1_n1157 , 1_n1158 , 1_n1159 , 1_n1160 , 1_n1161 , 1_n1162 , 1_n1163 , 1_n1164 , 1_n1166 , 1_n1167 , 1_n1168 , 1_n1169 , 1_n1170 , 1_n1171 , 1_n1172 , 1_n1173 , 1_n1174 , 1_n1175 , 1_n1176 , 1_n1177 , 1_n1178 , 1_n1179 , 1_n1180 , 1_n1182 , 1_n1183 , 1_n1184 , 1_n1185 , 1_n1186 , 1_n1187 , 1_n1188 , 1_n1189 , 1_n1190 , 1_n1191 , 1_n1192 , 1_n1193 , 1_n1194 , 1_n1195 , 1_n1196 , 1_n1197 , 1_n1199 , 1_n1200 , 1_n1201 , 1_n1202 , 1_n1203 , 1_n1204 , 1_n1205 , 1_n1206 , 1_n1207 , 1_n1208 , 1_n1209 , 1_n1210 , 1_n1211 , 1_n1212 , 1_n1213 , 1_n1214 , 1_n1215 , 1_n1216 , 1_n1217 , 1_n1218 , 1_n1219 , 1_n1220 , 1_n1221 , 1_n1222 , 1_n1223 , 1_n1224 , 1_n1225 , 1_n1226 , 1_n1227 , 1_n1228 , 1_n1229 , 1_n1230 , 1_n1232 , 1_n1233 , 1_n1234 , 1_n1235 , 1_n1236 , 1_n1237 , 1_n1238 , 1_n1239 , 1_n1240 , 1_n1241 , 1_n1242 , 1_n1243 , 1_n1244 , 1_n1245 , 1_n1246 , 1_n1247 , 1_n1248 , 1_n1249 , 1_n1250 , 1_n1251 , 1_n1252 , 1_n1253 , 1_n1254 , 1_n1255 , 1_n1256 , 1_n1257 , 1_n1258 , 1_n1259 , 1_n1260 , 1_n1261 , 1_n1262 , 1_n1263 , 1_n1264 , 1_n1265 , 1_n1266 , 1_n1267 , 1_n1268 , 1_n1269 , 1_n1270 , 1_n1271 , 1_n1272 , 1_n1273 , 1_n1274 , 1_n1275 , 1_n1276 , 1_n1277 , 1_n1278 , 1_n1279 , 1_n1280 , 1_n1281 , 1_n1282 , 1_n1283 , 1_n1284 , 1_n1285 , 1_n1286 , 1_n1287 , 1_n1288 , 1_n1289 , 1_n1290 , 1_n1291 , 1_n1292 , 1_n1293 , 1_n1294 , 1_n1295 , 1_n1296 , 1_n1297 , 1_n1298 , 1_n1299 , 1_n1300 , 1_n1301 , 1_n1303 , 1_n1304 , 1_n1305 , 1_n1306 , 1_n1308 , 1_n1309 , 1_n1310 , 1_n1311 , 1_n1312 , 1_n1313 , 1_n1314 , 1_n1315 , 1_n1316 , 1_n1317 , 1_n1318 , 1_n1319 , 1_n1320 , 1_n1321 , 1_n1322 , 1_n1323 , 1_n1324 , 1_n1325 , 1_n1326 , 1_n1327 , 1_n1328 , 1_n1329 , 1_n1330 , 1_n1331 , 1_n1332 , 1_n1333 , 1_n1334 , 1_n1335 , 1_n1336 , 1_n1337 , 1_n1338 , 1_n1339 , 1_n1340 , 1_n1341 , 1_n1342 , 1_n1343 , 1_n1344 , 1_n1345 , 1_n1346 , 1_n1347 , 1_n1348 , 1_n1349 , 1_n1350 , 1_n1351 , 1_n1352 , 1_n1353 , 1_n1354 , 1_n1355 , 1_n1356 , 1_n1357 , 1_n1358 , 1_n1359 , 1_n1360 , 1_n1361 , 1_n1362 , 1_n1363 , 1_n1365 , 1_n1366 , 1_n1367 , 1_n1368 , 1_n1369 , 1_n1370 , 1_n1371 , 1_n1372 , 1_n1373 , 1_n1374 , 1_n1375 , 1_n1376 , 1_n1377 , 1_n1378 , 1_n1379 , 1_n1380 , 1_n1381 , 1_n1382 , 1_n1383 , 1_n1384 , 1_n1385 , 1_n1386 , 1_n1387 , 1_n1388 , 1_n1389 , 1_n1390 , 1_n1391 , 1_n1393 , 1_n1394 , 1_n1395 , 1_n1396 , 1_n1397 , 1_n1398 , 1_n1399 , 1_n1400 , 1_n1402 , 1_n1403 , 1_n1404 , 1_n1405 , 1_n1406 , 1_n1407 , 1_n1408 , 1_n1409 , 1_n1410 , 1_n1411 , 1_n1412 , 1_n1413 , 1_n1414 , 1_n1415 , 1_n1416 , 1_n1417 , 1_n1418 , 1_n1419 , 1_n1420 , 1_n1421 , 1_n1422 , 1_n1423 , 1_n1424 , 1_n1425 , 1_n1426 , 1_n1427 , 1_n1428 , 1_n1429 , 1_n1430 , 1_n1431 , 1_n1432 , 1_n1433 , 1_n1434 , 1_n1435 , 1_n1436 , 1_n1437 , 1_n1438 , 1_n1439 , 1_n1440 , 1_n1441 , 1_n1442 , 1_n1443 , 1_n1444 , 1_n1445 , 1_n1446 , 1_n1447 , 1_n1448 , 1_n1449 , 1_n1450 , 1_n1451 , 1_n1452 , 1_n1453 , 1_n1454 , 1_n1455 , 1_n1456 , 1_n1457 , 1_n1458 , 1_n1459 , 1_n1460 , 1_n1461 , 1_n1462 , 1_n1463 , 1_n1464 , 1_n1465 , 1_n1466 , 1_n1467 , 1_n1468 , 1_n1469 , 1_n1470 , 1_n1471 , 1_n1472 , 1_n1473 , 1_n1474 , 1_n1475 , 1_n1476 , 1_n1477 , 1_n1478 , 1_n1479 , 1_n1480 , 1_n1481 , 1_n1482 , 1_n1483 , 1_n1484 , 1_n1485 , 1_n1486 , 1_n1488 , 1_n1489 , 1_n1490 , 1_n1491 , 1_n1492 , 1_n1493 , 1_n1494 , 1_n1495 , 1_n1496 , 1_n1497 , 1_n1498 , 1_n1499 , 1_n1500 , 1_n1501 , 1_n1502 , 1_n1503 , 1_n1504 , 1_n1505 , 1_n1506 , 1_n1507 , 1_n1508 , 1_n1509 , 1_n1510 , 1_n1511 , 1_n1512 , 1_n1513 , 1_n1514 , 1_n1515 , 1_n1516 , 1_n1517 , 1_n1518 , 1_n1519 , 1_n1520 , 1_n1521 , 1_n1522 , 1_n1523 , 1_n1524 , 1_n1525 , 1_n1526 , 1_n1527 , 1_n1528 , 1_n1529 , 1_n1530 , 1_n1531 , 1_n1532 , 1_n1533 , 1_n1534 , 1_n1535 , 1_n1536 , 1_n1537 , 1_n1538 , 1_n1539 , 1_n1540 , 1_n1541 , 1_n1542 , 1_n1543 , 1_n1544 , 1_n1545 , 1_n1546 , 1_n1547 , 1_n1548 , 1_n1549 , 1_n1550 , 1_n1551 , 1_n1552 , 1_n1553 , 1_n1554 , 1_n1555 , 1_n1556 , 1_n1557 , 1_n1558 , 1_n1559 , 1_n1560 , 1_n1562 , 1_n1563 , 1_n1564 , 1_n1565 , 1_n1566 , 1_n1567 , 1_n1568 , 1_n1569 , 1_n1570 , 1_n1571 , 1_n1572 , 1_n1573 , 1_n1574 , 1_n1575 , 1_n1576 , 1_n1577 , 1_n1578 , 1_n1579 , 1_n1580 , 1_n1581 , 1_n1582 , 1_n1583 , 1_n1584 , 1_n1585 , 1_n1586 , 1_n1587 , 1_n1588 , 1_n1589 , 1_n1590 , 1_n1591 , 1_n1592 , 1_n1593 , 1_n1594 , 1_n1595 , 1_n1596 , 1_n1597 , 1_n1598 , 1_n1599 , 1_n1600 , 1_n1601 , 1_n1602 , 1_n1603 , 1_n1604 , 1_n1605 , 1_n1606 , 1_n1607 , 1_n1608 , 1_n1609 , 1_n1610 , 1_n1611 , 1_n1612 , 1_n1613 , 1_n1614 , 1_n1615 , 1_n1616 , 1_n1617 , 1_n1618 , 1_n1619 , 1_n1620 , 1_n1621 , 1_n1622 , 1_n1623 , 1_n1624 , 1_n1625 , 1_n1626 , 1_n1627 , 1_n1628 , 1_n1629 , 1_n1630 , 1_n1631 , 1_n1632 , 1_n1633 , 1_n1634 , 1_n1635 , 1_n1637 , 1_n1638 , 1_n1639 , 1_n1640 , 1_n1641 , 1_n1642 , 1_n1643 , 1_n1644 , 1_n1645 , 1_n1646 , 1_n1647 , 1_n1648 , 1_n1649 , 1_n1651 , 1_n1652 , 1_n1653 , 1_n1654 , 1_n1655 , 1_n1656 , 1_n1657 , 1_n1658 , 1_n1659 , 1_n1660 , 1_n1661 , 1_n1662 , 1_n1663 , 1_n1664 , 1_n1665 , 1_n1666 , 1_n1667 , 1_n1668 , 1_n1669 , 1_n1670 , 1_n1671 , 1_n1672 , 1_n1673 , 1_n1674 , 1_n1675 , 1_n1676 , 1_n1677 , 1_n1678 , 1_n1679 , 1_n1680 , 1_n1681 , 1_n1682 , 1_n1683 , 1_n1684 , 1_n1685 , 1_n1686 , 1_n1687 , 1_n1688 , 1_n1689 , 1_n1690 , 1_n1691 , 1_n1692 , 1_n1693 , 1_n1694 , 1_n1695 , 1_n1696 , 1_n1697 , 1_n1698 , 1_n1699 , 1_n1700 , 1_n1701 , 1_n1702 , 1_n1703 , 1_n1704 , 1_n1705 , 1_n1706 , 1_n1707 , 1_n1708 , 1_n1710 , 1_n1711 , 1_n1712 , 1_n1713 , 1_n1714 , 1_n1715 , 1_n1716 , 1_n1717 , 1_n1718 , 1_n1719 , 1_n1720 , 1_n1721 , 1_n1722 , 1_n1723 , 1_n1725 , 1_n1726 , 1_n1727 , 1_n1728 , 1_n1729 , 1_n1730 , 1_n1731 , 1_n1732 , 1_n1733 , 1_n1734 , 1_n1735 , 1_n1736 , 1_n1737 , 1_n1738 , 1_n1739 , 1_n1740 , 1_n1741 , 1_n1742 , 1_n1743 , 1_n1744 , 1_n1745 , 1_n1746 , 1_n1747 , 1_n1748 , 1_n1749 , 1_n1750 , 1_n1751 , 1_n1752 , 1_n1753 , 1_n1754 , 1_n1755 , 1_n1756 , 1_n1758 , 1_n1759 , 1_n1760 , 1_n1761 , 1_n1762 , 1_n1763 , 1_n1764 , 1_n1765 , 1_n1766 , 1_n1767 , 1_n1768 , 1_n1769 , 1_n1770 , 1_n1771 , 1_n1772 , 1_n1773 , 1_n1774 , 1_n1775 , 1_n1776 , 1_n1777 , 1_n1778 , 1_n1779 , 1_n1780 , 1_n1781 , 1_n1782 , 1_n1783 , 1_n1784 , 1_n1785 , 1_n1786 , 1_n1787 , 1_n1788 , 1_n1789 , 1_n1790 , 1_n1791 , 1_n1792 , 1_n1793 , 1_n1794 , 1_n1795 , 1_n1796 , 1_n1797 , 1_n1798 , 1_n1799 , 1_n1800 , 1_n1801 , 1_n1802 , 1_n1803 , 1_n1804 , 1_n1805 , 1_n1807 , 1_n1808 , 1_n1809 , 1_n1810 , 1_n1811 , 1_n1812 , 1_n1813 , 1_n1814 , 1_n1815 , 1_n1816 , 1_n1817 , 1_n1818 , 1_n1819 , 1_n1820 , 1_n1821 , 1_n1822 , 1_n1823 , 1_n1824 , 1_n1825 , 1_n1826 , 1_n1827 , 1_n1828 , 1_n1829 , 1_n1830 , 1_n1831 , 1_n1832 , 1_n1833 , 1_n1834 , 1_n1835 , 1_n1836 , 1_n1837 , 1_n1838 , 1_n1839 , 1_n1840 , 1_n1841 , 1_n1842 , 1_n1843 , 1_n1844 , 1_n1845 , 1_n1846 , 1_n1847 , 1_n1848 , 1_n1849 , 1_n1850 , 1_n1851 , 1_n1852 , 1_n1853 , 1_n1854 , 1_n1855 , 1_n1856 , 1_n1857 , 1_n1858 , 1_n1859 , 1_n1861 , 1_n1862 , 1_n1863 , 1_n1864 , 1_n1865 , 1_n1866 , 1_n1867 , 1_n1868 , 1_n1869 , 1_n1870 , 1_n1871 , 1_n1872 , 1_n1873 , 1_n1874 , 1_n1875 , 1_n1876 , 1_n1877 , 1_n1878 , 1_n1879 , 1_n1880 , 1_n1881 , 1_n1882 , 1_n1883 , 1_n1884 , 1_n1885 , 1_n1886 , 1_n1887 , 1_n1888 , 1_n1889 , 1_n1890 , 1_n1891 , 1_n1892 , 1_n1893 , 1_n1894 , 1_n1895 , 1_n1896 , 1_n1897 , 1_n1898 , 1_n1899 , 1_n1900 , 1_n1901 , 1_n1902 , 1_n1903 , 1_n1904 , 1_n1905 , 1_n1906 , 1_n1907 , 1_n1908 , 1_n1909 , 1_n1910 , 1_n1911 , 1_n1913 , 1_n1914 , 1_n1915 , 1_n1917 , 1_n1918 , 1_n1919 , 1_n1920 , 1_n1921 , 1_n1922 , 1_n1923 , 1_n1924 , 1_n1925 , 1_n1926 , 1_n1927 , 1_n1928 , 1_n1929 , 1_n1930 , 1_n1931 , 1_n1932 , 1_n1933 , 1_n1934 , 1_n1935 , 1_n1936 , 1_n1938 , 1_n1939 , 1_n1940 , 1_n1941 , 1_n1942 , 1_n1943 , 1_n1944 , 1_n1945 , 1_n1946 , 1_n1947 , 1_n1948 , 1_n1949 , 1_n1950 , 1_n1951 , 1_n1952 , 1_n1953 , 1_n1954 , 1_n1955 , 1_n1956 , 1_n1957 , 1_n1958 , 1_n1959 , 1_n1960 , 1_n1961 , 1_n1962 , 1_n1963 , 1_n1964 , 1_n1965 , 1_n1966 , 1_n1967 , 1_n1968 , 1_n1969 , 1_n1970 , 1_n1971 , 1_n1972 , 1_n1973 , 1_n1974 , 1_n1975 , 1_n1976 , 1_n1977 , 1_n1978 , 1_n1979 , 1_n1980 , 1_n1981 , 1_n1983 , 1_n1984 , 1_n1985 , 1_n1986 , 1_n1987 , 1_n1988 , 1_n1989 , 1_n1990 , 1_n1991 , 1_n1992 , 1_n1993 , 1_n1994 , 1_n1995 , 1_n1996 , 1_n1997 , 1_n1998 , 1_n1999 , 1_n2000 , 1_n2001 , 1_n2002 , 1_n2003 , 1_n2004 , 1_n2005 , 1_n2006 , 1_n2007 , 1_n2008 , 1_n2009 , 1_n2010 , 1_n2011 , 1_n2012 , 1_n2013 , 1_n2014 , 1_n2015 , 1_n2016 , 1_n2017 , 1_n2018 , 1_n2019 , 1_n2020 , 1_n2021 , 1_n2022 , 1_n2023 , 1_n2024 , 1_n2025 , 1_n2026 , 1_n2027 , 1_n2028 , 1_n2029 , 1_n2030 , 1_n2031 , 1_n2032 , 1_n2033 , 1_n2034 , 1_n2035 , 1_n2036 , 1_n2037 , 1_n2038 , 1_n2039 , 1_n2040 , 1_n2041 , 1_n2042 , 1_n2043 , 1_n2044 , 1_n2045 , 1_n2046 , 1_n2047 , 1_n2048 , 1_n2049 , 1_n2050 , 1_n2051 , 1_n2052 , 1_n2053 , 1_n2054 , 1_n2055 , 1_n2056 , 1_n2058 , 1_n2059 , 1_n2060 , 1_n2062 , 1_n2063 , 1_n2064 , 1_n2065 , 1_n2066 , 1_n2067 , 1_n2069 , 1_n2070 , 1_n2071 , 1_n2072 , 1_n2073 , 1_n2074 , 1_n2075 , 1_n2076 , 1_n2077 , 1_n2078 , 1_n2079 , 1_n2080 , 1_n2081 , 1_n2082 , 1_n2083 , 1_n2084 , 1_n2085 , 1_n2086 , 1_n2087 , 1_n2088 , 1_n2089 , 1_n2090 , 1_n2091 , 1_n2092 , 1_n2093 , 1_n2094 , 1_n2095 , 1_n2096 , 1_n2097 , 1_n2098 , 1_n2099 , 1_n2100 , 1_n2101 , 1_n2102 , 1_n2103 , 1_n2104 , 1_n2105 , 1_n2106 , 1_n2107 , 1_n2108 , 1_n2109 , 1_n2110 , 1_n2111 , 1_n2112 , 1_n2113 , 1_n2114 , 1_n2115 , 1_n2116 , 1_n2117 , 1_n2118 , 1_n2119 , 1_n2120 , 1_n2121 , 1_n2122 , 1_n2123 , 1_n2124 , 1_n2125 , 1_n2126 , 1_n2127 , 1_n2128 , 1_n2129 , 1_n2130 , 1_n2131 , 1_n2132 , 1_n2133 , 1_n2134 , 1_n2135 , 1_n2136 , 1_n2137 , 1_n2138 , 1_n2139 , 1_n2140 , 1_n2141 , 1_n2142 , 1_n2143 , 1_n2144 , 1_n2145 , 1_n2146 , 1_n2147 , 1_n2148 , 1_n2149 , 1_n2150 , 1_n2151 , 1_n2152 , 1_n2153 , 1_n2154 , 1_n2155 , 1_n2156 , 1_n2157 , 1_n2158 , 1_n2159 , 1_n2160 , 1_n2161 , 1_n2162 , 1_n2163 , 1_n2164 , 1_n2165 , 1_n2166 , 1_n2167 , 1_n2168 , 1_n2169 , 1_n2170 , 1_n2171 , 1_n2172 , 1_n2173 , 1_n2175 , 1_n2176 , 1_n2177 , 1_n2178 , 1_n2179 , 1_n2180 , 1_n2181 , 1_n2182 , 1_n2183 , 1_n2184 , 1_n2185 , 1_n2186 , 1_n2187 , 1_n2188 , 1_n2189 , 1_n2191 , 1_n2192 , 1_n2193 , 1_n2194 , 1_n2195 , 1_n2196 , 1_n2197 , 1_n2198 , 1_n2199 , 1_n2200 , 1_n2201 , 1_n2202 , 1_n2203 , 1_n2204 , 1_n2205 , 1_n2206 , 1_n2207 , 1_n2208 , 1_n2209 , 1_n2210 , 1_n2211 , 1_n2212 , 1_n2213 , 1_n2214 , 1_n2215 , 1_n2216 , 1_n2217 , 1_n2218 , 1_n2219 , 1_n2220 , 1_n2221 , 1_n2222 , 1_n2223 , 1_n2224 , 1_n2225 , 1_n2226 , 1_n2227 , 1_n2228 , 1_n2229 , 1_n2230 , 1_n2231 , 1_n2232 , 1_n2233 , 1_n2234 , 1_n2236 , 1_n2237 , 1_n2238 , 1_n2239 , 1_n2240 , 1_n2241 , 1_n2242 , 1_n2243 , 1_n2244 , 1_n2245 , 1_n2246 , 1_n2247 , 1_n2248 , 1_n2249 , 1_n2250 , 1_n2251 , 1_n2253 , 1_n2254 , 1_n2255 , 1_n2256 , 1_n2257 , 1_n2258 , 1_n2259 , 1_n2260 , 1_n2261 , 1_n2262 , 1_n2263 , 1_n2264 , 1_n2265 , 1_n2266 , 1_n2267 , 1_n2268 , 1_n2269 , 1_n2270 , 1_n2271 , 1_n2272 , 1_n2273 , 1_n2274 , 1_n2275 , 1_n2276 , 1_n2277 , 1_n2278 , 1_n2279 , 1_n2280 , 1_n2281 , 1_n2282 , 1_n2283 , 1_n2284 , 1_n2285 , 1_n2286 , 1_n2287 , 1_n2288 , 1_n2289 , 1_n2290 , 1_n2291 , 1_n2292 , 1_n2293 , 1_n2294 , 1_n2296 , 1_n2297 , 1_n2298 , 1_n2299 , 1_n2300 , 1_n2301 , 1_n2302 , 1_n2303 , 1_n2304 , 1_n2305 , 1_n2306 , 1_n2307 , 1_n2308 , 1_n2309 , 1_n2310 , 1_n2311 , 1_n2312 , 1_n2313 , 1_n2314 , 1_n2315 , 1_n2316 , 1_n2317 , 1_n2318 , 1_n2319 , 1_n2320 , 1_n2321 , 1_n2322 , 1_n2323 , 1_n2324 , 1_n2325 , 1_n2326 , 1_n2327 , 1_n2328 , 1_n2329 , 1_n2330 , 1_n2331 , 1_n2332 , 1_n2333 , 1_n2334 , 1_n2335 , 1_n2336 , 1_n2337 , 1_n2338 , 1_n2340 , 1_n2342 , 1_n2343 , 1_n2344 , 1_n2345 , 1_n2346 , 1_n2347 , 1_n2348 , 1_n2349 , 1_n2350 , 1_n2351 , 1_n2352 , 1_n2353 , 1_n2354 , 1_n2355 , 1_n2356 , 1_n2357 , 1_n2358 , 1_n2359 , 1_n2360 , 1_n2361 , 1_n2362 , 1_n2363 , 1_n2364 , 1_n2365 , 1_n2366 , 1_n2367 , 1_n2368 , 1_n2369 , 1_n2370 , 1_n2371 , 1_n2372 , 1_n2373 , 1_n2374 , 1_n2375 , 1_n2376 , 1_n2377 , 1_n2378 , 1_n2379 , 1_n2380 , 1_n2381 , 1_n2382 , 1_n2383 , 1_n2384 , 1_n2385 , 1_n2386 , 1_n2387 , 1_n2388 , 1_n2389 , 1_n2390 , 1_n2391 , 1_n2392 , 1_n2393 , 1_n2394 , 1_n2395 , 1_n2396 , 1_n2397 , 1_n2398 , 1_n2399 , 1_n2400 , 1_n2401 , 1_n2402 , 1_n2403 , 1_n2404 , 1_n2405 , 1_n2406 , 1_n2407 , 1_n2408 , 1_n2409 , 1_n2410 , 1_n2411 , 1_n2412 , 1_n2413 , 1_n2414 , 1_n2415 , 1_n2416 , 1_n2417 , 1_n2418 , 1_n2419 , 1_n2420 , 1_n2421 , 1_n2422 , 1_n2423 , 1_n2424 , 1_n2425 , 1_n2426 , 1_n2427 , 1_n2428 , 1_n2429 , 1_n2430 , 1_n2431 , 1_n2432 , 1_n2433 , 1_n2434 , 1_n2435 , 1_n2436 , 1_n2437 , 1_n2438 , 1_n2439 , 1_n2440 , 1_n2441 , 1_n2442 , 1_n2443 , 1_n2444 , 1_n2445 , 1_n2446 , 1_n2447 , 1_n2448 , 1_n2449 , 1_n2450 , 1_n2451 , 1_n2452 , 1_n2453 , 1_n2454 , 1_n2455 , 1_n2456 , 1_n2457 , 1_n2459 , 1_n2460 , 1_n2461 , 1_n2462 , 1_n2463 , 1_n2464 , 1_n2465 , 1_n2466 , 1_n2467 , 1_n2468 , 1_n2469 , 1_n2470 , 1_n2471 , 1_n2472 , 1_n2473 , 1_n2474 , 1_n2475 , 1_n2476 , 1_n2477 , 1_n2478 , 1_n2479 , 1_n2480 , 1_n2481 , 1_n2483 , 1_n2484 , 1_n2485 , 1_n2486 , 1_n2487 , 1_n2488 , 1_n2489 , 1_n2490 , 1_n2491 , 1_n2492 , 1_n2493 , 1_n2494 , 1_n2495 , 1_n2496 , 1_n2497 , 1_n2499 , 1_n2500 , 1_n2501 , 1_n2502 , 1_n2503 , 1_n2504 , 1_n2505 , 1_n2506 , 1_n2507 , 1_n2508 , 1_n2509 , 1_n2510 , 1_n2511 , 1_n2512 , 1_n2513 , 1_n2514 , 1_n2515 , 1_n2516 , 1_n2517 , 1_n2518 , 1_n2519 , 1_n2520 , 1_n2521 , 1_n2522 , 1_n2523 , 1_n2524 , 1_n2525 , 1_n2526 , 1_n2527 , 1_n2528 , 1_n2529 , 1_n2530 , 1_n2531 , 1_n2532 , 1_n2533 , 1_n2534 , 1_n2535 , 1_n2536 , 1_n2537 , 1_n2538 , 1_n2539 , 1_n2540 , 1_n2541 , 1_n2542 , 1_n2543 , 1_n2544 , 1_n2545 , 1_n2546 , 1_n2547 , 1_n2548 , 1_n2550 , 1_n2551 , 1_n2552 , 1_n2553 , 1_n2554 , 1_n2555 , 1_n2556 , 1_n2557 , 1_n2558 , 1_n2559 , 1_n2560 , 1_n2561 , 1_n2562 , 1_n2563 , 1_n2564 , 1_n2565 , 1_n2566 , 1_n2567 , 1_n2568 , 1_n2569 , 1_n2570 , 1_n2571 , 1_n2572 , 1_n2573 , 1_n2574 , 1_n2575 , 1_n2576 , 1_n2577 , 1_n2578 , 1_n2579 , 1_n2580 , 1_n2581 , 1_n2582 , 1_n2583 , 1_n2584 , 1_n2585 , 1_n2586 , 1_n2587 , 1_n2588 , 1_n2589 , 1_n2591 , 1_n2593 , 1_n2594 , 1_n2595 , 1_n2596 , 1_n2597 , 1_n2598 , 1_n2599 , 1_n2600 , 1_n2601 , 1_n2602 , 1_n2603 , 1_n2604 , 1_n2605 , 1_n2606 , 1_n2607 , 1_n2608 , 1_n2609 , 1_n2610 , 1_n2611 , 1_n2612 , 1_n2613 , 1_n2614 , 1_n2615 , 1_n2616 , 1_n2617 , 1_n2618 , 1_n2619 , 1_n2620 , 1_n2621 , 1_n2622 , 1_n2623 , 1_n2624 , 1_n2625 , 1_n2626 , 1_n2627 , 1_n2628 , 1_n2629 , 1_n2630 , 1_n2631 , 1_n2632 , 1_n2633 , 1_n2634 , 1_n2635 , 1_n2636 , 1_n2637 , 1_n2638 , 1_n2639 , 1_n2640 , 1_n2641 , 1_n2642 , 1_n2643 , 1_n2644 , 1_n2645 , 1_n2646 , 1_n2647 , 1_n2648 , 1_n2649 , 1_n2650 , 1_n2651 , 1_n2652 , 1_n2653 , 1_n2654 , 1_n2655 , 1_n2656 , 1_n2657 , 1_n2658 , 1_n2659 , 1_n2660 , 1_n2661 , 1_n2662 , 1_n2663 , 1_n2664 , 1_n2665 , 1_n2667 , 1_n2668 , 1_n2669 , 1_n2670 , 1_n2671 , 1_n2672 , 1_n2673 , 1_n2674 , 1_n2675 , 1_n2676 , 1_n2677 , 1_n2678 , 1_n2679 , 1_n2680 , 1_n2681 , 1_n2682 , 1_n2683 , 1_n2684 , 1_n2685 , 1_n2686 , 1_n2687 , 1_n2688 , 1_n2689 , 1_n2690 , 1_n2691 , 1_n2692 , 1_n2693 , 1_n2694 , 1_n2695 , 1_n2696 , 1_n2697 , 1_n2698 , 1_n2699 , 1_n2700 , 1_n2701 , 1_n2702 , 1_n2703 , 1_n2704 , 1_n2705 , 1_n2706 , 1_n2707 , 1_n2708 , 1_n2710 , 1_n2711 , 1_n2712 , 1_n2713 , 1_n2714 , 1_n2715 , 1_n2716 , 1_n2717 , 1_n2718 , 1_n2719 , 1_n2720 , 1_n2721 , 1_n2722 , 1_n2723 , 1_n2724 , 1_n2725 , 1_n2726 , 1_n2727 , 1_n2728 , 1_n2729 , 1_n2730 , 1_n2731 , 1_n2732 , 1_n2733 , 1_n2734 , 1_n2735 , 1_n2736 , 1_n2738 , 1_n2739 , 1_n2740 , 1_n2741 , 1_n2742 , 1_n2743 , 1_n2744 , 1_n2745 , 1_n2746 , 1_n2747 , 1_n2748 , 1_n2749 , 1_n2750 , 1_n2751 , 1_n2752 , 1_n2753 , 1_n2754 , 1_n2755 , 1_n2756 , 1_n2757 , 1_n2759 , 1_n2760 , 1_n2761 , 1_n2762 , 1_n2763 , 1_n2764 , 1_n2765 , 1_n2766 , 1_n2767 , 1_n2768 , 1_n2769 , 1_n2770 , 1_n2772 , 1_n2773 , 1_n2774 , 1_n2775 , 1_n2776 , 1_n2778 , 1_n2779 , 1_n2780 , 1_n2781 , 1_n2782 , 1_n2783 , 1_n2784 , 1_n2785 , 1_n2786 , 1_n2787 , 1_n2788 , 1_n2789 , 1_n2790 , 1_n2791 , 1_n2792 , 1_n2793 , 1_n2794 , 1_n2795 , 1_n2796 , 1_n2797 , 1_n2798 , 1_n2799 , 1_n2800 , 1_n2801 , 1_n2802 , 1_n2803 , 1_n2804 , 1_n2806 , 1_n2807 , 1_n2808 , 1_n2809 , 1_n2810 , 1_n2811 , 1_n2812 , 1_n2813 , 1_n2814 , 1_n2815 , 1_n2816 , 1_n2817 , 1_n2818 , 1_n2819 , 1_n2820 , 1_n2821 , 1_n2822 , 1_n2823 , 1_n2824 , 1_n2825 , 1_n2826 , 1_n2827 , 1_n2828 , 1_n2829 , 1_n2830 , 1_n2831 , 1_n2832 , 1_n2833 , 1_n2834 , 1_n2835 , 1_n2836 , 1_n2837 , 1_n2838 , 1_n2839 , 1_n2840 , 1_n2841 , 1_n2842 , 1_n2843 , 1_n2844 , 1_n2845 , 1_n2846 , 1_n2847 , 1_n2848 , 1_n2849 , 1_n2850 , 1_n2851 , 1_n2852 , 1_n2853 , 1_n2854 , 1_n2855 , 1_n2856 , 1_n2857 , 1_n2858 , 1_n2859 , 1_n2860 , 1_n2861 , 1_n2862 , 1_n2863 , 1_n2864 , 1_n2865 , 1_n2866 , 1_n2867 , 1_n2868 , 1_n2869 , 1_n2870 , 1_n2871 , 1_n2872 , 1_n2873 , 1_n2874 , 1_n2875 , 1_n2876 , 1_n2877 , 1_n2878 , 1_n2879 , 1_n2880 , 1_n2881 , 1_n2883 , 1_n2884 , 1_n2885 , 1_n2886 , 1_n2887 , 1_n2888 , 1_n2889 , 1_n2890 , 1_n2891 , 1_n2892 , 1_n2893 , 1_n2894 , 1_n2895 , 1_n2896 , 1_n2897 , 1_n2898 , 1_n2899 , 1_n2900 , 1_n2901 , 1_n2902 , 1_n2903 , 1_n2905 , 1_n2906 , 1_n2907 , 1_n2908 , 1_n2909 , 1_n2910 , 1_n2911 , 1_n2912 , 1_n2913 , 1_n2914 , 1_n2915 , 1_n2916 , 1_n2917 , 1_n2918 , 1_n2919 , 1_n2920 , 1_n2921 , 1_n2922 , 1_n2923 , 1_n2924 , 1_n2925 , 1_n2926 , 1_n2927 , 1_n2928 , 1_n2929 , 1_n2930 , 1_n2931 , 1_n2932 , 1_n2933 , 1_n2935 , 1_n2936 , 1_n2937 , 1_n2938 , 1_n2939 , 1_n2940 , 1_n2941 , 1_n2942 , 1_n2943 , 1_n2944 , 1_n2945 , 1_n2946 , 1_n2947 , 1_n2948 , 1_n2949 , 1_n2950 , 1_n2951 , 1_n2952 , 1_n2953 , 1_n2954 , 1_n2955 , 1_n2956 , 1_n2957 , 1_n2958 , 1_n2959 , 1_n2960 , 1_n2961 , 1_n2962 , 1_n2963 , 1_n2964 , 1_n2965 , 1_n2966 , 1_n2967 , 1_n2968 , 1_n2969 , 1_n2970 , 1_n2971 , 1_n2972 , 1_n2973 , 1_n2974 , 1_n2975 , 1_n2976 , 1_n2977 , 1_n2978 , 1_n2979 , 1_n2980 , 1_n2981 , 1_n2982 , 1_n2983 , 1_n2984 , 1_n2985 , 1_n2986 , 1_n2987 , 1_n2988 , 1_n2989 , 1_n2990 , 1_n2991 , 1_n2992 , 1_n2993 , 1_n2994 , 1_n2995 , 1_n2996 , 1_n2997 , 1_n2998 , 1_n2999 , 1_n3000 , 1_n3001 , 1_n3002 , 1_n3003 , 1_n3004 , 1_n3005 , 1_n3007 , 1_n3008 , 1_n3009 , 1_n3010 , 1_n3011 , 1_n3012 , 1_n3013 , 1_n3014 , 1_n3015 , 1_n3016 , 1_n3017 , 1_n3018 , 1_n3019 , 1_n3020 , 1_n3021 , 1_n3022 , 1_n3023 , 1_n3024 , 1_n3025 , 1_n3026 , 1_n3027 , 1_n3028 , 1_n3029 , 1_n3030 , 1_n3031 , 1_n3032 , 1_n3033 , 1_n3034 , 1_n3035 , 1_n3036 , 1_n3037 , 1_n3038 , 1_n3039 , 1_n3040 , 1_n3041 , 1_n3042 , 1_n3043 , 1_n3044 , 1_n3045 , 1_n3046 , 1_n3047 , 1_n3048 , 1_n3049 , 1_n3050 , 1_n3051 , 1_n3052 , 1_n3053 , 1_n3054 , 1_n3055 , 1_n3056 , 1_n3057 , 1_n3058 , 1_n3059 , 1_n3060 , 1_n3061 , 1_n3062 , 1_n3063 , 1_n3064 , 1_n3065 , 1_n3066 , 1_n3067 , 1_n3068 , 1_n3069 , 1_n3070 , 1_n3071 , 1_n3072 , 1_n3073 , 1_n3074 , 1_n3075 , 1_n3077 , 1_n3078 , 1_n3079 , 1_n3080 , 1_n3081 , 1_n3082 , 1_n3083 , 1_n3084 , 1_n3086 , 1_n3087 , 1_n3088 , 1_n3089 , 1_n3090 , 1_n3091 , 1_n3092 , 1_n3093 , 1_n3094 , 1_n3095 , 1_n3096 , 1_n3097 , 1_n3098 , 1_n3099 , 1_n3100 , 1_n3101 , 1_n3102 , 1_n3103 , 1_n3104 , 1_n3105 , 1_n3106 , 1_n3107 , 1_n3108 , 1_n3109 , 1_n3110 , 1_n3111 , 1_n3113 , 1_n3114 , 1_n3115 , 1_n3116 , 1_n3117 , 1_n3118 , 1_n3119 , 1_n3120 , 1_n3121 , 1_n3122 , 1_n3123 , 1_n3124 , 1_n3125 , 1_n3126 , 1_n3127 , 1_n3128 , 1_n3129 , 1_n3131 , 1_n3132 , 1_n3133 , 1_n3134 , 1_n3135 , 1_n3136 , 1_n3137 , 1_n3138 , 1_n3139 , 1_n3140 , 1_n3141 , 1_n3142 , 1_n3143 , 1_n3144 , 1_n3145 , 1_n3146 , 1_n3147 , 1_n3148 , 1_n3149 , 1_n3150 , 1_n3151 , 1_n3152 , 1_n3153 , 1_n3154 , 1_n3155 , 1_n3156 , 1_n3157 , 1_n3158 , 1_n3159 , 1_n3160 , 1_n3161 , 1_n3162 , 1_n3163 , 1_n3164 , 1_n3165 , 1_n3166 , 1_n3167 , 1_n3168 , 1_n3169 , 1_n3170 , 1_n3171 , 1_n3172 , 1_n3173 , 1_n3174 , 1_n3175 , 1_n3176 , 1_n3177 , 1_n3179 , 1_n3180 , 1_n3181 , 1_n3182 , 1_n3183 , 1_n3184 , 1_n3185 , 1_n3186 , 1_n3187 , 1_n3188 , 1_n3189 , 1_n3190 , 1_n3191 , 1_n3192 , 1_n3193 , 1_n3194 , 1_n3195 , 1_n3196 , 1_n3197 , 1_n3198 , 1_n3199 , 1_n3200 , 1_n3201 , 1_n3202 , 1_n3203 , 1_n3204 , 1_n3205 , 1_n3206 , 1_n3207 , 1_n3208 , 1_n3209 , 1_n3210 , 1_n3211 , 1_n3212 , 1_n3213 , 1_n3214 , 1_n3215 , 1_n3216 , 1_n3217 , 1_n3218 , 1_n3219 , 1_n3220 , 1_n3221 , 1_n3222 , 1_n3223 , 1_n3224 , 1_n3225 , 1_n3226 , 1_n3227 , 1_n3228 , 1_n3229 , 1_n3230 , 1_n3231 , 1_n3232 , 1_n3233 , 1_n3234 , 1_n3235 , 1_n3236 , 1_n3237 , 1_n3238 , 1_n3239 , 1_n3240 , 1_n3241 , 1_n3242 , 1_n3243 , 1_n3244 , 1_n3245 , 1_n3246 , 1_n3247 , 1_n3248 , 1_n3249 , 1_n3250 , 1_n3251 , 1_n3252 , 1_n3253 , 1_n3254 , 1_n3255 , 1_n3256 , 1_n3257 , 1_n3258 , 1_n3259 , 1_n3260 , 1_n3261 , 1_n3263 , 1_n3264 , 1_n3265 , 1_n3266 , 1_n3267 , 1_n3268 , 1_n3269 , 1_n3270 , 1_n3271 , 1_n3272 , 1_n3273 , 1_n3274 , 1_n3275 , 1_n3276 , 1_n3277 , 1_n3278 , 1_n3279 , 1_n3280 , 1_n3281 , 1_n3282 , 1_n3283 , 1_n3284 , 1_n3285 , 1_n3286 , 1_n3287 , 1_n3288 , 1_n3289 , 1_n3290 , 1_n3291 , 1_n3292 , 1_n3293 , 1_n3294 , 1_n3295 , 1_n3296 , 1_n3297 , 1_n3298 , 1_n3299 , 1_n3300 , 1_n3301 , 1_n3302 , 1_n3303 , 1_n3304 , 1_n3305 , 1_n3306 , 1_n3307 , 1_n3308 , 1_n3309 , 1_n3310 , 1_n3312 , 1_n3313 , 1_n3314 , 1_n3315 , 1_n3316 , 1_n3317 , 1_n3318 , 1_n3319 , 1_n3320 , 1_n3321 , 1_n3322 , 1_n3324 , 1_n3325 , 1_n3326 , 1_n3327 , 1_n3328 , 1_n3329 , 1_n3330 , 1_n3331 , 1_n3332 , 1_n3333 , 1_n3334 , 1_n3335 , 1_n3336 , 1_n3337 , 1_n3338 , 1_n3339 , 1_n3340 , 1_n3341 , 1_n3342 , 1_n3343 , 1_n3344 , 1_n3345 , 1_n3346 , 1_n3347 , 1_n3348 , 1_n3349 , 1_n3350 , 1_n3351 , 1_n3352 , 1_n3353 , 1_n3354 , 1_n3355 , 1_n3356 , 1_n3357 , 1_n3358 , 1_n3359 , 1_n3360 , 1_n3361 , 1_n3363 , 1_n3364 , 1_n3365 , 1_n3366 , 1_n3367 , 1_n3368 , 1_n3369 , 1_n3370 , 1_n3371 , 1_n3372 , 1_n3373 , 1_n3374 , 1_n3375 , 1_n3376 , 1_n3377 , 1_n3378 , 1_n3379 , 1_n3380 , 1_n3381 , 1_n3382 , 1_n3383 , 1_n3384 , 1_n3385 , 1_n3386 , 1_n3387 , 1_n3388 , 1_n3389 , 1_n3390 , 1_n3391 , 1_n3392 , 1_n3393 , 1_n3394 , 1_n3395 , 1_n3396 , 1_n3397 , 1_n3398 , 1_n3399 , 1_n3400 , 1_n3401 , 1_n3402 , 1_n3403 , 1_n3404 , 1_n3405 , 1_n3406 , 1_n3407 , 1_n3408 , 1_n3410 , 1_n3411 , 1_n3412 , 1_n3413 , 1_n3414 , 1_n3415 , 1_n3416 , 1_n3417 , 1_n3418 , 1_n3419 , 1_n3420 , 1_n3421 , 1_n3422 , 1_n3423 , 1_n3424 , 1_n3425 , 1_n3426 , 1_n3427 , 1_n3428 , 1_n3429 , 1_n3430 , 1_n3431 , 1_n3432 , 1_n3433 , 1_n3434 , 1_n3435 , 1_n3436 , 1_n3437 , 1_n3438 , 1_n3439 , 1_n3440 , 1_n3441 , 1_n3442 , 1_n3443 , 1_n3444 , 1_n3445 , 1_n3446 , 1_n3447 , 1_n3448 , 1_n3449 , 1_n3450 , 1_n3451 , 1_n3452 , 1_n3453 , 1_n3454 , 1_n3455 , 1_n3456 , 1_n3457 , 1_n3458 , 1_n3459 , 1_n3460 , 1_n3461 , 1_n3462 , 1_n3463 , 1_n3464 , 1_n3465 , 1_n3466 , 1_n3467 , 1_n3468 , 1_n3469 , 1_n3470 , 1_n3471 , 1_n3472 , 1_n3473 , 1_n3474 , 1_n3475 , 1_n3476 , 1_n3477 , 1_n3478 , 1_n3479 , 1_n3480 , 1_n3481 , 1_n3482 , 1_n3483 , 1_n3484 , 1_n3485 , 1_n3486 , 1_n3487 , 1_n3488 , 1_n3489 , 1_n3490 , 1_n3491 , 1_n3492 , 1_n3493 , 1_n3494 , 1_n3495 , 1_n3496 , 1_n3497 , 1_n3498 , 1_n3499 , 1_n3500 , 1_n3501 , 1_n3502 , 1_n3503 , 1_n3504 , 1_n3505 , 1_n3506 , 1_n3507 , 1_n3508 , 1_n3509 , 1_n3510 , 1_n3511 , 1_n3512 , 1_n3513 , 1_n3514 , 1_n3515 , 1_n3516 , 1_n3517 , 1_n3518 , 1_n3519 , 1_n3520 , 1_n3521 , 1_n3522 , 1_n3523 , 1_n3524 , 1_n3525 , 1_n3526 , 1_n3527 , 1_n3528 , 1_n3529 , 1_n3530 , 1_n3531 , 1_n3532 , 1_n3533 , 1_n3534 , 1_n3535 , 1_n3536 , 1_n3537 , 1_n3538 , 1_n3539 , 1_n3540 , 1_n3541 , 1_n3542 , 1_n3543 , 1_n3544 , 1_n3545 , 1_n3546 , 1_n3547 , 1_n3548 , 1_n3549 , 1_n3550 , 1_n3551 , 1_n3552 , 1_n3553 , 1_n3554 , 1_n3555 , 1_n3556 , 1_n3557 , 1_n3558 , 1_n3559 , 1_n3560 , 1_n3561 , 1_n3562 , 1_n3563 , 1_n3564 , 1_n3565 , 1_n3566 , 1_n3567 , 1_n3568 , 1_n3569 , 1_n3570 , 1_n3571 , 1_n3572 , 1_n3573 , 1_n3574 , 1_n3575 , 1_n3576 , 1_n3577 , 1_n3578 , 1_n3579 , 1_n3580 , 1_n3581 , 1_n3582 , 1_n3583 , 1_n3584 , 1_n3585 , 1_n3586 , 1_n3587 , 1_n3588 , 1_n3589 , 1_n3590 , 1_n3592 , 1_n3593 , 1_n3594 , 1_n3595 , 1_n3596 , 1_n3597 , 1_n3598 , 1_n3599 , 1_n3600 , 1_n3601 , 1_n3602 , 1_n3603 , 1_n3604 , 1_n3605 , 1_n3606 , 1_n3607 , 1_n3608 , 1_n3609 , 1_n3610 , 1_n3611 , 1_n3612 , 1_n3613 , 1_n3614 , 1_n3615 , 1_n3616 , 1_n3617 , 1_n3618 , 1_n3619 , 1_n3620 , 1_n3621 , 1_n3622 , 1_n3623 , 1_n3624 , 1_n3625 , 1_n3626 , 1_n3627 , 1_n3628 , 1_n3629 , 1_n3630 , 1_n3631 , 1_n3632 , 1_n3633 , 1_n3634 , 1_n3635 , 1_n3636 , 1_n3637 , 1_n3638 , 1_n3639 , 1_n3640 , 1_n3642 , 1_n3643 , 1_n3644 , 1_n3645 , 1_n3646 , 1_n3647 , 1_n3648 , 1_n3649 , 1_n3650 , 1_n3651 , 1_n3652 , 1_n3653 , 1_n3654 , 1_n3655 , 1_n3656 , 1_n3657 , 1_n3658 , 1_n3659 , 1_n3660 , 1_n3661 , 1_n3662 , 1_n3663 , 1_n3664 , 1_n3665 , 1_n3666 , 1_n3667 , 1_n3668 , 1_n3670 , 1_n3671 , 1_n3672 , 1_n3673 , 1_n3674 , 1_n3675 , 1_n3676 , 1_n3678 , 1_n3679 , 1_n3680 , 1_n3681 , 1_n3682 , 1_n3683 , 1_n3684 , 1_n3685 , 1_n3686 , 1_n3687 , 1_n3688 , 1_n3689 , 1_n3690 , 1_n3691 , 1_n3692 , 1_n3693 , 1_n3694 , 1_n3695 , 1_n3696 , 1_n3697 , 1_n3698 , 1_n3699 , 1_n3700 , 1_n3701 , 1_n3702 , 1_n3703 , 1_n3704 , 1_n3705 , 1_n3706 , 1_n3707 , 1_n3708 , 1_n3709 , 1_n3710 , 1_n3711 , 1_n3712 , 1_n3713 , 1_n3714 , 1_n3715 , 1_n3716 , 1_n3717 , 1_n3718 , 1_n3719 , 1_n3720 , 1_n3721 , 1_n3722 , 1_n3723 , 1_n3724 , 1_n3725 , 1_n3726 , 1_n3727 , 1_n3728 , 1_n3729 , 1_n3730 , 1_n3731 , 1_n3732 , 1_n3733 , 1_n3734 , 1_n3735 , 1_n3736 , 1_n3737 , 1_n3738 , 1_n3739 , 1_n3740 , 1_n3741 , 1_n3742 , 1_n3743 , 1_n3744 , 1_n3745 , 1_n3746 , 1_n3747 , 1_n3749 , 1_n3750 , 1_n3751 , 1_n3752 , 1_n3753 , 1_n3754 , 1_n3755 , 1_n3756 , 1_n3757 , 1_n3758 , 1_n3759 , 1_n3760 , 1_n3761 , 1_n3762 , 1_n3763 , 1_n3764 , 1_n3765 , 1_n3766 , 1_n3767 , 1_n3768 , 1_n3770 , 1_n3771 , 1_n3772 , 1_n3773 , 1_n3774 , 1_n3775 , 1_n3776 , 1_n3777 , 1_n3778 , 1_n3779 , 1_n3780 , 1_n3781 , 1_n3782 , 1_n3783 , 1_n3784 , 1_n3785 , 1_n3786 , 1_n3787 , 1_n3788 , 1_n3789 , 1_n3791 , 1_n3792 , 1_n3793 , 1_n3794 , 1_n3795 , 1_n3796 , 1_n3797 , 1_n3798 , 1_n3799 , 1_n3800 , 1_n3801 , 1_n3802 , 1_n3803 , 1_n3804 , 1_n3805 , 1_n3806 , 1_n3807 , 1_n3808 , 1_n3809 , 1_n3810 , 1_n3811 , 1_n3812 , 1_n3813 , 1_n3814 , 1_n3816 , 1_n3817 , 1_n3818 , 1_n3819 , 1_n3820 , 1_n3821 , 1_n3822 , 1_n3823 , 1_n3824 , 1_n3825 , 1_n3826 , 1_n3827 , 1_n3828 , 1_n3829 , 1_n3830 , 1_n3831 , 1_n3833 , 1_n3834 , 1_n3835 , 1_n3836 , 1_n3837 , 1_n3838 , 1_n3839 , 1_n3840 , 1_n3841 , 1_n3842 , 1_n3843 , 1_n3844 , 1_n3845 , 1_n3846 , 1_n3847 , 1_n3848 , 1_n3849 , 1_n3850 , 1_n3851 , 1_n3852 , 1_n3853 , 1_n3854 , 1_n3855 , 1_n3856 , 1_n3857 , 1_n3858 , 1_n3859 , 1_n3860 , 1_n3861 , 1_n3862 , 1_n3863 , 1_n3864 , 1_n3865 , 1_n3866 , 1_n3867 , 1_n3868 , 1_n3869 , 1_n3870 , 1_n3871 , 1_n3872 , 1_n3873 , 1_n3874 , 1_n3875 , 1_n3876 , 1_n3877 , 1_n3878 , 1_n3879 , 1_n3880 , 1_n3881 , 1_n3882 , 1_n3883 , 1_n3884 , 1_n3885 , 1_n3886 , 1_n3887 , 1_n3888 , 1_n3889 , 1_n3890 , 1_n3891 , 1_n3892 , 1_n3893 , 1_n3894 , 1_n3895 , 1_n3896 , 1_n3897 , 1_n3898 , 1_n3899 , 1_n3900 , 1_n3901 , 1_n3902 , 1_n3903 , 1_n3904 , 1_n3905 , 1_n3906 , 1_n3907 , 1_n3908 , 1_n3909 , 1_n3910 , 1_n3911 , 1_n3912 , 1_n3913 , 1_n3914 , 1_n3915 , 1_n3916 , 1_n3917 , 1_n3918 , 1_n3919 , 1_n3920 , 1_n3921 , 1_n3922 , 1_n3923 , 1_n3924 , 1_n3925 , 1_n3926 , 1_n3927 , 1_n3928 , 1_n3929 , 1_n3930 , 1_n3931 , 1_n3932 , 1_n3933 , 1_n3934 , 1_n3935 , 1_n3936 , 1_n3937 , 1_n3938 , 1_n3939 , 1_n3940 , 1_n3941 , 1_n3942 , 1_n3943 , 1_n3944 , 1_n3945 , 1_n3947 , 1_n3948 , 1_n3949 , 1_n3950 , 1_n3951 , 1_n3952 , 1_n3953 , 1_n3954 , 1_n3955 , 1_n3956 , 1_n3957 , 1_n3958 , 1_n3959 , 1_n3960 , 1_n3961 , 1_n3962 , 1_n3963 , 1_n3964 , 1_n3965 , 1_n3966 , 1_n3967 , 1_n3968 , 1_n3969 , 1_n3970 , 1_n3971 , 1_n3972 , 1_n3973 , 1_n3974 , 1_n3975 , 1_n3976 , 1_n3977 , 1_n3978 , 1_n3979 , 1_n3980 , 1_n3981 , 1_n3982 , 1_n3983 , 1_n3984 , 1_n3985 , 1_n3986 , 1_n3987 , 1_n3988 , 1_n3989 , 1_n3990 , 1_n3991 , 1_n3992 , 1_n3993 , 1_n3994 , 1_n3995 , 1_n3996 , 1_n3997 , 1_n3998 , 1_n3999 , 1_n4000 , 1_n4001 , 1_n4002 , 1_n4003 , 1_n4004 , 1_n4005 , 1_n4007 , 1_n4008 , 1_n4009 , 1_n4010 , 1_n4011 , 1_n4012 , 1_n4013 , 1_n4014 , 1_n4015 , 1_n4016 , 1_n4017 , 1_n4018 , 1_n4019 , 1_n4020 , 1_n4021 , 1_n4022 , 1_n4023 , 1_n4024 , 1_n4025 , 1_n4026 , 1_n4027 , 1_n4028 , 1_n4029 , 1_n4030 , 1_n4031 , 1_n4032 , 1_n4033 , 1_n4034 , 1_n4035 , 1_n4036 , 1_n4037 , 1_n4038 , 1_n4039 , 1_n4040 , 1_n4041 , 1_n4042 , 1_n4043 , 1_n4044 , 1_n4045 , 1_n4046 , 1_n4047 , 1_n4048 , 1_n4049 , 1_n4050 , 1_n4051 , 1_n4052 , 1_n4053 , 1_n4054 , 1_n4055 , 1_n4056 , 1_n4057 , 1_n4058 , 1_n4060 , 1_n4061 , 1_n4062 , 1_n4063 , 1_n4064 , 1_n4065 , 1_n4066 , 1_n4067 , 1_n4068 , 1_n4069 , 1_n4070 , 1_n4071 , 1_n4072 , 1_n4073 , 1_n4074 , 1_n4076 , 1_n4077 , 1_n4078 , 1_n4079 , 1_n4080 , 1_n4081 , 1_n4082 , 1_n4083 , 1_n4084 , 1_n4085 , 1_n4086 , 1_n4087 , 1_n4088 , 1_n4089 , 1_n4090 , 1_n4091 , 1_n4092 , 1_n4093 , 1_n4094 , 1_n4095 , 1_n4096 , 1_n4097 , 1_n4098 , 1_n4099 , 1_n4100 , 1_n4101 , 1_n4102 , 1_n4103 , 1_n4104 , 1_n4105 , 1_n4106 , 1_n4107 , 1_n4108 , 1_n4109 , 1_n4110 , 1_n4111 , 1_n4112 , 1_n4113 , 1_n4115 , 1_n4116 , 1_n4117 , 1_n4118 , 1_n4119 , 1_n4120 , 1_n4121 , 1_n4123 , 1_n4124 , 1_n4125 , 1_n4126 , 1_n4127 , 1_n4128 , 1_n4129 , 1_n4130 , 1_n4131 , 1_n4132 , 1_n4133 , 1_n4134 , 1_n4135 , 1_n4136 , 1_n4137 , 1_n4138 , 1_n4139 , 1_n4140 , 1_n4142 , 1_n4143 , 1_n4144 , 1_n4145 , 1_n4146 , 1_n4147 , 1_n4148 , 1_n4149 , 1_n4150 , 1_n4151 , 1_n4152 , 1_n4153 , 1_n4154 , 1_n4155 , 1_n4156 , 1_n4157 , 1_n4158 , 1_n4159 , 1_n4160 , 1_n4161 , 1_n4162 , 1_n4163 , 1_n4164 , 1_n4165 , 1_n4166 , 1_n4167 , 1_n4168 , 1_n4169 , 1_n4170 , 1_n4171 , 1_n4172 , 1_n4173 , 1_n4174 , 1_n4175 , 1_n4176 , 1_n4177 , 1_n4178 , 1_n4179 , 1_n4180 , 1_n4181 , 1_n4182 , 1_n4183 , 1_n4184 , 1_n4185 , 1_n4186 , 1_n4187 , 1_n4188 , 1_n4189 , 1_n4190 , 1_n4191 , 1_n4192 , 1_n4193 , 1_n4194 , 1_n4195 , 1_n4196 , 1_n4197 , 1_n4198 , 1_n4199 , 1_n4200 , 1_n4201 , 1_n4203 , 1_n4204 , 1_n4205 , 1_n4206 , 1_n4207 , 1_n4208 , 1_n4209 , 1_n4210 , 1_n4211 , 1_n4212 , 1_n4213 , 1_n4214 , 1_n4215 , 1_n4216 , 1_n4217 , 1_n4218 , 1_n4219 , 1_n4220 , 1_n4221 , 1_n4222 , 1_n4223 , 1_n4224 , 1_n4225 , 1_n4226 , 1_n4227 , 1_n4228 , 1_n4229 , 1_n4230 , 1_n4231 , 1_n4232 , 1_n4233 , 1_n4234 , 1_n4235 , 1_n4236 , 1_n4237 , 1_n4238 , 1_n4239 , 1_n4240 , 1_n4241 , 1_n4242 , 1_n4243 , 1_n4244 , 1_n4245 , 1_n4246 , 1_n4247 , 1_n4248 , 1_n4249 , 1_n4250 , 1_n4251 , 1_n4252 , 1_n4253 , 1_n4254 , 1_n4255 , 1_n4256 , 1_n4257 , 1_n4258 , 1_n4259 , 1_n4260 , 1_n4261 , 1_n4262 , 1_n4263 , 1_n4264 , 1_n4265 , 1_n4266 , 1_n4267 , 1_n4268 , 1_n4269 , 1_n4270 , 1_n4271 , 1_n4272 , 1_n4273 , 1_n4274 , 1_n4275 , 1_n4276 , 1_n4277 , 1_n4278 , 1_n4279 , 1_n4280 , 1_n4281 , 1_n4282 , 1_n4283 , 1_n4284 , 1_n4285 , 1_n4286 , 1_n4287 , 1_n4288 , 1_n4289 , 1_n4290 , 1_n4291 , 1_n4292 , 1_n4293 , 1_n4294 , 1_n4295 , 1_n4296 , 1_n4297 , 1_n4298 , 1_n4299 , 1_n4300 , 1_n4301 , 1_n4302 , 1_n4303 , 1_n4304 , 1_n4305 , 1_n4306 , 1_n4307 , 1_n4308 , 1_n4309 , 1_n4310 , 1_n4311 , 1_n4312 , 1_n4313 , 1_n4314 , 1_n4315 , 1_n4316 , 1_n4317 , 1_n4318 , 1_n4319 , 1_n4320 , 1_n4321 , 1_n4322 , 1_n4323 , 1_n4324 , 1_n4325 , 1_n4326 , 1_n4327 , 1_n4328 , 1_n4329 , 1_n4331 , 1_n4332 , 1_n4333 , 1_n4334 , 1_n4336 , 1_n4337 , 1_n4338 , 1_n4339 , 1_n4340 , 1_n4341 , 1_n4342 , 1_n4343 , 1_n4344 , 1_n4345 , 1_n4346 , 1_n4347 , 1_n4348 , 1_n4349 , 1_n4350 , 1_n4351 , 1_n4352 , 1_n4353 , 1_n4354 , 1_n4355 , 1_n4356 , 1_n4358 , 1_n4359 , 1_n4360 , 1_n4361 , 1_n4362 , 1_n4363 , 1_n4364 , 1_n4365 , 1_n4366 , 1_n4367 , 1_n4368 , 1_n4369 , 1_n4370 , 1_n4371 , 1_n4372 , 1_n4373 , 1_n4374 , 1_n4375 , 1_n4376 , 1_n4377 , 1_n4378 , 1_n4379 , 1_n4380 , 1_n4381 , 1_n4383 , 1_n4384 , 1_n4385 , 1_n4386 , 1_n4387 , 1_n4388 , 1_n4389 , 1_n4390 , 1_n4391 , 1_n4392 , 1_n4393 , 1_n4394 , 1_n4395 , 1_n4396 , 1_n4397 , 1_n4398 , 1_n4399 , 1_n4400 , 1_n4401 , 1_n4402 , 1_n4403 , 1_n4404 , 1_n4405 , 1_n4406 , 1_n4407 , 1_n4408 , 1_n4409 , 1_n4410 , 1_n4411 , 1_n4412 , 1_n4413 , 1_n4414 , 1_n4415 , 1_n4416 , 1_n4417 , 1_n4418 , 1_n4420 , 1_n4421 , 1_n4422 , 1_n4423 , 1_n4424 , 1_n4425 , 1_n4426 , 1_n4427 , 1_n4428 , 1_n4429 , 1_n4430 , 1_n4431 , 1_n4432 , 1_n4433 , 1_n4434 , 1_n4435 , 1_n4436 , 1_n4437 , 1_n4438 , 1_n4439 , 1_n4440 , 1_n4441 , 1_n4442 , 1_n4443 , 1_n4444 , 1_n4445 , 1_n4446 , 1_n4447 , 1_n4448 , 1_n4449 , 1_n4450 , 1_n4451 , 1_n4453 , 1_n4454 , 1_n4455 , 1_n4456 , 1_n4457 , 1_n4458 , 1_n4459 , 1_n4460 , 1_n4461 , 1_n4462 , 1_n4463 , 1_n4464 , 1_n4465 , 1_n4466 , 1_n4467 , 1_n4468 , 1_n4469 , 1_n4471 , 1_n4472 , 1_n4473 , 1_n4474 , 1_n4475 , 1_n4476 , 1_n4477 , 1_n4478 , 1_n4479 , 1_n4480 , 1_n4481 , 1_n4482 , 1_n4483 , 1_n4484 , 1_n4485 , 1_n4486 , 1_n4487 , 1_n4488 , 1_n4489 , 1_n4490 , 1_n4491 , 1_n4492 , 1_n4493 , 1_n4494 , 1_n4495 , 1_n4496 , 1_n4497 , 1_n4498 , 1_n4499 , 1_n4500 , 1_n4501 , 1_n4502 , 1_n4503 , 1_n4504 , 1_n4505 , 1_n4506 , 1_n4507 , 1_n4508 , 1_n4509 , 1_n4510 , 1_n4511 , 1_n4512 , 1_n4513 , 1_n4514 , 1_n4515 , 1_n4516 , 1_n4517 , 1_n4518 , 1_n4519 , 1_n4520 , 1_n4521 , 1_n4522 , 1_n4523 , 1_n4524 , 1_n4525 , 1_n4526 , 1_n4527 , 1_n4528 , 1_n4529 , 1_n4530 , 1_n4531 , 1_n4532 , 1_n4533 , 1_n4534 , 1_n4535 , 1_n4536 , 1_n4537 , 1_n4538 , 1_n4539 , 1_n4540 , 1_n4541 , 1_n4542 , 1_n4543 , 1_n4544 , 1_n4545 , 1_n4546 , 1_n4547 , 1_n4548 , 1_n4549 , 1_n4550 , 1_n4551 , 1_n4552 , 1_n4554 , 1_n4555 , 1_n4556 , 1_n4557 , 1_n4558 , 1_n4559 , 1_n4560 , 1_n4561 , 1_n4562 , 1_n4563 , 1_n4564 , 1_n4565 , 1_n4566 , 1_n4567 , 1_n4568 , 1_n4569 , 1_n4570 , 1_n4571 , 1_n4572 , 1_n4573 , 1_n4574 , 1_n4575 , 1_n4576 , 1_n4577 , 1_n4578 , 1_n4579 , 1_n4580 , 1_n4581 , 1_n4582 , 1_n4583 , 1_n4584 , 1_n4585 , 1_n4586 , 1_n4587 , 1_n4588 , 1_n4589 , 1_n4590 , 1_n4591 , 1_n4592 , 1_n4593 , 1_n4594 , 1_n4595 , 1_n4596 , 1_n4597 , 1_n4598 , 1_n4599 , 1_n4600 , 1_n4601 , 1_n4602 , 1_n4603 , 1_n4604 , 1_n4605 , 1_n4606 , 1_n4607 , 1_n4608 , 1_n4609 , 1_n4610 , 1_n4611 , 1_n4612 , 1_n4613 , 1_n4614 , 1_n4615 , 1_n4616 , 1_n4617 , 1_n4618 , 1_n4619 , 1_n4620 , 1_n4621 , 1_n4622 , 1_n4623 , 1_n4624 , 1_n4625 , 1_n4626 , 1_n4627 , 1_n4628 , 1_n4629 , 1_n4630 , 1_n4631 , 1_n4632 , 1_n4633 , 1_n4634 , 1_n4635 , 1_n4636 , 1_n4637 , 1_n4638 , 1_n4639 , 1_n4640 , 1_n4641 , 1_n4642 , 1_n4643 , 1_n4644 , 1_n4645 , 1_n4646 , 1_n4647 , 1_n4648 , 1_n4649 , 1_n4650 , 1_n4651 , 1_n4652 , 1_n4653 , 1_n4654 , 1_n4655 , 1_n4656 , 1_n4657 , 1_n4658 , 1_n4659 , 1_n4660 , 1_n4661 , 1_n4662 , 1_n4663 , 1_n4664 , 1_n4665 , 1_n4666 , 1_n4667 , 1_n4668 , 1_n4669 , 1_n4670 , 1_n4671 , 1_n4672 , 1_n4673 , 1_n4674 , 1_n4675 , 1_n4676 , 1_n4677 , 1_n4678 , 1_n4679 , 1_n4680 , 1_n4681 , 1_n4682 , 1_n4683 , 1_n4684 , 1_n4685 , 1_n4686 , 1_n4687 , 1_n4688 , 1_n4689 , 1_n4690 , 1_n4691 , 1_n4692 , 1_n4693 , 1_n4694 , 1_n4695 , 1_n4696 , 1_n4697 , 1_n4698 , 1_n4699 , 1_n4700 , 1_n4701 , 1_n4702 , 1_n4703 , 1_n4704 , 1_n4705 , 1_n4706 , 1_n4707 , 1_n4708 , 1_n4709 , 1_n4710 , 1_n4711 , 1_n4712 , 1_n4713 , 1_n4714 , 1_n4715 , 1_n4716 , 1_n4717 , 1_n4718 , 1_n4719 , 1_n4720 , 1_n4721 , 1_n4722 , 1_n4723 , 1_n4724 , 1_n4725 , 1_n4726 , 1_n4727 , 1_n4728 , 1_n4729 , 1_n4730 , 1_n4731 , 1_n4732 , 1_n4733 , 1_n4734 , 1_n4735 , 1_n4736 , 1_n4737 , 1_n4738 , 1_n4739 , 1_n4740 , 1_n4741 , 1_n4742 , 1_n4744 , 1_n4745 , 1_n4746 , 1_n4747 , 1_n4749 , 1_n4750 , 1_n4751 , 1_n4752 , 1_n4753 , 1_n4754 , 1_n4755 , 1_n4756 , 1_n4757 , 1_n4758 , 1_n4759 , 1_n4760 , 1_n4761 , 1_n4762 , 1_n4763 , 1_n4764 , 1_n4765 , 1_n4766 , 1_n4767 , 1_n4768 , 1_n4769 , 1_n4770 , 1_n4771 , 1_n4772 , 1_n4773 , 1_n4774 , 1_n4775 , 1_n4776 , 1_n4778 , 1_n4779 , 1_n4780 , 1_n4781 , 1_n4782 , 1_n4783 , 1_n4784 , 1_n4785 , 1_n4786 , 1_n4787 , 1_n4788 , 1_n4789 , 1_n4790 , 1_n4791 , 1_n4792 , 1_n4793 , 1_n4794 , 1_n4795 , 1_n4796 , 1_n4797 , 1_n4798 , 1_n4799 , 1_n4800 , 1_n4801 , 1_n4802 , 1_n4803 , 1_n4804 , 1_n4805 , 1_n4806 , 1_n4807 , 1_n4808 , 1_n4809 , 1_n4810 , 1_n4811 , 1_n4812 , 1_n4813 , 1_n4814 , 1_n4815 , 1_n4816 , 1_n4817 , 1_n4818 , 1_n4819 , 1_n4820 , 1_n4821 , 1_n4822 , 1_n4823 , 1_n4825 , 1_n4826 , 1_n4827 , 1_n4828 , 1_n4829 , 1_n4830 , 1_n4831 , 1_n4832 , 1_n4833 , 1_n4834 , 1_n4835 , 1_n4836 , 1_n4837 , 1_n4838 , 1_n4839 , 1_n4840 , 1_n4841 , 1_n4842 , 1_n4843 , 1_n4844 , 1_n4845 , 1_n4846 , 1_n4847 , 1_n4848 , 1_n4849 , 1_n4850 , 1_n4851 , 1_n4852 , 1_n4853 , 1_n4854 , 1_n4855 , 1_n4856 , 1_n4857 , 1_n4858 , 1_n4859 , 1_n4860 , 1_n4861 , 1_n4863 , 1_n4865 , 1_n4866 , 1_n4867 , 1_n4868 , 1_n4869 , 1_n4870 , 1_n4871 , 1_n4872 , 1_n4873 , 1_n4874 , 1_n4875 , 1_n4876 , 1_n4877 , 1_n4878 , 1_n4879 , 1_n4880 , 1_n4881 , 1_n4882 , 1_n4883 , 1_n4884 , 1_n4885 , 1_n4886 , 1_n4887 , 1_n4888 , 1_n4889 , 1_n4890 , 1_n4891 , 1_n4892 , 1_n4893 , 1_n4894 , 1_n4895 , 1_n4896 , 1_n4897 , 1_n4898 , 1_n4899 , 1_n4900 , 1_n4901 , 1_n4902 , 1_n4903 , 1_n4904 , 1_n4905 , 1_n4906 , 1_n4907 , 1_n4908 , 1_n4909 , 1_n4910 , 1_n4911 , 1_n4912 , 1_n4913 , 1_n4914 , 1_n4915 , 1_n4916 , 1_n4917 , 1_n4918 , 1_n4919 , 1_n4920 , 1_n4921 , 1_n4922 , 1_n4923 , 1_n4924 , 1_n4925 , 1_n4926 , 1_n4927 , 1_n4928 , 1_n4929 , 1_n4930 , 1_n4931 , 1_n4932 , 1_n4933 , 1_n4934 , 1_n4935 , 1_n4936 , 1_n4937 , 1_n4938 , 1_n4939 , 1_n4940 , 1_n4941 , 1_n4942 , 1_n4943 , 1_n4944 , 1_n4945 , 1_n4946 , 1_n4947 , 1_n4948 , 1_n4949 , 1_n4950 , 1_n4951 , 1_n4952 , 1_n4953 , 1_n4954 , 1_n4955 , 1_n4956 , 1_n4957 , 1_n4958 , 1_n4959 , 1_n4960 , 1_n4961 , 1_n4962 , 1_n4963 , 1_n4965 , 1_n4966 , 1_n4967 , 1_n4968 , 1_n4969 , 1_n4970 , 1_n4971 , 1_n4972 , 1_n4973 , 1_n4974 , 1_n4975 , 1_n4976 , 1_n4977 , 1_n4978 , 1_n4979 , 1_n4980 , 1_n4981 , 1_n4982 , 1_n4983 , 1_n4984 , 1_n4985 , 1_n4986 , 1_n4987 , 1_n4988 , 1_n4989 , 1_n4990 , 1_n4991 , 1_n4992 , 1_n4993 , 1_n4994 , 1_n4995 , 1_n4996 , 1_n4997 , 1_n4999 , 1_n5000 , 1_n5001 , 1_n5002 , 1_n5004 , 1_n5005 , 1_n5006 , 1_n5007 , 1_n5008 , 1_n5009 , 1_n5010 , 1_n5011 , 1_n5012 , 1_n5013 , 1_n5014 , 1_n5015 , 1_n5016 , 1_n5017 , 1_n5018 , 1_n5019 , 1_n5020 , 1_n5021 , 1_n5022 , 1_n5023 , 1_n5024 , 1_n5025 , 1_n5026 , 1_n5027 , 1_n5028 , 1_n5029 , 1_n5030 , 1_n5032 , 1_n5033 , 1_n5034 , 1_n5035 , 1_n5036 , 1_n5037 , 1_n5038 , 1_n5039 , 1_n5040 , 1_n5041 , 1_n5042 , 1_n5043 , 1_n5044 , 1_n5045 , 1_n5046 , 1_n5047 , 1_n5048 , 1_n5049 , 1_n5050 , 1_n5051 , 1_n5052 , 1_n5053 , 1_n5054 , 1_n5055 , 1_n5056 , 1_n5057 , 1_n5058 , 1_n5059 , 1_n5061 , 1_n5062 , 1_n5063 , 1_n5064 , 1_n5066 , 1_n5067 , 1_n5068 , 1_n5069 , 1_n5070 , 1_n5071 , 1_n5072 , 1_n5073 , 1_n5074 , 1_n5075 , 1_n5076 , 1_n5077 , 1_n5078 , 1_n5079 , 1_n5080 , 1_n5081 , 1_n5082 , 1_n5083 , 1_n5084 , 1_n5085 , 1_n5086 , 1_n5087 , 1_n5088 , 1_n5089 , 1_n5090 , 1_n5091 , 1_n5092 , 1_n5093 , 1_n5094 , 1_n5095 , 1_n5096 , 1_n5097 , 1_n5098 , 1_n5099 , 1_n5100 , 1_n5101 , 1_n5102 , 1_n5103 , 1_n5104 , 1_n5105 , 1_n5106 , 1_n5107 , 1_n5108 , 1_n5109 , 1_n5110 , 1_n5111 , 1_n5112 , 1_n5113 , 1_n5114 , 1_n5115 , 1_n5116 , 1_n5117 , 1_n5118 , 1_n5119 , 1_n5120 , 1_n5121 , 1_n5122 , 1_n5123 , 1_n5124 , 1_n5125 , 1_n5126 , 1_n5127 , 1_n5128 , 1_n5129 , 1_n5130 , 1_n5131 , 1_n5132 , 1_n5133 , 1_n5134 , 1_n5135 , 1_n5136 , 1_n5137 , 1_n5138 , 1_n5139 , 1_n5140 , 1_n5141 , 1_n5142 , 1_n5143 , 1_n5144 , 1_n5145 , 1_n5146 , 1_n5147 , 1_n5148 , 1_n5149 , 1_n5150 , 1_n5151 , 1_n5152 , 1_n5153 , 1_n5154 , 1_n5155 , 1_n5156 , 1_n5157 , 1_n5158 , 1_n5159 , 1_n5160 , 1_n5161 , 1_n5162 , 1_n5163 , 1_n5164 , 1_n5165 , 1_n5166 , 1_n5168 , 1_n5169 , 1_n5170 , 1_n5171 , 1_n5172 , 1_n5173 , 1_n5174 , 1_n5175 , 1_n5176 , 1_n5177 , 1_n5178 , 1_n5179 , 1_n5180 , 1_n5181 , 1_n5182 , 1_n5183 , 1_n5184 , 1_n5185 , 1_n5186 , 1_n5187 , 1_n5188 , 1_n5190 , 1_n5191 , 1_n5192 , 1_n5193 , 1_n5194 , 1_n5195 , 1_n5196 , 1_n5197 , 1_n5198 , 1_n5199 , 1_n5200 , 1_n5201 , 1_n5202 , 1_n5203 , 1_n5204 , 1_n5205 , 1_n5206 , 1_n5207 , 1_n5208 , 1_n5209 , 1_n5210 , 1_n5211 , 1_n5212 , 1_n5213 , 1_n5215 , 1_n5216 , 1_n5217 , 1_n5218 , 1_n5219 , 1_n5220 , 1_n5221 , 1_n5222 , 1_n5223 , 1_n5224 , 1_n5225 , 1_n5226 , 1_n5227 , 1_n5228 , 1_n5229 , 1_n5230 , 1_n5231 , 1_n5232 , 1_n5233 , 1_n5234 , 1_n5235 , 1_n5236 , 1_n5237 , 1_n5238 , 1_n5239 , 1_n5240 , 1_n5241 , 1_n5242 , 1_n5243 , 1_n5244 , 1_n5245 , 1_n5246 , 1_n5247 , 1_n5248 , 1_n5249 , 1_n5250 , 1_n5251 , 1_n5252 , 1_n5253 , 1_n5254 , 1_n5255 , 1_n5256 , 1_n5257 , 1_n5258 , 1_n5259 , 1_n5260 , 1_n5261 , 1_n5262 , 1_n5263 , 1_n5264 , 1_n5265 , 1_n5266 , 1_n5267 , 1_n5268 , 1_n5269 , 1_n5270 , 1_n5271 , 1_n5272 , 1_n5273 , 1_n5274 , 1_n5275 , 1_n5276 , 1_n5277 , 1_n5278 , 1_n5279 , 1_n5280 , 1_n5281 , 1_n5282 , 1_n5283 , 1_n5284 , 1_n5285 , 1_n5286 , 1_n5287 , 1_n5288 , 1_n5289 , 1_n5290 , 1_n5291 , 1_n5292 , 1_n5293 , 1_n5294 , 1_n5295 , 1_n5296 , 1_n5297 , 1_n5298 , 1_n5299 , 1_n5300 , 1_n5301 , 1_n5302 , 1_n5303 , 1_n5304 , 1_n5305 , 1_n5306 , 1_n5307 , 1_n5308 , 1_n5309 , 1_n5310 , 1_n5311 , 1_n5312 , 1_n5313 , 1_n5314 , 1_n5315 , 1_n5316 , 1_n5317 , 1_n5318 , 1_n5319 , 1_n5321 , 1_n5322 , 1_n5323 , 1_n5324 , 1_n5325 , 1_n5326 , 1_n5327 , 1_n5328 , 1_n5329 , 1_n5330 , 1_n5331 , 1_n5332 , 1_n5333 , 1_n5334 , 1_n5335 , 1_n5336 , 1_n5337 , 1_n5338 , 1_n5339 , 1_n5340 , 1_n5341 , 1_n5342 , 1_n5343 , 1_n5344 , 1_n5345 , 1_n5346 , 1_n5347 , 1_n5348 , 1_n5349 , 1_n5350 , 1_n5351 , 1_n5352 , 1_n5353 , 1_n5354 , 1_n5355 , 1_n5357 , 1_n5358 , 1_n5359 , 1_n5360 , 1_n5361 , 1_n5362 , 1_n5363 , 1_n5365 , 1_n5366 , 1_n5367 , 1_n5368 , 1_n5369 , 1_n5370 , 1_n5371 , 1_n5372 , 1_n5373 , 1_n5374 , 1_n5375 , 1_n5376 , 1_n5377 , 1_n5378 , 1_n5379 , 1_n5380 , 1_n5381 , 1_n5382 , 1_n5383 , 1_n5384 , 1_n5385 , 1_n5386 , 1_n5387 , 1_n5388 , 1_n5389 , 1_n5390 , 1_n5391 , 1_n5392 , 1_n5393 , 1_n5394 , 1_n5395 , 1_n5396 , 1_n5397 , 1_n5398 , 1_n5399 , 1_n5400 , 1_n5401 , 1_n5402 , 1_n5403 , 1_n5404 , 1_n5405 , 1_n5406 , 1_n5407 , 1_n5408 , 1_n5409 , 1_n5410 , 1_n5411 , 1_n5412 , 1_n5413 , 1_n5414 , 1_n5415 , 1_n5416 , 1_n5417 , 1_n5418 , 1_n5419 , 1_n5420 , 1_n5421 , 1_n5422 , 1_n5423 , 1_n5424 , 1_n5425 , 1_n5426 , 1_n5428 , 1_n5429 , 1_n5430 , 1_n5431 , 1_n5432 , 1_n5433 , 1_n5434 , 1_n5435 , 1_n5436 , 1_n5437 , 1_n5438 , 1_n5439 , 1_n5440 , 1_n5441 , 1_n5442 , 1_n5443 , 1_n5444 , 1_n5445 , 1_n5446 , 1_n5447 , 1_n5448 , 1_n5449 , 1_n5450 , 1_n5451 , 1_n5452 , 1_n5453 , 1_n5454 , 1_n5455 , 1_n5456 , 1_n5457 , 1_n5458 , 1_n5459 , 1_n5460 , 1_n5461 , 1_n5462 , 1_n5463 , 1_n5464 , 1_n5465 , 1_n5466 , 1_n5467 , 1_n5468 , 1_n5469 , 1_n5471 , 1_n5472 , 1_n5473 , 1_n5474 , 1_n5475 , 1_n5476 , 1_n5477 , 1_n5478 , 1_n5479 , 1_n5480 , 1_n5481 , 1_n5482 , 1_n5483 , 1_n5484 , 1_n5485 , 1_n5486 , 1_n5487 , 1_n5488 , 1_n5489 , 1_n5490 , 1_n5491 , 1_n5492 , 1_n5493 , 1_n5494 , 1_n5495 , 1_n5496 , 1_n5497 , 1_n5498 , 1_n5499 , 1_n5500 , 1_n5501 , 1_n5502 , 1_n5503 , 1_n5504 , 1_n5505 , 1_n5506 , 1_n5507 , 1_n5508 , 1_n5509 , 1_n5510 , 1_n5511 , 1_n5512 , 1_n5513 , 1_n5514 , 1_n5515 , 1_n5516 , 1_n5517 , 1_n5518 , 1_n5519 , 1_n5520 , 1_n5521 , 1_n5522 , 1_n5523 , 1_n5524 , 1_n5525 , 1_n5526 , 1_n5527 , 1_n5528 , 1_n5529 , 1_n5530 , 1_n5531 , 1_n5532 , 1_n5533 , 1_n5534 , 1_n5535 , 1_n5537 , 1_n5538 , 1_n5539 , 1_n5540 , 1_n5541 , 1_n5542 , 1_n5543 , 1_n5544 , 1_n5545 , 1_n5546 , 1_n5547 , 1_n5550 , 1_n5551 , 1_n5552 , 1_n5553 , 1_n5554 , 1_n5555 , 1_n5556 , 1_n5558 , 1_n5559 , 1_n5560 , 1_n5561 , 1_n5562 , 1_n5563 , 1_n5564 , 1_n5565 , 1_n5566 , 1_n5567 , 1_n5569 , 1_n5570 , 1_n5571 , 1_n5572 , 1_n5573 , 1_n5574 , 1_n5575 , 1_n5576 , 1_n5577 , 1_n5578 , 1_n5579 , 1_n5580 , 1_n5581 , 1_n5582 , 1_n5583 , 1_n5584 , 1_n5585 , 1_n5587 , 1_n5588 , 1_n5589 , 1_n5590 , 1_n5591 , 1_n5592 , 1_n5593 , 1_n5594 , 1_n5595 , 1_n5596 , 1_n5597 , 1_n5598 , 1_n5599 , 1_n5600 , 1_n5601 , 1_n5602 , 1_n5603 , 1_n5604 , 1_n5605 , 1_n5606 , 1_n5607 , 1_n5608 , 1_n5610 , 1_n5611 , 1_n5612 , 1_n5613 , 1_n5614 , 1_n5615 , 1_n5616 , 1_n5617 , 1_n5618 , 1_n5619 , 1_n5620 , 1_n5621 , 1_n5622 , 1_n5623 , 1_n5624 , 1_n5625 , 1_n5626 , 1_n5627 , 1_n5628 , 1_n5629 , 1_n5630 , 1_n5631 , 1_n5632 , 1_n5633 , 1_n5634 , 1_n5635 , 1_n5636 , 1_n5637 , 1_n5638 , 1_n5639 , 1_n5640 , 1_n5641 , 1_n5642 , 1_n5643 , 1_n5644 , 1_n5645 , 1_n5646 , 1_n5647 , 1_n5648 , 1_n5649 , 1_n5650 , 1_n5651 , 1_n5652 , 1_n5653 , 1_n5654 , 1_n5655 , 1_n5656 , 1_n5657 , 1_n5658 , 1_n5659 , 1_n5660 , 1_n5661 , 1_n5662 , 1_n5663 , 1_n5664 , 1_n5665 , 1_n5666 , 1_n5667 , 1_n5668 , 1_n5669 , 1_n5670 , 1_n5672 , 1_n5673 , 1_n5674 , 1_n5675 , 1_n5676 , 1_n5677 , 1_n5678 , 1_n5679 , 1_n5680 , 1_n5681 , 1_n5682 , 1_n5683 , 1_n5685 , 1_n5686 , 1_n5687 , 1_n5688 , 1_n5689 , 1_n5690 , 1_n5691 , 1_n5692 , 1_n5693 , 1_n5694 , 1_n5695 , 1_n5696 , 1_n5697 , 1_n5698 , 1_n5699 , 1_n5700 , 1_n5701 , 1_n5702 , 1_n5703 , 1_n5704 , 1_n5705 , 1_n5706 , 1_n5707 , 1_n5708 , 1_n5709 , 1_n5710 , 1_n5711 , 1_n5712 , 1_n5713 , 1_n5714 , 1_n5716 , 1_n5717 , 1_n5718 , 1_n5719 , 1_n5720 , 1_n5721 , 1_n5722 , 1_n5723 , 1_n5724 , 1_n5725 , 1_n5726 , 1_n5727 , 1_n5728 , 1_n5730 , 1_n5731 , 1_n5732 , 1_n5733 , 1_n5734 , 1_n5735 , 1_n5736 , 1_n5737 , 1_n5738 , 1_n5739 , 1_n5740 , 1_n5741 , 1_n5742 , 1_n5743 , 1_n5744 , 1_n5745 , 1_n5746 , 1_n5747 , 1_n5748 , 1_n5749 , 1_n5750 , 1_n5751 , 1_n5752 , 1_n5753 , 1_n5754 , 1_n5755 , 1_n5756 , 1_n5757 , 1_n5759 , 1_n5760 , 1_n5761 , 1_n5762 , 1_n5763 , 1_n5764 , 1_n5765 , 1_n5766 , 1_n5767 , 1_n5768 , 1_n5769 , 1_n5770 , 1_n5771 , 1_n5772 , 1_n5773 , 1_n5774 , 1_n5775 , 1_n5776 , 1_n5777 , 1_n5778 , 1_n5779 , 1_n5780 , 1_n5781 , 1_n5782 , 1_n5783 , 1_n5784 , 1_n5785 , 1_n5786 , 1_n5787 , 1_n5788 , 1_n5789 , 1_n5790 , 1_n5791 , 1_n5792 , 1_n5793 , 1_n5794 , 1_n5795 , 1_n5796 , 1_n5797 , 1_n5798 , 1_n5799 , 1_n5800 , 1_n5802 , 1_n5803 , 1_n5804 , 1_n5805 , 1_n5806 , 1_n5807 , 1_n5808 , 1_n5809 , 1_n5810 , 1_n5811 , 1_n5812 , 1_n5813 , 1_n5814 , 1_n5815 , 1_n5816 , 1_n5817 , 1_n5818 , 1_n5819 , 1_n5820 , 1_n5821 , 1_n5822 , 1_n5823 , 1_n5824 , 1_n5825 , 1_n5826 , 1_n5827 , 1_n5828 , 1_n5829 , 1_n5830 , 1_n5831 , 1_n5832 , 1_n5833 , 1_n5834 , 1_n5835 , 1_n5836 , 1_n5837 , 1_n5838 , 1_n5839 , 1_n5840 , 1_n5841 , 1_n5842 , 1_n5843 , 1_n5844 , 1_n5845 , 1_n5846 , 1_n5847 , 1_n5848 , 1_n5849 , 1_n5850 , 1_n5851 , 1_n5852 , 1_n5853 , 1_n5854 , 1_n5855 , 1_n5856 , 1_n5857 , 1_n5858 , 1_n5859 , 1_n5860 , 1_n5861 , 1_n5862 , 1_n5863 , 1_n5864 , 1_n5865 , 1_n5866 , 1_n5867 , 1_n5868 , 1_n5869 , 1_n5870 , 1_n5871 , 1_n5872 , 1_n5873 , 1_n5874 , 1_n5875 , 1_n5876 , 1_n5877 , 1_n5878 , 1_n5879 , 1_n5880 , 1_n5881 , 1_n5883 , 1_n5885 , 1_n5886 , 1_n5887 , 1_n5888 , 1_n5889 , 1_n5890 , 1_n5891 , 1_n5892 , 1_n5893 , 1_n5894 , 1_n5895 , 1_n5896 , 1_n5897 , 1_n5898 , 1_n5899 , 1_n5900 , 1_n5901 , 1_n5902 , 1_n5903 , 1_n5904 , 1_n5905 , 1_n5906 , 1_n5907 , 1_n5908 , 1_n5909 , 1_n5910 , 1_n5911 , 1_n5912 , 1_n5913 , 1_n5914 , 1_n5915 , 1_n5916 , 1_n5917 , 1_n5918 , 1_n5919 , 1_n5921 , 1_n5922 , 1_n5923 , 1_n5924 , 1_n5925 , 1_n5926 , 1_n5927 , 1_n5928 , 1_n5929 , 1_n5930 , 1_n5931 , 1_n5932 , 1_n5933 , 1_n5934 , 1_n5935 , 1_n5936 , 1_n5937 , 1_n5938 , 1_n5939 , 1_n5940 , 1_n5941 , 1_n5942 , 1_n5943 , 1_n5944 , 1_n5945 , 1_n5946 , 1_n5947 , 1_n5948 , 1_n5949 , 1_n5950 , 1_n5951 , 1_n5952 , 1_n5953 , 1_n5954 , 1_n5955 , 1_n5956 , 1_n5957 , 1_n5958 , 1_n5959 , 1_n5960 , 1_n5961 , 1_n5963 , 1_n5964 , 1_n5965 , 1_n5966 , 1_n5967 , 1_n5968 , 1_n5970 , 1_n5971 , 1_n5972 , 1_n5973 , 1_n5974 , 1_n5975 , 1_n5976 , 1_n5977 , 1_n5978 , 1_n5979 , 1_n5980 , 1_n5981 , 1_n5982 , 1_n5983 , 1_n5984 , 1_n5985 , 1_n5986 , 1_n5987 , 1_n5988 , 1_n5989 , 1_n5990 , 1_n5991 , 1_n5992 , 1_n5993 , 1_n5994 , 1_n5995 , 1_n5996 , 1_n5997 , 1_n5998 , 1_n5999 , 1_n6000 , 1_n6001 , 1_n6002 , 1_n6003 , 1_n6004 , 1_n6005 , 1_n6006 , 1_n6007 , 1_n6008 , 1_n6009 , 1_n6010 , 1_n6011 , 1_n6012 , 1_n6013 , 1_n6014 , 1_n6015 , 1_n6016 , 1_n6017 , 1_n6018 , 1_n6020 , 1_n6021 , 1_n6022 , 1_n6024 , 1_n6025 , 1_n6026 , 1_n6027 , 1_n6028 , 1_n6029 , 1_n6030 , 1_n6031 , 1_n6032 , 1_n6033 , 1_n6034 , 1_n6035 , 1_n6036 , 1_n6037 , 1_n6038 , 1_n6039 , 1_n6040 , 1_n6041 , 1_n6042 , 1_n6043 , 1_n6044 , 1_n6045 , 1_n6046 , 1_n6047 , 1_n6048 , 1_n6049 , 1_n6050 , 1_n6051 , 1_n6052 , 1_n6053 , 1_n6054 , 1_n6055 , 1_n6056 , 1_n6057 , 1_n6058 , 1_n6059 , 1_n6060 , 1_n6061 , 1_n6062 , 1_n6063 , 1_n6064 , 1_n6065 , 1_n6066 , 1_n6067 , 1_n6068 , 1_n6069 , 1_n6070 , 1_n6071 , 1_n6072 , 1_n6073 , 1_n6074 , 1_n6075 , 1_n6076 , 1_n6077 , 1_n6078 , 1_n6079 , 1_n6080 , 1_n6081 , 1_n6082 , 1_n6083 , 1_n6084 , 1_n6086 , 1_n6087 , 1_n6088 , 1_n6089 , 1_n6090 , 1_n6091 , 1_n6092 , 1_n6093 , 1_n6094 , 1_n6095 , 1_n6096 , 1_n6097 , 1_n6098 , 1_n6099 , 1_n6100 , 1_n6101 , 1_n6102 , 1_n6104 , 1_n6105 , 1_n6106 , 1_n6107 , 1_n6108 , 1_n6110 , 1_n6111 , 1_n6112 , 1_n6113 , 1_n6114 , 1_n6115 , 1_n6116 , 1_n6117 , 1_n6118 , 1_n6119 , 1_n6120 , 1_n6121 , 1_n6122 , 1_n6123 , 1_n6124 , 1_n6125 , 1_n6126 , 1_n6127 , 1_n6128 , 1_n6129 , 1_n6130 , 1_n6131 , 1_n6132 , 1_n6133 , 1_n6134 , 1_n6135 , 1_n6136 , 1_n6137 , 1_n6138 , 1_n6139 , 1_n6140 , 1_n6141 , 1_n6142 , 1_n6143 , 1_n6144 , 1_n6145 , 1_n6146 , 1_n6147 , 1_n6148 , 1_n6150 , 1_n6151 , 1_n6152 , 1_n6153 , 1_n6154 , 1_n6155 , 1_n6156 , 1_n6157 , 1_n6158 , 1_n6159 , 1_n6160 , 1_n6161 , 1_n6162 , 1_n6163 , 1_n6164 , 1_n6165 , 1_n6166 , 1_n6167 , 1_n6169 , 1_n6170 , 1_n6171 , 1_n6172 , 1_n6173 , 1_n6174 , 1_n6175 , 1_n6176 , 1_n6177 , 1_n6178 , 1_n6179 , 1_n6180 , 1_n6181 , 1_n6182 , 1_n6183 , 1_n6184 , 1_n6185 , 1_n6186 , 1_n6187 , 1_n6188 , 1_n6189 , 1_n6190 , 1_n6191 , 1_n6192 , 1_n6193 , 1_n6194 , 1_n6195 , 1_n6196 , 1_n6197 , 1_n6198 , 1_n6199 , 1_n6200 , 1_n6201 , 1_n6202 , 1_n6203 , 1_n6204 , 1_n6205 , 1_n6206 , 1_n6207 , 1_n6208 , 1_n6209 , 1_n6210 , 1_n6211 , 1_n6212 , 1_n6213 , 1_n6214 , 1_n6215 , 1_n6216 , 1_n6217 , 1_n6218 , 1_n6219 , 1_n6220 , 1_n6221 , 1_n6222 , 1_n6223 , 1_n6224 , 1_n6225 , 1_n6226 , 1_n6227 , 1_n6228 , 1_n6229 , 1_n6230 , 1_n6231 , 1_n6232 , 1_n6233 , 1_n6234 , 1_n6235 , 1_n6236 , 1_n6237 , 1_n6238 , 1_n6239 , 1_n6240 , 1_n6241 , 1_n6242 , 1_n6243 , 1_n6244 , 1_n6245 , 1_n6246 , 1_n6247 , 1_n6248 , 1_n6249 , 1_n6250 , 1_n6251 , 1_n6252 , 1_n6253 , 1_n6254 , 1_n6255 , 1_n6256 , 1_n6257 , 1_n6258 , 1_n6259 , 1_n6260 , 1_n6261 , 1_n6262 , 1_n6263 , 1_n6264 , 1_n6265 , 1_n6266 , 1_n6267 , 1_n6268 , 1_n6269 , 1_n6270 , 1_n6271 , 1_n6272 , 1_n6273 , 1_n6274 , 1_n6275 , 1_n6276 , 1_n6277 , 1_n6278 , 1_n6279 , 1_n6280 , 1_n6281 , 1_n6282 , 1_n6283 , 1_n6284 , 1_n6285 , 1_n6286 , 1_n6287 , 1_n6288 , 1_n6289 , 1_n6290 , 1_n6291 , 1_n6292 , 1_n6293 , 1_n6294 , 1_n6295 , 1_n6296 , 1_n6298 , 1_n6299 , 1_n6300 , 1_n6302 , 1_n6303 , 1_n6304 , 1_n6305 , 1_n6306 , 1_n6307 , 1_n6308 , 1_n6309 , 1_n6310 , 1_n6311 , 1_n6312 , 1_n6313 , 1_n6314 , 1_n6315 , 1_n6316 , 1_n6317 , 1_n6318 , 1_n6319 , 1_n6320 , 1_n6321 , 1_n6322 , 1_n6323 , 1_n6324 , 1_n6325 , 1_n6326 , 1_n6327 , 1_n6328 , 1_n6329 , 1_n6330 , 1_n6331 , 1_n6332 , 1_n6334 , 1_n6335 , 1_n6336 , 1_n6337 , 1_n6338 , 1_n6339 , 1_n6340 , 1_n6341 , 1_n6342 , 1_n6343 , 1_n6344 , 1_n6345 , 1_n6346 , 1_n6347 , 1_n6348 , 1_n6349 , 1_n6350 , 1_n6351 , 1_n6352 , 1_n6353 , 1_n6354 , 1_n6355 , 1_n6356 , 1_n6357 , 1_n6358 , 1_n6359 , 1_n6360 , 1_n6361 , 1_n6362 , 1_n6363 , 1_n6364 , 1_n6365 , 1_n6366 , 1_n6367 , 1_n6368 , 1_n6369 , 1_n6370 , 1_n6371 , 1_n6372 , 1_n6373 , 1_n6374 , 1_n6375 , 1_n6376 , 1_n6377 , 1_n6378 , 1_n6379 , 1_n6380 , 1_n6381 , 1_n6382 , 1_n6383 , 1_n6384 , 1_n6385 , 1_n6386 , 1_n6387 , 1_n6388 , 1_n6389 , 1_n6390 , 1_n6391 , 1_n6393 , 1_n6394 , 1_n6395 , 1_n6396 , 1_n6397 , 1_n6398 , 1_n6399 , 1_n6400 , 1_n6401 , 1_n6402 , 1_n6403 , 1_n6404 , 1_n6405 , 1_n6406 , 1_n6407 , 1_n6408 , 1_n6410 , 1_n6411 , 1_n6412 , 1_n6413 , 1_n6414 , 1_n6415 , 1_n6416 , 1_n6417 , 1_n6418 , 1_n6419 , 1_n6420 , 1_n6421 , 1_n6422 , 1_n6423 , 1_n6424 , 1_n6425 , 1_n6426 , 1_n6427 , 1_n6428 , 1_n6429 , 1_n6430 , 1_n6431 , 1_n6432 , 1_n6433 , 1_n6435 , 1_n6436 , 1_n6437 , 1_n6438 , 1_n6439 , 1_n6440 , 1_n6441 , 1_n6442 , 1_n6443 , 1_n6444 , 1_n6445 , 1_n6446 , 1_n6447 , 1_n6448 , 1_n6449 , 1_n6450 , 1_n6451 , 1_n6452 , 1_n6453 , 1_n6454 , 1_n6455 , 1_n6456 , 1_n6457 , 1_n6458 , 1_n6459 , 1_n6460 , 1_n6461 , 1_n6462 , 1_n6463 , 1_n6464 , 1_n6465 , 1_n6466 , 1_n6467 , 1_n6468 , 1_n6469 , 1_n6470 , 1_n6471 , 1_n6472 , 1_n6473 , 1_n6474 , 1_n6475 , 1_n6476 , 1_n6477 , 1_n6478 , 1_n6479 , 1_n6480 , 1_n6481 , 1_n6482 , 1_n6483 , 1_n6484 , 1_n6485 , 1_n6486 , 1_n6487 , 1_n6488 , 1_n6489 , 1_n6490 , 1_n6491 , 1_n6492 , 1_n6493 , 1_n6494 , 1_n6495 , 1_n6496 , 1_n6497 , 1_n6498 , 1_n6499 , 1_n6500 , 1_n6501 , 1_n6502 , 1_n6503 , 1_n6504 , 1_n6505 , 1_n6506 , 1_n6507 , 1_n6508 , 1_n6509 , 1_n6510 , 1_n6511 , 1_n6512 , 1_n6513 , 1_n6514 , 1_n6515 , 1_n6516 , 1_n6517 , 1_n6518 , 1_n6519 , 1_n6520 , 1_n6521 , 1_n6522 , 1_n6523 , 1_n6524 , 1_n6525 , 1_n6526 , 1_n6527 , 1_n6528 , 1_n6529 , 1_n6530 , 1_n6531 , 1_n6532 , 1_n6533 , 1_n6534 , 1_n6535 , 1_n6536 , 1_n6537 , 1_n6538 , 1_n6539 , 1_n6540 , 1_n6541 , 1_n6542 , 1_n6543 , 1_n6544 , 1_n6545 , 1_n6546 , 1_n6547 , 1_n6548 , 1_n6549 , 1_n6550 , 1_n6551 , 1_n6552 , 1_n6553 , 1_n6554 , 1_n6555 , 1_n6556 , 1_n6557 , 1_n6558 , 1_n6559 , 1_n6560 , 1_n6561 , 1_n6562 , 1_n6563 , 1_n6564 , 1_n6565 , 1_n6566 , 1_n6567 , 1_n6568 , 1_n6569 , 1_n6570 , 1_n6571 , 1_n6572 , 1_n6573 , 1_n6574 , 1_n6575 , 1_n6576 , 1_n6577 , 1_n6578 , 1_n6579 , 1_n6580 , 1_n6581 , 1_n6582 , 1_n6583 , 1_n6584 , 1_n6585 , 1_n6587 , 1_n6588 , 1_n6589 , 1_n6590 , 1_n6591 , 1_n6592 , 1_n6593 , 1_n6594 , 1_n6595 , 1_n6596 , 1_n6597 , 1_n6598 , 1_n6599 , 1_n6600 , 1_n6601 , 1_n6602 , 1_n6603 , 1_n6604 , 1_n6605 , 1_n6606 , 1_n6607 , 1_n6608 , 1_n6609 , 1_n6610 , 1_n6611 , 1_n6612 , 1_n6613 , 1_n6614 , 1_n6615 , 1_n6616 , 1_n6617 , 1_n6618 , 1_n6619 , 1_n6620 , 1_n6621 , 1_n6622 , 1_n6623 , 1_n6624 , 1_n6625 , 1_n6626 , 1_n6627 , 1_n6628 , 1_n6629 , 1_n6630 , 1_n6631 , 1_n6632 , 1_n6633 , 1_n6634 , 1_n6635 , 1_n6636 , 1_n6637 , 1_n6638 , 1_n6639 , 1_n6640 , 1_n6641 , 1_n6642 , 1_n6643 , 1_n6644 , 1_n6645 , 1_n6646 , 1_n6647 , 1_n6648 , 1_n6649 , 1_n6650 , 1_n6651 , 1_n6652 , 1_n6653 , 1_n6654 , 1_n6656 , 1_n6657 , 1_n6658 , 1_n6659 , 1_n6660 , 1_n6661 , 1_n6662 , 1_n6663 , 1_n6664 , 1_n6665 , 1_n6666 , 1_n6667 , 1_n6669 , 1_n6670 , 1_n6671 , 1_n6672 , 1_n6673 , 1_n6674 , 1_n6675 , 1_n6676 , 1_n6677 , 1_n6678 , 1_n6679 , 1_n6680 , 1_n6681 , 1_n6682 , 1_n6684 , 1_n6685 , 1_n6686 , 1_n6687 , 1_n6688 , 1_n6689 , 1_n6690 , 1_n6691 , 1_n6692 , 1_n6693 , 1_n6694 , 1_n6695 , 1_n6696 , 1_n6697 , 1_n6698 , 1_n6699 , 1_n6700 , 1_n6701 , 1_n6702 , 1_n6703 , 1_n6704 , 1_n6705 , 1_n6706 , 1_n6707 , 1_n6708 , 1_n6709 , 1_n6710 , 1_n6711 , 1_n6712 , 1_n6713 , 1_n6714 , 1_n6715 , 1_n6716 , 1_n6717 , 1_n6718 , 1_n6719 , 1_n6720 , 1_n6721 , 1_n6722 , 1_n6723 , 1_n6724 , 1_n6725 , 1_n6726 , 1_n6727 , 1_n6728 , 1_n6729 , 1_n6730 , 1_n6731 , 1_n6732 , 1_n6733 , 1_n6734 , 1_n6735 , 1_n6736 , 1_n6737 , 1_n6738 , 1_n6739 , 1_n6740 , 1_n6741 , 1_n6742 , 1_n6743 , 1_n6744 , 1_n6745 , 1_n6746 , 1_n6747 , 1_n6748 , 1_n6749 , 1_n6750 , 1_n6751 , 1_n6752 , 1_n6753 , 1_n6754 , 1_n6755 , 1_n6756 , 1_n6757 , 1_n6758 , 1_n6759 , 1_n6760 , 1_n6761 , 1_n6762 , 1_n6763 , 1_n6764 , 1_n6765 , 1_n6766 , 1_n6767 , 1_n6768 , 1_n6769 , 1_n6770 , 1_n6771 , 1_n6772 , 1_n6773 , 1_n6774 , 1_n6775 , 1_n6776 , 1_n6777 , 1_n6778 , 1_n6779 , 1_n6780 , 1_n6781 , 1_n6782 , 1_n6783 , 1_n6784 , 1_n6785 , 1_n6786 , 1_n6787 , 1_n6788 , 1_n6789 , 1_n6790 , 1_n6791 , 1_n6792 , 1_n6793 , 1_n6794 , 1_n6795 , 1_n6796 , 1_n6797 , 1_n6798 , 1_n6799 , 1_n6800 , 1_n6801 , 1_n6802 , 1_n6803 , 1_n6804 , 1_n6805 , 1_n6806 , 1_n6807 , 1_n6808 , 1_n6809 , 1_n6810 , 1_n6811 , 1_n6812 , 1_n6813 , 1_n6814 , 1_n6815 , 1_n6816 , 1_n6817 , 1_n6819 , 1_n6820 , 1_n6821 , 1_n6822 , 1_n6823 , 1_n6824 , 1_n6825 , 1_n6827 , 1_n6828 , 1_n6829 , 1_n6830 , 1_n6831 , 1_n6832 , 1_n6833 , 1_n6834 , 1_n6835 , 1_n6836 , 1_n6837 , 1_n6838 , 1_n6839 , 1_n6840 , 1_n6841 , 1_n6842 , 1_n6844 , 1_n6845 , 1_n6846 , 1_n6847 , 1_n6848 , 1_n6849 , 1_n6850 , 1_n6851 , 1_n6852 , 1_n6853 , 1_n6854 , 1_n6855 , 1_n6856 , 1_n6857 , 1_n6858 , 1_n6859 , 1_n6860 , 1_n6861 , 1_n6863 , 1_n6864 , 1_n6865 , 1_n6866 , 1_n6867 , 1_n6868 , 1_n6869 , 1_n6870 , 1_n6871 , 1_n6872 , 1_n6873 , 1_n6874 , 1_n6875 , 1_n6876 , 1_n6877 , 1_n6878 , 1_n6879 , 1_n6880 , 1_n6881 , 1_n6882 , 1_n6883 , 1_n6884 , 1_n6885 , 1_n6886 , 1_n6887 , 1_n6888 , 1_n6889 , 1_n6890 , 1_n6891 , 1_n6892 , 1_n6893 , 1_n6894 , 1_n6895 , 1_n6896 , 1_n6897 , 1_n6898 , 1_n6899 , 1_n6900 , 1_n6901 , 1_n6902 , 1_n6903 , 1_n6904 , 1_n6905 , 1_n6906 , 1_n6907 , 1_n6908 , 1_n6909 , 1_n6910 , 1_n6911 , 1_n6912 , 1_n6913 , 1_n6914 , 1_n6915 , 1_n6916 , 1_n6917 , 1_n6918 , 1_n6919 , 1_n6920 , 1_n6921 , 1_n6922 , 1_n6923 , 1_n6924 , 1_n6925 , 1_n6926 , 1_n6927 , 1_n6928 , 1_n6929 , 1_n6930 , 1_n6931 , 1_n6932 , 1_n6933 , 1_n6934 , 1_n6935 , 1_n6936 , 1_n6938 , 1_n6939 , 1_n6940 , 1_n6941 , 1_n6942 , 1_n6943 , 1_n6944 , 1_n6945 , 1_n6946 , 1_n6947 , 1_n6948 , 1_n6949 , 1_n6950 , 1_n6951 , 1_n6952 , 1_n6953 , 1_n6954 , 1_n6955 , 1_n6956 , 1_n6957 , 1_n6958 , 1_n6959 , 1_n6960 , 1_n6961 , 1_n6962 , 1_n6963 , 1_n6964 , 1_n6965 , 1_n6966 , 1_n6967 , 1_n6968 , 1_n6969 , 1_n6970 , 1_n6971 , 1_n6972 , 1_n6973 , 1_n6974 , 1_n6975 , 1_n6976 , 1_n6977 , 1_n6978 , 1_n6979 , 1_n6980 , 1_n6981 , 1_n6982 , 1_n6983 , 1_n6984 , 1_n6985 , 1_n6986 , 1_n6987 , 1_n6988 , 1_n6989 , 1_n6990 , 1_n6991 , 1_n6992 , 1_n6993 , 1_n6994 , 1_n6995 , 1_n6996 , 1_n6997 , 1_n6998 , 1_n6999 , 1_n7000 , 1_n7001 , 1_n7002 , 1_n7003 , 1_n7004 , 1_n7005 , 1_n7006 , 1_n7007 , 1_n7008 , 1_n7009 , 1_n7010 , 1_n7011 , 1_n7012 , 1_n7013 , 1_n7014 , 1_n7015 , 1_n7016 , 1_n7017 , 1_n7018 , 1_n7019 , 1_n7020 , 1_n7021 , 1_n7022 , 1_n7023 , 1_n7024 , 1_n7025 , 1_n7026 , 1_n7027 , 1_n7028 , 1_n7029 , 1_n7030 , 1_n7031 , 1_n7032 , 1_n7033 , 1_n7035 , 1_n7036 , 1_n7037 , 1_n7038 , 1_n7039 , 1_n7040 , 1_n7041 , 1_n7042 , 1_n7043 , 1_n7044 , 1_n7045 , 1_n7046 , 1_n7047 , 1_n7048 , 1_n7049 , 1_n7050 , 1_n7051 , 1_n7052 , 1_n7053 , 1_n7054 , 1_n7055 , 1_n7056 , 1_n7057 , 1_n7058 , 1_n7059 , 1_n7060 , 1_n7062 , 1_n7063 , 1_n7064 , 1_n7065 , 1_n7066 , 1_n7067 , 1_n7068 , 1_n7069 , 1_n7070 , 1_n7071 , 1_n7072 , 1_n7073 , 1_n7074 , 1_n7075 , 1_n7076 , 1_n7077 , 1_n7078 , 1_n7079 , 1_n7080 , 1_n7081 , 1_n7082 , 1_n7083 , 1_n7084 , 1_n7085 , 1_n7086 , 1_n7087 , 1_n7088 , 1_n7089 , 1_n7090 , 1_n7091 , 1_n7092 , 1_n7093 , 1_n7094 , 1_n7095 , 1_n7096 , 1_n7097 , 1_n7098 , 1_n7099 , 1_n7100 , 1_n7101 , 1_n7102 , 1_n7103 , 1_n7104 , 1_n7105 , 1_n7106 , 1_n7107 , 1_n7108 , 1_n7109 , 1_n7110 , 1_n7112 , 1_n7114 , 1_n7115 , 1_n7116 , 1_n7117 , 1_n7118 , 1_n7119 , 1_n7120 , 1_n7121 , 1_n7122 , 1_n7123 , 1_n7124 , 1_n7125 , 1_n7126 , 1_n7127 , 1_n7128 , 1_n7129 , 1_n7130 , 1_n7131 , 1_n7133 , 1_n7134 , 1_n7135 , 1_n7136 , 1_n7137 , 1_n7138 , 1_n7139 , 1_n7140 , 1_n7141 , 1_n7142 , 1_n7143 , 1_n7144 , 1_n7145 , 1_n7146 , 1_n7147 , 1_n7148 , 1_n7149 , 1_n7150 , 1_n7151 , 1_n7152 , 1_n7153 , 1_n7154 , 1_n7155 , 1_n7156 , 1_n7157 , 1_n7158 , 1_n7159 , 1_n7160 , 1_n7162 , 1_n7163 , 1_n7164 , 1_n7165 , 1_n7166 , 1_n7167 , 1_n7168 , 1_n7169 , 1_n7170 , 1_n7171 , 1_n7172 , 1_n7173 , 1_n7174 , 1_n7175 , 1_n7176 , 1_n7177 , 1_n7178 , 1_n7179 , 1_n7180 , 1_n7181 , 1_n7182 , 1_n7183 , 1_n7184 , 1_n7185 , 1_n7186 , 1_n7187 , 1_n7188 , 1_n7189 , 1_n7190 , 1_n7191 , 1_n7192 , 1_n7193 , 1_n7194 , 1_n7195 , 1_n7196 , 1_n7197 , 1_n7198 , 1_n7199 , 1_n7200 , 1_n7201 , 1_n7202 , 1_n7203 , 1_n7204 , 1_n7205 , 1_n7206 , 1_n7207 , 1_n7208 , 1_n7209 , 1_n7210 , 1_n7211 , 1_n7212 , 1_n7213 , 1_n7214 , 1_n7215 , 1_n7216 , 1_n7217 , 1_n7218 , 1_n7219 , 1_n7220 , 1_n7221 , 1_n7222 , 1_n7223 , 1_n7224 , 1_n7225 , 1_n7226 , 1_n7227 , 1_n7228 , 1_n7229 , 1_n7230 , 1_n7231 , 1_n7232 , 1_n7233 , 1_n7234 , 1_n7235 , 1_n7236 , 1_n7237 , 1_n7238 , 1_n7239 , 1_n7240 , 1_n7242 , 1_n7243 , 1_n7244 , 1_n7245 , 1_n7246 , 1_n7247 , 1_n7248 , 1_n7249 , 1_n7250 , 1_n7251 , 1_n7252 , 1_n7253 , 1_n7254 , 1_n7255 , 1_n7256 , 1_n7257 , 1_n7258 , 1_n7259 , 1_n7260 , 1_n7261 , 1_n7262 , 1_n7263 , 1_n7264 , 1_n7265 , 1_n7266 , 1_n7267 , 1_n7268 , 1_n7269 , 1_n7270 , 1_n7271 , 1_n7272 , 1_n7273 , 1_n7274 , 1_n7275 , 1_n7276 , 1_n7277 , 1_n7278 , 1_n7279 , 1_n7280 , 1_n7281 , 1_n7282 , 1_n7283 , 1_n7284 , 1_n7285 , 1_n7286 , 1_n7287 , 1_n7288 , 1_n7289 , 1_n7290 , 1_n7291 , 1_n7292 , 1_n7293 , 1_n7294 , 1_n7295 , 1_n7296 , 1_n7297 , 1_n7298 , 1_n7299 , 1_n7300 , 1_n7301 , 1_n7302 , 1_n7303 , 1_n7304 , 1_n7305 , 1_n7306 , 1_n7307 , 1_n7308 , 1_n7309 , 1_n7310 , 1_n7311 , 1_n7312 , 1_n7313 , 1_n7314 , 1_n7315 , 1_n7316 , 1_n7317 , 1_n7318 , 1_n7319 , 1_n7320 , 1_n7321 , 1_n7322 , 1_n7323 , 1_n7324 , 1_n7325 , 1_n7326 , 1_n7327 , 1_n7328 , 1_n7329 , 1_n7330 , 1_n7331 , 1_n7332 , 1_n7333 , 1_n7334 , 1_n7335 , 1_n7336 , 1_n7337 , 1_n7338 , 1_n7339 , 1_n7340 , 1_n7341 , 1_n7342 , 1_n7343 , 1_n7344 , 1_n7345 , 1_n7346 , 1_n7347 , 1_n7348 , 1_n7349 , 1_n7350 , 1_n7351 , 1_n7352 , 1_n7353 , 1_n7354 , 1_n7355 , 1_n7356 , 1_n7357 , 1_n7358 , 1_n7359 , 1_n7360 , 1_n7361 , 1_n7362 , 1_n7363 , 1_n7364 , 1_n7365 , 1_n7366 , 1_n7367 , 1_n7368 , 1_n7369 , 1_n7370 , 1_n7371 , 1_n7372 , 1_n7373 , 1_n7375 , 1_n7376 , 1_n7377 , 1_n7378 , 1_n7379 , 1_n7380 , 1_n7381 , 1_n7382 , 1_n7383 , 1_n7384 , 1_n7385 , 1_n7386 , 1_n7387 , 1_n7388 , 1_n7389 , 1_n7390 , 1_n7391 , 1_n7392 , 1_n7393 , 1_n7394 , 1_n7395 , 1_n7396 , 1_n7397 , 1_n7398 , 1_n7399 , 1_n7400 , 1_n7401 , 1_n7402 , 1_n7403 , 1_n7404 , 1_n7405 , 1_n7406 , 1_n7407 , 1_n7408 , 1_n7409 , 1_n7410 , 1_n7412 , 1_n7413 , 1_n7414 , 1_n7415 , 1_n7416 , 1_n7417 , 1_n7418 , 1_n7419 , 1_n7420 , 1_n7421 , 1_n7422 , 1_n7423 , 1_n7424 , 1_n7425 , 1_n7426 , 1_n7427 , 1_n7428 , 1_n7429 , 1_n7430 , 1_n7431 , 1_n7432 , 1_n7433 , 1_n7434 , 1_n7435 , 1_n7436 , 1_n7437 , 1_n7438 , 1_n7439 , 1_n7440 , 1_n7441 , 1_n7442 , 1_n7443 , 1_n7444 , 1_n7445 , 1_n7446 , 1_n7447 , 1_n7448 , 1_n7449 , 1_n7450 , 1_n7451 , 1_n7452 , 1_n7453 , 1_n7454 , 1_n7455 , 1_n7456 , 1_n7457 , 1_n7458 , 1_n7459 , 1_n7460 , 1_n7461 , 1_n7462 , 1_n7463 , 1_n7464 , 1_n7465 , 1_n7466 , 1_n7467 , 1_n7468 , 1_n7469 , 1_n7470 , 1_n7471 , 1_n7472 , 1_n7473 , 1_n7474 , 1_n7475 , 1_n7476 , 1_n7477 , 1_n7478 , 1_n7479 , 1_n7480 , 1_n7481 , 1_n7482 , 1_n7483 , 1_n7484 , 1_n7485 , 1_n7486 , 1_n7487 , 1_n7488 , 1_n7489 , 1_n7490 , 1_n7491 , 1_n7492 , 1_n7493 , 1_n7494 , 1_n7495 , 1_n7496 , 1_n7497 , 1_n7498 , 1_n7499 , 1_n7500 , 1_n7501 , 1_n7502 , 1_n7503 , 1_n7504 , 1_n7505 , 1_n7506 , 1_n7507 , 1_n7508 , 1_n7509 , 1_n7510 , 1_n7511 , 1_n7512 , 1_n7513 , 1_n7514 , 1_n7515 , 1_n7516 , 1_n7517 , 1_n7518 , 1_n7519 , 1_n7520 , 1_n7521 , 1_n7522 , 1_n7523 , 1_n7524 , 1_n7525 , 1_n7526 , 1_n7527 , 1_n7528 , 1_n7530 , 1_n7531 , 1_n7532 , 1_n7533 , 1_n7534 , 1_n7535 , 1_n7536 , 1_n7537 , 1_n7538 , 1_n7539 , 1_n7540 , 1_n7541 , 1_n7542 , 1_n7543 , 1_n7544 , 1_n7545 , 1_n7546 , 1_n7547 , 1_n7548 , 1_n7549 , 1_n7550 , 1_n7551 , 1_n7552 , 1_n7554 , 1_n7555 , 1_n7556 , 1_n7557 , 1_n7558 , 1_n7559 , 1_n7560 , 1_n7561 , 1_n7562 , 1_n7563 , 1_n7564 , 1_n7565 , 1_n7566 , 1_n7567 , 1_n7568 , 1_n7569 , 1_n7570 , 1_n7571 , 1_n7572 , 1_n7573 , 1_n7574 , 1_n7575 , 1_n7576 , 1_n7577 , 1_n7578 , 1_n7579 , 1_n7580 , 1_n7581 , 1_n7583 , 1_n7584 , 1_n7585 , 1_n7586 , 1_n7587 , 1_n7588 , 1_n7589 , 1_n7590 , 1_n7591 , 1_n7592 , 1_n7593 , 1_n7594 , 1_n7595 , 1_n7596 , 1_n7597 , 1_n7598 , 1_n7599 , 1_n7600 , 1_n7601 , 1_n7602 , 1_n7603 , 1_n7604 , 1_n7605 , 1_n7606 , 1_n7607 , 1_n7608 , 1_n7609 , 1_n7610 , 1_n7611 , 1_n7612 , 1_n7613 , 1_n7614 , 1_n7615 , 1_n7616 , 1_n7617 , 1_n7618 , 1_n7619 , 1_n7620 , 1_n7621 , 1_n7622 , 1_n7623 , 1_n7624 , 1_n7625 , 1_n7626 , 1_n7627 , 1_n7628 , 1_n7629 , 1_n7630 , 1_n7631 , 1_n7632 , 1_n7633 , 1_n7634 , 1_n7635 , 1_n7636 , 1_n7637 , 1_n7638 , 1_n7639 , 1_n7640 , 1_n7641 , 1_n7642 , 1_n7643 , 1_n7644 , 1_n7645 , 1_n7646 , 1_n7647 , 1_n7648 , 1_n7649 , 1_n7650 , 1_n7651 , 1_n7652 , 1_n7653 , 1_n7654 , 1_n7655 , 1_n7656 , 1_n7657 , 1_n7658 , 1_n7660 , 1_n7661 , 1_n7662 , 1_n7663 , 1_n7664 , 1_n7665 , 1_n7666 , 1_n7667 , 1_n7668 , 1_n7669 , 1_n7670 , 1_n7671 , 1_n7672 , 1_n7673 , 1_n7674 , 1_n7675 , 1_n7676 , 1_n7677 , 1_n7678 , 1_n7679 , 1_n7680 , 1_n7681 , 1_n7682 , 1_n7683 , 1_n7684 , 1_n7685 , 1_n7686 , 1_n7688 , 1_n7689 , 1_n7690 , 1_n7691 , 1_n7692 , 1_n7693 , 1_n7694 , 1_n7695 , 1_n7696 , 1_n7697 , 1_n7698 , 1_n7699 , 1_n7700 , 1_n7701 , 1_n7702 , 1_n7703 , 1_n7704 , 1_n7705 , 1_n7706 , 1_n7707 , 1_n7708 , 1_n7709 , 1_n7710 , 1_n7711 , 1_n7712 , 1_n7713 , 1_n7714 , 1_n7716 , 1_n7717 , 1_n7718 , 1_n7719 , 1_n7721 , 1_n7722 , 1_n7723 , 1_n7724 , 1_n7725 , 1_n7726 , 1_n7727 , 1_n7728 , 1_n7730 , 1_n7731 , 1_n7732 , 1_n7733 , 1_n7734 , 1_n7735 , 1_n7736 , 1_n7737 , 1_n7738 , 1_n7739 , 1_n7740 , 1_n7741 , 1_n7742 , 1_n7743 , 1_n7744 , 1_n7745 , 1_n7746 , 1_n7747 , 1_n7748 , 1_n7749 , 1_n7750 , 1_n7751 , 1_n7752 , 1_n7753 , 1_n7754 , 1_n7756 , 1_n7757 , 1_n7758 , 1_n7759 , 1_n7760 , 1_n7761 , 1_n7762 , 1_n7763 , 1_n7764 , 1_n7765 , 1_n7766 , 1_n7767 , 1_n7768 , 1_n7769 , 1_n7770 , 1_n7771 , 1_n7773 , 1_n7774 , 1_n7775 , 1_n7776 , 1_n7777 , 1_n7778 , 1_n7779 , 1_n7780 , 1_n7781 , 1_n7782 , 1_n7783 , 1_n7784 , 1_n7785 , 1_n7786 , 1_n7787 , 1_n7788 , 1_n7789 , 1_n7791 , 1_n7792 , 1_n7793 , 1_n7794 , 1_n7795 , 1_n7796 , 1_n7797 , 1_n7798 , 1_n7799 , 1_n7800 , 1_n7801 , 1_n7802 , 1_n7803 , 1_n7804 , 1_n7805 , 1_n7806 , 1_n7807 , 1_n7808 , 1_n7809 , 1_n7810 , 1_n7811 , 1_n7813 , 1_n7814 , 1_n7815 , 1_n7816 , 1_n7817 , 1_n7818 , 1_n7819 , 1_n7820 , 1_n7821 , 1_n7822 , 1_n7823 , 1_n7824 , 1_n7825 , 1_n7826 , 1_n7827 , 1_n7828 , 1_n7829 , 1_n7830 , 1_n7831 , 1_n7832 , 1_n7833 , 1_n7834 , 1_n7835 , 1_n7836 , 1_n7837 , 1_n7838 , 1_n7839 , 1_n7840 , 1_n7841 , 1_n7842 , 1_n7843 , 1_n7844 , 1_n7845 , 1_n7846 , 1_n7847 , 1_n7848 , 1_n7849 , 1_n7850 , 1_n7851 , 1_n7852 , 1_n7853 , 1_n7854 , 1_n7855 , 1_n7856 , 1_n7857 , 1_n7859 , 1_n7861 , 1_n7862 , 1_n7863 , 1_n7864 , 1_n7865 , 1_n7866 , 1_n7867 , 1_n7868 , 1_n7869 , 1_n7870 , 1_n7871 , 1_n7872 , 1_n7873 , 1_n7874 , 1_n7875 , 1_n7876 , 1_n7877 , 1_n7878 , 1_n7879 , 1_n7880 , 1_n7881 , 1_n7882 , 1_n7883 , 1_n7884 , 1_n7885 , 1_n7886 , 1_n7887 , 1_n7888 , 1_n7889 , 1_n7890 , 1_n7891 , 1_n7892 , 1_n7893 , 1_n7894 , 1_n7895 , 1_n7896 , 1_n7897 , 1_n7898 , 1_n7899 , 1_n7900 , 1_n7901 , 1_n7902 , 1_n7903 , 1_n7904 , 1_n7905 , 1_n7906 , 1_n7907 , 1_n7908 , 1_n7909 , 1_n7910 , 1_n7911 , 1_n7912 , 1_n7913 , 1_n7914 , 1_n7915 , 1_n7916 , 1_n7917 , 1_n7918 , 1_n7919 , 1_n7920 , 1_n7921 , 1_n7922 , 1_n7923 , 1_n7924 , 1_n7925 , 1_n7926 , 1_n7927 , 1_n7928 , 1_n7929 , 1_n7930 , 1_n7931 , 1_n7932 , 1_n7933 , 1_n7934 , 1_n7935 , 1_n7936 , 1_n7937 , 1_n7938 , 1_n7939 , 1_n7940 , 1_n7941 , 1_n7942 , 1_n7943 , 1_n7944 , 1_n7945 , 1_n7946 , 1_n7947 , 1_n7948 , 1_n7949 , 1_n7950 , 1_n7951 , 1_n7952 , 1_n7953 , 1_n7954 , 1_n7955 , 1_n7956 , 1_n7957 , 1_n7958 , 1_n7959 , 1_n7960 , 1_n7961 , 1_n7962 , 1_n7963 , 1_n7964 , 1_n7965 , 1_n7966 , 1_n7967 , 1_n7969 , 1_n7970 , 1_n7971 , 1_n7972 , 1_n7973 , 1_n7975 , 1_n7976 , 1_n7977 , 1_n7978 , 1_n7979 , 1_n7980 , 1_n7981 , 1_n7982 , 1_n7983 , 1_n7984 , 1_n7985 , 1_n7986 , 1_n7987 , 1_n7988 , 1_n7989 , 1_n7990 , 1_n7991 , 1_n7992 , 1_n7993 , 1_n7994 , 1_n7995 , 1_n7996 , 1_n7997 , 1_n7998 , 1_n7999 , 1_n8000 , 1_n8001 , 1_n8002 , 1_n8003 , 1_n8004 , 1_n8005 , 1_n8006 , 1_n8007 , 1_n8008 , 1_n8009 , 1_n8010 , 1_n8011 , 1_n8012 , 1_n8013 , 1_n8014 , 1_n8015 , 1_n8016 , 1_n8017 , 1_n8018 , 1_n8019 , 1_n8020 , 1_n8021 , 1_n8022 , 1_n8023 , 1_n8024 , 1_n8025 , 1_n8026 , 1_n8027 , 1_n8028 , 1_n8029 , 1_n8030 , 1_n8031 , 1_n8032 , 1_n8033 , 1_n8034 , 1_n8035 , 1_n8036 , 1_n8037 , 1_n8038 , 1_n8039 , 1_n8040 , 1_n8041 , 1_n8042 , 1_n8043 , 1_n8044 , 1_n8045 , 1_n8046 , 1_n8047 , 1_n8048 , 1_n8049 , 1_n8050 , 1_n8051 , 1_n8052 , 1_n8053 , 1_n8054 , 1_n8055 , 1_n8056 , 1_n8057 , 1_n8058 , 1_n8059 , 1_n8060 , 1_n8061 , 1_n8062 , 1_n8063 , 1_n8064 , 1_n8065 , 1_n8066 , 1_n8067 , 1_n8068 , 1_n8069 , 1_n8070 , 1_n8071 , 1_n8072 , 1_n8073 , 1_n8074 , 1_n8075 , 1_n8076 , 1_n8077 , 1_n8078 , 1_n8079 , 1_n8080 , 1_n8081 , 1_n8082 , 1_n8083 , 1_n8084 , 1_n8085 , 1_n8086 , 1_n8087 , 1_n8088 , 1_n8089 , 1_n8090 , 1_n8091 , 1_n8092 , 1_n8093 , 1_n8094 , 1_n8095 , 1_n8096 , 1_n8097 , 1_n8098 , 1_n8099 , 1_n8100 , 1_n8101 , 1_n8102 , 1_n8103 , 1_n8104 , 1_n8105 , 1_n8106 , 1_n8107 , 1_n8108 , 1_n8109 , 1_n8110 , 1_n8111 , 1_n8112 , 1_n8113 , 1_n8114 , 1_n8115 , 1_n8116 , 1_n8117 , 1_n8118 , 1_n8119 , 1_n8120 , 1_n8121 , 1_n8122 , 1_n8123 , 1_n8124 , 1_n8125 , 1_n8126 , 1_n8127 , 1_n8128 , 1_n8129 , 1_n8130 , 1_n8131 , 1_n8132 , 1_n8133 , 1_n8134 , 1_n8135 , 1_n8136 , 1_n8137 , 1_n8138 , 1_n8140 , 1_n8141 , 1_n8142 , 1_n8143 , 1_n8144 , 1_n8145 , 1_n8146 , 1_n8147 , 1_n8148 , 1_n8149 , 1_n8150 , 1_n8151 , 1_n8152 , 1_n8153 , 1_n8154 , 1_n8155 , 1_n8156 , 1_n8157 , 1_n8158 , 1_n8159 , 1_n8160 , 1_n8161 , 1_n8162 , 1_n8164 , 1_n8165 , 1_n8166 , 1_n8167 , 1_n8168 , 1_n8169 , 1_n8170 , 1_n8171 , 1_n8173 , 1_n8174 , 1_n8175 , 1_n8176 , 1_n8177 , 1_n8178 , 1_n8179 , 1_n8180 , 1_n8181 , 1_n8182 , 1_n8184 , 1_n8185 , 1_n8186 , 1_n8187 , 1_n8188 , 1_n8189 , 1_n8190 , 1_n8191 , 1_n8192 , 1_n8193 , 1_n8194 , 1_n8195 , 1_n8196 , 1_n8197 , 1_n8198 , 1_n8199 , 1_n8200 , 1_n8201 , 1_n8202 , 1_n8203 , 1_n8204 , 1_n8205 , 1_n8206 , 1_n8207 , 1_n8208 , 1_n8209 , 1_n8210 , 1_n8211 , 1_n8212 , 1_n8213 , 1_n8214 , 1_n8215 , 1_n8216 , 1_n8217 , 1_n8218 , 1_n8220 , 1_n8221 , 1_n8222 , 1_n8223 , 1_n8224 , 1_n8225 , 1_n8226 , 1_n8227 , 1_n8229 , 1_n8231 , 1_n8232 , 1_n8234 , 1_n8235 , 1_n8236 , 1_n8237 , 1_n8238 , 1_n8239 , 1_n8240 , 1_n8241 , 1_n8242 , 1_n8243 , 1_n8244 , 1_n8245 , 1_n8246 , 1_n8247 , 1_n8248 , 1_n8249 , 1_n8250 , 1_n8251 , 1_n8252 , 1_n8253 , 1_n8254 , 1_n8255 , 1_n8256 , 1_n8257 , 1_n8258 , 1_n8259 , 1_n8260 , 1_n8261 , 1_n8262 , 1_n8263 , 1_n8264 , 1_n8266 , 1_n8267 , 1_n8268 , 1_n8269 , 1_n8270 , 1_n8271 , 1_n8272 , 1_n8273 , 1_n8274 , 1_n8275 , 1_n8276 , 1_n8277 , 1_n8278 , 1_n8279 , 1_n8280 , 1_n8281 , 1_n8282 , 1_n8283 , 1_n8284 , 1_n8285 , 1_n8286 , 1_n8287 , 1_n8288 , 1_n8289 , 1_n8291 , 1_n8292 , 1_n8293 , 1_n8294 , 1_n8295 , 1_n8296 , 1_n8297 , 1_n8298 , 1_n8299 , 1_n8300 , 1_n8301 , 1_n8302 , 1_n8303 , 1_n8304 , 1_n8305 , 1_n8306 , 1_n8307 , 1_n8309 , 1_n8310 , 1_n8311 , 1_n8312 , 1_n8313 , 1_n8314 , 1_n8315 , 1_n8316 , 1_n8317 , 1_n8318 , 1_n8319 , 1_n8320 , 1_n8321 , 1_n8322 , 1_n8323 , 1_n8324 , 1_n8325 , 1_n8326 , 1_n8327 , 1_n8328 , 1_n8329 , 1_n8330 , 1_n8331 , 1_n8333 , 1_n8334 , 1_n8335 , 1_n8337 , 1_n8338 , 1_n8339 , 1_n8340 , 1_n8341 , 1_n8342 , 1_n8343 , 1_n8344 , 1_n8345 , 1_n8346 , 1_n8347 , 1_n8348 , 1_n8349 , 1_n8350 , 1_n8351 , 1_n8352 , 1_n8353 , 1_n8354 , 1_n8355 , 1_n8356 , 1_n8357 , 1_n8358 , 1_n8359 , 1_n8360 , 1_n8361 , 1_n8362 , 1_n8363 , 1_n8364 , 1_n8365 , 1_n8366 , 1_n8367 , 1_n8368 , 1_n8369 , 1_n8370 , 1_n8371 , 1_n8372 , 1_n8373 , 1_n8374 , 1_n8375 , 1_n8376 , 1_n8377 , 1_n8378 , 1_n8379 , 1_n8380 , 1_n8381 , 1_n8382 , 1_n8383 , 1_n8384 , 1_n8385 , 1_n8386 , 1_n8387 , 1_n8388 , 1_n8389 , 1_n8390 , 1_n8391 , 1_n8392 , 1_n8393 , 1_n8394 , 1_n8395 , 1_n8396 , 1_n8397 , 1_n8398 , 1_n8399 , 1_n8400 , 1_n8401 , 1_n8402 , 1_n8403 , 1_n8404 , 1_n8405 , 1_n8406 , 1_n8407 , 1_n8408 , 1_n8409 , 1_n8410 , 1_n8411 , 1_n8412 , 1_n8413 , 1_n8414 , 1_n8415 , 1_n8416 , 1_n8417 , 1_n8418 , 1_n8419 , 1_n8420 , 1_n8421 , 1_n8422 , 1_n8423 , 1_n8424 , 1_n8425 , 1_n8426 , 1_n8427 , 1_n8428 , 1_n8429 , 1_n8430 , 1_n8431 , 1_n8432 , 1_n8433 , 1_n8434 , 1_n8435 , 1_n8436 , 1_n8437 , 1_n8438 , 1_n8439 , 1_n8440 , 1_n8441 , 1_n8442 , 1_n8443 , 1_n8444 , 1_n8445 , 1_n8446 , 1_n8447 , 1_n8448 , 1_n8449 , 1_n8450 , 1_n8451 , 1_n8452 , 1_n8453 , 1_n8454 , 1_n8455 , 1_n8456 , 1_n8457 , 1_n8458 , 1_n8459 , 1_n8460 , 1_n8461 , 1_n8462 , 1_n8463 , 1_n8464 , 1_n8465 , 1_n8467 , 1_n8469 , 1_n8470 , 1_n8471 , 1_n8472 , 1_n8473 , 1_n8474 , 1_n8475 , 1_n8476 , 1_n8477 , 1_n8478 , 1_n8479 , 1_n8480 , 1_n8481 , 1_n8482 , 1_n8483 , 1_n8484 , 1_n8485 , 1_n8486 , 1_n8487 , 1_n8488 , 1_n8489 , 1_n8490 , 1_n8491 , 1_n8492 , 1_n8493 , 1_n8494 , 1_n8495 , 1_n8496 , 1_n8497 , 1_n8498 , 1_n8499 , 1_n8500 , 1_n8501 , 1_n8502 , 1_n8503 , 1_n8504 , 1_n8505 , 1_n8507 , 1_n8508 , 1_n8509 , 1_n8510 , 1_n8511 , 1_n8512 , 1_n8513 , 1_n8514 , 1_n8515 , 1_n8517 , 1_n8518 , 1_n8519 , 1_n8520 , 1_n8521 , 1_n8523 , 1_n8524 , 1_n8525 , 1_n8526 , 1_n8527 , 1_n8528 , 1_n8529 , 1_n8530 , 1_n8531 , 1_n8532 , 1_n8533 , 1_n8534 , 1_n8535 , 1_n8536 , 1_n8537 , 1_n8538 , 1_n8539 , 1_n8540 , 1_n8541 , 1_n8542 , 1_n8543 , 1_n8544 , 1_n8545 , 1_n8546 , 1_n8547 , 1_n8548 , 1_n8549 , 1_n8550 , 1_n8551 , 1_n8552 , 1_n8553 , 1_n8554 , 1_n8555 , 1_n8556 , 1_n8557 , 1_n8558 , 1_n8559 , 1_n8560 , 1_n8561 , 1_n8562 , 1_n8563 , 1_n8564 , 1_n8565 , 1_n8566 , 1_n8567 , 1_n8568 , 1_n8569 , 1_n8570 , 1_n8571 , 1_n8572 , 1_n8573 , 1_n8574 , 1_n8575 , 1_n8576 , 1_n8577 , 1_n8578 , 1_n8579 , 1_n8580 , 1_n8581 , 1_n8582 , 1_n8583 , 1_n8584 , 1_n8585 , 1_n8586 , 1_n8587 , 1_n8588 , 1_n8589 , 1_n8590 , 1_n8591 , 1_n8592 , 1_n8593 , 1_n8594 , 1_n8595 , 1_n8596 , 1_n8597 , 1_n8598 , 1_n8599 , 1_n8600 , 1_n8601 , 1_n8602 , 1_n8603 , 1_n8604 , 1_n8605 , 1_n8606 , 1_n8607 , 1_n8608 , 1_n8609 , 1_n8610 , 1_n8611 , 1_n8612 , 1_n8613 , 1_n8614 , 1_n8615 , 1_n8616 , 1_n8617 , 1_n8618 , 1_n8619 , 1_n8620 , 1_n8621 , 1_n8622 , 1_n8623 , 1_n8624 , 1_n8625 , 1_n8626 , 1_n8627 , 1_n8628 , 1_n8629 , 1_n8630 , 1_n8631 , 1_n8632 , 1_n8633 , 1_n8634 , 1_n8635 , 1_n8636 , 1_n8637 , 1_n8638 , 1_n8639 , 1_n8640 , 1_n8641 , 1_n8642 , 1_n8643 , 1_n8644 , 1_n8645 , 1_n8646 , 1_n8647 , 1_n8648 , 1_n8649 , 1_n8650 , 1_n8651 , 1_n8652 , 1_n8653 , 1_n8654 , 1_n8655 , 1_n8656 , 1_n8657 , 1_n8658 , 1_n8659 , 1_n8660 , 1_n8661 , 1_n8662 , 1_n8663 , 1_n8664 , 1_n8665 , 1_n8666 , 1_n8667 , 1_n8668 , 1_n8669 , 1_n8670 , 1_n8671 , 1_n8672 , 1_n8673 , 1_n8674 , 1_n8675 , 1_n8676 , 1_n8677 , 1_n8678 , 1_n8679 , 1_n8680 , 1_n8681 , 1_n8682 , 1_n8683 , 1_n8684 , 1_n8685 , 1_n8686 , 1_n8687 , 1_n8688 , 1_n8689 , 1_n8690 , 1_n8691 , 1_n8692 , 1_n8693 , 1_n8694 , 1_n8695 , 1_n8696 , 1_n8697 , 1_n8698 , 1_n8699 , 1_n8700 , 1_n8702 , 1_n8703 , 1_n8704 , 1_n8705 , 1_n8706 , 1_n8707 , 1_n8708 , 1_n8709 , 1_n8710 , 1_n8711 , 1_n8712 , 1_n8713 , 1_n8714 , 1_n8715 , 1_n8717 , 1_n8718 , 1_n8719 , 1_n8720 , 1_n8721 , 1_n8722 , 1_n8723 , 1_n8724 , 1_n8725 , 1_n8726 , 1_n8727 , 1_n8728 , 1_n8729 , 1_n8730 , 1_n8731 , 1_n8732 , 1_n8733 , 1_n8734 , 1_n8735 , 1_n8736 , 1_n8737 , 1_n8738 , 1_n8739 , 1_n8740 , 1_n8741 , 1_n8742 , 1_n8743 , 1_n8744 , 1_n8745 , 1_n8746 , 1_n8747 , 1_n8748 , 1_n8749 , 1_n8750 , 1_n8751 , 1_n8752 , 1_n8753 , 1_n8754 , 1_n8755 , 1_n8756 , 1_n8757 , 1_n8758 , 1_n8759 , 1_n8760 , 1_n8761 , 1_n8762 , 1_n8763 , 1_n8764 , 1_n8765 , 1_n8766 , 1_n8767 , 1_n8769 , 1_n8770 , 1_n8771 , 1_n8772 , 1_n8773 , 1_n8774 , 1_n8775 , 1_n8776 , 1_n8777 , 1_n8778 , 1_n8779 , 1_n8780 , 1_n8781 , 1_n8782 , 1_n8783 , 1_n8784 , 1_n8785 , 1_n8786 , 1_n8787 , 1_n8788 , 1_n8789 , 1_n8790 , 1_n8791 , 1_n8792 , 1_n8793 , 1_n8794 , 1_n8795 , 1_n8796 , 1_n8797 , 1_n8798 , 1_n8799 , 1_n8800 , 1_n8801 , 1_n8802 , 1_n8803 , 1_n8804 , 1_n8805 , 1_n8806 , 1_n8807 , 1_n8808 , 1_n8809 , 1_n8810 , 1_n8811 , 1_n8812 , 1_n8813 , 1_n8814 , 1_n8815 , 1_n8816 , 1_n8817 , 1_n8818 , 1_n8819 , 1_n8821 , 1_n8822 , 1_n8823 , 1_n8824 , 1_n8825 , 1_n8826 , 1_n8827 , 1_n8828 , 1_n8829 , 1_n8830 , 1_n8831 , 1_n8832 , 1_n8833 , 1_n8834 , 1_n8835 , 1_n8836 , 1_n8837 , 1_n8838 , 1_n8839 , 1_n8840 , 1_n8841 , 1_n8842 , 1_n8843 , 1_n8844 , 1_n8845 , 1_n8846 , 1_n8847 , 1_n8848 , 1_n8849 , 1_n8850 , 1_n8851 , 1_n8852 , 1_n8853 , 1_n8854 , 1_n8855 , 1_n8856 , 1_n8857 , 1_n8858 , 1_n8861 , 1_n8862 , 1_n8863 , 1_n8864 , 1_n8865 , 1_n8866 , 1_n8867 , 1_n8868 , 1_n8869 , 1_n8870 , 1_n8871 , 1_n8872 , 1_n8873 , 1_n8874 , 1_n8875 , 1_n8876 , 1_n8877 , 1_n8878 , 1_n8879 , 1_n8880 , 1_n8881 , 1_n8882 , 1_n8883 , 1_n8884 , 1_n8885 , 1_n8886 , 1_n8887 , 1_n8888 , 1_n8889 , 1_n8890 , 1_n8891 , 1_n8892 , 1_n8893 , 1_n8894 , 1_n8895 , 1_n8896 , 1_n8897 , 1_n8898 , 1_n8899 , 1_n8900 , 1_n8901 , 1_n8902 , 1_n8903 , 1_n8904 , 1_n8905 , 1_n8906 , 1_n8907 , 1_n8908 , 1_n8909 , 1_n8910 , 1_n8911 , 1_n8912 , 1_n8913 , 1_n8914 , 1_n8915 , 1_n8916 , 1_n8917 , 1_n8918 , 1_n8919 , 1_n8920 , 1_n8921 , 1_n8922 , 1_n8923 , 1_n8924 , 1_n8925 , 1_n8926 , 1_n8927 , 1_n8928 , 1_n8929 , 1_n8930 , 1_n8931 , 1_n8932 , 1_n8933 , 1_n8934 , 1_n8935 , 1_n8936 , 1_n8937 , 1_n8938 , 1_n8939 , 1_n8941 , 1_n8942 , 1_n8943 , 1_n8944 , 1_n8945 , 1_n8946 , 1_n8947 , 1_n8948 , 1_n8949 , 1_n8950 , 1_n8951 , 1_n8952 , 1_n8953 , 1_n8954 , 1_n8955 , 1_n8956 , 1_n8957 , 1_n8958 , 1_n8959 , 1_n8960 , 1_n8961 , 1_n8962 , 1_n8963 , 1_n8964 , 1_n8965 , 1_n8966 , 1_n8967 , 1_n8968 , 1_n8969 , 1_n8970 , 1_n8971 , 1_n8972 , 1_n8973 , 1_n8974 , 1_n8975 , 1_n8976 , 1_n8977 , 1_n8978 , 1_n8979 , 1_n8980 , 1_n8981 , 1_n8982 , 1_n8983 , 1_n8984 , 1_n8985 , 1_n8986 , 1_n8987 , 1_n8988 , 1_n8989 , 1_n8990 , 1_n8991 , 1_n8992 , 1_n8993 , 1_n8994 , 1_n8995 , 1_n8996 , 1_n8997 , 1_n8998 , 1_n8999 , 1_n9000 , 1_n9001 , 1_n9002 , 1_n9003 , 1_n9004 , 1_n9005 , 1_n9006 , 1_n9007 , 1_n9008 , 1_n9009 , 1_n9010 , 1_n9011 , 1_n9012 , 1_n9013 , 1_n9014 , 1_n9015 , 1_n9016 , 1_n9017 , 1_n9018 , 1_n9019 , 1_n9020 , 1_n9021 , 1_n9022 , 1_n9023 , 1_n9024 , 1_n9025 , 1_n9026 , 1_n9027 , 1_n9028 , 1_n9029 , 1_n9030 , 1_n9031 , 1_n9032 , 1_n9033 , 1_n9034 , 1_n9035 , 1_n9036 , 1_n9037 , 1_n9038 , 1_n9039 , 1_n9040 , 1_n9042 , 1_n9043 , 1_n9044 , 1_n9045 , 1_n9046 , 1_n9047 , 1_n9048 , 1_n9049 , 1_n9050 , 1_n9051 , 1_n9052 , 1_n9053 , 1_n9054 , 1_n9055 , 1_n9056 , 1_n9057 , 1_n9058 , 1_n9059 , 1_n9060 , 1_n9061 , 1_n9062 , 1_n9063 , 1_n9064 , 1_n9065 , 1_n9066 , 1_n9067 , 1_n9068 , 1_n9069 , 1_n9070 , 1_n9071 , 1_n9072 , 1_n9073 , 1_n9074 , 1_n9075 , 1_n9076 , 1_n9077 , 1_n9078 , 1_n9079 , 1_n9080 , 1_n9081 , 1_n9082 , 1_n9083 , 1_n9084 , 1_n9085 , 1_n9086 , 1_n9087 , 1_n9088 , 1_n9089 , 1_n9090 , 1_n9091 , 1_n9092 , 1_n9094 , 1_n9095 , 1_n9096 , 1_n9097 , 1_n9098 , 1_n9099 , 1_n9101 , 1_n9102 , 1_n9103 , 1_n9104 , 1_n9105 , 1_n9106 , 1_n9107 , 1_n9108 , 1_n9109 , 1_n9110 , 1_n9111 , 1_n9112 , 1_n9113 , 1_n9114 , 1_n9115 , 1_n9116 , 1_n9117 , 1_n9118 , 1_n9119 , 1_n9120 , 1_n9121 , 1_n9122 , 1_n9123 , 1_n9124 , 1_n9125 , 1_n9126 , 1_n9127 , 1_n9128 , 1_n9129 , 1_n9130 , 1_n9131 , 1_n9132 , 1_n9133 , 1_n9134 , 1_n9135 , 1_n9136 , 1_n9137 , 1_n9138 , 1_n9139 , 1_n9140 , 1_n9141 , 1_n9142 , 1_n9143 , 1_n9144 , 1_n9145 , 1_n9146 , 1_n9147 , 1_n9148 , 1_n9149 , 1_n9150 , 1_n9151 , 1_n9152 , 1_n9153 , 1_n9154 , 1_n9155 , 1_n9156 , 1_n9157 , 1_n9158 , 1_n9159 , 1_n9160 , 1_n9161 , 1_n9162 , 1_n9163 , 1_n9164 , 1_n9165 , 1_n9166 , 1_n9167 , 1_n9168 , 1_n9169 , 1_n9170 , 1_n9171 , 1_n9172 , 1_n9173 , 1_n9174 , 1_n9175 , 1_n9176 , 1_n9177 , 1_n9178 , 1_n9179 , 1_n9180 , 1_n9181 , 1_n9182 , 1_n9183 , 1_n9184 , 1_n9185 , 1_n9186 , 1_n9188 , 1_n9189 , 1_n9190 , 1_n9191 , 1_n9192 , 1_n9193 , 1_n9194 , 1_n9195 , 1_n9196 , 1_n9197 , 1_n9198 , 1_n9199 , 1_n9200 , 1_n9201 , 1_n9202 , 1_n9203 , 1_n9204 , 1_n9205 , 1_n9206 , 1_n9207 , 1_n9208 , 1_n9209 , 1_n9210 , 1_n9211 , 1_n9212 , 1_n9213 , 1_n9214 , 1_n9215 , 1_n9217 , 1_n9218 , 1_n9219 , 1_n9220 , 1_n9221 , 1_n9222 , 1_n9223 , 1_n9224 , 1_n9225 , 1_n9226 , 1_n9227 , 1_n9228 , 1_n9229 , 1_n9230 , 1_n9231 , 1_n9232 , 1_n9233 , 1_n9234 , 1_n9235 , 1_n9236 , 1_n9237 , 1_n9238 , 1_n9239 , 1_n9240 , 1_n9241 , 1_n9242 , 1_n9243 , 1_n9244 , 1_n9245 , 1_n9246 , 1_n9247 , 1_n9248 , 1_n9249 , 1_n9250 , 1_n9251 , 1_n9252 , 1_n9253 , 1_n9254 , 1_n9255 , 1_n9256 , 1_n9257 , 1_n9258 , 1_n9259 , 1_n9260 , 1_n9261 , 1_n9262 , 1_n9263 , 1_n9264 , 1_n9265 , 1_n9266 , 1_n9267 , 1_n9268 , 1_n9269 , 1_n9270 , 1_n9271 , 1_n9272 , 1_n9273 , 1_n9274 , 1_n9275 , 1_n9276 , 1_n9277 , 1_n9278 , 1_n9279 , 1_n9280 , 1_n9281 , 1_n9282 , 1_n9283 , 1_n9284 , 1_n9285 , 1_n9286 , 1_n9287 , 1_n9288 , 1_n9289 , 1_n9290 , 1_n9291 , 1_n9292 , 1_n9293 , 1_n9294 , 1_n9295 , 1_n9296 , 1_n9297 , 1_n9298 , 1_n9299 , 1_n9301 , 1_n9302 , 1_n9303 , 1_n9304 , 1_n9305 , 1_n9306 , 1_n9307 , 1_n9308 , 1_n9309 , 1_n9310 , 1_n9311 , 1_n9312 , 1_n9313 , 1_n9314 , 1_n9315 , 1_n9316 , 1_n9317 , 1_n9318 , 1_n9319 , 1_n9320 , 1_n9321 , 1_n9322 , 1_n9323 , 1_n9324 , 1_n9325 , 1_n9326 , 1_n9327 , 1_n9328 , 1_n9330 , 1_n9331 , 1_n9332 , 1_n9333 , 1_n9334 , 1_n9335 , 1_n9336 , 1_n9337 , 1_n9338 , 1_n9339 , 1_n9340 , 1_n9341 , 1_n9342 , 1_n9343 , 1_n9344 , 1_n9345 , 1_n9346 , 1_n9347 , 1_n9348 , 1_n9349 , 1_n9350 , 1_n9351 , 1_n9352 , 1_n9354 , 1_n9355 , 1_n9356 , 1_n9357 , 1_n9358 , 1_n9359 , 1_n9360 , 1_n9361 , 1_n9362 , 1_n9363 , 1_n9364 , 1_n9365 , 1_n9366 , 1_n9367 , 1_n9368 , 1_n9369 , 1_n9370 , 1_n9371 , 1_n9372 , 1_n9373 , 1_n9374 , 1_n9375 , 1_n9376 , 1_n9377 , 1_n9378 , 1_n9379 , 1_n9380 , 1_n9381 , 1_n9382 , 1_n9383 , 1_n9384 , 1_n9385 , 1_n9386 , 1_n9387 , 1_n9388 , 1_n9389 , 1_n9390 , 1_n9391 , 1_n9392 , 1_n9393 , 1_n9394 , 1_n9395 , 1_n9396 , 1_n9397 , 1_n9398 , 1_n9399 , 1_n9400 , 1_n9401 , 1_n9402 , 1_n9403 , 1_n9404 , 1_n9405 , 1_n9406 , 1_n9407 , 1_n9408 , 1_n9409 , 1_n9410 , 1_n9411 , 1_n9412 , 1_n9413 , 1_n9414 , 1_n9415 , 1_n9416 , 1_n9417 , 1_n9418 , 1_n9419 , 1_n9420 , 1_n9421 , 1_n9422 , 1_n9423 , 1_n9424 , 1_n9425 , 1_n9426 , 1_n9427 , 1_n9428 , 1_n9429 , 1_n9430 , 1_n9431 , 1_n9432 , 1_n9433 , 1_n9434 , 1_n9435 , 1_n9436 , 1_n9437 , 1_n9438 , 1_n9439 , 1_n9440 , 1_n9441 , 1_n9442 , 1_n9443 , 1_n9444 , 1_n9445 , 1_n9446 , 1_n9447 , 1_n9448 , 1_n9449 , 1_n9450 , 1_n9451 , 1_n9452 , 1_n9453 , 1_n9454 , 1_n9455 , 1_n9456 , 1_n9457 , 1_n9458 , 1_n9459 , 1_n9460 , 1_n9461 , 1_n9462 , 1_n9463 , 1_n9464 , 1_n9465 , 1_n9466 , 1_n9467 , 1_n9468 , 1_n9469 , 1_n9470 , 1_n9471 , 1_n9472 , 1_n9473 , 1_n9474 , 1_n9476 , 1_n9477 , 1_n9478 , 1_n9479 , 1_n9480 , 1_n9481 , 1_n9482 , 1_n9483 , 1_n9484 , 1_n9485 , 1_n9486 , 1_n9487 , 1_n9488 , 1_n9489 , 1_n9490 , 1_n9491 , 1_n9492 , 1_n9493 , 1_n9494 , 1_n9495 , 1_n9496 , 1_n9497 , 1_n9498 , 1_n9499 , 1_n9500 , 1_n9501 , 1_n9502 , 1_n9503 , 1_n9504 , 1_n9505 , 1_n9506 , 1_n9507 , 1_n9508 , 1_n9509 , 1_n9510 , 1_n9511 , 1_n9512 , 1_n9513 , 1_n9514 , 1_n9515 , 1_n9516 , 1_n9517 , 1_n9518 , 1_n9519 , 1_n9520 , 1_n9521 , 1_n9522 , 1_n9523 , 1_n9524 , 1_n9525 , 1_n9526 , 1_n9527 , 1_n9529 , 1_n9530 , 1_n9532 , 1_n9533 , 1_n9534 , 1_n9535 , 1_n9536 , 1_n9537 , 1_n9538 , 1_n9539 , 1_n9540 , 1_n9541 , 1_n9542 , 1_n9543 , 1_n9544 , 1_n9545 , 1_n9546 , 1_n9547 , 1_n9548 , 1_n9549 , 1_n9550 , 1_n9551 , 1_n9552 , 1_n9553 , 1_n9554 , 1_n9555 , 1_n9556 , 1_n9557 , 1_n9558 , 1_n9559 , 1_n9560 , 1_n9561 , 1_n9562 , 1_n9563 , 1_n9564 , 1_n9565 , 1_n9566 , 1_n9567 , 1_n9568 , 1_n9569 , 1_n9571 , 1_n9572 , 1_n9573 , 1_n9574 , 1_n9575 , 1_n9576 , 1_n9577 , 1_n9578 , 1_n9579 , 1_n9580 , 1_n9581 , 1_n9582 , 1_n9583 , 1_n9584 , 1_n9585 , 1_n9586 , 1_n9587 , 1_n9588 , 1_n9589 , 1_n9590 , 1_n9592 , 1_n9593 , 1_n9594 , 1_n9595 , 1_n9596 , 1_n9597 , 1_n9598 , 1_n9599 , 1_n9600 , 1_n9601 , 1_n9602 , 1_n9603 , 1_n9604 , 1_n9605 , 1_n9606 , 1_n9607 , 1_n9608 , 1_n9609 , 1_n9610 , 1_n9611 , 1_n9612 , 1_n9613 , 1_n9614 , 1_n9615 , 1_n9616 , 1_n9617 , 1_n9618 , 1_n9619 , 1_n9621 , 1_n9622 , 1_n9623 , 1_n9624 , 1_n9625 , 1_n9626 , 1_n9627 , 1_n9628 , 1_n9629 , 1_n9630 , 1_n9631 , 1_n9632 , 1_n9633 , 1_n9634 , 1_n9635 , 1_n9636 , 1_n9637 , 1_n9638 , 1_n9639 , 1_n9640 , 1_n9641 , 1_n9642 , 1_n9643 , 1_n9644 , 1_n9645 , 1_n9646 , 1_n9647 , 1_n9648 , 1_n9649 , 1_n9650 , 1_n9651 , 1_n9652 , 1_n9653 , 1_n9654 , 1_n9655 , 1_n9656 , 1_n9657 , 1_n9658 , 1_n9659 , 1_n9660 , 1_n9661 , 1_n9662 , 1_n9663 , 1_n9664 , 1_n9665 , 1_n9666 , 1_n9667 , 1_n9668 , 1_n9670 , 1_n9671 , 1_n9672 , 1_n9673 , 1_n9674 , 1_n9675 , 1_n9676 , 1_n9677 , 1_n9678 , 1_n9679 , 1_n9680 , 1_n9681 , 1_n9682 , 1_n9683 , 1_n9684 , 1_n9685 , 1_n9686 , 1_n9687 , 1_n9688 , 1_n9689 , 1_n9690 , 1_n9691 , 1_n9692 , 1_n9693 , 1_n9694 , 1_n9695 , 1_n9696 , 1_n9697 , 1_n9698 , 1_n9699 , 1_n9700 , 1_n9701 , 1_n9702 , 1_n9703 , 1_n9704 , 1_n9705 , 1_n9706 , 1_n9707 , 1_n9708 , 1_n9709 , 1_n9710 , 1_n9711 , 1_n9712 , 1_n9713 , 1_n9714 , 1_n9715 , 1_n9716 , 1_n9717 , 1_n9718 , 1_n9719 , 1_n9720 , 1_n9721 , 1_n9722 , 1_n9723 , 1_n9724 , 1_n9725 , 1_n9726 , 1_n9727 , 1_n9728 , 1_n9729 , 1_n9730 , 1_n9731 , 1_n9733 , 1_n9734 , 1_n9735 , 1_n9736 , 1_n9737 , 1_n9738 , 1_n9739 , 1_n9740 , 1_n9741 , 1_n9742 , 1_n9743 , 1_n9744 , 1_n9745 , 1_n9746 , 1_n9748 , 1_n9749 , 1_n9750 , 1_n9751 , 1_n9752 , 1_n9753 , 1_n9754 , 1_n9755 , 1_n9756 , 1_n9757 , 1_n9758 , 1_n9759 , 1_n9760 , 1_n9761 , 1_n9762 , 1_n9763 , 1_n9764 , 1_n9765 , 1_n9766 , 1_n9767 , 1_n9768 , 1_n9769 , 1_n9770 , 1_n9771 , 1_n9772 , 1_n9773 , 1_n9774 , 1_n9775 , 1_n9776 , 1_n9777 , 1_n9778 , 1_n9779 , 1_n9780 , 1_n9781 , 1_n9782 , 1_n9783 , 1_n9784 , 1_n9785 , 1_n9786 , 1_n9787 , 1_n9788 , 1_n9789 , 1_n9790 , 1_n9791 , 1_n9792 , 1_n9793 , 1_n9794 , 1_n9795 , 1_n9796 , 1_n9797 , 1_n9798 , 1_n9799 , 1_n9800 , 1_n9801 , 1_n9802 , 1_n9803 , 1_n9804 , 1_n9805 , 1_n9806 , 1_n9807 , 1_n9808 , 1_n9809 , 1_n9810 , 1_n9811 , 1_n9812 , 1_n9813 , 1_n9814 , 1_n9815 , 1_n9816 , 1_n9817 , 1_n9818 , 1_n9819 , 1_n9820 , 1_n9821 , 1_n9822 , 1_n9823 , 1_n9824 , 1_n9825 , 1_n9826 , 1_n9827 , 1_n9828 , 1_n9829 , 1_n9830 , 1_n9831 , 1_n9832 , 1_n9833 , 1_n9834 , 1_n9835 , 1_n9836 , 1_n9837 , 1_n9838 , 1_n9839 , 1_n9840 , 1_n9841 , 1_n9842 , 1_n9843 , 1_n9844 , 1_n9845 , 1_n9847 , 1_n9848 , 1_n9849 , 1_n9850 , 1_n9851 , 1_n9852 , 1_n9853 , 1_n9854 , 1_n9855 , 1_n9856 , 1_n9857 , 1_n9858 , 1_n9859 , 1_n9860 , 1_n9861 , 1_n9862 , 1_n9863 , 1_n9864 , 1_n9865 , 1_n9867 , 1_n9868 , 1_n9869 , 1_n9870 , 1_n9871 , 1_n9873 , 1_n9874 , 1_n9875 , 1_n9876 , 1_n9877 , 1_n9878 , 1_n9879 , 1_n9880 , 1_n9881 , 1_n9882 , 1_n9883 , 1_n9884 , 1_n9885 , 1_n9886 , 1_n9888 , 1_n9889 , 1_n9890 , 1_n9891 , 1_n9892 , 1_n9893 , 1_n9894 , 1_n9895 , 1_n9896 , 1_n9897 , 1_n9898 , 1_n9899 , 1_n9900 , 1_n9901 , 1_n9902 , 1_n9903 , 1_n9904 , 1_n9905 , 1_n9907 , 1_n9908 , 1_n9909 , 1_n9910 , 1_n9911 , 1_n9912 , 1_n9913 , 1_n9914 , 1_n9916 , 1_n9917 , 1_n9918 , 1_n9919 , 1_n9920 , 1_n9921 , 1_n9922 , 1_n9923 , 1_n9924 , 1_n9925 , 1_n9926 , 1_n9927 , 1_n9928 , 1_n9929 , 1_n9930 , 1_n9931 , 1_n9932 , 1_n9933 , 1_n9934 , 1_n9935 , 1_n9936 , 1_n9937 , 1_n9938 , 1_n9939 , 1_n9940 , 1_n9941 , 1_n9942 , 1_n9943 , 1_n9944 , 1_n9945 , 1_n9946 , 1_n9947 , 1_n9948 , 1_n9949 , 1_n9950 , 1_n9951 , 1_n9952 , 1_n9953 , 1_n9954 , 1_n9955 , 1_n9956 , 1_n9957 , 1_n9958 , 1_n9959 , 1_n9960 , 1_n9961 , 1_n9962 , 1_n9963 , 1_n9964 , 1_n9965 , 1_n9966 , 1_n9967 , 1_n9968 , 1_n9969 , 1_n9970 , 1_n9971 , 1_n9972 , 1_n9973 , 1_n9974 , 1_n9975 , 1_n9976 , 1_n9977 , 1_n9978 , 1_n9979 , 1_n9980 , 1_n9981 , 1_n9982 , 1_n9983 , 1_n9984 , 1_n9985 , 1_n9986 , 1_n9987 , 1_n9988 , 1_n9989 , 1_n9990 , 1_n9991 , 1_n9992 , 1_n9993 , 1_n9994 , 1_n9995 , 1_n9996 , 1_n9997 , 1_n9998 , 1_n9999 , 1_n10000 , 1_n10001 , 1_n10002 , 1_n10003 , 1_n10004 , 1_n10005 , 1_n10006 , 1_n10007 , 1_n10008 , 1_n10009 , 1_n10010 , 1_n10011 , 1_n10012 , 1_n10013 , 1_n10014 , 1_n10015 , 1_n10016 , 1_n10017 , 1_n10018 , 1_n10019 , 1_n10020 , 1_n10021 , 1_n10022 , 1_n10023 , 1_n10024 , 1_n10025 , 1_n10026 , 1_n10027 , 1_n10028 , 1_n10029 , 1_n10030 , 1_n10031 , 1_n10032 , 1_n10033 , 1_n10034 , 1_n10035 , 1_n10036 , 1_n10037 , 1_n10038 , 1_n10039 , 1_n10040 , 1_n10041 , 1_n10042 , 1_n10043 , 1_n10044 , 1_n10045 , 1_n10046 , 1_n10047 , 1_n10048 , 1_n10049 , 1_n10050 , 1_n10051 , 1_n10052 , 1_n10053 , 1_n10054 , 1_n10055 , 1_n10056 , 1_n10057 , 1_n10058 , 1_n10059 , 1_n10060 , 1_n10061 , 1_n10062 , 1_n10064 , 1_n10065 , 1_n10066 , 1_n10067 , 1_n10068 , 1_n10069 , 1_n10070 , 1_n10071 , 1_n10072 , 1_n10073 , 1_n10074 , 1_n10075 , 1_n10076 , 1_n10077 , 1_n10078 , 1_n10079 , 1_n10080 , 1_n10081 , 1_n10082 , 1_n10083 , 1_n10084 , 1_n10085 , 1_n10086 , 1_n10087 , 1_n10088 , 1_n10089 , 1_n10090 , 1_n10091 , 1_n10092 , 1_n10093 , 1_n10094 , 1_n10095 , 1_n10096 , 1_n10097 , 1_n10098 , 1_n10099 , 1_n10100 , 1_n10102 , 1_n10103 , 1_n10104 , 1_n10105 , 1_n10106 , 1_n10107 , 1_n10108 , 1_n10109 , 1_n10110 , 1_n10111 , 1_n10112 , 1_n10114 , 1_n10115 , 1_n10116 , 1_n10117 , 1_n10118 , 1_n10119 , 1_n10120 , 1_n10121 , 1_n10123 , 1_n10124 , 1_n10125 , 1_n10126 , 1_n10127 , 1_n10128 , 1_n10129 , 1_n10130 , 1_n10131 , 1_n10132 , 1_n10133 , 1_n10134 , 1_n10135 , 1_n10136 , 1_n10137 , 1_n10138 , 1_n10139 , 1_n10140 , 1_n10141 , 1_n10143 , 1_n10144 , 1_n10145 , 1_n10146 , 1_n10147 , 1_n10148 , 1_n10149 , 1_n10150 , 1_n10151 , 1_n10152 , 1_n10153 , 1_n10154 , 1_n10155 , 1_n10156 , 1_n10157 , 1_n10158 , 1_n10159 , 1_n10160 , 1_n10161 , 1_n10163 , 1_n10164 , 1_n10165 , 1_n10166 , 1_n10167 , 1_n10169 , 1_n10170 , 1_n10171 , 1_n10172 , 1_n10173 , 1_n10174 , 1_n10175 , 1_n10176 , 1_n10177 , 1_n10178 , 1_n10179 , 1_n10180 , 1_n10181 , 1_n10182 , 1_n10183 , 1_n10184 , 1_n10185 , 1_n10186 , 1_n10187 , 1_n10188 , 1_n10189 , 1_n10190 , 1_n10191 , 1_n10192 , 1_n10193 , 1_n10194 , 1_n10195 , 1_n10196 , 1_n10197 , 1_n10198 , 1_n10199 , 1_n10200 , 1_n10201 , 1_n10202 , 1_n10203 , 1_n10204 , 1_n10205 , 1_n10206 , 1_n10207 , 1_n10208 , 1_n10209 , 1_n10210 , 1_n10211 , 1_n10212 , 1_n10213 , 1_n10214 , 1_n10215 , 1_n10216 , 1_n10217 , 1_n10218 , 1_n10219 , 1_n10220 , 1_n10221 , 1_n10222 , 1_n10223 , 1_n10224 , 1_n10225 , 1_n10226 , 1_n10227 , 1_n10228 , 1_n10229 , 1_n10230 , 1_n10231 , 1_n10232 , 1_n10233 , 1_n10234 , 1_n10235 , 1_n10236 , 1_n10237 , 1_n10238 , 1_n10239 , 1_n10240 , 1_n10241 , 1_n10242 , 1_n10244 , 1_n10245 , 1_n10246 , 1_n10247 , 1_n10248 , 1_n10249 , 1_n10250 , 1_n10251 , 1_n10252 , 1_n10253 , 1_n10254 , 1_n10255 , 1_n10256 , 1_n10257 , 1_n10258 , 1_n10259 , 1_n10260 , 1_n10261 , 1_n10262 , 1_n10263 , 1_n10264 , 1_n10265 , 1_n10266 , 1_n10267 , 1_n10268 , 1_n10269 , 1_n10270 , 1_n10271 , 1_n10272 , 1_n10273 , 1_n10274 , 1_n10275 , 1_n10276 , 1_n10277 , 1_n10278 , 1_n10279 , 1_n10280 , 1_n10281 , 1_n10282 , 1_n10283 , 1_n10284 , 1_n10285 , 1_n10286 , 1_n10287 , 1_n10288 , 1_n10289 , 1_n10290 , 1_n10291 , 1_n10292 , 1_n10293 , 1_n10294 , 1_n10295 , 1_n10296 , 1_n10297 , 1_n10298 , 1_n10299 , 1_n10300 , 1_n10301 , 1_n10302 , 1_n10303 , 1_n10304 , 1_n10305 , 1_n10306 , 1_n10307 , 1_n10308 , 1_n10309 , 1_n10310 , 1_n10311 , 1_n10312 , 1_n10313 , 1_n10314 , 1_n10315 , 1_n10316 , 1_n10317 , 1_n10318 , 1_n10319 , 1_n10320 , 1_n10321 , 1_n10322 , 1_n10323 , 1_n10324 , 1_n10325 , 1_n10326 , 1_n10327 , 1_n10328 , 1_n10329 , 1_n10330 , 1_n10331 , 1_n10332 , 1_n10333 , 1_n10334 , 1_n10335 , 1_n10336 , 1_n10337 , 1_n10338 , 1_n10339 , 1_n10340 , 1_n10341 , 1_n10342 , 1_n10343 , 1_n10344 , 1_n10345 , 1_n10346 , 1_n10347 , 1_n10348 , 1_n10349 , 1_n10350 , 1_n10351 , 1_n10352 , 1_n10353 , 1_n10354 , 1_n10355 , 1_n10356 , 1_n10357 , 1_n10358 , 1_n10359 , 1_n10360 , 1_n10361 , 1_n10362 , 1_n10363 , 1_n10364 , 1_n10365 , 1_n10366 , 1_n10367 , 1_n10368 , 1_n10369 , 1_n10370 , 1_n10371 , 1_n10372 , 1_n10373 , 1_n10374 , 1_n10375 , 1_n10376 , 1_n10377 , 1_n10378 , 1_n10379 , 1_n10380 , 1_n10381 , 1_n10382 , 1_n10383 , 1_n10384 , 1_n10385 , 1_n10386 , 1_n10387 , 1_n10388 , 1_n10389 , 1_n10390 , 1_n10391 , 1_n10392 , 1_n10393 , 1_n10394 , 1_n10395 , 1_n10396 , 1_n10397 , 1_n10398 , 1_n10399 , 1_n10400 , 1_n10401 , 1_n10402 , 1_n10403 , 1_n10404 , 1_n10405 , 1_n10406 , 1_n10407 , 1_n10409 , 1_n10410 , 1_n10411 , 1_n10412 , 1_n10413 , 1_n10414 , 1_n10415 , 1_n10417 , 1_n10418 , 1_n10419 , 1_n10420 , 1_n10421 , 1_n10422 , 1_n10423 , 1_n10424 , 1_n10425 , 1_n10426 , 1_n10427 , 1_n10428 , 1_n10429 , 1_n10430 , 1_n10431 , 1_n10432 , 1_n10433 , 1_n10434 , 1_n10435 , 1_n10436 , 1_n10437 , 1_n10438 , 1_n10439 , 1_n10440 , 1_n10441 , 1_n10442 , 1_n10443 , 1_n10444 , 1_n10445 , 1_n10446 , 1_n10447 , 1_n10448 , 1_n10449 , 1_n10450 , 1_n10452 , 1_n10454 , 1_n10455 , 1_n10456 , 1_n10457 , 1_n10458 , 1_n10459 , 1_n10460 , 1_n10461 , 1_n10462 , 1_n10463 , 1_n10464 , 1_n10465 , 1_n10466 , 1_n10467 , 1_n10468 , 1_n10469 , 1_n10470 , 1_n10471 , 1_n10472 , 1_n10473 , 1_n10474 , 1_n10475 , 1_n10476 , 1_n10477 , 1_n10478 , 1_n10479 , 1_n10480 , 1_n10481 , 1_n10482 , 1_n10483 , 1_n10484 , 1_n10485 , 1_n10486 , 1_n10487 , 1_n10488 , 1_n10489 , 1_n10490 , 1_n10491 , 1_n10492 , 1_n10493 , 1_n10494 , 1_n10495 , 1_n10496 , 1_n10497 , 1_n10498 , 1_n10499 , 1_n10500 , 1_n10501 , 1_n10502 , 1_n10503 , 1_n10504 , 1_n10505 , 1_n10506 , 1_n10507 , 1_n10508 , 1_n10509 , 1_n10510 , 1_n10511 , 1_n10512 , 1_n10513 , 1_n10514 , 1_n10515 , 1_n10516 , 1_n10517 , 1_n10518 , 1_n10519 , 1_n10520 , 1_n10521 , 1_n10523 , 1_n10525 , 1_n10526 , 1_n10527 , 1_n10528 , 1_n10529 , 1_n10530 , 1_n10531 , 1_n10532 , 1_n10533 , 1_n10534 , 1_n10535 , 1_n10536 , 1_n10537 , 1_n10538 , 1_n10539 , 1_n10540 , 1_n10541 , 1_n10542 , 1_n10543 , 1_n10544 , 1_n10545 , 1_n10546 , 1_n10547 , 1_n10548 , 1_n10549 , 1_n10550 , 1_n10551 , 1_n10552 , 1_n10553 , 1_n10554 , 1_n10555 , 1_n10556 , 1_n10557 , 1_n10558 , 1_n10559 , 1_n10561 , 1_n10562 , 1_n10563 , 1_n10564 , 1_n10565 , 1_n10566 , 1_n10567 , 1_n10568 , 1_n10569 , 1_n10570 , 1_n10571 , 1_n10572 , 1_n10573 , 1_n10574 , 1_n10575 , 1_n10576 , 1_n10577 , 1_n10578 , 1_n10579 , 1_n10580 , 1_n10581 , 1_n10582 , 1_n10583 , 1_n10584 , 1_n10585 , 1_n10586 , 1_n10587 , 1_n10588 , 1_n10589 , 1_n10590 , 1_n10591 , 1_n10592 , 1_n10593 , 1_n10595 , 1_n10596 , 1_n10597 , 1_n10598 , 1_n10599 , 1_n10600 , 1_n10601 , 1_n10602 , 1_n10603 , 1_n10604 , 1_n10605 , 1_n10607 , 1_n10608 , 1_n10609 , 1_n10610 , 1_n10611 , 1_n10612 , 1_n10613 , 1_n10614 , 1_n10615 , 1_n10616 , 1_n10617 , 1_n10618 , 1_n10619 , 1_n10620 , 1_n10621 , 1_n10622 , 1_n10623 , 1_n10624 , 1_n10625 , 1_n10626 , 1_n10627 , 1_n10629 , 1_n10630 , 1_n10631 , 1_n10632 , 1_n10633 , 1_n10634 , 1_n10635 , 1_n10636 , 1_n10637 , 1_n10638 , 1_n10639 , 1_n10640 , 1_n10641 , 1_n10643 , 1_n10644 , 1_n10645 , 1_n10646 , 1_n10647 , 1_n10648 , 1_n10649 , 1_n10650 , 1_n10651 , 1_n10652 , 1_n10653 , 1_n10654 , 1_n10655 , 1_n10656 , 1_n10658 , 1_n10659 , 1_n10660 , 1_n10661 , 1_n10662 , 1_n10663 , 1_n10664 , 1_n10665 , 1_n10666 , 1_n10667 , 1_n10668 , 1_n10669 , 1_n10670 , 1_n10671 , 1_n10672 , 1_n10673 , 1_n10674 , 1_n10675 , 1_n10676 , 1_n10677 , 1_n10678 , 1_n10679 , 1_n10680 , 1_n10681 , 1_n10682 , 1_n10683 , 1_n10684 , 1_n10685 , 1_n10686 , 1_n10687 , 1_n10688 , 1_n10689 , 1_n10690 , 1_n10691 , 1_n10692 , 1_n10693 , 1_n10694 , 1_n10695 , 1_n10696 , 1_n10697 , 1_n10698 , 1_n10699 , 1_n10700 , 1_n10701 , 1_n10702 , 1_n10703 , 1_n10704 , 1_n10705 , 1_n10706 , 1_n10707 , 1_n10708 , 1_n10709 , 1_n10710 , 1_n10711 , 1_n10712 , 1_n10713 , 1_n10714 , 1_n10715 , 1_n10716 , 1_n10717 , 1_n10718 , 1_n10719 , 1_n10720 , 1_n10721 , 1_n10722 , 1_n10723 , 1_n10724 , 1_n10725 , 1_n10726 , 1_n10727 , 1_n10728 , 1_n10729 , 1_n10730 , 1_n10731 , 1_n10732 , 1_n10733 , 1_n10734 , 1_n10735 , 1_n10737 , 1_n10738 , 1_n10739 , 1_n10740 , 1_n10741 , 1_n10742 , 1_n10743 , 1_n10744 , 1_n10745 , 1_n10746 , 1_n10747 , 1_n10748 , 1_n10749 , 1_n10750 , 1_n10751 , 1_n10752 , 1_n10753 , 1_n10754 , 1_n10755 , 1_n10756 , 1_n10757 , 1_n10758 , 1_n10759 , 1_n10760 , 1_n10761 , 1_n10762 , 1_n10763 , 1_n10764 , 1_n10765 , 1_n10766 , 1_n10767 , 1_n10768 , 1_n10769 , 1_n10771 , 1_n10772 , 1_n10773 , 1_n10774 , 1_n10775 , 1_n10776 , 1_n10777 , 1_n10778 , 1_n10779 , 1_n10780 , 1_n10781 , 1_n10782 , 1_n10783 , 1_n10784 , 1_n10785 , 1_n10786 , 1_n10787 , 1_n10788 , 1_n10789 , 1_n10790 , 1_n10791 , 1_n10792 , 1_n10793 , 1_n10794 , 1_n10795 , 1_n10796 , 1_n10798 , 1_n10799 , 1_n10800 , 1_n10801 , 1_n10802 , 1_n10803 , 1_n10804 , 1_n10806 , 1_n10807 , 1_n10808 , 1_n10809 , 1_n10810 , 1_n10811 , 1_n10812 , 1_n10813 , 1_n10814 , 1_n10815 , 1_n10816 , 1_n10817 , 1_n10818 , 1_n10819 , 1_n10820 , 1_n10821 , 1_n10822 , 1_n10823 , 1_n10824 , 1_n10825 , 1_n10826 , 1_n10827 , 1_n10828 , 1_n10829 , 1_n10830 , 1_n10831 , 1_n10832 , 1_n10833 , 1_n10834 , 1_n10835 , 1_n10836 , 1_n10837 , 1_n10838 , 1_n10839 , 1_n10840 , 1_n10841 , 1_n10842 , 1_n10843 , 1_n10844 , 1_n10845 , 1_n10846 , 1_n10847 , 1_n10848 , 1_n10849 , 1_n10850 , 1_n10851 , 1_n10852 , 1_n10853 , 1_n10854 , 1_n10855 , 1_n10856 , 1_n10857 , 1_n10858 , 1_n10859 , 1_n10860 , 1_n10861 , 1_n10862 , 1_n10863 , 1_n10864 , 1_n10865 , 1_n10867 , 1_n10868 , 1_n10869 , 1_n10870 , 1_n10871 , 1_n10872 , 1_n10873 , 1_n10875 , 1_n10876 , 1_n10877 , 1_n10878 , 1_n10879 , 1_n10880 , 1_n10881 , 1_n10882 , 1_n10883 , 1_n10884 , 1_n10885 , 1_n10886 , 1_n10887 , 1_n10888 , 1_n10889 , 1_n10890 , 1_n10891 , 1_n10892 , 1_n10893 , 1_n10894 , 1_n10895 , 1_n10896 , 1_n10897 , 1_n10898 , 1_n10899 , 1_n10900 , 1_n10901 , 1_n10902 , 1_n10903 , 1_n10904 , 1_n10905 , 1_n10906 , 1_n10907 , 1_n10909 , 1_n10910 , 1_n10911 , 1_n10912 , 1_n10913 , 1_n10914 , 1_n10915 , 1_n10916 , 1_n10917 , 1_n10918 , 1_n10919 , 1_n10920 , 1_n10921 , 1_n10922 , 1_n10923 , 1_n10924 , 1_n10925 , 1_n10926 , 1_n10927 , 1_n10928 , 1_n10929 , 1_n10930 , 1_n10931 , 1_n10932 , 1_n10933 , 1_n10934 , 1_n10935 , 1_n10936 , 1_n10937 , 1_n10938 , 1_n10939 , 1_n10940 , 1_n10941 , 1_n10942 , 1_n10943 , 1_n10944 , 1_n10945 , 1_n10946 , 1_n10947 , 1_n10948 , 1_n10949 , 1_n10950 , 1_n10951 , 1_n10952 , 1_n10953 , 1_n10954 , 1_n10955 , 1_n10956 , 1_n10957 , 1_n10958 , 1_n10959 , 1_n10960 , 1_n10961 , 1_n10962 , 1_n10963 , 1_n10964 , 1_n10965 , 1_n10966 , 1_n10967 , 1_n10968 , 1_n10969 , 1_n10970 , 1_n10971 , 1_n10972 , 1_n10973 , 1_n10974 , 1_n10975 , 1_n10976 , 1_n10977 , 1_n10978 , 1_n10979 , 1_n10980 , 1_n10981 , 1_n10982 , 1_n10983 , 1_n10984 , 1_n10985 , 1_n10986 , 1_n10987 , 1_n10988 , 1_n10989 , 1_n10990 , 1_n10991 , 1_n10992 , 1_n10993 , 1_n10994 , 1_n10995 , 1_n10996 , 1_n10997 , 1_n10998 , 1_n10999 , 1_n11000 , 1_n11001 , 1_n11002 , 1_n11003 , 1_n11004 , 1_n11005 , 1_n11006 , 1_n11007 , 1_n11008 , 1_n11009 , 1_n11010 , 1_n11011 , 1_n11012 , 1_n11013 , 1_n11014 , 1_n11015 , 1_n11016 , 1_n11017 , 1_n11018 , 1_n11019 , 1_n11020 , 1_n11021 , 1_n11022 , 1_n11023 , 1_n11024 , 1_n11025 , 1_n11026 , 1_n11027 , 1_n11028 , 1_n11029 , 1_n11031 , 1_n11032 , 1_n11033 , 1_n11034 , 1_n11035 , 1_n11036 , 1_n11037 , 1_n11038 , 1_n11039 , 1_n11040 , 1_n11041 , 1_n11042 , 1_n11043 , 1_n11044 , 1_n11045 , 1_n11046 , 1_n11047 , 1_n11048 , 1_n11049 , 1_n11050 , 1_n11051 , 1_n11052 , 1_n11053 , 1_n11054 , 1_n11055 , 1_n11056 , 1_n11059 , 1_n11060 , 1_n11062 , 1_n11063 , 1_n11064 , 1_n11065 , 1_n11066 , 1_n11067 , 1_n11068 , 1_n11069 , 1_n11070 , 1_n11071 , 1_n11072 , 1_n11073 , 1_n11074 , 1_n11075 , 1_n11076 , 1_n11078 , 1_n11079 , 1_n11080 , 1_n11081 , 1_n11082 , 1_n11083 , 1_n11084 , 1_n11085 , 1_n11086 , 1_n11087 , 1_n11088 , 1_n11089 , 1_n11090 , 1_n11091 , 1_n11092 , 1_n11093 , 1_n11094 , 1_n11095 , 1_n11096 , 1_n11097 , 1_n11098 , 1_n11099 , 1_n11100 , 1_n11101 , 1_n11102 , 1_n11103 , 1_n11104 , 1_n11105 , 1_n11106 , 1_n11107 , 1_n11108 , 1_n11110 , 1_n11112 , 1_n11113 , 1_n11114 , 1_n11115 , 1_n11116 , 1_n11117 , 1_n11118 , 1_n11119 , 1_n11120 , 1_n11121 , 1_n11122 , 1_n11123 , 1_n11124 , 1_n11125 , 1_n11126 , 1_n11127 , 1_n11128 , 1_n11129 , 1_n11130 , 1_n11131 , 1_n11132 , 1_n11133 , 1_n11134 , 1_n11135 , 1_n11136 , 1_n11137 , 1_n11138 , 1_n11139 , 1_n11141 , 1_n11142 , 1_n11143 , 1_n11144 , 1_n11145 , 1_n11146 , 1_n11148 , 1_n11149 , 1_n11150 , 1_n11151 , 1_n11152 , 1_n11153 , 1_n11154 , 1_n11155 , 1_n11156 , 1_n11157 , 1_n11158 , 1_n11159 , 1_n11160 , 1_n11161 , 1_n11162 , 1_n11163 , 1_n11164 , 1_n11165 , 1_n11166 , 1_n11167 , 1_n11168 , 1_n11169 , 1_n11170 , 1_n11171 , 1_n11172 , 1_n11173 , 1_n11174 , 1_n11175 , 1_n11176 , 1_n11177 , 1_n11178 , 1_n11179 , 1_n11181 , 1_n11182 , 1_n11183 , 1_n11184 , 1_n11185 , 1_n11186 , 1_n11187 , 1_n11188 , 1_n11189 , 1_n11190 , 1_n11191 , 1_n11192 , 1_n11193 , 1_n11194 , 1_n11195 , 1_n11196 , 1_n11197 , 1_n11198 , 1_n11199 , 1_n11200 , 1_n11201 , 1_n11202 , 1_n11203 , 1_n11204 , 1_n11205 , 1_n11206 , 1_n11207 , 1_n11208 , 1_n11209 , 1_n11210 , 1_n11211 , 1_n11212 , 1_n11213 , 1_n11214 , 1_n11215 , 1_n11216 , 1_n11217 , 1_n11218 , 1_n11219 , 1_n11220 , 1_n11221 , 1_n11223 , 1_n11224 , 1_n11225 , 1_n11226 , 1_n11227 , 1_n11228 , 1_n11229 , 1_n11230 , 1_n11231 , 1_n11232 , 1_n11233 , 1_n11234 , 1_n11235 , 1_n11237 , 1_n11238 , 1_n11239 , 1_n11240 , 1_n11241 , 1_n11242 , 1_n11243 , 1_n11244 , 1_n11245 , 1_n11246 , 1_n11247 , 1_n11248 , 1_n11249 , 1_n11250 , 1_n11251 , 1_n11253 , 1_n11254 , 1_n11255 , 1_n11256 , 1_n11257 , 1_n11258 , 1_n11259 , 1_n11260 , 1_n11261 , 1_n11262 , 1_n11263 , 1_n11265 , 1_n11266 , 1_n11267 , 1_n11268 , 1_n11269 , 1_n11270 , 1_n11271 , 1_n11272 , 1_n11273 , 1_n11274 , 1_n11275 , 1_n11276 , 1_n11277 , 1_n11278 , 1_n11279 , 1_n11280 , 1_n11281 , 1_n11282 , 1_n11283 , 1_n11284 , 1_n11285 , 1_n11286 , 1_n11287 , 1_n11288 , 1_n11289 , 1_n11290 , 1_n11291 , 1_n11292 , 1_n11293 , 1_n11294 , 1_n11295 , 1_n11296 , 1_n11297 , 1_n11298 , 1_n11299 , 1_n11300 , 1_n11301 , 1_n11302 , 1_n11303 , 1_n11304 , 1_n11305 , 1_n11306 , 1_n11307 , 1_n11308 , 1_n11309 , 1_n11310 , 1_n11311 , 1_n11312 , 1_n11313 , 1_n11314 , 1_n11315 , 1_n11316 , 1_n11317 , 1_n11318 , 1_n11319 , 1_n11320 , 1_n11321 , 1_n11322 , 1_n11323 , 1_n11325 , 1_n11326 , 1_n11327 , 1_n11328 , 1_n11329 , 1_n11330 , 1_n11331 , 1_n11332 , 1_n11333 , 1_n11334 , 1_n11335 , 1_n11336 , 1_n11337 , 1_n11338 , 1_n11339 , 1_n11340 , 1_n11341 , 1_n11342 , 1_n11343 , 1_n11344 , 1_n11345 , 1_n11346 , 1_n11347 , 1_n11348 , 1_n11349 , 1_n11351 , 1_n11352 , 1_n11353 , 1_n11354 , 1_n11355 , 1_n11356 , 1_n11357 , 1_n11358 , 1_n11359 , 1_n11360 , 1_n11361 , 1_n11362 , 1_n11363 , 1_n11364 , 1_n11365 , 1_n11366 , 1_n11367 , 1_n11368 , 1_n11369 , 1_n11370 , 1_n11371 , 1_n11372 , 1_n11373 , 1_n11374 , 1_n11375 , 1_n11376 , 1_n11377 , 1_n11378 , 1_n11379 , 1_n11380 , 1_n11381 , 1_n11382 , 1_n11383 , 1_n11384 , 1_n11385 , 1_n11386 , 1_n11387 , 1_n11388 , 1_n11389 , 1_n11390 , 1_n11391 , 1_n11392 , 1_n11393 , 1_n11394 , 1_n11395 , 1_n11397 , 1_n11398 , 1_n11399 , 1_n11400 , 1_n11401 , 1_n11402 , 1_n11403 , 1_n11404 , 1_n11405 , 1_n11406 , 1_n11407 , 1_n11408 , 1_n11409 , 1_n11410 , 1_n11412 , 1_n11413 , 1_n11414 , 1_n11415 , 1_n11416 , 1_n11417 , 1_n11418 , 1_n11419 , 1_n11420 , 1_n11421 , 1_n11422 , 1_n11423 , 1_n11424 , 1_n11425 , 1_n11426 , 1_n11427 , 1_n11428 , 1_n11430 , 1_n11431 , 1_n11432 , 1_n11433 , 1_n11434 , 1_n11435 , 1_n11436 , 1_n11437 , 1_n11438 , 1_n11439 , 1_n11440 , 1_n11441 , 1_n11442 , 1_n11443 , 1_n11444 , 1_n11445 , 1_n11446 , 1_n11447 , 1_n11448 , 1_n11449 , 1_n11450 , 1_n11451 , 1_n11452 , 1_n11453 , 1_n11454 , 1_n11455 , 1_n11456 , 1_n11457 , 1_n11458 , 1_n11459 , 1_n11460 , 1_n11461 , 1_n11462 , 1_n11463 , 1_n11464 , 1_n11465 , 1_n11466 , 1_n11467 , 1_n11468 , 1_n11469 , 1_n11470 , 1_n11471 , 1_n11472 , 1_n11473 , 1_n11474 , 1_n11475 , 1_n11476 , 1_n11477 , 1_n11478 , 1_n11479 , 1_n11480 , 1_n11481 , 1_n11482 , 1_n11483 , 1_n11485 , 1_n11486 , 1_n11487 , 1_n11489 , 1_n11490 , 1_n11491 , 1_n11492 , 1_n11493 , 1_n11494 , 1_n11495 , 1_n11496 , 1_n11497 , 1_n11498 , 1_n11499 , 1_n11500 , 1_n11501 , 1_n11502 , 1_n11503 , 1_n11504 , 1_n11505 , 1_n11506 , 1_n11507 , 1_n11508 , 1_n11509 , 1_n11510 , 1_n11511 , 1_n11512 , 1_n11513 , 1_n11514 , 1_n11515 , 1_n11516 , 1_n11517 , 1_n11518 , 1_n11519 , 1_n11520 , 1_n11521 , 1_n11522 , 1_n11523 , 1_n11524 , 1_n11525 , 1_n11526 , 1_n11527 , 1_n11528 , 1_n11529 , 1_n11530 , 1_n11531 , 1_n11532 , 1_n11533 , 1_n11534 , 1_n11535 , 1_n11536 , 1_n11538 , 1_n11539 , 1_n11540 , 1_n11541 , 1_n11542 , 1_n11543 , 1_n11544 , 1_n11545 , 1_n11546 , 1_n11547 , 1_n11548 , 1_n11549 , 1_n11550 , 1_n11551 , 1_n11552 , 1_n11553 , 1_n11554 , 1_n11555 , 1_n11556 , 1_n11557 , 1_n11558 , 1_n11559 , 1_n11560 , 1_n11561 , 1_n11562 , 1_n11563 , 1_n11564 , 1_n11565 , 1_n11566 , 1_n11567 , 1_n11568 , 1_n11569 , 1_n11570 , 1_n11571 , 1_n11572 , 1_n11573 , 1_n11575 , 1_n11576 , 1_n11577 , 1_n11578 , 1_n11579 , 1_n11580 , 1_n11581 , 1_n11582 , 1_n11583 , 1_n11584 , 1_n11585 , 1_n11586 , 1_n11587 , 1_n11588 , 1_n11589 , 1_n11590 , 1_n11591 , 1_n11592 , 1_n11593 , 1_n11594 , 1_n11595 , 1_n11596 , 1_n11597 , 1_n11598 , 1_n11599 , 1_n11600 , 1_n11601 , 1_n11602 , 1_n11603 , 1_n11604 , 1_n11605 , 1_n11606 , 1_n11607 , 1_n11608 , 1_n11609 , 1_n11610 , 1_n11611 , 1_n11612 , 1_n11613 , 1_n11614 , 1_n11615 , 1_n11616 , 1_n11617 , 1_n11618 , 1_n11619 , 1_n11620 , 1_n11621 , 1_n11622 , 1_n11623 , 1_n11624 , 1_n11625 , 1_n11626 , 1_n11627 , 1_n11628 , 1_n11629 , 1_n11630 , 1_n11631 , 1_n11632 , 1_n11633 , 1_n11635 , 1_n11636 , 1_n11637 , 1_n11638 , 1_n11639 , 1_n11640 , 1_n11641 , 1_n11642 , 1_n11643 , 1_n11644 , 1_n11645 , 1_n11646 , 1_n11647 , 1_n11648 , 1_n11649 , 1_n11650 , 1_n11651 , 1_n11652 , 1_n11653 , 1_n11654 , 1_n11655 , 1_n11656 , 1_n11657 , 1_n11658 , 1_n11659 , 1_n11660 , 1_n11661 , 1_n11662 , 1_n11663 , 1_n11664 , 1_n11666 , 1_n11668 , 1_n11669 , 1_n11670 , 1_n11671 , 1_n11672 , 1_n11673 , 1_n11674 , 1_n11675 , 1_n11676 , 1_n11677 , 1_n11678 , 1_n11679 , 1_n11680 , 1_n11681 , 1_n11682 , 1_n11683 , 1_n11684 , 1_n11685 , 1_n11686 , 1_n11687 , 1_n11688 , 1_n11689 , 1_n11690 , 1_n11691 , 1_n11692 , 1_n11693 , 1_n11694 , 1_n11695 , 1_n11696 , 1_n11697 , 1_n11698 , 1_n11699 , 1_n11700 , 1_n11701 , 1_n11702 , 1_n11703 , 1_n11704 , 1_n11705 , 1_n11706 , 1_n11707 , 1_n11708 , 1_n11709 , 1_n11710 , 1_n11711 , 1_n11712 , 1_n11713 , 1_n11714 , 1_n11715 , 1_n11716 , 1_n11717 , 1_n11718 , 1_n11719 , 1_n11720 , 1_n11721 , 1_n11722 , 1_n11723 , 1_n11724 , 1_n11725 , 1_n11726 , 1_n11727 , 1_n11728 , 1_n11729 , 1_n11730 , 1_n11731 , 1_n11733 , 1_n11735 , 1_n11736 , 1_n11737 , 1_n11738 , 1_n11739 , 1_n11740 , 1_n11741 , 1_n11742 , 1_n11743 , 1_n11744 , 1_n11745 , 1_n11746 , 1_n11747 , 1_n11748 , 1_n11749 , 1_n11750 , 1_n11751 , 1_n11752 , 1_n11753 , 1_n11754 , 1_n11755 , 1_n11756 , 1_n11757 , 1_n11758 , 1_n11759 , 1_n11760 , 1_n11761 , 1_n11762 , 1_n11763 , 1_n11764 , 1_n11765 , 1_n11766 , 1_n11767 , 1_n11768 , 1_n11769 , 1_n11770 , 1_n11771 , 1_n11772 , 1_n11773 , 1_n11774 , 1_n11775 , 1_n11776 , 1_n11777 , 1_n11779 , 1_n11780 , 1_n11781 , 1_n11782 , 1_n11783 , 1_n11784 , 1_n11785 , 1_n11786 , 1_n11787 , 1_n11788 , 1_n11789 , 1_n11790 , 1_n11791 , 1_n11793 , 1_n11794 , 1_n11795 , 1_n11796 , 1_n11797 , 1_n11798 , 1_n11799 , 1_n11800 , 1_n11801 , 1_n11802 , 1_n11803 , 1_n11804 , 1_n11805 , 1_n11806 , 1_n11807 , 1_n11808 , 1_n11809 , 1_n11810 , 1_n11811 , 1_n11812 , 1_n11813 , 1_n11814 , 1_n11815 , 1_n11816 , 1_n11817 , 1_n11818 , 1_n11819 , 1_n11820 , 1_n11821 , 1_n11822 , 1_n11823 , 1_n11824 , 1_n11825 , 1_n11826 , 1_n11827 , 1_n11828 , 1_n11829 , 1_n11830 , 1_n11831 , 1_n11832 , 1_n11833 , 1_n11834 , 1_n11836 , 1_n11837 , 1_n11838 , 1_n11839 , 1_n11840 , 1_n11841 , 1_n11842 , 1_n11843 , 1_n11844 , 1_n11845 , 1_n11846 , 1_n11847 , 1_n11848 , 1_n11849 , 1_n11850 , 1_n11851 , 1_n11852 , 1_n11853 , 1_n11854 , 1_n11855 , 1_n11856 , 1_n11857 , 1_n11858 , 1_n11859 , 1_n11860 , 1_n11861 , 1_n11862 , 1_n11863 , 1_n11864 , 1_n11865 , 1_n11866 , 1_n11867 , 1_n11868 , 1_n11869 , 1_n11870 , 1_n11871 , 1_n11872 , 1_n11873 , 1_n11874 , 1_n11875 , 1_n11876 , 1_n11877 , 1_n11878 , 1_n11880 , 1_n11881 , 1_n11883 , 1_n11884 , 1_n11885 , 1_n11886 , 1_n11887 , 1_n11888 , 1_n11889 , 1_n11890 , 1_n11892 , 1_n11893 , 1_n11894 , 1_n11896 , 1_n11897 , 1_n11898 , 1_n11899 , 1_n11900 , 1_n11901 , 1_n11902 , 1_n11903 , 1_n11904 , 1_n11905 , 1_n11906 , 1_n11907 , 1_n11908 , 1_n11909 , 1_n11910 , 1_n11911 , 1_n11912 , 1_n11913 , 1_n11914 , 1_n11915 , 1_n11916 , 1_n11917 , 1_n11918 , 1_n11919 , 1_n11920 , 1_n11921 , 1_n11922 , 1_n11923 , 1_n11924 , 1_n11925 , 1_n11926 , 1_n11927 , 1_n11928 , 1_n11929 , 1_n11930 , 1_n11931 , 1_n11932 , 1_n11933 , 1_n11934 , 1_n11935 , 1_n11936 , 1_n11937 , 1_n11938 , 1_n11939 , 1_n11940 , 1_n11941 , 1_n11942 , 1_n11943 , 1_n11944 , 1_n11945 , 1_n11946 , 1_n11947 , 1_n11948 , 1_n11949 , 1_n11950 , 1_n11951 , 1_n11952 , 1_n11953 , 1_n11954 , 1_n11955 , 1_n11956 , 1_n11957 , 1_n11958 , 1_n11959 , 1_n11960 , 1_n11961 , 1_n11962 , 1_n11963 , 1_n11964 , 1_n11965 , 1_n11966 , 1_n11967 , 1_n11968 , 1_n11969 , 1_n11970 , 1_n11971 , 1_n11972 , 1_n11973 , 1_n11974 , 1_n11975 , 1_n11976 , 1_n11977 , 1_n11978 , 1_n11979 , 1_n11980 , 1_n11981 , 1_n11982 , 1_n11983 , 1_n11984 , 1_n11985 , 1_n11986 , 1_n11987 , 1_n11988 , 1_n11989 , 1_n11990 , 1_n11991 , 1_n11992 , 1_n11993 , 1_n11994 , 1_n11995 , 1_n11996 , 1_n11997 , 1_n11998 , 1_n11999 , 1_n12000 , 1_n12001 , 1_n12002 , 1_n12004 , 1_n12005 , 1_n12006 , 1_n12007 , 1_n12008 , 1_n12009 , 1_n12010 , 1_n12011 , 1_n12012 , 1_n12013 , 1_n12014 , 1_n12015 , 1_n12016 , 1_n12017 , 1_n12018 , 1_n12019 , 1_n12020 , 1_n12021 , 1_n12022 , 1_n12023 , 1_n12024 , 1_n12025 , 1_n12026 , 1_n12027 , 1_n12028 , 1_n12029 , 1_n12030 , 1_n12031 , 1_n12032 , 1_n12033 , 1_n12034 , 1_n12035 , 1_n12036 , 1_n12037 , 1_n12038 , 1_n12039 , 1_n12040 , 1_n12041 , 1_n12042 , 1_n12043 , 1_n12044 , 1_n12045 , 1_n12046 , 1_n12047 , 1_n12048 , 1_n12049 , 1_n12050 , 1_n12051 , 1_n12052 , 1_n12053 , 1_n12054 , 1_n12055 , 1_n12056 , 1_n12057 , 1_n12058 , 1_n12060 , 1_n12061 , 1_n12062 , 1_n12063 , 1_n12064 , 1_n12066 , 1_n12068 , 1_n12069 , 1_n12070 , 1_n12071 , 1_n12072 , 1_n12073 , 1_n12074 , 1_n12075 , 1_n12076 , 1_n12077 , 1_n12078 , 1_n12079 , 1_n12080 , 1_n12081 , 1_n12082 , 1_n12083 , 1_n12084 , 1_n12085 , 1_n12086 , 1_n12087 , 1_n12088 , 1_n12089 , 1_n12090 , 1_n12091 , 1_n12092 , 1_n12093 , 1_n12094 , 1_n12095 , 1_n12096 , 1_n12097 , 1_n12098 , 1_n12099 , 1_n12100 , 1_n12101 , 1_n12102 , 1_n12103 , 1_n12104 , 1_n12105 , 1_n12106 , 1_n12107 , 1_n12108 , 1_n12109 , 1_n12110 , 1_n12111 , 1_n12112 , 1_n12113 , 1_n12114 , 1_n12115 , 1_n12116 , 1_n12117 , 1_n12118 , 1_n12119 , 1_n12120 , 1_n12121 , 1_n12122 , 1_n12123 , 1_n12124 , 1_n12125 , 1_n12126 , 1_n12127 , 1_n12128 , 1_n12129 , 1_n12130 , 1_n12131 , 1_n12132 , 1_n12133 , 1_n12134 , 1_n12135 , 1_n12136 , 1_n12137 , 1_n12138 , 1_n12139 , 1_n12140 , 1_n12141 , 1_n12142 , 1_n12143 , 1_n12144 , 1_n12145 , 1_n12146 , 1_n12147 , 1_n12148 , 1_n12149 , 1_n12150 , 1_n12151 , 1_n12152 , 1_n12153 , 1_n12154 , 1_n12155 , 1_n12156 , 1_n12157 , 1_n12158 , 1_n12159 , 1_n12160 , 1_n12161 , 1_n12162 , 1_n12163 , 1_n12164 , 1_n12165 , 1_n12166 , 1_n12167 , 1_n12168 , 1_n12169 , 1_n12170 , 1_n12171 , 1_n12172 , 1_n12173 , 1_n12174 , 1_n12175 , 1_n12176 , 1_n12177 , 1_n12178 , 1_n12179 , 1_n12180 , 1_n12181 , 1_n12182 , 1_n12183 , 1_n12184 , 1_n12185 , 1_n12186 , 1_n12188 , 1_n12189 , 1_n12190 , 1_n12191 , 1_n12192 , 1_n12193 , 1_n12194 , 1_n12195 , 1_n12196 , 1_n12197 , 1_n12198 , 1_n12199 , 1_n12200 , 1_n12201 , 1_n12202 , 1_n12203 , 1_n12204 , 1_n12205 , 1_n12206 , 1_n12207 , 1_n12208 , 1_n12209 , 1_n12210 , 1_n12211 , 1_n12212 , 1_n12213 , 1_n12214 , 1_n12215 , 1_n12216 , 1_n12217 , 1_n12218 , 1_n12219 , 1_n12220 , 1_n12221 , 1_n12222 , 1_n12223 , 1_n12224 , 1_n12225 , 1_n12226 , 1_n12227 , 1_n12228 , 1_n12229 , 1_n12230 , 1_n12231 , 1_n12232 , 1_n12233 , 1_n12234 , 1_n12235 , 1_n12236 , 1_n12237 , 1_n12238 , 1_n12239 , 1_n12240 , 1_n12241 , 1_n12242 , 1_n12243 , 1_n12244 , 1_n12245 , 1_n12246 , 1_n12247 , 1_n12248 , 1_n12249 , 1_n12250 , 1_n12251 , 1_n12252 , 1_n12253 , 1_n12254 , 1_n12255 , 1_n12256 , 1_n12257 , 1_n12258 , 1_n12259 , 1_n12260 , 1_n12261 , 1_n12262 , 1_n12264 , 1_n12265 , 1_n12266 , 1_n12267 , 1_n12268 , 1_n12269 , 1_n12270 , 1_n12271 , 1_n12272 , 1_n12273 , 1_n12274 , 1_n12275 , 1_n12276 , 1_n12277 , 1_n12278 , 1_n12279 , 1_n12280 , 1_n12281 , 1_n12282 , 1_n12283 , 1_n12285 , 1_n12286 , 1_n12287 , 1_n12288 , 1_n12290 , 1_n12291 , 1_n12292 , 1_n12293 , 1_n12294 , 1_n12295 , 1_n12296 , 1_n12297 , 1_n12298 , 1_n12299 , 1_n12300 , 1_n12301 , 1_n12302 , 1_n12303 , 1_n12304 , 1_n12305 , 1_n12307 , 1_n12308 , 1_n12309 , 1_n12310 , 1_n12311 , 1_n12312 , 1_n12313 , 1_n12314 , 1_n12315 , 1_n12316 , 1_n12317 , 1_n12318 , 1_n12319 , 1_n12320 , 1_n12321 , 1_n12322 , 1_n12323 , 1_n12324 , 1_n12325 , 1_n12326 , 1_n12327 , 1_n12328 , 1_n12329 , 1_n12330 , 1_n12331 , 1_n12332 , 1_n12333 , 1_n12335 , 1_n12336 , 1_n12337 , 1_n12338 , 1_n12339 , 1_n12340 , 1_n12341 , 1_n12342 , 1_n12343 , 1_n12344 , 1_n12345 , 1_n12346 , 1_n12347 , 1_n12349 , 1_n12350 , 1_n12351 , 1_n12353 , 1_n12354 , 1_n12355 , 1_n12356 , 1_n12357 , 1_n12358 , 1_n12359 , 1_n12360 , 1_n12361 , 1_n12362 , 1_n12363 , 1_n12364 , 1_n12365 , 1_n12366 , 1_n12367 , 1_n12368 , 1_n12369 , 1_n12370 , 1_n12371 , 1_n12373 , 1_n12374 , 1_n12375 , 1_n12376 , 1_n12377 , 1_n12378 , 1_n12379 , 1_n12380 , 1_n12381 , 1_n12382 , 1_n12383 , 1_n12384 , 1_n12385 , 1_n12386 , 1_n12387 , 1_n12388 , 1_n12389 , 1_n12390 , 1_n12391 , 1_n12392 , 1_n12393 , 1_n12394 , 1_n12395 , 1_n12396 , 1_n12397 , 1_n12398 , 1_n12399 , 1_n12400 , 1_n12401 , 1_n12402 , 1_n12403 , 1_n12404 , 1_n12405 , 1_n12407 , 1_n12409 , 1_n12410 , 1_n12411 , 1_n12412 , 1_n12413 , 1_n12414 , 1_n12415 , 1_n12416 , 1_n12417 , 1_n12418 , 1_n12419 , 1_n12420 , 1_n12421 , 1_n12422 , 1_n12423 , 1_n12424 , 1_n12425 , 1_n12426 , 1_n12427 , 1_n12428 , 1_n12429 , 1_n12430 , 1_n12431 , 1_n12432 , 1_n12433 , 1_n12434 , 1_n12435 , 1_n12436 , 1_n12437 , 1_n12438 , 1_n12439 , 1_n12440 , 1_n12441 , 1_n12442 , 1_n12443 , 1_n12444 , 1_n12445 , 1_n12446 , 1_n12447 , 1_n12448 , 1_n12449 , 1_n12450 , 1_n12451 , 1_n12452 , 1_n12453 , 1_n12454 , 1_n12455 , 1_n12456 , 1_n12457 , 1_n12458 , 1_n12459 , 1_n12460 , 1_n12461 , 1_n12462 , 1_n12464 , 1_n12465 , 1_n12466 , 1_n12467 , 1_n12468 , 1_n12469 , 1_n12470 , 1_n12471 , 1_n12472 , 1_n12473 , 1_n12474 , 1_n12475 , 1_n12476 , 1_n12477 , 1_n12478 , 1_n12479 , 1_n12480 , 1_n12481 , 1_n12483 , 1_n12484 , 1_n12485 , 1_n12486 , 1_n12487 , 1_n12488 , 1_n12489 , 1_n12490 , 1_n12491 , 1_n12492 , 1_n12493 , 1_n12494 , 1_n12495 , 1_n12496 , 1_n12497 , 1_n12498 , 1_n12499 , 1_n12500 , 1_n12501 , 1_n12502 , 1_n12504 , 1_n12505 , 1_n12506 , 1_n12507 , 1_n12508 , 1_n12509 , 1_n12510 , 1_n12511 , 1_n12512 , 1_n12513 , 1_n12514 , 1_n12516 , 1_n12517 , 1_n12518 , 1_n12519 , 1_n12520 , 1_n12521 , 1_n12522 , 1_n12523 , 1_n12524 , 1_n12525 , 1_n12526 , 1_n12527 , 1_n12528 , 1_n12529 , 1_n12530 , 1_n12531 , 1_n12532 , 1_n12533 , 1_n12534 , 1_n12535 , 1_n12536 , 1_n12537 , 1_n12538 , 1_n12539 , 1_n12540 , 1_n12541 , 1_n12542 , 1_n12543 , 1_n12544 , 1_n12545 , 1_n12546 , 1_n12547 , 1_n12548 , 1_n12549 , 1_n12550 , 1_n12551 , 1_n12552 , 1_n12553 , 1_n12554 , 1_n12555 , 1_n12556 , 1_n12557 , 1_n12558 , 1_n12559 , 1_n12560 , 1_n12561 , 1_n12562 , 1_n12563 , 1_n12564 , 1_n12565 , 1_n12566 , 1_n12567 , 1_n12568 , 1_n12569 , 1_n12570 , 1_n12571 , 1_n12572 , 1_n12573 , 1_n12574 , 1_n12575 , 1_n12576 , 1_n12577 , 1_n12578 , 1_n12580 , 1_n12581 , 1_n12582 , 1_n12583 , 1_n12584 , 1_n12585 , 1_n12586 , 1_n12587 , 1_n12588 , 1_n12589 , 1_n12590 , 1_n12591 , 1_n12593 , 1_n12594 , 1_n12595 , 1_n12596 , 1_n12597 , 1_n12598 , 1_n12599 , 1_n12600 , 1_n12601 , 1_n12602 , 1_n12603 , 1_n12604 , 1_n12606 , 1_n12607 , 1_n12608 , 1_n12609 , 1_n12610 , 1_n12611 , 1_n12612 , 1_n12613 , 1_n12614 , 1_n12615 , 1_n12617 , 1_n12618 , 1_n12619 , 1_n12620 , 1_n12621 , 1_n12622 , 1_n12623 , 1_n12624 , 1_n12625 , 1_n12626 , 1_n12627 , 1_n12628 , 1_n12629 , 1_n12630 , 1_n12631 , 1_n12632 , 1_n12633 , 1_n12634 , 1_n12635 , 1_n12636 , 1_n12637 , 1_n12638 , 1_n12639 , 1_n12640 , 1_n12641 , 1_n12642 , 1_n12643 , 1_n12644 , 1_n12645 , 1_n12646 , 1_n12647 , 1_n12648 , 1_n12649 , 1_n12650 , 1_n12652 , 1_n12653 , 1_n12654 , 1_n12655 , 1_n12656 , 1_n12657 , 1_n12658 , 1_n12659 , 1_n12660 , 1_n12661 , 1_n12662 , 1_n12663 , 1_n12664 , 1_n12665 , 1_n12666 , 1_n12667 , 1_n12668 , 1_n12669 , 1_n12670 , 1_n12671 , 1_n12672 , 1_n12673 , 1_n12674 , 1_n12675 , 1_n12676 , 1_n12677 , 1_n12678 , 1_n12679 , 1_n12680 , 1_n12681 , 1_n12682 , 1_n12683 , 1_n12684 , 1_n12685 , 1_n12686 , 1_n12687 , 1_n12688 , 1_n12689 , 1_n12690 , 1_n12691 , 1_n12692 , 1_n12694 , 1_n12695 , 1_n12696 , 1_n12697 , 1_n12698 , 1_n12699 , 1_n12700 , 1_n12701 , 1_n12702 , 1_n12703 , 1_n12704 , 1_n12705 , 1_n12706 , 1_n12707 , 1_n12708 , 1_n12709 , 1_n12710 , 1_n12711 , 1_n12712 , 1_n12713 , 1_n12714 , 1_n12715 , 1_n12716 , 1_n12717 , 1_n12718 , 1_n12719 , 1_n12720 , 1_n12721 , 1_n12722 , 1_n12723 , 1_n12724 , 1_n12725 , 1_n12726 , 1_n12727 , 1_n12728 , 1_n12729 , 1_n12730 , 1_n12731 , 1_n12732 , 1_n12733 , 1_n12734 , 1_n12735 , 1_n12736 , 1_n12737 , 1_n12738 , 1_n12739 , 1_n12740 , 1_n12741 , 1_n12742 , 1_n12743 , 1_n12744 , 1_n12745 , 1_n12746 , 1_n12747 , 1_n12748 , 1_n12749 , 1_n12751 , 1_n12752 , 1_n12753 , 1_n12754 , 1_n12755 , 1_n12756 , 1_n12757 , 1_n12758 , 1_n12759 , 1_n12760 , 1_n12761 , 1_n12762 , 1_n12763 , 1_n12764 , 1_n12765 , 1_n12766 , 1_n12767 , 1_n12768 , 1_n12769 , 1_n12770 , 1_n12771 , 1_n12772 , 1_n12773 , 1_n12774 , 1_n12775 , 1_n12776 , 1_n12777 , 1_n12778 , 1_n12779 , 1_n12780 , 1_n12781 , 1_n12782 , 1_n12783 , 1_n12784 , 1_n12785 , 1_n12786 , 1_n12787 , 1_n12788 , 1_n12789 , 1_n12790 , 1_n12791 , 1_n12792 , 1_n12793 , 1_n12794 , 1_n12795 , 1_n12796 , 1_n12797 , 1_n12798 , 1_n12799 , 1_n12800 , 1_n12801 , 1_n12802 , 1_n12803 , 1_n12804 , 1_n12805 , 1_n12806 , 1_n12807 , 1_n12808 , 1_n12809 , 1_n12810 , 1_n12811 , 1_n12812 , 1_n12813 , 1_n12814 , 1_n12815 , 1_n12816 , 1_n12817 , 1_n12818 , 1_n12819 , 1_n12820 , 1_n12821 , 1_n12822 , 1_n12823 , 1_n12824 , 1_n12825 , 1_n12826 , 1_n12827 , 1_n12828 , 1_n12829 , 1_n12830 , 1_n12831 , 1_n12832 , 1_n12833 , 1_n12834 , 1_n12835 , 1_n12836 , 1_n12837 , 1_n12838 , 1_n12840 , 1_n12841 , 1_n12842 , 1_n12843 , 1_n12844 , 1_n12845 , 1_n12846 , 1_n12847 , 1_n12848 , 1_n12849 , 1_n12850 , 1_n12851 , 1_n12852 , 1_n12854 , 1_n12855 , 1_n12856 , 1_n12857 , 1_n12858 , 1_n12859 , 1_n12860 , 1_n12861 , 1_n12862 , 1_n12863 , 1_n12864 , 1_n12865 , 1_n12866 , 1_n12867 , 1_n12868 , 1_n12869 , 1_n12870 , 1_n12871 , 1_n12872 , 1_n12873 , 1_n12874 , 1_n12875 , 1_n12876 , 1_n12877 , 1_n12878 , 1_n12879 , 1_n12880 , 1_n12881 , 1_n12882 , 1_n12883 , 1_n12884 , 1_n12885 , 1_n12886 , 1_n12887 , 1_n12888 , 1_n12889 , 1_n12890 , 1_n12891 , 1_n12892 , 1_n12893 , 1_n12894 , 1_n12895 , 1_n12896 , 1_n12897 , 1_n12898 , 1_n12899 , 1_n12900 , 1_n12901 , 1_n12902 , 1_n12903 , 1_n12904 , 1_n12905 , 1_n12906 , 1_n12907 , 1_n12908 , 1_n12909 , 1_n12910 , 1_n12911 , 1_n12913 , 1_n12914 , 1_n12915 , 1_n12916 , 1_n12917 , 1_n12918 , 1_n12919 , 1_n12920 , 1_n12921 , 1_n12922 , 1_n12923 , 1_n12924 , 1_n12925 , 1_n12926 , 1_n12927 , 1_n12928 , 1_n12929 , 1_n12930 , 1_n12931 , 1_n12932 , 1_n12933 , 1_n12934 , 1_n12935 , 1_n12936 , 1_n12937 , 1_n12938 , 1_n12939 , 1_n12940 , 1_n12941 , 1_n12942 , 1_n12943 , 1_n12944 , 1_n12945 , 1_n12946 , 1_n12947 , 1_n12948 , 1_n12949 , 1_n12950 , 1_n12951 , 1_n12952 , 1_n12953 , 1_n12954 , 1_n12955 , 1_n12956 , 1_n12957 , 1_n12958 , 1_n12959 , 1_n12960 , 1_n12961 , 1_n12962 , 1_n12963 , 1_n12964 , 1_n12966 , 1_n12967 , 1_n12969 , 1_n12970 , 1_n12971 , 1_n12972 , 1_n12973 , 1_n12974 , 1_n12975 , 1_n12976 , 1_n12977 , 1_n12978 , 1_n12979 , 1_n12980 , 1_n12981 , 1_n12982 , 1_n12983 , 1_n12984 , 1_n12985 , 1_n12986 , 1_n12987 , 1_n12988 , 1_n12989 , 1_n12990 , 1_n12991 , 1_n12992 , 1_n12993 , 1_n12994 , 1_n12995 , 1_n12996 , 1_n12997 , 1_n12998 , 1_n12999 , 1_n13000 , 1_n13001 , 1_n13003 , 1_n13004 , 1_n13005 , 1_n13006 , 1_n13007 , 1_n13008 , 1_n13009 , 1_n13010 , 1_n13011 , 1_n13012 , 1_n13013 , 1_n13014 , 1_n13015 , 1_n13016 , 1_n13017 , 1_n13018 , 1_n13019 , 1_n13020 , 1_n13021 , 1_n13022 , 1_n13023 , 1_n13024 , 1_n13025 , 1_n13026 , 1_n13027 , 1_n13028 , 1_n13029 , 1_n13030 , 1_n13031 , 1_n13032 , 1_n13033 , 1_n13034 , 1_n13036 , 1_n13037 , 1_n13038 , 1_n13039 , 1_n13040 , 1_n13041 , 1_n13042 , 1_n13043 , 1_n13044 , 1_n13045 , 1_n13046 , 1_n13047 , 1_n13048 , 1_n13049 , 1_n13050 , 1_n13051 , 1_n13052 , 1_n13053 , 1_n13054 , 1_n13055 , 1_n13056 , 1_n13057 , 1_n13059 , 1_n13061 , 1_n13062 , 1_n13063 , 1_n13064 , 1_n13065 , 1_n13066 , 1_n13067 , 1_n13068 , 1_n13069 , 1_n13070 , 1_n13071 , 1_n13072 , 1_n13073 , 1_n13074 , 1_n13075 , 1_n13076 , 1_n13077 , 1_n13078 , 1_n13079 , 1_n13080 , 1_n13081 , 1_n13082 , 1_n13083 , 1_n13084 , 1_n13085 , 1_n13086 , 1_n13087 , 1_n13088 , 1_n13089 , 1_n13090 , 1_n13091 , 1_n13092 , 1_n13093 , 1_n13094 , 1_n13095 , 1_n13096 , 1_n13097 , 1_n13098 , 1_n13099 , 1_n13100 , 1_n13101 , 1_n13102 , 1_n13103 , 1_n13104 , 1_n13105 , 1_n13106 , 1_n13107 , 1_n13108 , 1_n13109 , 1_n13110 , 1_n13111 , 1_n13112 , 1_n13113 , 1_n13114 , 1_n13115 , 1_n13116 , 1_n13117 , 1_n13118 , 1_n13119 , 1_n13120 , 1_n13121 , 1_n13122 , 1_n13123 , 1_n13124 , 1_n13125 , 1_n13126 , 1_n13127 , 1_n13128 , 1_n13129 , 1_n13130 , 1_n13131 , 1_n13132 , 1_n13133 , 1_n13134 , 1_n13135 , 1_n13136 , 1_n13137 , 1_n13138 , 1_n13139 , 1_n13140 , 1_n13141 , 1_n13142 , 1_n13143 , 1_n13144 , 1_n13145 , 1_n13146 , 1_n13147 , 1_n13148 , 1_n13149 , 1_n13150 , 1_n13151 , 1_n13152 , 1_n13153 , 1_n13154 , 1_n13155 , 1_n13156 , 1_n13157 , 1_n13158 , 1_n13159 , 1_n13160 , 1_n13161 , 1_n13162 , 1_n13163 , 1_n13164 , 1_n13165 , 1_n13166 , 1_n13167 , 1_n13168 , 1_n13169 , 1_n13170 , 1_n13171 , 1_n13172 , 1_n13173 , 1_n13174 , 1_n13175 , 1_n13176 , 1_n13177 , 1_n13178 , 1_n13179 , 1_n13180 , 1_n13181 , 1_n13182 , 1_n13183 , 1_n13184 , 1_n13185 , 1_n13186 , 1_n13187 , 1_n13188 , 1_n13189 , 1_n13190 , 1_n13191 , 1_n13192 , 1_n13193 , 1_n13194 , 1_n13195 , 1_n13196 , 1_n13197 , 1_n13198 , 1_n13199 , 1_n13200 , 1_n13202 , 1_n13203 , 1_n13204 , 1_n13205 , 1_n13206 , 1_n13207 , 1_n13208 , 1_n13209 , 1_n13210 , 1_n13211 , 1_n13212 , 1_n13213 , 1_n13214 , 1_n13215 , 1_n13216 , 1_n13217 , 1_n13218 , 1_n13219 , 1_n13220 , 1_n13221 , 1_n13222 , 1_n13223 , 1_n13224 , 1_n13225 , 1_n13226 , 1_n13227 , 1_n13228 , 1_n13229 , 1_n13230 , 1_n13231 , 1_n13232 , 1_n13233 , 1_n13234 , 1_n13235 , 1_n13236 , 1_n13237 , 1_n13238 , 1_n13239 , 1_n13240 , 1_n13241 , 1_n13242 , 1_n13243 ;
assign 1_n3523 = 1_n7151 & 1_n6767;
assign 1_n1818 = ~(1_n11618 ^ 1_n10125);
assign 1_n6666 = 1_n1354 | 1_n6635;
assign 1_n13003 = 1_n10781 | 1_n8348;
assign 1_n8017 = 1_n995 | 1_n12970;
assign 1_n9879 = 1_n4074 & 1_n12255;
assign 1_n849 = ~(1_n1713 ^ 1_n1158);
assign 1_n837 = ~(1_n3701 | 1_n2651);
assign 1_n3470 = ~(1_n12726 ^ 1_n4668);
assign 1_n6673 = ~(1_n2914 ^ 1_n655);
assign 1_n8353 = ~(1_n3258 ^ 1_n2954);
assign 1_n1644 = 1_n7660 | 1_n10173;
assign 1_n4458 = ~(1_n11074 ^ 1_n9291);
assign 1_n4154 = 1_n12552 | 1_n10871;
assign 1_n5448 = ~1_n13203;
assign 1_n938 = 1_n2711 | 1_n11144;
assign 1_n9174 = ~1_n72;
assign 1_n6954 = 1_n3044 | 1_n11894;
assign 1_n224 = ~(1_n10835 ^ 1_n2683);
assign 1_n7171 = ~1_n2309;
assign 1_n1343 = ~(1_n8789 | 1_n7265);
assign 1_n3099 = ~1_n5324;
assign 1_n12128 = ~1_n5568;
assign 1_n12514 = ~(1_n5673 | 1_n13166);
assign 1_n5497 = 1_n10761 | 1_n6732;
assign 1_n6006 = 1_n3747 & 1_n4857;
assign 1_n8827 = ~(1_n6431 ^ 1_n7145);
assign 1_n9763 = 1_n7126 & 1_n2227;
assign 1_n11908 = 1_n4316 | 1_n2924;
assign 1_n2161 = ~(1_n11270 ^ 1_n1874);
assign 1_n618 = ~(1_n7815 ^ 1_n4460);
assign 1_n1422 = ~1_n12965;
assign 1_n9158 = ~(1_n601 ^ 1_n9373);
assign 1_n9135 = 1_n1550 | 1_n2209;
assign 1_n12910 = 1_n1958 & 1_n4654;
assign 1_n13069 = 1_n10439 | 1_n12388;
assign 1_n13000 = ~(1_n4381 ^ 1_n10298);
assign 1_n12582 = ~(1_n1459 ^ 1_n1950);
assign 1_n1273 = ~(1_n8182 ^ 1_n8861);
assign 1_n11174 = ~1_n485;
assign 1_n5045 = ~1_n5586;
assign 1_n7486 = 1_n6079 | 1_n4448;
assign 1_n9434 = 1_n6006 | 1_n9735;
assign 1_n6268 = 1_n7700 | 1_n1026;
assign 1_n11498 = 1_n6991 | 1_n11644;
assign 1_n1005 = ~1_n10373;
assign 1_n10206 = ~1_n6964;
assign 1_n746 = ~(1_n4418 ^ 1_n496);
assign 1_n12707 = 1_n7675 | 1_n1144;
assign 1_n11383 = 1_n5865 | 1_n5242;
assign 1_n12636 = ~1_n9701;
assign 1_n6506 = ~1_n3311;
assign 1_n5217 = 1_n7939 | 1_n1337;
assign 1_n6028 = ~1_n12482;
assign 1_n7328 = ~(1_n6204 ^ 1_n12282);
assign 1_n3430 = 1_n12568 | 1_n12847;
assign 1_n13217 = ~(1_n8937 ^ 1_n9105);
assign 1_n7035 = ~(1_n3487 ^ 1_n1164);
assign 1_n11295 = 1_n10032 | 1_n7254;
assign 1_n734 = ~1_n11411;
assign 1_n11278 = ~(1_n9811 ^ 1_n9427);
assign 1_n10946 = ~(1_n12215 ^ 1_n3738);
assign 1_n610 = ~(1_n10055 ^ 1_n774);
assign 1_n10496 = ~(1_n10728 ^ 1_n13055);
assign 1_n12601 = ~(1_n3959 ^ 1_n9631);
assign 1_n10620 = 1_n6939 | 1_n9159;
assign 1_n5216 = ~1_n1426;
assign 1_n3802 = ~(1_n596 ^ 1_n1088);
assign 1_n12895 = 1_n13027 | 1_n10662;
assign 1_n11521 = ~1_n9732;
assign 1_n4884 = ~1_n3670;
assign 1_n9741 = ~1_n8078;
assign 1_n1826 = 1_n6083 ^ 1_n7616;
assign 1_n3658 = ~(1_n12111 ^ 1_n4323);
assign 1_n6851 = 1_n11030 & 1_n12289;
assign 1_n10227 = ~(1_n10752 ^ 1_n594);
assign 1_n11559 = 1_n6226 ^ 1_n4888;
assign 1_n127 = 1_n10882 | 1_n11551;
assign 1_n8256 = 1_n7819 | 1_n10043;
assign 1_n10029 = 1_n8852;
assign 1_n4473 = ~1_n2295;
assign 1_n10956 = ~1_n5729;
assign 1_n3456 = ~1_n11682;
assign 1_n9718 = ~1_n6670;
assign 1_n7609 = 1_n8188 | 1_n4490;
assign 1_n10187 = ~(1_n330 | 1_n12782);
assign 1_n5538 = 1_n4081 & 1_n9186;
assign 1_n1464 = ~(1_n520 ^ 1_n7499);
assign 1_n9928 = ~(1_n4616 ^ 1_n9260);
assign 1_n1570 = 1_n12471;
assign 1_n1525 = ~(1_n8885 ^ 1_n10490);
assign 1_n3435 = 1_n3669 & 1_n834;
assign 1_n11902 = 1_n2848 | 1_n12501;
assign 1_n2414 = 1_n4258 | 1_n10106;
assign 1_n252 = 1_n10338 & 1_n6627;
assign 1_n9289 = 1_n1168 | 1_n7723;
assign 1_n12010 = 1_n5480 | 1_n2796;
assign 1_n13046 = ~(1_n6622 ^ 1_n10271);
assign 1_n12280 = 1_n683 | 1_n9080;
assign 1_n7727 = 1_n7912 | 1_n13118;
assign 1_n8096 = ~(1_n8582 ^ 1_n10826);
assign 1_n9186 = 1_n5455 | 1_n4724;
assign 1_n4933 = ~(1_n5944 ^ 1_n5560);
assign 1_n7994 = ~(1_n2528 ^ 1_n8607);
assign 1_n10128 = ~1_n11891;
assign 1_n1597 = 1_n3186 | 1_n3500;
assign 1_n12870 = ~(1_n1824 | 1_n10842);
assign 1_n11470 = 1_n1782 & 1_n10313;
assign 1_n5626 = ~1_n7556;
assign 1_n5131 = ~(1_n7739 ^ 1_n3051);
assign 1_n425 = 1_n1907 & 1_n9672;
assign 1_n7539 = ~(1_n9415 ^ 1_n9935);
assign 1_n3425 = 1_n10761 | 1_n8702;
assign 1_n8270 = ~(1_n465 ^ 1_n727);
assign 1_n12783 = 1_n7695 & 1_n9404;
assign 1_n3269 = ~(1_n6985 ^ 1_n12644);
assign 1_n12026 = 1_n3006 & 1_n6149;
assign 1_n12042 = ~1_n10925;
assign 1_n9682 = ~1_n11324;
assign 1_n10094 = 1_n4795 & 1_n8792;
assign 1_n8499 = ~1_n10451;
assign 1_n12046 = 1_n10812 | 1_n2937;
assign 1_n2932 = ~(1_n4047 ^ 1_n10504);
assign 1_n3026 = 1_n3135 & 1_n5808;
assign 1_n12849 = 1_n8207 & 1_n1545;
assign 1_n4076 = ~(1_n12132 ^ 1_n965);
assign 1_n7769 = 1_n7041 | 1_n12695;
assign 1_n11615 = ~(1_n1868 ^ 1_n639);
assign 1_n12282 = ~(1_n6713 ^ 1_n6848);
assign 1_n4146 = 1_n8868 | 1_n2958;
assign 1_n12518 = ~1_n2646;
assign 1_n4928 = 1_n2430 & 1_n13186;
assign 1_n2372 = ~(1_n8740 ^ 1_n9673);
assign 1_n1964 = ~(1_n12106 ^ 1_n11044);
assign 1_n2158 = 1_n5607 | 1_n9431;
assign 1_n12165 = 1_n12737 | 1_n5956;
assign 1_n9096 = 1_n11398 & 1_n5467;
assign 1_n6181 = 1_n5378 & 1_n7277;
assign 1_n10765 = ~(1_n5090 ^ 1_n5825);
assign 1_n10235 = 1_n7933 | 1_n7244;
assign 1_n10691 = 1_n4755 | 1_n10289;
assign 1_n11500 = ~(1_n7563 ^ 1_n3718);
assign 1_n2741 = ~(1_n10187 ^ 1_n4817);
assign 1_n12881 = ~1_n4470;
assign 1_n8882 = 1_n48 | 1_n4947;
assign 1_n12252 = 1_n5759 & 1_n664;
assign 1_n11017 = ~(1_n5932 ^ 1_n284);
assign 1_n8688 = 1_n2580 | 1_n7533;
assign 1_n6625 = 1_n7931 | 1_n11255;
assign 1_n7215 = 1_n11183 | 1_n7859;
assign 1_n10018 = ~1_n8468;
assign 1_n3622 = 1_n8063 & 1_n3371;
assign 1_n11049 = ~(1_n2108 ^ 1_n7715);
assign 1_n7369 = ~(1_n2074 | 1_n6239);
assign 1_n7264 = ~(1_n3499 ^ 1_n5493);
assign 1_n15 = ~(1_n2867 | 1_n11302);
assign 1_n6977 = 1_n7625 & 1_n3577;
assign 1_n1657 = ~(1_n1414 ^ 1_n11594);
assign 1_n8071 = 1_n11471 & 1_n3006;
assign 1_n8822 = 1_n2106 & 1_n10607;
assign 1_n8482 = ~(1_n8706 ^ 1_n9916);
assign 1_n6836 = 1_n6039 & 1_n5862;
assign 1_n8910 = ~(1_n745 | 1_n1899);
assign 1_n6581 = ~1_n12682;
assign 1_n4969 = 1_n264 & 1_n10423;
assign 1_n4875 = ~1_n1198;
assign 1_n7723 = 1_n10879;
assign 1_n4889 = 1_n10680 & 1_n4121;
assign 1_n1511 = ~1_n12263;
assign 1_n10200 = 1_n5671 & 1_n8233;
assign 1_n9518 = 1_n6162 & 1_n8361;
assign 1_n3167 = ~1_n2840;
assign 1_n12055 = 1_n9429 | 1_n12501;
assign 1_n3747 = ~(1_n8035 ^ 1_n9201);
assign 1_n1459 = ~(1_n1525 ^ 1_n4142);
assign 1_n7157 = ~(1_n2593 ^ 1_n8114);
assign 1_n2025 = 1_n4595 | 1_n11343;
assign 1_n8315 = ~1_n772;
assign 1_n5117 = 1_n8183 & 1_n10606;
assign 1_n10969 = ~(1_n2741 ^ 1_n7724);
assign 1_n9023 = 1_n1365 | 1_n11162;
assign 1_n11207 = ~(1_n4982 ^ 1_n12583);
assign 1_n8844 = ~(1_n9406 ^ 1_n3154);
assign 1_n5897 = ~(1_n405 ^ 1_n1808);
assign 1_n9959 = 1_n5670 | 1_n10135;
assign 1_n5651 = ~(1_n3346 ^ 1_n1154);
assign 1_n2272 = 1_n965 | 1_n7619;
assign 1_n12545 = ~(1_n6303 ^ 1_n2855);
assign 1_n6019 = ~(1_n1466 ^ 1_n5895);
assign 1_n7748 = ~1_n772;
assign 1_n1773 = 1_n5605 | 1_n5868;
assign 1_n5741 = ~(1_n123 ^ 1_n5069);
assign 1_n8776 = ~1_n401;
assign 1_n6970 = 1_n7597 | 1_n6265;
assign 1_n7467 = ~(1_n2424 ^ 1_n5326);
assign 1_n1797 = 1_n11535 & 1_n8925;
assign 1_n663 = ~1_n12379;
assign 1_n3064 = ~(1_n4914 ^ 1_n10942);
assign 1_n3127 = ~1_n6818;
assign 1_n5021 = 1_n11125 | 1_n998;
assign 1_n7406 = ~(1_n13149 ^ 1_n9556);
assign 1_n7055 = ~1_n10418;
assign 1_n5403 = ~(1_n9797 ^ 1_n1532);
assign 1_n8895 = ~(1_n4557 ^ 1_n11784);
assign 1_n12945 = ~(1_n681 | 1_n8347);
assign 1_n6336 = 1_n6743 | 1_n4936;
assign 1_n9803 = 1_n59 | 1_n5406;
assign 1_n8253 = 1_n10998 & 1_n11890;
assign 1_n1039 = ~1_n224;
assign 1_n12475 = 1_n7125 & 1_n12365;
assign 1_n1123 = ~(1_n11737 ^ 1_n2953);
assign 1_n4878 = 1_n3122 | 1_n10100;
assign 1_n12483 = ~1_n12853;
assign 1_n11066 = ~(1_n9898 ^ 1_n2);
assign 1_n9060 = 1_n454 | 1_n2192;
assign 1_n6801 = ~(1_n2647 ^ 1_n58);
assign 1_n11464 = 1_n4808 | 1_n2133;
assign 1_n56 = ~1_n12893;
assign 1_n3394 = 1_n2109 | 1_n2232;
assign 1_n8591 = ~(1_n5698 ^ 1_n3242);
assign 1_n12397 = 1_n2986 & 1_n1262;
assign 1_n5936 = 1_n11482 | 1_n8822;
assign 1_n12536 = 1_n3346 | 1_n10828;
assign 1_n182 = 1_n7840 & 1_n12178;
assign 1_n5374 = 1_n8977 | 1_n6404;
assign 1_n5665 = 1_n5260 | 1_n7302;
assign 1_n6797 = 1_n1329 | 1_n12847;
assign 1_n11384 = 1_n10300 & 1_n5027;
assign 1_n544 = ~1_n7328;
assign 1_n9948 = 1_n13239 & 1_n826;
assign 1_n7302 = ~(1_n972 | 1_n10692);
assign 1_n12985 = ~(1_n12564 ^ 1_n295);
assign 1_n6934 = 1_n4842 | 1_n1686;
assign 1_n10213 = ~1_n11488;
assign 1_n4065 = ~(1_n9986 ^ 1_n9694);
assign 1_n4118 = ~(1_n4117 | 1_n3250);
assign 1_n548 = ~(1_n3150 ^ 1_n6695);
assign 1_n11717 = 1_n850 | 1_n6339;
assign 1_n10634 = ~(1_n641 ^ 1_n12418);
assign 1_n2885 = ~(1_n8464 ^ 1_n9392);
assign 1_n7889 = 1_n6250 | 1_n479;
assign 1_n10884 = 1_n5639 & 1_n7441;
assign 1_n4336 = 1_n6699 | 1_n9784;
assign 1_n7686 = ~(1_n4311 ^ 1_n7280);
assign 1_n4585 = 1_n6714 & 1_n12135;
assign 1_n5941 = ~(1_n7983 ^ 1_n10957);
assign 1_n2699 = ~(1_n2064 ^ 1_n6719);
assign 1_n1667 = 1_n12621 | 1_n12695;
assign 1_n1128 = 1_n5597 | 1_n5846;
assign 1_n7241 = ~(1_n1858 ^ 1_n8884);
assign 1_n4706 = 1_n7207 | 1_n6789;
assign 1_n12100 = ~(1_n8789 ^ 1_n11047);
assign 1_n1720 = ~1_n854;
assign 1_n1727 = 1_n7903 | 1_n12768;
assign 1_n2694 = 1_n3859 & 1_n10391;
assign 1_n11269 = 1_n10950 | 1_n7723;
assign 1_n12665 = 1_n3311 & 1_n854;
assign 1_n9038 = ~(1_n4915 ^ 1_n11245);
assign 1_n7103 = 1_n8280 ^ 1_n7205;
assign 1_n11224 = ~(1_n1700 ^ 1_n6224);
assign 1_n10194 = ~(1_n7726 ^ 1_n9611);
assign 1_n8063 = 1_n7571 | 1_n9749;
assign 1_n9003 = 1_n1986 | 1_n5515;
assign 1_n2603 = ~(1_n11198 ^ 1_n9001);
assign 1_n12041 = ~(1_n12652 | 1_n12699);
assign 1_n10243 = ~(1_n9664 ^ 1_n5837);
assign 1_n8126 = ~(1_n3976 | 1_n3723);
assign 1_n509 = ~(1_n11533 ^ 1_n8434);
assign 1_n926 = ~(1_n10067 | 1_n11759);
assign 1_n3428 = ~1_n772;
assign 1_n6790 = 1_n10770 & 1_n8290;
assign 1_n7120 = ~(1_n10782 ^ 1_n12379);
assign 1_n1432 = 1_n10770 & 1_n8506;
assign 1_n3993 = ~(1_n3936 | 1_n4810);
assign 1_n8434 = 1_n10287 | 1_n4724;
assign 1_n10369 = 1_n2036 & 1_n2434;
assign 1_n2820 = ~(1_n5750 ^ 1_n5873);
assign 1_n11906 = ~(1_n11583 ^ 1_n11939);
assign 1_n10844 = ~(1_n6507 | 1_n5848);
assign 1_n5991 = ~(1_n11605 ^ 1_n3565);
assign 1_n3182 = ~(1_n12290 ^ 1_n207);
assign 1_n1127 = 1_n6084 & 1_n8061;
assign 1_n8535 = ~(1_n7139 ^ 1_n886);
assign 1_n6715 = 1_n8625 & 1_n9970;
assign 1_n12405 = ~(1_n9026 ^ 1_n1435);
assign 1_n12489 = 1_n869 & 1_n11564;
assign 1_n10275 = 1_n12829 | 1_n6461;
assign 1_n6766 = ~(1_n10996 | 1_n12420);
assign 1_n895 = 1_n11793 | 1_n4354;
assign 1_n6200 = ~(1_n1966 ^ 1_n3658);
assign 1_n5125 = 1_n7216 | 1_n4947;
assign 1_n8232 = 1_n2916 & 1_n4466;
assign 1_n3698 = ~1_n3085;
assign 1_n9623 = 1_n4884 & 1_n1116;
assign 1_n5759 = ~(1_n11271 ^ 1_n1944);
assign 1_n7298 = 1_n12955 | 1_n8360;
assign 1_n13065 = ~(1_n11051 ^ 1_n5718);
assign 1_n4814 = 1_n3158 | 1_n2133;
assign 1_n12076 = 1_n10448 | 1_n11101;
assign 1_n3499 = 1_n9170 & 1_n4661;
assign 1_n7258 = ~1_n966;
assign 1_n5466 = ~1_n9831;
assign 1_n9354 = 1_n6964 | 1_n1211;
assign 1_n684 = 1_n156 & 1_n2342;
assign 1_n13035 = ~(1_n680 ^ 1_n2364);
assign 1_n1952 = 1_n10369 | 1_n12854;
assign 1_n7505 = 1_n9975 & 1_n5700;
assign 1_n1378 = ~(1_n7408 ^ 1_n893);
assign 1_n3432 = ~(1_n4910 | 1_n2820);
assign 1_n7681 = 1_n11391 & 1_n516;
assign 1_n1009 = ~(1_n4594 ^ 1_n11293);
assign 1_n11528 = ~(1_n12916 ^ 1_n2735);
assign 1_n5451 = 1_n3049 | 1_n11137;
assign 1_n870 = ~(1_n5330 ^ 1_n8870);
assign 1_n11889 = 1_n11092 | 1_n8712;
assign 1_n274 = ~(1_n10086 | 1_n1322);
assign 1_n1816 = ~(1_n5099 | 1_n364);
assign 1_n8711 = 1_n3488 & 1_n5835;
assign 1_n8045 = ~(1_n11306 ^ 1_n1909);
assign 1_n5854 = ~1_n9654;
assign 1_n4148 = 1_n6718 & 1_n8567;
assign 1_n6276 = ~1_n7969;
assign 1_n2215 = ~1_n10264;
assign 1_n10363 = 1_n2785 | 1_n10802;
assign 1_n3736 = 1_n4029 | 1_n12800;
assign 1_n392 = ~1_n10805;
assign 1_n1523 = ~(1_n8333 ^ 1_n2906);
assign 1_n5909 = 1_n11344 | 1_n9480;
assign 1_n9058 = ~(1_n7915 ^ 1_n4106);
assign 1_n6101 = ~1_n6080;
assign 1_n4479 = 1_n1320 | 1_n4237;
assign 1_n1323 = ~1_n9887;
assign 1_n2727 = 1_n7455 | 1_n7734;
assign 1_n3146 = 1_n1527 & 1_n6961;
assign 1_n8865 = ~(1_n4591 | 1_n1885);
assign 1_n3829 = ~1_n6124;
assign 1_n3233 = ~(1_n11991 ^ 1_n7273);
assign 1_n8698 = ~(1_n11223 ^ 1_n9998);
assign 1_n11480 = ~(1_n9789 ^ 1_n5206);
assign 1_n4666 = 1_n8675 | 1_n7127;
assign 1_n6098 = 1_n7657 | 1_n11608;
assign 1_n3812 = 1_n1475 | 1_n1714;
assign 1_n10472 = ~(1_n13151 ^ 1_n5156);
assign 1_n2397 = ~(1_n8743 ^ 1_n408);
assign 1_n4537 = ~1_n10866;
assign 1_n7474 = 1_n5126 & 1_n7225;
assign 1_n7175 = ~(1_n4591 ^ 1_n9284);
assign 1_n10810 = 1_n17 & 1_n11460;
assign 1_n6935 = ~(1_n3991 ^ 1_n12749);
assign 1_n2867 = ~(1_n8207 | 1_n1545);
assign 1_n12294 = 1_n560 | 1_n7530;
assign 1_n5141 = 1_n10109 | 1_n62;
assign 1_n5614 = 1_n8289 & 1_n5294;
assign 1_n11789 = ~(1_n996 ^ 1_n11902);
assign 1_n8977 = ~1_n1650;
assign 1_n8289 = ~(1_n4193 ^ 1_n12634);
assign 1_n230 = 1_n7395 | 1_n8535;
assign 1_n3147 = ~(1_n10089 ^ 1_n6641);
assign 1_n3582 = 1_n8074 | 1_n7668;
assign 1_n3248 = 1_n8976 & 1_n13179;
assign 1_n5393 = ~(1_n513 ^ 1_n651);
assign 1_n4574 = 1_n6295 | 1_n12188;
assign 1_n12391 = ~1_n6155;
assign 1_n533 = ~(1_n6504 | 1_n9459);
assign 1_n51 = 1_n3260 | 1_n10823;
assign 1_n10044 = 1_n6949 | 1_n7524;
assign 1_n8003 = ~(1_n8072 ^ 1_n4549);
assign 1_n2402 = ~(1_n10052 ^ 1_n10264);
assign 1_n1561 = ~(1_n11576 ^ 1_n12742);
assign 1_n2185 = 1_n11102 ^ 1_n12014;
assign 1_n8205 = ~(1_n5664 ^ 1_n3556);
assign 1_n5438 = 1_n694 | 1_n6635;
assign 1_n11137 = ~1_n9475;
assign 1_n4718 = ~(1_n7818 ^ 1_n7274);
assign 1_n2290 = 1_n10375 & 1_n1128;
assign 1_n9296 = ~1_n5770;
assign 1_n2386 = ~1_n5136;
assign 1_n1843 = 1_n2767 & 1_n10584;
assign 1_n9720 = ~1_n7330;
assign 1_n855 = ~1_n11473;
assign 1_n332 = 1_n67 & 1_n2774;
assign 1_n10445 = 1_n13234 & 1_n2257;
assign 1_n1752 = ~(1_n10102 ^ 1_n11894);
assign 1_n12259 = 1_n4272 | 1_n12847;
assign 1_n429 = ~(1_n13177 ^ 1_n2844);
assign 1_n9627 = ~(1_n9654 | 1_n11323);
assign 1_n3695 = 1_n13082 | 1_n12273;
assign 1_n2591 = 1_n7718 | 1_n5242;
assign 1_n90 = 1_n8339 & 1_n8542;
assign 1_n1663 = ~1_n8137;
assign 1_n8095 = ~(1_n12747 | 1_n10337);
assign 1_n7881 = ~(1_n12896 | 1_n3312);
assign 1_n10569 = ~(1_n12468 ^ 1_n1255);
assign 1_n7775 = ~(1_n1632 | 1_n12013);
assign 1_n1531 = ~(1_n13132 | 1_n3777);
assign 1_n9569 = ~1_n4712;
assign 1_n6228 = 1_n761 & 1_n834;
assign 1_n3946 = ~(1_n11968 ^ 1_n12523);
assign 1_n9352 = 1_n4745 & 1_n12411;
assign 1_n2675 = 1_n5045;
assign 1_n9577 = 1_n2486 ^ 1_n11084;
assign 1_n6099 = ~1_n287;
assign 1_n4341 = ~(1_n4533 ^ 1_n12320);
assign 1_n1594 = 1_n3613 | 1_n9130;
assign 1_n8671 = ~1_n5800;
assign 1_n6873 = 1_n10501 | 1_n12959;
assign 1_n178 = 1_n10343 | 1_n9182;
assign 1_n13113 = 1_n3453 & 1_n5335;
assign 1_n11699 = ~(1_n9176 ^ 1_n3054);
assign 1_n6311 = ~(1_n3400 ^ 1_n1203);
assign 1_n11801 = 1_n1406 | 1_n8534;
assign 1_n7251 = 1_n4994 & 1_n10077;
assign 1_n12189 = 1_n2853 & 1_n2854;
assign 1_n5069 = 1_n2850 & 1_n8526;
assign 1_n1955 = 1_n3068 | 1_n6732;
assign 1_n5377 = ~1_n10405;
assign 1_n4152 = ~1_n3918;
assign 1_n6769 = 1_n9272;
assign 1_n5399 = 1_n3607 & 1_n8996;
assign 1_n2997 = ~(1_n4593 | 1_n6096);
assign 1_n10914 = 1_n3415 & 1_n11558;
assign 1_n2496 = ~(1_n5094 ^ 1_n7517);
assign 1_n11981 = 1_n7543 & 1_n931;
assign 1_n739 = 1_n9793 | 1_n12789;
assign 1_n3519 = 1_n2107 & 1_n8548;
assign 1_n1193 = ~1_n11325;
assign 1_n12300 = 1_n1213 | 1_n7682;
assign 1_n5727 = ~(1_n11867 ^ 1_n421);
assign 1_n11662 = 1_n1735 | 1_n10674;
assign 1_n11301 = ~(1_n6653 | 1_n7490);
assign 1_n7195 = 1_n4016 | 1_n4095;
assign 1_n1514 = 1_n1090 | 1_n1292;
assign 1_n2389 = ~(1_n2023 ^ 1_n5824);
assign 1_n2911 = ~(1_n10278 | 1_n1441);
assign 1_n8704 = 1_n2615 | 1_n2871;
assign 1_n5375 = ~1_n7877;
assign 1_n2898 = ~(1_n4861 ^ 1_n8377);
assign 1_n4381 = ~(1_n3291 ^ 1_n3601);
assign 1_n7605 = 1_n12568 | 1_n12273;
assign 1_n4105 = 1_n4539 | 1_n11234;
assign 1_n3697 = ~(1_n7549 | 1_n2597);
assign 1_n463 = ~(1_n3247 ^ 1_n3560);
assign 1_n2596 = 1_n8613 | 1_n7312;
assign 1_n2478 = ~1_n11468;
assign 1_n13056 = 1_n6489 ^ 1_n2342;
assign 1_n2996 = 1_n1375 & 1_n12097;
assign 1_n9031 = ~(1_n377 ^ 1_n10083);
assign 1_n3689 = ~(1_n5030 | 1_n12908);
assign 1_n4506 = 1_n4044 | 1_n12672;
assign 1_n1419 = 1_n3534 | 1_n4947;
assign 1_n8101 = 1_n2609 & 1_n5342;
assign 1_n3043 = ~(1_n6049 ^ 1_n8427);
assign 1_n5126 = ~(1_n10506 ^ 1_n10151);
assign 1_n3081 = ~(1_n12492 ^ 1_n7263);
assign 1_n11804 = ~(1_n7304 | 1_n11649);
assign 1_n3982 = 1_n9882 | 1_n4373;
assign 1_n2457 = 1_n4001 ^ 1_n9692;
assign 1_n3511 = ~(1_n10667 ^ 1_n11474);
assign 1_n4502 = ~(1_n7870 | 1_n5043);
assign 1_n1971 = 1_n6668 & 1_n12853;
assign 1_n399 = 1_n3544 | 1_n1702;
assign 1_n9564 = 1_n7095 & 1_n4211;
assign 1_n6266 = ~(1_n10405 | 1_n608);
assign 1_n12834 = ~1_n5758;
assign 1_n9321 = ~1_n5094;
assign 1_n5198 = ~(1_n2237 | 1_n9953);
assign 1_n12272 = ~1_n983;
assign 1_n7857 = 1_n4004 | 1_n9549;
assign 1_n7666 = ~(1_n3916 ^ 1_n4907);
assign 1_n1115 = ~(1_n5410 ^ 1_n2779);
assign 1_n5408 = ~(1_n3985 ^ 1_n885);
assign 1_n10498 = 1_n10013 ^ 1_n12578;
assign 1_n6375 = ~1_n469;
assign 1_n3083 = 1_n10188 | 1_n3963;
assign 1_n10718 = ~(1_n10888 ^ 1_n4826);
assign 1_n8854 = ~(1_n11573 ^ 1_n9844);
assign 1_n210 = 1_n1934 & 1_n1234;
assign 1_n11453 = 1_n4467 | 1_n12142;
assign 1_n11636 = 1_n6355 | 1_n3890;
assign 1_n10322 = 1_n4382 & 1_n1636;
assign 1_n292 = 1_n13229 & 1_n7849;
assign 1_n9220 = 1_n5005 & 1_n13110;
assign 1_n1930 = ~1_n7374;
assign 1_n9271 = ~(1_n1880 ^ 1_n6551);
assign 1_n4672 = ~(1_n10482 ^ 1_n4254);
assign 1_n2409 = 1_n8661 & 1_n5568;
assign 1_n10371 = ~(1_n10940 ^ 1_n5821);
assign 1_n9032 = 1_n78 & 1_n116;
assign 1_n7027 = ~(1_n11092 ^ 1_n8712);
assign 1_n7525 = ~(1_n5996 ^ 1_n6844);
assign 1_n6474 = 1_n1514 & 1_n8318;
assign 1_n7432 = 1_n241 | 1_n9070;
assign 1_n10678 = 1_n3299 | 1_n7741;
assign 1_n2549 = ~(1_n4889 ^ 1_n1122);
assign 1_n2497 = ~(1_n2176 ^ 1_n10951);
assign 1_n6026 = ~(1_n12553 ^ 1_n4350);
assign 1_n6046 = ~1_n11830;
assign 1_n1271 = ~1_n972;
assign 1_n3381 = ~(1_n10378 | 1_n4249);
assign 1_n11526 = ~(1_n11658 ^ 1_n5101);
assign 1_n5339 = ~(1_n6859 ^ 1_n4823);
assign 1_n933 = 1_n2263 & 1_n1443;
assign 1_n10111 = 1_n12972 & 1_n3927;
assign 1_n3969 = ~(1_n988 ^ 1_n4873);
assign 1_n3765 = ~(1_n3214 ^ 1_n7173);
assign 1_n2361 = 1_n1175 & 1_n8084;
assign 1_n4052 = ~(1_n10931 ^ 1_n13164);
assign 1_n6662 = ~(1_n6515 ^ 1_n8755);
assign 1_n765 = ~1_n9;
assign 1_n6541 = 1_n13109 & 1_n12435;
assign 1_n9259 = 1_n5545 & 1_n2025;
assign 1_n9554 = ~(1_n2044 ^ 1_n13048);
assign 1_n11395 = 1_n11331 & 1_n2881;
assign 1_n11489 = 1_n5440 | 1_n2244;
assign 1_n8091 = 1_n3047 | 1_n12273;
assign 1_n8203 = ~(1_n5798 ^ 1_n6252);
assign 1_n6681 = ~(1_n3205 ^ 1_n9751);
assign 1_n8349 = 1_n8206 | 1_n2059;
assign 1_n7052 = ~1_n8253;
assign 1_n7594 = ~(1_n3504 | 1_n13045);
assign 1_n12464 = ~(1_n12628 | 1_n5484);
assign 1_n5388 = ~(1_n9095 | 1_n3813);
assign 1_n4931 = ~(1_n12021 ^ 1_n6893);
assign 1_n10179 = 1_n2623;
assign 1_n2164 = ~(1_n228 ^ 1_n6127);
assign 1_n7297 = 1_n12050 | 1_n4899;
assign 1_n2307 = ~1_n3496;
assign 1_n1474 = 1_n2247 & 1_n12928;
assign 1_n12274 = 1_n3099 | 1_n3074;
assign 1_n4948 = ~(1_n5561 ^ 1_n2060);
assign 1_n9880 = 1_n9722 | 1_n9974;
assign 1_n8188 = ~1_n761;
assign 1_n1910 = 1_n2425 & 1_n2380;
assign 1_n1330 = ~(1_n4977 ^ 1_n1221);
assign 1_n6567 = ~(1_n2732 | 1_n11081);
assign 1_n5706 = ~(1_n3305 ^ 1_n9368);
assign 1_n8665 = ~1_n4743;
assign 1_n6879 = 1_n1059 & 1_n6856;
assign 1_n5417 = ~(1_n4427 | 1_n5663);
assign 1_n2569 = 1_n11617 & 1_n11630;
assign 1_n150 = 1_n10943 | 1_n6511;
assign 1_n5642 = ~(1_n1143 ^ 1_n6994);
assign 1_n2342 = 1_n1364 & 1_n3815;
assign 1_n10507 = 1_n7669 | 1_n9101;
assign 1_n5389 = 1_n10253 ^ 1_n12182;
assign 1_n13198 = ~1_n4337;
assign 1_n8336 = ~(1_n7491 ^ 1_n1362);
assign 1_n11164 = 1_n4625 & 1_n9331;
assign 1_n9237 = 1_n8386 | 1_n615;
assign 1_n6491 = 1_n9702 | 1_n1571;
assign 1_n8204 = 1_n228 & 1_n2829;
assign 1_n1520 = 1_n1270 | 1_n6903;
assign 1_n11777 = ~(1_n13180 ^ 1_n3624);
assign 1_n2242 = ~(1_n2014 ^ 1_n13224);
assign 1_n11936 = ~(1_n9678 ^ 1_n9999);
assign 1_n3480 = 1_n2156 & 1_n7971;
assign 1_n3327 = 1_n8653 & 1_n2808;
assign 1_n986 = ~(1_n6761 | 1_n2571);
assign 1_n649 = 1_n1769 & 1_n12117;
assign 1_n10528 = ~(1_n5421 | 1_n9376);
assign 1_n5825 = ~(1_n7638 ^ 1_n3728);
assign 1_n7667 = 1_n12246 & 1_n888;
assign 1_n5062 = ~(1_n10288 ^ 1_n1014);
assign 1_n809 = 1_n10434 | 1_n12723;
assign 1_n2516 = 1_n12930 | 1_n1144;
assign 1_n12791 = 1_n10558 | 1_n12273;
assign 1_n5917 = ~1_n1707;
assign 1_n10134 = 1_n11635 & 1_n2482;
assign 1_n3524 = ~1_n4574;
assign 1_n4204 = 1_n5842 | 1_n10761;
assign 1_n10913 = ~(1_n8382 ^ 1_n4813);
assign 1_n9727 = 1_n4275 | 1_n9842;
assign 1_n501 = ~(1_n11461 ^ 1_n2444);
assign 1_n3544 = 1_n13218 & 1_n9420;
assign 1_n3000 = 1_n10097 & 1_n12071;
assign 1_n379 = ~1_n5536;
assign 1_n12648 = ~1_n1982;
assign 1_n107 = ~1_n10537;
assign 1_n11887 = ~1_n4479;
assign 1_n1666 = ~(1_n10902 ^ 1_n12198);
assign 1_n9122 = 1_n12324 | 1_n2133;
assign 1_n3828 = 1_n8077 & 1_n9720;
assign 1_n2725 = ~1_n4688;
assign 1_n3496 = ~(1_n5593 ^ 1_n5055);
assign 1_n10149 = 1_n12832 ^ 1_n1174;
assign 1_n5725 = 1_n3352 ^ 1_n3435;
assign 1_n8495 = 1_n12643 & 1_n11888;
assign 1_n10348 = ~(1_n535 ^ 1_n7178);
assign 1_n1388 = ~1_n9428;
assign 1_n5130 = 1_n3928 | 1_n1985;
assign 1_n2031 = ~(1_n11266 ^ 1_n3774);
assign 1_n5562 = ~1_n10408;
assign 1_n3645 = 1_n10416 & 1_n12306;
assign 1_n12119 = 1_n9323 | 1_n1797;
assign 1_n3302 = 1_n1919 | 1_n4373;
assign 1_n10622 = ~(1_n10688 ^ 1_n9990);
assign 1_n6263 = ~(1_n2363 ^ 1_n11420);
assign 1_n39 = ~1_n4240;
assign 1_n2081 = ~1_n9794;
assign 1_n3477 = 1_n12563 | 1_n4949;
assign 1_n4950 = 1_n7457 & 1_n3117;
assign 1_n1220 = 1_n5583 | 1_n6017;
assign 1_n1176 = 1_n10037 | 1_n4373;
assign 1_n502 = ~(1_n4486 ^ 1_n8345);
assign 1_n5047 = 1_n1208 & 1_n7264;
assign 1_n45 = ~1_n1084;
assign 1_n9656 = 1_n5297 | 1_n11619;
assign 1_n5033 = 1_n3752 & 1_n6153;
assign 1_n2712 = 1_n2849 | 1_n2793;
assign 1_n11275 = 1_n5058 & 1_n1922;
assign 1_n13171 = ~(1_n9972 ^ 1_n9555);
assign 1_n672 = ~1_n192;
assign 1_n9274 = ~(1_n8133 ^ 1_n3302);
assign 1_n11590 = ~(1_n11954 ^ 1_n12210);
assign 1_n11495 = 1_n60 & 1_n5230;
assign 1_n2905 = ~(1_n5034 | 1_n4222);
assign 1_n5159 = ~(1_n1062 ^ 1_n3947);
assign 1_n9641 = ~1_n988;
assign 1_n7598 = 1_n11987 | 1_n3019;
assign 1_n2616 = ~(1_n5929 | 1_n10215);
assign 1_n188 = 1_n9059 | 1_n4089;
assign 1_n9469 = ~(1_n5736 ^ 1_n3986);
assign 1_n6938 = 1_n2024 & 1_n6508;
assign 1_n1448 = 1_n1263 | 1_n4058;
assign 1_n3772 = 1_n10189 & 1_n7743;
assign 1_n11589 = ~(1_n87 ^ 1_n7373);
assign 1_n1943 = 1_n6583 & 1_n7231;
assign 1_n12342 = 1_n6816 | 1_n4551;
assign 1_n10636 = ~1_n7845;
assign 1_n5678 = ~(1_n2644 ^ 1_n6709);
assign 1_n4456 = 1_n11449 | 1_n8348;
assign 1_n4644 = 1_n10603 & 1_n6540;
assign 1_n7554 = ~(1_n7099 ^ 1_n2620);
assign 1_n459 = ~(1_n9851 ^ 1_n5144);
assign 1_n7349 = ~(1_n7484 | 1_n3848);
assign 1_n11018 = ~1_n4006;
assign 1_n12926 = ~1_n12867;
assign 1_n7704 = 1_n7232 & 1_n8733;
assign 1_n6699 = ~1_n5189;
assign 1_n3956 = 1_n2289 | 1_n3538;
assign 1_n10422 = 1_n2457 | 1_n8964;
assign 1_n4266 = ~(1_n12250 | 1_n8692);
assign 1_n3169 = ~1_n10908;
assign 1_n6909 = 1_n518 & 1_n7776;
assign 1_n10542 = ~(1_n5695 ^ 1_n7339);
assign 1_n1094 = ~1_n5244;
assign 1_n4697 = ~(1_n12184 | 1_n10030);
assign 1_n9731 = 1_n1360 | 1_n3972;
assign 1_n12155 = 1_n6177 & 1_n5857;
assign 1_n594 = ~(1_n13187 ^ 1_n12641);
assign 1_n10143 = ~1_n9570;
assign 1_n11515 = 1_n2246 | 1_n6145;
assign 1_n3713 = ~(1_n6058 ^ 1_n2976);
assign 1_n13109 = 1_n1131 | 1_n1153;
assign 1_n2260 = ~(1_n3272 | 1_n12869);
assign 1_n6139 = 1_n12485 | 1_n9192;
assign 1_n8594 = 1_n4515 | 1_n10681;
assign 1_n1229 = 1_n599 & 1_n876;
assign 1_n8019 = ~1_n8410;
assign 1_n11928 = ~1_n6826;
assign 1_n2766 = 1_n1438 | 1_n1985;
assign 1_n6868 = ~(1_n3260 ^ 1_n1913);
assign 1_n8169 = ~(1_n3448 | 1_n8317);
assign 1_n2393 = 1_n2458 & 1_n3409;
assign 1_n3007 = 1_n9450 | 1_n12623;
assign 1_n5048 = ~1_n3085;
assign 1_n9266 = 1_n6254 | 1_n8326;
assign 1_n4453 = ~1_n951;
assign 1_n10011 = 1_n4088 & 1_n7043;
assign 1_n10056 = 1_n8108 | 1_n10179;
assign 1_n6860 = ~(1_n4528 | 1_n12906);
assign 1_n3010 = ~(1_n3366 ^ 1_n570);
assign 1_n11130 = ~1_n180;
assign 1_n1338 = ~(1_n8368 | 1_n9441);
assign 1_n2371 = ~(1_n7879 ^ 1_n6997);
assign 1_n3974 = ~(1_n4113 ^ 1_n1707);
assign 1_n10043 = ~1_n3085;
assign 1_n6331 = 1_n1936 & 1_n4383;
assign 1_n8636 = 1_n4148 | 1_n900;
assign 1_n3218 = ~(1_n8042 | 1_n2533);
assign 1_n6755 = ~1_n8768;
assign 1_n1336 = ~(1_n11262 ^ 1_n5379);
assign 1_n954 = 1_n11355 & 1_n7774;
assign 1_n8211 = 1_n8843 | 1_n4640;
assign 1_n3813 = ~1_n5073;
assign 1_n5895 = ~(1_n11448 ^ 1_n9226);
assign 1_n644 = ~1_n3669;
assign 1_n10737 = ~(1_n10735 ^ 1_n5276);
assign 1_n11979 = ~(1_n129 ^ 1_n2929);
assign 1_n4557 = 1_n428 & 1_n5117;
assign 1_n9241 = ~(1_n798 ^ 1_n7603);
assign 1_n1227 = 1_n3965 | 1_n5460;
assign 1_n12060 = 1_n11203 | 1_n3926;
assign 1_n3483 = 1_n1712 | 1_n12784;
assign 1_n279 = ~(1_n1801 | 1_n2477);
assign 1_n10673 = ~1_n6956;
assign 1_n6206 = ~(1_n8926 ^ 1_n9469);
assign 1_n9026 = 1_n4980 | 1_n2875;
assign 1_n6117 = ~(1_n91 | 1_n7641);
assign 1_n8847 = 1_n53 | 1_n10761;
assign 1_n9255 = 1_n2973 | 1_n5646;
assign 1_n27 = ~(1_n9633 ^ 1_n12887);
assign 1_n11775 = 1_n6140 & 1_n3031;
assign 1_n3768 = 1_n5922 | 1_n7874;
assign 1_n9249 = 1_n11591 | 1_n10319;
assign 1_n741 = 1_n3077 & 1_n2687;
assign 1_n9369 = 1_n12262 & 1_n3227;
assign 1_n7999 = 1_n5401 | 1_n13039;
assign 1_n3665 = 1_n9392 | 1_n8464;
assign 1_n5046 = ~(1_n12899 ^ 1_n6899);
assign 1_n5929 = ~(1_n10865 ^ 1_n3010);
assign 1_n11044 = ~(1_n7929 ^ 1_n7735);
assign 1_n1542 = 1_n6606 | 1_n8504;
assign 1_n12327 = 1_n12798 | 1_n12240;
assign 1_n8181 = ~(1_n9059 ^ 1_n4089);
assign 1_n5402 = ~1_n7841;
assign 1_n1298 = ~(1_n9307 ^ 1_n9097);
assign 1_n7463 = 1_n7296 & 1_n8914;
assign 1_n8970 = ~(1_n2205 ^ 1_n2654);
assign 1_n985 = ~(1_n6362 ^ 1_n7772);
assign 1_n393 = ~(1_n576 ^ 1_n3757);
assign 1_n7286 = ~1_n6347;
assign 1_n12809 = 1_n5806 | 1_n121;
assign 1_n8944 = ~(1_n7786 | 1_n9562);
assign 1_n1592 = 1_n7086 & 1_n666;
assign 1_n11884 = ~(1_n9047 | 1_n12231);
assign 1_n11342 = 1_n11842 & 1_n10197;
assign 1_n722 = ~(1_n10007 ^ 1_n9337);
assign 1_n357 = 1_n9927 | 1_n10493;
assign 1_n9798 = ~(1_n4930 ^ 1_n3070);
assign 1_n6461 = ~(1_n9610 ^ 1_n6456);
assign 1_n9210 = ~(1_n13150 ^ 1_n2396);
assign 1_n2113 = ~(1_n5699 ^ 1_n3604);
assign 1_n209 = ~1_n7888;
assign 1_n7931 = 1_n10043 | 1_n2675;
assign 1_n616 = ~(1_n4263 | 1_n1649);
assign 1_n4758 = 1_n4382 & 1_n12284;
assign 1_n7029 = 1_n11311 | 1_n5712;
assign 1_n5960 = ~(1_n1041 ^ 1_n10910);
assign 1_n3749 = 1_n6220 | 1_n894;
assign 1_n7186 = ~(1_n600 | 1_n12425);
assign 1_n12746 = 1_n860 ^ 1_n5393;
assign 1_n10843 = 1_n9513 & 1_n1400;
assign 1_n8782 = ~(1_n11589 ^ 1_n6312);
assign 1_n6356 = ~(1_n9025 | 1_n11374);
assign 1_n3705 = ~(1_n7320 ^ 1_n8267);
assign 1_n569 = ~1_n2758;
assign 1_n7199 = ~1_n2787;
assign 1_n946 = ~1_n5427;
assign 1_n6939 = ~1_n4330;
assign 1_n10464 = ~(1_n5537 ^ 1_n11629);
assign 1_n11596 = 1_n8801 | 1_n4644;
assign 1_n7728 = 1_n875 & 1_n4509;
assign 1_n3797 = 1_n10757 & 1_n467;
assign 1_n623 = 1_n6326 | 1_n12543;
assign 1_n1940 = 1_n2048 | 1_n9682;
assign 1_n5287 = 1_n778 & 1_n10704;
assign 1_n7446 = 1_n10472 & 1_n12172;
assign 1_n7434 = 1_n4037 | 1_n7495;
assign 1_n4168 = ~(1_n13163 ^ 1_n5143);
assign 1_n4197 = ~(1_n12455 | 1_n12161);
assign 1_n12162 = 1_n6721 | 1_n5076;
assign 1_n592 = ~(1_n3541 ^ 1_n2587);
assign 1_n7031 = 1_n12362 | 1_n3987;
assign 1_n4268 = 1_n10780 | 1_n8268;
assign 1_n3629 = ~(1_n2739 | 1_n9232);
assign 1_n5038 = 1_n11640 ^ 1_n3830;
assign 1_n11553 = 1_n338 | 1_n2544;
assign 1_n8402 = 1_n9238 | 1_n12166;
assign 1_n12856 = ~1_n1369;
assign 1_n439 = ~(1_n8815 ^ 1_n7622);
assign 1_n3532 = 1_n2899 | 1_n1570;
assign 1_n11799 = ~1_n10033;
assign 1_n4101 = ~(1_n7181 ^ 1_n13103);
assign 1_n5414 = ~1_n10770;
assign 1_n2998 = ~(1_n9022 | 1_n10038);
assign 1_n10067 = ~(1_n4695 ^ 1_n9504);
assign 1_n10513 = 1_n1436 | 1_n9159;
assign 1_n3707 = ~(1_n2149 ^ 1_n2085);
assign 1_n2620 = ~(1_n108 ^ 1_n2892);
assign 1_n6561 = ~(1_n4513 ^ 1_n9267);
assign 1_n8476 = ~(1_n11321 ^ 1_n748);
assign 1_n13184 = 1_n1258 & 1_n4971;
assign 1_n8721 = 1_n1025 ^ 1_n8760;
assign 1_n455 = ~(1_n1904 ^ 1_n6974);
assign 1_n6788 = ~(1_n631 ^ 1_n11724);
assign 1_n1487 = 1_n8253 ^ 1_n7584;
assign 1_n10920 = 1_n13170 | 1_n6404;
assign 1_n10261 = 1_n13012 | 1_n1985;
assign 1_n7017 = 1_n860 | 1_n8371;
assign 1_n921 = 1_n13194 | 1_n4947;
assign 1_n6257 = 1_n8894 & 1_n5898;
assign 1_n12770 = 1_n1892 | 1_n1679;
assign 1_n44 = ~1_n11109;
assign 1_n2761 = ~(1_n4153 ^ 1_n7032);
assign 1_n2359 = 1_n808 | 1_n4621;
assign 1_n9541 = ~(1_n10571 ^ 1_n3798);
assign 1_n6212 = 1_n6182 | 1_n2059;
assign 1_n7045 = ~1_n6610;
assign 1_n2344 = ~(1_n7705 | 1_n5239);
assign 1_n11714 = 1_n1883 | 1_n6404;
assign 1_n2076 = 1_n1451 | 1_n2059;
assign 1_n9848 = 1_n234 | 1_n3843;
assign 1_n7843 = 1_n6768 | 1_n4455;
assign 1_n4258 = ~1_n499;
assign 1_n1175 = ~1_n5845;
assign 1_n7911 = 1_n2238 | 1_n9586;
assign 1_n11948 = ~(1_n2301 ^ 1_n7524);
assign 1_n11444 = ~(1_n7797 ^ 1_n7525);
assign 1_n12081 = ~(1_n12230 ^ 1_n9542);
assign 1_n11587 = ~(1_n5640 ^ 1_n9746);
assign 1_n12317 = ~(1_n550 | 1_n6594);
assign 1_n11406 = ~(1_n8758 ^ 1_n2629);
assign 1_n9771 = ~(1_n2820 ^ 1_n4646);
assign 1_n12520 = 1_n7591 & 1_n4547;
assign 1_n431 = 1_n4782 & 1_n12793;
assign 1_n4665 = ~1_n5884;
assign 1_n574 = ~(1_n1759 | 1_n11382);
assign 1_n3652 = ~1_n3203;
assign 1_n4946 = ~(1_n3251 ^ 1_n8686);
assign 1_n12676 = 1_n6166 | 1_n9195;
assign 1_n5868 = ~(1_n7317 ^ 1_n3261);
assign 1_n9319 = 1_n3914 & 1_n8017;
assign 1_n1335 = ~1_n5969;
assign 1_n9597 = 1_n11087 | 1_n542;
assign 1_n2668 = 1_n66 & 1_n4111;
assign 1_n4119 = ~(1_n4814 ^ 1_n2891);
assign 1_n12135 = 1_n4741 | 1_n177;
assign 1_n3140 = ~(1_n12399 ^ 1_n10706);
assign 1_n3867 = ~1_n11647;
assign 1_n5886 = ~(1_n296 ^ 1_n1083);
assign 1_n1481 = ~(1_n11909 ^ 1_n4125);
assign 1_n3944 = 1_n1897 | 1_n1832;
assign 1_n6015 = ~1_n11482;
assign 1_n10292 = ~1_n3358;
assign 1_n7905 = ~(1_n12486 ^ 1_n892);
assign 1_n6297 = ~(1_n3000 ^ 1_n5751);
assign 1_n13095 = ~(1_n6517 ^ 1_n6493);
assign 1_n8981 = 1_n448 & 1_n10345;
assign 1_n2636 = ~1_n4460;
assign 1_n9491 = ~(1_n3271 | 1_n10677);
assign 1_n4124 = ~(1_n9437 | 1_n779);
assign 1_n3165 = ~1_n2569;
assign 1_n3315 = 1_n6224 | 1_n7186;
assign 1_n4087 = ~1_n3251;
assign 1_n3795 = 1_n11505 | 1_n2367;
assign 1_n12386 = ~(1_n5687 ^ 1_n3300);
assign 1_n1632 = ~1_n8222;
assign 1_n9548 = ~(1_n5220 | 1_n11636);
assign 1_n12899 = ~1_n6783;
assign 1_n12255 = 1_n2592 & 1_n8860;
assign 1_n4863 = 1_n1737 | 1_n8534;
assign 1_n9893 = ~1_n42;
assign 1_n65 = 1_n4598 & 1_n5843;
assign 1_n7806 = ~(1_n2834 ^ 1_n5298);
assign 1_n8065 = ~1_n7309;
assign 1_n10998 = ~1_n9087;
assign 1_n11147 = ~(1_n4315 ^ 1_n12278);
assign 1_n6253 = 1_n558 & 1_n9294;
assign 1_n668 = 1_n6419 | 1_n8030;
assign 1_n3628 = ~(1_n6771 ^ 1_n7268);
assign 1_n6746 = 1_n6919 & 1_n1559;
assign 1_n1805 = 1_n5401 | 1_n617;
assign 1_n2052 = ~(1_n13128 ^ 1_n12609);
assign 1_n12371 = ~1_n6312;
assign 1_n6800 = 1_n5323 & 1_n4094;
assign 1_n1019 = 1_n8058 & 1_n2285;
assign 1_n7622 = 1_n1571 | 1_n2675;
assign 1_n2461 = ~(1_n4332 | 1_n11200);
assign 1_n8025 = 1_n2475 & 1_n6513;
assign 1_n4717 = 1_n2352 | 1_n7049;
assign 1_n4362 = 1_n9711 | 1_n9195;
assign 1_n8301 = ~1_n5729;
assign 1_n7442 = 1_n4428 & 1_n786;
assign 1_n476 = 1_n12653 | 1_n3884;
assign 1_n2980 = 1_n8306 | 1_n8563;
assign 1_n11793 = 1_n11920 | 1_n8348;
assign 1_n4855 = ~1_n443;
assign 1_n4029 = 1_n10991 | 1_n7723;
assign 1_n11544 = ~1_n12115;
assign 1_n6661 = ~(1_n2986 ^ 1_n7744);
assign 1_n12612 = 1_n8940 & 1_n7720;
assign 1_n7327 = 1_n13031 & 1_n9399;
assign 1_n8088 = 1_n11150 | 1_n2034;
assign 1_n2256 = ~(1_n3430 ^ 1_n7557);
assign 1_n5810 = ~(1_n1213 ^ 1_n8886);
assign 1_n8667 = ~(1_n11958 ^ 1_n3469);
assign 1_n10025 = 1_n5243 & 1_n10234;
assign 1_n6804 = ~(1_n8930 | 1_n8103);
assign 1_n4576 = 1_n6333 & 1_n2295;
assign 1_n1897 = ~1_n3964;
assign 1_n9980 = 1_n5448 | 1_n5487;
assign 1_n3410 = ~(1_n4050 ^ 1_n5305);
assign 1_n1185 = 1_n12671 | 1_n5242;
assign 1_n914 = 1_n11854 & 1_n8644;
assign 1_n12154 = ~(1_n7646 ^ 1_n1464);
assign 1_n4175 = 1_n2771 & 1_n2758;
assign 1_n11370 = ~1_n3591;
assign 1_n6088 = 1_n3157 | 1_n10471;
assign 1_n7272 = ~1_n9336;
assign 1_n2764 = 1_n4792 | 1_n10573;
assign 1_n48 = ~1_n12284;
assign 1_n8840 = ~1_n10622;
assign 1_n4833 = ~(1_n11838 ^ 1_n9296);
assign 1_n3951 = 1_n3062 | 1_n6769;
assign 1_n4582 = 1_n9129 | 1_n3459;
assign 1_n5336 = 1_n4363 & 1_n12888;
assign 1_n11391 = 1_n12964 | 1_n2679;
assign 1_n2533 = 1_n10465 | 1_n4949;
assign 1_n8781 = ~(1_n10743 | 1_n3399);
assign 1_n577 = ~(1_n1787 ^ 1_n10399);
assign 1_n5081 = ~(1_n5993 ^ 1_n1298);
assign 1_n4445 = 1_n11612 | 1_n12328;
assign 1_n9511 = ~1_n287;
assign 1_n8214 = ~(1_n11382 ^ 1_n1759);
assign 1_n2612 = ~(1_n11909 | 1_n10595);
assign 1_n12920 = 1_n2729 | 1_n76;
assign 1_n811 = ~(1_n3540 ^ 1_n7909);
assign 1_n11753 = 1_n5966 & 1_n8257;
assign 1_n11982 = ~1_n3130;
assign 1_n6482 = ~1_n170;
assign 1_n8273 = ~(1_n13139 ^ 1_n4318);
assign 1_n5435 = 1_n9891 | 1_n6973;
assign 1_n4698 = ~1_n948;
assign 1_n6151 = 1_n1674 & 1_n5274;
assign 1_n6663 = 1_n8211 & 1_n6111;
assign 1_n10505 = ~(1_n302 ^ 1_n2300);
assign 1_n9142 = ~(1_n12457 ^ 1_n3449);
assign 1_n2975 = ~1_n446;
assign 1_n2493 = ~1_n12219;
assign 1_n9441 = 1_n1887 | 1_n6635;
assign 1_n4275 = 1_n3537 | 1_n8490;
assign 1_n11100 = 1_n3344 | 1_n6635;
assign 1_n5950 = ~(1_n5738 | 1_n11403);
assign 1_n8580 = ~1_n10276;
assign 1_n5823 = 1_n12581 | 1_n5836;
assign 1_n3384 = ~1_n2798;
assign 1_n1223 = 1_n6758 & 1_n5930;
assign 1_n8748 = ~(1_n502 | 1_n3319);
assign 1_n7202 = 1_n13051 | 1_n8383;
assign 1_n9337 = ~(1_n9388 | 1_n7520);
assign 1_n5636 = 1_n7798 | 1_n2133;
assign 1_n12971 = 1_n6841 | 1_n11609;
assign 1_n311 = 1_n4927 | 1_n11100;
assign 1_n5400 = ~1_n10504;
assign 1_n11468 = ~1_n1742;
assign 1_n5905 = ~1_n5083;
assign 1_n7981 = ~(1_n2081 | 1_n12810);
assign 1_n12019 = ~1_n9585;
assign 1_n5795 = 1_n5713 | 1_n1463;
assign 1_n6122 = ~(1_n5300 ^ 1_n3125);
assign 1_n7079 = ~(1_n6605 ^ 1_n6020);
assign 1_n1792 = 1_n1677 & 1_n9814;
assign 1_n9239 = 1_n11061 & 1_n287;
assign 1_n5915 = ~1_n9833;
assign 1_n7050 = ~(1_n10420 ^ 1_n7466);
assign 1_n2600 = ~1_n1254;
assign 1_n1857 = ~1_n1110;
assign 1_n6280 = 1_n12213 & 1_n6045;
assign 1_n7814 = ~1_n7537;
assign 1_n7210 = 1_n10400 | 1_n4724;
assign 1_n7109 = 1_n11262 | 1_n2992;
assign 1_n3801 = ~(1_n5805 | 1_n9786);
assign 1_n3841 = ~(1_n7153 ^ 1_n13166);
assign 1_n9501 = ~(1_n8369 | 1_n3286);
assign 1_n5429 = ~(1_n7085 ^ 1_n1266);
assign 1_n11233 = ~(1_n13236 ^ 1_n4734);
assign 1_n5053 = ~(1_n7938 | 1_n11204);
assign 1_n11035 = 1_n12052 | 1_n4253;
assign 1_n2216 = ~(1_n7183 ^ 1_n6604);
assign 1_n4847 = 1_n1498 ^ 1_n9623;
assign 1_n2972 = 1_n1135 | 1_n5264;
assign 1_n9490 = ~1_n6892;
assign 1_n11025 = ~(1_n3273 ^ 1_n1780);
assign 1_n2507 = 1_n6603 | 1_n362;
assign 1_n6508 = 1_n8646 | 1_n6732;
assign 1_n3426 = ~(1_n7210 ^ 1_n12499);
assign 1_n12768 = ~1_n3085;
assign 1_n1457 = 1_n4022 | 1_n4936;
assign 1_n11 = 1_n4041 | 1_n12404;
assign 1_n12724 = 1_n6684 & 1_n2971;
assign 1_n3916 = 1_n7522 | 1_n3703;
assign 1_n407 = ~1_n7294;
assign 1_n1001 = 1_n5503 | 1_n1452;
assign 1_n10966 = ~1_n6085;
assign 1_n11904 = ~(1_n7271 ^ 1_n8618);
assign 1_n8086 = ~(1_n3765 | 1_n10734);
assign 1_n4956 = ~(1_n3278 | 1_n12385);
assign 1_n12303 = ~1_n1195;
assign 1_n8871 = 1_n8995 | 1_n7863;
assign 1_n4596 = ~(1_n9058 ^ 1_n4687);
assign 1_n6920 = 1_n10770 & 1_n8233;
assign 1_n902 = ~1_n8230;
assign 1_n1945 = ~1_n10671;
assign 1_n6537 = 1_n7076 | 1_n9223;
assign 1_n12553 = ~(1_n12168 ^ 1_n904);
assign 1_n4519 = 1_n12481 & 1_n8750;
assign 1_n5607 = ~1_n3357;
assign 1_n5900 = 1_n11629 | 1_n7768;
assign 1_n4995 = 1_n1451 | 1_n121;
assign 1_n8832 = 1_n10714 | 1_n10474;
assign 1_n8325 = ~1_n4122;
assign 1_n9404 = ~(1_n13240 ^ 1_n7285);
assign 1_n12071 = 1_n2646 | 1_n9381;
assign 1_n12557 = 1_n542 | 1_n8702;
assign 1_n1374 = ~(1_n3931 ^ 1_n1790);
assign 1_n6651 = 1_n69 | 1_n8534;
assign 1_n9788 = ~1_n12692;
assign 1_n11421 = 1_n4403 & 1_n1828;
assign 1_n7499 = ~(1_n11478 ^ 1_n12208);
assign 1_n12800 = 1_n4334 & 1_n1777;
assign 1_n9786 = ~1_n5868;
assign 1_n3023 = 1_n10845 & 1_n200;
assign 1_n10296 = ~(1_n6615 | 1_n450);
assign 1_n10547 = 1_n6120 & 1_n4783;
assign 1_n376 = 1_n12099 & 1_n11866;
assign 1_n7910 = ~(1_n8161 ^ 1_n38);
assign 1_n3637 = 1_n2109 | 1_n2726;
assign 1_n3500 = 1_n11849 & 1_n3778;
assign 1_n12777 = 1_n9400 | 1_n11107;
assign 1_n7507 = ~(1_n6445 | 1_n3845);
assign 1_n5692 = ~1_n6068;
assign 1_n8255 = 1_n5535 | 1_n9847;
assign 1_n4917 = ~(1_n9487 ^ 1_n4870);
assign 1_n9793 = ~1_n11734;
assign 1_n255 = 1_n7473 | 1_n196;
assign 1_n10386 = 1_n2710 | 1_n1871;
assign 1_n3734 = ~(1_n5961 ^ 1_n8190);
assign 1_n5739 = 1_n7484 & 1_n3848;
assign 1_n1619 = ~(1_n3193 ^ 1_n5803);
assign 1_n6194 = ~1_n9343;
assign 1_n3380 = ~1_n2597;
assign 1_n1243 = ~(1_n3150 | 1_n6839);
assign 1_n1276 = ~(1_n7592 ^ 1_n11299);
assign 1_n12399 = ~(1_n2103 | 1_n12325);
assign 1_n174 = 1_n9588 | 1_n10708;
assign 1_n4113 = 1_n9736 & 1_n10667;
assign 1_n11483 = ~(1_n11233 | 1_n12498);
assign 1_n5633 = 1_n11235 | 1_n6113;
assign 1_n894 = ~1_n12853;
assign 1_n3541 = ~(1_n1839 ^ 1_n11409);
assign 1_n2884 = ~1_n497;
assign 1_n3030 = 1_n2484 | 1_n8383;
assign 1_n9831 = 1_n9283 & 1_n7220;
assign 1_n4522 = ~1_n11434;
assign 1_n12418 = 1_n4028 & 1_n6851;
assign 1_n1517 = ~(1_n13185 | 1_n10309);
assign 1_n9526 = ~(1_n6898 | 1_n6027);
assign 1_n3846 = 1_n7827 & 1_n10549;
assign 1_n2816 = ~1_n10642;
assign 1_n4301 = ~1_n6639;
assign 1_n12936 = ~(1_n10593 ^ 1_n5576);
assign 1_n12828 = 1_n1982 & 1_n11488;
assign 1_n11428 = ~(1_n4995 ^ 1_n7551);
assign 1_n12860 = ~(1_n4711 | 1_n10787);
assign 1_n6470 = ~(1_n7745 ^ 1_n3844);
assign 1_n705 = 1_n564 & 1_n9596;
assign 1_n900 = ~(1_n8947 | 1_n12176);
assign 1_n13123 = 1_n12432 | 1_n3417;
assign 1_n8632 = ~1_n6668;
assign 1_n4575 = 1_n9426 | 1_n3053;
assign 1_n6653 = 1_n798 & 1_n8331;
assign 1_n12240 = ~1_n3472;
assign 1_n216 = 1_n1472 ^ 1_n2652;
assign 1_n8809 = ~1_n10126;
assign 1_n5902 = ~(1_n6401 ^ 1_n9798);
assign 1_n6376 = 1_n6131 | 1_n9757;
assign 1_n4317 = 1_n13154 | 1_n12273;
assign 1_n10110 = 1_n2183 | 1_n6635;
assign 1_n2815 = ~(1_n6248 | 1_n8968);
assign 1_n10293 = ~1_n6536;
assign 1_n10975 = ~1_n9616;
assign 1_n5570 = ~(1_n3002 ^ 1_n8698);
assign 1_n712 = ~1_n865;
assign 1_n9582 = 1_n8502 & 1_n5720;
assign 1_n2434 = 1_n1447 | 1_n206;
assign 1_n10165 = 1_n6847 & 1_n8994;
assign 1_n6992 = 1_n8169 | 1_n10407;
assign 1_n12209 = ~(1_n10110 ^ 1_n11195);
assign 1_n2384 = ~(1_n5013 ^ 1_n12238);
assign 1_n8662 = 1_n8280 | 1_n11016;
assign 1_n2046 = 1_n10421 | 1_n7935;
assign 1_n11967 = 1_n10469 | 1_n4404;
assign 1_n1754 = 1_n9424 & 1_n6619;
assign 1_n11677 = ~1_n6765;
assign 1_n6791 = 1_n8236 & 1_n3184;
assign 1_n13147 = 1_n6668 & 1_n5729;
assign 1_n11892 = ~(1_n8316 ^ 1_n12353);
assign 1_n100 = 1_n444 | 1_n3383;
assign 1_n6056 = ~1_n10142;
assign 1_n12635 = 1_n8436 | 1_n1155;
assign 1_n6038 = 1_n4513 & 1_n3309;
assign 1_n12540 = ~(1_n6354 ^ 1_n8707);
assign 1_n5742 = ~1_n4348;
assign 1_n10124 = ~(1_n4048 ^ 1_n827);
assign 1_n11670 = 1_n3304 & 1_n4916;
assign 1_n3590 = ~(1_n11925 | 1_n11342);
assign 1_n161 = ~1_n7974;
assign 1_n4510 = ~(1_n2036 ^ 1_n5925);
assign 1_n6918 = 1_n8294 | 1_n10685;
assign 1_n2523 = 1_n5105 | 1_n11772;
assign 1_n1908 = ~1_n11454;
assign 1_n12854 = 1_n4975 & 1_n10520;
assign 1_n10854 = ~(1_n10933 | 1_n10799);
assign 1_n3451 = ~(1_n10405 ^ 1_n7393);
assign 1_n2738 = ~1_n3815;
assign 1_n10795 = ~1_n10002;
assign 1_n12737 = 1_n11810 | 1_n8268;
assign 1_n6849 = ~(1_n10356 | 1_n8809);
assign 1_n1688 = ~1_n8522;
assign 1_n2521 = ~(1_n2826 | 1_n10965);
assign 1_n1242 = 1_n7907 & 1_n10108;
assign 1_n9993 = 1_n1364 & 1_n124;
assign 1_n3943 = ~(1_n10273 | 1_n5198);
assign 1_n8547 = 1_n6399 | 1_n5063;
assign 1_n12032 = ~1_n817;
assign 1_n6278 = 1_n3926 & 1_n11203;
assign 1_n1814 = 1_n8707 & 1_n6354;
assign 1_n8460 = 1_n11457 | 1_n5349;
assign 1_n9766 = ~(1_n9881 ^ 1_n1740);
assign 1_n9262 = ~(1_n12181 ^ 1_n12130);
assign 1_n11838 = ~1_n4312;
assign 1_n4245 = 1_n2763 & 1_n9366;
assign 1_n8953 = ~(1_n2465 ^ 1_n11615);
assign 1_n8796 = ~(1_n4685 | 1_n1045);
assign 1_n13073 = ~1_n7982;
assign 1_n12196 = 1_n4731 | 1_n210;
assign 1_n1425 = ~(1_n10857 ^ 1_n4577);
assign 1_n5553 = ~(1_n9895 ^ 1_n384);
assign 1_n8421 = 1_n8450 | 1_n5669;
assign 1_n8329 = ~1_n6843;
assign 1_n2772 = ~1_n6822;
assign 1_n11089 = ~(1_n7901 ^ 1_n8955);
assign 1_n7048 = ~(1_n1766 | 1_n1358);
assign 1_n9639 = 1_n13201 & 1_n5548;
assign 1_n9294 = ~(1_n6636 ^ 1_n1660);
assign 1_n8842 = ~(1_n7842 ^ 1_n6147);
assign 1_n11847 = 1_n6229 | 1_n1417;
assign 1_n6267 = ~1_n1203;
assign 1_n3300 = 1_n4612 | 1_n3949;
assign 1_n12597 = 1_n8356 | 1_n8918;
assign 1_n8136 = ~(1_n6535 ^ 1_n4064);
assign 1_n8226 = 1_n240 & 1_n8734;
assign 1_n9057 = ~(1_n6478 | 1_n11678);
assign 1_n8823 = ~(1_n4571 ^ 1_n3823);
assign 1_n5910 = ~(1_n3561 | 1_n12830);
assign 1_n652 = ~1_n9093;
assign 1_n9375 = ~1_n3876;
assign 1_n8297 = ~1_n10728;
assign 1_n3272 = ~(1_n11570 | 1_n4239);
assign 1_n348 = ~(1_n8539 ^ 1_n2293);
assign 1_n64 = ~1_n6087;
assign 1_n9303 = 1_n10113 & 1_n10451;
assign 1_n2122 = ~1_n8399;
assign 1_n9010 = ~1_n469;
assign 1_n4858 = ~(1_n9959 ^ 1_n8896);
assign 1_n688 = ~(1_n10327 | 1_n6711);
assign 1_n10215 = 1_n9748 & 1_n12895;
assign 1_n1182 = ~(1_n7934 ^ 1_n289);
assign 1_n110 = 1_n9273 | 1_n9686;
assign 1_n10072 = ~(1_n11930 | 1_n3924);
assign 1_n4770 = 1_n10872 & 1_n12308;
assign 1_n7208 = 1_n828 ^ 1_n5483;
assign 1_n1190 = 1_n1952 & 1_n2601;
assign 1_n9273 = 1_n2496 & 1_n4988;
assign 1_n5802 = ~1_n1874;
assign 1_n12370 = ~1_n6897;
assign 1_n4525 = 1_n9917 | 1_n10049;
assign 1_n1562 = 1_n7794 | 1_n7563;
assign 1_n10532 = 1_n626 & 1_n7887;
assign 1_n6306 = ~1_n2590;
assign 1_n9182 = ~1_n11280;
assign 1_n1823 = 1_n10984 & 1_n3404;
assign 1_n118 = ~1_n13192;
assign 1_n12029 = 1_n1259 & 1_n297;
assign 1_n6058 = 1_n2604 & 1_n12358;
assign 1_n5180 = 1_n7146 | 1_n5076;
assign 1_n2454 = ~(1_n1517 ^ 1_n430);
assign 1_n3237 = ~(1_n10643 | 1_n3633);
assign 1_n2794 = 1_n9788 & 1_n9989;
assign 1_n12410 = ~(1_n3321 ^ 1_n10190);
assign 1_n8058 = ~1_n5304;
assign 1_n851 = 1_n5491 & 1_n10171;
assign 1_n6579 = ~1_n6226;
assign 1_n7339 = 1_n4608 & 1_n1918;
assign 1_n12170 = ~1_n7813;
assign 1_n5004 = 1_n1436 | 1_n4640;
assign 1_n11900 = 1_n12033 | 1_n4416;
assign 1_n1833 = 1_n13112 & 1_n12851;
assign 1_n9840 = ~(1_n12528 ^ 1_n2694);
assign 1_n11760 = 1_n2003 & 1_n9237;
assign 1_n12880 = ~(1_n1896 | 1_n11005);
assign 1_n6754 = ~(1_n8272 ^ 1_n11062);
assign 1_n701 = 1_n3682 | 1_n7013;
assign 1_n7402 = ~(1_n10444 | 1_n8586);
assign 1_n4171 = 1_n7969 ^ 1_n6433;
assign 1_n12463 = ~(1_n1192 ^ 1_n13029);
assign 1_n3283 = ~(1_n9067 ^ 1_n7341);
assign 1_n11560 = 1_n7247 | 1_n2228;
assign 1_n11740 = ~1_n8358;
assign 1_n11431 = ~1_n12428;
assign 1_n10893 = ~1_n2758;
assign 1_n7502 = 1_n11322 & 1_n11662;
assign 1_n6486 = ~1_n1231;
assign 1_n4225 = 1_n6051 | 1_n11998;
assign 1_n8980 = 1_n7052 & 1_n2219;
assign 1_n4957 = 1_n2540 ^ 1_n9013;
assign 1_n4999 = ~(1_n3909 ^ 1_n698);
assign 1_n12995 = ~1_n441;
assign 1_n1729 = 1_n12551 | 1_n5781;
assign 1_n4334 = 1_n12997 | 1_n2133;
assign 1_n8641 = ~(1_n9734 | 1_n8523);
assign 1_n4446 = 1_n3416 | 1_n4474;
assign 1_n2399 = ~(1_n668 | 1_n6663);
assign 1_n3539 = 1_n5656 | 1_n11538;
assign 1_n3671 = ~1_n5684;
assign 1_n11869 = ~1_n6515;
assign 1_n699 = ~(1_n11859 ^ 1_n6877);
assign 1_n7421 = ~1_n4572;
assign 1_n7071 = ~(1_n374 | 1_n5225);
assign 1_n12454 = ~(1_n5509 | 1_n12875);
assign 1_n1008 = ~1_n8932;
assign 1_n10648 = ~(1_n2973 ^ 1_n5646);
assign 1_n12656 = 1_n559 | 1_n4947;
assign 1_n11197 = 1_n12602 | 1_n3902;
assign 1_n7111 = ~(1_n2212 ^ 1_n9768);
assign 1_n13182 = ~1_n9669;
assign 1_n10052 = 1_n9172 & 1_n4231;
assign 1_n3294 = 1_n6744 & 1_n347;
assign 1_n8398 = ~(1_n5530 ^ 1_n2138);
assign 1_n1568 = ~(1_n5636 ^ 1_n152);
assign 1_n1489 = ~(1_n1657 ^ 1_n2828);
assign 1_n9336 = ~(1_n1465 ^ 1_n12973);
assign 1_n2237 = ~(1_n12897 ^ 1_n10216);
assign 1_n11565 = 1_n10908 & 1_n854;
assign 1_n12320 = 1_n5964 & 1_n2270;
assign 1_n4191 = 1_n2937 & 1_n10812;
assign 1_n11632 = 1_n10809 & 1_n4342;
assign 1_n5701 = ~(1_n2474 ^ 1_n12017);
assign 1_n7465 = ~(1_n3024 ^ 1_n2119);
assign 1_n368 = ~(1_n12410 ^ 1_n1027);
assign 1_n259 = 1_n2806 & 1_n2189;
assign 1_n2479 = 1_n4792 | 1_n3454;
assign 1_n3875 = ~(1_n12269 ^ 1_n1519);
assign 1_n12554 = ~(1_n10450 ^ 1_n5201);
assign 1_n2550 = ~1_n471;
assign 1_n5281 = ~(1_n10806 ^ 1_n5977);
assign 1_n11448 = ~(1_n282 ^ 1_n8916);
assign 1_n4125 = ~(1_n3869 ^ 1_n8717);
assign 1_n7537 = 1_n4370 | 1_n6635;
assign 1_n346 = 1_n1647 & 1_n4402;
assign 1_n12705 = 1_n3024 | 1_n2119;
assign 1_n12070 = 1_n9968 | 1_n9850;
assign 1_n10912 = 1_n628 | 1_n10106;
assign 1_n4010 = 1_n11664 | 1_n9795;
assign 1_n4235 = 1_n12093 | 1_n12847;
assign 1_n5623 = 1_n7538 & 1_n2782;
assign 1_n6811 = ~1_n4387;
assign 1_n8734 = 1_n4251 | 1_n3079;
assign 1_n10183 = 1_n8053 | 1_n2675;
assign 1_n10051 = ~1_n3298;
assign 1_n8338 = ~(1_n1375 | 1_n12097);
assign 1_n1372 = 1_n6904 | 1_n5915;
assign 1_n3555 = ~1_n9188;
assign 1_n4492 = 1_n11318 & 1_n8880;
assign 1_n12900 = 1_n5252 & 1_n2573;
assign 1_n7599 = ~(1_n11193 ^ 1_n6705);
assign 1_n8415 = ~(1_n9790 | 1_n10831);
assign 1_n7722 = 1_n6333 & 1_n834;
assign 1_n9622 = ~1_n6392;
assign 1_n728 = ~(1_n3271 ^ 1_n1776);
assign 1_n5129 = 1_n8969 | 1_n9141;
assign 1_n228 = ~(1_n5725 ^ 1_n5928);
assign 1_n10763 = ~(1_n149 ^ 1_n6773);
assign 1_n6784 = ~(1_n4359 ^ 1_n12775);
assign 1_n4104 = 1_n1567 | 1_n12400;
assign 1_n1048 = 1_n9675 | 1_n6265;
assign 1_n12199 = ~(1_n8891 ^ 1_n3182);
assign 1_n1158 = 1_n3225 | 1_n6265;
assign 1_n9537 = ~1_n11324;
assign 1_n2388 = 1_n4732 | 1_n4230;
assign 1_n12173 = ~(1_n4000 ^ 1_n8477);
assign 1_n7542 = 1_n11087 | 1_n2449;
assign 1_n7184 = ~1_n12579;
assign 1_n5589 = 1_n7085 | 1_n1781;
assign 1_n587 = ~(1_n6572 ^ 1_n6546);
assign 1_n11452 = ~1_n5174;
assign 1_n9366 = 1_n11335 | 1_n2123;
assign 1_n13087 = 1_n13243 & 1_n7003;
assign 1_n9572 = 1_n12877 & 1_n12288;
assign 1_n7548 = ~(1_n10477 | 1_n8965);
assign 1_n2449 = 1_n10240;
assign 1_n5386 = ~(1_n6887 ^ 1_n13024);
assign 1_n4108 = 1_n13117 | 1_n10871;
assign 1_n9905 = 1_n420 & 1_n1798;
assign 1_n575 = 1_n8067 & 1_n10817;
assign 1_n11909 = 1_n334 | 1_n12948;
assign 1_n8972 = 1_n10761 | 1_n1570;
assign 1_n9203 = 1_n4099 & 1_n10691;
assign 1_n5526 = 1_n2195 | 1_n3523;
assign 1_n11135 = ~(1_n6195 | 1_n1900);
assign 1_n9610 = ~(1_n2992 ^ 1_n1336);
assign 1_n6377 = 1_n8688 & 1_n548;
assign 1_n8453 = ~1_n7165;
assign 1_n13138 = 1_n10756 | 1_n9195;
assign 1_n10001 = ~(1_n3822 ^ 1_n1613);
assign 1_n2092 = 1_n7339 & 1_n5695;
assign 1_n11644 = ~(1_n11881 | 1_n9535);
assign 1_n7968 = 1_n9705 ^ 1_n12101;
assign 1_n10341 = 1_n1113 | 1_n1144;
assign 1_n5609 = ~(1_n5914 ^ 1_n12729);
assign 1_n10239 = ~(1_n279 | 1_n11338);
assign 1_n4694 = ~1_n1543;
assign 1_n3653 = 1_n6188 & 1_n12922;
assign 1_n1996 = 1_n5711 & 1_n5085;
assign 1_n301 = ~(1_n1617 ^ 1_n5596);
assign 1_n5404 = ~(1_n528 ^ 1_n5870);
assign 1_n10356 = ~(1_n1553 ^ 1_n7964);
assign 1_n4589 = ~1_n6601;
assign 1_n1095 = ~(1_n4197 | 1_n4697);
assign 1_n3443 = 1_n11608 & 1_n7657;
assign 1_n1637 = ~(1_n2242 ^ 1_n9073);
assign 1_n9733 = 1_n1983 | 1_n6255;
assign 1_n9228 = ~1_n10162;
assign 1_n10757 = ~1_n2703;
assign 1_n8410 = 1_n9622 | 1_n4420;
assign 1_n2288 = ~(1_n6902 ^ 1_n10750);
assign 1_n2534 = 1_n7981 | 1_n6089;
assign 1_n8801 = 1_n2919 | 1_n12388;
assign 1_n9590 = 1_n6423 & 1_n593;
assign 1_n12689 = 1_n6206 | 1_n11097;
assign 1_n6313 = ~1_n11993;
assign 1_n7917 = 1_n5949 | 1_n6635;
assign 1_n10198 = ~1_n9943;
assign 1_n929 = 1_n4334 | 1_n1777;
assign 1_n2355 = 1_n8994 | 1_n6847;
assign 1_n5155 = 1_n4418 | 1_n6926;
assign 1_n12841 = ~1_n9475;
assign 1_n3019 = 1_n2162 & 1_n4678;
assign 1_n7936 = ~(1_n12085 ^ 1_n2071);
assign 1_n6428 = 1_n4809 | 1_n3632;
assign 1_n8967 = ~(1_n3625 ^ 1_n6871);
assign 1_n6527 = ~(1_n11743 | 1_n12727);
assign 1_n12622 = 1_n2266 & 1_n3743;
assign 1_n2993 = 1_n11120 | 1_n5885;
assign 1_n7708 = ~1_n7585;
assign 1_n8345 = ~(1_n1735 ^ 1_n10164);
assign 1_n12548 = 1_n12141 | 1_n10513;
assign 1_n4394 = ~(1_n5445 ^ 1_n5681);
assign 1_n4380 = ~(1_n10186 ^ 1_n8151);
assign 1_n3468 = ~1_n10150;
assign 1_n8803 = 1_n7128 ^ 1_n4078;
assign 1_n9027 = ~(1_n3833 ^ 1_n3754);
assign 1_n298 = 1_n3821 | 1_n12755;
assign 1_n4223 = 1_n5510 & 1_n5795;
assign 1_n4271 = ~(1_n5762 ^ 1_n2501);
assign 1_n9209 = ~1_n9843;
assign 1_n5315 = 1_n8668 & 1_n8381;
assign 1_n6536 = ~(1_n9831 ^ 1_n11025);
assign 1_n9900 = 1_n2613 | 1_n12233;
assign 1_n10031 = ~(1_n4713 | 1_n11441);
assign 1_n10431 = ~(1_n2167 | 1_n7535);
assign 1_n949 = 1_n7675 | 1_n9195;
assign 1_n10045 = ~1_n3076;
assign 1_n2683 = ~(1_n1400 ^ 1_n9513);
assign 1_n7976 = ~(1_n11131 | 1_n1137);
assign 1_n6162 = 1_n5867 & 1_n8088;
assign 1_n2907 = 1_n8816 & 1_n11999;
assign 1_n3587 = ~1_n1084;
assign 1_n3138 = ~(1_n1009 ^ 1_n3678);
assign 1_n5190 = 1_n2903 & 1_n8803;
assign 1_n4703 = 1_n11324 & 1_n1724;
assign 1_n11865 = ~(1_n8551 ^ 1_n1249);
assign 1_n7338 = ~(1_n11095 | 1_n6390);
assign 1_n2895 = ~(1_n1975 ^ 1_n356);
assign 1_n5989 = 1_n644 | 1_n542;
assign 1_n12820 = 1_n8600 ^ 1_n3137;
assign 1_n1643 = ~(1_n2817 | 1_n1299);
assign 1_n3004 = 1_n4313 | 1_n3487;
assign 1_n4012 = ~(1_n1223 | 1_n7673);
assign 1_n63 = ~1_n9531;
assign 1_n13093 = 1_n7276 & 1_n3106;
assign 1_n4866 = ~1_n2038;
assign 1_n5791 = 1_n5371 & 1_n3097;
assign 1_n3503 = ~(1_n1607 ^ 1_n2745);
assign 1_n5863 = 1_n3408 | 1_n11086;
assign 1_n12718 = ~1_n11537;
assign 1_n1210 = 1_n1072 | 1_n2851;
assign 1_n4940 = 1_n11269 | 1_n8196;
assign 1_n4205 = 1_n4612 | 1_n8563;
assign 1_n10572 = ~(1_n12419 ^ 1_n3196);
assign 1_n5416 = 1_n4668 | 1_n12726;
assign 1_n2968 = ~(1_n374 ^ 1_n11992);
assign 1_n4185 = ~1_n9887;
assign 1_n10712 = 1_n1571 | 1_n6265;
assign 1_n3673 = ~(1_n1752 | 1_n11106);
assign 1_n7001 = ~1_n8273;
assign 1_n11185 = ~1_n1278;
assign 1_n4296 = ~(1_n6118 ^ 1_n1229);
assign 1_n9230 = ~(1_n10412 ^ 1_n4031);
assign 1_n8990 = ~(1_n3874 | 1_n7198);
assign 1_n3729 = ~1_n7238;
assign 1_n8501 = ~(1_n8289 ^ 1_n1502);
assign 1_n1418 = 1_n9942 & 1_n890;
assign 1_n7621 = ~(1_n8632 | 1_n9913);
assign 1_n7774 = ~(1_n5642 ^ 1_n4422);
assign 1_n6372 = 1_n10761 | 1_n6404;
assign 1_n8685 = 1_n4878 & 1_n10141;
assign 1_n1704 = 1_n519 & 1_n11896;
assign 1_n9856 = ~(1_n5093 ^ 1_n2506);
assign 1_n11922 = ~1_n1923;
assign 1_n3710 = ~(1_n4192 ^ 1_n7114);
assign 1_n6373 = ~(1_n7101 ^ 1_n1132);
assign 1_n11415 = 1_n470 & 1_n8370;
assign 1_n8174 = ~1_n11835;
assign 1_n8604 = ~(1_n99 ^ 1_n10416);
assign 1_n309 = 1_n11876 & 1_n1657;
assign 1_n9781 = 1_n3478 | 1_n5537;
assign 1_n9829 = ~1_n3894;
assign 1_n12175 = 1_n8757 | 1_n6404;
assign 1_n4673 = 1_n1184 & 1_n11188;
assign 1_n4252 = 1_n959 ^ 1_n4758;
assign 1_n8448 = 1_n10448 | 1_n5076;
assign 1_n8625 = 1_n4208 | 1_n1144;
assign 1_n10396 = ~(1_n6651 ^ 1_n9657);
assign 1_n9128 = ~(1_n7581 ^ 1_n9973);
assign 1_n896 = 1_n9225 | 1_n3023;
assign 1_n7095 = 1_n5019 | 1_n6141;
assign 1_n4966 = ~(1_n1549 | 1_n5753);
assign 1_n472 = ~(1_n12133 ^ 1_n7595);
assign 1_n3848 = 1_n4272 | 1_n5797;
assign 1_n3806 = ~(1_n1178 ^ 1_n10489);
assign 1_n3592 = 1_n3096 | 1_n542;
assign 1_n6667 = 1_n1968 | 1_n12745;
assign 1_n2732 = 1_n1160 & 1_n2446;
assign 1_n7894 = 1_n9911 | 1_n1843;
assign 1_n1954 = ~1_n10398;
assign 1_n12148 = ~(1_n12172 ^ 1_n5223);
assign 1_n11582 = 1_n12904 & 1_n12427;
assign 1_n1139 = 1_n9901 & 1_n11801;
assign 1_n10129 = 1_n7934 | 1_n289;
assign 1_n11227 = ~1_n6868;
assign 1_n6161 = ~(1_n7978 ^ 1_n1129);
assign 1_n3376 = 1_n8873 & 1_n4804;
assign 1_n10085 = ~1_n5969;
assign 1_n4110 = 1_n2223 & 1_n4706;
assign 1_n10425 = ~1_n727;
assign 1_n4707 = 1_n9776 ^ 1_n4037;
assign 1_n10637 = 1_n2463 | 1_n10871;
assign 1_n5016 = ~1_n10563;
assign 1_n5328 = ~1_n9747;
assign 1_n9168 = 1_n5671 & 1_n3769;
assign 1_n1265 = 1_n13170 | 1_n12388;
assign 1_n7242 = ~1_n6195;
assign 1_n1660 = ~(1_n11272 ^ 1_n10087);
assign 1_n10479 = 1_n12673 & 1_n7761;
assign 1_n8083 = 1_n3647 & 1_n5098;
assign 1_n8147 = ~(1_n12389 ^ 1_n6138);
assign 1_n7426 = ~(1_n12817 ^ 1_n12872);
assign 1_n155 = 1_n652 | 1_n2544;
assign 1_n5887 = ~(1_n6425 | 1_n13091);
assign 1_n12502 = ~(1_n11392 ^ 1_n9760);
assign 1_n2229 = 1_n7715 & 1_n12306;
assign 1_n10927 = ~1_n5334;
assign 1_n10548 = ~(1_n9270 ^ 1_n2422);
assign 1_n6204 = 1_n8040 & 1_n7464;
assign 1_n12805 = 1_n10641 | 1_n11152;
assign 1_n8587 = 1_n5601 & 1_n10265;
assign 1_n4401 = 1_n6304 | 1_n539;
assign 1_n10819 = 1_n7609 & 1_n11924;
assign 1_n2648 = 1_n9464 & 1_n9191;
assign 1_n6158 = ~(1_n3526 ^ 1_n350);
assign 1_n6833 = 1_n5517 & 1_n12559;
assign 1_n303 = 1_n2091 | 1_n3597;
assign 1_n9079 = ~(1_n7406 ^ 1_n1182);
assign 1_n13240 = 1_n698 & 1_n3909;
assign 1_n6289 = ~(1_n6893 | 1_n948);
assign 1_n13230 = ~(1_n10496 ^ 1_n5159);
assign 1_n2425 = 1_n9089 | 1_n7760;
assign 1_n9305 = ~1_n5189;
assign 1_n11592 = ~(1_n3105 ^ 1_n6410);
assign 1_n3093 = ~(1_n7438 ^ 1_n3732);
assign 1_n10887 = ~(1_n7448 ^ 1_n194);
assign 1_n1024 = 1_n2057 & 1_n834;
assign 1_n8542 = 1_n8228 & 1_n411;
assign 1_n8951 = ~1_n486;
assign 1_n2532 = ~(1_n293 | 1_n7150);
assign 1_n11806 = ~1_n9376;
assign 1_n11243 = ~(1_n9365 ^ 1_n636);
assign 1_n9666 = 1_n7208 ^ 1_n11846;
assign 1_n4288 = 1_n3000 | 1_n9971;
assign 1_n12875 = 1_n4725 & 1_n2265;
assign 1_n10607 = 1_n8922 | 1_n5389;
assign 1_n2054 = ~(1_n8990 ^ 1_n3675);
assign 1_n11509 = ~1_n4441;
assign 1_n798 = ~(1_n217 ^ 1_n3889);
assign 1_n4091 = 1_n953 & 1_n8107;
assign 1_n10007 = ~(1_n1564 | 1_n512);
assign 1_n8729 = ~1_n7411;
assign 1_n6808 = ~1_n323;
assign 1_n12757 = ~(1_n9958 | 1_n3719);
assign 1_n9022 = ~(1_n12974 | 1_n11587);
assign 1_n2004 = ~(1_n3484 | 1_n13189);
assign 1_n8611 = ~(1_n11383 ^ 1_n8396);
assign 1_n4316 = 1_n5461 | 1_n2449;
assign 1_n648 = ~(1_n10568 ^ 1_n12520);
assign 1_n9438 = 1_n11370 | 1_n5797;
assign 1_n4521 = 1_n7626 | 1_n5340;
assign 1_n7522 = ~1_n2737;
assign 1_n13001 = 1_n5218 | 1_n496;
assign 1_n12721 = ~1_n3130;
assign 1_n12455 = 1_n18 | 1_n11668;
assign 1_n790 = 1_n7537 ^ 1_n3211;
assign 1_n9394 = ~(1_n9364 ^ 1_n10058);
assign 1_n5699 = ~(1_n11312 ^ 1_n7812);
assign 1_n11501 = 1_n11037 | 1_n2059;
assign 1_n5350 = 1_n12150 | 1_n4145;
assign 1_n13004 = ~(1_n5720 ^ 1_n8502);
assign 1_n4806 = ~(1_n9894 ^ 1_n5210);
assign 1_n3161 = ~(1_n4834 ^ 1_n11934);
assign 1_n2309 = ~(1_n8362 ^ 1_n4011);
assign 1_n4019 = ~(1_n4941 ^ 1_n2628);
assign 1_n9044 = 1_n6003 | 1_n10579;
assign 1_n9651 = ~1_n10709;
assign 1_n5373 = 1_n3557 & 1_n6742;
assign 1_n11923 = ~(1_n5778 ^ 1_n2381);
assign 1_n11508 = 1_n4398 & 1_n8997;
assign 1_n8894 = ~(1_n6273 ^ 1_n12144);
assign 1_n1576 = ~(1_n10620 ^ 1_n1569);
assign 1_n4144 = ~1_n4470;
assign 1_n3775 = 1_n9888 & 1_n6394;
assign 1_n9103 = ~(1_n7012 ^ 1_n1160);
assign 1_n12059 = ~(1_n7324 ^ 1_n7996);
assign 1_n10755 = ~1_n6196;
assign 1_n12701 = 1_n2268 & 1_n3245;
assign 1_n8992 = 1_n1871 & 1_n2710;
assign 1_n10729 = ~(1_n8922 ^ 1_n11759);
assign 1_n6919 = 1_n5212 & 1_n6802;
assign 1_n4991 = ~(1_n10766 ^ 1_n2078);
assign 1_n13025 = ~1_n443;
assign 1_n227 = ~1_n8290;
assign 1_n9330 = 1_n1340 | 1_n8435;
assign 1_n3220 = ~(1_n10344 | 1_n266);
assign 1_n10433 = ~1_n9620;
assign 1_n2208 = ~(1_n3218 | 1_n6437);
assign 1_n6394 = 1_n8940 & 1_n6392;
assign 1_n9358 = ~(1_n5479 ^ 1_n2951);
assign 1_n5094 = 1_n6680 | 1_n7306;
assign 1_n10335 = 1_n7184 | 1_n8268;
assign 1_n8191 = ~(1_n6499 ^ 1_n7343);
assign 1_n4299 = ~(1_n5941 ^ 1_n4972);
assign 1_n2143 = ~(1_n5585 ^ 1_n8092);
assign 1_n4902 = ~(1_n1454 ^ 1_n9185);
assign 1_n3636 = 1_n569 | 1_n9195;
assign 1_n12699 = 1_n10830 | 1_n6732;
assign 1_n10764 = ~1_n10408;
assign 1_n10644 = ~1_n12550;
assign 1_n4214 = ~(1_n6898 ^ 1_n10146);
assign 1_n5149 = 1_n9980 & 1_n11424;
assign 1_n8319 = 1_n9217 & 1_n3688;
assign 1_n2621 = 1_n7240 & 1_n1528;
assign 1_n2112 = 1_n190 & 1_n12063;
assign 1_n9297 = 1_n10781 | 1_n8268;
assign 1_n5573 = ~(1_n4550 | 1_n3968);
assign 1_n13127 = 1_n9476 | 1_n3772;
assign 1_n5608 = 1_n2802 | 1_n12410;
assign 1_n558 = ~1_n212;
assign 1_n11654 = 1_n584 | 1_n10029;
assign 1_n9947 = ~(1_n1393 ^ 1_n5442);
assign 1_n3230 = 1_n12976 & 1_n4533;
assign 1_n1586 = 1_n8480 | 1_n10012;
assign 1_n4803 = ~(1_n5358 ^ 1_n7027);
assign 1_n10377 = ~(1_n10115 | 1_n9799);
assign 1_n12248 = ~(1_n8842 ^ 1_n5984);
assign 1_n7571 = 1_n4657 | 1_n10179;
assign 1_n760 = 1_n9878 & 1_n3030;
assign 1_n5443 = ~(1_n7454 | 1_n7099);
assign 1_n2261 = 1_n13012 | 1_n11107;
assign 1_n5507 = ~(1_n12593 | 1_n350);
assign 1_n10211 = ~1_n12356;
assign 1_n911 = ~(1_n8135 | 1_n6822);
assign 1_n6258 = ~(1_n7460 | 1_n4450);
assign 1_n2060 = ~(1_n1864 ^ 1_n10712);
assign 1_n4840 = 1_n12378 & 1_n11059;
assign 1_n12125 = ~(1_n8284 ^ 1_n4543);
assign 1_n11932 = ~(1_n9206 ^ 1_n2645);
assign 1_n8379 = ~(1_n9948 ^ 1_n6288);
assign 1_n816 = ~1_n8071;
assign 1_n3939 = 1_n9710 & 1_n11846;
assign 1_n2326 = 1_n11492 | 1_n8711;
assign 1_n8413 = ~1_n7376;
assign 1_n8674 = ~(1_n2442 ^ 1_n8634);
assign 1_n12799 = 1_n3003 | 1_n4662;
assign 1_n4352 = ~1_n6085;
assign 1_n5574 = ~(1_n2786 ^ 1_n669);
assign 1_n1490 = 1_n2556 | 1_n4230;
assign 1_n10592 = ~(1_n1131 ^ 1_n8192);
assign 1_n324 = ~(1_n6396 | 1_n11425);
assign 1_n13044 = 1_n9966 & 1_n4720;
assign 1_n10503 = 1_n5847 | 1_n7515;
assign 1_n9568 = 1_n5921 & 1_n8571;
assign 1_n8655 = ~1_n1626;
assign 1_n5973 = ~1_n12284;
assign 1_n5708 = 1_n6580 & 1_n8942;
assign 1_n6519 = ~1_n2339;
assign 1_n7592 = ~(1_n1763 ^ 1_n5132);
assign 1_n9516 = ~(1_n8979 ^ 1_n10320);
assign 1_n9757 = 1_n2427 & 1_n2178;
assign 1_n4530 = ~1_n832;
assign 1_n11311 = 1_n2736 & 1_n2659;
assign 1_n2346 = ~1_n12579;
assign 1_n10756 = ~1_n3409;
assign 1_n614 = 1_n1553 | 1_n7964;
assign 1_n9381 = 1_n9468 & 1_n11919;
assign 1_n11929 = ~1_n9906;
assign 1_n12122 = 1_n7805 | 1_n2059;
assign 1_n11496 = ~(1_n7114 | 1_n4192);
assign 1_n8209 = 1_n5275 & 1_n3109;
assign 1_n4702 = ~(1_n7693 | 1_n5977);
assign 1_n4851 = 1_n11587 & 1_n12974;
assign 1_n199 = 1_n7026 & 1_n10964;
assign 1_n943 = 1_n3109 | 1_n5275;
assign 1_n1719 = 1_n11498 & 1_n458;
assign 1_n3798 = 1_n12788 & 1_n6900;
assign 1_n3603 = ~(1_n7958 ^ 1_n2682);
assign 1_n5308 = ~(1_n10538 | 1_n5650);
assign 1_n2210 = ~(1_n7345 | 1_n11613);
assign 1_n4918 = ~(1_n5110 ^ 1_n1217);
assign 1_n8730 = 1_n794 & 1_n2980;
assign 1_n7647 = ~(1_n10666 | 1_n10752);
assign 1_n7408 = ~(1_n12728 ^ 1_n9139);
assign 1_n1130 = 1_n2104 & 1_n10808;
assign 1_n1966 = ~(1_n6545 ^ 1_n4131);
assign 1_n4483 = ~(1_n3007 ^ 1_n8847);
assign 1_n12691 = ~(1_n998 ^ 1_n1399);
assign 1_n8288 = ~(1_n7938 ^ 1_n12966);
assign 1_n2924 = 1_n7152 | 1_n1570;
assign 1_n9834 = 1_n2204 | 1_n1546;
assign 1_n11477 = ~(1_n4181 ^ 1_n11013);
assign 1_n867 = 1_n8850 | 1_n9907;
assign 1_n1401 = 1_n66 ^ 1_n4111;
assign 1_n818 = 1_n13173 & 1_n1388;
assign 1_n2018 = ~1_n10866;
assign 1_n2759 = 1_n10662 & 1_n13027;
assign 1_n9256 = 1_n1474 | 1_n5450;
assign 1_n8038 = ~1_n2771;
assign 1_n11816 = ~(1_n10961 ^ 1_n6552);
assign 1_n1527 = 1_n6063 | 1_n2544;
assign 1_n2652 = 1_n5586 & 1_n12263;
assign 1_n2219 = ~(1_n4574 ^ 1_n12340);
assign 1_n12752 = ~1_n6032;
assign 1_n8300 = ~(1_n4648 ^ 1_n11155);
assign 1_n8862 = 1_n321 | 1_n3981;
assign 1_n7871 = 1_n11827 & 1_n9395;
assign 1_n7929 = 1_n11231 & 1_n9202;
assign 1_n6125 = 1_n2641 | 1_n6404;
assign 1_n2539 = 1_n10099 & 1_n10275;
assign 1_n12402 = 1_n9910 | 1_n9741;
assign 1_n10545 = 1_n7915 & 1_n5395;
assign 1_n10046 = ~(1_n3238 | 1_n9242);
assign 1_n7602 = ~1_n8822;
assign 1_n9253 = 1_n4876 | 1_n769;
assign 1_n10135 = ~1_n2758;
assign 1_n4541 = ~(1_n1928 ^ 1_n8089);
assign 1_n4344 = ~(1_n3585 | 1_n5779);
assign 1_n7196 = 1_n5477 | 1_n5174;
assign 1_n6621 = ~(1_n8976 ^ 1_n13179);
assign 1_n11901 = 1_n3892 | 1_n7935;
assign 1_n8857 = ~1_n7116;
assign 1_n9447 = ~(1_n791 ^ 1_n2376);
assign 1_n3556 = 1_n2848 | 1_n479;
assign 1_n5076 = 1_n218;
assign 1_n2554 = ~(1_n8272 | 1_n3337);
assign 1_n8197 = ~(1_n364 ^ 1_n5178);
assign 1_n8496 = 1_n9519 | 1_n6541;
assign 1_n1199 = ~1_n12289;
assign 1_n12487 = ~(1_n4797 | 1_n1405);
assign 1_n6563 = ~1_n5284;
assign 1_n10676 = 1_n11562 | 1_n7335;
assign 1_n9778 = 1_n12220 & 1_n2100;
assign 1_n11285 = ~(1_n5945 ^ 1_n13199);
assign 1_n111 = ~1_n11433;
assign 1_n3584 = ~1_n4630;
assign 1_n11114 = ~1_n10594;
assign 1_n8117 = ~(1_n7680 ^ 1_n12818);
assign 1_n9408 = 1_n10427 & 1_n3424;
assign 1_n5931 = ~(1_n8631 | 1_n9752);
assign 1_n12894 = ~(1_n3819 ^ 1_n10295);
assign 1_n7262 = ~1_n4682;
assign 1_n6975 = 1_n7216 | 1_n8563;
assign 1_n4639 = 1_n334 | 1_n3225;
assign 1_n2964 = ~(1_n4475 ^ 1_n6999);
assign 1_n166 = ~(1_n7639 ^ 1_n4327);
assign 1_n9229 = 1_n5227 & 1_n6391;
assign 1_n10578 = 1_n9701 & 1_n10457;
assign 1_n12925 = ~(1_n12777 ^ 1_n13210);
assign 1_n5270 = 1_n1757 & 1_n9669;
assign 1_n94 = ~(1_n6549 ^ 1_n9167);
assign 1_n6321 = 1_n7595 & 1_n12133;
assign 1_n11465 = 1_n5308 | 1_n9379;
assign 1_n6521 = ~(1_n3322 | 1_n4913);
assign 1_n83 = ~(1_n7376 ^ 1_n1567);
assign 1_n589 = 1_n11635 & 1_n3006;
assign 1_n6910 = ~(1_n6471 | 1_n4955);
assign 1_n9602 = ~(1_n5345 | 1_n11727);
assign 1_n2271 = ~1_n1646;
assign 1_n10401 = ~(1_n5380 ^ 1_n7417);
assign 1_n7920 = ~(1_n197 | 1_n8785);
assign 1_n12560 = 1_n4366 | 1_n6635;
assign 1_n6848 = ~(1_n9700 ^ 1_n4652);
assign 1_n6764 = ~1_n564;
assign 1_n3497 = 1_n1739 & 1_n11462;
assign 1_n3472 = ~(1_n11280 ^ 1_n8000);
assign 1_n1012 = ~1_n11488;
assign 1_n4973 = ~(1_n2258 ^ 1_n4017);
assign 1_n1153 = 1_n6970 & 1_n4445;
assign 1_n1973 = ~1_n9032;
assign 1_n5737 = 1_n9310 | 1_n6040;
assign 1_n8753 = 1_n6004 | 1_n12443;
assign 1_n462 = 1_n5261 | 1_n5242;
assign 1_n8545 = 1_n9809 | 1_n1094;
assign 1_n1161 = 1_n8305 & 1_n9695;
assign 1_n4137 = 1_n2027 | 1_n6728;
assign 1_n7307 = 1_n685 & 1_n8068;
assign 1_n144 = 1_n2381 | 1_n5778;
assign 1_n12593 = ~(1_n3526 | 1_n12933);
assign 1_n5987 = ~(1_n6531 ^ 1_n1717);
assign 1_n3945 = 1_n12376 | 1_n6081;
assign 1_n694 = ~1_n772;
assign 1_n2681 = ~1_n5735;
assign 1_n3513 = 1_n11419 & 1_n943;
assign 1_n5332 = ~(1_n3209 ^ 1_n8721);
assign 1_n6608 = ~1_n1972;
assign 1_n3406 = ~(1_n12431 ^ 1_n3782);
assign 1_n12584 = 1_n8463 | 1_n7306;
assign 1_n11136 = ~(1_n11935 ^ 1_n3811);
assign 1_n8141 = 1_n13159 | 1_n3981;
assign 1_n7331 = 1_n1398 | 1_n11616;
assign 1_n12641 = 1_n162 & 1_n8051;
assign 1_n1157 = 1_n5459 & 1_n5474;
assign 1_n5952 = ~(1_n8521 ^ 1_n2577);
assign 1_n3676 = ~1_n937;
assign 1_n8893 = ~(1_n11379 ^ 1_n11995);
assign 1_n5162 = 1_n484 & 1_n7618;
assign 1_n13156 = ~(1_n10583 | 1_n5241);
assign 1_n6246 = ~(1_n1225 ^ 1_n8583);
assign 1_n11262 = 1_n160 ^ 1_n6585;
assign 1_n5988 = 1_n12776 | 1_n11603;
assign 1_n5264 = ~1_n411;
assign 1_n11576 = 1_n2624 & 1_n5135;
assign 1_n1283 = ~(1_n10658 ^ 1_n11579);
assign 1_n721 = 1_n667 & 1_n5693;
assign 1_n4017 = 1_n8239 & 1_n12500;
assign 1_n6552 = ~(1_n8394 ^ 1_n5310);
assign 1_n9785 = ~(1_n4717 ^ 1_n5115);
assign 1_n11409 = ~(1_n6189 ^ 1_n5685);
assign 1_n6113 = 1_n10772 | 1_n4947;
assign 1_n12219 = 1_n10044 & 1_n1376;
assign 1_n5476 = ~(1_n12885 | 1_n2629);
assign 1_n10943 = 1_n10761 | 1_n12328;
assign 1_n8477 = ~(1_n5795 ^ 1_n5510);
assign 1_n12001 = 1_n6359 | 1_n6014;
assign 1_n7306 = ~1_n5920;
assign 1_n7483 = 1_n8609 | 1_n12174;
assign 1_n6838 = 1_n4186 & 1_n1269;
assign 1_n2221 = ~1_n6392;
assign 1_n3613 = 1_n1002 & 1_n5390;
assign 1_n11388 = ~(1_n6811 ^ 1_n11364);
assign 1_n12904 = 1_n10279 | 1_n9754;
assign 1_n4292 = ~(1_n9584 ^ 1_n7948);
assign 1_n11485 = ~1_n5784;
assign 1_n6420 = ~1_n959;
assign 1_n12261 = ~(1_n10313 ^ 1_n1782);
assign 1_n5584 = 1_n4269 & 1_n8293;
assign 1_n9397 = 1_n995 & 1_n12970;
assign 1_n12730 = ~(1_n11669 ^ 1_n7936);
assign 1_n3805 = ~1_n9915;
assign 1_n1896 = 1_n12955 | 1_n488;
assign 1_n4184 = 1_n3963 | 1_n9492;
assign 1_n1041 = ~1_n9508;
assign 1_n10973 = 1_n9277 ^ 1_n6269;
assign 1_n5809 = 1_n3575 & 1_n2700;
assign 1_n9386 = ~(1_n7426 | 1_n5080);
assign 1_n6022 = ~(1_n3530 ^ 1_n5676);
assign 1_n4442 = ~1_n6668;
assign 1_n9363 = ~(1_n10703 | 1_n4905);
assign 1_n6189 = 1_n1971 & 1_n939;
assign 1_n7557 = 1_n10426 & 1_n2098;
assign 1_n11727 = ~(1_n1294 | 1_n12975);
assign 1_n942 = ~(1_n3721 ^ 1_n4053);
assign 1_n12430 = 1_n12535 & 1_n2271;
assign 1_n5726 = 1_n8592 & 1_n8579;
assign 1_n8789 = 1_n2744 & 1_n12424;
assign 1_n12885 = ~1_n8758;
assign 1_n5322 = ~(1_n5603 ^ 1_n1176);
assign 1_n12787 = 1_n5054 & 1_n1574;
assign 1_n1696 = ~1_n761;
assign 1_n12009 = ~1_n7729;
assign 1_n11053 = 1_n6451 | 1_n8032;
assign 1_n7591 = 1_n12767 | 1_n10445;
assign 1_n2814 = ~(1_n12286 ^ 1_n113);
assign 1_n11818 = 1_n7317 | 1_n3261;
assign 1_n7358 = ~1_n3669;
assign 1_n5488 = ~(1_n6156 ^ 1_n12403);
assign 1_n7132 = ~(1_n8822 ^ 1_n1162);
assign 1_n1755 = ~(1_n2928 ^ 1_n3228);
assign 1_n2108 = ~(1_n11228 ^ 1_n7529);
assign 1_n9698 = ~1_n11930;
assign 1_n13208 = ~(1_n9164 ^ 1_n3256);
assign 1_n1545 = 1_n10437 | 1_n2544;
assign 1_n7454 = ~(1_n108 | 1_n2892);
assign 1_n306 = 1_n3070 & 1_n4930;
assign 1_n3510 = ~1_n3974;
assign 1_n3005 = ~(1_n11718 ^ 1_n5081);
assign 1_n1211 = ~1_n10186;
assign 1_n3098 = ~(1_n6813 ^ 1_n3284);
assign 1_n1676 = 1_n377 & 1_n6930;
assign 1_n6863 = 1_n4433 & 1_n9964;
assign 1_n6247 = 1_n3512 & 1_n5794;
assign 1_n10244 = ~1_n1974;
assign 1_n11504 = 1_n7033 | 1_n10213;
assign 1_n11564 = 1_n11192 | 1_n9199;
assign 1_n12245 = ~(1_n11657 ^ 1_n10176);
assign 1_n5821 = 1_n5455 | 1_n4373;
assign 1_n10148 = ~(1_n6525 | 1_n12730);
assign 1_n7091 = ~1_n6763;
assign 1_n4905 = ~(1_n8442 ^ 1_n221);
assign 1_n6360 = ~1_n11584;
assign 1_n12109 = ~1_n1165;
assign 1_n11682 = ~(1_n1090 ^ 1_n7835);
assign 1_n7877 = ~1_n7281;
assign 1_n8494 = ~1_n7844;
assign 1_n9050 = ~(1_n4898 ^ 1_n3028);
assign 1_n4008 = ~(1_n4496 ^ 1_n3370);
assign 1_n3329 = 1_n7156 & 1_n1932;
assign 1_n3834 = 1_n10883 | 1_n10319;
assign 1_n1390 = ~1_n4135;
assign 1_n5644 = 1_n1139 | 1_n6216;
assign 1_n3321 = 1_n6295 | 1_n2637;
assign 1_n8533 = ~1_n3439;
assign 1_n354 = 1_n9579 & 1_n5233;
assign 1_n5119 = ~1_n7734;
assign 1_n6444 = 1_n3958 | 1_n2846;
assign 1_n1737 = ~1_n8290;
assign 1_n1014 = ~(1_n3893 ^ 1_n1993);
assign 1_n6385 = 1_n2673 & 1_n5726;
assign 1_n2298 = 1_n3928 | 1_n10871;
assign 1_n12466 = ~(1_n12864 | 1_n2110);
assign 1_n1248 = ~(1_n8308 | 1_n5214);
assign 1_n13101 = 1_n1941 | 1_n4640;
assign 1_n12578 = 1_n8308 & 1_n9669;
assign 1_n1293 = ~(1_n6738 ^ 1_n9486);
assign 1_n2276 = ~1_n8183;
assign 1_n2470 = ~(1_n3654 ^ 1_n12070);
assign 1_n7038 = ~(1_n2764 ^ 1_n4123);
assign 1_n1508 = ~1_n6471;
assign 1_n2176 = ~(1_n8659 ^ 1_n9755);
assign 1_n6419 = ~1_n7113;
assign 1_n682 = ~(1_n3695 | 1_n5723);
assign 1_n830 = 1_n4153 | 1_n10973;
assign 1_n3240 = 1_n12851 | 1_n13112;
assign 1_n5539 = ~(1_n114 | 1_n10866);
assign 1_n7259 = ~(1_n13000 ^ 1_n9753);
assign 1_n8059 = ~(1_n10326 ^ 1_n7793);
assign 1_n4082 = ~(1_n540 ^ 1_n8760);
assign 1_n2212 = 1_n7662 & 1_n1006;
assign 1_n1981 = ~(1_n10564 | 1_n7521);
assign 1_n2151 = 1_n11840 & 1_n12036;
assign 1_n2007 = ~(1_n12716 | 1_n7785);
assign 1_n12585 = 1_n6801 | 1_n4062;
assign 1_n192 = ~1_n4821;
assign 1_n5877 = 1_n9159 | 1_n5076;
assign 1_n2398 = 1_n4456 & 1_n5353;
assign 1_n6740 = ~(1_n2310 ^ 1_n7605);
assign 1_n6389 = 1_n7154 & 1_n8898;
assign 1_n416 = ~(1_n6104 ^ 1_n9053);
assign 1_n846 = ~(1_n7779 ^ 1_n2482);
assign 1_n11591 = ~1_n854;
assign 1_n6042 = ~(1_n3061 | 1_n13192);
assign 1_n1212 = 1_n5168 | 1_n10029;
assign 1_n10780 = ~1_n3112;
assign 1_n10947 = 1_n6303 | 1_n10601;
assign 1_n11577 = ~(1_n12756 | 1_n8557);
assign 1_n5804 = ~(1_n8919 ^ 1_n167);
assign 1_n4741 = ~1_n11634;
assign 1_n3413 = ~1_n684;
assign 1_n2427 = 1_n2357 | 1_n11857;
assign 1_n7919 = ~(1_n7467 ^ 1_n1476);
assign 1_n2731 = 1_n9721 & 1_n7606;
assign 1_n1148 = 1_n11225 | 1_n4373;
assign 1_n12412 = 1_n7172 | 1_n11978;
assign 1_n5074 = 1_n12256 & 1_n10353;
assign 1_n7065 = ~(1_n4458 ^ 1_n11083);
assign 1_n5406 = 1_n11195 & 1_n10110;
assign 1_n6381 = ~1_n9906;
assign 1_n4920 = 1_n5279 & 1_n10305;
assign 1_n9373 = ~(1_n4507 ^ 1_n1342);
assign 1_n2075 = ~(1_n8420 ^ 1_n12064);
assign 1_n9688 = ~(1_n656 ^ 1_n3685);
assign 1_n1975 = 1_n7707 | 1_n121;
assign 1_n6185 = ~(1_n9728 ^ 1_n11555);
assign 1_n8532 = ~1_n4335;
assign 1_n11524 = ~(1_n1225 | 1_n6716);
assign 1_n2428 = 1_n7889 | 1_n2685;
assign 1_n3547 = 1_n3520 | 1_n6377;
assign 1_n424 = 1_n10256 | 1_n10871;
assign 1_n11423 = 1_n1571 | 1_n6404;
assign 1_n218 = ~1_n7715;
assign 1_n4656 = ~(1_n4491 ^ 1_n7733);
assign 1_n5201 = ~(1_n9462 ^ 1_n11795);
assign 1_n11209 = 1_n2236 & 1_n5774;
assign 1_n6108 = 1_n4310 & 1_n13205;
assign 1_n5807 = 1_n9479 | 1_n8883;
assign 1_n8792 = 1_n10712 | 1_n1864;
assign 1_n10298 = ~(1_n8288 ^ 1_n10442);
assign 1_n9338 = ~(1_n8497 | 1_n7400);
assign 1_n1861 = ~(1_n9227 | 1_n9207);
assign 1_n3196 = ~(1_n790 ^ 1_n7528);
assign 1_n10365 = ~(1_n12157 ^ 1_n6070);
assign 1_n1732 = ~1_n7617;
assign 1_n5731 = ~(1_n11681 ^ 1_n13065);
assign 1_n4061 = 1_n3132 | 1_n5286;
assign 1_n4165 = 1_n2589 & 1_n12806;
assign 1_n7413 = 1_n3898 | 1_n3981;
assign 1_n4735 = ~(1_n749 | 1_n7756);
assign 1_n9291 = ~(1_n4685 ^ 1_n12443);
assign 1_n11201 = ~(1_n10070 ^ 1_n10663);
assign 1_n6703 = ~(1_n13220 | 1_n3232);
assign 1_n8736 = 1_n13149 | 1_n13113;
assign 1_n12287 = 1_n2281 & 1_n973;
assign 1_n6097 = ~1_n1718;
assign 1_n988 = ~(1_n2169 ^ 1_n8624);
assign 1_n4781 = ~(1_n3153 ^ 1_n3806);
assign 1_n7256 = ~(1_n6523 ^ 1_n9241);
assign 1_n641 = 1_n6939 | 1_n9195;
assign 1_n1163 = ~(1_n2090 ^ 1_n11305);
assign 1_n9212 = 1_n677 & 1_n5703;
assign 1_n2094 = ~(1_n11655 | 1_n870);
assign 1_n6021 = ~(1_n8908 ^ 1_n8376);
assign 1_n1074 = ~(1_n1746 | 1_n262);
assign 1_n3466 = 1_n4857 | 1_n3747;
assign 1_n6749 = ~1_n103;
assign 1_n737 = ~1_n8163;
assign 1_n9968 = 1_n3746 & 1_n10913;
assign 1_n5401 = ~1_n4998;
assign 1_n6464 = ~1_n9705;
assign 1_n7564 = 1_n2861 | 1_n206;
assign 1_n5146 = ~1_n603;
assign 1_n3931 = ~1_n7455;
assign 1_n217 = ~(1_n2476 ^ 1_n10707);
assign 1_n10710 = 1_n5035 | 1_n859;
assign 1_n11446 = ~1_n411;
assign 1_n6485 = ~(1_n3888 ^ 1_n7828);
assign 1_n12031 = ~1_n344;
assign 1_n6380 = ~1_n4773;
assign 1_n11782 = ~(1_n9640 ^ 1_n12158);
assign 1_n2456 = ~(1_n6366 | 1_n6871);
assign 1_n12529 = 1_n1941 | 1_n10106;
assign 1_n7351 = 1_n8329 | 1_n4724;
assign 1_n7895 = 1_n5772 & 1_n7899;
assign 1_n5551 = ~(1_n7426 ^ 1_n635);
assign 1_n1902 = ~(1_n7401 ^ 1_n5852);
assign 1_n12323 = 1_n6259 | 1_n3461;
assign 1_n9860 = 1_n3630 | 1_n2675;
assign 1_n4227 = ~1_n502;
assign 1_n12389 = ~(1_n10608 ^ 1_n12898);
assign 1_n2248 = 1_n9679 | 1_n11137;
assign 1_n3378 = ~(1_n7354 ^ 1_n501);
assign 1_n861 = 1_n6388 | 1_n8461;
assign 1_n2961 = 1_n6568 | 1_n6290;
assign 1_n2680 = 1_n4128 | 1_n9982;
assign 1_n12260 = ~(1_n11685 ^ 1_n6124);
assign 1_n222 = 1_n3816 | 1_n4682;
assign 1_n1706 = ~1_n10167;
assign 1_n3012 = 1_n3901 & 1_n12326;
assign 1_n4543 = 1_n2318 & 1_n12046;
assign 1_n104 = 1_n9769 | 1_n6044;
assign 1_n12194 = ~(1_n11918 | 1_n6962);
assign 1_n10842 = 1_n4105 & 1_n9354;
assign 1_n12407 = ~(1_n10513 ^ 1_n1550);
assign 1_n5946 = 1_n4988 | 1_n2496;
assign 1_n9963 = ~(1_n7811 ^ 1_n6179);
assign 1_n1441 = 1_n9040 & 1_n4381;
assign 1_n3197 = 1_n5018 | 1_n4477;
assign 1_n11946 = 1_n12394 | 1_n8367;
assign 1_n9145 = ~1_n1641;
assign 1_n3888 = 1_n7780 | 1_n10871;
assign 1_n9484 = 1_n628 | 1_n9195;
assign 1_n461 = ~(1_n10132 ^ 1_n1779);
assign 1_n1813 = ~1_n6661;
assign 1_n5723 = 1_n12812 & 1_n602;
assign 1_n213 = ~(1_n6043 ^ 1_n12423);
assign 1_n2077 = ~(1_n11261 | 1_n4216);
assign 1_n11844 = ~(1_n7882 | 1_n1923);
assign 1_n10521 = 1_n6591 & 1_n11385;
assign 1_n6304 = ~(1_n11937 | 1_n2920);
assign 1_n1118 = ~(1_n7933 ^ 1_n7244);
assign 1_n10161 = ~1_n2164;
assign 1_n4274 = 1_n7414 | 1_n8845;
assign 1_n8138 = 1_n4201 | 1_n2059;
assign 1_n6064 = 1_n2482 & 1_n6149;
assign 1_n9138 = ~(1_n2024 ^ 1_n12006);
assign 1_n13016 = 1_n3783 | 1_n10818;
assign 1_n692 = 1_n8062 | 1_n99;
assign 1_n4410 = ~(1_n10476 ^ 1_n8809);
assign 1_n8647 = 1_n3282 & 1_n7196;
assign 1_n3601 = ~(1_n1766 ^ 1_n976);
assign 1_n4002 = 1_n4506 & 1_n3617;
assign 1_n10476 = ~1_n10356;
assign 1_n9380 = ~1_n12820;
assign 1_n3069 = 1_n1733 | 1_n7079;
assign 1_n8079 = ~1_n9620;
assign 1_n168 = ~1_n6386;
assign 1_n4089 = 1_n11661 & 1_n9525;
assign 1_n6693 = ~(1_n8048 ^ 1_n11210);
assign 1_n3038 = ~1_n5572;
assign 1_n5925 = ~(1_n2434 ^ 1_n12854);
assign 1_n8312 = ~(1_n9347 ^ 1_n10933);
assign 1_n2199 = ~1_n5336;
assign 1_n3465 = ~(1_n492 ^ 1_n5894);
assign 1_n3778 = 1_n4432 | 1_n6119;
assign 1_n6037 = ~(1_n13226 | 1_n13064);
assign 1_n8772 = ~(1_n9877 ^ 1_n7777);
assign 1_n191 = 1_n8065 & 1_n2157;
assign 1_n1469 = 1_n4982 & 1_n3652;
assign 1_n8855 = ~1_n1192;
assign 1_n1348 = ~(1_n3771 ^ 1_n158);
assign 1_n7020 = 1_n1504 & 1_n11669;
assign 1_n12141 = 1_n7291 | 1_n2287;
assign 1_n3985 = 1_n12620 & 1_n6170;
assign 1_n9996 = 1_n8486 & 1_n3141;
assign 1_n9165 = ~(1_n10941 ^ 1_n7407);
assign 1_n11588 = ~(1_n7307 ^ 1_n1818);
assign 1_n852 = 1_n11869 & 1_n8755;
assign 1_n11876 = 1_n1377 | 1_n6760;
assign 1_n5050 = 1_n10923 | 1_n804;
assign 1_n2281 = 1_n6625 & 1_n9346;
assign 1_n9630 = ~(1_n7225 | 1_n5126);
assign 1_n559 = ~1_n5920;
assign 1_n1294 = 1_n1051 | 1_n1144;
assign 1_n2435 = ~(1_n942 ^ 1_n2084);
assign 1_n6762 = ~(1_n12124 ^ 1_n12205);
assign 1_n9842 = ~(1_n7177 ^ 1_n12265);
assign 1_n5672 = 1_n6365 ^ 1_n872;
assign 1_n2542 = ~1_n6668;
assign 1_n4443 = 1_n11427 & 1_n2021;
assign 1_n4170 = ~(1_n7714 | 1_n7338);
assign 1_n12304 = ~1_n5951;
assign 1_n525 = 1_n8637 | 1_n3686;
assign 1_n11880 = 1_n5694 | 1_n10319;
assign 1_n2791 = ~1_n9358;
assign 1_n7382 = ~(1_n3033 ^ 1_n11207);
assign 1_n9364 = ~(1_n6202 ^ 1_n8897);
assign 1_n10653 = ~(1_n11248 ^ 1_n5179);
assign 1_n5063 = ~(1_n4242 | 1_n598);
assign 1_n6035 = 1_n2338 | 1_n10319;
assign 1_n1476 = ~(1_n3780 ^ 1_n8685);
assign 1_n9692 = ~(1_n7051 ^ 1_n9380);
assign 1_n8546 = 1_n13159 | 1_n10319;
assign 1_n1557 = 1_n3791 | 1_n10008;
assign 1_n6398 = ~(1_n226 | 1_n12075);
assign 1_n9095 = ~1_n8330;
assign 1_n3320 = 1_n1959 & 1_n11139;
assign 1_n9861 = 1_n8585 | 1_n5076;
assign 1_n5169 = ~1_n2771;
assign 1_n5606 = ~(1_n419 | 1_n6577);
assign 1_n7711 = ~(1_n50 ^ 1_n11782);
assign 1_n9075 = 1_n16;
assign 1_n8920 = ~(1_n6804 ^ 1_n8372);
assign 1_n6460 = ~(1_n699 ^ 1_n6798);
assign 1_n7021 = ~(1_n1123 ^ 1_n7967);
assign 1_n5152 = ~1_n9093;
assign 1_n13008 = ~(1_n7797 | 1_n5996);
assign 1_n12882 = ~1_n1307;
assign 1_n6633 = 1_n5017 & 1_n1019;
assign 1_n8425 = 1_n434 | 1_n3787;
assign 1_n10449 = ~(1_n1840 ^ 1_n8844);
assign 1_n9525 = 1_n10566 | 1_n11877;
assign 1_n6573 = ~(1_n12041 | 1_n2635);
assign 1_n3290 = ~(1_n4749 ^ 1_n9044);
assign 1_n6631 = ~(1_n3288 ^ 1_n5291);
assign 1_n11516 = ~(1_n1568 ^ 1_n11043);
assign 1_n2103 = ~(1_n5799 | 1_n9645);
assign 1_n2866 = ~(1_n299 ^ 1_n10773);
assign 1_n3830 = 1_n5031 & 1_n8233;
assign 1_n6179 = 1_n5634 | 1_n3981;
assign 1_n4598 = 1_n8976 | 1_n13179;
assign 1_n13185 = 1_n1728 & 1_n5551;
assign 1_n6586 = ~(1_n9381 ^ 1_n10192);
assign 1_n3325 = 1_n7393 | 1_n6266;
assign 1_n4106 = ~(1_n5395 ^ 1_n11639);
assign 1_n5799 = 1_n6332 | 1_n6404;
assign 1_n2701 = ~1_n10451;
assign 1_n1915 = 1_n7149 & 1_n6098;
assign 1_n5278 = 1_n8095 | 1_n4932;
assign 1_n1488 = ~(1_n243 ^ 1_n4863);
assign 1_n12893 = ~(1_n4802 ^ 1_n1149);
assign 1_n7596 = ~(1_n931 ^ 1_n7543);
assign 1_n2537 = ~(1_n8357 ^ 1_n6865);
assign 1_n7041 = ~1_n2339;
assign 1_n2486 = 1_n1671 & 1_n11642;
assign 1_n10752 = ~(1_n10651 ^ 1_n6876);
assign 1_n2744 = ~1_n11096;
assign 1_n12027 = 1_n9048 | 1_n3635;
assign 1_n13223 = ~(1_n8407 ^ 1_n4247);
assign 1_n3333 = 1_n9962 | 1_n9195;
assign 1_n1668 = 1_n5799 & 1_n9645;
assign 1_n550 = 1_n4086 & 1_n6064;
assign 1_n4529 = ~(1_n2908 | 1_n6060);
assign 1_n1478 = ~(1_n4244 | 1_n5961);
assign 1_n10477 = ~(1_n1507 ^ 1_n7097);
assign 1_n11778 = ~(1_n8560 ^ 1_n5672);
assign 1_n7977 = ~1_n8970;
assign 1_n13042 = ~(1_n2164 ^ 1_n7090);
assign 1_n4441 = 1_n6056 | 1_n12164;
assign 1_n1150 = 1_n8556 | 1_n10871;
assign 1_n11435 = ~(1_n9559 ^ 1_n9704);
assign 1_n4436 = ~(1_n11526 ^ 1_n12347);
assign 1_n11721 = 1_n10603 | 1_n6540;
assign 1_n6680 = ~1_n9732;
assign 1_n4820 = ~(1_n1185 ^ 1_n5059);
assign 1_n8928 = 1_n11379 | 1_n8841;
assign 1_n11159 = ~(1_n294 ^ 1_n6648);
assign 1_n2538 = ~1_n10408;
assign 1_n4040 = 1_n1635 | 1_n1572;
assign 1_n2987 = 1_n6487 ^ 1_n826;
assign 1_n7371 = ~1_n11872;
assign 1_n11837 = ~(1_n6385 ^ 1_n2836);
assign 1_n10583 = ~(1_n12790 | 1_n9807);
assign 1_n12927 = ~(1_n6933 | 1_n7562);
assign 1_n11823 = ~1_n1176;
assign 1_n1486 = 1_n4822 & 1_n830;
assign 1_n5454 = 1_n2965 ^ 1_n6704;
assign 1_n3301 = ~1_n2962;
assign 1_n10203 = ~1_n11201;
assign 1_n9349 = 1_n2799 | 1_n2451;
assign 1_n4872 = ~(1_n1351 ^ 1_n4205);
assign 1_n9997 = 1_n8720 | 1_n3703;
assign 1_n1671 = ~1_n10547;
assign 1_n5600 = 1_n11729 | 1_n8348;
assign 1_n8116 = 1_n265 & 1_n6657;
assign 1_n438 = ~1_n1007;
assign 1_n5398 = ~(1_n9432 ^ 1_n9263);
assign 1_n13110 = 1_n333 | 1_n2222;
assign 1_n1516 = 1_n1962 & 1_n3685;
assign 1_n6876 = ~(1_n11070 ^ 1_n3503);
assign 1_n5582 = 1_n11094 | 1_n8490;
assign 1_n6948 = ~(1_n2418 ^ 1_n2139);
assign 1_n7794 = 1_n5923 | 1_n7935;
assign 1_n9302 = ~(1_n12719 | 1_n10778);
assign 1_n7110 = ~1_n6574;
assign 1_n6750 = ~1_n2734;
assign 1_n4971 = 1_n4257 & 1_n12988;
assign 1_n1566 = 1_n12510 & 1_n619;
assign 1_n10871 = 1_n4517;
assign 1_n5578 = ~(1_n10683 ^ 1_n12393);
assign 1_n9702 = ~1_n5758;
assign 1_n3476 = ~(1_n7549 ^ 1_n3380);
assign 1_n1313 = 1_n5303 | 1_n2032;
assign 1_n7032 = 1_n11797 & 1_n12311;
assign 1_n5370 = 1_n12052 | 1_n6635;
assign 1_n4020 = 1_n10716 & 1_n9813;
assign 1_n2246 = 1_n5010 & 1_n8943;
assign 1_n9494 = 1_n1353 | 1_n1144;
assign 1_n77 = ~(1_n4007 ^ 1_n6665);
assign 1_n10174 = 1_n39 | 1_n3103;
assign 1_n2028 = ~1_n7273;
assign 1_n11424 = 1_n4558 | 1_n1811;
assign 1_n8110 = ~(1_n10713 ^ 1_n1692);
assign 1_n1748 = ~(1_n12030 ^ 1_n6748);
assign 1_n7102 = ~1_n12683;
assign 1_n4497 = 1_n4157 | 1_n4326;
assign 1_n3031 = ~1_n12953;
assign 1_n240 = 1_n4496 | 1_n1247;
assign 1_n6195 = ~(1_n3037 ^ 1_n11390);
assign 1_n11377 = ~(1_n12633 ^ 1_n8309);
assign 1_n4677 = 1_n2598 | 1_n13151;
assign 1_n12902 = 1_n4372 | 1_n1678;
assign 1_n11170 = 1_n4719 & 1_n1096;
assign 1_n12432 = 1_n79 | 1_n4640;
assign 1_n4650 = ~(1_n4624 | 1_n11495);
assign 1_n9551 = ~(1_n7975 ^ 1_n7523);
assign 1_n4415 = 1_n12004 & 1_n7738;
assign 1_n3549 = 1_n12848 & 1_n9466;
assign 1_n1595 = 1_n8115 & 1_n11041;
assign 1_n1363 = ~(1_n7225 ^ 1_n12359);
assign 1_n6822 = 1_n367 | 1_n12566;
assign 1_n8960 = 1_n6402 & 1_n9918;
assign 1_n10164 = ~(1_n10674 ^ 1_n6837);
assign 1_n13216 = 1_n12054 | 1_n5392;
assign 1_n1494 = 1_n10383 | 1_n7723;
assign 1_n7792 = 1_n333 | 1_n10956;
assign 1_n8987 = ~1_n5989;
assign 1_n3267 = ~(1_n4444 ^ 1_n8589);
assign 1_n7273 = 1_n13174 & 1_n1596;
assign 1_n13165 = 1_n5568 & 1_n10451;
assign 1_n1207 = 1_n11466 | 1_n10106;
assign 1_n12308 = ~1_n7035;
assign 1_n3298 = 1_n8971 & 1_n8936;
assign 1_n7767 = ~(1_n11828 | 1_n3452);
assign 1_n2713 = 1_n4291 | 1_n2562;
assign 1_n12686 = ~1_n9124;
assign 1_n9029 = 1_n2250 | 1_n10701;
assign 1_n6127 = ~(1_n2829 ^ 1_n8128);
assign 1_n12586 = ~(1_n1098 | 1_n2311);
assign 1_n2323 = ~1_n10134;
assign 1_n8912 = ~1_n11061;
assign 1_n4313 = 1_n7419 ^ 1_n9619;
assign 1_n515 = ~(1_n4673 | 1_n292);
assign 1_n3048 = 1_n10026 & 1_n4542;
assign 1_n897 = 1_n5037 & 1_n9651;
assign 1_n6299 = ~(1_n8271 ^ 1_n10626);
assign 1_n12296 = 1_n9310 | 1_n1571;
assign 1_n4478 = 1_n13077 | 1_n4640;
assign 1_n5058 = ~1_n11850;
assign 1_n2930 = ~1_n4426;
assign 1_n8775 = ~1_n3365;
assign 1_n6318 = 1_n4693 | 1_n814;
assign 1_n5111 = 1_n9614 | 1_n1581;
assign 1_n8416 = 1_n10476 | 1_n10126;
assign 1_n10591 = ~1_n7720;
assign 1_n10355 = 1_n1887 | 1_n8348;
assign 1_n7827 = ~1_n3693;
assign 1_n10615 = 1_n4206 & 1_n9023;
assign 1_n7878 = ~1_n7659;
assign 1_n6320 = 1_n2377 | 1_n6860;
assign 1_n6350 = ~(1_n11705 ^ 1_n4662);
assign 1_n7576 = ~(1_n966 ^ 1_n7336);
assign 1_n4852 = 1_n1096 | 1_n4719;
assign 1_n8221 = 1_n8487 | 1_n11822;
assign 1_n159 = ~1_n8150;
assign 1_n2289 = 1_n8904 | 1_n8030;
assign 1_n5086 = ~1_n103;
assign 1_n12220 = 1_n10591 | 1_n8534;
assign 1_n115 = ~1_n499;
assign 1_n10567 = ~(1_n7147 ^ 1_n397);
assign 1_n11911 = ~(1_n5185 | 1_n1734);
assign 1_n11080 = 1_n2872 | 1_n10029;
assign 1_n6156 = ~1_n3042;
assign 1_n10303 = ~(1_n13081 ^ 1_n11263);
assign 1_n9063 = ~(1_n9188 ^ 1_n1815);
assign 1_n3715 = 1_n10783 & 1_n125;
assign 1_n4816 = ~1_n4285;
assign 1_n2720 = 1_n7493 & 1_n2553;
assign 1_n903 = ~(1_n8402 ^ 1_n2783);
assign 1_n7314 = ~(1_n11486 ^ 1_n9410);
assign 1_n11256 = 1_n8161 & 1_n6651;
assign 1_n3139 = 1_n3572 | 1_n10352;
assign 1_n2475 = ~(1_n1523 ^ 1_n6197);
assign 1_n11420 = 1_n3225 | 1_n6732;
assign 1_n8902 = ~(1_n1411 ^ 1_n476);
assign 1_n11294 = 1_n13201 & 1_n11058;
assign 1_n7595 = 1_n5031 & 1_n287;
assign 1_n7820 = 1_n6005 & 1_n1150;
assign 1_n8799 = 1_n7730 | 1_n650;
assign 1_n11145 = ~(1_n11423 ^ 1_n3408);
assign 1_n9483 = 1_n2321 | 1_n3999;
assign 1_n12753 = ~(1_n7958 | 1_n5864);
assign 1_n9701 = 1_n9510 & 1_n11525;
assign 1_n6917 = ~1_n745;
assign 1_n422 = 1_n3284 | 1_n6813;
assign 1_n10395 = ~(1_n10026 ^ 1_n9802);
assign 1_n8487 = 1_n8744 | 1_n4179;
assign 1_n6109 = ~(1_n2112 ^ 1_n8501);
assign 1_n5662 = 1_n10127 & 1_n6645;
assign 1_n13013 = ~1_n937;
assign 1_n8879 = 1_n11333 | 1_n2942;
assign 1_n9975 = ~(1_n7702 ^ 1_n5989);
assign 1_n13191 = ~1_n6948;
assign 1_n727 = 1_n8406 & 1_n6076;
assign 1_n11814 = 1_n10304 & 1_n9517;
assign 1_n6199 = ~(1_n3481 | 1_n9338);
assign 1_n10284 = 1_n2095 | 1_n11810;
assign 1_n11334 = ~(1_n12696 ^ 1_n648);
assign 1_n10979 = 1_n7119 | 1_n12328;
assign 1_n9328 = 1_n6125 | 1_n9608;
assign 1_n10845 = 1_n7550 | 1_n9518;
assign 1_n653 = 1_n2280 & 1_n11102;
assign 1_n172 = 1_n8843 | 1_n12501;
assign 1_n2750 = ~(1_n10889 ^ 1_n4425);
assign 1_n4921 = 1_n7011 | 1_n7117;
assign 1_n12262 = 1_n2296 | 1_n10029;
assign 1_n11593 = ~1_n6650;
assign 1_n71 = 1_n784 & 1_n2433;
assign 1_n12840 = 1_n6355 | 1_n1696;
assign 1_n7364 = ~(1_n10625 | 1_n10160);
assign 1_n6103 = ~(1_n4023 ^ 1_n474);
assign 1_n1380 = ~(1_n2016 | 1_n2050);
assign 1_n11148 = ~1_n4382;
assign 1_n1107 = ~(1_n1798 ^ 1_n420);
assign 1_n10786 = ~1_n8675;
assign 1_n5483 = 1_n3178 & 1_n5548;
assign 1_n7961 = ~1_n1364;
assign 1_n7403 = 1_n6245 | 1_n3698;
assign 1_n3562 = ~(1_n8156 ^ 1_n10170);
assign 1_n10060 = 1_n6309 | 1_n6037;
assign 1_n945 = ~(1_n5269 ^ 1_n4939);
assign 1_n563 = 1_n7102 & 1_n1054;
assign 1_n8556 = ~1_n12306;
assign 1_n8267 = ~(1_n5942 ^ 1_n7334);
assign 1_n24 = 1_n11536 | 1_n911;
assign 1_n11657 = ~(1_n11407 ^ 1_n9550);
assign 1_n6884 = ~(1_n1854 ^ 1_n1273);
assign 1_n9647 = 1_n9557 | 1_n4686;
assign 1_n2000 = ~(1_n7840 ^ 1_n9435);
assign 1_n9374 = ~(1_n5230 ^ 1_n9636);
assign 1_n12512 = 1_n998 & 1_n11125;
assign 1_n562 = ~(1_n3929 | 1_n1853);
assign 1_n11206 = ~(1_n3057 ^ 1_n10863);
assign 1_n10541 = 1_n6225 | 1_n5414;
assign 1_n2969 = 1_n7429 & 1_n9567;
assign 1_n11393 = ~(1_n12143 | 1_n3793);
assign 1_n8176 = ~1_n8768;
assign 1_n6050 = ~(1_n12451 ^ 1_n2402);
assign 1_n1701 = 1_n1278 | 1_n3712;
assign 1_n11029 = ~1_n1876;
assign 1_n8663 = ~1_n10697;
assign 1_n3789 = ~(1_n502 ^ 1_n11588);
assign 1_n9091 = 1_n1584 & 1_n11572;
assign 1_n11879 = ~(1_n9418 ^ 1_n1057);
assign 1_n12568 = ~1_n497;
assign 1_n9383 = ~1_n5356;
assign 1_n13202 = ~(1_n6021 | 1_n1186);
assign 1_n9576 = ~(1_n4239 ^ 1_n11570);
assign 1_n759 = ~1_n2939;
assign 1_n7892 = ~(1_n4731 ^ 1_n5790);
assign 1_n4606 = ~1_n12488;
assign 1_n10858 = ~1_n12609;
assign 1_n1841 = 1_n2148 | 1_n1043;
assign 1_n5700 = 1_n10017 | 1_n12388;
assign 1_n2239 = ~(1_n6799 ^ 1_n7826);
assign 1_n2913 = ~(1_n8356 ^ 1_n456);
assign 1_n10065 = 1_n2677 | 1_n10912;
assign 1_n604 = ~(1_n6015 | 1_n7602);
assign 1_n3352 = 1_n3225 | 1_n10900;
assign 1_n7639 = ~(1_n11791 ^ 1_n269);
assign 1_n1810 = ~(1_n9951 ^ 1_n3495);
assign 1_n4646 = ~(1_n10537 ^ 1_n5049);
assign 1_n549 = ~1_n1254;
assign 1_n4372 = 1_n7821 & 1_n5039;
assign 1_n6399 = 1_n13000 & 1_n8981;
assign 1_n5972 = ~(1_n3958 ^ 1_n2846);
assign 1_n11940 = ~1_n8466;
assign 1_n4062 = ~(1_n10004 | 1_n3358);
assign 1_n381 = ~(1_n6657 ^ 1_n265);
assign 1_n2168 = 1_n7467 | 1_n2249;
assign 1_n3538 = 1_n12432 & 1_n3417;
assign 1_n435 = 1_n5767 | 1_n6589;
assign 1_n1162 = ~(1_n6015 ^ 1_n1529);
assign 1_n1067 = ~1_n7613;
assign 1_n8732 = 1_n476 & 1_n1411;
assign 1_n3045 = 1_n2232 | 1_n6814;
assign 1_n11291 = ~1_n9300;
assign 1_n11831 = ~(1_n214 | 1_n4378);
assign 1_n2790 = 1_n1212 & 1_n13061;
assign 1_n10980 = 1_n11130 & 1_n5208;
assign 1_n6459 = ~(1_n9567 ^ 1_n7429);
assign 1_n7392 = ~(1_n2337 ^ 1_n8277);
assign 1_n5852 = ~(1_n11343 ^ 1_n4595);
assign 1_n3278 = 1_n10582 & 1_n11887;
assign 1_n2029 = ~(1_n1310 ^ 1_n5632);
assign 1_n3260 = 1_n12948 | 1_n6265;
assign 1_n8597 = 1_n11706 & 1_n1379;
assign 1_n5020 = 1_n10366 & 1_n10328;
assign 1_n2127 = 1_n10566 & 1_n11877;
assign 1_n4704 = 1_n8998 | 1_n12132;
assign 1_n12538 = ~(1_n13203 ^ 1_n5487);
assign 1_n10639 = ~(1_n12313 ^ 1_n522);
assign 1_n1247 = 1_n3079 & 1_n4251;
assign 1_n9119 = ~1_n11059;
assign 1_n7344 = 1_n4668 & 1_n12726;
assign 1_n12339 = 1_n10860 & 1_n1347;
assign 1_n12265 = ~(1_n147 ^ 1_n10094);
assign 1_n3654 = ~(1_n6082 | 1_n12542);
assign 1_n6802 = 1_n5164 | 1_n7412;
assign 1_n5185 = ~(1_n4971 ^ 1_n6597);
assign 1_n5800 = ~(1_n13184 ^ 1_n6891);
assign 1_n2970 = ~1_n10642;
assign 1_n2167 = 1_n11643 & 1_n7378;
assign 1_n345 = ~(1_n4157 ^ 1_n2317);
assign 1_n2551 = ~1_n9929;
assign 1_n12581 = 1_n10530 & 1_n12938;
assign 1_n2259 = 1_n3940 | 1_n2637;
assign 1_n2868 = 1_n941 & 1_n12599;
assign 1_n9552 = 1_n1241 | 1_n11817;
assign 1_n7424 = ~1_n4141;
assign 1_n935 = ~1_n287;
assign 1_n8677 = 1_n4478 & 1_n1599;
assign 1_n6756 = ~1_n4597;
assign 1_n4157 = 1_n4077 | 1_n9638;
assign 1_n7998 = ~1_n9475;
assign 1_n6959 = 1_n12790 & 1_n9807;
assign 1_n3309 = ~(1_n12567 ^ 1_n8465);
assign 1_n4134 = 1_n1125 | 1_n4606;
assign 1_n8637 = 1_n6739 & 1_n9279;
assign 1_n5668 = 1_n12592 & 1_n3076;
assign 1_n3389 = ~(1_n8031 ^ 1_n4450);
assign 1_n8032 = 1_n7324 & 1_n6682;
assign 1_n631 = ~(1_n7298 ^ 1_n8266);
assign 1_n5983 = 1_n7195 & 1_n311;
assign 1_n5766 = ~1_n9856;
assign 1_n3774 = 1_n6407 | 1_n6732;
assign 1_n10207 = ~(1_n8208 ^ 1_n3873);
assign 1_n2564 = 1_n13201 & 1_n9915;
assign 1_n9725 = 1_n11347 | 1_n824;
assign 1_n6763 = ~(1_n2335 ^ 1_n12892);
assign 1_n1416 = ~1_n5320;
assign 1_n1672 = ~1_n5780;
assign 1_n480 = ~(1_n6701 ^ 1_n7844);
assign 1_n11440 = ~(1_n6427 ^ 1_n5886);
assign 1_n781 = 1_n7247 | 1_n10059;
assign 1_n12614 = 1_n1571 | 1_n2718;
assign 1_n9643 = ~(1_n96 | 1_n10390);
assign 1_n11020 = 1_n1790 | 1_n11686;
assign 1_n4839 = ~(1_n5552 ^ 1_n7367);
assign 1_n260 = ~(1_n11874 | 1_n2716);
assign 1_n6511 = 1_n12795 | 1_n8490;
assign 1_n8551 = ~(1_n1940 ^ 1_n11880);
assign 1_n6599 = ~(1_n1862 | 1_n6180);
assign 1_n11733 = ~(1_n12833 ^ 1_n4005);
assign 1_n11039 = 1_n2254 | 1_n8534;
assign 1_n7357 = 1_n1587 | 1_n3890;
assign 1_n7503 = 1_n6724 | 1_n7221;
assign 1_n5226 = ~1_n2498;
assign 1_n2477 = ~(1_n4572 ^ 1_n981);
assign 1_n9588 = 1_n3553 | 1_n4640;
assign 1_n11738 = ~1_n4847;
assign 1_n12465 = ~1_n5189;
assign 1_n3239 = ~1_n11390;
assign 1_n12013 = 1_n12104 & 1_n12018;
assign 1_n12191 = 1_n2338 | 1_n13148;
assign 1_n10195 = ~1_n9684;
assign 1_n966 = ~(1_n11095 ^ 1_n11243);
assign 1_n11271 = ~(1_n232 ^ 1_n1870);
assign 1_n13180 = ~(1_n9082 ^ 1_n9687);
assign 1_n4327 = ~(1_n10672 ^ 1_n11442);
assign 1_n11116 = ~(1_n6899 | 1_n7214);
assign 1_n3948 = ~(1_n8361 ^ 1_n6162);
assign 1_n9768 = ~(1_n1988 ^ 1_n6143);
assign 1_n4242 = ~(1_n8981 | 1_n13000);
assign 1_n4678 = 1_n9195 | 1_n1144;
assign 1_n202 = ~1_n12306;
assign 1_n8787 = 1_n4727 | 1_n13196;
assign 1_n7028 = ~(1_n1727 ^ 1_n4060);
assign 1_n10878 = 1_n1370 | 1_n4640;
assign 1_n1616 = 1_n10527 | 1_n12188;
assign 1_n1980 = ~(1_n7313 ^ 1_n3500);
assign 1_n12157 = ~(1_n2020 | 1_n5267);
assign 1_n10236 = ~(1_n10081 ^ 1_n7282);
assign 1_n8187 = 1_n8182 | 1_n3716;
assign 1_n11317 = ~(1_n8770 ^ 1_n2284);
assign 1_n12205 = 1_n8938 & 1_n8164;
assign 1_n2314 = 1_n7667 ^ 1_n12961;
assign 1_n10746 = 1_n4149 & 1_n7147;
assign 1_n3061 = ~(1_n11530 ^ 1_n9589);
assign 1_n4455 = ~1_n2771;
assign 1_n4540 = ~1_n7113;
assign 1_n1633 = ~(1_n1826 | 1_n9871);
assign 1_n7762 = 1_n11780 & 1_n5869;
assign 1_n1859 = ~(1_n6345 ^ 1_n8879);
assign 1_n9499 = 1_n12730 & 1_n6525;
assign 1_n7228 = ~(1_n1540 | 1_n8150);
assign 1_n1602 = 1_n11800 & 1_n5424;
assign 1_n7318 = 1_n5865 | 1_n4947;
assign 1_n2770 = ~(1_n1578 ^ 1_n8597);
assign 1_n4431 = ~(1_n7480 | 1_n11052);
assign 1_n5492 = ~(1_n4066 | 1_n12622);
assign 1_n11735 = 1_n10123 & 1_n10822;
assign 1_n2649 = 1_n13097 & 1_n1577;
assign 1_n12550 = 1_n3130 & 1_n12284;
assign 1_n81 = 1_n11581 | 1_n3328;
assign 1_n541 = 1_n10947 & 1_n2862;
assign 1_n6556 = 1_n6283 | 1_n11173;
assign 1_n7683 = ~1_n5889;
assign 1_n282 = 1_n13165 & 1_n8322;
assign 1_n4978 = 1_n5845 ^ 1_n8084;
assign 1_n3053 = 1_n12051 & 1_n2086;
assign 1_n11546 = 1_n11682 ^ 1_n5355;
assign 1_n6741 = 1_n8803 | 1_n2903;
assign 1_n856 = 1_n3646 | 1_n12273;
assign 1_n8113 = 1_n10973 & 1_n4153;
assign 1_n1076 = 1_n10447 | 1_n4979;
assign 1_n2362 = 1_n6024 | 1_n4915;
assign 1_n9871 = ~1_n10627;
assign 1_n4025 = 1_n2028 & 1_n5468;
assign 1_n1662 = 1_n693 & 1_n11453;
assign 1_n9890 = ~(1_n8648 ^ 1_n8774);
assign 1_n3114 = 1_n9832 & 1_n3683;
assign 1_n12373 = ~(1_n7437 ^ 1_n6762);
assign 1_n12954 = ~1_n5801;
assign 1_n6230 = ~(1_n12698 | 1_n2051);
assign 1_n10976 = ~(1_n11944 ^ 1_n4299);
assign 1_n6114 = ~(1_n10505 ^ 1_n6161);
assign 1_n5926 = 1_n8863 | 1_n4640;
assign 1_n3319 = 1_n11554 | 1_n1156;
assign 1_n11310 = 1_n5431 & 1_n440;
assign 1_n4432 = 1_n4464 | 1_n4640;
assign 1_n1056 = 1_n6914 | 1_n9615;
assign 1_n3682 = 1_n9017 | 1_n7723;
assign 1_n6013 = ~(1_n10820 ^ 1_n10763);
assign 1_n12951 = ~(1_n11327 | 1_n394);
assign 1_n13197 = ~(1_n1891 ^ 1_n10084);
assign 1_n804 = 1_n1644 & 1_n12646;
assign 1_n97 = ~1_n9887;
assign 1_n4439 = ~(1_n12511 ^ 1_n2966);
assign 1_n7363 = ~(1_n4659 ^ 1_n11507);
assign 1_n9894 = 1_n7135 | 1_n7075;
assign 1_n10230 = ~1_n10294;
assign 1_n12477 = ~(1_n4231 ^ 1_n2073);
assign 1_n10114 = ~1_n39;
assign 1_n1760 = ~(1_n2426 ^ 1_n9912);
assign 1_n8333 = ~(1_n5912 ^ 1_n1982);
assign 1_n6870 = 1_n7084 | 1_n2675;
assign 1_n9222 = ~(1_n9925 ^ 1_n6361);
assign 1_n1808 = ~(1_n1394 ^ 1_n3233);
assign 1_n8673 = 1_n425 & 1_n6205;
assign 1_n1994 = ~(1_n1286 ^ 1_n2617);
assign 1_n4022 = ~1_n12693;
assign 1_n11154 = 1_n5031 & 1_n1916;
assign 1_n5157 = ~1_n1364;
assign 1_n8010 = 1_n464 | 1_n1466;
assign 1_n13064 = ~(1_n4560 ^ 1_n12923);
assign 1_n2662 = 1_n3434 & 1_n4021;
assign 1_n10250 = ~1_n9535;
assign 1_n999 = ~(1_n4857 ^ 1_n9735);
assign 1_n9705 = 1_n8225 | 1_n1985;
assign 1_n2338 = ~1_n9906;
assign 1_n6629 = ~1_n3641;
assign 1_n3405 = ~(1_n5151 | 1_n7843);
assign 1_n10931 = 1_n9428 ^ 1_n13173;
assign 1_n11248 = 1_n5569 | 1_n4373;
assign 1_n404 = ~(1_n704 ^ 1_n11516);
assign 1_n977 = 1_n8174 | 1_n9075;
assign 1_n6412 = 1_n9581 | 1_n4230;
assign 1_n8681 = ~1_n7374;
assign 1_n9001 = 1_n115 | 1_n10871;
assign 1_n7587 = ~(1_n2794 | 1_n1467);
assign 1_n13186 = ~1_n12121;
assign 1_n10409 = ~(1_n11274 ^ 1_n10559);
assign 1_n4201 = ~1_n3677;
assign 1_n10632 = ~(1_n4879 ^ 1_n563);
assign 1_n6690 = 1_n8492 & 1_n6120;
assign 1_n7216 = ~1_n1724;
assign 1_n1921 = 1_n8453 & 1_n4825;
assign 1_n5832 = ~1_n6873;
assign 1_n7493 = 1_n9909 | 1_n7803;
assign 1_n11856 = ~(1_n4211 | 1_n7095);
assign 1_n1571 = 1_n438;
assign 1_n4685 = 1_n8173 | 1_n121;
assign 1_n5475 = ~(1_n5647 ^ 1_n1837);
assign 1_n12075 = ~(1_n8080 | 1_n10140);
assign 1_n9004 = ~(1_n3106 ^ 1_n7276);
assign 1_n10885 = 1_n2685 & 1_n7889;
assign 1_n10581 = 1_n6984 & 1_n1297;
assign 1_n808 = ~1_n5320;
assign 1_n8472 = ~1_n4862;
assign 1_n12983 = ~(1_n9082 | 1_n13074);
assign 1_n3604 = ~(1_n8949 ^ 1_n6637);
assign 1_n8375 = 1_n8401 & 1_n337;
assign 1_n8062 = ~(1_n10416 | 1_n11030);
assign 1_n2593 = ~(1_n5833 ^ 1_n10370);
assign 1_n12661 = 1_n1938 ^ 1_n12932;
assign 1_n5227 = 1_n3563 | 1_n11870;
assign 1_n1978 = 1_n2449 | 1_n8702;
assign 1_n12616 = ~(1_n3372 ^ 1_n7577);
assign 1_n10389 = 1_n2493 & 1_n4203;
assign 1_n5479 = ~1_n3894;
assign 1_n12798 = ~1_n10019;
assign 1_n3475 = ~(1_n10247 ^ 1_n2756);
assign 1_n11643 = ~1_n7516;
assign 1_n10945 = ~(1_n2389 ^ 1_n2051);
assign 1_n2842 = 1_n12224 | 1_n1144;
assign 1_n10103 = ~1_n61;
assign 1_n3454 = ~1_n8230;
assign 1_n5073 = 1_n8978 & 1_n9733;
assign 1_n9070 = ~1_n3192;
assign 1_n9399 = 1_n5871 ^ 1_n8974;
assign 1_n492 = 1_n2015 & 1_n1701;
assign 1_n9054 = 1_n13073 | 1_n3426;
assign 1_n1031 = ~(1_n529 ^ 1_n8705);
assign 1_n10251 = ~(1_n9375 ^ 1_n10204);
assign 1_n12966 = 1_n10512 ^ 1_n5827;
assign 1_n4562 = 1_n1998 & 1_n5357;
assign 1_n4773 = 1_n5214 & 1_n4330;
assign 1_n1317 = ~(1_n6418 | 1_n1738);
assign 1_n295 = 1_n7219 & 1_n7222;
assign 1_n2608 = 1_n172 | 1_n4973;
assign 1_n4003 = 1_n11227 & 1_n2676;
assign 1_n5354 = 1_n3078 & 1_n6952;
assign 1_n12395 = ~1_n8183;
assign 1_n484 = 1_n9810 | 1_n542;
assign 1_n3089 = ~(1_n605 | 1_n11395);
assign 1_n4769 = ~(1_n710 ^ 1_n3376);
assign 1_n9758 = ~(1_n3117 ^ 1_n7457);
assign 1_n304 = ~(1_n6144 | 1_n11621);
assign 1_n4368 = ~(1_n6643 ^ 1_n2845);
assign 1_n2084 = ~(1_n6465 ^ 1_n9647);
assign 1_n3363 = 1_n8621 | 1_n9935;
assign 1_n6824 = ~(1_n11824 | 1_n10658);
assign 1_n2401 = 1_n8173 | 1_n12395;
assign 1_n326 = ~(1_n1988 | 1_n10035);
assign 1_n2128 = ~(1_n4937 ^ 1_n6192);
assign 1_n3960 = 1_n5231 & 1_n7227;
assign 1_n3002 = ~(1_n10456 ^ 1_n7664);
assign 1_n7117 = 1_n3293 | 1_n947;
assign 1_n470 = 1_n7354 | 1_n5743;
assign 1_n7459 = 1_n1718 | 1_n7567;
assign 1_n6316 = 1_n3407 | 1_n1026;
assign 1_n7888 = ~1_n11123;
assign 1_n7221 = 1_n11940;
assign 1_n7313 = 1_n9729 ^ 1_n6758;
assign 1_n7918 = 1_n10005 | 1_n10117;
assign 1_n9234 = 1_n10465 | 1_n1463;
assign 1_n6284 = 1_n723 & 1_n10506;
assign 1_n8390 = 1_n5683 | 1_n12721;
assign 1_n7906 = 1_n121 | 1_n1869;
assign 1_n3635 = ~(1_n7328 | 1_n6025);
assign 1_n7469 = 1_n11420 | 1_n2363;
assign 1_n1404 = 1_n9760 & 1_n11392;
assign 1_n780 = ~(1_n4742 ^ 1_n3837);
assign 1_n12696 = ~(1_n10344 ^ 1_n70);
assign 1_n233 = 1_n621 | 1_n3246;
assign 1_n2481 = 1_n4400 & 1_n12285;
assign 1_n545 = ~1_n5594;
assign 1_n3291 = ~(1_n1901 ^ 1_n11874);
assign 1_n1953 = 1_n8466 & 1_n8233;
assign 1_n6899 = 1_n7906;
assign 1_n4801 = ~(1_n7131 ^ 1_n11136);
assign 1_n8524 = 1_n5748 & 1_n11221;
assign 1_n200 = 1_n8361 | 1_n6162;
assign 1_n2871 = 1_n9949 & 1_n11889;
assign 1_n12547 = ~(1_n386 ^ 1_n3369);
assign 1_n2570 = 1_n12836 | 1_n1819;
assign 1_n409 = ~(1_n10613 | 1_n10711);
assign 1_n511 = 1_n2872 | 1_n9159;
assign 1_n4682 = 1_n10981 & 1_n5187;
assign 1_n3724 = ~1_n11953;
assign 1_n10850 = ~(1_n6717 ^ 1_n291);
assign 1_n5826 = 1_n12490 | 1_n2059;
assign 1_n1237 = 1_n2018 & 1_n854;
assign 1_n5828 = 1_n2329 | 1_n1026;
assign 1_n5100 = ~(1_n3914 ^ 1_n8503);
assign 1_n5424 = 1_n5905 & 1_n6727;
assign 1_n8271 = 1_n11537 & 1_n9915;
assign 1_n6895 = ~(1_n7774 ^ 1_n11355);
assign 1_n3929 = ~(1_n12270 | 1_n12076);
assign 1_n10077 = 1_n8306 | 1_n11982;
assign 1_n10354 = 1_n5913 & 1_n6412;
assign 1_n7006 = 1_n10908 & 1_n8468;
assign 1_n2282 = 1_n845 | 1_n8563;
assign 1_n11568 = ~(1_n10850 ^ 1_n1486);
assign 1_n5293 = ~(1_n8674 ^ 1_n1403);
assign 1_n3467 = 1_n12357 | 1_n13133;
assign 1_n11599 = 1_n3281 | 1_n3981;
assign 1_n7572 = 1_n4267 & 1_n6152;
assign 1_n9018 = ~1_n11906;
assign 1_n6355 = ~1_n817;
assign 1_n2643 = 1_n11871 | 1_n3225;
assign 1_n8193 = 1_n6481 | 1_n3651;
assign 1_n8777 = ~1_n5962;
assign 1_n3229 = 1_n5004 & 1_n4314;
assign 1_n6016 = 1_n11542 | 1_n12695;
assign 1_n940 = 1_n712 | 1_n9136;
assign 1_n10385 = 1_n8210 & 1_n10310;
assign 1_n13108 = ~1_n761;
assign 1_n196 = ~1_n8134;
assign 1_n3936 = 1_n5086 | 1_n1741;
assign 1_n6906 = ~1_n4687;
assign 1_n879 = 1_n1823 | 1_n7704;
assign 1_n758 = ~(1_n3715 ^ 1_n8831);
assign 1_n2650 = ~(1_n2196 ^ 1_n1295);
assign 1_n4910 = ~1_n6244;
assign 1_n4272 = ~1_n11350;
assign 1_n11620 = 1_n10317 | 1_n12361;
assign 1_n12138 = 1_n10752 & 1_n10666;
assign 1_n10540 = ~(1_n1219 | 1_n4567);
assign 1_n8890 = 1_n5694 | 1_n5242;
assign 1_n752 = 1_n3428 | 1_n12695;
assign 1_n3625 = ~(1_n40 ^ 1_n7873);
assign 1_n350 = 1_n1588 & 1_n12536;
assign 1_n2664 = ~(1_n8328 ^ 1_n10434);
assign 1_n4602 = 1_n1335 | 1_n1089;
assign 1_n8100 = ~(1_n2911 ^ 1_n11506);
assign 1_n8440 = 1_n12294 | 1_n7435;
assign 1_n7611 = 1_n2443 & 1_n11641;
assign 1_n403 = ~(1_n6892 ^ 1_n9952);
assign 1_n10981 = 1_n8495 | 1_n8929;
assign 1_n4064 = 1_n9104 & 1_n4852;
assign 1_n2244 = ~(1_n862 ^ 1_n7895);
assign 1_n2232 = ~1_n4862;
assign 1_n10456 = ~(1_n8080 ^ 1_n1576);
assign 1_n909 = 1_n1757 & 1_n3409;
assign 1_n3917 = ~(1_n10242 | 1_n10050);
assign 1_n11309 = ~(1_n8683 ^ 1_n10208);
assign 1_n10915 = ~(1_n5690 | 1_n4032);
assign 1_n10171 = 1_n6412 | 1_n5913;
assign 1_n5070 = 1_n379 | 1_n12273;
assign 1_n6542 = ~(1_n11063 ^ 1_n8862);
assign 1_n9931 = ~1_n12482;
assign 1_n6705 = ~(1_n13054 ^ 1_n12084);
assign 1_n12604 = ~1_n9620;
assign 1_n11381 = 1_n7160 & 1_n4374;
assign 1_n10099 = 1_n7688 | 1_n12524;
assign 1_n6776 = 1_n3115 | 1_n597;
assign 1_n5290 = 1_n10032 | 1_n8030;
assign 1_n7864 = ~1_n2072;
assign 1_n10833 = ~(1_n3001 ^ 1_n12179);
assign 1_n5115 = 1_n5146 | 1_n3981;
assign 1_n4460 = 1_n12274 & 1_n5111;
assign 1_n918 = ~(1_n2900 ^ 1_n6793);
assign 1_n10309 = ~(1_n1655 | 1_n1482);
assign 1_n7438 = 1_n44 | 1_n3981;
assign 1_n5937 = ~(1_n3730 ^ 1_n9932);
assign 1_n2030 = 1_n4943 & 1_n2124;
assign 1_n1744 = ~1_n8203;
assign 1_n5027 = 1_n89 & 1_n1813;
assign 1_n1822 = ~(1_n1481 | 1_n7848);
assign 1_n4667 = ~(1_n11490 ^ 1_n6282);
assign 1_n11748 = 1_n7658 & 1_n8512;
assign 1_n4539 = 1_n12560 ^ 1_n7854;
assign 1_n11071 = ~(1_n472 ^ 1_n5260);
assign 1_n7691 = 1_n13024 & 1_n6887;
assign 1_n2734 = ~(1_n11663 ^ 1_n8269);
assign 1_n2556 = ~1_n8506;
assign 1_n23 = ~(1_n4629 ^ 1_n2643);
assign 1_n5824 = ~(1_n2874 ^ 1_n8635);
assign 1_n8391 = ~1_n2501;
assign 1_n12734 = ~1_n5371;
assign 1_n6760 = ~1_n13076;
assign 1_n9226 = ~(1_n6822 ^ 1_n10776);
assign 1_n1580 = ~(1_n12130 | 1_n12181);
assign 1_n9609 = 1_n19 & 1_n3549;
assign 1_n9687 = ~(1_n4074 ^ 1_n6232);
assign 1_n9691 = 1_n2165 | 1_n5409;
assign 1_n12972 = 1_n1943 | 1_n12519;
assign 1_n6123 = 1_n1052 | 1_n8563;
assign 1_n8040 = ~1_n4933;
assign 1_n12759 = 1_n6454 & 1_n1975;
assign 1_n1901 = ~1_n10459;
assign 1_n9799 = ~(1_n4934 | 1_n5084);
assign 1_n7684 = 1_n5163 | 1_n5242;
assign 1_n1049 = ~(1_n2260 ^ 1_n4446);
assign 1_n447 = 1_n6671 & 1_n6441;
assign 1_n5269 = ~(1_n5213 | 1_n12687);
assign 1_n8586 = 1_n3687 & 1_n1800;
assign 1_n9204 = 1_n3157 | 1_n8206;
assign 1_n2844 = 1_n3705 ^ 1_n5938;
assign 1_n7366 = 1_n6629 | 1_n1985;
assign 1_n8128 = 1_n7649 & 1_n7031;
assign 1_n3264 = 1_n4114 & 1_n11222;
assign 1_n10323 = ~(1_n2187 | 1_n2612);
assign 1_n2948 = 1_n5562 | 1_n3981;
assign 1_n11153 = 1_n10018 | 1_n121;
assign 1_n588 = ~1_n1393;
assign 1_n10487 = ~(1_n5020 | 1_n1512);
assign 1_n11772 = ~1_n8230;
assign 1_n1733 = ~1_n12627;
assign 1_n522 = ~(1_n2193 ^ 1_n4167);
assign 1_n5268 = ~1_n1160;
assign 1_n1006 = 1_n235 | 1_n4285;
assign 1_n13229 = ~1_n5543;
assign 1_n12234 = ~1_n7336;
assign 1_n13227 = ~(1_n9161 ^ 1_n1726);
assign 1_n4638 = 1_n1361 | 1_n6910;
assign 1_n9695 = 1_n5890 | 1_n4373;
assign 1_n7552 = ~(1_n10731 ^ 1_n7540);
assign 1_n2728 = 1_n11722 | 1_n7502;
assign 1_n4054 = 1_n6526 | 1_n1951;
assign 1_n55 = ~(1_n1223 ^ 1_n8189);
assign 1_n6529 = ~(1_n10479 ^ 1_n4522);
assign 1_n10597 = ~1_n6654;
assign 1_n5840 = 1_n2834 | 1_n5298;
assign 1_n1867 = 1_n11303 | 1_n4990;
assign 1_n9802 = ~(1_n4542 ^ 1_n12259);
assign 1_n646 = ~(1_n7696 ^ 1_n13230);
assign 1_n4825 = 1_n9889 & 1_n4841;
assign 1_n6193 = ~1_n8716;
assign 1_n9895 = 1_n5974 & 1_n3655;
assign 1_n8595 = ~(1_n1306 | 1_n1682);
assign 1_n2041 = ~1_n5729;
assign 1_n4990 = ~(1_n4789 | 1_n8467);
assign 1_n13034 = ~(1_n9158 ^ 1_n2288);
assign 1_n7304 = 1_n4338 & 1_n13093;
assign 1_n7484 = 1_n11542 | 1_n4373;
assign 1_n5777 = ~(1_n1489 ^ 1_n5281);
assign 1_n8819 = 1_n9284 & 1_n11660;
assign 1_n1178 = 1_n9702 | 1_n3225;
assign 1_n11124 = 1_n12473 | 1_n2530;
assign 1_n9109 = 1_n8758 | 1_n10285;
assign 1_n1475 = ~(1_n8590 ^ 1_n3035);
assign 1_n2624 = 1_n2111 | 1_n3162;
assign 1_n8343 = ~(1_n6042 | 1_n6829);
assign 1_n6322 = ~(1_n1074 ^ 1_n4893);
assign 1_n6979 = 1_n1268 | 1_n6885;
assign 1_n9965 = 1_n3514 & 1_n8191;
assign 1_n12673 = ~1_n3040;
assign 1_n10961 = 1_n6979 & 1_n57;
assign 1_n11703 = 1_n9389 | 1_n5061;
assign 1_n8962 = ~(1_n5385 ^ 1_n8636);
assign 1_n2227 = 1_n2542 | 1_n2287;
assign 1_n7512 = ~(1_n6947 ^ 1_n4511);
assign 1_n1360 = ~1_n4998;
assign 1_n9615 = 1_n534 & 1_n5416;
assign 1_n11051 = ~(1_n7782 ^ 1_n13038);
assign 1_n11845 = ~(1_n12861 ^ 1_n6440);
assign 1_n12678 = ~(1_n10296 ^ 1_n5145);
assign 1_n4709 = 1_n1252 ^ 1_n13165;
assign 1_n7661 = ~1_n2882;
assign 1_n5247 = 1_n7856 | 1_n9873;
assign 1_n5172 = 1_n12772 | 1_n4991;
assign 1_n6431 = ~(1_n61 ^ 1_n9896);
assign 1_n7326 = ~(1_n4392 ^ 1_n12893);
assign 1_n2915 = ~1_n7515;
assign 1_n9696 = ~(1_n591 | 1_n7554);
assign 1_n10984 = ~(1_n11862 ^ 1_n4129);
assign 1_n10562 = ~(1_n6235 ^ 1_n8802);
assign 1_n5873 = ~(1_n7162 ^ 1_n3672);
assign 1_n10628 = ~(1_n8071 ^ 1_n7799);
assign 1_n6142 = ~1_n10799;
assign 1_n3659 = ~(1_n6530 ^ 1_n9758);
assign 1_n7963 = ~1_n1497;
assign 1_n1440 = 1_n8724 | 1_n12064;
assign 1_n2894 = ~(1_n6855 ^ 1_n8832);
assign 1_n11394 = ~(1_n3175 ^ 1_n10769);
assign 1_n5079 = ~1_n9187;
assign 1_n878 = 1_n26 & 1_n1239;
assign 1_n3738 = ~(1_n10220 ^ 1_n5387);
assign 1_n11897 = ~(1_n6349 ^ 1_n11309);
assign 1_n802 = ~(1_n12457 | 1_n2810);
assign 1_n7677 = ~(1_n7573 ^ 1_n9219);
assign 1_n11595 = 1_n4986 | 1_n4694;
assign 1_n6709 = ~(1_n3657 ^ 1_n7650);
assign 1_n8330 = 1_n11049 ^ 1_n4320;
assign 1_n12190 = 1_n1286 | 1_n12736;
assign 1_n11040 = ~1_n5705;
assign 1_n12485 = ~(1_n9969 ^ 1_n6249);
assign 1_n7907 = ~1_n4909;
assign 1_n939 = 1_n8230 & 1_n9531;
assign 1_n10996 = ~(1_n8396 | 1_n11383);
assign 1_n6978 = 1_n8871 & 1_n7139;
assign 1_n5490 = ~1_n11190;
assign 1_n12364 = ~(1_n524 ^ 1_n5617);
assign 1_n12785 = 1_n1285 & 1_n12055;
assign 1_n11550 = 1_n2678 | 1_n5076;
assign 1_n12769 = ~(1_n13107 ^ 1_n5619);
assign 1_n7970 = 1_n7501 ^ 1_n9063;
assign 1_n4282 = ~(1_n509 ^ 1_n4882);
assign 1_n11977 = ~(1_n8099 ^ 1_n12766);
assign 1_n25 = ~(1_n4879 ^ 1_n8760);
assign 1_n4891 = ~1_n9738;
assign 1_n11364 = ~1_n726;
assign 1_n12886 = ~1_n1900;
assign 1_n7651 = ~(1_n11118 ^ 1_n6214);
assign 1_n60 = ~1_n9636;
assign 1_n8747 = ~(1_n2835 | 1_n6833);
assign 1_n11621 = ~1_n362;
assign 1_n3379 = ~(1_n12574 ^ 1_n5951);
assign 1_n3965 = ~1_n12605;
assign 1_n8579 = 1_n1908 & 1_n11279;
assign 1_n6767 = 1_n9144 | 1_n6870;
assign 1_n4764 = ~(1_n8772 ^ 1_n506);
assign 1_n814 = 1_n9140 & 1_n174;
assign 1_n387 = ~(1_n1060 ^ 1_n10159);
assign 1_n704 = ~(1_n463 ^ 1_n9961);
assign 1_n10245 = ~1_n4828;
assign 1_n5461 = ~1_n11537;
assign 1_n9703 = ~(1_n10051 | 1_n1140);
assign 1_n13164 = ~(1_n1903 ^ 1_n8375);
assign 1_n7334 = ~(1_n5892 ^ 1_n2030);
assign 1_n3017 = ~1_n8715;
assign 1_n10020 = 1_n8510 | 1_n12718;
assign 1_n8915 = 1_n11472 | 1_n6882;
assign 1_n11503 = 1_n5360 ^ 1_n7970;
assign 1_n1433 = 1_n9482 & 1_n12323;
assign 1_n9978 = 1_n4109 | 1_n964;
assign 1_n11839 = ~(1_n2034 ^ 1_n11150);
assign 1_n9125 = ~1_n11673;
assign 1_n12577 = ~(1_n7688 ^ 1_n12524);
assign 1_n8108 = ~1_n1165;
assign 1_n12943 = 1_n12595 & 1_n1881;
assign 1_n5395 = ~(1_n8846 ^ 1_n4440);
assign 1_n10918 = 1_n3126 | 1_n2958;
assign 1_n783 = ~1_n8841;
assign 1_n11921 = ~(1_n2432 ^ 1_n3521);
assign 1_n2587 = ~(1_n3964 ^ 1_n6879);
assign 1_n5128 = ~(1_n3568 ^ 1_n5641);
assign 1_n220 = ~(1_n3679 ^ 1_n7600);
assign 1_n11189 = ~(1_n8157 ^ 1_n9576);
assign 1_n742 = ~(1_n11012 | 1_n3674);
assign 1_n12700 = 1_n4397 & 1_n8165;
assign 1_n12814 = ~1_n4862;
assign 1_n11098 = ~(1_n7795 | 1_n3803);
assign 1_n12924 = ~(1_n10114 | 1_n11332);
assign 1_n11360 = 1_n9316 | 1_n10072;
assign 1_n7291 = ~1_n5729;
assign 1_n6913 = ~1_n5185;
assign 1_n11554 = ~(1_n12661 | 1_n10321);
assign 1_n6229 = 1_n6407 | 1_n6404;
assign 1_n11759 = ~1_n5389;
assign 1_n5613 = 1_n9289 | 1_n7831;
assign 1_n11542 = ~1_n9846;
assign 1_n7170 = 1_n321 | 1_n10319;
assign 1_n1863 = ~(1_n10183 | 1_n1949);
assign 1_n8516 = ~(1_n7959 ^ 1_n2529);
assign 1_n10314 = ~1_n2737;
assign 1_n10302 = ~(1_n11645 | 1_n2);
assign 1_n8351 = ~1_n1764;
assign 1_n8449 = 1_n10914 | 1_n7185;
assign 1_n2940 = ~(1_n7862 ^ 1_n7166);
assign 1_n13224 = ~(1_n678 ^ 1_n166);
assign 1_n7150 = ~(1_n612 | 1_n9986);
assign 1_n7890 = ~1_n5470;
assign 1_n6780 = ~(1_n2962 ^ 1_n1415);
assign 1_n89 = ~1_n6675;
assign 1_n8381 = 1_n5445 | 1_n5681;
assign 1_n6628 = ~(1_n12843 ^ 1_n8988);
assign 1_n6138 = ~1_n7539;
assign 1_n5619 = ~(1_n5280 | 1_n8439);
assign 1_n8976 = ~(1_n1418 ^ 1_n10875);
assign 1_n5383 = ~1_n8887;
assign 1_n7741 = ~1_n12853;
assign 1_n5880 = ~(1_n11715 ^ 1_n2968);
assign 1_n7047 = ~(1_n10120 | 1_n346);
assign 1_n8828 = ~(1_n2550 | 1_n9472);
assign 1_n10267 = ~(1_n6754 | 1_n8094);
assign 1_n6024 = 1_n2449 | 1_n6404;
assign 1_n2383 = 1_n3532 | 1_n9190;
assign 1_n8376 = 1_n11957 & 1_n4958;
assign 1_n10347 = ~(1_n10817 ^ 1_n8067);
assign 1_n2433 = 1_n11851 | 1_n157;
assign 1_n2851 = ~(1_n12545 ^ 1_n6631);
assign 1_n2568 = ~(1_n8124 | 1_n4262);
assign 1_n11068 = 1_n8987 & 1_n3508;
assign 1_n3552 = ~1_n1503;
assign 1_n11382 = 1_n1688 | 1_n1463;
assign 1_n1225 = ~(1_n7611 ^ 1_n6570);
assign 1_n12048 = ~(1_n8714 | 1_n11853);
assign 1_n8465 = ~(1_n6336 ^ 1_n8752);
assign 1_n4609 = ~(1_n695 | 1_n7483);
assign 1_n8619 = 1_n8599 | 1_n6468;
assign 1_n12332 = 1_n6875 | 1_n4373;
assign 1_n10593 = 1_n12914 | 1_n5917;
assign 1_n7939 = ~1_n9138;
assign 1_n7249 = ~1_n6385;
assign 1_n5194 = 1_n7135 | 1_n9195;
assign 1_n3979 = ~(1_n7064 | 1_n4250);
assign 1_n6454 = ~(1_n1598 ^ 1_n2273);
assign 1_n8363 = ~1_n3321;
assign 1_n273 = ~(1_n11674 ^ 1_n7092);
assign 1_n8052 = 1_n12412 & 1_n4174;
assign 1_n5495 = ~(1_n1764 | 1_n2213);
assign 1_n8469 = 1_n1594 & 1_n7337;
assign 1_n2236 = 1_n7880 | 1_n4230;
assign 1_n11027 = 1_n12225 | 1_n9012;
assign 1_n6301 = ~(1_n11452 ^ 1_n6815);
assign 1_n3722 = 1_n2057 & 1_n2882;
assign 1_n1941 = ~1_n6149;
assign 1_n11307 = 1_n10499 | 1_n6893;
assign 1_n1649 = ~1_n11816;
assign 1_n12779 = ~(1_n8882 ^ 1_n1850);
assign 1_n1670 = ~(1_n1240 ^ 1_n12630);
assign 1_n3935 = 1_n2581 | 1_n13108;
assign 1_n1605 = ~1_n951;
assign 1_n3886 = ~(1_n8229 | 1_n4633);
assign 1_n1807 = ~1_n10548;
assign 1_n3490 = 1_n6488 | 1_n12388;
assign 1_n11251 = 1_n8179 | 1_n7140;
assign 1_n7856 = 1_n8400 | 1_n5242;
assign 1_n3029 = 1_n1325 | 1_n5423;
assign 1_n2 = 1_n4365 & 1_n2507;
assign 1_n3271 = 1_n3932 & 1_n7015;
assign 1_n13075 = 1_n6132 | 1_n8783;
assign 1_n3558 = 1_n6378 & 1_n9325;
assign 1_n11131 = 1_n2386 & 1_n6899;
assign 1_n5767 = 1_n11274 & 1_n12993;
assign 1_n2853 = 1_n6928 & 1_n1711;
assign 1_n5012 = ~(1_n12976 ^ 1_n4341);
assign 1_n7243 = ~1_n8288;
assign 1_n8626 = ~1_n12916;
assign 1_n8186 = 1_n7376 | 1_n2455;
assign 1_n1880 = ~(1_n8565 ^ 1_n4938);
assign 1_n5618 = ~(1_n13093 ^ 1_n2436);
assign 1_n12496 = 1_n5611 | 1_n2544;
assign 1_n7957 = 1_n2963 & 1_n8010;
assign 1_n4234 = ~(1_n3496 ^ 1_n12862);
assign 1_n157 = 1_n9854 & 1_n11193;
assign 1_n3349 = ~(1_n3594 ^ 1_n4632);
assign 1_n5746 = ~1_n6904;
assign 1_n7902 = 1_n10045 | 1_n7935;
assign 1_n12704 = 1_n9905 & 1_n173;
assign 1_n871 = ~1_n12085;
assign 1_n2136 = ~1_n1130;
assign 1_n6337 = 1_n9730 | 1_n11479;
assign 1_n5066 = ~1_n7710;
assign 1_n12239 = ~(1_n12162 ^ 1_n511);
assign 1_n12484 = ~1_n5408;
assign 1_n836 = 1_n10279 ^ 1_n9447;
assign 1_n3819 = ~1_n10563;
assign 1_n9587 = ~(1_n1284 ^ 1_n12369);
assign 1_n5698 = ~(1_n10073 ^ 1_n731);
assign 1_n12892 = ~(1_n2913 ^ 1_n10747);
assign 1_n9676 = ~(1_n3307 ^ 1_n11326);
assign 1_n6364 = ~1_n11488;
assign 1_n1951 = ~(1_n2937 ^ 1_n7764);
assign 1_n8599 = 1_n5949 | 1_n4230;
assign 1_n5351 = 1_n6883 | 1_n4947;
assign 1_n11003 = ~1_n3264;
assign 1_n193 = ~1_n2220;
assign 1_n6604 = 1_n81 & 1_n9884;
assign 1_n3764 = ~1_n9898;
assign 1_n5234 = 1_n9430 & 1_n2579;
assign 1_n9824 = ~(1_n1866 ^ 1_n2075);
assign 1_n5179 = 1_n10780 | 1_n8348;
assign 1_n7008 = 1_n7862 & 1_n9861;
assign 1_n4248 = 1_n2418 & 1_n9945;
assign 1_n12385 = ~(1_n729 | 1_n4700);
assign 1_n1423 = ~(1_n6280 ^ 1_n8121);
assign 1_n11617 = 1_n10901 | 1_n10687;
assign 1_n2303 = ~(1_n8489 ^ 1_n7853);
assign 1_n6068 = 1_n10587 | 1_n10871;
assign 1_n3663 = ~(1_n11997 ^ 1_n10062);
assign 1_n12285 = 1_n6129 | 1_n9075;
assign 1_n8948 = ~1_n7895;
assign 1_n8798 = ~(1_n2433 ^ 1_n5064);
assign 1_n6922 = ~1_n11350;
assign 1_n2145 = ~1_n938;
assign 1_n10695 = ~(1_n5131 ^ 1_n10397);
assign 1_n8358 = 1_n7950 | 1_n4936;
assign 1_n7835 = ~(1_n8957 ^ 1_n581);
assign 1_n7951 = 1_n1207 | 1_n7008;
assign 1_n11708 = 1_n9161 & 1_n6372;
assign 1_n4397 = 1_n7372 | 1_n4107;
assign 1_n284 = ~(1_n11283 ^ 1_n349);
assign 1_n8770 = 1_n12249 | 1_n5242;
assign 1_n2936 = ~(1_n3027 | 1_n3717);
assign 1_n4210 = ~(1_n484 ^ 1_n960);
assign 1_n1129 = ~(1_n2776 ^ 1_n6201);
assign 1_n3751 = ~(1_n1682 ^ 1_n4347);
assign 1_n7776 = 1_n12434 | 1_n479;
assign 1_n5099 = ~1_n3354;
assign 1_n11754 = 1_n895 & 1_n1639;
assign 1_n1312 = 1_n1296 | 1_n4936;
assign 1_n4021 = 1_n4540 | 1_n1463;
assign 1_n992 = 1_n10230 | 1_n8283;
assign 1_n8576 = 1_n2264 | 1_n11144;
assign 1_n1771 = 1_n8139 & 1_n6826;
assign 1_n5864 = 1_n8693 & 1_n709;
assign 1_n11357 = 1_n12528 | 1_n2694;
assign 1_n13038 = ~(1_n11915 ^ 1_n4133);
assign 1_n8539 = 1_n1416 | 1_n8868;
assign 1_n2837 = ~(1_n5503 ^ 1_n1452);
assign 1_n2855 = ~(1_n2842 ^ 1_n9484);
assign 1_n681 = ~(1_n1173 | 1_n3628);
assign 1_n6252 = ~(1_n2016 ^ 1_n9685);
assign 1_n9473 = ~(1_n10811 ^ 1_n10008);
assign 1_n10557 = ~(1_n3045 | 1_n8577);
assign 1_n6840 = 1_n1729 & 1_n6745;
assign 1_n7447 = ~(1_n8671 ^ 1_n1624);
assign 1_n3667 = ~(1_n4681 ^ 1_n11979);
assign 1_n797 = 1_n10527 | 1_n1463;
assign 1_n8231 = ~1_n346;
assign 1_n7093 = 1_n9967 & 1_n1442;
assign 1_n815 = 1_n313 & 1_n4212;
assign 1_n11994 = 1_n569 | 1_n2544;
assign 1_n3293 = ~1_n9475;
assign 1_n9742 = ~(1_n2585 ^ 1_n11238);
assign 1_n7287 = 1_n971 | 1_n5242;
assign 1_n2682 = ~(1_n5307 ^ 1_n709);
assign 1_n8490 = 1_n2557;
assign 1_n5597 = 1_n9069 | 1_n8534;
assign 1_n5482 = ~(1_n6165 | 1_n2448);
assign 1_n9810 = ~1_n401;
assign 1_n3274 = ~(1_n8223 ^ 1_n6520);
assign 1_n5718 = ~(1_n7953 ^ 1_n2871);
assign 1_n6144 = ~1_n6603;
assign 1_n12045 = ~1_n1771;
assign 1_n3338 = ~1_n4043;
assign 1_n12618 = ~(1_n11924 ^ 1_n7609);
assign 1_n5874 = 1_n4209 | 1_n7846;
assign 1_n3448 = 1_n4043 ^ 1_n1171;
assign 1_n9694 = ~(1_n1620 ^ 1_n2743);
assign 1_n11570 = 1_n4722 | 1_n8563;
assign 1_n7816 = ~(1_n9731 ^ 1_n674);
assign 1_n4151 = ~(1_n8675 ^ 1_n6429);
assign 1_n9141 = 1_n12674 & 1_n1001;
assign 1_n12202 = ~(1_n11084 | 1_n4931);
assign 1_n10886 = ~1_n11324;
assign 1_n2349 = ~(1_n12218 ^ 1_n10283);
assign 1_n4133 = 1_n9266 & 1_n5822;
assign 1_n4659 = 1_n9808 | 1_n542;
assign 1_n12228 = ~(1_n7982 ^ 1_n3426);
assign 1_n7 = 1_n6033 | 1_n13242;
assign 1_n1866 = ~(1_n2496 ^ 1_n6696);
assign 1_n6593 = ~(1_n12662 ^ 1_n6691);
assign 1_n436 = ~1_n10048;
assign 1_n8134 = 1_n10958 | 1_n792;
assign 1_n2625 = ~1_n13014;
assign 1_n7482 = ~(1_n5700 ^ 1_n8278);
assign 1_n4147 = ~(1_n11281 | 1_n4702);
assign 1_n9083 = 1_n2129 | 1_n12062;
assign 1_n11184 = ~(1_n10001 ^ 1_n6673);
assign 1_n5707 = ~1_n4885;
assign 1_n7575 = 1_n9924 ^ 1_n5668;
assign 1_n4572 = ~(1_n3797 ^ 1_n4705);
assign 1_n7082 = ~1_n4249;
assign 1_n1393 = ~(1_n8924 ^ 1_n3439);
assign 1_n1250 = 1_n9767 | 1_n9195;
assign 1_n1195 = ~(1_n11717 ^ 1_n8608);
assign 1_n11193 = 1_n7422 | 1_n9178;
assign 1_n10524 = ~(1_n5253 ^ 1_n4860);
assign 1_n4081 = 1_n6638 | 1_n6635;
assign 1_n10412 = 1_n9511 | 1_n8348;
assign 1_n4202 = ~(1_n170 ^ 1_n12547);
assign 1_n7380 = ~(1_n5354 | 1_n1831);
assign 1_n1567 = ~(1_n1683 ^ 1_n12557);
assign 1_n11978 = ~(1_n299 | 1_n967);
assign 1_n13128 = 1_n11284 | 1_n1043;
assign 1_n5816 = ~(1_n7747 ^ 1_n1183);
assign 1_n12351 = ~(1_n2568 | 1_n1608);
assign 1_n9806 = 1_n11114 | 1_n12188;
assign 1_n5595 = ~1_n8332;
assign 1_n4083 = ~(1_n10847 ^ 1_n10061);
assign 1_n7693 = ~(1_n10806 | 1_n1489);
assign 1_n11878 = 1_n11861 | 1_n8016;
assign 1_n5425 = 1_n5146 | 1_n5242;
assign 1_n11419 = 1_n10859 | 1_n8209;
assign 1_n5314 = 1_n5935 | 1_n4854;
assign 1_n12334 = ~(1_n6248 ^ 1_n1016);
assign 1_n12093 = ~1_n9887;
assign 1_n9650 = ~1_n1734;
assign 1_n5108 = 1_n2971 | 1_n6684;
assign 1_n10050 = ~(1_n7850 | 1_n3329);
assign 1_n11380 = 1_n5163 | 1_n9223;
assign 1_n6583 = ~(1_n7028 ^ 1_n10542);
assign 1_n10332 = ~1_n4439;
assign 1_n11791 = ~(1_n7497 | 1_n3386);
assign 1_n8355 = 1_n8629 | 1_n1161;
assign 1_n6450 = ~(1_n6750 ^ 1_n7653);
assign 1_n10361 = ~1_n1758;
assign 1_n12960 = ~(1_n12703 ^ 1_n13046);
assign 1_n7451 = ~(1_n11714 ^ 1_n1772);
assign 1_n8659 = 1_n12155 | 1_n10362;
assign 1_n3337 = 1_n3382 & 1_n10640;
assign 1_n5545 = 1_n7401 | 1_n7855;
assign 1_n2321 = ~1_n3311;
assign 1_n11094 = ~1_n12372;
assign 1_n266 = 1_n5787 & 1_n735;
assign 1_n7476 = ~(1_n12619 ^ 1_n6115);
assign 1_n6217 = 1_n533 | 1_n1287;
assign 1_n9163 = ~(1_n10153 ^ 1_n9183);
assign 1_n163 = ~(1_n7463 | 1_n11884);
assign 1_n8397 = 1_n790 | 1_n12419;
assign 1_n1066 = ~(1_n2227 ^ 1_n7126);
assign 1_n5405 = ~(1_n4757 ^ 1_n11450);
assign 1_n26 = ~1_n4747;
assign 1_n3512 = ~(1_n6299 ^ 1_n1882);
assign 1_n5158 = ~1_n2343;
assign 1_n5297 = ~(1_n5380 | 1_n6524);
assign 1_n6091 = 1_n12656 & 1_n10807;
assign 1_n10801 = ~(1_n11698 ^ 1_n7492);
assign 1_n9426 = 1_n12495 & 1_n4772;
assign 1_n3078 = ~1_n8149;
assign 1_n62 = ~(1_n9334 ^ 1_n8456);
assign 1_n11675 = ~(1_n4614 ^ 1_n8014);
assign 1_n5015 = 1_n1989 | 1_n7377;
assign 1_n9693 = ~1_n8689;
assign 1_n1641 = ~(1_n1939 ^ 1_n381);
assign 1_n9822 = 1_n12665 & 1_n11091;
assign 1_n5289 = ~1_n2731;
assign 1_n4612 = ~1_n12065;
assign 1_n922 = ~(1_n7957 ^ 1_n9566);
assign 1_n6005 = 1_n6858 & 1_n3665;
assign 1_n4254 = ~(1_n5998 ^ 1_n724);
assign 1_n12723 = ~(1_n8328 | 1_n12508);
assign 1_n11368 = ~(1_n4651 | 1_n10210);
assign 1_n4377 = 1_n8661 & 1_n7529;
assign 1_n11385 = 1_n12462 | 1_n5092;
assign 1_n131 = ~(1_n12237 ^ 1_n9506);
assign 1_n4914 = ~(1_n10348 ^ 1_n7590);
assign 1_n1375 = 1_n13036 | 1_n10871;
assign 1_n1016 = ~(1_n120 ^ 1_n12028);
assign 1_n6029 = 1_n8412 | 1_n273;
assign 1_n6830 = 1_n2002 | 1_n2308;
assign 1_n3976 = ~(1_n1984 ^ 1_n4483);
assign 1_n4457 = 1_n9706 & 1_n412;
assign 1_n685 = 1_n5038 | 1_n11368;
assign 1_n9935 = ~(1_n4128 ^ 1_n9982);
assign 1_n10078 = 1_n7715 & 1_n3409;
assign 1_n3585 = ~(1_n10774 | 1_n11777);
assign 1_n2983 = ~(1_n10238 ^ 1_n6286);
assign 1_n7848 = 1_n343 & 1_n9750;
assign 1_n4997 = ~(1_n6835 ^ 1_n3476);
assign 1_n2641 = ~1_n10805;
assign 1_n3068 = ~1_n2341;
assign 1_n285 = ~(1_n12632 | 1_n3990);
assign 1_n7478 = ~(1_n9970 ^ 1_n8625);
assign 1_n9654 = 1_n7087 ^ 1_n3008;
assign 1_n5138 = 1_n13231 | 1_n6128;
assign 1_n11450 = 1_n1695 | 1_n6635;
assign 1_n6987 = 1_n11213 & 1_n11241;
assign 1_n5018 = 1_n7925 | 1_n5242;
assign 1_n5879 = ~(1_n6455 ^ 1_n2724);
assign 1_n1299 = ~(1_n10799 ^ 1_n4097);
assign 1_n13077 = ~1_n9093;
assign 1_n9035 = 1_n11184 & 1_n7503;
assign 1_n12126 = ~1_n9531;
assign 1_n9356 = 1_n11933 | 1_n8702;
assign 1_n121 = 1_n12335;
assign 1_n8891 = 1_n3498 | 1_n905;
assign 1_n8041 = 1_n2961 & 1_n9142;
assign 1_n3714 = 1_n12732 | 1_n9075;
assign 1_n4465 = ~1_n287;
assign 1_n10701 = 1_n11065 & 1_n8708;
assign 1_n269 = ~(1_n12505 | 1_n9787);
assign 1_n9193 = ~(1_n1265 ^ 1_n8804);
assign 1_n7535 = ~(1_n1628 | 1_n3202);
assign 1_n2445 = 1_n2469 & 1_n2383;
assign 1_n6982 = 1_n6850 & 1_n4229;
assign 1_n4775 = ~(1_n7235 ^ 1_n7703);
assign 1_n1428 = 1_n2670 | 1_n546;
assign 1_n2395 = ~(1_n3942 ^ 1_n3089);
assign 1_n621 = 1_n1040 & 1_n5564;
assign 1_n8078 = 1_n609 & 1_n4677;
assign 1_n6140 = 1_n10168 & 1_n12263;
assign 1_n7714 = ~(1_n636 | 1_n9365);
assign 1_n6559 = ~1_n11134;
assign 1_n11562 = 1_n493 | 1_n1144;
assign 1_n5341 = ~1_n7036;
assign 1_n13059 = 1_n5120 & 1_n8474;
assign 1_n8294 = ~(1_n8052 ^ 1_n11038);
assign 1_n9116 = ~(1_n8422 | 1_n7407);
assign 1_n7360 = ~(1_n6311 ^ 1_n11568);
assign 1_n9084 = 1_n6710 | 1_n1197;
assign 1_n10440 = ~1_n3438;
assign 1_n1692 = 1_n5957 & 1_n8808;
assign 1_n6578 = ~1_n12186;
assign 1_n6966 = ~1_n9258;
assign 1_n3913 = 1_n8637 ^ 1_n10569;
assign 1_n10397 = ~(1_n2079 ^ 1_n11153);
assign 1_n2830 = ~(1_n7580 ^ 1_n4985);
assign 1_n3446 = ~(1_n786 ^ 1_n5484);
assign 1_n13172 = 1_n9340 & 1_n142;
assign 1_n2078 = ~(1_n1742 ^ 1_n6893);
assign 1_n1241 = 1_n12410 & 1_n2802;
assign 1_n11070 = ~(1_n1443 ^ 1_n6496);
assign 1_n1858 = ~1_n4636;
assign 1_n7470 = 1_n12575 | 1_n5623;
assign 1_n13195 = 1_n7481 & 1_n10644;
assign 1_n1111 = 1_n7686 & 1_n4508;
assign 1_n4166 = ~1_n1198;
assign 1_n3536 = 1_n9245 & 1_n12866;
assign 1_n6943 = 1_n406 | 1_n11446;
assign 1_n10279 = 1_n9628 & 1_n7459;
assign 1_n4555 = 1_n2512 & 1_n12237;
assign 1_n5330 = ~(1_n1481 ^ 1_n11848);
assign 1_n5805 = ~1_n5605;
assign 1_n11128 = ~(1_n7601 | 1_n3779);
assign 1_n10804 = 1_n5540 & 1_n1917;
assign 1_n6512 = 1_n1056 & 1_n3582;
assign 1_n9782 = 1_n10281 | 1_n2675;
assign 1_n9589 = ~(1_n2492 ^ 1_n250);
assign 1_n8076 = ~(1_n6763 | 1_n10440);
assign 1_n1236 = ~1_n7378;
assign 1_n645 = ~1_n4570;
assign 1_n12434 = ~1_n8522;
assign 1_n9006 = ~(1_n2072 ^ 1_n12283);
assign 1_n4404 = ~(1_n8970 ^ 1_n12701);
assign 1_n3299 = ~1_n7061;
assign 1_n5140 = ~(1_n2912 ^ 1_n4900);
assign 1_n2831 = 1_n7707 | 1_n4947;
assign 1_n7197 = 1_n9712 & 1_n1592;
assign 1_n5082 = ~1_n8794;
assign 1_n3033 = 1_n8081 & 1_n13191;
assign 1_n4974 = ~1_n6655;
assign 1_n5641 = ~(1_n13169 ^ 1_n3083);
assign 1_n9013 = 1_n8940 & 1_n287;
assign 1_n8263 = 1_n8039 | 1_n360;
assign 1_n9221 = 1_n10586 | 1_n1199;
assign 1_n10144 = 1_n2720 | 1_n4160;
assign 1_n1327 = 1_n11076 ^ 1_n412;
assign 1_n12629 = ~1_n1198;
assign 1_n9509 = 1_n11736 | 1_n2695;
assign 1_n5663 = ~(1_n141 | 1_n13195);
assign 1_n10265 = 1_n13116 | 1_n3709;
assign 1_n1796 = 1_n4654 | 1_n1958;
assign 1_n3822 = 1_n3972 | 1_n11152;
assign 1_n8695 = 1_n5220 & 1_n11636;
assign 1_n4079 = 1_n2437 | 1_n6652;
assign 1_n2035 = ~(1_n3270 ^ 1_n13143);
assign 1_n5183 = ~(1_n11374 ^ 1_n9025);
assign 1_n10609 = 1_n7900 | 1_n8030;
assign 1_n12492 = ~(1_n5553 ^ 1_n3);
assign 1_n365 = 1_n9397 | 1_n9319;
assign 1_n10922 = ~(1_n8803 ^ 1_n12787);
assign 1_n7589 = 1_n6343 | 1_n10788;
assign 1_n10832 = 1_n1732 & 1_n10502;
assign 1_n2558 = ~(1_n8760 | 1_n3209);
assign 1_n12594 = ~(1_n2262 ^ 1_n4535);
assign 1_n8883 = 1_n6271 | 1_n7723;
assign 1_n7746 = ~(1_n3285 | 1_n7381);
assign 1_n7944 = ~(1_n12252 | 1_n5573);
assign 1_n9533 = ~(1_n10318 | 1_n530);
assign 1_n12307 = ~(1_n12681 ^ 1_n6685);
assign 1_n1827 = 1_n694 | 1_n12717;
assign 1_n11032 = 1_n7244 & 1_n7933;
assign 1_n8779 = 1_n737 | 1_n6404;
assign 1_n1962 = 1_n3713 | 1_n7962;
assign 1_n6658 = ~1_n6023;
assign 1_n355 = ~(1_n12168 | 1_n1890);
assign 1_n1718 = 1_n3431 ^ 1_n9717;
assign 1_n4308 = 1_n8254 | 1_n11107;
assign 1_n3054 = 1_n9131 | 1_n8030;
assign 1_n12006 = ~(1_n6508 ^ 1_n4199);
assign 1_n3879 = 1_n7265 & 1_n8789;
assign 1_n7699 = 1_n7742 | 1_n5076;
assign 1_n5811 = 1_n3809 | 1_n2290;
assign 1_n5519 = ~(1_n9817 ^ 1_n4014);
assign 1_n9604 = ~(1_n4130 | 1_n1627);
assign 1_n7441 = 1_n1779 | 1_n10132;
assign 1_n10137 = ~1_n11222;
assign 1_n1572 = ~(1_n6990 | 1_n974);
assign 1_n11255 = 1_n3425 & 1_n1028;
assign 1_n11974 = ~1_n25;
assign 1_n7022 = 1_n3419 | 1_n2035;
assign 1_n2274 = ~(1_n12867 ^ 1_n11079);
assign 1_n7879 = ~(1_n9819 ^ 1_n10555);
assign 1_n9085 = 1_n9693 | 1_n4325;
assign 1_n4239 = 1_n12009 | 1_n9223;
assign 1_n7793 = ~(1_n11050 ^ 1_n11401);
assign 1_n11747 = 1_n25 ^ 1_n10724;
assign 1_n1977 = 1_n12049 | 1_n7935;
assign 1_n5271 = ~1_n11634;
assign 1_n5940 = 1_n12456 | 1_n7180;
assign 1_n11653 = 1_n11356 | 1_n177;
assign 1_n11764 = ~(1_n4502 ^ 1_n9458);
assign 1_n7514 = ~(1_n7841 ^ 1_n5149);
assign 1_n5814 = 1_n11653 | 1_n13042;
assign 1_n9730 = ~1_n2555;
assign 1_n3865 = ~(1_n12042 ^ 1_n4256);
assign 1_n79 = ~1_n9531;
assign 1_n9974 = ~(1_n1299 ^ 1_n8312);
assign 1_n7206 = ~(1_n2371 ^ 1_n3269);
assign 1_n2999 = 1_n5563 | 1_n11032;
assign 1_n3958 = 1_n3761 | 1_n1014;
assign 1_n11074 = ~(1_n11780 ^ 1_n11758);
assign 1_n2201 = ~(1_n9363 | 1_n1566);
assign 1_n12908 = ~1_n6987;
assign 1_n8098 = ~1_n1683;
assign 1_n2491 = 1_n477 | 1_n5024;
assign 1_n5717 = 1_n9240 | 1_n7002;
assign 1_n9460 = ~1_n9115;
assign 1_n4805 = 1_n10113 & 1_n7113;
assign 1_n7721 = ~(1_n3659 | 1_n8260);
assign 1_n12073 = ~(1_n12740 ^ 1_n1748);
assign 1_n8615 = ~1_n8233;
assign 1_n6270 = ~(1_n9534 | 1_n3192);
assign 1_n9904 = 1_n10966 | 1_n2958;
assign 1_n433 = 1_n5248 | 1_n10299;
assign 1_n11150 = 1_n7868 | 1_n8348;
assign 1_n11750 = ~1_n4889;
assign 1_n12495 = ~(1_n551 ^ 1_n2142);
assign 1_n206 = 1_n2557;
assign 1_n10008 = ~1_n836;
assign 1_n10196 = 1_n11547 | 1_n3689;
assign 1_n10318 = ~1_n5972;
assign 1_n10272 = ~1_n10630;
assign 1_n11638 = 1_n12919 & 1_n10533;
assign 1_n340 = ~(1_n1888 ^ 1_n3464);
assign 1_n489 = 1_n7501 | 1_n11359;
assign 1_n2749 = ~(1_n1200 | 1_n7645);
assign 1_n1956 = 1_n10837 & 1_n1015;
assign 1_n9493 = 1_n7563 & 1_n7794;
assign 1_n12654 = 1_n9873 & 1_n7856;
assign 1_n12398 = ~(1_n4262 ^ 1_n8124);
assign 1_n5122 = 1_n2500 | 1_n1371;
assign 1_n5888 = 1_n4473 | 1_n8490;
assign 1_n12929 = ~(1_n2980 ^ 1_n794);
assign 1_n9432 = ~(1_n2978 | 1_n10443);
assign 1_n3520 = ~(1_n11671 | 1_n9062);
assign 1_n1998 = ~1_n3887;
assign 1_n7821 = 1_n9540 ^ 1_n9510;
assign 1_n7616 = 1_n7914 & 1_n12949;
assign 1_n8558 = 1_n4964 & 1_n1916;
assign 1_n6061 = ~(1_n7117 ^ 1_n7170);
assign 1_n12662 = ~(1_n1775 ^ 1_n6316);
assign 1_n2986 = ~(1_n5272 ^ 1_n5856);
assign 1_n5295 = 1_n11127 & 1_n2355;
assign 1_n11023 = ~(1_n4379 | 1_n2897);
assign 1_n11985 = 1_n4997 | 1_n3237;
assign 1_n5284 = 1_n1511 | 1_n7935;
assign 1_n3989 = ~(1_n6071 ^ 1_n10829);
assign 1_n7795 = ~(1_n12322 | 1_n12374);
assign 1_n9148 = ~1_n8916;
assign 1_n8934 = ~1_n11217;
assign 1_n9958 = ~(1_n7236 ^ 1_n2099);
assign 1_n8462 = 1_n8042 & 1_n2533;
assign 1_n516 = 1_n1319 | 1_n3984;
assign 1_n2552 = 1_n7607 & 1_n3501;
assign 1_n673 = 1_n4220 | 1_n4360;
assign 1_n10006 = 1_n12656 | 1_n10807;
assign 1_n6546 = ~(1_n5888 ^ 1_n9549);
assign 1_n4742 = ~1_n10105;
assign 1_n12677 = 1_n7880 | 1_n8348;
assign 1_n3924 = ~1_n4023;
assign 1_n8601 = 1_n2473 | 1_n11770;
assign 1_n586 = 1_n1449 & 1_n7852;
assign 1_n7510 = 1_n2468 | 1_n12489;
assign 1_n5528 = 1_n5959 | 1_n12889;
assign 1_n13166 = ~(1_n7686 ^ 1_n12436);
assign 1_n4683 = ~(1_n3741 | 1_n3551);
assign 1_n10672 = ~(1_n5680 | 1_n7200);
assign 1_n10427 = 1_n928 | 1_n3287;
assign 1_n10793 = ~1_n13020;
assign 1_n7058 = ~(1_n5929 ^ 1_n10215);
assign 1_n5655 = 1_n107 | 1_n5049;
assign 1_n11629 = 1_n4657 | 1_n6404;
assign 1_n11223 = 1_n6008 & 1_n10268;
assign 1_n6196 = 1_n8251 & 1_n12821;
assign 1_n4183 = ~(1_n6511 ^ 1_n10943);
assign 1_n10023 = 1_n9955 | 1_n10570;
assign 1_n7521 = 1_n12940 & 1_n7496;
assign 1_n5142 = 1_n12982 | 1_n3497;
assign 1_n3018 = 1_n5990 | 1_n4230;
assign 1_n6989 = ~(1_n6382 | 1_n10175);
assign 1_n13137 = ~(1_n10113 | 1_n1757);
assign 1_n6928 = 1_n1977 | 1_n9149;
assign 1_n3313 = 1_n8249 | 1_n6635;
assign 1_n5982 = ~(1_n6618 | 1_n10986);
assign 1_n11969 = ~1_n12923;
assign 1_n4892 = ~(1_n8749 ^ 1_n8761);
assign 1_n5134 = 1_n10944 | 1_n6706;
assign 1_n6585 = 1_n2057 & 1_n3076;
assign 1_n8508 = ~1_n8155;
assign 1_n9479 = 1_n227 | 1_n8268;
assign 1_n6781 = ~(1_n5794 ^ 1_n11753);
assign 1_n3354 = 1_n11157 | 1_n1463;
assign 1_n5029 = ~(1_n10485 | 1_n11856);
assign 1_n8149 = ~(1_n4905 ^ 1_n7757);
assign 1_n6429 = ~(1_n376 ^ 1_n3921);
assign 1_n4192 = 1_n7084 | 1_n9784;
assign 1_n1512 = ~(1_n11912 | 1_n9715);
assign 1_n219 = ~(1_n6065 | 1_n10852);
assign 1_n6925 = 1_n12856 & 1_n6821;
assign 1_n2468 = 1_n1714 & 1_n1475;
assign 1_n12741 = ~1_n13060;
assign 1_n696 = ~(1_n2479 ^ 1_n5078);
assign 1_n7880 = ~1_n5536;
assign 1_n11466 = ~1_n4006;
assign 1_n11492 = ~(1_n9869 ^ 1_n7168);
assign 1_n3364 = ~1_n5758;
assign 1_n3737 = ~(1_n10967 ^ 1_n13189);
assign 1_n2155 = 1_n5937 | 1_n4165;
assign 1_n971 = ~1_n389;
assign 1_n4131 = ~(1_n10339 | 1_n7005);
assign 1_n2619 = ~1_n4281;
assign 1_n9329 = ~(1_n91 ^ 1_n9196);
assign 1_n8616 = ~(1_n6610 ^ 1_n4069);
assign 1_n9988 = ~1_n824;
assign 1_n140 = ~(1_n2881 ^ 1_n2751);
assign 1_n9762 = 1_n3231 & 1_n4175;
assign 1_n12763 = 1_n10237 & 1_n6472;
assign 1_n4067 = ~(1_n5502 | 1_n11452);
assign 1_n998 = ~(1_n8629 ^ 1_n1852);
assign 1_n824 = 1_n9157 & 1_n11595;
assign 1_n5730 = ~(1_n7666 ^ 1_n2984);
assign 1_n7813 = 1_n4524 & 1_n9697;
assign 1_n6845 = 1_n13062 | 1_n6176;
assign 1_n9372 = 1_n37 & 1_n5224;
assign 1_n1661 = 1_n1329 | 1_n7723;
assign 1_n1584 = 1_n3166 & 1_n8687;
assign 1_n6627 = 1_n9930 | 1_n3980;
assign 1_n9957 = ~(1_n1699 ^ 1_n3731);
assign 1_n9566 = ~(1_n8351 ^ 1_n2213);
assign 1_n865 = 1_n10622 ^ 1_n13157;
assign 1_n12325 = ~(1_n10056 | 1_n1668);
assign 1_n826 = 1_n2306 & 1_n9247;
assign 1_n6692 = ~(1_n3510 | 1_n11906);
assign 1_n11927 = ~1_n12390;
assign 1_n5369 = 1_n2619 | 1_n8012;
assign 1_n3154 = ~(1_n4764 ^ 1_n7138);
assign 1_n3835 = 1_n8937 & 1_n1141;
assign 1_n8115 = 1_n8795 | 1_n2959;
assign 1_n11728 = 1_n2479 | 1_n8292;
assign 1_n10494 = ~(1_n6205 ^ 1_n425);
assign 1_n10748 = ~1_n8954;
assign 1_n561 = ~1_n3144;
assign 1_n1333 = ~1_n5984;
assign 1_n5559 = ~1_n4691;
assign 1_n8697 = ~1_n10867;
assign 1_n7984 = ~(1_n3478 ^ 1_n10464);
assign 1_n195 = ~(1_n5577 ^ 1_n12251);
assign 1_n11757 = ~1_n22;
assign 1_n1382 = ~(1_n3988 ^ 1_n2445);
assign 1_n1622 = ~(1_n32 ^ 1_n4020);
assign 1_n6408 = 1_n4521 & 1_n13099;
assign 1_n11669 = ~(1_n31 ^ 1_n5051);
assign 1_n4925 = ~(1_n7435 ^ 1_n7088);
assign 1_n1869 = ~1_n854;
assign 1_n9052 = ~(1_n5513 ^ 1_n10251);
assign 1_n2512 = ~(1_n11233 ^ 1_n7736);
assign 1_n2571 = ~(1_n4277 | 1_n3046);
assign 1_n12500 = 1_n4298 | 1_n8582;
assign 1_n3478 = 1_n5461 | 1_n6769;
assign 1_n471 = ~(1_n9401 ^ 1_n3930);
assign 1_n5191 = ~(1_n1493 | 1_n8624);
assign 1_n7114 = 1_n644 | 1_n7152;
assign 1_n9021 = ~(1_n9835 ^ 1_n804);
assign 1_n9546 = 1_n11633 & 1_n5829;
assign 1_n6089 = 1_n12336 & 1_n1267;
assign 1_n181 = 1_n588 | 1_n7585;
assign 1_n9224 = 1_n7110 | 1_n9052;
assign 1_n1104 = 1_n3381 | 1_n4819;
assign 1_n1889 = ~1_n11049;
assign 1_n2962 = 1_n8666 & 1_n6204;
assign 1_n10256 = ~1_n4470;
assign 1_n10367 = 1_n10717 & 1_n12874;
assign 1_n13061 = ~(1_n2771 ^ 1_n6168);
assign 1_n6090 = ~(1_n8785 ^ 1_n197);
assign 1_n6008 = ~1_n13006;
assign 1_n8419 = ~1_n7932;
assign 1_n9170 = ~1_n8713;
assign 1_n468 = ~(1_n3744 ^ 1_n9184);
assign 1_n6999 = 1_n5412 & 1_n10340;
assign 1_n2220 = 1_n1058 | 1_n12847;
assign 1_n8247 = ~(1_n7421 | 1_n981);
assign 1_n3119 = ~(1_n6794 | 1_n5812);
assign 1_n1510 = ~(1_n548 ^ 1_n2369);
assign 1_n8867 = ~(1_n2151 ^ 1_n105);
assign 1_n3897 = ~(1_n10905 ^ 1_n3626);
assign 1_n12944 = 1_n9396 | 1_n9311;
assign 1_n5588 = ~1_n10594;
assign 1_n8157 = 1_n11683 | 1_n11144;
assign 1_n8463 = ~1_n10142;
assign 1_n4229 = 1_n4271 | 1_n9348;
assign 1_n4094 = 1_n11078 | 1_n7837;
assign 1_n10435 = 1_n1145 | 1_n10892;
assign 1_n10266 = ~1_n12605;
assign 1_n11067 = 1_n5675 & 1_n4559;
assign 1_n7787 = ~1_n5453;
assign 1_n7128 = 1_n10402 | 1_n10319;
assign 1_n3234 = ~(1_n10785 ^ 1_n429);
assign 1_n3839 = 1_n11447 & 1_n12765;
assign 1_n11756 = 1_n5069 & 1_n123;
assign 1_n9536 = ~(1_n4663 ^ 1_n8056);
assign 1_n10855 = ~(1_n7920 | 1_n11034);
assign 1_n6623 = ~(1_n12039 ^ 1_n4182);
assign 1_n4844 = ~1_n10606;
assign 1_n6914 = 1_n7668 & 1_n8074;
assign 1_n13041 = 1_n4785 | 1_n7615;
assign 1_n6359 = 1_n10462 | 1_n4724;
assign 1_n6452 = 1_n552 | 1_n3376;
assign 1_n263 = 1_n971 | 1_n2958;
assign 1_n7644 = ~(1_n7690 ^ 1_n199);
assign 1_n3382 = 1_n4290 | 1_n6364;
assign 1_n11287 = ~(1_n8812 | 1_n5287);
assign 1_n12980 = 1_n6155 ^ 1_n10670;
assign 1_n6825 = ~1_n11112;
assign 1_n3020 = 1_n5194 | 1_n5272;
assign 1_n11033 = 1_n8529 | 1_n6404;
assign 1_n1000 = ~1_n1600;
assign 1_n7608 = ~1_n13060;
assign 1_n1286 = 1_n11096 ^ 1_n12424;
assign 1_n8097 = ~1_n2920;
assign 1_n9677 = ~1_n3121;
assign 1_n6601 = 1_n7561 & 1_n4970;
assign 1_n2223 = 1_n8379 | 1_n5273;
assign 1_n9540 = 1_n2420 | 1_n2287;
assign 1_n5376 = ~(1_n1507 | 1_n3519);
assign 1_n11046 = ~(1_n2184 ^ 1_n5486);
assign 1_n8861 = ~(1_n6688 ^ 1_n8471);
assign 1_n4042 = 1_n7791 & 1_n6469;
assign 1_n92 = ~(1_n823 ^ 1_n7928);
assign 1_n11037 = ~1_n5065;
assign 1_n6660 = ~(1_n1398 ^ 1_n1946);
assign 1_n5754 = ~(1_n6359 ^ 1_n4255);
assign 1_n10534 = ~(1_n7709 | 1_n3165);
assign 1_n7410 = ~1_n8735;
assign 1_n3110 = 1_n5249 & 1_n3614;
assign 1_n838 = ~(1_n6021 ^ 1_n8227);
assign 1_n4759 = 1_n391 | 1_n12978;
assign 1_n6555 = ~(1_n3171 ^ 1_n9665);
assign 1_n7790 = ~(1_n10904 ^ 1_n10777);
assign 1_n9522 = ~(1_n8881 ^ 1_n3596);
assign 1_n12764 = 1_n9162 | 1_n8702;
assign 1_n8013 = ~(1_n6740 ^ 1_n9141);
assign 1_n9878 = 1_n5152 | 1_n4495;
assign 1_n5334 = 1_n5990 | 1_n7221;
assign 1_n6309 = ~1_n11900;
assign 1_n3077 = 1_n182 | 1_n5295;
assign 1_n885 = ~(1_n477 ^ 1_n8554);
assign 1_n5859 = ~(1_n3441 | 1_n6909);
assign 1_n996 = 1_n5670 | 1_n7642;
assign 1_n4232 = 1_n11946 & 1_n11481;
assign 1_n12110 = ~(1_n2043 ^ 1_n5995);
assign 1_n13043 = ~1_n9941;
assign 1_n5806 = ~1_n1724;
assign 1_n6816 = ~(1_n7546 ^ 1_n3610);
assign 1_n4961 = ~(1_n8864 | 1_n2422);
assign 1_n539 = 1_n4594 & 1_n7588;
assign 1_n4730 = ~(1_n2304 | 1_n10961);
assign 1_n1491 = 1_n8455 ^ 1_n2229;
assign 1_n6387 = 1_n7599 & 1_n9037;
assign 1_n4244 = 1_n2883 & 1_n1506;
assign 1_n11918 = 1_n7041 | 1_n8348;
assign 1_n661 = 1_n373 & 1_n12309;
assign 1_n11659 = 1_n3628 & 1_n1173;
assign 1_n7234 = ~1_n12263;
assign 1_n4993 = ~(1_n7575 ^ 1_n8145);
assign 1_n9466 = 1_n5870 & 1_n528;
assign 1_n7737 = ~(1_n577 | 1_n2117);
assign 1_n1405 = ~(1_n7095 ^ 1_n9117);
assign 1_n4162 = ~(1_n2792 ^ 1_n12911);
assign 1_n3791 = ~1_n10811;
assign 1_n12442 = 1_n12384 & 1_n7383;
assign 1_n5775 = 1_n2769 & 1_n9660;
assign 1_n308 = ~1_n2539;
assign 1_n3107 = ~(1_n11865 ^ 1_n4895);
assign 1_n12901 = 1_n7890 | 1_n10761;
assign 1_n5077 = 1_n3839 | 1_n11346;
assign 1_n10862 = 1_n4021 | 1_n3434;
assign 1_n12987 = ~(1_n2940 ^ 1_n5741);
assign 1_n6665 = ~(1_n1095 ^ 1_n9028);
assign 1_n4635 = 1_n8882 | 1_n1850;
assign 1_n13071 = ~1_n4349;
assign 1_n13086 = ~1_n11537;
assign 1_n12120 = 1_n9590 & 1_n6509;
assign 1_n2535 = ~(1_n10373 ^ 1_n10091);
assign 1_n5195 = ~(1_n3050 ^ 1_n3170);
assign 1_n4390 = 1_n10462 | 1_n2133;
assign 1_n7254 = ~1_n11488;
assign 1_n7752 = 1_n11941 | 1_n8348;
assign 1_n7649 = 1_n11159 | 1_n10040;
assign 1_n4070 = ~(1_n9641 | 1_n4873);
assign 1_n4578 = ~(1_n11444 ^ 1_n3198);
assign 1_n8014 = ~(1_n455 ^ 1_n5104);
assign 1_n12857 = ~(1_n9830 ^ 1_n4283);
assign 1_n9251 = ~(1_n6505 | 1_n13037);
assign 1_n8786 = ~1_n862;
assign 1_n7292 = ~(1_n1807 | 1_n6281);
assign 1_n8245 = 1_n2332 | 1_n177;
assign 1_n10311 = 1_n9933 & 1_n7193;
assign 1_n10906 = 1_n8672 | 1_n9195;
assign 1_n8341 = ~1_n11079;
assign 1_n10087 = ~(1_n5181 ^ 1_n9295);
assign 1_n2865 = ~(1_n5102 ^ 1_n4051);
assign 1_n4072 = 1_n5695 | 1_n7339;
assign 1_n6216 = 1_n4850 & 1_n2499;
assign 1_n8302 = 1_n755 | 1_n12967;
assign 1_n12761 = ~(1_n10774 ^ 1_n5779);
assign 1_n4681 = ~(1_n10547 ^ 1_n7323);
assign 1_n5583 = ~1_n3152;
assign 1_n12233 = 1_n11137 | 1_n10319;
assign 1_n4979 = ~1_n6168;
assign 1_n7678 = ~1_n12025;
assign 1_n7875 = ~(1_n2435 ^ 1_n12554);
assign 1_n11848 = ~(1_n9750 ^ 1_n504);
assign 1_n11239 = ~1_n9531;
assign 1_n9439 = 1_n2736 | 1_n2659;
assign 1_n11254 = 1_n13001 & 1_n5155;
assign 1_n3013 = 1_n12786 | 1_n8534;
assign 1_n8061 = 1_n5595 | 1_n7530;
assign 1_n7959 = 1_n3945 & 1_n10495;
assign 1_n9655 = 1_n2482 & 1_n12853;
assign 1_n8949 = 1_n13012 | 1_n12188;
assign 1_n2821 = 1_n8183 & 1_n6085;
assign 1_n9248 = ~(1_n2813 ^ 1_n4691);
assign 1_n8648 = 1_n935 | 1_n2133;
assign 1_n4100 = ~(1_n4377 ^ 1_n5439);
assign 1_n1222 = 1_n1801 & 1_n2477;
assign 1_n4490 = ~1_n9915;
assign 1_n4448 = 1_n9486 & 1_n6738;
assign 1_n3744 = 1_n12469 | 1_n12957;
assign 1_n12131 = ~(1_n1580 | 1_n9463);
assign 1_n5298 = ~(1_n8651 ^ 1_n2951);
assign 1_n5343 = 1_n10142 & 1_n5962;
assign 1_n13112 = 1_n11336 & 1_n5318;
assign 1_n10022 = 1_n6016 | 1_n8782;
assign 1_n1832 = ~1_n6879;
assign 1_n7024 = ~(1_n5233 ^ 1_n12934);
assign 1_n6956 = 1_n10761 | 1_n4936;
assign 1_n2191 = 1_n1795 | 1_n8543;
assign 1_n3932 = 1_n11196 | 1_n9533;
assign 1_n7394 = 1_n2992 & 1_n11262;
assign 1_n1839 = ~(1_n3749 ^ 1_n801);
assign 1_n2672 = 1_n11576 & 1_n8839;
assign 1_n12974 = 1_n2902 & 1_n1189;
assign 1_n8424 = 1_n7191 | 1_n5939;
assign 1_n4056 = ~(1_n1025 | 1_n4482);
assign 1_n1140 = ~(1_n12229 ^ 1_n4019);
assign 1_n1787 = ~1_n10002;
assign 1_n1948 = ~(1_n10538 ^ 1_n5650);
assign 1_n10964 = 1_n667 | 1_n5693;
assign 1_n13014 = 1_n4981 | 1_n9110;
assign 1_n9649 = 1_n8060 | 1_n3229;
assign 1_n9452 = ~(1_n3458 ^ 1_n2964);
assign 1_n10664 = ~(1_n12204 | 1_n12235);
assign 1_n12206 = 1_n4039 | 1_n9188;
assign 1_n12312 = 1_n12483 | 1_n4194;
assign 1_n40 = ~(1_n6013 ^ 1_n5232);
assign 1_n11196 = ~(1_n159 ^ 1_n6154);
assign 1_n10414 = 1_n5200 & 1_n12979;
assign 1_n12842 = 1_n11624 & 1_n5338;
assign 1_n2517 = ~(1_n6310 | 1_n4414);
assign 1_n12329 = ~(1_n6460 ^ 1_n5362);
assign 1_n10796 = ~(1_n12707 ^ 1_n10699);
assign 1_n9279 = 1_n12092 | 1_n10982;
assign 1_n10716 = 1_n1925 | 1_n4407;
assign 1_n9120 = 1_n2480 & 1_n5877;
assign 1_n6000 = 1_n3354 | 1_n6730;
assign 1_n8423 = ~(1_n8742 | 1_n4816);
assign 1_n1608 = 1_n5665 & 1_n8454;
assign 1_n5803 = 1_n1589 | 1_n2133;
assign 1_n9344 = 1_n5732 & 1_n5504;
assign 1_n5236 = ~(1_n7697 ^ 1_n4615);
assign 1_n5067 = 1_n151 & 1_n7078;
assign 1_n5455 = ~1_n11429;
assign 1_n9301 = ~(1_n10865 | 1_n1004);
assign 1_n4628 = 1_n7437 & 1_n12124;
assign 1_n8162 = ~(1_n1469 | 1_n7054);
assign 1_n8006 = ~1_n5969;
assign 1_n5898 = 1_n2742 | 1_n90;
assign 1_n11059 = 1_n2085 & 1_n2149;
assign 1_n4174 = 1_n5322 | 1_n5222;
assign 1_n10772 = ~1_n12965;
assign 1_n3753 = 1_n10437 | 1_n11107;
assign 1_n10066 = ~1_n7945;
assign 1_n7185 = ~(1_n9508 | 1_n10910);
assign 1_n3369 = ~(1_n3192 ^ 1_n8515);
assign 1_n2942 = ~1_n11061;
assign 1_n1252 = 1_n7642 | 1_n479;
assign 1_n2363 = 1_n9305 | 1_n10179;
assign 1_n5468 = ~1_n11991;
assign 1_n7193 = 1_n2884 | 1_n5797;
assign 1_n546 = ~1_n6236;
assign 1_n4761 = 1_n9402 | 1_n4333;
assign 1_n3836 = 1_n4179 | 1_n2059;
assign 1_n5500 = 1_n2460 & 1_n4750;
assign 1_n547 = ~(1_n7161 | 1_n1144);
assign 1_n12818 = 1_n10233 & 1_n6218;
assign 1_n1126 = ~1_n9097;
assign 1_n8927 = 1_n1222 | 1_n10239;
assign 1_n10739 = ~1_n2023;
assign 1_n5789 = ~(1_n11711 | 1_n41);
assign 1_n3833 = 1_n5492 | 1_n13135;
assign 1_n7996 = 1_n6682 ^ 1_n6451;
assign 1_n799 = 1_n11512 & 1_n4869;
assign 1_n7461 = 1_n6401 | 1_n306;
assign 1_n11535 = ~1_n2595;
assign 1_n8562 = ~1_n3409;
assign 1_n6057 = 1_n349 | 1_n11283;
assign 1_n6225 = ~1_n4335;
assign 1_n4994 = ~(1_n8932 ^ 1_n9204);
assign 1_n9157 = 1_n689 | 1_n4626;
assign 1_n2373 = 1_n823 | 1_n4405;
assign 1_n9258 = 1_n3588 & 1_n5967;
assign 1_n11225 = ~1_n2174;
assign 1_n3809 = 1_n6222 & 1_n3101;
assign 1_n2638 = ~(1_n8920 ^ 1_n12678);
assign 1_n10820 = 1_n13141 & 1_n11088;
assign 1_n3348 = 1_n542 | 1_n2675;
assign 1_n6227 = ~(1_n386 | 1_n6482);
assign 1_n6686 = ~(1_n8850 ^ 1_n632);
assign 1_n2870 = 1_n7385 | 1_n12794;
assign 1_n1053 = ~(1_n2975 | 1_n12056);
assign 1_n12948 = ~1_n834;
assign 1_n771 = 1_n9129 | 1_n6404;
assign 1_n5907 = 1_n10182 & 1_n12532;
assign 1_n6004 = ~1_n4685;
assign 1_n10434 = 1_n8876 ^ 1_n3180;
assign 1_n6568 = ~1_n2233;
assign 1_n9392 = 1_n10893 | 1_n1144;
assign 1_n2835 = ~(1_n12553 | 1_n4350);
assign 1_n5845 = 1_n2462 | 1_n8563;
assign 1_n8077 = ~1_n11760;
assign 1_n10373 = 1_n4161 | 1_n7221;
assign 1_n8994 = 1_n2129 | 1_n7221;
assign 1_n9040 = 1_n7243 | 1_n11232;
assign 1_n12668 = 1_n12963 | 1_n4812;
assign 1_n12774 = 1_n9620 & 1_n8716;
assign 1_n2105 = 1_n9703 | 1_n9064;
assign 1_n1999 = ~1_n2445;
assign 1_n11881 = ~(1_n6467 ^ 1_n11112);
assign 1_n12887 = ~(1_n5394 ^ 1_n4140);
assign 1_n5423 = ~1_n8233;
assign 1_n1316 = ~(1_n11023 | 1_n3462);
assign 1_n12883 = ~(1_n3976 ^ 1_n1884);
assign 1_n2296 = ~1_n12289;
assign 1_n6224 = ~(1_n3623 ^ 1_n8917);
assign 1_n11732 = ~(1_n9258 ^ 1_n4234);
assign 1_n1769 = ~1_n12594;
assign 1_n5447 = ~(1_n1494 ^ 1_n9297);
assign 1_n8318 = 1_n8957 | 1_n581;
assign 1_n8249 = ~1_n5536;
assign 1_n4660 = ~1_n11607;
assign 1_n10962 = 1_n2851 & 1_n1072;
assign 1_n5327 = ~(1_n9150 | 1_n8743);
assign 1_n8974 = 1_n2068 & 1_n11109;
assign 1_n4016 = 1_n7396 | 1_n4230;
assign 1_n5628 = ~(1_n1408 ^ 1_n2239);
assign 1_n12710 = ~(1_n2143 | 1_n8527);
assign 1_n6312 = 1_n3827 & 1_n5021;
assign 1_n8563 = 1_n3169;
assign 1_n6087 = ~(1_n11371 ^ 1_n2336);
assign 1_n3646 = ~1_n3769;
assign 1_n302 = ~(1_n11590 ^ 1_n11205);
assign 1_n9188 = ~(1_n8412 ^ 1_n273);
assign 1_n7633 = ~(1_n3581 | 1_n6331);
assign 1_n950 = ~1_n7448;
assign 1_n9480 = ~(1_n3818 ^ 1_n12040);
assign 1_n8682 = ~(1_n11436 | 1_n5053);
assign 1_n6347 = ~(1_n12428 ^ 1_n4435);
assign 1_n13100 = ~(1_n8738 | 1_n5997);
assign 1_n6483 = ~(1_n6619 ^ 1_n637);
assign 1_n300 = 1_n4464 | 1_n11107;
assign 1_n2522 = ~(1_n11223 | 1_n3002);
assign 1_n11101 = ~1_n6668;
assign 1_n5547 = ~1_n9906;
assign 1_n12572 = 1_n8839 | 1_n11576;
assign 1_n2604 = ~1_n9412;
assign 1_n10689 = ~1_n10027;
assign 1_n11162 = ~(1_n12121 ^ 1_n10458);
assign 1_n7628 = ~(1_n9033 ^ 1_n12743);
assign 1_n864 = 1_n761 & 1_n11058;
assign 1_n3720 = 1_n11116 | 1_n7976;
assign 1_n795 = ~1_n11411;
assign 1_n573 = 1_n1065 ^ 1_n7238;
assign 1_n3340 = ~1_n7541;
assign 1_n9578 = 1_n1505 & 1_n2482;
assign 1_n2599 = ~1_n8290;
assign 1_n8568 = ~(1_n12518 | 1_n3041);
assign 1_n4520 = ~(1_n7311 ^ 1_n12438);
assign 1_n11088 = ~1_n5228;
assign 1_n5107 = ~1_n401;
assign 1_n5685 = ~1_n9092;
assign 1_n3314 = ~(1_n5523 ^ 1_n2818);
assign 1_n498 = 1_n7257 & 1_n3450;
assign 1_n11624 = 1_n12802 | 1_n4295;
assign 1_n4276 = 1_n11226 | 1_n10106;
assign 1_n3709 = 1_n8541 & 1_n1264;
assign 1_n534 = 1_n12971 | 1_n7344;
assign 1_n12470 = 1_n6313 & 1_n7321;
assign 1_n5681 = 1_n11847 & 1_n7469;
assign 1_n1099 = 1_n3553 | 1_n2544;
assign 1_n10219 = 1_n1370 | 1_n7075;
assign 1_n12078 = 1_n2416 | 1_n2133;
assign 1_n1057 = 1_n1214 ^ 1_n11861;
assign 1_n4958 = 1_n1394 | 1_n3233;
assign 1_n6176 = 1_n8510 | 1_n177;
assign 1_n1085 = 1_n7167 | 1_n7935;
assign 1_n7081 = 1_n3453 | 1_n5335;
assign 1_n13228 = ~1_n2898;
assign 1_n2179 = 1_n11674 | 1_n7092;
assign 1_n5837 = ~(1_n7554 ^ 1_n140);
assign 1_n1836 = 1_n2255 ^ 1_n9652;
assign 1_n2405 = ~(1_n7448 | 1_n194);
assign 1_n5994 = ~(1_n5730 ^ 1_n6122);
assign 1_n1610 = 1_n2326 & 1_n2267;
assign 1_n7756 = ~(1_n8001 | 1_n7352);
assign 1_n1781 = ~1_n2668;
assign 1_n5752 = 1_n6769 | 1_n6404;
assign 1_n8106 = 1_n11903 & 1_n5765;
assign 1_n2919 = ~1_n834;
assign 1_n8876 = 1_n12343 & 1_n768;
assign 1_n2420 = ~1_n2758;
assign 1_n1435 = 1_n7119 | 1_n1570;
assign 1_n8021 = ~(1_n7245 ^ 1_n7007);
assign 1_n6523 = 1_n1976 & 1_n7586;
assign 1_n12534 = ~(1_n4215 ^ 1_n3983);
assign 1_n477 = ~(1_n4016 ^ 1_n843);
assign 1_n10053 = 1_n997 & 1_n970;
assign 1_n7668 = ~(1_n7279 ^ 1_n4532);
assign 1_n405 = 1_n9569 & 1_n10746;
assign 1_n9745 = ~1_n287;
assign 1_n5093 = 1_n5801 & 1_n9475;
assign 1_n4514 = ~1_n3130;
assign 1_n2017 = ~(1_n1847 | 1_n10090);
assign 1_n12979 = ~(1_n2918 ^ 1_n7259);
assign 1_n3880 = 1_n5705 ^ 1_n10078;
assign 1_n5080 = ~1_n635;
assign 1_n10732 = ~(1_n3219 | 1_n739);
assign 1_n6184 = 1_n2678 | 1_n9195;
assign 1_n2257 = 1_n6503 | 1_n310;
assign 1_n8888 = 1_n8139 & 1_n5920;
assign 1_n7565 = 1_n11437 | 1_n10693;
assign 1_n4278 = 1_n4886 & 1_n7810;
assign 1_n4399 = 1_n8704 & 1_n10529;
assign 1_n7975 = 1_n9305 | 1_n7530;
assign 1_n3323 = ~(1_n486 ^ 1_n1341);
assign 1_n2269 = 1_n1234 | 1_n1934;
assign 1_n9428 = 1_n10761 | 1_n10433;
assign 1_n6974 = 1_n946 | 1_n1985;
assign 1_n8461 = ~(1_n8125 ^ 1_n1138);
assign 1_n12180 = ~1_n3860;
assign 1_n12479 = 1_n12592 & 1_n2882;
assign 1_n595 = ~(1_n10384 | 1_n384);
assign 1_n10713 = 1_n4132 | 1_n12847;
assign 1_n8918 = 1_n2204 & 1_n1546;
assign 1_n283 = 1_n13062 & 1_n6176;
assign 1_n9406 = ~(1_n3155 | 1_n8656);
assign 1_n4901 = 1_n1524 | 1_n9778;
assign 1_n1010 = ~(1_n1862 ^ 1_n1283);
assign 1_n5945 = ~(1_n10859 ^ 1_n11631);
assign 1_n8327 = 1_n12899 & 1_n7710;
assign 1_n10894 = 1_n9806 | 1_n7224;
assign 1_n6946 = 1_n11195 | 1_n10110;
assign 1_n6718 = ~(1_n10543 ^ 1_n10955);
assign 1_n3212 = ~(1_n2160 ^ 1_n6198);
assign 1_n1477 = ~1_n7359;
assign 1_n2637 = ~1_n11030;
assign 1_n10033 = ~(1_n6925 ^ 1_n9394);
assign 1_n6275 = 1_n3669 & 1_n3085;
assign 1_n149 = 1_n12159 | 1_n8374;
assign 1_n3207 = ~(1_n10198 ^ 1_n2832);
assign 1_n9883 = ~(1_n4170 ^ 1_n1631);
assign 1_n9908 = ~(1_n5331 ^ 1_n2518);
assign 1_n4269 = 1_n10113 & 1_n12853;
assign 1_n892 = 1_n5088 & 1_n5814;
assign 1_n2150 = 1_n11899 & 1_n383;
assign 1_n2715 = 1_n12592 & 1_n11058;
assign 1_n8724 = 1_n1866 & 1_n8420;
assign 1_n9264 = 1_n5176 | 1_n7868;
assign 1_n11078 = ~1_n6168;
assign 1_n12362 = 1_n12741 | 1_n8702;
assign 1_n2365 = ~(1_n5193 ^ 1_n5643);
assign 1_n12988 = 1_n3829 & 1_n11685;
assign 1_n3355 = 1_n12268 | 1_n12401;
assign 1_n11245 = 1_n2688 | 1_n10179;
assign 1_n1529 = 1_n8102 ^ 1_n7717;
assign 1_n13094 = ~1_n1983;
assign 1_n7601 = ~(1_n8284 | 1_n4543);
assign 1_n12062 = ~1_n2590;
assign 1_n628 = ~1_n12289;
assign 1_n2785 = 1_n10730 | 1_n479;
assign 1_n9184 = 1_n1188 | 1_n4230;
assign 1_n3342 = 1_n6333 & 1_n10063;
assign 1_n11794 = 1_n7502 & 1_n11722;
assign 1_n1682 = ~(1_n10255 ^ 1_n12985);
assign 1_n10982 = ~1_n11027;
assign 1_n12649 = ~(1_n7472 | 1_n10723);
assign 1_n12680 = ~1_n1660;
assign 1_n9263 = 1_n11523 | 1_n6230;
assign 1_n1159 = ~(1_n10786 | 1_n7452);
assign 1_n12177 = ~(1_n7051 | 1_n12820);
assign 1_n466 = ~(1_n7904 ^ 1_n6);
assign 1_n1819 = ~(1_n5453 | 1_n9293);
assign 1_n2722 = ~1_n9163;
assign 1_n883 = 1_n6671 | 1_n6441;
assign 1_n10415 = ~(1_n10917 ^ 1_n4163);
assign 1_n6220 = ~1_n7812;
assign 1_n9315 = ~(1_n4667 ^ 1_n7423);
assign 1_n3777 = ~(1_n8595 | 1_n7753);
assign 1_n3954 = ~(1_n1714 ^ 1_n3788);
assign 1_n8146 = 1_n7408 | 1_n8869;
assign 1_n5986 = ~(1_n10656 | 1_n9292);
assign 1_n12204 = ~1_n1253;
assign 1_n6694 = 1_n11696 & 1_n7854;
assign 1_n9155 = 1_n4727 & 1_n13196;
assign 1_n12494 = ~(1_n6491 ^ 1_n8699);
assign 1_n4500 = ~(1_n12564 | 1_n295);
assign 1_n4603 = ~(1_n10533 ^ 1_n12919);
assign 1_n12156 = 1_n10199 & 1_n5579;
assign 1_n1837 = ~(1_n7673 ^ 1_n55);
assign 1_n4297 = ~(1_n1679 ^ 1_n7042);
assign 1_n2111 = 1_n4411 ^ 1_n388;
assign 1_n4255 = 1_n2491 & 1_n3529;
assign 1_n2471 = 1_n7674 | 1_n532;
assign 1_n3211 = 1_n11665 & 1_n2737;
assign 1_n12697 = 1_n5478 | 1_n479;
assign 1_n9658 = ~1_n2987;
assign 1_n4190 = ~(1_n1279 ^ 1_n5831);
assign 1_n4975 = 1_n10592 | 1_n1404;
assign 1_n11038 = ~(1_n11182 ^ 1_n2932);
assign 1_n1607 = 1_n7507 | 1_n3320;
assign 1_n3651 = ~1_n3875;
assign 1_n8628 = 1_n5568 & 1_n7113;
assign 1_n4556 = ~(1_n12631 | 1_n2421);
assign 1_n8783 = ~(1_n11561 | 1_n1423);
assign 1_n5017 = ~1_n12245;
assign 1_n257 = ~(1_n2429 ^ 1_n7014);
assign 1_n3365 = 1_n5838 | 1_n9587;
assign 1_n12522 = ~1_n1535;
assign 1_n10090 = ~1_n9419;
assign 1_n8354 = 1_n11334 & 1_n8627;
assign 1_n5123 = ~(1_n11699 ^ 1_n4806);
assign 1_n1728 = ~1_n646;
assign 1_n9309 = ~1_n5536;
assign 1_n2640 = ~1_n137;
assign 1_n2214 = 1_n10447 | 1_n5076;
assign 1_n5193 = ~(1_n7189 ^ 1_n5195);
assign 1_n12163 = 1_n4605 & 1_n4134;
assign 1_n647 = ~(1_n9425 ^ 1_n1146);
assign 1_n10366 = ~(1_n5706 ^ 1_n403);
assign 1_n5397 = ~(1_n9677 ^ 1_n2541);
assign 1_n1420 = ~1_n10333;
assign 1_n5957 = 1_n9890 | 1_n4343;
assign 1_n1746 = 1_n10306 & 1_n5114;
assign 1_n7316 = 1_n3338 & 1_n1171;
assign 1_n6847 = 1_n9783 & 1_n7391;
assign 1_n5653 = 1_n10839 | 1_n368;
assign 1_n679 = 1_n7522 | 1_n8268;
assign 1_n5098 = 1_n12871 | 1_n6265;
assign 1_n7559 = 1_n8310 & 1_n7187;
assign 1_n10419 = 1_n6756 & 1_n9565;
assign 1_n6926 = 1_n13221 ^ 1_n78;
assign 1_n6886 = 1_n5968 | 1_n8702;
assign 1_n686 = 1_n12881 | 1_n9195;
assign 1_n9683 = 1_n592 & 1_n914;
assign 1_n3115 = ~(1_n6492 ^ 1_n8217);
assign 1_n4360 = ~1_n5596;
assign 1_n8274 = 1_n12636 & 1_n7009;
assign 1_n11293 = ~(1_n2920 ^ 1_n11937);
assign 1_n8567 = 1_n10322 & 1_n4604;
assign 1_n6574 = ~(1_n1922 ^ 1_n11850);
assign 1_n9502 = 1_n4974 | 1_n12188;
assign 1_n8368 = 1_n6519 | 1_n12273;
assign 1_n8309 = ~(1_n5857 ^ 1_n6177);
assign 1_n7733 = 1_n4627 & 1_n3279;
assign 1_n4328 = ~(1_n4533 | 1_n12976);
assign 1_n5068 = ~(1_n9890 ^ 1_n8117);
assign 1_n10009 = ~(1_n5956 ^ 1_n6803);
assign 1_n10661 = ~1_n5404;
assign 1_n1060 = ~(1_n11773 ^ 1_n5026);
assign 1_n5390 = 1_n3970 | 1_n320;
assign 1_n7638 = 1_n5152 | 1_n10552;
assign 1_n9343 = ~(1_n1425 ^ 1_n4613);
assign 1_n4343 = 1_n12818 & 1_n7680;
assign 1_n12491 = ~1_n608;
assign 1_n11220 = ~(1_n10026 | 1_n4542);
assign 1_n4513 = 1_n5047 | 1_n10364;
assign 1_n10138 = 1_n12872 & 1_n12817;
assign 1_n6829 = 1_n7991 & 1_n3899;
assign 1_n9130 = ~(1_n246 | 1_n11942);
assign 1_n9496 = 1_n3534 | 1_n5242;
assign 1_n4731 = ~(1_n7011 ^ 1_n6061);
assign 1_n3632 = 1_n6466 & 1_n5512;
assign 1_n10782 = ~(1_n5799 ^ 1_n4721);
assign 1_n2877 = ~1_n12263;
assign 1_n776 = ~1_n10451;
assign 1_n5646 = ~(1_n7035 ^ 1_n4906);
assign 1_n1689 = ~(1_n7110 ^ 1_n7614);
assign 1_n2178 = 1_n3191 | 1_n3423;
assign 1_n10626 = 1_n951 & 1_n10063;
assign 1_n5769 = 1_n5365 & 1_n8749;
assign 1_n5208 = 1_n12813 & 1_n2361;
assign 1_n9626 = ~(1_n10236 | 1_n12438);
assign 1_n3016 = ~(1_n7550 ^ 1_n3948);
assign 1_n2598 = 1_n5611 | 1_n9159;
assign 1_n12796 = ~(1_n5669 ^ 1_n5568);
assign 1_n6110 = ~1_n649;
assign 1_n12621 = ~1_n3769;
assign 1_n2547 = 1_n6333 & 1_n3085;
assign 1_n5041 = ~1_n10168;
assign 1_n3618 = ~1_n12898;
assign 1_n9930 = 1_n11808 | 1_n6770;
assign 1_n10274 = 1_n11272 & 1_n5181;
assign 1_n8572 = ~(1_n8467 ^ 1_n1263);
assign 1_n12149 = ~(1_n4374 ^ 1_n7160);
assign 1_n5871 = 1_n12203 | 1_n9075;
assign 1_n11616 = 1_n9120 & 1_n1099;
assign 1_n4625 = 1_n3225 | 1_n12388;
assign 1_n2440 = ~1_n5143;
assign 1_n1485 = ~(1_n6171 | 1_n5532);
assign 1_n12066 = ~1_n11267;
assign 1_n10514 = ~(1_n3293 | 1_n10866);
assign 1_n1174 = ~(1_n4715 ^ 1_n913);
assign 1_n12144 = ~(1_n11335 ^ 1_n1280);
assign 1_n423 = ~1_n691;
assign 1_n7778 = 1_n5879 ^ 1_n13176;
assign 1_n7629 = 1_n2545 | 1_n9495;
assign 1_n9327 = ~(1_n11460 ^ 1_n4962);
assign 1_n3457 = ~(1_n8165 ^ 1_n12191);
assign 1_n9862 = ~(1_n1855 ^ 1_n11315);
assign 1_n9563 = ~(1_n191 ^ 1_n3378);
assign 1_n1368 = ~(1_n11963 | 1_n1924);
assign 1_n7007 = ~(1_n4346 | 1_n1643);
assign 1_n3407 = ~1_n11396;
assign 1_n3059 = ~(1_n1983 ^ 1_n4672);
assign 1_n6610 = 1_n7089 & 1_n12624;
assign 1_n4426 = ~1_n9621;
assign 1_n10104 = 1_n5359 | 1_n6987;
assign 1_n5267 = ~(1_n8513 | 1_n10750);
assign 1_n6489 = 1_n1089 | 1_n2449;
assign 1_n12823 = 1_n9298 & 1_n8127;
assign 1_n8265 = ~(1_n6317 ^ 1_n6134);
assign 1_n8715 = 1_n2449 | 1_n12328;
assign 1_n319 = ~(1_n7065 ^ 1_n2526);
assign 1_n9164 = ~(1_n10280 | 1_n8649);
assign 1_n9595 = 1_n1260 & 1_n8418;
assign 1_n3853 = ~1_n11055;
assign 1_n1873 = 1_n8788 ^ 1_n9202;
assign 1_n3199 = 1_n12668 & 1_n6449;
assign 1_n390 = 1_n3248 | 1_n65;
assign 1_n4221 = ~1_n5470;
assign 1_n4421 = ~(1_n408 | 1_n5472);
assign 1_n10738 = 1_n11664 | 1_n10715;
assign 1_n12012 = 1_n11003 | 1_n8044;
assign 1_n11091 = 1_n8139 & 1_n854;
assign 1_n7985 = ~(1_n11836 ^ 1_n5396);
assign 1_n11499 = 1_n5157 | 1_n6769;
assign 1_n12600 = 1_n9146 | 1_n11802;
assign 1_n12743 = ~(1_n5843 ^ 1_n6621);
assign 1_n4355 = ~(1_n10890 | 1_n4090);
assign 1_n6697 = 1_n5433 | 1_n8348;
assign 1_n1946 = ~(1_n1099 ^ 1_n9120);
assign 1_n7852 = 1_n9019 | 1_n12695;
assign 1_n6728 = 1_n13049 & 1_n13115;
assign 1_n857 = ~(1_n12055 ^ 1_n12900);
assign 1_n2789 = ~1_n10568;
assign 1_n5765 = ~(1_n9929 ^ 1_n5501);
assign 1_n5745 = 1_n1324 | 1_n4315;
assign 1_n12507 = ~(1_n7412 ^ 1_n5164);
assign 1_n4220 = ~1_n1617;
assign 1_n1524 = ~1_n3303;
assign 1_n3980 = 1_n6883 | 1_n10319;
assign 1_n2148 = ~1_n9591;
assign 1_n12050 = 1_n3259 | 1_n4936;
assign 1_n11075 = 1_n1034 & 1_n12777;
assign 1_n7458 = ~(1_n10262 ^ 1_n11504);
assign 1_n4649 = ~1_n5920;
assign 1_n11739 = ~(1_n5127 ^ 1_n10976);
assign 1_n9523 = ~(1_n9264 ^ 1_n2400);
assign 1_n10321 = ~1_n13053;
assign 1_n7496 = ~(1_n4770 ^ 1_n5777);
assign 1_n7763 = ~(1_n12192 ^ 1_n5571);
assign 1_n8279 = 1_n4798 & 1_n10519;
assign 1_n1303 = ~(1_n3214 | 1_n7173);
assign 1_n1905 = 1_n3599 | 1_n773;
assign 1_n12293 = 1_n1052 | 1_n3963;
assign 1_n3125 = ~(1_n7944 ^ 1_n8726);
assign 1_n12606 = ~(1_n12085 | 1_n2071);
assign 1_n12350 = ~(1_n1812 ^ 1_n3567);
assign 1_n8084 = 1_n5801 & 1_n5920;
assign 1_n5571 = 1_n11113 | 1_n2059;
assign 1_n4664 = 1_n9796 | 1_n11794;
assign 1_n1496 = 1_n1696 | 1_n1571;
assign 1_n1290 = ~1_n8328;
assign 1_n6241 = 1_n8889 | 1_n12068;
assign 1_n9815 = ~(1_n9529 ^ 1_n5963);
assign 1_n6471 = ~(1_n878 ^ 1_n6087);
assign 1_n3094 = ~1_n6292;
assign 1_n12023 = ~1_n401;
assign 1_n10300 = ~1_n9446;
assign 1_n4324 = ~(1_n12960 ^ 1_n611);
assign 1_n13118 = 1_n7295 & 1_n9530;
assign 1_n2578 = 1_n9004 | 1_n9946;
assign 1_n4580 = 1_n7957 | 1_n5495;
assign 1_n689 = 1_n4694 & 1_n4986;
assign 1_n1383 = 1_n6335 & 1_n6221;
assign 1_n3210 = ~1_n12943;
assign 1_n6441 = 1_n8315 | 1_n8348;
assign 1_n12666 = 1_n6556 & 1_n4635;
assign 1_n907 = 1_n9675 | 1_n12388;
assign 1_n11744 = 1_n8532 | 1_n7723;
assign 1_n1054 = 1_n8710 | 1_n10933;
assign 1_n478 = 1_n4316 & 1_n2924;
assign 1_n12917 = ~(1_n4241 | 1_n1794);
assign 1_n3553 = ~1_n12651;
assign 1_n11175 = 1_n11785 | 1_n639;
assign 1_n3050 = ~(1_n4159 | 1_n11532);
assign 1_n11709 = ~(1_n6962 ^ 1_n11918);
assign 1_n5450 = ~(1_n491 | 1_n2990);
assign 1_n579 = ~1_n12701;
assign 1_n5449 = 1_n586 | 1_n1770;
assign 1_n7913 = 1_n1491 | 1_n8242;
assign 1_n3962 = ~1_n3832;
assign 1_n6874 = 1_n3700 & 1_n7750;
assign 1_n6708 = ~(1_n10912 ^ 1_n572);
assign 1_n9101 = 1_n2420 | 1_n9159;
assign 1_n4793 = ~(1_n6880 ^ 1_n2957);
assign 1_n11805 = ~(1_n3212 ^ 1_n918);
assign 1_n1503 = 1_n2777 & 1_n9570;
assign 1_n6796 = 1_n12014 | 1_n653;
assign 1_n421 = 1_n2848 | 1_n1463;
assign 1_n12997 = ~1_n8506;
assign 1_n7311 = ~1_n10236;
assign 1_n2390 = 1_n5899 | 1_n8578;
assign 1_n10685 = ~(1_n3711 | 1_n7573);
assign 1_n11563 = ~(1_n6203 | 1_n2154);
assign 1_n12295 = ~1_n5065;
assign 1_n11264 = ~(1_n4682 ^ 1_n5985);
assign 1_n3785 = ~(1_n10441 | 1_n1355);
assign 1_n3395 = 1_n991 | 1_n8030;
assign 1_n9891 = ~1_n10643;
assign 1_n7239 = ~1_n12319;
assign 1_n10154 = 1_n8212 | 1_n9380;
assign 1_n6231 = ~1_n3112;
assign 1_n6940 = 1_n10938 | 1_n1841;
assign 1_n4454 = ~1_n510;
assign 1_n12113 = 1_n2952 & 1_n7444;
assign 1_n7865 = ~1_n4862;
assign 1_n7986 = ~1_n4711;
assign 1_n4339 = ~1_n386;
assign 1_n11752 = ~(1_n3011 ^ 1_n4935);
assign 1_n12877 = 1_n4802 | 1_n8493;
assign 1_n7368 = ~(1_n5090 | 1_n7638);
assign 1_n4212 = 1_n5766 | 1_n6080;
assign 1_n12804 = 1_n11928 | 1_n2059;
assign 1_n3701 = 1_n8285 & 1_n10933;
assign 1_n7129 = 1_n12736 & 1_n1286;
assign 1_n4630 = 1_n6707 ^ 1_n3760;
assign 1_n8236 = 1_n4561 | 1_n8607;
assign 1_n3479 = ~(1_n7830 ^ 1_n3875);
assign 1_n8222 = ~(1_n12333 ^ 1_n9194);
assign 1_n386 = ~(1_n7464 ^ 1_n4933);
assign 1_n6048 = ~(1_n8134 ^ 1_n2537);
assign 1_n1492 = ~(1_n5428 | 1_n11421);
assign 1_n1235 = ~(1_n12913 ^ 1_n10675);
assign 1_n7372 = ~1_n10657;
assign 1_n3845 = ~(1_n10184 ^ 1_n3391);
assign 1_n6711 = 1_n1345 | 1_n8632;
assign 1_n12474 = ~(1_n10328 ^ 1_n9715);
assign 1_n3564 = ~1_n4748;
assign 1_n101 = 1_n2951 | 1_n8651;
assign 1_n3623 = 1_n10761 | 1_n7530;
assign 1_n11609 = ~1_n10408;
assign 1_n6152 = 1_n7001 | 1_n8520;
assign 1_n11163 = 1_n2674 | 1_n10482;
assign 1_n9341 = ~(1_n2386 ^ 1_n12193);
assign 1_n12915 = 1_n10908 & 1_n5962;
assign 1_n11611 = ~1_n885;
assign 1_n10410 = 1_n1722 & 1_n4393;
assign 1_n3149 = ~1_n11324;
assign 1_n9137 = 1_n2771 & 1_n9093;
assign 1_n10255 = ~(1_n7910 ^ 1_n13092);
assign 1_n9089 = 1_n6861 & 1_n5465;
assign 1_n11850 = ~(1_n1235 ^ 1_n10494);
assign 1_n9598 = ~(1_n4489 | 1_n6462);
assign 1_n3404 = 1_n9867 | 1_n10029;
assign 1_n1522 = 1_n12367 | 1_n3673;
assign 1_n12458 = ~1_n4331;
assign 1_n1642 = ~(1_n8354 | 1_n6319);
assign 1_n5005 = 1_n5713 | 1_n9195;
assign 1_n299 = 1_n3392 & 1_n7979;
assign 1_n12685 = ~(1_n1150 ^ 1_n6005);
assign 1_n9573 = 1_n7266 | 1_n7060;
assign 1_n1181 = ~(1_n11852 ^ 1_n2876);
assign 1_n9624 = 1_n2229 & 1_n2207;
assign 1_n2010 = 1_n10015 & 1_n6608;
assign 1_n12181 = 1_n2641 | 1_n12657;
assign 1_n12822 = 1_n8993 & 1_n8250;
assign 1_n6045 = 1_n1521 | 1_n10272;
assign 1_n11578 = ~(1_n1449 ^ 1_n6702);
assign 1_n4688 = 1_n7226 & 1_n6912;
assign 1_n13157 = 1_n2404 & 1_n10325;
assign 1_n2799 = ~(1_n1506 ^ 1_n2883);
assign 1_n4679 = 1_n1434 | 1_n12657;
assign 1_n9211 = 1_n808 | 1_n1720;
assign 1_n9513 = 1_n12490 | 1_n8563;
assign 1_n3066 = ~(1_n1212 ^ 1_n4546);
assign 1_n2703 = 1_n5050 & 1_n5820;
assign 1_n9376 = ~(1_n1460 ^ 1_n6050);
assign 1_n9333 = ~(1_n11610 ^ 1_n12543);
assign 1_n4218 = 1_n3753 | 1_n6819;
assign 1_n9637 = 1_n3854 | 1_n4936;
assign 1_n327 = ~1_n9578;
assign 1_n9099 = 1_n9620 & 1_n3815;
assign 1_n5543 = 1_n2378 & 1_n8346;
assign 1_n4551 = 1_n30 & 1_n1419;
assign 1_n7937 = 1_n9367 & 1_n1357;
assign 1_n555 = ~(1_n1312 ^ 1_n12939);
assign 1_n8831 = ~(1_n10613 ^ 1_n10357);
assign 1_n6882 = ~(1_n3264 | 1_n1762);
assign 1_n10467 = 1_n4393 | 1_n1722;
assign 1_n4783 = ~1_n9125;
assign 1_n2085 = 1_n10560 & 1_n1724;
assign 1_n4385 = ~1_n5758;
assign 1_n3972 = ~1_n8506;
assign 1_n11737 = ~(1_n9613 ^ 1_n12534);
assign 1_n3525 = 1_n7416 & 1_n6722;
assign 1_n5484 = 1_n11566 & 1_n453;
assign 1_n4155 = ~(1_n3766 ^ 1_n12890);
assign 1_n4117 = 1_n10916 & 1_n11402;
assign 1_n10088 = ~(1_n8911 ^ 1_n7357);
assign 1_n3188 = ~(1_n17 ^ 1_n9327);
assign 1_n1028 = 1_n392 | 1_n177;
assign 1_n8385 = ~(1_n939 ^ 1_n1971);
assign 1_n1891 = ~(1_n11786 ^ 1_n2070);
assign 1_n10388 = 1_n6247 | 1_n11753;
assign 1_n8629 = ~(1_n585 ^ 1_n12835);
assign 1_n6215 = ~1_n5189;
assign 1_n9912 = ~(1_n3917 ^ 1_n7631);
assign 1_n12033 = 1_n9563 & 1_n12216;
assign 1_n12158 = ~(1_n10365 ^ 1_n10556);
assign 1_n3529 = 1_n3204 | 1_n4729;
assign 1_n5241 = ~(1_n10284 | 1_n6959);
assign 1_n11551 = ~(1_n1267 ^ 1_n9779);
assign 1_n9100 = ~(1_n5747 ^ 1_n3006);
assign 1_n11527 = ~(1_n2231 | 1_n9295);
assign 1_n11369 = ~1_n1472;
assign 1_n711 = ~(1_n6647 ^ 1_n6908);
assign 1_n3518 = ~(1_n1496 | 1_n5844);
assign 1_n982 = ~(1_n2898 ^ 1_n4688);
assign 1_n7266 = 1_n7905 & 1_n359;
assign 1_n2686 = ~(1_n10567 | 1_n2131);
assign 1_n12368 = ~1_n5352;
assign 1_n10439 = ~1_n3832;
assign 1_n2313 = ~(1_n4336 ^ 1_n12222);
assign 1_n7560 = ~1_n5197;
assign 1_n2263 = ~1_n6496;
assign 1_n2069 = ~(1_n12053 | 1_n8910);
assign 1_n12922 = 1_n7543 | 1_n931;
assign 1_n12555 = 1_n6880 | 1_n5072;
assign 1_n1471 = ~(1_n7650 | 1_n3657);
assign 1_n11195 = 1_n1820 | 1_n12273;
assign 1_n1251 = ~1_n1956;
assign 1_n1513 = ~(1_n1757 | 1_n10416);
assign 1_n2642 = ~(1_n7488 ^ 1_n4738);
assign 1_n9664 = 1_n11053 & 1_n4790;
assign 1_n7541 = 1_n6769 | 1_n10179;
assign 1_n6243 = 1_n7300 & 1_n11156;
assign 1_n12861 = 1_n3598 | 1_n9195;
assign 1_n2218 = ~(1_n10257 ^ 1_n2879);
assign 1_n3084 = 1_n10637 & 1_n9234;
assign 1_n4864 = ~(1_n481 ^ 1_n923);
assign 1_n11347 = ~1_n6107;
assign 1_n11479 = ~(1_n9123 ^ 1_n380);
assign 1_n1886 = 1_n123 | 1_n5069;
assign 1_n11671 = ~(1_n9826 ^ 1_n6090);
assign 1_n11478 = ~(1_n12931 ^ 1_n8641);
assign 1_n2147 = ~(1_n10882 ^ 1_n12906);
assign 1_n2879 = ~(1_n6121 ^ 1_n8282);
assign 1_n732 = ~(1_n9597 | 1_n9372);
assign 1_n4295 = 1_n2922 & 1_n281;
assign 1_n9816 = ~(1_n2523 | 1_n6237);
assign 1_n10759 = 1_n6996 & 1_n6614;
assign 1_n13081 = 1_n1406 | 1_n5797;
assign 1_n11810 = ~1_n8506;
assign 1_n7046 = 1_n4391 | 1_n6102;
assign 1_n135 = ~(1_n5903 ^ 1_n11955);
assign 1_n3998 = ~1_n8345;
assign 1_n8694 = 1_n11370 | 1_n7221;
assign 1_n2529 = ~(1_n11953 ^ 1_n6048);
assign 1_n1985 = 1_n3058;
assign 1_n318 = ~1_n9187;
assign 1_n147 = 1_n1587 | 1_n11668;
assign 1_n7204 = 1_n1629 | 1_n13020;
assign 1_n2033 = ~(1_n5844 ^ 1_n1496);
assign 1_n2576 = 1_n8582 & 1_n4298;
assign 1_n12933 = ~(1_n9142 ^ 1_n7740);
assign 1_n1093 = ~(1_n5342 ^ 1_n2609);
assign 1_n9097 = 1_n2781 & 1_n8440;
assign 1_n10875 = ~(1_n3767 ^ 1_n11257);
assign 1_n729 = ~(1_n4397 ^ 1_n3457);
assign 1_n12786 = ~1_n3769;
assign 1_n2788 = 1_n3528 | 1_n10918;
assign 1_n11346 = 1_n4189 & 1_n1799;
assign 1_n280 = 1_n3460 | 1_n10016;
assign 1_n2808 = 1_n8330 | 1_n5073;
assign 1_n9972 = ~1_n2037;
assign 1_n10777 = ~(1_n6357 ^ 1_n12602);
assign 1_n7163 = ~1_n10013;
assign 1_n7494 = 1_n12028 & 1_n120;
assign 1_n2048 = ~1_n6937;
assign 1_n2292 = 1_n11245 | 1_n9737;
assign 1_n5170 = 1_n8228 & 1_n13058;
assign 1_n10598 = 1_n2993 & 1_n10480;
assign 1_n11543 = 1_n7864 | 1_n3939;
assign 1_n43 = ~(1_n8571 ^ 1_n925);
assign 1_n5790 = ~(1_n1234 ^ 1_n1934);
assign 1_n7025 = ~1_n1143;
assign 1_n117 = 1_n1609 | 1_n11911;
assign 1_n893 = ~(1_n5007 ^ 1_n6977);
assign 1_n9724 = 1_n10432 | 1_n10403;
assign 1_n850 = 1_n10829 & 1_n6071;
assign 1_n1355 = ~(1_n4962 | 1_n10810);
assign 1_n9461 = ~1_n9277;
assign 1_n8607 = 1_n1314 & 1_n8177;
assign 1_n13194 = ~1_n4862;
assign 1_n3824 = ~(1_n3706 ^ 1_n1407);
assign 1_n2863 = 1_n11610 | 1_n1456;
assign 1_n12413 = 1_n3404 | 1_n10984;
assign 1_n1156 = 1_n1196 & 1_n2345;
assign 1_n7023 = 1_n12000 | 1_n8912;
assign 1_n6995 = 1_n8623 | 1_n10581;
assign 1_n1772 = 1_n9016 | 1_n1026;
assign 1_n10694 = ~(1_n4926 | 1_n5710);
assign 1_n748 = ~(1_n12745 ^ 1_n4092);
assign 1_n5439 = 1_n6810 | 1_n12501;
assign 1_n6609 = ~(1_n2477 ^ 1_n1801);
assign 1_n916 = ~(1_n2240 ^ 1_n1023);
assign 1_n398 = ~(1_n11217 | 1_n9601);
assign 1_n6403 = 1_n12220 | 1_n2100;
assign 1_n12821 = 1_n2215 & 1_n10052;
assign 1_n9685 = 1_n8959 & 1_n7106;
assign 1_n1347 = ~1_n1085;
assign 1_n5056 = ~(1_n7634 ^ 1_n9442);
assign 1_n165 = 1_n5874 | 1_n9122;
assign 1_n1717 = 1_n1548 & 1_n4176;
assign 1_n11960 = ~1_n9906;
assign 1_n11726 = ~(1_n6509 ^ 1_n9590);
assign 1_n7141 = ~(1_n6155 ^ 1_n179);
assign 1_n10026 = 1_n785 | 1_n8268;
assign 1_n6147 = ~(1_n3682 ^ 1_n4259);
assign 1_n6187 = 1_n7028 | 1_n2092;
assign 1_n1295 = ~(1_n12531 ^ 1_n2241);
assign 1_n3095 = 1_n6231 | 1_n1043;
assign 1_n5696 = 1_n3835 | 1_n10521;
assign 1_n1444 = ~(1_n4711 ^ 1_n8540);
assign 1_n4949 = ~1_n11030;
assign 1_n5175 = ~(1_n10869 ^ 1_n8359);
assign 1_n9284 = ~(1_n2334 ^ 1_n2316);
assign 1_n10656 = 1_n2432 & 1_n11637;
assign 1_n11941 = ~1_n510;
assign 1_n2047 = ~(1_n10090 ^ 1_n3086);
assign 1_n3217 = 1_n6483 & 1_n9448;
assign 1_n10000 = ~(1_n608 ^ 1_n3451);
assign 1_n6558 = 1_n8082 | 1_n12388;
assign 1_n10337 = ~(1_n12139 ^ 1_n3306);
assign 1_n3390 = 1_n9803 & 1_n6946;
assign 1_n9603 = 1_n6422 & 1_n11260;
assign 1_n4428 = ~(1_n366 ^ 1_n301);
assign 1_n6814 = ~1_n8183;
assign 1_n9867 = ~1_n7659;
assign 1_n7590 = ~(1_n11327 ^ 1_n394);
assign 1_n542 = 1_n3185;
assign 1_n11575 = 1_n12434 | 1_n2544;
assign 1_n9850 = ~(1_n12341 | 1_n7487);
assign 1_n1319 = 1_n11808 | 1_n3999;
assign 1_n2228 = ~1_n9915;
assign 1_n2586 = ~(1_n820 ^ 1_n4295);
assign 1_n953 = 1_n2748 | 1_n7353;
assign 1_n12226 = ~(1_n4117 ^ 1_n8321);
assign 1_n5555 = ~(1_n12194 ^ 1_n7727);
assign 1_n11469 = ~(1_n4650 ^ 1_n13102);
assign 1_n3794 = 1_n6945 & 1_n5108;
assign 1_n10338 = 1_n3714 | 1_n8552;
assign 1_n3614 = 1_n6448 | 1_n11806;
assign 1_n10374 = 1_n11150 & 1_n2034;
assign 1_n12871 = ~1_n10805;
assign 1_n5616 = 1_n1945 | 1_n1927;
assign 1_n5013 = 1_n2701 | 1_n8038;
assign 1_n1102 = 1_n771 | 1_n478;
assign 1_n2949 = 1_n11823 & 1_n4499;
assign 1_n2431 = 1_n3534 | 1_n121;
assign 1_n13083 = ~1_n9307;
assign 1_n9176 = 1_n4540 | 1_n10029;
assign 1_n1620 = ~(1_n4570 ^ 1_n3600);
assign 1_n12627 = 1_n64 & 1_n878;
assign 1_n8505 = ~1_n11030;
assign 1_n1033 = ~(1_n8550 | 1_n13119);
assign 1_n3131 = 1_n10024 & 1_n9481;
assign 1_n5103 = 1_n2661 | 1_n2575;
assign 1_n6700 = ~(1_n2753 ^ 1_n10846);
assign 1_n2061 = ~(1_n1637 ^ 1_n1844);
assign 1_n9939 = ~(1_n969 | 1_n7762);
assign 1_n5637 = ~(1_n4886 ^ 1_n7810);
assign 1_n9307 = ~(1_n7445 ^ 1_n9876);
assign 1_n11600 = 1_n4248 | 1_n3513;
assign 1_n5347 = 1_n9123 & 1_n8240;
assign 1_n1890 = 1_n5625 & 1_n9539;
assign 1_n162 = 1_n6954 | 1_n1556;
assign 1_n532 = 1_n5874 & 1_n9122;
assign 1_n7860 = ~(1_n1610 ^ 1_n6678);
assign 1_n1027 = ~(1_n2802 ^ 1_n11817);
assign 1_n12004 = 1_n8204 | 1_n8128;
assign 1_n4036 = 1_n3130 & 1_n1724;
assign 1_n5604 = 1_n12113 & 1_n8008;
assign 1_n6435 = ~(1_n6113 ^ 1_n11235);
assign 1_n5517 = 1_n8935 | 1_n12858;
assign 1_n11403 = 1_n8298 & 1_n1821;
assign 1_n8213 = ~(1_n4118 | 1_n8321);
assign 1_n1244 = 1_n616 | 1_n6117;
assign 1_n2807 = 1_n6519 | 1_n8534;
assign 1_n10747 = ~(1_n7856 ^ 1_n9873);
assign 1_n2231 = ~(1_n5181 | 1_n11272);
assign 1_n1230 = 1_n10314 | 1_n1043;
assign 1_n9123 = ~(1_n2384 ^ 1_n2873);
assign 1_n8322 = ~1_n1252;
assign 1_n3731 = 1_n13182 | 1_n5939;
assign 1_n7765 = ~1_n9905;
assign 1_n6346 = 1_n3594 | 1_n4632;
assign 1_n12851 = 1_n10756 | 1_n10871;
assign 1_n9417 = ~1_n4803;
assign 1_n2038 = 1_n317 & 1_n1557;
assign 1_n5958 = ~(1_n11039 | 1_n521);
assign 1_n2762 = 1_n3634 | 1_n8268;
assign 1_n11292 = 1_n1894 & 1_n6191;
assign 1_n6386 = ~(1_n12122 ^ 1_n11788);
assign 1_n6894 = 1_n7255 | 1_n5315;
assign 1_n1189 = ~1_n7706;
assign 1_n11547 = ~(1_n4740 ^ 1_n11952);
assign 1_n4645 = ~(1_n11050 ^ 1_n5046);
assign 1_n6260 = ~1_n7259;
assign 1_n12346 = 1_n13019 | 1_n507;
assign 1_n8454 = 1_n472 | 1_n1271;
assign 1_n11761 = 1_n8836 & 1_n8766;
assign 1_n10340 = 1_n8488 | 1_n8642;
assign 1_n5422 = ~(1_n1768 ^ 1_n6626);
assign 1_n3400 = 1_n9461 & 1_n6269;
assign 1_n4643 = ~1_n11158;
assign 1_n2123 = ~1_n6273;
assign 1_n6592 = 1_n12999 & 1_n4923;
assign 1_n49 = ~(1_n7039 ^ 1_n2105);
assign 1_n10707 = ~(1_n1085 ^ 1_n10860);
assign 1_n11702 = 1_n10281 | 1_n1026;
assign 1_n6549 = ~(1_n8373 ^ 1_n5519);
assign 1_n11321 = 1_n56 & 1_n4392;
assign 1_n12117 = 1_n11926 & 1_n8657;
assign 1_n3215 = 1_n12019 | 1_n6660;
assign 1_n8714 = ~(1_n1239 ^ 1_n4747);
assign 1_n1815 = ~1_n4039;
assign 1_n12057 = 1_n8043 | 1_n7270;
assign 1_n9202 = 1_n12348 & 1_n6937;
assign 1_n3685 = ~(1_n2530 ^ 1_n9545);
assign 1_n3561 = ~(1_n5052 | 1_n11325);
assign 1_n4524 = ~1_n9483;
assign 1_n6888 = 1_n9538 & 1_n7942;
assign 1_n12684 = 1_n3467 & 1_n5577;
assign 1_n3135 = ~(1_n6222 ^ 1_n6931);
assign 1_n12200 = ~(1_n1478 | 1_n6547);
assign 1_n453 = 1_n4252 | 1_n9554;
assign 1_n6262 = ~(1_n1611 ^ 1_n8894);
assign 1_n11491 = ~1_n3967;
assign 1_n13175 = ~(1_n10993 ^ 1_n8159);
assign 1_n7757 = ~(1_n10703 ^ 1_n1566);
assign 1_n5363 = 1_n8550 & 1_n13119;
assign 1_n8000 = ~(1_n2473 ^ 1_n910);
assign 1_n5174 = 1_n11360 & 1_n11330;
assign 1_n1903 = 1_n5645 | 1_n7935;
assign 1_n9722 = ~1_n3895;
assign 1_n1267 = 1_n4762 | 1_n4375;
assign 1_n2203 = 1_n6506 | 1_n8360;
assign 1_n2809 = ~1_n2540;
assign 1_n10570 = ~1_n3562;
assign 1_n5203 = ~(1_n10424 | 1_n13076);
assign 1_n12216 = ~(1_n7832 ^ 1_n9230);
assign 1_n8293 = ~1_n11366;
assign 1_n8455 = 1_n9606 | 1_n2544;
assign 1_n9674 = ~1_n12468;
assign 1_n582 = 1_n7500 ^ 1_n567;
assign 1_n2745 = ~(1_n5987 ^ 1_n6447);
assign 1_n6481 = ~1_n7830;
assign 1_n1270 = 1_n3244 & 1_n8457;
assign 1_n6921 = 1_n9353 & 1_n3815;
assign 1_n6432 = ~(1_n8237 ^ 1_n3638);
assign 1_n7149 = 1_n3443 | 1_n6795;
assign 1_n1716 = ~(1_n5737 ^ 1_n9262);
assign 1_n7146 = ~1_n12651;
assign 1_n5985 = ~(1_n5062 ^ 1_n6957);
assign 1_n12497 = ~(1_n3554 ^ 1_n4108);
assign 1_n10453 = ~(1_n7452 ^ 1_n4151);
assign 1_n7433 = 1_n7311 | 1_n6251;
assign 1_n4429 = ~(1_n440 ^ 1_n6827);
assign 1_n9080 = ~1_n10451;
assign 1_n7538 = 1_n2764 | 1_n7504;
assign 1_n3691 = 1_n3720 & 1_n4079;
assign 1_n8503 = ~(1_n12970 ^ 1_n995);
assign 1_n133 = 1_n6777 | 1_n10205;
assign 1_n10197 = ~(1_n4928 ^ 1_n3064);
assign 1_n8875 = 1_n1912 & 1_n11634;
assign 1_n7324 = 1_n4236 & 1_n11989;
assign 1_n11107 = 1_n917;
assign 1_n7014 = ~(1_n12704 | 1_n10267);
assign 1_n11302 = ~(1_n10438 | 1_n12849);
assign 1_n8051 = 1_n7329 | 1_n12350;
assign 1_n777 = 1_n3910 ^ 1_n9666;
assign 1_n10108 = ~1_n3310;
assign 1_n7389 = 1_n4903 & 1_n9015;
assign 1_n10095 = ~(1_n12317 ^ 1_n9902);
assign 1_n9455 = 1_n9087 & 1_n2453;
assign 1_n10762 = 1_n6988 | 1_n7430;
assign 1_n526 = ~1_n3862;
assign 1_n2645 = ~(1_n11520 ^ 1_n7370);
assign 1_n4552 = ~(1_n7494 | 1_n2815);
assign 1_n828 = 1_n4198 | 1_n7221;
assign 1_n6505 = ~(1_n6884 | 1_n6424);
assign 1_n11367 = ~(1_n5125 ^ 1_n12077);
assign 1_n3521 = ~(1_n3351 ^ 1_n1956);
assign 1_n8291 = 1_n3006 & 1_n7411;
assign 1_n4395 = 1_n73 & 1_n2634;
assign 1_n377 = 1_n5168 | 1_n9159;
assign 1_n9110 = ~(1_n6737 | 1_n4245);
assign 1_n905 = ~1_n2771;
assign 1_n10116 = 1_n8866 & 1_n8620;
assign 1_n4786 = ~1_n4020;
assign 1_n3281 = ~1_n469;
assign 1_n8304 = ~(1_n4728 | 1_n10414);
assign 1_n7475 = 1_n6349 | 1_n2408;
assign 1_n9545 = 1_n12473 ^ 1_n11149;
assign 1_n576 = ~(1_n8059 ^ 1_n10722);
assign 1_n4038 = 1_n4144 | 1_n8030;
assign 1_n11356 = ~1_n1650;
assign 1_n2692 = ~1_n7729;
assign 1_n8845 = 1_n1648 & 1_n8952;
assign 1_n2095 = ~1_n12605;
assign 1_n99 = 1_n9793 | 1_n1144;
assign 1_n9121 = ~(1_n1072 ^ 1_n10473);
assign 1_n4850 = 1_n4830 | 1_n12089;
assign 1_n9945 = 1_n938 ^ 1_n7006;
assign 1_n9507 = 1_n5164 & 1_n7412;
assign 1_n5249 = 1_n4523 | 1_n10528;
assign 1_n1043 = 1_n3858;
assign 1_n566 = 1_n9479 & 1_n8883;
assign 1_n1310 = ~(1_n12466 ^ 1_n10742);
assign 1_n9470 = 1_n11018 | 1_n10213;
assign 1_n1829 = 1_n6687 & 1_n432;
assign 1_n4342 = ~1_n11901;
assign 1_n12939 = 1_n2449 | 1_n1026;
assign 1_n5088 = 1_n10755 | 1_n12831;
assign 1_n9412 = ~(1_n1285 ^ 1_n857);
assign 1_n9167 = ~(1_n5858 ^ 1_n7206);
assign 1_n1301 = ~1_n2592;
assign 1_n11426 = 1_n3907 & 1_n10413;
assign 1_n4653 = ~1_n13160;
assign 1_n10336 = 1_n12663 | 1_n10535;
assign 1_n3034 = ~(1_n2120 ^ 1_n3808);
assign 1_n4846 = ~1_n8314;
assign 1_n1634 = ~1_n5167;
assign 1_n5908 = ~(1_n3891 ^ 1_n2833);
assign 1_n9175 = ~(1_n6603 ^ 1_n10079);
assign 1_n7448 = ~(1_n9441 ^ 1_n8368);
assign 1_n4880 = 1_n7002 & 1_n9240;
assign 1_n7899 = 1_n5025 | 1_n3893;
assign 1_n13162 = 1_n7878 | 1_n2893;
assign 1_n13218 = 1_n4232 | 1_n6692;
assign 1_n859 = ~(1_n3978 ^ 1_n8270);
assign 1_n10960 = 1_n9487 | 1_n4870;
assign 1_n10859 = ~(1_n9318 ^ 1_n10970);
assign 1_n5355 = 1_n3167 & 1_n2995;
assign 1_n8033 = ~1_n10789;
assign 1_n8441 = ~(1_n7439 ^ 1_n10963);
assign 1_n8622 = 1_n8863 | 1_n10573;
assign 1_n8617 = ~1_n9708;
assign 1_n6774 = ~1_n1418;
assign 1_n10783 = 1_n9643 | 1_n2775;
assign 1_n4886 = ~(1_n4991 ^ 1_n12980);
assign 1_n11507 = ~(1_n3151 ^ 1_n11033);
assign 1_n13187 = ~(1_n6389 ^ 1_n2869);
assign 1_n68 = 1_n10460 & 1_n5589;
assign 1_n1651 = ~1_n9300;
assign 1_n5724 = 1_n6346 & 1_n1745;
assign 1_n4345 = 1_n3315 & 1_n5760;
assign 1_n4564 = ~1_n4862;
assign 1_n4267 = 1_n4156 | 1_n10907;
assign 1_n6292 = 1_n10481 | 1_n4514;
assign 1_n6463 = ~1_n6058;
assign 1_n10158 = ~1_n3145;
assign 1_n9944 = ~(1_n1656 | 1_n5376);
assign 1_n226 = 1_n1569 & 1_n7883;
assign 1_n5640 = ~(1_n4800 ^ 1_n9103);
assign 1_n12107 = ~1_n6456;
assign 1_n3826 = ~1_n11891;
assign 1_n4745 = 1_n6890 & 1_n6584;
assign 1_n6933 = ~(1_n6864 | 1_n4977);
assign 1_n450 = ~(1_n4210 | 1_n6150);
assign 1_n2787 = ~(1_n1019 ^ 1_n12245);
assign 1_n1533 = 1_n1041 | 1_n3824;
assign 1_n11594 = ~(1_n9918 ^ 1_n11339);
assign 1_n4095 = 1_n4927 & 1_n11100;
assign 1_n6810 = ~1_n6149;
assign 1_n10812 = 1_n6223 | 1_n10029;
assign 1_n5674 = 1_n9994 & 1_n7811;
assign 1_n6972 = ~(1_n8627 | 1_n11334);
assign 1_n1109 = 1_n7486 & 1_n6159;
assign 1_n12411 = 1_n8562 | 1_n10106;
assign 1_n3166 = 1_n12759 | 1_n356;
assign 1_n3486 = 1_n8625 | 1_n9970;
assign 1_n9472 = 1_n6323 & 1_n10510;
assign 1_n4854 = 1_n4089 & 1_n9059;
assign 1_n4284 = ~(1_n9096 ^ 1_n1110);
assign 1_n3921 = ~(1_n4630 ^ 1_n4380);
assign 1_n540 = ~(1_n10019 ^ 1_n3472);
assign 1_n9250 = ~(1_n11621 ^ 1_n9175);
assign 1_n9673 = 1_n5806 | 1_n2276;
assign 1_n4593 = ~(1_n6701 | 1_n7844);
assign 1_n1179 = ~(1_n9612 ^ 1_n12677);
assign 1_n10662 = ~(1_n8888 ^ 1_n9707);
assign 1_n10264 = ~(1_n8023 ^ 1_n12363);
assign 1_n6369 = ~1_n6550;
assign 1_n247 = ~(1_n4384 | 1_n2210);
assign 1_n9636 = 1_n932 & 1_n4494;
assign 1_n571 = ~(1_n4709 ^ 1_n7781);
assign 1_n3052 = ~(1_n8087 ^ 1_n3403);
assign 1_n4015 = ~(1_n11010 ^ 1_n9046);
assign 1_n3859 = 1_n12861 | 1_n9661;
assign 1_n2194 = 1_n517 | 1_n1229;
assign 1_n9082 = ~(1_n695 ^ 1_n6411);
assign 1_n8922 = ~1_n10067;
assign 1_n11765 = ~(1_n6599 | 1_n1108);
assign 1_n13 = 1_n4077 | 1_n8348;
assign 1_n1356 = ~1_n2658;
assign 1_n8790 = ~1_n4353;
assign 1_n4661 = 1_n12995 & 1_n8433;
assign 1_n2284 = 1_n11113 | 1_n4947;
assign 1_n8638 = ~(1_n12329 ^ 1_n12);
assign 1_n7642 = ~1_n9093;
assign 1_n11042 = ~(1_n3479 ^ 1_n11084);
assign 1_n1556 = ~(1_n7329 ^ 1_n12350);
assign 1_n10488 = 1_n11333 | 1_n3676;
assign 1_n8850 = 1_n2718 | 1_n6769;
assign 1_n402 = ~(1_n4196 | 1_n2004);
assign 1_n5496 = 1_n6658 | 1_n4373;
assign 1_n2483 = ~(1_n12409 ^ 1_n743);
assign 1_n706 = ~(1_n3360 ^ 1_n2234);
assign 1_n12638 = ~(1_n11571 ^ 1_n12271);
assign 1_n4325 = 1_n1216 & 1_n8452;
assign 1_n6514 = ~(1_n1177 ^ 1_n9449);
assign 1_n6416 = ~1_n4862;
assign 1_n5856 = ~(1_n5194 ^ 1_n5623);
assign 1_n12469 = ~1_n9591;
assign 1_n5313 = ~1_n1465;
assign 1_n5930 = ~1_n9729;
assign 1_n12626 = 1_n9493 | 1_n9114;
assign 1_n9971 = ~(1_n6820 | 1_n2915);
assign 1_n458 = 1_n3906 | 1_n10250;
assign 1_n666 = ~1_n2750;
assign 1_n2589 = 1_n5719 & 1_n6057;
assign 1_n5196 = 1_n9102 & 1_n10368;
assign 1_n2721 = 1_n8723 & 1_n2151;
assign 1_n9869 = 1_n6387 | 1_n7071;
assign 1_n9435 = ~(1_n12178 ^ 1_n5295);
assign 1_n2197 = ~(1_n11971 | 1_n9068);
assign 1_n2540 = 1_n542 | 1_n206;
assign 1_n9977 = 1_n1419 | 1_n30;
assign 1_n12387 = 1_n4937 & 1_n978;
assign 1_n11678 = ~(1_n12081 | 1_n12116);
assign 1_n11519 = ~1_n12284;
assign 1_n9488 = 1_n10792 | 1_n5087;
assign 1_n2982 = 1_n3864 | 1_n7218;
assign 1_n4375 = ~(1_n7992 | 1_n6554);
assign 1_n4318 = ~(1_n2188 ^ 1_n6955);
assign 1_n6782 = ~(1_n4827 ^ 1_n916);
assign 1_n5257 = 1_n10081 | 1_n7282;
assign 1_n2526 = ~(1_n3860 ^ 1_n7352);
assign 1_n4501 = ~(1_n7018 ^ 1_n3328);
assign 1_n8220 = 1_n2088 & 1_n5851;
assign 1_n6839 = 1_n2945 & 1_n8559;
assign 1_n10910 = ~1_n3824;
assign 1_n5575 = 1_n2559 & 1_n4921;
assign 1_n2499 = 1_n1842 | 1_n6697;
assign 1_n1169 = 1_n12868 & 1_n2755;
assign 1_n1315 = 1_n12924 | 1_n492;
assign 1_n11858 = ~1_n5750;
assign 1_n1793 = ~(1_n6558 ^ 1_n9782);
assign 1_n5319 = ~(1_n12184 ^ 1_n2588);
assign 1_n2524 = ~(1_n9358 | 1_n4645);
assign 1_n5885 = 1_n5351 & 1_n12659;
assign 1_n11505 = 1_n4861 & 1_n5447;
assign 1_n10625 = 1_n10877 | 1_n8702;
assign 1_n6787 = 1_n4834 & 1_n12580;
assign 1_n7375 = 1_n4385 | 1_n6769;
assign 1_n1071 = ~(1_n4479 ^ 1_n10582);
assign 1_n2954 = ~(1_n1031 ^ 1_n1412);
assign 1_n8988 = ~(1_n8398 ^ 1_n1190);
assign 1_n9845 = ~(1_n11220 | 1_n10953);
assign 1_n5934 = ~(1_n351 ^ 1_n4833);
assign 1_n1680 = 1_n1199 | 1_n8030;
assign 1_n11758 = ~(1_n3263 ^ 1_n12045);
assign 1_n5933 = 1_n9181 | 1_n4237;
assign 1_n9207 = 1_n3814 & 1_n12504;
assign 1_n11809 = ~(1_n7383 ^ 1_n5068);
assign 1_n10376 = 1_n10908 & 1_n469;
assign 1_n8030 = 1_n5654;
assign 1_n7809 = 1_n11340 | 1_n4601;
assign 1_n1470 = ~(1_n12947 ^ 1_n43);
assign 1_n13199 = ~(1_n2950 ^ 1_n3143);
assign 1_n2800 = ~1_n11068;
assign 1_n4403 = 1_n11291 | 1_n12328;
assign 1_n12105 = 1_n7406 | 1_n11860;
assign 1_n1552 = ~(1_n7892 ^ 1_n9818);
assign 1_n7270 = ~(1_n13061 ^ 1_n3066);
assign 1_n6783 = ~1_n9822;
assign 1_n10294 = 1_n6330 & 1_n3387;
assign 1_n4674 = ~(1_n7096 | 1_n8340);
assign 1_n5861 = 1_n1756 & 1_n4773;
assign 1_n10448 = ~1_n12289;
assign 1_n5485 = ~1_n7540;
assign 1_n11155 = 1_n3616 | 1_n12328;
assign 1_n9973 = ~(1_n5606 ^ 1_n13129);
assign 1_n8722 = 1_n12677 | 1_n9612;
assign 1_n3235 = ~1_n6302;
assign 1_n8518 = 1_n12112 ^ 1_n11513;
assign 1_n1059 = 1_n11905 | 1_n3782;
assign 1_n10091 = 1_n542 | 1_n4936;
assign 1_n11820 = ~(1_n11632 | 1_n4683);
assign 1_n7217 = 1_n1038 ^ 1_n8191;
assign 1_n12599 = 1_n7742 | 1_n12188;
assign 1_n11460 = 1_n4722 | 1_n9075;
assign 1_n8194 = ~1_n6167;
assign 1_n12229 = ~(1_n11221 ^ 1_n1382);
assign 1_n13211 = ~(1_n11691 ^ 1_n11072);
assign 1_n13152 = ~(1_n8298 | 1_n1821);
assign 1_n1284 = ~(1_n8049 ^ 1_n5214);
assign 1_n8624 = ~(1_n6027 ^ 1_n4214);
assign 1_n5165 = 1_n6084 | 1_n8061;
assign 1_n114 = ~1_n10606;
assign 1_n10951 = ~(1_n3765 ^ 1_n10734);
assign 1_n11693 = ~(1_n12715 ^ 1_n3465);
assign 1_n10177 = ~(1_n3319 ^ 1_n3789);
assign 1_n8229 = 1_n11913 & 1_n3642;
assign 1_n8180 = 1_n6375 | 1_n11144;
assign 1_n1534 = ~(1_n2894 ^ 1_n806);
assign 1_n239 = 1_n2752 | 1_n7010;
assign 1_n2710 = 1_n11779 | 1_n9195;
assign 1_n12281 = ~1_n424;
assign 1_n11252 = ~(1_n3355 ^ 1_n12364);
assign 1_n10310 = 1_n1446 & 1_n11652;
assign 1_n2508 = ~(1_n7940 | 1_n2152);
assign 1_n5202 = 1_n4827 & 1_n2240;
assign 1_n2605 = ~1_n5237;
assign 1_n4610 = ~1_n7659;
assign 1_n2297 = 1_n10418 & 1_n3094;
assign 1_n9859 = ~(1_n6012 | 1_n8797);
assign 1_n7747 = 1_n2771 & 1_n9531;
assign 1_n7832 = 1_n1390 & 1_n12612;
assign 1_n112 = 1_n5976 & 1_n1372;
assign 1_n4746 = ~(1_n6495 ^ 1_n2374);
assign 1_n6066 = 1_n9658 | 1_n11809;
assign 1_n9362 = 1_n1605 | 1_n6944;
assign 1_n11373 = 1_n12728 | 1_n11209;
assign 1_n2160 = 1_n13036 | 1_n5076;
assign 1_n6203 = 1_n2135 | 1_n12881;
assign 1_n1500 = ~(1_n11907 | 1_n12327);
assign 1_n5331 = 1_n10021 | 1_n7837;
assign 1_n4226 = 1_n11476 & 1_n7398;
assign 1_n9634 = 1_n3487 & 1_n4313;
assign 1_n1812 = ~(1_n9946 ^ 1_n12731);
assign 1_n2991 = ~(1_n1063 ^ 1_n5147);
assign 1_n7057 = ~(1_n6259 ^ 1_n3461);
assign 1_n6530 = 1_n12159 | 1_n650;
assign 1_n1929 = ~(1_n6024 ^ 1_n9038);
assign 1_n3874 = ~(1_n13009 | 1_n7105);
assign 1_n10950 = ~1_n9570;
assign 1_n622 = ~1_n11618;
assign 1_n6534 = ~(1_n3469 | 1_n11958);
assign 1_n4960 = ~1_n411;
assign 1_n5478 = ~1_n12306;
assign 1_n10285 = ~1_n2629;
assign 1_n7495 = 1_n8587 & 1_n9776;
assign 1_n2190 = ~(1_n3709 ^ 1_n11769);
assign 1_n7523 = 1_n3225 | 1_n8702;
assign 1_n1318 = ~(1_n6107 ^ 1_n444);
assign 1_n4857 = 1_n2332 | 1_n4936;
assign 1_n4384 = 1_n4557 & 1_n4703;
assign 1_n7130 = ~1_n12935;
assign 1_n4780 = ~1_n1902;
assign 1_n11073 = ~(1_n414 ^ 1_n945);
assign 1_n1288 = 1_n12799 & 1_n5361;
assign 1_n10224 = ~(1_n276 ^ 1_n10454);
assign 1_n1453 = 1_n7752 | 1_n10360;
assign 1_n4776 = 1_n12993 | 1_n11274;
assign 1_n8757 = ~1_n9300;
assign 1_n2606 = ~(1_n12603 | 1_n1910);
assign 1_n12811 = ~(1_n645 | 1_n3600);
assign 1_n11198 = ~(1_n13153 | 1_n4674);
assign 1_n7176 = 1_n10135 | 1_n8030;
assign 1_n6991 = ~(1_n10842 ^ 1_n10347);
assign 1_n1407 = ~(1_n2822 ^ 1_n9658);
assign 1_n7285 = ~(1_n8091 ^ 1_n10382);
assign 1_n697 = ~(1_n6766 ^ 1_n4292);
assign 1_n5664 = 1_n12153 | 1_n7825;
assign 1_n1589 = ~1_n8290;
assign 1_n5581 = 1_n10516 & 1_n4171;
assign 1_n1611 = 1_n2591 ^ 1_n11202;
assign 1_n1446 = 1_n4964 & 1_n8506;
assign 1_n9108 = 1_n2547 & 1_n7471;
assign 1_n317 = 1_n8469 | 1_n961;
assign 1_n4563 = 1_n2681 & 1_n9344;
assign 1_n1549 = ~1_n4946;
assign 1_n6893 = 1_n13214;
assign 1_n8666 = ~1_n12282;
assign 1_n12637 = 1_n1536 | 1_n6265;
assign 1_n5953 = 1_n8761 | 1_n5769;
assign 1_n102 = 1_n12037 & 1_n10467;
assign 1_n8037 = 1_n6452 & 1_n7190;
assign 1_n11028 = 1_n8597 & 1_n1578;
assign 1_n4740 = 1_n10193 | 1_n5631;
assign 1_n11713 = ~1_n641;
assign 1_n313 = ~(1_n600 ^ 1_n11224);
assign 1_n10679 = ~(1_n2113 ^ 1_n9024);
assign 1_n2889 = ~1_n6085;
assign 1_n11601 = ~(1_n2019 | 1_n7696);
assign 1_n5204 = 1_n1099 | 1_n9120;
assign 1_n229 = ~(1_n5208 ^ 1_n180);
assign 1_n695 = 1_n2723 | 1_n12786;
assign 1_n1884 = ~(1_n5284 ^ 1_n818);
assign 1_n6235 = 1_n10128 | 1_n12501;
assign 1_n6003 = 1_n10070 & 1_n10053;
assign 1_n664 = 1_n3211 & 1_n7814;
assign 1_n4230 = 1_n482;
assign 1_n9864 = 1_n8764 & 1_n10880;
assign 1_n4486 = 1_n1697 & 1_n12932;
assign 1_n1685 = ~(1_n11636 ^ 1_n5220);
assign 1_n1674 = ~1_n11296;
assign 1_n7101 = 1_n11757 | 1_n6265;
assign 1_n5903 = ~(1_n2171 | 1_n10665);
assign 1_n8055 = ~1_n9136;
assign 1_n3996 = 1_n2283 | 1_n3762;
assign 1_n10633 = 1_n7715 & 1_n7411;
assign 1_n11888 = 1_n2660 | 1_n6317;
assign 1_n382 = ~(1_n1294 ^ 1_n11480);
assign 1_n10939 = 1_n7133 | 1_n12695;
assign 1_n1548 = 1_n10184 | 1_n3391;
assign 1_n11999 = 1_n8594 | 1_n12804;
assign 1_n8837 = ~1_n10185;
assign 1_n12839 = ~(1_n9514 ^ 1_n9688);
assign 1_n4236 = 1_n6143 | 1_n326;
assign 1_n3773 = 1_n12354 | 1_n11414;
assign 1_n6532 = 1_n9909 ^ 1_n3108;
assign 1_n5057 = 1_n437 | 1_n87;
assign 1_n7330 = ~(1_n2823 ^ 1_n11962);
assign 1_n10306 = ~(1_n5288 ^ 1_n2274);
assign 1_n9503 = ~(1_n3532 ^ 1_n10935);
assign 1_n676 = ~(1_n527 ^ 1_n3992);
assign 1_n3374 = 1_n11050 & 1_n457;
assign 1_n2951 = 1_n10497;
assign 1_n7322 = 1_n195 | 1_n8198;
assign 1_n600 = 1_n6325 & 1_n2006;
assign 1_n10069 = ~(1_n11439 ^ 1_n9667);
assign 1_n10106 = 1_n8640;
assign 1_n5625 = 1_n5328 | 1_n10871;
assign 1_n7090 = 1_n10870 & 1_n3937;
assign 1_n2971 = 1_n4732 | 1_n7221;
assign 1_n4496 = ~(1_n2613 ^ 1_n2172);
assign 1_n6001 = ~1_n6085;
assign 1_n4982 = ~(1_n4130 ^ 1_n1201);
assign 1_n5299 = 1_n2884 | 1_n10016;
assign 1_n8605 = ~(1_n9563 | 1_n12216);
assign 1_n7183 = ~(1_n12361 ^ 1_n4526);
assign 1_n3727 = ~1_n3061;
assign 1_n8872 = ~(1_n2505 ^ 1_n6340);
assign 1_n12968 = ~(1_n3488 ^ 1_n7965);
assign 1_n11679 = 1_n9392 & 1_n8464;
assign 1_n29 = ~(1_n5878 | 1_n708);
assign 1_n9899 = ~1_n10577;
assign 1_n1029 = 1_n2551 | 1_n5501;
assign 1_n13203 = 1_n11972 & 1_n11583;
assign 1_n8646 = ~1_n22;
assign 1_n4622 = ~(1_n3088 | 1_n6184);
assign 1_n11990 = 1_n3634 | 1_n8348;
assign 1_n11337 = ~(1_n2066 ^ 1_n12007);
assign 1_n1635 = ~(1_n9607 | 1_n1837);
assign 1_n1218 = ~1_n10408;
assign 1_n613 = 1_n11657 | 1_n7579;
assign 1_n13141 = ~1_n3330;
assign 1_n8810 = ~(1_n2897 ^ 1_n4379);
assign 1_n11580 = 1_n2974 | 1_n5240;
assign 1_n3341 = 1_n8760 | 1_n540;
assign 1_n959 = 1_n9010 | 1_n4947;
assign 1_n7549 = ~1_n5266;
assign 1_n12338 = ~(1_n5572 ^ 1_n9762);
assign 1_n1436 = ~1_n12289;
assign 1_n1677 = 1_n13079 | 1_n6474;
assign 1_n7341 = ~(1_n1378 ^ 1_n9021);
assign 1_n1942 = 1_n6184 & 1_n3088;
assign 1_n375 = 1_n4709 | 1_n526;
assign 1_n12527 = ~(1_n1389 ^ 1_n11942);
assign 1_n4782 = 1_n11371 | 1_n11292;
assign 1_n1784 = 1_n7932 | 1_n12998;
assign 1_n3175 = 1_n11167 | 1_n3485;
assign 1_n4528 = ~(1_n6036 ^ 1_n1641);
assign 1_n12036 = ~1_n6522;
assign 1_n6497 = ~(1_n473 | 1_n1662);
assign 1_n12007 = 1_n11803 & 1_n7886;
assign 1_n9632 = ~1_n9591;
assign 1_n3187 = 1_n4523 ^ 1_n11031;
assign 1_n7652 = 1_n8848 | 1_n8227;
assign 1_n5939 = ~1_n8230;
assign 1_n567 = ~(1_n2246 ^ 1_n3234);
assign 1_n8471 = 1_n3866 | 1_n11668;
assign 1_n2573 = 1_n4224 | 1_n9864;
assign 1_n1246 = ~1_n5180;
assign 1_n9144 = 1_n10059 | 1_n12388;
assign 1_n1928 = ~(1_n12828 | 1_n10732);
assign 1_n3725 = 1_n1135 | 1_n12164;
assign 1_n4527 = ~1_n7341;
assign 1_n12083 = ~1_n13214;
assign 1_n4222 = ~(1_n6555 | 1_n8437);
assign 1_n7783 = ~1_n2882;
assign 1_n7076 = ~1_n411;
assign 1_n10937 = 1_n5681 & 1_n5445;
assign 1_n536 = 1_n11810 | 1_n12273;
assign 1_n1387 = 1_n6587 | 1_n10179;
assign 1_n6828 = ~(1_n1136 ^ 1_n7956);
assign 1_n11341 = ~1_n6790;
assign 1_n4309 = ~(1_n6356 | 1_n6989);
assign 1_n10098 = ~1_n11441;
assign 1_n2417 = ~(1_n1793 ^ 1_n8178);
assign 1_n12583 = ~(1_n3203 ^ 1_n7054);
assign 1_n4989 = ~(1_n5808 ^ 1_n13209);
assign 1_n12195 = 1_n2866 & 1_n12825;
assign 1_n2716 = 1_n10541 & 1_n4260;
assign 1_n12688 = ~(1_n6943 | 1_n3637);
assign 1_n10517 = 1_n9946 & 1_n9004;
assign 1_n1020 = 1_n147 | 1_n10094;
assign 1_n12751 = ~(1_n7567 ^ 1_n6097);
assign 1_n3631 = ~(1_n3298 ^ 1_n1140);
assign 1_n10237 = 1_n1501 | 1_n3971;
assign 1_n5762 = ~(1_n10389 ^ 1_n1964);
assign 1_n6092 = ~(1_n11192 ^ 1_n9199);
assign 1_n4370 = ~1_n12408;
assign 1_n9462 = ~(1_n12299 | 1_n324);
assign 1_n1172 = ~(1_n8581 ^ 1_n10330);
assign 1_n4298 = 1_n4143 | 1_n12501;
assign 1_n5256 = 1_n7622 | 1_n8815;
assign 1_n10602 = ~(1_n5290 ^ 1_n5214);
assign 1_n8733 = 1_n12262 | 1_n3227;
assign 1_n1887 = ~1_n1307;
assign 1_n4785 = 1_n493 | 1_n5169;
assign 1_n725 = 1_n6649 & 1_n9770;
assign 1_n6487 = ~(1_n4046 ^ 1_n4603);
assign 1_n8478 = ~(1_n5850 | 1_n638);
assign 1_n5154 = 1_n5151 & 1_n7843;
assign 1_n2861 = ~1_n2498;
assign 1_n12958 = ~(1_n1777 ^ 1_n4029);
assign 1_n10107 = ~(1_n11314 ^ 1_n1037);
assign 1_n10865 = 1_n445 | 1_n3949;
assign 1_n2165 = ~1_n5678;
assign 1_n4340 = ~(1_n8241 | 1_n4807);
assign 1_n10201 = 1_n3110 | 1_n1462;
assign 1_n11318 = 1_n6099 | 1_n8268;
assign 1_n6173 = ~1_n10606;
assign 1_n12343 = 1_n2965 | 1_n12561;
assign 1_n5891 = ~(1_n10839 ^ 1_n3559);
assign 1_n7735 = 1_n5142 & 1_n4945;
assign 1_n7005 = ~(1_n1414 | 1_n8960);
assign 1_n7260 = 1_n3893 & 1_n5025;
assign 1_n6734 = 1_n5568 & 1_n3006;
assign 1_n12080 = 1_n10500 | 1_n11063;
assign 1_n11840 = 1_n5568 & 1_n4470;
assign 1_n10048 = ~(1_n9994 ^ 1_n9963);
assign 1_n7956 = ~(1_n6870 ^ 1_n9144);
assign 1_n1851 = ~(1_n12661 ^ 1_n1196);
assign 1_n9801 = 1_n8648 | 1_n6436;
assign 1_n5721 = ~1_n2010;
assign 1_n980 = ~1_n4377;
assign 1_n5235 = 1_n2960 & 1_n3240;
assign 1_n981 = 1_n9054 & 1_n11825;
assign 1_n7267 = ~(1_n9957 ^ 1_n11036);
assign 1_n10808 = 1_n1364 & 1_n9915;
assign 1_n4790 = 1_n6682 | 1_n7324;
assign 1_n8998 = 1_n5460 | 1_n6306;
assign 1_n2904 = ~(1_n2668 ^ 1_n5429);
assign 1_n8166 = ~1_n9611;
assign 1_n10972 = 1_n11345 | 1_n5250;
assign 1_n11741 = 1_n9216 & 1_n5962;
assign 1_n9464 = ~1_n2279;
assign 1_n1693 = 1_n4185 | 1_n13181;
assign 1_n11646 = 1_n12151 | 1_n1814;
assign 1_n4900 = ~(1_n2536 ^ 1_n4821);
assign 1_n7168 = ~(1_n7286 ^ 1_n12377);
assign 1_n10715 = ~1_n4877;
assign 1_n1931 = 1_n1159 | 1_n6429;
assign 1_n2908 = 1_n8720 | 1_n11300;
assign 1_n5230 = ~(1_n770 ^ 1_n7115);
assign 1_n10907 = ~(1_n8273 | 1_n12986);
assign 1_n57 = 1_n12042 | 1_n1836;
assign 1_n680 = ~(1_n11739 ^ 1_n4324);
assign 1_n7965 = 1_n5835 ^ 1_n11492;
assign 1_n8438 = ~1_n6669;
assign 1_n6858 = 1_n686 | 1_n11679;
assign 1_n11862 = 1_n2771 & 1_n12289;
assign 1_n6072 = ~(1_n6744 | 1_n347);
assign 1_n6962 = 1_n12882 | 1_n4373;
assign 1_n11103 = ~(1_n1626 ^ 1_n11694);
assign 1_n5820 = 1_n9835 | 1_n1378;
assign 1_n6074 = 1_n9061 | 1_n8364;
assign 1_n2064 = ~(1_n6510 | 1_n5160);
assign 1_n3743 = 1_n4102 | 1_n5002;
assign 1_n1598 = 1_n8139 & 1_n9475;
assign 1_n1106 = ~(1_n1545 ^ 1_n10438);
assign 1_n6892 = ~(1_n9494 ^ 1_n11976);
assign 1_n7436 = ~1_n11565;
assign 1_n12711 = 1_n10775 & 1_n9956;
assign 1_n10068 = ~1_n1242;
assign 1_n4463 = 1_n2712 & 1_n5640;
assign 1_n2912 = 1_n2669 | 1_n8268;
assign 1_n1365 = 1_n899 | 1_n12501;
assign 1_n2360 = ~(1_n5958 | 1_n5426);
assign 1_n9642 = 1_n3537 | 1_n12388;
assign 1_n5981 = 1_n3892 | 1_n6404;
assign 1_n8199 = ~1_n8571;
assign 1_n3339 = 1_n5749 | 1_n2133;
assign 1_n1799 = 1_n4659 | 1_n3151;
assign 1_n7083 = ~(1_n7552 ^ 1_n13020);
assign 1_n1116 = 1_n6160 & 1_n10010;
assign 1_n10963 = 1_n208 & 1_n9716;
assign 1_n11441 = 1_n5077 & 1_n12702;
assign 1_n4084 = 1_n7772 & 1_n12289;
assign 1_n9581 = ~1_n9591;
assign 1_n13116 = ~1_n11971;
assign 1_n12866 = 1_n4799 & 1_n9074;
assign 1_n10461 = 1_n8973 & 1_n2132;
assign 1_n4512 = ~(1_n7932 ^ 1_n6677);
assign 1_n11857 = 1_n3191 & 1_n3423;
assign 1_n3373 = ~1_n2464;
assign 1_n6448 = ~1_n5421;
assign 1_n4710 = 1_n7890 | 1_n2919;
assign 1_n9721 = 1_n7379 | 1_n9116;
assign 1_n5338 = 1_n820 | 1_n4832;
assign 1_n8380 = 1_n4686 | 1_n4796;
assign 1_n3660 = 1_n3784 | 1_n3981;
assign 1_n6898 = 1_n2655 & 1_n12479;
assign 1_n13106 = 1_n117 & 1_n1749;
assign 1_n12266 = 1_n5875 | 1_n12721;
assign 1_n11139 = 1_n8903 | 1_n5432;
assign 1_n7201 = ~(1_n4184 ^ 1_n11855);
assign 1_n5999 = ~1_n11061;
assign 1_n6967 = ~1_n5969;
assign 1_n12462 = 1_n11864 | 1_n12328;
assign 1_n10438 = 1_n4258 | 1_n12501;
assign 1_n4904 = 1_n5070 & 1_n5438;
assign 1_n7430 = ~1_n10408;
assign 1_n4652 = 1_n10610 & 1_n12525;
assign 1_n0 = ~1_n7720;
assign 1_n1906 = 1_n12913 | 1_n11351;
assign 1_n8242 = ~(1_n7821 ^ 1_n4767);
assign 1_n5924 = 1_n5291 & 1_n3288;
assign 1_n2291 = 1_n11605 | 1_n7288;
assign 1_n11093 = ~(1_n2314 | 1_n1042);
assign 1_n9709 = ~1_n11236;
assign 1_n1722 = 1_n5352 ^ 1_n7044;
assign 1_n11181 = ~(1_n856 ^ 1_n2560);
assign 1_n3895 = ~1_n11974;
assign 1_n5566 = 1_n12354 & 1_n11414;
assign 1_n9046 = ~(1_n9146 ^ 1_n11802);
assign 1_n1927 = 1_n5709 ^ 1_n10343;
assign 1_n12298 = 1_n8334 & 1_n11717;
assign 1_n8957 = 1_n5226 | 1_n177;
assign 1_n10405 = ~(1_n10655 ^ 1_n224);
assign 1_n3517 = 1_n4462 | 1_n6265;
assign 1_n8160 = ~1_n12592;
assign 1_n6332 = ~1_n2882;
assign 1_n1913 = ~(1_n11273 ^ 1_n3957);
assign 1_n1574 = 1_n3683 | 1_n9832;
assign 1_n10965 = 1_n3826 | 1_n4194;
assign 1_n2032 = 1_n179 & 1_n9740;
assign 1_n4768 = ~(1_n4545 | 1_n1834);
assign 1_n10924 = ~1_n11546;
assign 1_n7059 = ~(1_n7604 ^ 1_n531);
assign 1_n744 = 1_n7059 ^ 1_n8997;
assign 1_n4071 = ~(1_n12599 ^ 1_n10350);
assign 1_n7133 = ~1_n2666;
assign 1_n9770 = 1_n4874 | 1_n9419;
assign 1_n5916 = 1_n9765 | 1_n7491;
assign 1_n9066 = 1_n7872 | 1_n9075;
assign 1_n6998 = 1_n8556 | 1_n1144;
assign 1_n8411 = ~(1_n12405 ^ 1_n4951);
assign 1_n12052 = ~1_n8860;
assign 1_n2192 = 1_n12677 & 1_n9612;
assign 1_n10014 = ~1_n3100;
assign 1_n6341 = 1_n11075 | 1_n13210;
assign 1_n7325 = 1_n3430 | 1_n7557;
assign 1_n9037 = ~(1_n10980 ^ 1_n3181);
assign 1_n847 = ~(1_n4145 ^ 1_n12150);
assign 1_n7702 = 1_n1571 | 1_n5841;
assign 1_n8500 = ~1_n7065;
assign 1_n8705 = ~(1_n6334 ^ 1_n9719);
assign 1_n12551 = 1_n8407 & 1_n12321;
assign 1_n6132 = 1_n3160 & 1_n10435;
assign 1_n753 = ~(1_n11138 ^ 1_n10801);
assign 1_n6751 = ~1_n9531;
assign 1_n5260 = ~(1_n4265 ^ 1_n2715);
assign 1_n12630 = 1_n4290 | 1_n9195;
assign 1_n10550 = ~(1_n3384 | 1_n4670);
assign 1_n9544 = ~(1_n6904 ^ 1_n1875);
assign 1_n1398 = ~(1_n12669 ^ 1_n8230);
assign 1_n11984 = ~(1_n10518 ^ 1_n7943);
assign 1_n5569 = ~1_n3112;
assign 1_n1761 = 1_n3243 | 1_n8702;
assign 1_n4654 = 1_n2452 | 1_n12501;
assign 1_n12021 = ~(1_n6327 ^ 1_n10499);
assign 1_n4211 = ~(1_n11666 ^ 1_n2626);
assign 1_n7645 = 1_n9632 | 1_n11354;
assign 1_n10659 = 1_n8073 & 1_n5247;
assign 1_n1083 = ~(1_n9713 ^ 1_n12136);
assign 1_n7582 = 1_n9455 | 1_n8253;
assign 1_n10153 = ~(1_n2661 ^ 1_n8195);
assign 1_n6993 = ~(1_n5114 | 1_n10306);
assign 1_n10860 = 1_n245 & 1_n9099;
assign 1_n3575 = ~(1_n7516 ^ 1_n10779);
assign 1_n5841 = ~1_n1364;
assign 1_n12755 = ~(1_n7822 | 1_n9603);
assign 1_n10841 = 1_n614 & 1_n133;
assign 1_n10719 = 1_n6344 | 1_n2234;
assign 1_n8159 = 1_n3217 | 1_n10246;
assign 1_n7456 = 1_n8264 | 1_n10834;
assign 1_n5552 = ~(1_n12639 ^ 1_n7698);
assign 1_n11899 = ~(1_n10638 ^ 1_n606);
assign 1_n7833 = ~1_n3091;
assign 1_n537 = ~(1_n8319 ^ 1_n711);
assign 1_n3757 = ~(1_n11276 ^ 1_n4801);
assign 1_n1655 = 1_n9020 & 1_n5771;
assign 1_n10870 = 1_n11021 | 1_n6999;
assign 1_n7623 = 1_n11519 | 1_n9282;
assign 1_n3209 = ~(1_n5397 ^ 1_n10933);
assign 1_n5059 = 1_n2373 & 1_n782;
assign 1_n12634 = ~(1_n2143 ^ 1_n8527);
assign 1_n2869 = ~(1_n4338 ^ 1_n5618);
assign 1_n7116 = ~(1_n10825 ^ 1_n2052);
assign 1_n7884 = 1_n11397 & 1_n12558;
assign 1_n13005 = ~1_n2068;
assign 1_n6924 = ~1_n4002;
assign 1_n8237 = 1_n10926 | 1_n6564;
assign 1_n10327 = 1_n6220 | 1_n4144;
assign 1_n8978 = 1_n3491 | 1_n4672;
assign 1_n7640 = 1_n1817 & 1_n5904;
assign 1_n8382 = ~(1_n10269 ^ 1_n5570);
assign 1_n6807 = 1_n2219 | 1_n7052;
assign 1_n8219 = ~(1_n7572 ^ 1_n6450);
assign 1_n5703 = 1_n10713 | 1_n2994;
assign 1_n9323 = ~1_n5709;
assign 1_n6588 = 1_n6562 | 1_n2201;
assign 1_n6077 = ~(1_n12332 ^ 1_n4771);
assign 1_n8707 = 1_n51 & 1_n671;
assign 1_n872 = 1_n621 ^ 1_n9836;
assign 1_n6367 = ~1_n1724;
assign 1_n9998 = 1_n11821 & 1_n8132;
assign 1_n5813 = ~(1_n9186 ^ 1_n4081);
assign 1_n553 = ~(1_n10034 | 1_n5089);
assign 1_n3766 = ~1_n6660;
assign 1_n9345 = ~1_n6174;
assign 1_n12982 = 1_n12074 & 1_n1873;
assign 1_n8254 = ~1_n9669;
assign 1_n4604 = ~1_n10225;
assign 1_n11973 = ~1_n8967;
assign 1_n6745 = 1_n12321 | 1_n8407;
assign 1_n5733 = ~1_n5065;
assign 1_n12164 = ~1_n854;
assign 1_n11008 = ~1_n3134;
assign 1_n3359 = 1_n5316 | 1_n9290;
assign 1_n12835 = ~(1_n6441 ^ 1_n6671);
assign 1_n3780 = 1_n3962 | 1_n8490;
assign 1_n11312 = 1_n9739 | 1_n11101;
assign 1_n8784 = 1_n7690 | 1_n199;
assign 1_n7829 = 1_n8166 & 1_n5434;
assign 1_n2378 = 1_n6463 | 1_n2976;
assign 1_n10588 = 1_n5816 & 1_n136;
assign 1_n1855 = 1_n1111 | 1_n4207;
assign 1_n6190 = 1_n9166 & 1_n4284;
assign 1_n11138 = ~(1_n6088 ^ 1_n5610);
assign 1_n10312 = ~(1_n6801 ^ 1_n4476);
assign 1_n3322 = ~(1_n1527 | 1_n6961);
assign 1_n2628 = 1_n2778 & 1_n12433;
assign 1_n10280 = ~(1_n9296 | 1_n11838);
assign 1_n6687 = 1_n8658 | 1_n6891;
assign 1_n7619 = 1_n8998 & 1_n12132;
assign 1_n4026 = 1_n1623 & 1_n5001;
assign 1_n7472 = 1_n12106 & 1_n7929;
assign 1_n6128 = 1_n199 & 1_n7690;
assign 1_n1702 = ~(1_n12936 | 1_n12538);
assign 1_n7248 = ~(1_n3152 ^ 1_n6017);
assign 1_n10811 = ~(1_n7220 ^ 1_n12373);
assign 1_n13006 = 1_n11320 | 1_n5076;
assign 1_n4310 = ~(1_n9656 ^ 1_n1948);
assign 1_n4055 = ~1_n5332;
assign 1_n9171 = ~(1_n1611 | 1_n8834);
assign 1_n10573 = ~1_n11030;
assign 1_n9678 = ~(1_n1227 ^ 1_n4647);
assign 1_n4723 = ~1_n4064;
assign 1_n5812 = ~1_n2977;
assign 1_n10643 = ~(1_n3398 ^ 1_n9480);
assign 1_n3047 = ~1_n510;
assign 1_n1101 = ~1_n2758;
assign 1_n8189 = 1_n1597 & 1_n10618;
assign 1_n3577 = 1_n5070 | 1_n5438;
assign 1_n6744 = 1_n10974 | 1_n8268;
assign 1_n8451 = ~(1_n3140 ^ 1_n5398);
assign 1_n275 = ~1_n10963;
assign 1_n11934 = ~(1_n12580 ^ 1_n4669);
assign 1_n12114 = ~1_n92;
assign 1_n12973 = ~(1_n8890 ^ 1_n5955);
assign 1_n12919 = 1_n7297 & 1_n303;
assign 1_n7143 = 1_n8329 | 1_n12847;
assign 1_n11767 = ~(1_n1873 ^ 1_n3497);
assign 1_n7742 = ~1_n2252;
assign 1_n1025 = 1_n1945 & 1_n8601;
assign 1_n7064 = 1_n9238 | 1_n2059;
assign 1_n12437 = ~(1_n12815 | 1_n2874);
assign 1_n12503 = ~(1_n8218 ^ 1_n3059);
assign 1_n9629 = 1_n12680 & 1_n6636;
assign 1_n839 = 1_n8245 | 1_n12039;
assign 1_n820 = 1_n6381 | 1_n10886;
assign 1_n11768 = 1_n5863 & 1_n5436;
assign 1_n4289 = 1_n10177 | 1_n8075;
assign 1_n6054 = ~(1_n5214 | 1_n2771);
assign 1_n3350 = 1_n3313 | 1_n14;
assign 1_n2566 = 1_n13177 & 1_n3705;
assign 1_n5860 = 1_n7839 & 1_n3552;
assign 1_n6654 = 1_n11352 | 1_n2544;
assign 1_n6418 = 1_n9974 & 1_n9323;
assign 1_n1831 = 1_n5462 & 1_n11716;
assign 1_n2774 = 1_n5970 & 1_n1687;
assign 1_n5627 = ~(1_n8856 | 1_n4340);
assign 1_n9942 = ~1_n7209;
assign 1_n6551 = ~(1_n6018 ^ 1_n280);
assign 1_n2153 = 1_n359 | 1_n7905;
assign 1_n11774 = 1_n8466 & 1_n11222;
assign 1_n20 = ~(1_n37 | 1_n5224);
assign 1_n12807 = 1_n9646 | 1_n12984;
assign 1_n3885 = ~1_n8043;
assign 1_n12607 = ~(1_n2233 | 1_n1421);
assign 1_n4307 = ~(1_n2368 ^ 1_n10107);
assign 1_n12090 = 1_n121 | 1_n11609;
assign 1_n138 = ~1_n1912;
assign 1_n11308 = ~1_n7517;
assign 1_n4651 = 1_n3340 & 1_n1953;
assign 1_n11063 = 1_n12841 | 1_n9075;
assign 1_n8198 = ~(1_n9336 | 1_n4152);
assign 1_n4447 = 1_n1251 & 1_n3351;
assign 1_n1922 = 1_n1039 & 1_n10655;
assign 1_n6009 = ~(1_n5726 ^ 1_n1552);
assign 1_n10781 = ~1_n497;
assign 1_n3905 = ~(1_n12901 ^ 1_n8047);
assign 1_n1991 = ~(1_n9443 ^ 1_n4261);
assign 1_n10473 = 1_n2999 & 1_n10235;
assign 1_n2730 = ~(1_n11805 ^ 1_n1969);
assign 1_n9190 = ~(1_n7 ^ 1_n10231);
assign 1_n11640 = 1_n4808 | 1_n12847;
assign 1_n6244 = ~1_n4646;
assign 1_n9382 = ~1_n6034;
assign 1_n1578 = 1_n6383 | 1_n10179;
assign 1_n7750 = 1_n4863 | 1_n243;
assign 1_n11296 = ~(1_n8557 ^ 1_n3704);
assign 1_n8939 = ~(1_n13156 ^ 1_n11186);
assign 1_n4434 = ~(1_n4408 ^ 1_n5910);
assign 1_n2881 = ~(1_n12760 ^ 1_n5012);
assign 1_n8298 = 1_n8681 | 1_n4373;
assign 1_n6033 = ~1_n3815;
assign 1_n3317 = ~(1_n4216 ^ 1_n6668);
assign 1_n6417 = 1_n10049 | 1_n9223;
assign 1_n6528 = ~1_n11394;
assign 1_n1331 = ~1_n3409;
assign 1_n6040 = ~1_n3085;
assign 1_n2974 = ~(1_n9317 ^ 1_n2458);
assign 1_n7732 = 1_n4352 | 1_n9682;
assign 1_n10510 = 1_n7731 | 1_n4596;
assign 1_n7713 = ~(1_n3512 ^ 1_n6781);
assign 1_n7990 = 1_n4046 | 1_n11638;
assign 1_n3902 = ~(1_n6357 | 1_n2325);
assign 1_n6679 = ~(1_n10832 | 1_n13007);
assign 1_n5751 = ~(1_n5847 ^ 1_n2915);
assign 1_n5779 = 1_n435 & 1_n4776;
assign 1_n442 = ~1_n6453;
assign 1_n8246 = ~(1_n2640 | 1_n1858);
assign 1_n1197 = ~1_n854;
assign 1_n10848 = 1_n7908 | 1_n5302;
assign 1_n10619 = 1_n9649 & 1_n2096;
assign 1_n5317 = 1_n10157 & 1_n400;
assign 1_n1588 = 1_n6368 | 1_n1154;
assign 1_n12517 = 1_n2574 | 1_n11228;
assign 1_n4407 = 1_n11945 & 1_n3773;
assign 1_n6544 = 1_n12196 & 1_n2269;
assign 1_n12461 = ~(1_n10548 ^ 1_n6281);
assign 1_n1934 = 1_n11119 & 1_n9900;
assign 1_n7868 = ~1_n4335;
assign 1_n5224 = 1_n8006 | 1_n12242;
assign 1_n5008 = 1_n8379 & 1_n5273;
assign 1_n3096 = ~1_n4419;
assign 1_n9391 = ~(1_n10308 | 1_n12917);
assign 1_n3950 = ~(1_n4439 ^ 1_n10177);
assign 1_n3573 = ~(1_n2924 ^ 1_n771);
assign 1_n9648 = 1_n11868 | 1_n8030;
assign 1_n3292 = ~(1_n1911 ^ 1_n9862);
assign 1_n3189 = ~(1_n5833 | 1_n3095);
assign 1_n13124 = ~(1_n5648 ^ 1_n7420);
assign 1_n7036 = ~(1_n10895 ^ 1_n4183);
assign 1_n8386 = 1_n5990 | 1_n7723;
assign 1_n6211 = 1_n8176 | 1_n2221;
assign 1_n1257 = 1_n12533 | 1_n283;
assign 1_n10125 = ~(1_n6727 ^ 1_n5083);
assign 1_n12681 = 1_n2221 | 1_n7723;
assign 1_n2492 = 1_n3068 | 1_n7530;
assign 1_n12363 = ~(1_n8488 ^ 1_n8642);
assign 1_n9849 = 1_n11376 ^ 1_n10200;
assign 1_n3852 = 1_n10686 | 1_n1895;
assign 1_n3223 = ~(1_n12588 ^ 1_n9302);
assign 1_n1279 = ~(1_n574 | 1_n9405);
assign 1_n2702 = 1_n10936 | 1_n10028;
assign 1_n3158 = ~1_n12482;
assign 1_n1925 = 1_n8811 & 1_n7284;
assign 1_n5743 = 1_n2444 & 1_n11461;
assign 1_n1708 = ~(1_n3707 ^ 1_n1371);
assign 1_n8470 = ~1_n5535;
assign 1_n9907 = 1_n2046 & 1_n12637;
assign 1_n11314 = ~(1_n2801 ^ 1_n7993);
assign 1_n7180 = 1_n4616 & 1_n8255;
assign 1_n9706 = ~1_n11076;
assign 1_n5755 = ~(1_n12477 ^ 1_n9404);
assign 1_n10290 = ~1_n1650;
assign 1_n3270 = 1_n7062 | 1_n7221;
assign 1_n9820 = ~(1_n11120 ^ 1_n12459);
assign 1_n7597 = ~1_n3815;
assign 1_n13129 = ~(1_n4887 ^ 1_n10523);
assign 1_n4821 = 1_n3509 | 1_n7723;
assign 1_n7690 = 1_n5265 | 1_n4640;
assign 1_n5412 = 1_n8023 | 1_n11569;
assign 1_n3649 = 1_n6916 & 1_n1664;
assign 1_n5580 = ~(1_n3597 ^ 1_n12050);
assign 1_n6406 = ~(1_n9133 ^ 1_n5113);
assign 1_n11438 = 1_n4301 & 1_n344;
assign 1_n1872 = ~(1_n8291 | 1_n783);
assign 1_n11538 = 1_n5367 & 1_n8496;
assign 1_n11518 = 1_n1308 & 1_n4498;
assign 1_n6650 = ~(1_n1501 ^ 1_n6256);
assign 1_n9813 = 1_n7284 | 1_n8811;
assign 1_n8793 = 1_n7176 & 1_n8366;
assign 1_n5509 = ~(1_n5637 ^ 1_n8193);
assign 1_n7214 = 1_n2670 ^ 1_n12665;
assign 1_n3151 = 1_n1571 | 1_n1570;
assign 1_n10398 = 1_n10770 & 1_n510;
assign 1_n9064 = ~(1_n2141 | 1_n10841);
assign 1_n3807 = 1_n9810 | 1_n3805;
assign 1_n6383 = ~1_n12263;
assign 1_n12355 = 1_n12093 | 1_n12273;
assign 1_n6596 = ~1_n10522;
assign 1_n12675 = 1_n1130 & 1_n12088;
assign 1_n10774 = 1_n2880 & 1_n11154;
assign 1_n8210 = ~1_n12414;
assign 1_n5430 = ~1_n13058;
assign 1_n7799 = ~(1_n11134 ^ 1_n10687);
assign 1_n3128 = ~1_n4982;
assign 1_n3533 = 1_n3407 | 1_n177;
assign 1_n4424 = ~(1_n395 ^ 1_n9659);
assign 1_n2474 = 1_n12441 | 1_n9223;
assign 1_n4913 = ~(1_n9938 | 1_n3146);
assign 1_n11336 = 1_n3385 | 1_n2005;
assign 1_n11952 = ~(1_n8137 ^ 1_n10954);
assign 1_n7952 = ~(1_n7160 | 1_n4374);
assign 1_n8550 = 1_n5688 | 1_n5076;
assign 1_n2012 = ~(1_n11117 ^ 1_n3093);
assign 1_n8489 = ~(1_n7048 | 1_n11265);
assign 1_n860 = 1_n11069 & 1_n4158;
assign 1_n10499 = 1_n7281;
assign 1_n597 = 1_n11555 & 1_n9728;
assign 1_n1788 = ~(1_n8448 ^ 1_n12496);
assign 1_n10726 = ~1_n5871;
assign 1_n2222 = ~1_n11030;
assign 1_n7177 = ~(1_n4041 ^ 1_n7392);
assign 1_n2557 = ~1_n9353;
assign 1_n5530 = ~(1_n2460 ^ 1_n10987);
assign 1_n10181 = ~(1_n5980 ^ 1_n4238);
assign 1_n8132 = 1_n12172 | 1_n10472;
assign 1_n9401 = 1_n6906 & 1_n6186;
assign 1_n3569 = ~(1_n12582 ^ 1_n1204);
assign 1_n12104 = 1_n2790 | 1_n4546;
assign 1_n12645 = ~(1_n12276 ^ 1_n1094);
assign 1_n10188 = ~1_n8468;
assign 1_n3092 = ~1_n3087;
assign 1_n877 = 1_n6590 | 1_n5076;
assign 1_n8712 = 1_n4406 & 1_n5165;
assign 1_n7211 = 1_n6629 | 1_n11107;
assign 1_n3263 = 1_n2321 | 1_n7998;
assign 1_n2543 = ~(1_n6111 ^ 1_n8211);
assign 1_n9471 = 1_n9154 | 1_n4640;
assign 1_n12906 = ~1_n11551;
assign 1_n10834 = 1_n8849 | 1_n6635;
assign 1_n5610 = 1_n6367 | 1_n11521;
assign 1_n3356 = ~(1_n2343 | 1_n3861);
assign 1_n4794 = ~(1_n4321 ^ 1_n11749);
assign 1_n8989 = ~1_n5553;
assign 1_n491 = 1_n410 & 1_n8662;
assign 1_n1923 = 1_n110 & 1_n5946;
assign 1_n7707 = ~1_n6826;
assign 1_n12819 = 1_n4114 & 1_n2339;
assign 1_n169 = 1_n5007 | 1_n6977;
assign 1_n7352 = 1_n623 & 1_n2863;
assign 1_n5720 = 1_n12563 | 1_n4640;
assign 1_n5215 = ~1_n4146;
assign 1_n12404 = 1_n8277 & 1_n2337;
assign 1_n9506 = 1_n6318 & 1_n12057;
assign 1_n7635 = ~(1_n10053 | 1_n10070);
assign 1_n3568 = ~(1_n1560 ^ 1_n1654);
assign 1_n8846 = 1_n4114 & 1_n1916;
assign 1_n6188 = 1_n8380 | 1_n11981;
assign 1_n5246 = 1_n12697 | 1_n7640;
assign 1_n3205 = ~(1_n13206 | 1_n5473);
assign 1_n6100 = ~1_n1964;
assign 1_n1629 = ~1_n7552;
assign 1_n6237 = 1_n10327 & 1_n6711;
assign 1_n271 = 1_n2352 | 1_n4352;
assign 1_n10896 = 1_n7917 | 1_n2049;
assign 1_n8570 = 1_n5939 | 1_n9159;
assign 1_n4422 = 1_n10710 & 1_n7665;
assign 1_n10283 = ~(1_n6373 ^ 1_n3663);
assign 1_n7840 = ~(1_n10139 ^ 1_n1093);
assign 1_n3914 = 1_n11277 | 1_n71;
assign 1_n2189 = 1_n6365 | 1_n8560;
assign 1_n7632 = 1_n5826 | 1_n2831;
assign 1_n5240 = 1_n10526 & 1_n9892;
assign 1_n7067 = ~(1_n675 ^ 1_n12345);
assign 1_n10905 = ~(1_n5978 | 1_n8126);
assign 1_n5087 = ~1_n3085;
assign 1_n6081 = ~(1_n7010 ^ 1_n9663);
assign 1_n12671 = ~1_n6937;
assign 1_n2275 = ~(1_n8880 ^ 1_n7789);
assign 1_n12542 = 1_n8700 & 1_n8382;
assign 1_n936 = 1_n12330 | 1_n2731;
assign 1_n4879 = ~1_n3121;
assign 1_n6837 = 1_n5182 | 1_n3981;
assign 1_n2902 = ~1_n679;
assign 1_n12095 = ~1_n12101;
assign 1_n3371 = 1_n5752 | 1_n2177;
assign 1_n3741 = ~(1_n307 ^ 1_n2033);
assign 1_n5089 = 1_n4369 & 1_n2951;
assign 1_n364 = ~1_n6730;
assign 1_n11436 = ~(1_n11248 | 1_n8200);
assign 1_n11231 = ~1_n8788;
assign 1_n794 = 1_n5683 | 1_n3949;
assign 1_n2279 = 1_n6236 & 1_n11565;
assign 1_n2840 = ~(1_n3348 ^ 1_n1167);
assign 1_n3 = 1_n8154 & 1_n8975;
assign 1_n12642 = 1_n1358 & 1_n1766;
assign 1_n4760 = 1_n4875 | 1_n7935;
assign 1_n7145 = ~(1_n5479 ^ 1_n2648);
assign 1_n8896 = 1_n6768 | 1_n4442;
assign 1_n2423 = ~(1_n7395 ^ 1_n2131);
assign 1_n3258 = ~(1_n7267 ^ 1_n11413);
assign 1_n10549 = 1_n5692 & 1_n5834;
assign 1_n9422 = 1_n8242 & 1_n1491;
assign 1_n7220 = 1_n7636 & 1_n4562;
assign 1_n1069 = ~(1_n307 | 1_n3422);
assign 1_n12251 = ~(1_n7465 ^ 1_n12357);
assign 1_n8164 = 1_n2066 | 1_n12007;
assign 1_n6672 = ~1_n772;
assign 1_n417 = 1_n7394 | 1_n5379;
assign 1_n2063 = ~(1_n1740 | 1_n9881);
assign 1_n3121 = ~1_n4426;
assign 1_n9936 = ~(1_n6302 ^ 1_n9032);
assign 1_n5749 = ~1_n5536;
assign 1_n9672 = 1_n9513 | 1_n1400;
assign 1_n11688 = 1_n13183 | 1_n1570;
assign 1_n4616 = 1_n4537 & 1_n10408;
assign 1_n9510 = 1_n6668 & 1_n4470;
assign 1_n1421 = 1_n13178 & 1_n6576;
assign 1_n829 = ~1_n6818;
assign 1_n8571 = 1_n3962 | 1_n7935;
assign 1_n9519 = 1_n4741 | 1_n12328;
assign 1_n11627 = ~(1_n7746 ^ 1_n3856);
assign 1_n13135 = 1_n3280 & 1_n3844;
assign 1_n8555 = ~(1_n143 ^ 1_n7237);
assign 1_n12795 = ~1_n10805;
assign 1_n2211 = ~1_n6362;
assign 1_n8145 = 1_n7568 & 1_n6376;
assign 1_n9760 = 1_n8187 & 1_n3620;
assign 1_n3011 = ~(1_n1960 ^ 1_n8939);
assign 1_n7524 = 1_n4664 & 1_n2728;
assign 1_n4090 = ~(1_n3250 ^ 1_n12226);
assign 1_n1712 = ~1_n1752;
assign 1_n6857 = ~(1_n7660 ^ 1_n8709);
assign 1_n2685 = 1_n8421 & 1_n5150;
assign 1_n1988 = ~(1_n7137 ^ 1_n8096);
assign 1_n9776 = ~(1_n7809 ^ 1_n13232);
assign 1_n9966 = 1_n3433 | 1_n3649;
assign 1_n10692 = ~1_n472;
assign 1_n9521 = ~(1_n11448 | 1_n3082);
assign 1_n1233 = ~(1_n2600 ^ 1_n5000);
assign 1_n12610 = 1_n10792 | 1_n2449;
assign 1_n1394 = 1_n7223 | 1_n9223;
assign 1_n9112 = ~1_n5065;
assign 1_n4767 = ~(1_n5039 ^ 1_n1678);
assign 1_n19 = ~1_n11151;
assign 1_n598 = 1_n896 & 1_n11620;
assign 1_n10807 = 1_n12814 | 1_n5242;
assign 1_n6952 = 1_n2199 & 1_n2385;
assign 1_n6319 = ~(1_n6972 | 1_n12694);
assign 1_n2945 = ~1_n1623;
assign 1_n10126 = ~(1_n9134 ^ 1_n2035);
assign 1_n5042 = ~(1_n7489 ^ 1_n10836);
assign 1_n9925 = ~(1_n220 ^ 1_n2548);
assign 1_n10736 = ~(1_n7885 ^ 1_n1010);
assign 1_n201 = ~(1_n8304 ^ 1_n7347);
assign 1_n9917 = ~1_n4743;
assign 1_n5780 = ~(1_n11318 ^ 1_n2275);
assign 1_n10596 = ~(1_n3590 ^ 1_n9256);
assign 1_n898 = 1_n12126 | 1_n1144;
assign 1_n8526 = 1_n11994 | 1_n331;
assign 1_n989 = ~(1_n2521 | 1_n6792);
assign 1_n12242 = ~1_n1364;
assign 1_n7333 = 1_n6677 | 1_n12714;
assign 1_n11458 = ~(1_n4428 ^ 1_n3446);
assign 1_n552 = 1_n11500 & 1_n710;
assign 1_n6986 = ~1_n4862;
assign 1_n98 = ~1_n11634;
assign 1_n11525 = ~1_n9540;
assign 1_n10378 = ~(1_n6805 ^ 1_n5386);
assign 1_n12049 = ~1_n834;
assign 1_n4877 = ~1_n12083;
assign 1_n4285 = 1_n10914 ^ 1_n5960;
assign 1_n4944 = ~(1_n11546 | 1_n7199);
assign 1_n10788 = ~(1_n7382 | 1_n10461);
assign 1_n8679 = ~1_n1915;
assign 1_n412 = 1_n10291 & 1_n11439;
assign 1_n6957 = 1_n7069 ^ 1_n5124;
assign 1_n10320 = 1_n2452 | 1_n11522;
assign 1_n3421 = ~(1_n348 | 1_n4219);
assign 1_n7002 = ~(1_n3090 ^ 1_n13095);
assign 1_n5838 = ~1_n1935;
assign 1_n2422 = ~(1_n1510 ^ 1_n11298);
assign 1_n655 = 1_n3736 & 1_n929;
assign 1_n10233 = 1_n7789 | 1_n4492;
assign 1_n1103 = 1_n12353 & 1_n8316;
assign 1_n9791 = 1_n8648 & 1_n6436;
assign 1_n609 = 1_n3067 | 1_n10985;
assign 1_n4970 = 1_n7242 | 1_n12886;
assign 1_n12549 = ~(1_n3030 ^ 1_n9878);
assign 1_n10262 = 1_n10112 | 1_n5521;
assign 1_n7916 = 1_n9675 | 1_n1570;
assign 1_n10649 = ~(1_n2784 ^ 1_n1838);
assign 1_n8190 = ~(1_n4244 ^ 1_n6547);
assign 1_n5092 = 1_n10277 & 1_n3297;
assign 1_n6249 = ~(1_n7732 ^ 1_n6035);
assign 1_n7926 = ~(1_n11447 ^ 1_n12277);
assign 1_n8053 = ~1_n353;
assign 1_n10714 = ~1_n8468;
assign 1_n6815 = 1_n5502 ^ 1_n11319;
assign 1_n5772 = 1_n7260 | 1_n523;
assign 1_n8964 = ~(1_n8654 | 1_n8951);
assign 1_n7716 = ~1_n11016;
assign 1_n9633 = ~(1_n6598 ^ 1_n12439);
assign 1_n4547 = 1_n565 | 1_n8593;
assign 1_n2801 = 1_n3364 | 1_n6033;
assign 1_n8011 = ~1_n8135;
assign 1_n2270 = 1_n3880 | 1_n8953;
assign 1_n13074 = 1_n13021 & 1_n6232;
assign 1_n9410 = ~(1_n10487 ^ 1_n3904);
assign 1_n6626 = 1_n8415 | 1_n11959;
assign 1_n6049 = 1_n399 & 1_n2596;
assign 1_n643 = ~(1_n12806 ^ 1_n2589);
assign 1_n5961 = ~(1_n7043 ^ 1_n8136);
assign 1_n3926 = 1_n2302 & 1_n844;
assign 1_n13167 = ~1_n13217;
assign 1_n9308 = ~1_n2466;
assign 1_n2301 = 1_n11683 | 1_n3981;
assign 1_n4085 = 1_n1659 | 1_n10574;
assign 1_n7385 = ~(1_n12315 | 1_n6495);
assign 1_n12481 = ~(1_n4592 ^ 1_n5889);
assign 1_n2896 = ~(1_n11455 ^ 1_n11839);
assign 1_n9178 = 1_n3833 & 1_n2946;
assign 1_n1834 = ~(1_n10020 | 1_n12884);
assign 1_n7396 = ~1_n3769;
assign 1_n4968 = ~(1_n7155 ^ 1_n9825);
assign 1_n3881 = ~(1_n9670 ^ 1_n7902);
assign 1_n6357 = ~(1_n12358 ^ 1_n9412);
assign 1_n5593 = 1_n3006 & 1_n12289;
assign 1_n11539 = 1_n2485 | 1_n6032;
assign 1_n8060 = 1_n7291 | 1_n8030;
assign 1_n7444 = 1_n9161 | 1_n6372;
assign 1_n11118 = ~(1_n6569 | 1_n7169);
assign 1_n10826 = ~(1_n4298 ^ 1_n8262);
assign 1_n4451 = 1_n2825 | 1_n12388;
assign 1_n754 = 1_n3606 ^ 1_n12632;
assign 1_n232 = ~(1_n10284 ^ 1_n12513);
assign 1_n11217 = 1_n1731 ^ 1_n4443;
assign 1_n1325 = ~1_n11061;
assign 1_n11461 = 1_n10017 | 1_n8490;
assign 1_n1037 = ~(1_n4351 ^ 1_n3482);
assign 1_n2858 = ~1_n11937;
assign 1_n5876 = ~(1_n6765 ^ 1_n2572);
assign 1_n10259 = ~(1_n5637 | 1_n8193);
assign 1_n9534 = ~(1_n8762 ^ 1_n1397);
assign 1_n8299 = ~(1_n11211 ^ 1_n5422);
assign 1_n383 = 1_n7074 | 1_n9223;
assign 1_n5919 = ~(1_n11953 | 1_n578);
assign 1_n3961 = 1_n207 & 1_n12290;
assign 1_n3535 = ~(1_n12996 ^ 1_n6514);
assign 1_n7904 = ~(1_n8643 | 1_n7954);
assign 1_n7218 = ~(1_n2112 | 1_n5614);
assign 1_n75 = ~1_n13060;
assign 1_n7705 = ~(1_n4397 | 1_n8165);
assign 1_n12072 = 1_n10500 & 1_n11063;
assign 1_n1664 = 1_n1578 | 1_n8597;
assign 1_n5239 = ~(1_n12191 | 1_n12700);
assign 1_n12523 = ~(1_n8714 ^ 1_n7677);
assign 1_n2254 = ~1_n8860;
assign 1_n7786 = ~(1_n5120 | 1_n8474);
assign 1_n11455 = 1_n10037 | 1_n8534;
assign 1_n7428 = ~(1_n4931 ^ 1_n9577);
assign 1_n6869 = ~(1_n7362 | 1_n12609);
assign 1_n460 = ~(1_n4273 ^ 1_n7985);
assign 1_n1261 = ~1_n2882;
assign 1_n12803 = ~(1_n4275 ^ 1_n76);
assign 1_n8202 = 1_n3101 | 1_n1789;
assign 1_n10047 = ~(1_n9108 ^ 1_n7036);
assign 1_n10856 = ~1_n4586;
assign 1_n9751 = 1_n3911 | 1_n4947;
assign 1_n3297 = 1_n3517 | 1_n3571;
assign 1_n10169 = ~(1_n4314 ^ 1_n5004);
assign 1_n6639 = 1_n6275 & 1_n9993;
assign 1_n10863 = ~(1_n12137 ^ 1_n3213);
assign 1_n4136 = ~1_n7307;
assign 1_n7725 = ~(1_n10025 ^ 1_n12079);
assign 1_n13238 = ~1_n10770;
assign 1_n6255 = ~1_n8218;
assign 1_n7122 = 1_n5261 | 1_n3981;
assign 1_n9430 = ~1_n5815;
assign 1_n12565 = 1_n7435 & 1_n12294;
assign 1_n4909 = ~(1_n10864 ^ 1_n1757);
assign 1_n9298 = 1_n4352 | 1_n4947;
assign 1_n12722 = 1_n2150 | 1_n3177;
assign 1_n5658 = ~1_n6791;
assign 1_n6175 = ~1_n6780;
assign 1_n12450 = 1_n3469 & 1_n11958;
assign 1_n7662 = 1_n9920 | 1_n8423;
assign 1_n12136 = 1_n543 | 1_n6982;
assign 1_n5415 = 1_n8549 & 1_n8919;
assign 1_n12123 = ~(1_n6832 ^ 1_n13124);
assign 1_n4599 = 1_n2080 | 1_n2463;
assign 1_n1122 = ~(1_n8518 ^ 1_n6081);
assign 1_n10102 = 1_n7980 & 1_n3846;
assign 1_n3386 = ~(1_n5403 | 1_n11387);
assign 1_n5513 = 1_n13089 | 1_n6207;
assign 1_n3742 = ~(1_n884 ^ 1_n11251);
assign 1_n10234 = ~1_n10409;
assign 1_n6727 = 1_n3830 & 1_n4098;
assign 1_n6472 = 1_n3018 | 1_n6951;
assign 1_n3253 = ~1_n6222;
assign 1_n1202 = 1_n7358 | 1_n6769;
assign 1_n10936 = 1_n87 & 1_n437;
assign 1_n3755 = ~1_n6643;
assign 1_n7789 = 1_n6028 | 1_n7221;
assign 1_n7882 = ~(1_n11501 ^ 1_n8611);
assign 1_n8366 = 1_n11466 | 1_n4640;
assign 1_n12683 = 1_n11511 & 1_n9621;
assign 1_n12451 = ~(1_n2333 ^ 1_n11830);
assign 1_n12643 = 1_n2382 | 1_n3546;
assign 1_n2639 = ~1_n5189;
assign 1_n11686 = ~(1_n3931 | 1_n5119);
assign 1_n11166 = 1_n1735 & 1_n10674;
assign 1_n1300 = ~1_n1075;
assign 1_n7391 = 1_n5452 | 1_n12681;
assign 1_n10818 = 1_n34 & 1_n701;
assign 1_n6733 = ~1_n5189;
assign 1_n6271 = ~1_n9591;
assign 1_n1456 = ~(1_n6454 ^ 1_n2895);
assign 1_n5127 = ~(1_n4027 ^ 1_n10952);
assign 1_n1047 = ~1_n3605;
assign 1_n7225 = 1_n6433 & 1_n6276;
assign 1_n1184 = ~1_n7387;
assign 1_n1040 = 1_n8838 | 1_n6078;
assign 1_n1565 = ~(1_n12801 | 1_n9604);
assign 1_n113 = ~(1_n5734 ^ 1_n6886);
assign 1_n7255 = 1_n1653 & 1_n6479;
assign 1_n4182 = ~(1_n8245 ^ 1_n3632);
assign 1_n3228 = ~(1_n11268 ^ 1_n298);
assign 1_n2184 = ~(1_n4599 ^ 1_n9361);
assign 1_n4531 = 1_n7188 | 1_n8534;
assign 1_n9415 = 1_n1105 & 1_n3136;
assign 1_n4293 = ~1_n12391;
assign 1_n11358 = ~(1_n10261 ^ 1_n8820);
assign 1_n6675 = 1_n6725 & 1_n10862;
assign 1_n9767 = ~1_n9093;
assign 1_n9051 = 1_n8200 | 1_n2216;
assign 1_n3361 = 1_n13077 | 1_n3454;
assign 1_n2632 = ~(1_n7731 ^ 1_n4596);
assign 1_n5783 = 1_n882 | 1_n8655;
assign 1_n3335 = 1_n11061 & 1_n3769;
assign 1_n11344 = ~1_n3398;
assign 1_n288 = ~(1_n4941 | 1_n12229);
assign 1_n736 = ~(1_n274 ^ 1_n7318);
assign 1_n4873 = 1_n3060 & 1_n7046;
assign 1_n1501 = 1_n3047 | 1_n11354;
assign 1_n12521 = 1_n1933 | 1_n9407;
assign 1_n1540 = ~1_n5897;
assign 1_n642 = ~(1_n11904 ^ 1_n6788);
assign 1_n2193 = 1_n1725 | 1_n6769;
assign 1_n6495 = ~(1_n10036 ^ 1_n3072);
assign 1_n4715 = ~1_n11837;
assign 1_n2786 = 1_n6178 | 1_n5048;
assign 1_n11099 = ~1_n8476;
assign 1_n2860 = 1_n11618 | 1_n4136;
assign 1_n4493 = 1_n6336 | 1_n8752;
assign 1_n4611 = 1_n10287 | 1_n12695;
assign 1_n974 = 1_n1786 & 1_n254;
assign 1_n4373 = 1_n12537;
assign 1_n10081 = 1_n10229 | 1_n6288;
assign 1_n9377 = ~(1_n3227 ^ 1_n12262);
assign 1_n4129 = 1_n6168 & 1_n5729;
assign 1_n8749 = 1_n2768 | 1_n8268;
assign 1_n6303 = 1_n8301 | 1_n6166;
assign 1_n7088 = ~(1_n12294 ^ 1_n5067);
assign 1_n9557 = ~1_n1724;
assign 1_n10037 = ~1_n8233;
assign 1_n10136 = 1_n12841 | 1_n121;
assign 1_n874 = ~(1_n8703 ^ 1_n4965);
assign 1_n7278 = 1_n7775 | 1_n11483;
assign 1_n6632 = 1_n203 & 1_n4218;
assign 1_n3595 = 1_n1326 | 1_n5476;
assign 1_n1768 = ~(1_n4555 | 1_n2450);
assign 1_n11798 = 1_n5533 & 1_n5621;
assign 1_n2253 = 1_n475 | 1_n12942;
assign 1_n6492 = 1_n6439 | 1_n6306;
assign 1_n7479 = 1_n12445 & 1_n1681;
assign 1_n8824 = 1_n3852 & 1_n10363;
assign 1_n9454 = 1_n3360 | 1_n10511;
assign 1_n11522 = ~1_n8230;
assign 1_n4992 = ~(1_n8211 | 1_n6111);
assign 1_n5342 = 1_n5947 | 1_n7723;
assign 1_n12509 = ~(1_n6540 ^ 1_n10603);
assign 1_n2765 = ~(1_n5937 ^ 1_n643);
assign 1_n2429 = ~(1_n5283 | 1_n2554);
assign 1_n8303 = ~(1_n13027 ^ 1_n3653);
assign 1_n5444 = ~(1_n9886 ^ 1_n2218);
assign 1_n7165 = ~(1_n6718 ^ 1_n2847);
assign 1_n10083 = 1_n4753 & 1_n8570;
assign 1_n4811 = 1_n2516 | 1_n9155;
assign 1_n554 = 1_n11142 | 1_n3792;
assign 1_n223 = ~(1_n9743 ^ 1_n7946);
assign 1_n2367 = 1_n6776 & 1_n12708;
assign 1_n7387 = ~(1_n592 ^ 1_n4845);
assign 1_n4813 = 1_n5909 & 1_n12792;
assign 1_n11475 = 1_n12300 & 1_n10972;
assign 1_n11797 = 1_n1256 | 1_n6285;
assign 1_n2810 = 1_n8485 & 1_n12078;
assign 1_n9571 = 1_n7333 & 1_n1784;
assign 1_n8070 = 1_n9215 & 1_n10927;
assign 1_n13222 = ~(1_n2524 | 1_n3691);
assign 1_n6896 = ~(1_n9594 ^ 1_n3621);
assign 1_n620 = 1_n11580 & 1_n9937;
assign 1_n843 = ~(1_n11100 ^ 1_n4927);
assign 1_n10123 = 1_n12545 | 1_n5924;
assign 1_n5827 = ~1_n8200;
assign 1_n10049 = ~1_n5962;
assign 1_n10773 = ~(1_n5322 ^ 1_n7172);
assign 1_n8593 = 1_n10172 ^ 1_n9137;
assign 1_n7337 = 1_n1389 | 1_n3014;
assign 1_n9832 = 1_n3851 & 1_n12382;
assign 1_n8404 = ~(1_n7402 ^ 1_n2331);
assign 1_n11523 = ~(1_n10739 | 1_n5824);
assign 1_n5318 = 1_n7828 | 1_n3888;
assign 1_n7490 = ~(1_n3855 | 1_n1046);
assign 1_n419 = ~(1_n5678 | 1_n8684);
assign 1_n9379 = 1_n9656 & 1_n10848;
assign 1_n4406 = 1_n4663 | 1_n1127;
assign 1_n9911 = 1_n12732 | 1_n10319;
assign 1_n4550 = ~(1_n664 | 1_n5759);
assign 1_n4732 = ~1_n2737;
assign 1_n2819 = ~(1_n7989 ^ 1_n977);
assign 1_n917 = ~1_n3006;
assign 1_n5442 = ~(1_n972 ^ 1_n11071);
assign 1_n6014 = ~(1_n345 ^ 1_n8054);
assign 1_n10352 = ~1_n2758;
assign 1_n12318 = 1_n920 | 1_n9079;
assign 1_n5835 = ~(1_n1645 ^ 1_n6169);
assign 1_n13031 = ~(1_n4832 ^ 1_n2586);
assign 1_n12447 = ~(1_n6338 | 1_n5739);
assign 1_n10869 = ~(1_n2931 ^ 1_n1980);
assign 1_n4207 = ~(1_n12735 | 1_n11432);
assign 1_n4597 = ~(1_n4793 ^ 1_n11622);
assign 1_n5557 = ~(1_n9920 ^ 1_n9991);
assign 1_n7417 = ~(1_n10824 ^ 1_n8147);
assign 1_n4287 = ~(1_n288 | 1_n2628);
assign 1_n3840 = 1_n12222 & 1_n4336;
assign 1_n5182 = ~1_n12965;
assign 1_n2133 = 1_n1301;
assign 1_n5259 = ~(1_n5906 ^ 1_n1100);
assign 1_n1042 = ~(1_n5731 | 1_n11108);
assign 1_n635 = 1_n6069 | 1_n11067;
assign 1_n4972 = ~(1_n13131 ^ 1_n7108);
assign 1_n2714 = 1_n9690 & 1_n10741;
assign 1_n4911 = ~(1_n11269 ^ 1_n8196);
assign 1_n5426 = ~(1_n2935 | 1_n31);
assign 1_n1849 = 1_n12107 & 1_n8907;
assign 1_n5161 = ~(1_n6396 ^ 1_n7425);
assign 1_n11607 = ~(1_n9079 ^ 1_n10934);
assign 1_n10247 = ~(1_n11090 ^ 1_n468);
assign 1_n4046 = ~(1_n1747 ^ 1_n11145);
assign 1_n1219 = 1_n9115 & 1_n6538;
assign 1_n10684 = ~(1_n2785 ^ 1_n1895);
assign 1_n12186 = 1_n5707 & 1_n1432;
assign 1_n2967 = ~1_n3954;
assign 1_n5788 = ~(1_n5216 | 1_n3751);
assign 1_n78 = 1_n951 & 1_n3085;
assign 1_n4444 = ~(1_n3740 ^ 1_n9599);
assign 1_n9478 = ~1_n9747;
assign 1_n116 = ~1_n13221;
assign 1_n12844 = 1_n8351 | 1_n6532;
assign 1_n9143 = ~(1_n11901 ^ 1_n10809);
assign 1_n12271 = 1_n8020 | 1_n206;
assign 1_n10424 = ~(1_n1098 ^ 1_n9766);
assign 1_n3174 = 1_n5040 | 1_n11144;
assign 1_n1023 = 1_n8472 | 1_n3981;
assign 1_n3247 = 1_n12837 | 1_n1325;
assign 1_n5166 = 1_n3770 | 1_n3084;
assign 1_n8272 = 1_n2135 | 1_n894;
assign 1_n2653 = ~(1_n9994 | 1_n7811);
assign 1_n4842 = ~(1_n12971 ^ 1_n3470);
assign 1_n12989 = 1_n8176 | 1_n11122;
assign 1_n6136 = 1_n1077 | 1_n3960;
assign 1_n5145 = 1_n10031 | 1_n4226;
assign 1_n4332 = 1_n9228 | 1_n3817;
assign 1_n8751 = 1_n3105 | 1_n6746;
assign 1_n9783 = 1_n6685 | 1_n1458;
assign 1_n11047 = 1_n2299 & 1_n12190;
assign 1_n762 = ~(1_n12943 ^ 1_n2839);
assign 1_n8414 = 1_n3175 & 1_n8731;
assign 1_n862 = ~(1_n1951 ^ 1_n12739);
assign 1_n2752 = ~1_n1055;
assign 1_n709 = ~1_n4036;
assign 1_n5506 = 1_n12451 | 1_n2402;
assign 1_n5294 = ~1_n1502;
assign 1_n9797 = 1_n406 | 1_n11950;
assign 1_n7788 = ~(1_n10585 ^ 1_n2696);
assign 1_n6410 = ~(1_n1559 ^ 1_n6919);
assign 1_n1825 = 1_n6051 & 1_n11998;
assign 1_n11637 = ~1_n3521;
assign 1_n10677 = 1_n12056 & 1_n2975;
assign 1_n8512 = 1_n10085 | 1_n7530;
assign 1_n12970 = ~(1_n471 ^ 1_n9472);
assign 1_n2110 = ~(1_n10064 | 1_n760);
assign 1_n5011 = 1_n8712 & 1_n11092;
assign 1_n2262 = ~(1_n11183 ^ 1_n10791);
assign 1_n9476 = 1_n7445 & 1_n216;
assign 1_n3200 = ~(1_n9505 ^ 1_n10596);
assign 1_n2037 = ~1_n3244;
assign 1_n8284 = ~(1_n8812 ^ 1_n9532);
assign 1_n8261 = 1_n197 & 1_n8785;
assign 1_n7749 = ~1_n9347;
assign 1_n3825 = ~1_n510;
assign 1_n4073 = 1_n6348 & 1_n6936;
assign 1_n10466 = ~1_n10390;
assign 1_n2376 = ~(1_n7556 ^ 1_n12291);
assign 1_n7099 = 1_n6279 & 1_n4634;
assign 1_n12801 = ~(1_n2925 | 1_n4583);
assign 1_n1396 = 1_n5888 | 1_n6572;
assign 1_n2419 = 1_n9216 & 1_n411;
assign 1_n11513 = 1_n5568 & 1_n12853;
assign 1_n8670 = 1_n3969 & 1_n10945;
assign 1_n10758 = ~(1_n9234 ^ 1_n10637);
assign 1_n11422 = 1_n12635 & 1_n9922;
assign 1_n9789 = 1_n8598 | 1_n1985;
assign 1_n10276 = 1_n9265 & 1_n9286;
assign 1_n4425 = ~(1_n10498 ^ 1_n5515);
assign 1_n10176 = ~(1_n2027 ^ 1_n6728);
assign 1_n6637 = 1_n449 | 1_n10302;
assign 1_n7768 = 1_n3478 & 1_n5537;
assign 1_n4491 = 1_n11037 | 1_n9223;
assign 1_n2438 = ~(1_n10709 ^ 1_n4413);
assign 1_n12994 = ~1_n5642;
assign 1_n5761 = ~(1_n7881 ^ 1_n11477);
assign 1_n4176 = 1_n6778 | 1_n12110;
assign 1_n12249 = ~1_n11180;
assign 1_n10003 = ~(1_n12216 ^ 1_n9563);
assign 1_n8365 = ~(1_n1359 ^ 1_n2438);
assign 1_n12640 = 1_n11707 & 1_n6358;
assign 1_n11108 = 1_n12396 | 1_n6978;
assign 1_n207 = 1_n1345 | 1_n10029;
assign 1_n11190 = ~(1_n6417 ^ 1_n8399);
assign 1_n12022 = 1_n3127 | 1_n8563;
assign 1_n9991 = ~(1_n235 ^ 1_n4816);
assign 1_n9808 = ~1_n11537;
assign 1_n8812 = 1_n5688 | 1_n8030;
assign 1_n6907 = 1_n7918 & 1_n1470;
assign 1_n7205 = ~(1_n4139 ^ 1_n6698);
assign 1_n910 = 1_n12683 | 1_n10617;
assign 1_n6073 = ~(1_n1774 ^ 1_n83);
assign 1_n9231 = 1_n8167 & 1_n3341;
assign 1_n12931 = ~(1_n13200 | 1_n6779);
assign 1_n1648 = 1_n1023 | 1_n5202;
assign 1_n264 = ~(1_n8593 ^ 1_n8921);
assign 1_n1498 = ~(1_n7000 ^ 1_n4394);
assign 1_n12264 = 1_n2768 | 1_n4230;
assign 1_n179 = ~(1_n2010 ^ 1_n7685);
assign 1_n9030 = ~(1_n5612 | 1_n5413);
assign 1_n10481 = ~1_n1636;
assign 1_n1675 = 1_n10509 | 1_n4844;
assign 1_n3640 = ~1_n5536;
assign 1_n10229 = ~1_n9948;
assign 1_n2555 = 1_n7171 & 1_n11684;
assign 1_n12736 = ~(1_n3244 ^ 1_n7107);
assign 1_n4462 = ~1_n9915;
assign 1_n4014 = ~(1_n8473 ^ 1_n3410);
assign 1_n590 = ~(1_n3115 ^ 1_n6185);
assign 1_n10204 = ~1_n1327;
assign 1_n3978 = 1_n13025 | 1_n3981;
assign 1_n7543 = 1_n4621 | 1_n121;
assign 1_n4304 = ~(1_n10183 ^ 1_n11931);
assign 1_n2575 = 1_n5922 & 1_n7874;
assign 1_n2946 = 1_n1957 | 1_n5408;
assign 1_n11610 = 1_n12417 ^ 1_n10376;
assign 1_n8389 = 1_n5086 | 1_n4515;
assign 1_n3684 = 1_n8106 | 1_n5317;
assign 1_n4865 = 1_n10619 & 1_n300;
assign 1_n10062 = ~(1_n85 ^ 1_n2857);
assign 1_n551 = 1_n6571 & 1_n11124;
assign 1_n6051 = 1_n3225 | 1_n7935;
assign 1_n5026 = ~(1_n8620 ^ 1_n8866);
assign 1_n1483 = 1_n8325 | 1_n1043;
assign 1_n10919 = 1_n2614 | 1_n1463;
assign 1_n5630 = ~1_n8394;
assign 1_n11328 = ~1_n7040;
assign 1_n12016 = 1_n11754 & 1_n8426;
assign 1_n12738 = ~1_n9367;
assign 1_n7845 = 1_n12174 | 1_n1043;
assign 1_n3180 = ~(1_n4797 ^ 1_n9311);
assign 1_n9169 = 1_n2128 | 1_n12910;
assign 1_n3062 = ~1_n12352;
assign 1_n10544 = 1_n8941 | 1_n10016;
assign 1_n9843 = ~(1_n1232 ^ 1_n10946);
assign 1_n10665 = ~(1_n1984 | 1_n8963);
assign 1_n1328 = 1_n5190 | 1_n12787;
assign 1_n13220 = ~(1_n8579 ^ 1_n4008);
assign 1_n6055 = ~1_n3286;
assign 1_n995 = ~(1_n4302 ^ 1_n2539);
assign 1_n4280 = ~(1_n5417 ^ 1_n4541);
assign 1_n10704 = 1_n2217 | 1_n479;
assign 1_n10064 = 1_n12153 | 1_n776;
assign 1_n4379 = 1_n7672 | 1_n4373;
assign 1_n3203 = 1_n2145 & 1_n7006;
assign 1_n7997 = ~(1_n622 | 1_n7307);
assign 1_n2779 = ~(1_n1316 ^ 1_n8395);
assign 1_n2200 = ~(1_n6298 ^ 1_n12529);
assign 1_n904 = ~(1_n9539 ^ 1_n5625);
assign 1_n4766 = 1_n10664 | 1_n8519;
assign 1_n7688 = 1_n9281 | 1_n6623;
assign 1_n965 = 1_n8498 | 1_n8268;
assign 1_n3758 = ~(1_n7896 | 1_n851);
assign 1_n1408 = ~(1_n12131 ^ 1_n12223);
assign 1_n6538 = ~1_n12452;
assign 1_n4532 = 1_n3311 & 1_n10408;
assign 1_n7893 = ~(1_n7542 | 1_n4534);
assign 1_n12097 = 1_n1191 | 1_n1463;
assign 1_n11618 = ~(1_n2021 ^ 1_n12937);
assign 1_n2011 = 1_n9282 | 1_n7158;
assign 1_n7126 = 1_n6250 | 1_n9159;
assign 1_n12493 = ~1_n11574;
assign 1_n5394 = ~(1_n6211 ^ 1_n8388);
assign 1_n6932 = ~(1_n7284 ^ 1_n4407);
assign 1_n4472 = 1_n250 & 1_n2492;
assign 1_n12576 = ~1_n5600;
assign 1_n6234 = 1_n10092 & 1_n3368;
assign 1_n4726 = ~(1_n2344 ^ 1_n4956);
assign 1_n4912 = 1_n2254 | 1_n237;
assign 1_n2530 = 1_n6074 & 1_n11191;
assign 1_n7962 = ~1_n9514;
assign 1_n10543 = ~(1_n348 ^ 1_n4177);
assign 1_n11533 = 1_n1634 | 1_n12621;
assign 1_n5948 = 1_n2786 | 1_n8972;
assign 1_n69 = ~1_n772;
assign 1_n2024 = 1_n3854 | 1_n6404;
assign 1_n5822 = 1_n7319 | 1_n12764;
assign 1_n10734 = 1_n5840 & 1_n101;
assign 1_n5932 = 1_n6439 | 1_n12273;
assign 1_n3779 = 1_n11650 & 1_n1121;
assign 1_n6315 = 1_n5927 | 1_n10292;
assign 1_n7964 = ~(1_n6777 ^ 1_n10205);
assign 1_n7692 = 1_n9995 & 1_n7598;
assign 1_n10590 = ~1_n6782;
assign 1_n7427 = 1_n6182 | 1_n9223;
assign 1_n3420 = 1_n2726 | 1_n3949;
assign 1_n5598 = ~(1_n2706 ^ 1_n687);
assign 1_n3898 = ~1_n11180;
assign 1_n2411 = ~1_n12156;
assign 1_n9514 = 1_n11197 & 1_n1078;
assign 1_n9796 = ~(1_n9930 ^ 1_n2565);
assign 1_n10141 = 1_n2563 | 1_n1509;
assign 1_n10751 = ~(1_n4948 ^ 1_n268);
assign 1_n7506 = 1_n12778 | 1_n11922;
assign 1_n4590 = ~(1_n7709 ^ 1_n10000);
assign 1_n3971 = 1_n3018 & 1_n6951;
assign 1_n10754 = 1_n12402 & 1_n10456;
assign 1_n5670 = ~1_n7812;
assign 1_n3071 = 1_n2381 & 1_n5778;
assign 1_n6777 = 1_n10334 | 1_n10179;
assign 1_n11010 = 1_n4642 | 1_n2626;
assign 1_n2325 = ~1_n10904;
assign 1_n9769 = 1_n4289 & 1_n8878;
assign 1_n1431 = 1_n2558 | 1_n4056;
assign 1_n1640 = ~(1_n10782 | 1_n12379);
assign 1_n6343 = 1_n11207 & 1_n3033;
assign 1_n5878 = 1_n10988 & 1_n4831;
assign 1_n5002 = ~1_n7697;
assign 1_n12235 = ~(1_n3687 ^ 1_n10803);
assign 1_n12846 = ~1_n892;
assign 1_n1332 = 1_n5205 | 1_n2907;
assign 1_n3504 = ~(1_n95 | 1_n146);
assign 1_n9838 = ~1_n12020;
assign 1_n3892 = ~1_n2498;
assign 1_n2527 = 1_n5942 & 1_n5892;
assign 1_n8528 = ~(1_n7845 ^ 1_n13098);
assign 1_n6102 = ~(1_n7713 ^ 1_n5311);
assign 1_n6618 = 1_n11341 & 1_n1954;
assign 1_n10575 = ~(1_n1667 ^ 1_n11372);
assign 1_n6635 = 1_n4696;
assign 1_n2742 = ~1_n1611;
assign 1_n12789 = ~1_n11030;
assign 1_n11651 = 1_n4185 | 1_n8268;
assign 1_n9450 = ~1_n10805;
assign 1_n2021 = 1_n3092 & 1_n11740;
assign 1_n7624 = ~(1_n5938 | 1_n2410);
assign 1_n3941 = ~(1_n3189 | 1_n682);
assign 1_n4762 = 1_n4759 & 1_n2665;
assign 1_n5409 = ~1_n8684;
assign 1_n5542 = 1_n4995 | 1_n9792;
assign 1_n10930 = ~(1_n3880 ^ 1_n11670);
assign 1_n1558 = 1_n2994 & 1_n10713;
assign 1_n2473 = ~1_n10343;
assign 1_n10042 = ~(1_n7369 ^ 1_n7808);
assign 1_n2688 = ~1_n817;
assign 1_n608 = 1_n10580 | 1_n815;
assign 1_n105 = ~(1_n4038 ^ 1_n4424);
assign 1_n6980 = 1_n6479 | 1_n1653;
assign 1_n12664 = 1_n2175 | 1_n7873;
assign 1_n4729 = 1_n10682 & 1_n10896;
assign 1_n3362 = ~(1_n3633 ^ 1_n12863);
assign 1_n9181 = ~1_n1636;
assign 1_n4186 = 1_n139 & 1_n3853;
assign 1_n1079 = ~(1_n3919 | 1_n12108);
assign 1_n3909 = 1_n5671 & 1_n8290;
assign 1_n10997 = 1_n4087 | 1_n8686;
assign 1_n11359 = ~(1_n1815 | 1_n3555);
assign 1_n12140 = 1_n4104 & 1_n8186;
assign 1_n1281 = ~(1_n4589 ^ 1_n11503);
assign 1_n6598 = ~(1_n11378 ^ 1_n1661);
assign 1_n5309 = ~(1_n2186 ^ 1_n92);
assign 1_n3781 = 1_n5500 | 1_n11475;
assign 1_n7039 = ~(1_n1809 | 1_n4287);
assign 1_n1240 = 1_n6721 | 1_n1144;
assign 1_n6617 = ~(1_n10584 ^ 1_n9911);
assign 1_n821 = ~1_n6357;
assign 1_n5563 = ~(1_n3333 ^ 1_n7478);
assign 1_n889 = 1_n5999 | 1_n2599;
assign 1_n3236 = ~(1_n9042 | 1_n10612);
assign 1_n4283 = 1_n6486 | 1_n4640;
assign 1_n9283 = ~1_n12373;
assign 1_n4613 = ~(1_n12697 ^ 1_n7640);
assign 1_n5291 = 1_n12253 & 1_n3486;
assign 1_n5896 = 1_n9113 | 1_n8490;
assign 1_n12273 = 1_n5550;
assign 1_n12867 = ~(1_n4400 ^ 1_n3994);
assign 1_n10904 = 1_n934 & 1_n6674;
assign 1_n6582 = 1_n8085 & 1_n4679;
assign 1_n6657 = 1_n13168 | 1_n12188;
assign 1_n7119 = ~1_n3076;
assign 1_n10902 = ~(1_n8986 | 1_n11601);
assign 1_n2708 = ~(1_n12355 ^ 1_n12264);
assign 1_n9492 = ~1_n411;
assign 1_n11387 = 1_n9718 & 1_n5933;
assign 1_n4224 = 1_n8672 | 1_n12188;
assign 1_n7643 = 1_n12130 & 1_n12181;
assign 1_n1280 = 1_n6644 ^ 1_n2547;
assign 1_n11531 = 1_n10491 & 1_n13180;
assign 1_n11365 = ~1_n1717;
assign 1_n5306 = 1_n1671 | 1_n7323;
assign 1_n7584 = ~(1_n2219 ^ 1_n7509);
assign 1_n10353 = 1_n207 | 1_n12290;
assign 1_n12993 = 1_n2762 ^ 1_n11154;
assign 1_n1862 = ~(1_n8690 ^ 1_n6995);
assign 1_n5537 = 1_n2228 | 1_n1570;
assign 1_n519 = 1_n8050 | 1_n663;
assign 1_n8767 = 1_n12667 & 1_n1787;
assign 1_n11442 = 1_n3071 | 1_n341;
assign 1_n3122 = 1_n6769 | 1_n6265;
assign 1_n11972 = ~1_n11939;
assign 1_n13214 = 1_n10681 | 1_n12596;
assign 1_n5498 = ~(1_n1603 ^ 1_n3455);
assign 1_n5839 = ~1_n8311;
assign 1_n7181 = 1_n3908 | 1_n1144;
assign 1_n1731 = ~(1_n10911 ^ 1_n8201);
assign 1_n3540 = ~(1_n4147 ^ 1_n1981);
assign 1_n11354 = ~1_n10642;
assign 1_n10585 = 1_n10586 | 1_n12126;
assign 1_n6449 = 1_n6753 | 1_n8573;
assign 1_n11272 = ~(1_n7398 ^ 1_n8287);
assign 1_n11766 = ~(1_n9341 ^ 1_n2161);
assign 1_n30 = 1_n554 & 1_n3975;
assign 1_n3611 = ~(1_n7767 ^ 1_n10372);
assign 1_n11009 = 1_n7780 | 1_n10106;
assign 1_n12815 = 1_n1070 & 1_n12169;
assign 1_n7015 = 1_n5972 | 1_n4987;
assign 1_n7709 = ~1_n9515;
assign 1_n10460 = 1_n106 | 1_n1266;
assign 1_n5446 = ~1_n6707;
assign 1_n12116 = 1_n1973 & 1_n6302;
assign 1_n4632 = ~(1_n12670 ^ 1_n10971);
assign 1_n6707 = 1_n1402 | 1_n9223;
assign 1_n8534 = 1_n6596;
assign 1_n11540 = ~1_n8745;
assign 1_n8334 = 1_n10924 | 1_n2787;
assign 1_n8713 = ~(1_n3796 ^ 1_n5325);
assign 1_n11698 = ~(1_n11733 ^ 1_n9815);
assign 1_n3612 = ~(1_n8814 ^ 1_n9560);
assign 1_n4080 = ~1_n497;
assign 1_n8069 = ~(1_n3810 ^ 1_n4918);
assign 1_n6648 = ~(1_n9331 ^ 1_n4625);
assign 1_n822 = 1_n7926 & 1_n1334;
assign 1_n4196 = 1_n1391 & 1_n10967;
assign 1_n12695 = 1_n2278;
assign 1_n6533 = ~1_n4188;
assign 1_n6605 = ~(1_n2312 ^ 1_n12685);
assign 1_n11235 = 1_n1402 | 1_n2059;
assign 1_n2917 = 1_n8751 & 1_n8344;
assign 1_n4577 = ~(1_n8366 ^ 1_n7176);
assign 1_n9402 = ~1_n7896;
assign 1_n5797 = 1_n2278;
assign 1_n9586 = ~1_n12248;
assign 1_n2144 = 1_n2538 | 1_n3949;
assign 1_n13066 = 1_n6908 | 1_n5819;
assign 1_n3843 = 1_n5900 & 1_n9781;
assign 1_n5596 = 1_n1332 & 1_n11463;
assign 1_n9443 = 1_n7068 | 1_n9159;
assign 1_n12171 = ~1_n4651;
assign 1_n4571 = ~(1_n12981 | 1_n6272);
assign 1_n5244 = ~(1_n7869 ^ 1_n754);
assign 1_n9106 = 1_n12322 & 1_n12374;
assign 1_n6213 = ~(1_n7926 ^ 1_n236);
assign 1_n8835 = ~1_n2577;
assign 1_n6951 = 1_n12469 | 1_n12273;
assign 1_n164 = 1_n4761 & 1_n6013;
assign 1_n12310 = 1_n10775 | 1_n9956;
assign 1_n8373 = ~(1_n12073 ^ 1_n8003);
assign 1_n3761 = ~1_n10288;
assign 1_n4279 = 1_n7966 | 1_n6404;
assign 1_n1803 = ~(1_n5399 | 1_n7405);
assign 1_n9134 = 1_n1652 & 1_n10419;
assign 1_n10035 = ~1_n2212;
assign 1_n8559 = 1_n6595 | 1_n7935;
assign 1_n10192 = ~(1_n12518 ^ 1_n12024);
assign 1_n9580 = 1_n3365 ^ 1_n11819;
assign 1_n3733 = ~(1_n3868 | 1_n11143);
assign 1_n12311 = 1_n5803 | 1_n3193;
assign 1_n158 = ~(1_n13050 ^ 1_n5106);
assign 1_n3786 = 1_n4451 | 1_n5725;
assign 1_n8843 = ~1_n1302;
assign 1_n5867 = 1_n11455 | 1_n10374;
assign 1_n825 = ~(1_n11562 ^ 1_n12497);
assign 1_n10443 = ~(1_n12437 | 1_n3799);
assign 1_n267 = 1_n10314 | 1_n12959;
assign 1_n2500 = 1_n5207 & 1_n3707;
assign 1_n10564 = 1_n11014 & 1_n4770;
assign 1_n4938 = 1_n7283 | 1_n12273;
assign 1_n4388 = ~(1_n4500 | 1_n1);
assign 1_n2345 = 1_n3619 | 1_n13053;
assign 1_n10263 = ~1_n10162;
assign 1_n2370 = 1_n1218 | 1_n5242;
assign 1_n2387 = ~1_n6168;
assign 1_n5199 = 1_n13063 | 1_n5493;
assign 1_n10519 = ~1_n12078;
assign 1_n11194 = 1_n7091 | 1_n3438;
assign 1_n1417 = 1_n11420 & 1_n2363;
assign 1_n11817 = 1_n3750 & 1_n11399;
assign 1_n2019 = ~(1_n10496 | 1_n5159);
assign 1_n5248 = 1_n3325 & 1_n4942;
assign 1_n1068 = 1_n10979 ^ 1_n8875;
assign 1_n8642 = 1_n11703 & 1_n8853;
assign 1_n976 = 1_n2717 & 1_n6920;
assign 1_n3484 = ~(1_n10967 | 1_n1391);
assign 1_n9351 = ~(1_n11602 ^ 1_n8100);
assign 1_n11437 = ~(1_n5621 | 1_n5533);
assign 1_n7203 = ~(1_n6656 | 1_n10036);
assign 1_n13070 = ~(1_n914 | 1_n592);
assign 1_n2939 = 1_n9253 & 1_n7972;
assign 1_n3304 = 1_n696 | 1_n9352;
assign 1_n8111 = ~1_n1792;
assign 1_n408 = 1_n5968 | 1_n10179;
assign 1_n7457 = 1_n1554 | 1_n6133;
assign 1_n6565 = 1_n9757 & 1_n6131;
assign 1_n120 = ~(1_n12035 ^ 1_n2939);
assign 1_n10638 = ~(1_n8487 ^ 1_n10394);
assign 1_n8056 = ~(1_n8061 ^ 1_n6084);
assign 1_n9007 = ~(1_n1282 ^ 1_n11529);
assign 1_n10790 = ~(1_n2650 ^ 1_n3569);
assign 1_n2796 = ~(1_n6536 | 1_n4866);
assign 1_n10666 = ~1_n594;
assign 1_n5143 = ~(1_n8942 ^ 1_n6632);
assign 1_n1414 = ~(1_n5850 ^ 1_n187);
assign 1_n2667 = 1_n4205 & 1_n1351;
assign 1_n9631 = ~(1_n9708 ^ 1_n684);
assign 1_n11210 = 1_n13194 | 1_n10319;
assign 1_n13183 = ~1_n2295;
assign 1_n1245 = 1_n1018 & 1_n764;
assign 1_n88 = ~(1_n7583 ^ 1_n6168);
assign 1_n10610 = 1_n5944 | 1_n7305;
assign 1_n8561 = ~1_n9093;
assign 1_n4894 = ~(1_n7657 ^ 1_n6795);
assign 1_n565 = 1_n5588 | 1_n10029;
assign 1_n10646 = 1_n1434 | 1_n3459;
assign 1_n156 = ~1_n6489;
assign 1_n10954 = ~(1_n12622 ^ 1_n6470);
assign 1_n12246 = ~1_n2765;
assign 1_n9985 = ~(1_n4368 | 1_n7716);
assign 1_n10504 = ~(1_n3122 ^ 1_n6477);
assign 1_n5503 = 1_n7532 | 1_n6635;
assign 1_n11261 = ~(1_n6668 | 1_n7812);
assign 1_n3222 = ~1_n4457;
assign 1_n2617 = 1_n4929 & 1_n12060;
assign 1_n1591 = ~(1_n676 ^ 1_n6432);
assign 1_n9252 = 1_n3224 & 1_n1888;
assign 1_n11471 = ~1_n5747;
assign 1_n1164 = ~(1_n4313 ^ 1_n12029);
assign 1_n9756 = ~(1_n11160 ^ 1_n8069);
assign 1_n10156 = ~(1_n1380 ^ 1_n5254);
assign 1_n10351 = 1_n10587 | 1_n9159;
assign 1_n11822 = 1_n10136 & 1_n3174;
assign 1_n5337 = 1_n5558 | 1_n13043;
assign 1_n10558 = ~1_n12579;
assign 1_n3186 = 1_n2931 & 1_n7313;
assign 1_n12991 = ~(1_n331 ^ 1_n11994);
assign 1_n3075 = ~(1_n12381 | 1_n4589);
assign 1_n9033 = ~1_n5498;
assign 1_n10383 = ~1_n2174;
assign 1_n2938 = 1_n10631 & 1_n10329;
assign 1_n535 = ~(1_n10327 ^ 1_n10074);
assign 1_n2139 = ~(1_n9945 ^ 1_n3513);
assign 1_n12907 = ~(1_n6273 | 1_n12145);
assign 1_n12034 = ~(1_n9039 ^ 1_n2775);
assign 1_n1970 = 1_n513 | 1_n9027;
assign 1_n11305 = ~(1_n3834 ^ 1_n9411);
assign 1_n8015 = ~(1_n9870 ^ 1_n1104);
assign 1_n7669 = 1_n11781 | 1_n902;
assign 1_n8644 = ~1_n9474;
assign 1_n7321 = 1_n1126 & 1_n13083;
assign 1_n493 = ~1_n12853;
assign 1_n4812 = 1_n12569 & 1_n7508;
assign 1_n10806 = 1_n9619 & 1_n5382;
assign 1_n2250 = 1_n2753 & 1_n7593;
assign 1_n5494 = ~1_n6043;
assign 1_n2023 = 1_n2725 & 1_n13228;
assign 1_n12776 = ~(1_n7316 ^ 1_n4510);
assign 1_n11303 = ~(1_n2656 ^ 1_n323);
assign 1_n1263 = ~1_n4789;
assign 1_n7420 = 1_n1485 | 1_n5931;
assign 1_n8813 = ~(1_n11278 ^ 1_n8482);
assign 1_n7013 = ~1_n4259;
assign 1_n4 = 1_n11242 | 1_n2133;
assign 1_n8825 = 1_n2504 | 1_n8563;
assign 1_n12812 = ~1_n10654;
assign 1_n2909 = ~(1_n2069 ^ 1_n9030);
assign 1_n7637 = ~(1_n8358 ^ 1_n3087);
assign 1_n10525 = ~1_n1988;
assign 1_n7764 = ~(1_n10812 ^ 1_n5074);
assign 1_n1121 = ~(1_n6555 ^ 1_n12338);
assign 1_n8654 = ~1_n9580;
assign 1_n5998 = 1_n5659 ^ 1_n11988;
assign 1_n4145 = 1_n8510 | 1_n8702;
assign 1_n13009 = 1_n10558 | 1_n7723;
assign 1_n9553 = ~(1_n7555 ^ 1_n2864);
assign 1_n4389 = 1_n11249 & 1_n13207;
assign 1_n11115 = 1_n5574 | 1_n5604;
assign 1_n1583 = ~(1_n6305 ^ 1_n984);
assign 1_n2751 = 1_n1905 & 1_n2608;
assign 1_n8026 = ~1_n1498;
assign 1_n10988 = ~1_n13034;
assign 1_n3678 = ~(1_n2431 ^ 1_n11169);
assign 1_n2580 = ~1_n11671;
assign 1_n4626 = ~(1_n7585 ^ 1_n9947);
assign 1_n2888 = ~(1_n4035 ^ 1_n8902);
assign 1_n7771 = ~1_n12340;
assign 1_n1794 = 1_n12230 & 1_n4204;
assign 1_n8668 = 1_n7000 | 1_n10937;
assign 1_n8459 = ~(1_n11899 ^ 1_n2926);
assign 1_n2015 = 1_n2031 | 1_n10130;
assign 1_n3326 = 1_n950 | 1_n3257;
assign 1_n2613 = 1_n10474 | 1_n5782;
assign 1_n7700 = ~1_n13060;
assign 1_n7353 = 1_n5883 & 1_n7653;
assign 1_n3179 = ~(1_n10259 | 1_n12454);
assign 1_n5441 = 1_n5973 | 1_n8563;
assign 1_n3995 = 1_n103 & 1_n10408;
assign 1_n5233 = 1_n9606 | 1_n12188;
assign 1_n3559 = 1_n6135 & 1_n4859;
assign 1_n3334 = ~1_n11386;
assign 1_n10074 = ~(1_n6711 ^ 1_n2523);
assign 1_n10096 = 1_n6726 | 1_n7530;
assign 1_n9126 = ~(1_n6431 | 1_n8826);
assign 1_n4060 = ~(1_n5098 ^ 1_n3647);
assign 1_n1200 = 1_n13181 | 1_n1589;
assign 1_n7105 = 1_n6658 | 1_n7221;
assign 1_n3716 = 1_n8471 & 1_n6688;
assign 1_n9657 = 1_n11313 & 1_n883;
assign 1_n3717 = ~(1_n4710 | 1_n3840);
assign 1_n9118 = ~1_n5962;
assign 1_n5139 = 1_n6595 | 1_n7903;
assign 1_n5722 = 1_n10144 & 1_n8545;
assign 1_n6739 = 1_n3465 | 1_n10222;
assign 1_n9765 = ~1_n4968;
assign 1_n10576 = ~(1_n12994 | 1_n4422);
assign 1_n3748 = ~(1_n9151 ^ 1_n2664);
assign 1_n4240 = ~(1_n1116 ^ 1_n3670);
assign 1_n1868 = 1_n8392 | 1_n9159;
assign 1_n11361 = 1_n1360 | 1_n3531;
assign 1_n8834 = ~1_n90;
assign 1_n7212 = ~(1_n7427 ^ 1_n9203);
assign 1_n9697 = ~1_n2011;
assign 1_n12930 = ~1_n4470;
assign 1_n6413 = ~(1_n2739 ^ 1_n975);
assign 1_n1993 = ~(1_n5025 ^ 1_n523);
assign 1_n12650 = ~(1_n9974 ^ 1_n11747);
assign 1_n11242 = ~1_n12408;
assign 1_n3702 = 1_n13163 & 1_n2440;
assign 1_n8504 = ~1_n429;
assign 1_n2442 = 1_n813 | 1_n10029;
assign 1_n10271 = ~(1_n6539 ^ 1_n12257);
assign 1_n8039 = ~1_n5513;
assign 1_n4623 = ~(1_n9168 ^ 1_n9639);
assign 1_n2630 = 1_n11366 ^ 1_n4269;
assign 1_n9265 = ~1_n10231;
assign 1_n11781 = ~1_n4470;
assign 1_n5713 = ~1_n12651;
assign 1_n7657 = 1_n6733 | 1_n1570;
assign 1_n10957 = ~(1_n8417 | 1_n10011);
assign 1_n9025 = 1_n7184 | 1_n6635;
assign 1_n13242 = ~1_n11537;
assign 1_n4680 = ~1_n3447;
assign 1_n7577 = 1_n5544 ^ 1_n10149;
assign 1_n11462 = 1_n10429 | 1_n252;
assign 1_n9817 = ~(1_n12797 ^ 1_n4726);
assign 1_n11882 = ~(1_n8520 ^ 1_n4329);
assign 1_n5384 = ~(1_n8811 ^ 1_n6932);
assign 1_n10851 = 1_n2985 | 1_n9704;
assign 1_n12040 = ~(1_n8794 ^ 1_n11814);
assign 1_n8001 = 1_n7065 & 1_n12180;
assign 1_n6768 = ~1_n4006;
assign 1_n2531 = ~(1_n12710 | 1_n4193);
assign 1_n7346 = ~1_n5933;
assign 1_n6281 = 1_n3363 & 1_n2680;
assign 1_n6197 = 1_n10796 ^ 1_n12058;
assign 1_n1136 = 1_n10900 | 1_n2449;
assign 1_n6421 = ~1_n7670;
assign 1_n585 = ~1_n1432;
assign 1_n6294 = ~(1_n6130 ^ 1_n8780);
assign 1_n9295 = 1_n7269 & 1_n9342;
assign 1_n7850 = 1_n5595 | 1_n2875;
assign 1_n5927 = ~1_n10004;
assign 1_n11604 = ~(1_n11655 ^ 1_n738);
assign 1_n3856 = 1_n7941 | 1_n4868;
assign 1_n5711 = 1_n3697 | 1_n7655;
assign 1_n4246 = ~(1_n11987 ^ 1_n3019);
assign 1_n1088 = ~(1_n11998 ^ 1_n6051);
assign 1_n617 = ~1_n8233;
assign 1_n12644 = ~(1_n15 ^ 1_n3056);
assign 1_n5411 = 1_n2013 | 1_n6484;
assign 1_n8566 = 1_n11258 & 1_n11967;
assign 1_n4753 = 1_n7124 | 1_n11550;
assign 1_n4965 = 1_n13084 | 1_n12501;
assign 1_n2943 = ~1_n13058;
assign 1_n4954 = 1_n3128 & 1_n3203;
assign 1_n6476 = ~(1_n3627 ^ 1_n13212);
assign 1_n8269 = ~(1_n10999 ^ 1_n10342);
assign 1_n8618 = 1_n4584 | 1_n4373;
assign 1_n415 = ~(1_n9261 ^ 1_n11977);
assign 1_n12335 = ~1_n12003;
assign 1_n11208 = ~(1_n1205 | 1_n2649);
assign 1_n3952 = ~(1_n12362 ^ 1_n3987);
assign 1_n7983 = ~(1_n1395 | 1_n8781);
assign 1_n3482 = ~(1_n10371 ^ 1_n13015);
assign 1_n2700 = 1_n579 & 1_n7977;
assign 1_n9884 = 1_n7018 | 1_n3016;
assign 1_n1656 = ~(1_n2107 | 1_n8548);
assign 1_n452 = 1_n216 | 1_n7445;
assign 1_n241 = ~1_n9534;
assign 1_n13169 = 1_n2711 | 1_n9268;
assign 1_n8004 = ~(1_n12186 | 1_n6163);
assign 1_n12422 = 1_n7919 ^ 1_n11056;
assign 1_n4818 = ~1_n1612;
assign 1_n4927 = 1_n5666 | 1_n12273;
assign 1_n12923 = ~(1_n8889 ^ 1_n6022);
assign 1_n2792 = 1_n5923 | 1_n1026;
assign 1_n6835 = 1_n3347 | 1_n5036;
assign 1_n11142 = 1_n4514 | 1_n11244;
assign 1_n1888 = 1_n1621 | 1_n2133;
assign 1_n1152 = ~1_n10451;
assign 1_n10316 = 1_n3587 | 1_n9223;
assign 1_n7000 = ~(1_n8028 ^ 1_n4162);
assign 1_n3850 = ~(1_n3628 ^ 1_n9218);
assign 1_n2941 = ~1_n5066;
assign 1_n6012 = 1_n11886 & 1_n4025;
assign 1_n8839 = ~(1_n4876 ^ 1_n769);
assign 1_n8445 = 1_n3732 & 1_n7438;
assign 1_n7429 = 1_n9332 & 1_n5818;
assign 1_n6712 = 1_n5890 | 1_n8534;
assign 1_n11315 = 1_n12514 | 1_n514;
assign 1_n3955 = ~(1_n11306 | 1_n8432);
assign 1_n11605 = ~1_n7326;
assign 1_n1536 = ~1_n8332;
assign 1_n1455 = ~(1_n9236 ^ 1_n5023);
assign 1_n10526 = 1_n12517 & 1_n7303;
assign 1_n11319 = ~(1_n8800 ^ 1_n7628);
assign 1_n12018 = 1_n13061 | 1_n1212;
assign 1_n7142 = ~1_n1198;
assign 1_n5923 = ~1_n5189;
assign 1_n7798 = ~1_n2339;
assign 1_n2900 = 1_n8556 | 1_n11772;
assign 1_n12014 = 1_n1268 ^ 1_n3865;
assign 1_n9686 = 1_n11943 & 1_n2305;
assign 1_n581 = 1_n4737 & 1_n1785;
assign 1_n11192 = 1_n2689 | 1_n8702;
assign 1_n432 = 1_n8141 | 1_n11510;
assign 1_n8125 = 1_n8183 & 1_n5920;
assign 1_n6562 = 1_n4905 & 1_n10703;
assign 1_n2400 = 1_n1406 | 1_n5999;
assign 1_n5890 = ~1_n2737;
assign 1_n1782 = 1_n3266 & 1_n2224;
assign 1_n2096 = 1_n5004 | 1_n4314;
assign 1_n10554 = ~(1_n10921 ^ 1_n11675);
assign 1_n8836 = ~1_n3116;
assign 1_n3550 = 1_n1669 & 1_n1185;
assign 1_n2921 = ~(1_n2439 ^ 1_n1049);
assign 1_n12406 = ~(1_n1655 ^ 1_n10082);
assign 1_n12505 = ~(1_n12867 | 1_n11079);
assign 1_n7717 = ~(1_n6009 ^ 1_n9055);
assign 1_n8664 = ~1_n7090;
assign 1_n4538 = 1_n7142 | 1_n2675;
assign 1_n6602 = 1_n8697 | 1_n10648;
assign 1_n4097 = 1_n6988 | 1_n11591;
assign 1_n9644 = ~(1_n3848 ^ 1_n7484);
assign 1_n7425 = ~(1_n11189 ^ 1_n6512);
assign 1_n11069 = 1_n10954 | 1_n4504;
assign 1_n6484 = 1_n6132 ^ 1_n6094;
assign 1_n9183 = ~(1_n4224 ^ 1_n9864);
assign 1_n2561 = ~(1_n6690 ^ 1_n7141);
assign 1_n3908 = ~1_n6655;
assign 1_n10024 = 1_n10800 & 1_n8019;
assign 1_n7422 = ~(1_n744 | 1_n12484);
assign 1_n8020 = ~1_n1709;
assign 1_n2723 = ~1_n8768;
assign 1_n11706 = 1_n1387 | 1_n4565;
assign 1_n12552 = ~1_n11891;
assign 1_n4319 = ~(1_n9213 ^ 1_n7651);
assign 1_n9828 = ~1_n1573;
assign 1_n6831 = ~(1_n4146 ^ 1_n4623);
assign 1_n10720 = ~(1_n9519 ^ 1_n6541);
assign 1_n7063 = ~(1_n4012 | 1_n8189);
assign 1_n6192 = ~(1_n978 ^ 1_n11009);
assign 1_n5459 = 1_n11718 | 1_n5081;
assign 1_n10330 = ~(1_n7763 ^ 1_n5578);
assign 1_n10210 = ~1_n7637;
assign 1_n948 = ~(1_n10795 ^ 1_n12667);
assign 1_n4826 = 1_n12441 | 1_n4063;
assign 1_n1232 = 1_n1420 & 1_n8387;
assign 1_n137 = ~(1_n3069 ^ 1_n8365);
assign 1_n8807 = ~(1_n12472 ^ 1_n1926);
assign 1_n3041 = ~1_n9381;
assign 1_n5147 = ~(1_n2814 ^ 1_n12123);
assign 1_n5511 = 1_n9422 | 1_n1109;
assign 1_n11390 = ~(1_n7002 ^ 1_n7308);
assign 1_n10157 = 1_n11903 | 1_n5765;
assign 1_n3814 = 1_n555 | 1_n5677;
assign 1_n6645 = ~1_n3645;
assign 1_n1324 = ~1_n4233;
assign 1_n5243 = ~1_n741;
assign 1_n1406 = ~1_n9887;
assign 1_n400 = 1_n2566 | 1_n7624;
assign 1_n8689 = 1_n1495 ^ 1_n4518;
assign 1_n3057 = ~(1_n3394 ^ 1_n12392);
assign 1_n12053 = ~(1_n672 | 1_n2912);
assign 1_n1779 = 1_n9767 | 1_n8030;
assign 1_n12456 = ~(1_n8470 | 1_n5469);
assign 1_n1361 = 1_n10232 & 1_n9520;
assign 1_n12099 = ~1_n9849;
assign 1_n3545 = 1_n3369 | 1_n6227;
assign 1_n70 = ~(1_n7240 ^ 1_n735);
assign 1_n5649 = 1_n12834 | 1_n2449;
assign 1_n5677 = 1_n8663 & 1_n6476;
assign 1_n12133 = 1_n8466 & 1_n7720;
assign 1_n1100 = ~(1_n6842 ^ 1_n86);
assign 1_n3439 = 1_n7377 | 1_n9075;
assign 1_n3481 = 1_n12418 & 1_n11713;
assign 1_n10492 = ~1_n12389;
assign 1_n12726 = 1_n10772 | 1_n11144;
assign 1_n1249 = ~(1_n9056 ^ 1_n7612);
assign 1_n1208 = ~(1_n12824 ^ 1_n6897);
assign 1_n3509 = ~1_n3112;
assign 1_n11156 = 1_n7891 | 1_n8048;
assign 1_n5178 = ~(1_n3354 ^ 1_n10367);
assign 1_n4700 = 1_n12838 & 1_n4479;
assign 1_n6159 = 1_n6738 | 1_n9486;
assign 1_n80 = ~1_n951;
assign 1_n4128 = 1_n10281 | 1_n206;
assign 1_n7568 = 1_n8035 | 1_n6565;
assign 1_n6310 = ~(1_n4277 ^ 1_n9908);
assign 1_n6453 = 1_n7033 | 1_n5521;
assign 1_n6219 = ~1_n841;
assign 1_n2826 = 1_n79 | 1_n4442;
assign 1_n6953 = 1_n12000 | 1_n4253;
assign 1_n6748 = 1_n3892 | 1_n12069;
assign 1_n11001 = ~(1_n10918 ^ 1_n3528);
assign 1_n7663 = ~(1_n4772 ^ 1_n12495);
assign 1_n8958 = ~(1_n11064 ^ 1_n5237);
assign 1_n1344 = 1_n3602 & 1_n6807;
assign 1_n2070 = 1_n8950 | 1_n6635;
assign 1_n13134 = 1_n5520 | 1_n10761;
assign 1_n10359 = 1_n1706 | 1_n4643;
assign 1_n356 = 1_n8221 & 1_n7261;
assign 1_n276 = ~(1_n9456 | 1_n1754);
assign 1_n8089 = ~(1_n10690 ^ 1_n10095);
assign 1_n8285 = ~1_n6142;
assign 1_n8971 = ~1_n253;
assign 1_n6706 = ~1_n1486;
assign 1_n2195 = 1_n13056 & 1_n385;
assign 1_n2935 = 1_n521 & 1_n11039;
assign 1_n876 = 1_n5125 | 1_n12077;
assign 1_n12369 = ~(1_n7889 ^ 1_n2685);
assign 1_n11106 = ~1_n12784;
assign 1_n11894 = ~(1_n2851 ^ 1_n9121);
assign 1_n6890 = 1_n11009 | 1_n12387;
assign 1_n374 = 1_n7017 & 1_n1970;
assign 1_n11762 = ~(1_n921 ^ 1_n10650);
assign 1_n7712 = ~(1_n9448 | 1_n6483);
assign 1_n6622 = ~(1_n6208 ^ 1_n352);
assign 1_n8620 = 1_n6846 | 1_n3703;
assign 1_n9854 = 1_n12084 | 1_n13054;
assign 1_n2719 = ~(1_n13223 ^ 1_n12822);
assign 1_n47 = ~1_n5551;
assign 1_n9716 = 1_n1903 | 1_n10931;
assign 1_n1460 = 1_n7047 | 1_n12783;
assign 1_n2928 = ~(1_n6527 ^ 1_n7278);
assign 1_n12848 = ~1_n13120;
assign 1_n325 = 1_n5031 & 1_n8506;
assign 1_n8683 = 1_n2232 | 1_n2958;
assign 1_n8344 = 1_n1559 | 1_n6919;
assign 1_n1683 = 1_n1571 | 1_n7530;
assign 1_n9069 = ~1_n6392;
assign 1_n38 = 1_n6672 | 1_n13238;
assign 1_n6723 = 1_n5943 | 1_n8730;
assign 1_n3876 = ~(1_n3536 ^ 1_n6857);
assign 1_n4553 = ~(1_n10790 ^ 1_n4083);
assign 1_n2202 = ~(1_n12394 ^ 1_n11863);
assign 1_n7861 = 1_n7620 | 1_n9195;
assign 1_n4320 = 1_n7529 & 1_n7772;
assign 1_n12694 = 1_n231 & 1_n8906;
assign 1_n8592 = ~1_n4008;
assign 1_n2320 = ~(1_n12260 | 1_n11433);
assign 1_n5009 = 1_n4184 | 1_n12725;
assign 1_n12742 = 1_n8839 ^ 1_n1281;
assign 1_n6806 = 1_n11599 | 1_n7892;
assign 1_n8409 = ~(1_n3642 ^ 1_n5196);
assign 1_n5176 = ~1_n8768;
assign 1_n2415 = ~1_n4740;
assign 1_n4788 = 1_n4803 ^ 1_n256;
assign 1_n523 = 1_n12918 & 1_n5246;
assign 1_n7487 = ~(1_n10913 | 1_n3746);
assign 1_n3498 = ~1_n4470;
assign 1_n12005 = 1_n10851 & 1_n3275;
assign 1_n5781 = 1_n9509 & 1_n357;
assign 1_n8991 = ~(1_n9448 ^ 1_n7389);
assign 1_n8403 = ~(1_n4654 ^ 1_n1958);
assign 1_n3891 = ~(1_n7474 | 1_n4068);
assign 1_n4417 = ~(1_n9554 ^ 1_n3849);
assign 1_n440 = 1_n12871 | 1_n12388;
assign 1_n3087 = 1_n6769 | 1_n1026;
assign 1_n10079 = 1_n7331 & 1_n5204;
assign 1_n8436 = ~1_n12603;
assign 1_n4835 = 1_n13215 & 1_n150;
assign 1_n11725 = ~(1_n9523 ^ 1_n11656);
assign 1_n7706 = 1_n6724 | 1_n7723;
assign 1_n3370 = ~(1_n4251 ^ 1_n3079);
assign 1_n10986 = ~1_n11445;
assign 1_n4614 = ~(1_n4101 ^ 1_n9357);
assign 1_n2207 = ~1_n8455;
assign 1_n5296 = 1_n4667 & 1_n10546;
assign 1_n3901 = 1_n7884 | 1_n12426;
assign 1_n9933 = 1_n10228 & 1_n3915;
assign 1_n9821 = ~1_n8036;
assign 1_n10399 = ~(1_n10499 ^ 1_n6893);
assign 1_n1763 = 1_n3299 | 1_n8301;
assign 1_n3324 = ~(1_n6294 ^ 1_n3034);
assign 1_n13045 = ~(1_n5505 | 1_n13171);
assign 1_n8672 = ~1_n9669;
assign 1_n4361 = ~1_n1228;
assign 1_n1770 = 1_n5314 & 1_n188;
assign 1_n4687 = 1_n9153 & 1_n12001;
assign 1_n2266 = 1_n8528 | 1_n13237;
assign 1_n5105 = ~1_n4006;
assign 1_n11746 = 1_n9928 & 1_n9445;
assign 1_n7159 = ~1_n3064;
assign 1_n12628 = ~(1_n786 | 1_n4428);
assign 1_n632 = ~(1_n12637 ^ 1_n2046);
assign 1_n3025 = ~1_n7316;
assign 1_n46 = 1_n2826 & 1_n10965;
assign 1_n1743 = ~(1_n8689 ^ 1_n6516);
assign 1_n1618 = ~1_n7720;
assign 1_n10319 = 1_n13005;
assign 1_n833 = ~(1_n2088 | 1_n5851);
assign 1_n6594 = ~(1_n12707 | 1_n5333);
assign 1_n3783 = ~1_n7360;
assign 1_n12771 = 1_n11171 | 1_n12273;
assign 1_n2152 = 1_n3345 & 1_n8112;
assign 1_n8818 = ~(1_n10920 ^ 1_n5975);
assign 1_n3132 = ~1_n3711;
assign 1_n1856 = ~(1_n10033 | 1_n8669);
assign 1_n5071 = 1_n2652 & 1_n11369;
assign 1_n1226 = ~1_n1312;
assign 1_n7528 = 1_n8146 & 1_n169;
assign 1_n485 = 1_n2535 ^ 1_n11741;
assign 1_n12956 = ~(1_n11567 ^ 1_n4999);
assign 1_n4093 = 1_n10760 & 1_n5330;
assign 1_n1750 = ~1_n8228;
assign 1_n504 = 1_n3445 & 1_n6581;
assign 1_n7213 = 1_n7249 | 1_n2836;
assign 1_n11989 = 1_n10525 | 1_n2212;
assign 1_n4143 = ~1_n7113;
assign 1_n323 = 1_n508 & 1_n6393;
assign 1_n7043 = ~(1_n10743 ^ 1_n6529);
assign 1_n7588 = 1_n2858 | 1_n8097;
assign 1_n3070 = 1_n1571 | 1_n12388;
assign 1_n10516 = ~(1_n11893 ^ 1_n6350);
assign 1_n11276 = ~(1_n1547 ^ 1_n466);
assign 1_n10940 = 1_n1930 | 1_n8348;
assign 1_n9542 = ~(1_n4204 ^ 1_n4241);
assign 1_n5311 = 1_n4096 & 1_n9072;
assign 1_n2302 = 1_n4692 | 1_n2351;
assign 1_n11846 = 1_n9216 & 1_n13058;
assign 1_n4433 = 1_n6713 | 1_n2989;
assign 1_n3227 = 1_n9723 | 1_n8030;
assign 1_n7112 = 1_n4430 | 1_n68;
assign 1_n6283 = ~(1_n36 ^ 1_n5219);
assign 1_n6794 = ~(1_n1935 ^ 1_n9587);
assign 1_n8627 = 1_n1021 & 1_n8628;
assign 1_n7740 = ~(1_n2233 ^ 1_n1421);
assign 1_n3681 = ~1_n8543;
assign 1_n3683 = 1_n10481 | 1_n9075;
assign 1_n637 = ~(1_n382 ^ 1_n3967);
assign 1_n6897 = ~(1_n5188 ^ 1_n13022);
assign 1_n7630 = 1_n8396 & 1_n11383;
assign 1_n1322 = ~(1_n8539 | 1_n3525);
assign 1_n12672 = 1_n7894 & 1_n6300;
assign 1_n12457 = ~(1_n3345 ^ 1_n580);
assign 1_n7658 = 1_n1571 | 1_n8702;
assign 1_n5367 = 1_n5810 | 1_n3133;
assign 1_n10291 = ~1_n9667;
assign 1_n5144 = 1_n3516 | 1_n5547;
assign 1_n11796 = 1_n4870 & 1_n9487;
assign 1_n3963 = ~1_n3130;
assign 1_n2283 = 1_n7223 | 1_n3981;
assign 1_n10442 = 1_n5644 & 1_n7179;
assign 1_n6079 = ~(1_n7669 ^ 1_n10767);
assign 1_n1321 = ~1_n2630;
assign 1_n10877 = ~1_n4357;
assign 1_n12225 = 1_n1797 & 1_n9722;
assign 1_n12511 = 1_n7771 & 1_n3524;
assign 1_n11014 = ~1_n5777;
assign 1_n3823 = ~(1_n12675 | 1_n3629);
assign 1_n7824 = ~1_n4543;
assign 1_n10436 = 1_n993 & 1_n6353;
assign 1_n750 = ~(1_n1442 ^ 1_n9967);
assign 1_n2966 = ~(1_n877 ^ 1_n12991);
assign 1_n2735 = ~(1_n13172 ^ 1_n2567);
assign 1_n7167 = ~1_n11634;
assign 1_n4560 = 1_n4779 & 1_n7832;
assign 1_n9743 = 1_n9822 | 1_n634;
assign 1_n10329 = 1_n2914 | 1_n655;
assign 1_n11297 = ~1_n10633;
assign 1_n9868 = ~1_n9570;
assign 1_n11433 = 1_n6915 | 1_n1710;
assign 1_n11267 = 1_n4532 & 1_n7279;
assign 1_n4262 = ~(1_n6321 ^ 1_n5780);
assign 1_n6095 = 1_n3420 | 1_n6123;
assign 1_n12459 = ~(1_n12659 ^ 1_n5351);
assign 1_n12794 = ~(1_n4112 | 1_n4389);
assign 1_n8841 = ~(1_n6384 ^ 1_n13142);
assign 1_n2251 = ~(1_n11775 | 1_n12139);
assign 1_n2319 = 1_n8802 & 1_n6235;
assign 1_n9431 = ~1_n3012;
assign 1_n2582 = ~1_n9887;
assign 1_n4926 = ~(1_n9624 | 1_n4914);
assign 1_n8955 = ~(1_n7264 ^ 1_n1208);
assign 1_n7859 = 1_n1680 & 1_n451;
assign 1_n8435 = 1_n2694 & 1_n12528;
assign 1_n2934 = ~(1_n8495 ^ 1_n11048);
assign 1_n50 = ~(1_n10695 ^ 1_n12331);
assign 1_n3163 = 1_n6774 | 1_n10875;
assign 1_n12946 = ~(1_n3345 | 1_n8112);
assign 1_n6121 = ~(1_n9548 | 1_n1124);
assign 1_n1543 = 1_n11174 & 1_n13052;
assign 1_n8581 = ~(1_n8652 ^ 1_n658);
assign 1_n11016 = 1_n3442 & 1_n2191;
assign 1_n9268 = ~1_n9732;
assign 1_n13131 = ~(1_n833 | 1_n12706);
assign 1_n9515 = 1_n841 ^ 1_n6734;
assign 1_n11329 = 1_n4022 | 1_n206;
assign 1_n5947 = ~1_n8860;
assign 1_n3387 = ~1_n7436;
assign 1_n8750 = ~(1_n12979 ^ 1_n12589);
assign 1_n7097 = ~(1_n8548 ^ 1_n2107);
assign 1_n1801 = ~(1_n3436 ^ 1_n1157);
assign 1_n4050 = ~(1_n9629 | 1_n6253);
assign 1_n2020 = 1_n9158 & 1_n6902;
assign 1_n129 = 1_n7987 & 1_n12556;
assign 1_n10698 = 1_n12009 | 1_n4947;
assign 1_n11545 = ~1_n3361;
assign 1_n6603 = ~(1_n6654 ^ 1_n5180);
assign 1_n9826 = 1_n4620 | 1_n6265;
assign 1_n183 = 1_n11473 ^ 1_n2047;
assign 1_n6065 = 1_n6332 | 1_n2675;
assign 1_n8394 = ~(1_n7822 ^ 1_n9603);
assign 1_n8350 = 1_n1816 | 1_n10367;
assign 1_n6308 = ~1_n9394;
assign 1_n11630 = 1_n11134 | 1_n816;
assign 1_n5106 = ~(1_n9859 ^ 1_n5830);
assign 1_n12134 = 1_n2330 & 1_n7320;
assign 1_n6867 = ~(1_n3289 ^ 1_n8765);
assign 1_n329 = 1_n10877 | 1_n2675;
assign 1_n5819 = ~(1_n6647 | 1_n6052);
assign 1_n7851 = ~(1_n5273 ^ 1_n8379);
assign 1_n8286 = 1_n12264 | 1_n12355;
assign 1_n13130 = ~(1_n11002 | 1_n3930);
assign 1_n6473 = 1_n4914 & 1_n9624;
assign 1_n2689 = ~1_n2498;
assign 1_n4172 = 1_n5597 & 1_n5846;
assign 1_n12094 = ~(1_n4554 ^ 1_n8927);
assign 1_n9547 = ~(1_n3404 ^ 1_n7704);
assign 1_n4935 = ~(1_n8737 ^ 1_n1244);
assign 1_n11230 = ~1_n8616;
assign 1_n12159 = ~1_n12605;
assign 1_n990 = 1_n6493 & 1_n6517;
assign 1_n9779 = ~(1_n2081 ^ 1_n9681);
assign 1_n10531 = 1_n3393 & 1_n6812;
assign 1_n7365 = ~(1_n1821 ^ 1_n8298);
assign 1_n636 = 1_n7900 | 1_n4640;
assign 1_n13226 = ~1_n10733;
assign 1_n3596 = 1_n7133 | 1_n1043;
assign 1_n3607 = ~(1_n6413 ^ 1_n12562);
assign 1_n360 = ~(1_n10204 | 1_n3876);
assign 1_n7179 = 1_n11801 | 1_n1901;
assign 1_n6736 = ~(1_n5071 ^ 1_n1133);
assign 1_n1742 = 1_n6950 & 1_n10002;
assign 1_n8150 = 1_n9617 & 1_n10359;
assign 1_n6516 = ~(1_n9833 ^ 1_n9544);
assign 1_n221 = ~(1_n10745 ^ 1_n5457);
assign 1_n11007 = ~1_n834;
assign 1_n11246 = ~(1_n3308 ^ 1_n2349);
assign 1_n2746 = 1_n12911 & 1_n2792;
assign 1_n11729 = ~1_n2737;
assign 1_n5928 = ~(1_n4451 ^ 1_n2308);
assign 1_n12963 = 1_n8573 & 1_n6753;
assign 1_n8785 = 1_n11933 | 1_n206;
assign 1_n9739 = ~1_n11734;
assign 1_n10614 = ~(1_n5319 ^ 1_n12005);
assign 1_n12379 = 1_n9848 & 1_n7807;
assign 1_n6236 = 1_n691 | 1_n2941;
assign 1_n11113 = ~1_n12065;
assign 1_n3086 = ~(1_n4874 ^ 1_n7692);
assign 1_n770 = 1_n8905 & 1_n12625;
assign 1_n11964 = ~(1_n12083 | 1_n2478);
assign 1_n11585 = ~(1_n3668 ^ 1_n6560);
assign 1_n8087 = ~(1_n8170 ^ 1_n662);
assign 1_n3287 = 1_n6187 & 1_n4072;
assign 1_n3308 = ~(1_n8025 | 1_n9865);
assign 1_n2519 = ~(1_n7558 ^ 1_n5682);
assign 1_n12625 = ~1_n9903;
assign 1_n11751 = ~1_n8768;
assign 1_n10952 = ~(1_n12440 ^ 1_n1541);
assign 1_n12708 = 1_n9728 | 1_n11555;
assign 1_n10307 = ~(1_n6479 ^ 1_n5315);
assign 1_n6570 = ~(1_n5660 ^ 1_n10562);
assign 1_n9047 = ~(1_n8914 | 1_n7296);
assign 1_n6912 = 1_n11168 | 1_n590;
assign 1_n9314 = ~(1_n2294 | 1_n12228);
assign 1_n7460 = ~1_n8031;
assign 1_n6469 = ~1_n4217;
assign 1_n7760 = 1_n3492 & 1_n8286;
assign 1_n5858 = ~(1_n1534 ^ 1_n3292);
assign 1_n10888 = 1_n5086 | 1_n12814;
assign 1_n9934 = ~1_n11634;
assign 1_n2488 = ~(1_n9571 ^ 1_n12149);
assign 1_n2947 = 1_n10166 | 1_n6497;
assign 1_n2404 = ~1_n1929;
assign 1_n10993 = 1_n154 | 1_n776;
assign 1_n3507 = 1_n4880 | 1_n10659;
assign 1_n10015 = 1_n9353 & 1_n834;
assign 1_n5893 = 1_n8660 | 1_n2938;
assign 1_n3144 = 1_n10392 & 1_n9655;
assign 1_n6317 = 1_n1931 & 1_n4666;
assign 1_n343 = ~1_n504;
assign 1_n718 = ~(1_n2307 | 1_n9258);
assign 1_n10130 = ~(1_n3973 | 1_n11185);
assign 1_n3565 = ~1_n7288;
assign 1_n1177 = ~(1_n9050 ^ 1_n10080);
assign 1_n7869 = 1_n4944 | 1_n12298;
assign 1_n3193 = 1_n9632 | 1_n8268;
assign 1_n4963 = 1_n618 | 1_n9858;
assign 1_n8706 = ~(1_n6072 | 1_n10840);
assign 1_n10076 = ~(1_n12699 ^ 1_n11363);
assign 1_n4896 = 1_n6578 & 1_n6712;
assign 1_n7982 = 1_n4527 & 1_n9067;
assign 1_n448 = ~1_n13003;
assign 1_n5188 = ~(1_n5574 ^ 1_n5764);
assign 1_n12978 = 1_n12283 & 1_n11543;
assign 1_n9423 = ~(1_n10568 | 1_n12520);
assign 1_n2467 = ~(1_n3367 ^ 1_n3938);
assign 1_n1756 = 1_n4129 & 1_n11862;
assign 1_n4149 = ~1_n397;
assign 1_n7841 = ~(1_n498 ^ 1_n9459);
assign 1_n11214 = ~(1_n1942 | 1_n2115);
assign 1_n11050 = ~(1_n7214 ^ 1_n1237);
assign 1_n778 = 1_n13036 | 1_n4640;
assign 1_n3674 = ~1_n3411;
assign 1_n6510 = 1_n7798 | 1_n8268;
assign 1_n11167 = ~(1_n865 | 1_n8055);
assign 1_n7780 = ~1_n10594;
assign 1_n8961 = 1_n3660 | 1_n8958;
assign 1_n4591 = 1_n9313 ^ 1_n764;
assign 1_n8073 = 1_n2913 | 1_n12654;
assign 1_n6010 = ~(1_n12809 | 1_n12066);
assign 1_n6640 = 1_n4625 | 1_n9331;
assign 1_n3620 = 1_n8471 | 1_n6688;
assign 1_n342 = 1_n3163 & 1_n286;
assign 1_n86 = ~(1_n11831 ^ 1_n10647);
assign 1_n426 = ~(1_n4986 ^ 1_n4626);
assign 1_n3246 = ~(1_n624 | 1_n12752);
assign 1_n3074 = ~(1_n9614 ^ 1_n1581);
assign 1_n12145 = ~1_n11335;
assign 1_n12480 = ~(1_n4309 ^ 1_n8999);
assign 1_n997 = 1_n4382 & 1_n1724;
assign 1_n11412 = ~(1_n1096 ^ 1_n5575);
assign 1_n1304 = ~(1_n11917 ^ 1_n1339);
assign 1_n6344 = 1_n10511 & 1_n3360;
assign 1_n12243 = ~1_n9315;
assign 1_n3040 = 1_n6056 | 1_n9492;
assign 1_n1454 = ~(1_n1921 | 1_n933);
assign 1_n2188 = ~(1_n1340 ^ 1_n9840);
assign 1_n6468 = 1_n9228 | 1_n12273;
assign 1_n12089 = 1_n1842 & 1_n6697;
assign 1_n9984 = 1_n9659 & 1_n395;
assign 1_n10640 = 1_n10021 | 1_n2222;
assign 1_n4058 = ~1_n8467;
assign 1_n204 = ~1_n9762;
assign 1_n8085 = 1_n1089 | 1_n8143;
assign 1_n5326 = ~(1_n3571 ^ 1_n3517);
assign 1_n8802 = 1_n63 | 1_n2544;
assign 1_n13107 = ~(1_n13008 | 1_n4637);
assign 1_n12879 = 1_n185 | 1_n4431;
assign 1_n8795 = 1_n7162 & 1_n7769;
assign 1_n6415 = ~(1_n7157 ^ 1_n9742);
assign 1_n3433 = 1_n5188 & 1_n9637;
assign 1_n6171 = ~1_n7829;
assign 1_n7098 = 1_n3643 | 1_n6544;
assign 1_n4173 = 1_n868 | 1_n8269;
assign 1_n4641 = ~(1_n10762 | 1_n1675);
assign 1_n12658 = 1_n2606 | 1_n11422;
assign 1_n11965 = ~1_n5320;
assign 1_n9444 = ~1_n6392;
assign 1_n7934 = 1_n3460 | 1_n6635;
assign 1_n12124 = 1_n7074 | 1_n5242;
assign 1_n11054 = ~1_n4006;
assign 1_n1050 = 1_n13090 | 1_n12415;
assign 1_n3415 = 1_n3142 | 1_n2320;
assign 1_n6503 = 1_n7825 | 1_n10029;
assign 1_n2992 = ~(1_n13056 ^ 1_n3021);
assign 1_n10246 = ~(1_n7712 | 1_n7389);
assign 1_n13151 = ~(1_n2602 ^ 1_n13147);
assign 1_n4804 = 1_n2854 | 1_n2853;
assign 1_n3726 = ~1_n9887;
assign 1_n3831 = 1_n9216 & 1_n5920;
assign 1_n4634 = 1_n8671 | 1_n5796;
assign 1_n12663 = ~1_n8923;
assign 1_n4209 = ~1_n287;
assign 1_n624 = ~(1_n12267 ^ 1_n9495);
assign 1_n12602 = 1_n9061 ^ 1_n5876;
assign 1_n8252 = 1_n6958 | 1_n12360;
assign 1_n5223 = 1_n6634 & 1_n7547;
assign 1_n194 = 1_n1413 & 1_n9398;
assign 1_n6576 = 1_n4814 | 1_n8584;
assign 1_n12937 = ~(1_n5752 ^ 1_n12827);
assign 1_n4392 = 1_n168 & 1_n1245;
assign 1_n12396 = ~(1_n4788 | 1_n8122);
assign 1_n10604 = ~(1_n656 | 1_n9514);
assign 1_n486 = 1_n9653 & 1_n1979;
assign 1_n1370 = ~1_n11734;
assign 1_n12921 = 1_n354 | 1_n12934;
assign 1_n4636 = 1_n809 & 1_n7404;
assign 1_n1939 = ~(1_n10351 ^ 1_n1788);
assign 1_n5687 = 1_n9010 | 1_n121;
assign 1_n7563 = ~(1_n12774 ^ 1_n6228);
assign 1_n5579 = 1_n12124 | 1_n7437;
assign 1_n5116 = ~(1_n2665 ^ 1_n7992);
assign 1_n4615 = ~(1_n4102 ^ 1_n8528);
assign 1_n8104 = 1_n12419 & 1_n790;
assign 1_n6198 = 1_n1191 | 1_n2544;
assign 1_n2426 = ~(1_n4279 ^ 1_n7348);
assign 1_n12558 = 1_n3428 | 1_n4230;
assign 1_n10254 = 1_n5310 & 1_n5630;
assign 1_n2353 = 1_n186 | 1_n7551;
assign 1_n316 = 1_n7529 & 1_n5729;
assign 1_n9133 = 1_n2692 | 1_n5242;
assign 1_n3330 = 1_n13013 | 1_n4454;
assign 1_n4474 = 1_n7973 & 1_n4963;
assign 1_n8578 = ~1_n1423;
assign 1_n3704 = ~(1_n12756 ^ 1_n9408);
assign 1_n12015 = ~(1_n9927 ^ 1_n10493);
assign 1_n8908 = ~(1_n4025 ^ 1_n11886);
assign 1_n5104 = ~(1_n11445 ^ 1_n3055);
assign 1_n6770 = ~1_n10408;
assign 1_n11855 = ~(1_n2831 ^ 1_n5826);
assign 1_n10571 = 1_n11680 | 1_n9195;
assign 1_n3688 = 1_n2630 | 1_n561;
assign 1_n11860 = 1_n289 & 1_n7934;
assign 1_n2634 = 1_n2950 | 1_n5945;
assign 1_n12086 = ~1_n5659;
assign 1_n6327 = ~1_n10105;
assign 1_n6186 = ~1_n9058;
assign 1_n887 = 1_n5731 ^ 1_n2314;
assign 1_n3202 = 1_n7253 & 1_n8531;
assign 1_n9468 = 1_n8575 | 1_n12423;
assign 1_n9424 = 1_n4778 | 1_n11491;
assign 1_n5118 = 1_n10202 | 1_n8226;
assign 1_n3703 = ~1_n10642;
assign 1_n9885 = ~1_n2350;
assign 1_n2926 = ~(1_n383 ^ 1_n3177);
assign 1_n1600 = ~(1_n2812 ^ 1_n3207);
assign 1_n4291 = ~(1_n5365 ^ 1_n4892);
assign 1_n6390 = 1_n636 & 1_n9365;
assign 1_n1575 = 1_n11114 | 1_n1012;
assign 1_n4686 = ~1_n8139;
assign 1_n5486 = ~(1_n1079 ^ 1_n1616);
assign 1_n2950 = 1_n10188 | 1_n2958;
assign 1_n912 = 1_n5430 | 1_n9075;
assign 1_n3526 = 1_n7130 & 1_n5489;
assign 1_n2235 = ~(1_n1543 ^ 1_n426);
assign 1_n11152 = ~1_n2590;
assign 1_n10579 = ~(1_n7635 | 1_n12087);
assign 1_n12445 = 1_n10588 | 1_n9744;
assign 1_n10668 = 1_n10253 | 1_n6703;
assign 1_n5254 = ~(1_n6588 ^ 1_n1115);
assign 1_n8773 = ~(1_n10069 | 1_n5419);
assign 1_n10238 = ~(1_n4837 ^ 1_n8013);
assign 1_n9952 = 1_n9552 & 1_n5608;
assign 1_n7100 = 1_n4377 & 1_n10633;
assign 1_n9393 = ~(1_n4952 | 1_n1133);
assign 1_n7189 = ~(1_n8300 ^ 1_n148);
assign 1_n1479 = ~(1_n891 ^ 1_n2082);
assign 1_n9278 = ~(1_n5879 | 1_n13176);
assign 1_n3597 = 1_n1571 | 1_n1026;
assign 1_n9357 = ~(1_n4306 ^ 1_n4362);
assign 1_n2931 = ~(1_n10984 ^ 1_n9547);
assign 1_n3882 = ~(1_n4035 | 1_n3912);
assign 1_n12646 = 1_n1230 | 1_n9699;
assign 1_n12575 = 1_n5272 & 1_n5194;
assign 1_n7412 = 1_n8472 | 1_n8563;
assign 1_n10297 = ~(1_n11603 ^ 1_n12776);
assign 1_n10535 = ~1_n7479;
assign 1_n8123 = 1_n1912 & 1_n12263;
assign 1_n10667 = 1_n7410 & 1_n8070;
assign 1_n12278 = ~(1_n4233 ^ 1_n8966);
assign 1_n177 = 1_n6210;
assign 1_n6363 = 1_n4221 | 1_n6769;
assign 1_n7135 = ~1_n10594;
assign 1_n12056 = ~(1_n3444 ^ 1_n838);
assign 1_n9162 = ~1_n8332;
assign 1_n4411 = 1_n11701 & 1_n11194;
assign 1_n9456 = ~(1_n382 | 1_n3967);
assign 1_n8808 = 1_n7680 | 1_n12818;
assign 1_n993 = 1_n3195 | 1_n10470;
assign 1_n12669 = ~(1_n11550 ^ 1_n2458);
assign 1_n10080 = ~(1_n1765 ^ 1_n8393);
assign 1_n1381 = ~(1_n10148 | 1_n8232);
assign 1_n3661 = 1_n11080 | 1_n10155;
assign 1_n2340 = ~(1_n10609 ^ 1_n13126);
assign 1_n9403 = 1_n5853 | 1_n5658;
assign 1_n2238 = 1_n7672 | 1_n7221;
assign 1_n6256 = ~(1_n6951 ^ 1_n3018);
assign 1_n9964 = 1_n9700 | 1_n4652;
assign 1_n4573 = 1_n2504 | 1_n2276;
assign 1_n6726 = ~1_n8859;
assign 1_n11937 = 1_n3516 | 1_n559;
assign 1_n8024 = ~1_n1364;
assign 1_n3471 = ~(1_n778 | 1_n10704);
assign 1_n5039 = 1_n11018 | 1_n9159;
assign 1_n9425 = ~(1_n13171 ^ 1_n5555);
assign 1_n205 = ~1_n6484;
assign 1_n1652 = ~1_n2000;
assign 1_n11697 = ~1_n3352;
assign 1_n2225 = 1_n8729 | 1_n9159;
assign 1_n2336 = ~(1_n6191 ^ 1_n1894);
assign 1_n2412 = ~1_n9924;
assign 1_n3194 = ~1_n11709;
assign 1_n11323 = ~1_n13172;
assign 1_n599 = 1_n9676 | 1_n5817;
assign 1_n10184 = 1_n10616 | 1_n11578;
assign 1_n5984 = 1_n4756 & 1_n2901;
assign 1_n4728 = 1_n6260 & 1_n2918;
assign 1_n3088 = ~(1_n11030 ^ 1_n11488);
assign 1_n7437 = ~(1_n6283 ^ 1_n12779);
assign 1_n2053 = 1_n5348 & 1_n6523;
assign 1_n334 = ~1_n401;
assign 1_n2476 = ~(1_n5649 ^ 1_n1685);
assign 1_n11520 = ~(1_n7197 | 1_n4447);
assign 1_n1465 = 1_n10975 & 1_n6352;
assign 1_n5432 = 1_n5988 & 1_n6992;
assign 1_n9809 = ~1_n12276;
assign 1_n12837 = ~1_n12482;
assign 1_n6286 = 1_n10719 & 1_n9454;
assign 1_n2724 = ~(1_n7360 ^ 1_n10818);
assign 1_n8942 = ~(1_n7823 ^ 1_n9875);
assign 1_n481 = 1_n13066 & 1_n4468;
assign 1_n11885 = 1_n6772 & 1_n8574;
assign 1_n6691 = ~(1_n9391 ^ 1_n9057);
assign 1_n10889 = ~(1_n5816 ^ 1_n6642);
assign 1_n6799 = ~(1_n12008 | 1_n1863);
assign 1_n7650 = 1_n10334 | 1_n11668;
assign 1_n8429 = ~(1_n5599 | 1_n6613);
assign 1_n3953 = ~(1_n6114 ^ 1_n4839);
assign 1_n3940 = ~1_n12651;
assign 1_n8328 = ~(1_n12627 ^ 1_n7079);
assign 1_n10387 = ~(1_n259 | 1_n12138);
assign 1_n7949 = 1_n2140 | 1_n620;
assign 1_n1764 = ~(1_n11684 ^ 1_n2309);
assign 1_n1528 = 1_n5214 & 1_n3409;
assign 1_n5935 = ~(1_n3013 ^ 1_n11410);
assign 1_n281 = 1_n9969 | 1_n7732;
assign 1_n5396 = ~(1_n3475 ^ 1_n11932);
assign 1_n9549 = 1_n11646 & 1_n9976;
assign 1_n8034 = 1_n9288 & 1_n10006;
assign 1_n2310 = 1_n2669 | 1_n6635;
assign 1_n9017 = ~1_n11222;
assign 1_n4619 = 1_n12926 | 1_n8341;
assign 1_n6116 = ~(1_n11059 ^ 1_n13091);
assign 1_n3782 = 1_n10241 & 1_n10959;
assign 1_n5605 = ~(1_n6518 ^ 1_n557);
assign 1_n6589 = 1_n5531 & 1_n5602;
assign 1_n5329 = ~(1_n3159 ^ 1_n12507);
assign 1_n3241 = 1_n9465 | 1_n9772;
assign 1_n7252 = 1_n8560 & 1_n6365;
assign 1_n9712 = ~1_n3850;
assign 1_n1544 = ~1_n6570;
assign 1_n11157 = ~1_n7411;
assign 1_n8531 = 1_n5095 | 1_n2205;
assign 1_n9836 = ~(1_n2485 ^ 1_n12752);
assign 1_n11821 = 1_n7446 | 1_n5223;
assign 1_n7636 = ~1_n1384;
assign 1_n3316 = 1_n481 | 1_n10899;
assign 1_n708 = 1_n6238 & 1_n2137;
assign 1_n12424 = 1_n4964 & 1_n2339;
assign 1_n10853 = ~(1_n9965 ^ 1_n10831);
assign 1_n3598 = ~1_n12853;
assign 1_n4369 = ~(1_n11401 ^ 1_n6899);
assign 1_n11241 = 1_n3496 | 1_n6966;
assign 1_n10837 = 1_n7809 | 1_n13232;
assign 1_n5245 = ~1_n11064;
assign 1_n7265 = ~(1_n9530 ^ 1_n13057);
assign 1_n6903 = 1_n4901 & 1_n6403;
assign 1_n7229 = 1_n7608 | 1_n6404;
assign 1_n1581 = ~(1_n9315 ^ 1_n4399);
assign 1_n11171 = ~1_n1916;
assign 1_n8112 = 1_n2942 | 1_n1618;
assign 1_n3036 = ~1_n6075;
assign 1_n7625 = 1_n1490 | 1_n4904;
assign 1_n4658 = 1_n3461 & 1_n6259;
assign 1_n1878 = 1_n7193 | 1_n9933;
assign 1_n7810 = 1_n12476 | 1_n5184;
assign 1_n9270 = 1_n4488 & 1_n3036;
assign 1_n7673 = ~(1_n3368 ^ 1_n7576);
assign 1_n8479 = 1_n8108 | 1_n8702;
assign 1_n5349 = ~(1_n7326 | 1_n3565);
assign 1_n6500 = ~(1_n10423 ^ 1_n3276);
assign 1_n9555 = 1_n8849 | 1_n5414;
assign 1_n6043 = ~(1_n2482 ^ 1_n10113);
assign 1_n7758 = 1_n7133 | 1_n12847;
assign 1_n10733 = 1_n10751 ^ 1_n1032;
assign 1_n6649 = 1_n2017 | 1_n7692;
assign 1_n8725 = ~(1_n11417 ^ 1_n11019);
assign 1_n961 = ~(1_n10811 | 1_n836);
assign 1_n1705 = 1_n2144 | 1_n12421;
assign 1_n11199 = 1_n6308 & 1_n6925;
assign 1_n4747 = ~(1_n2516 ^ 1_n5728);
assign 1_n6430 = 1_n4355 | 1_n8933;
assign 1_n74 = 1_n2724 & 1_n6455;
assign 1_n12283 = ~(1_n10697 ^ 1_n2366);
assign 1_n8898 = ~1_n1812;
assign 1_n8092 = 1_n7450 & 1_n7867;
assign 1_n7315 = 1_n7409 | 1_n2714;
assign 1_n11244 = ~1_n13058;
assign 1_n7030 = ~(1_n3637 ^ 1_n12047);
assign 1_n7224 = 1_n6566 & 1_n155;
assign 1_n3752 = ~1_n2392;
assign 1_n3502 = 1_n4033 & 1_n1503;
assign 1_n5292 = 1_n3250 & 1_n4117;
assign 1_n9477 = 1_n4946 | 1_n4139;
assign 1_n8633 = ~(1_n11970 ^ 1_n2502);
assign 1_n7648 = 1_n9049 & 1_n2827;
assign 1_n5572 = 1_n12563 | 1_n10029;
assign 1_n10205 = ~(1_n28 ^ 1_n253);
assign 1_n2955 = 1_n6624 & 1_n7575;
assign 1_n1413 = 1_n6787 | 1_n4669;
assign 1_n3656 = 1_n3270 | 1_n13143;
assign 1_n10057 = ~1_n5962;
assign 1_n10552 = ~1_n6668;
assign 1_n5704 = 1_n1887 | 1_n1043;
assign 1_n2050 = ~(1_n5798 | 1_n9276);
assign 1_n5643 = ~(1_n4781 ^ 1_n8633);
assign 1_n9421 = ~1_n11574;
assign 1_n11363 = 1_n161 | 1_n10179;
assign 1_n4620 = ~1_n2295;
assign 1_n4705 = ~(1_n5759 ^ 1_n12038);
assign 1_n2584 = ~(1_n2125 ^ 1_n10118);
assign 1_n7169 = ~(1_n11530 | 1_n4472);
assign 1_n9048 = 1_n3545 & 1_n13140;
assign 1_n4219 = 1_n7055 & 1_n6292;
assign 1_n4363 = 1_n994 | 1_n1433;
assign 1_n7808 = ~(1_n6199 ^ 1_n3147);
assign 1_n1758 = ~(1_n4531 ^ 1_n6077);
assign 1_n3686 = ~(1_n12468 | 1_n2202);
assign 1_n9414 = 1_n308 & 1_n4302;
assign 1_n310 = 1_n8392 | 1_n8030;
assign 1_n8919 = 1_n8887 ^ 1_n5270;
assign 1_n6698 = ~(1_n1549 ^ 1_n12611);
assign 1_n12563 = ~1_n12306;
assign 1_n2337 = 1_n8335 | 1_n6265;
assign 1_n1377 = ~1_n10424;
assign 1_n8903 = 1_n12776 & 1_n11603;
assign 1_n13119 = 1_n318 | 1_n10106;
assign 1_n9723 = ~1_n7659;
assign 1_n10225 = 1_n9112 | 1_n4947;
assign 1_n4045 = 1_n1995 | 1_n1081;
assign 1_n2073 = ~(1_n9389 ^ 1_n9551);
assign 1_n7950 = ~1_n9915;
assign 1_n8121 = ~(1_n9436 ^ 1_n3674);
assign 1_n11970 = ~(1_n494 ^ 1_n11329);
assign 1_n7838 = ~(1_n7294 ^ 1_n10111);
assign 1_n2828 = ~(1_n10424 ^ 1_n13076);
assign 1_n11800 = ~1_n3838;
assign 1_n5061 = 1_n7523 & 1_n7975;
assign 1_n1186 = ~1_n8227;
assign 1_n1725 = ~1_n6409;
assign 1_n12137 = 1_n7372 | 1_n11628;
assign 1_n6908 = ~(1_n1313 ^ 1_n3667);
assign 1_n5732 = 1_n7529 & 1_n10451;
assign 1_n5160 = 1_n7283 | 1_n7723;
assign 1_n10040 = 1_n3987 & 1_n12362;
assign 1_n3871 = 1_n6975 | 1_n7871;
assign 1_n160 = 1_n9934 | 1_n2675;
assign 1_n9247 = 1_n2715 & 1_n4265;
assign 1_n5024 = 1_n4729 & 1_n3204;
assign 1_n1255 = ~1_n2202;
assign 1_n7781 = ~(1_n4337 ^ 1_n10478);
assign 1_n7958 = ~(1_n12716 ^ 1_n9322);
assign 1_n4302 = ~(1_n1849 ^ 1_n5594);
assign 1_n10506 = ~(1_n3741 ^ 1_n9143);
assign 1_n3589 = ~1_n589;
assign 1_n6094 = ~(1_n11561 ^ 1_n8578);
assign 1_n1519 = ~(1_n4356 ^ 1_n10499);
assign 1_n6855 = 1_n8400 | 1_n13148;
assign 1_n930 = ~1_n12577;
assign 1_n2610 = 1_n9945 | 1_n2418;
assign 1_n9937 = 1_n9892 | 1_n10526;
assign 1_n12030 = 1_n3259 | 1_n80;
assign 1_n9465 = ~1_n4507;
assign 1_n1045 = ~1_n12443;
assign 1_n5756 = ~(1_n10341 ^ 1_n3636);
assign 1_n3516 = ~1_n3311;
assign 1_n11916 = ~(1_n3728 | 1_n8537);
assign 1_n8250 = 1_n12055 | 1_n1285;
assign 1_n8763 = 1_n12737 & 1_n5956;
assign 1_n8658 = ~1_n13184;
assign 1_n2406 = ~1_n2458;
assign 1_n6543 = ~1_n12641;
assign 1_n4561 = 1_n7924 & 1_n2528;
assign 1_n4941 = 1_n2412 & 1_n5668;
assign 1_n5303 = 1_n6690 & 1_n12772;
assign 1_n7613 = ~(1_n2514 ^ 1_n13160);
assign 1_n4738 = 1_n74 | 1_n9278;
assign 1_n12916 = 1_n424 ^ 1_n1698;
assign 1_n2509 = 1_n8008 | 1_n12113;
assign 1_n396 = ~(1_n9292 ^ 1_n11921);
assign 1_n3055 = ~(1_n6446 ^ 1_n4178);
assign 1_n52 = 1_n6849 | 1_n12526;
assign 1_n456 = ~(1_n1546 ^ 1_n2204);
assign 1_n11808 = ~1_n11324;
assign 1_n8826 = 1_n2648 & 1_n9829;
assign 1_n7192 = 1_n5040 | 1_n6370;
assign 1_n3884 = ~(1_n1676 | 1_n10083);
assign 1_n7855 = 1_n4595 & 1_n11343;
assign 1_n1515 = 1_n12139 & 1_n11775;
assign 1_n2937 = ~(1_n4175 ^ 1_n3231);
assign 1_n197 = 1_n10290 | 1_n11668;
assign 1_n5815 = 1_n8093 & 1_n7019;
assign 1_n10600 = ~(1_n145 | 1_n853);
assign 1_n11265 = ~(1_n12642 | 1_n3291);
assign 1_n8287 = ~(1_n4713 ^ 1_n11441);
assign 1_n13178 = 1_n11626 | 1_n2891;
assign 1_n3219 = ~(1_n11488 | 1_n1982);
assign 1_n3997 = 1_n724 & 1_n11163;
assign 1_n8195 = ~(1_n7874 ^ 1_n5922);
assign 1_n8484 = ~(1_n12610 ^ 1_n13067);
assign 1_n367 = ~(1_n5556 | 1_n13198);
assign 1_n9918 = 1_n1320 | 1_n2671;
assign 1_n5365 = 1_n5423 | 1_n2133;
assign 1_n12058 = 1_n4622 | 1_n11214;
assign 1_n6595 = ~1_n13060;
assign 1_n2177 = 1_n1883 | 1_n6732;
assign 1_n8560 = 1_n1522 & 1_n3483;
assign 1_n2922 = 1_n6035 | 1_n11146;
assign 1_n747 = 1_n626 | 1_n7887;
assign 1_n2813 = ~(1_n1256 ^ 1_n1619);
assign 1_n3973 = 1_n2198 & 1_n193;
assign 1_n11712 = 1_n11690 & 1_n12743;
assign 1_n2439 = ~(1_n1803 ^ 1_n7587);
assign 1_n8901 = 1_n11320 | 1_n6293;
assign 1_n2335 = 1_n2747 & 1_n8762;
assign 1_n3863 = ~(1_n9371 ^ 1_n8323);
assign 1_n3251 = 1_n9828 & 1_n10804;
assign 1_n5221 = ~(1_n4968 | 1_n11700);
assign 1_n11603 = ~(1_n2513 ^ 1_n11578);
assign 1_n13020 = ~(1_n3878 ^ 1_n7248);
assign 1_n10217 = ~(1_n5407 ^ 1_n2708);
assign 1_n1144 = 1_n8569;
assign 1_n449 = ~(1_n3764 | 1_n2888);
assign 1_n12587 = ~(1_n232 | 1_n3580);
assign 1_n6240 = 1_n683 | 1_n4144;
assign 1_n7148 = ~(1_n13193 ^ 1_n2642);
assign 1_n12530 = 1_n154 | 1_n9962;
assign 1_n7121 = ~(1_n6184 ^ 1_n2115);
assign 1_n11986 = ~1_n12417;
assign 1_n9242 = 1_n1582 & 1_n5706;
assign 1_n9535 = 1_n660 | 1_n1530;
assign 1_n1141 = ~(1_n880 ^ 1_n2856);
assign 1_n6809 = ~(1_n11518 ^ 1_n10337);
assign 1_n441 = ~(1_n12737 ^ 1_n10009);
assign 1_n8699 = 1_n6726 | 1_n206;
assign 1_n7174 = 1_n9094 | 1_n6605;
assign 1_n8921 = ~(1_n565 ^ 1_n10445);
assign 1_n10362 = 1_n1539 & 1_n12633;
assign 1_n13062 = 1_n1296 | 1_n8702;
assign 1_n3904 = ~(1_n1461 ^ 1_n2303);
assign 1_n5834 = 1_n2482 & 1_n12289;
assign 1_n1337 = ~1_n11254;
assign 1_n3080 = ~(1_n6805 | 1_n7691);
assign 1_n10270 = ~(1_n1744 | 1_n315);
assign 1_n6984 = ~(1_n10134 ^ 1_n183);
assign 1_n2329 = ~1_n7974;
assign 1_n3767 = 1_n11291 | 1_n7530;
assign 1_n1326 = 1_n3473 & 1_n8337;
assign 1_n1287 = ~(1_n5402 | 1_n5149);
assign 1_n11877 = 1_n10263 | 1_n12695;
assign 1_n12712 = 1_n5365 | 1_n8749;
assign 1_n1538 = ~1_n12418;
assign 1_n8127 = 1_n5667 | 1_n5242;
assign 1_n2118 = ~1_n12408;
assign 1_n13143 = ~(1_n10409 ^ 1_n741);
assign 1_n8047 = 1_n9450 | 1_n6968;
assign 1_n9092 = 1_n2458 & 1_n9669;
assign 1_n9208 = ~(1_n5702 | 1_n7866);
assign 1_n5697 = ~1_n13098;
assign 1_n3870 = ~1_n825;
assign 1_n1741 = ~1_n10606;
assign 1_n2204 = 1_n7158 | 1_n2059;
assign 1_n8863 = ~1_n3409;
assign 1_n10004 = 1_n4964 & 1_n11222;
assign 1_n10971 = ~(1_n12812 ^ 1_n2983);
assign 1_n10191 = 1_n545 & 1_n1849;
assign 1_n5237 = 1_n5118 & 1_n6806;
assign 1_n2120 = ~(1_n2807 ^ 1_n10355);
assign 1_n11843 = ~(1_n11673 | 1_n42);
assign 1_n1987 = 1_n7869 & 1_n3606;
assign 1_n3310 = 1_n10871 | 1_n1463;
assign 1_n6178 = ~1_n11537;
assign 1_n4427 = 1_n4708 & 1_n12550;
assign 1_n394 = 1_n12902 & 1_n1684;
assign 1_n4001 = 1_n433 & 1_n9224;
assign 1_n2665 = ~(1_n10483 ^ 1_n6782);
assign 1_n7680 = 1_n10143 | 1_n12847;
assign 1_n336 = 1_n93 & 1_n7772;
assign 1_n11439 = 1_n6164 & 1_n413;
assign 1_n12760 = 1_n1030 & 1_n4243;
assign 1_n5366 = 1_n5926 | 1_n10884;
assign 1_n12341 = 1_n11985 & 1_n5435;
assign 1_n13111 = ~(1_n6179 | 1_n5674);
assign 1_n8292 = 1_n11548 | 1_n9159;
assign 1_n11795 = 1_n6010 | 1_n11746;
assign 1_n5262 = 1_n9646 & 1_n12984;
assign 1_n10663 = ~(1_n10053 ^ 1_n12087);
assign 1_n8678 = ~(1_n5114 ^ 1_n3506);
assign 1_n9995 = 1_n6498 | 1_n258;
assign 1_n4648 = 1_n10290 | 1_n6265;
assign 1_n5951 = ~(1_n5935 ^ 1_n8181);
assign 1_n54 = ~(1_n5438 ^ 1_n5070);
assign 1_n4903 = 1_n12397 | 1_n5235;
assign 1_n703 = 1_n10990 | 1_n13032;
assign 1_n12215 = ~(1_n3296 ^ 1_n5458);
assign 1_n13150 = ~(1_n10163 | 1_n4344);
assign 1_n13121 = 1_n855 & 1_n2047;
assign 1_n11652 = 1_n8940 & 1_n5536;
assign 1_n10384 = ~1_n9895;
assign 1_n9282 = ~1_n8139;
assign 1_n5650 = ~1_n5302;
assign 1_n10515 = ~(1_n149 | 1_n8152);
assign 1_n10703 = 1_n5270 & 1_n5383;
assign 1_n7144 = 1_n4848 & 1_n4984;
assign 1_n3450 = ~1_n6700;
assign 1_n4799 = 1_n4114 & 1_n8506;
assign 1_n8907 = ~1_n9610;
assign 1_n2583 = 1_n12592 & 1_n3085;
assign 1_n9090 = ~(1_n2630 ^ 1_n2561);
assign 1_n13019 = ~(1_n10048 | 1_n12842);
assign 1_n7761 = 1_n8183 & 1_n9475;
assign 1_n1917 = 1_n3998 & 1_n4486;
assign 1_n7561 = 1_n4411 | 1_n11135;
assign 1_n969 = ~(1_n3263 | 1_n12045);
assign 1_n529 = ~(1_n4264 ^ 1_n6287);
assign 1_n132 = 1_n9567 | 1_n7429;
assign 1_n7074 = ~1_n469;
assign 1_n4929 = 1_n9553 | 1_n6278;
assign 1_n444 = ~(1_n11433 ^ 1_n12214);
assign 1_n12490 = ~1_n9475;
assign 1_n7520 = ~(1_n6800 | 1_n13236);
assign 1_n2614 = ~1_n1302;
assign 1_n4976 = 1_n9181 | 1_n5740;
assign 1_n7012 = 1_n5890 | 1_n2133;
assign 1_n3491 = ~(1_n13094 | 1_n8218);
assign 1_n13040 = 1_n4618 & 1_n1232;
assign 1_n6080 = 1_n6421 & 1_n13088;
assign 1_n4412 = ~1_n1753;
assign 1_n12788 = 1_n12855 | 1_n9088;
assign 1_n4321 = 1_n2877 | 1_n7903;
assign 1_n4047 = 1_n3342 & 1_n8606;
assign 1_n6488 = ~1_n3076;
assign 1_n10990 = ~(1_n2431 | 1_n10178);
assign 1_n972 = 1_n12043 & 1_n1005;
assign 1_n8244 = 1_n189 | 1_n11929;
assign 1_n5210 = 1_n1331 | 1_n4455;
assign 1_n5211 = ~(1_n4021 ^ 1_n6863);
assign 1_n3172 = 1_n11582 | 1_n3801;
assign 1_n10651 = 1_n233 & 1_n11539;
assign 1_n4011 = ~(1_n7277 ^ 1_n5378);
assign 1_n4942 = 1_n5377 | 1_n12491;
assign 1_n6288 = ~(1_n1092 ^ 1_n1479);
assign 1_n4601 = ~(1_n10802 ^ 1_n10684);
assign 1_n1933 = 1_n8532 | 1_n12273;
assign 1_n185 = ~(1_n6264 | 1_n11458);
assign 1_n12111 = ~(1_n2063 | 1_n12586);
assign 1_n4784 = 1_n2130 | 1_n8465;
assign 1_n2802 = 1_n6768 | 1_n9195;
assign 1_n3444 = 1_n7228 | 1_n1383;
assign 1_n8364 = ~(1_n6765 | 1_n10744);
assign 1_n378 = ~(1_n12374 ^ 1_n12322);
assign 1_n7399 = ~(1_n11763 ^ 1_n8021);
assign 1_n7388 = ~1_n6417;
assign 1_n10417 = 1_n10708 & 1_n9588;
assign 1_n9606 = ~1_n4748;
assign 1_n8513 = ~(1_n6902 | 1_n9158);
assign 1_n7817 = ~1_n720;
assign 1_n6335 = 1_n5897 | 1_n159;
assign 1_n1082 = ~1_n12564;
assign 1_n5392 = ~(1_n2334 | 1_n3468);
assign 1_n4139 = ~1_n5753;
assign 1_n6785 = ~(1_n3951 ^ 1_n5896);
assign 1_n12319 = ~(1_n4369 ^ 1_n9805);
assign 1_n9992 = ~1_n1521;
assign 1_n6846 = ~1_n12482;
assign 1_n3284 = 1_n10761 | 1_n12388;
assign 1_n3890 = ~1_n9620;
assign 1_n10308 = ~(1_n12230 | 1_n4204);
assign 1_n6146 = 1_n1359 | 1_n2438;
assign 1_n9792 = ~(1_n2011 ^ 1_n9483);
assign 1_n4386 = ~(1_n6097 | 1_n11416);
assign 1_n11454 = ~(1_n10500 ^ 1_n6542);
assign 1_n505 = 1_n5107 | 1_n1571;
assign 1_n2631 = 1_n7011 & 1_n7117;
assign 1_n10916 = ~1_n3395;
assign 1_n12478 = ~1_n4318;
assign 1_n7240 = 1_n10948 & 1_n9137;
assign 1_n9081 = ~(1_n6242 ^ 1_n10276);
assign 1_n7075 = ~1_n6168;
assign 1_n5212 = 1_n3159 | 1_n9507;
assign 1_n9892 = 1_n12748 | 1_n12188;
assign 1_n3750 = 1_n6172 | 1_n7610;
assign 1_n11122 = ~1_n7720;
assign 1_n10073 = ~(1_n5299 ^ 1_n13072);
assign 1_n9115 = 1_n3435 & 1_n11697;
assign 1_n13139 = 1_n8835 & 1_n8521;
assign 1_n978 = 1_n652 | 1_n5076;
assign 1_n8936 = ~1_n28;
assign 1_n363 = ~(1_n1675 ^ 1_n4573);
assign 1_n13011 = 1_n6590 | 1_n1985;
assign 1_n7547 = 1_n6509 | 1_n9590;
assign 1_n9199 = 1_n4736 & 1_n5256;
assign 1_n9240 = 1_n9489 | 1_n5242;
assign 1_n4057 = ~(1_n4840 | 1_n5887);
assign 1_n10172 = 1_n4495 | 1_n8499;
assign 1_n11583 = 1_n8026 & 1_n9623;
assign 1_n9818 = ~(1_n11599 ^ 1_n8226);
assign 1_n13052 = ~1_n5965;
assign 1_n2098 = 1_n7418 | 1_n11744;
assign 1_n6630 = ~1_n497;
assign 1_n8983 = 1_n4164 & 1_n5441;
assign 1_n5974 = ~1_n9212;
assign 1_n10155 = 1_n12552 | 1_n8030;
assign 1_n4883 = 1_n5370 | 1_n5983;
assign 1_n5993 = 1_n8646 | 1_n177;
assign 1_n9910 = ~1_n7671;
assign 1_n7452 = 1_n6533 & 1_n427;
assign 1_n5522 = ~1_n7919;
assign 1_n5358 = ~(1_n6254 ^ 1_n4367);
assign 1_n3693 = ~(1_n3770 ^ 1_n10758);
assign 1_n11895 = ~(1_n9578 ^ 1_n213);
assign 1_n10146 = 1_n10388 & 1_n10700;
assign 1_n3063 = ~1_n5576;
assign 1_n3987 = 1_n11596 & 1_n11721;
assign 1_n5346 = 1_n6943 & 1_n3637;
assign 1_n8660 = 1_n5776 & 1_n924;
assign 1_n1614 = ~(1_n2379 | 1_n690);
assign 1_n7516 = ~(1_n3138 ^ 1_n7058);
assign 1_n7872 = ~1_n11109;
assign 1_n10882 = ~1_n4528;
assign 1_n3579 = 1_n3564 | 1_n10871;
assign 1_n10288 = 1_n6194 & 1_n2721;
assign 1_n3984 = 1_n2889 | 1_n10319;
assign 1_n2663 = 1_n9695 | 1_n8305;
assign 1_n12859 = ~1_n12670;
assign 1_n7885 = 1_n11878 & 1_n7390;
assign 1_n3295 = ~(1_n5742 | 1_n12170);
assign 1_n3357 = ~(1_n7751 ^ 1_n750);
assign 1_n10446 = 1_n9017 | 1_n8534;
assign 1_n1072 = 1_n8131 | 1_n1985;
assign 1_n4189 = 1_n11033 | 1_n2126;
assign 1_n4714 = ~1_n2856;
assign 1_n6036 = 1_n8248 & 1_n7155;
assign 1_n2374 = ~(1_n7496 ^ 1_n9981);
assign 1_n844 = 1_n1715 | 1_n8313;
assign 1_n9272 = ~1_n10063;
assign 1_n1138 = 1_n10142 & 1_n13058;
assign 1_n1051 = ~1_n7113;
assign 1_n4358 = 1_n5592 & 1_n4607;
assign 1_n12037 = 1_n10410 | 1_n4073;
assign 1_n6251 = ~(1_n3145 ^ 1_n1583);
assign 1_n9014 = 1_n10943 & 1_n6511;
assign 1_n8396 = 1_n6129 | 1_n4947;
assign 1_n2873 = ~(1_n5926 ^ 1_n10884);
assign 1_n3257 = ~1_n194;
assign 1_n4808 = ~1_n4335;
assign 1_n812 = ~1_n3431;
assign 1_n9585 = 1_n7772 & 1_n7411;
assign 1_n12709 = 1_n6605 & 1_n9094;
assign 1_n12775 = 1_n10421 | 1_n12388;
assign 1_n87 = ~(1_n2658 ^ 1_n10396);
assign 1_n2674 = ~1_n5998;
assign 1_n6577 = 1_n9691 & 1_n217;
assign 1_n1003 = 1_n5097 & 1_n8002;
assign 1_n4876 = 1_n3301 | 1_n1415;
assign 1_n12313 = ~(1_n11560 ^ 1_n10646);
assign 1_n3849 = ~(1_n4252 ^ 1_n12666);
assign 1_n10794 = ~1_n13087;
assign 1_n8444 = 1_n5720 | 1_n8502;
assign 1_n10189 = 1_n6148 | 1_n11494;
assign 1_n3184 = 1_n2528 | 1_n7924;
assign 1_n8760 = 1_n11123;
assign 1_n5654 = ~1_n8308;
assign 1_n5032 = ~(1_n589 ^ 1_n7217);
assign 1_n6480 = 1_n5266 | 1_n3380;
assign 1_n8728 = ~1_n1495;
assign 1_n7655 = 1_n6480 & 1_n6835;
assign 1_n12990 = 1_n3225 | 1_n7530;
assign 1_n1409 = ~(1_n4760 ^ 1_n12516);
assign 1_n9285 = 1_n8389 & 1_n7192;
assign 1_n3198 = ~(1_n4042 ^ 1_n2271);
assign 1_n7124 = ~(1_n2458 | 1_n8230);
assign 1_n7473 = ~1_n8357;
assign 1_n8184 = ~(1_n6961 ^ 1_n1527);
assign 1_n11410 = ~(1_n5353 ^ 1_n4456);
assign 1_n5514 = 1_n7234 | 1_n12718;
assign 1_n9312 = ~(1_n9883 ^ 1_n8404);
assign 1_n13154 = ~1_n287;
assign 1_n11298 = ~(1_n12816 ^ 1_n8037);
assign 1_n2149 = 1_n10908 & 1_n6937;
assign 1_n11963 = 1_n3503 & 1_n11070;
assign 1_n11529 = ~(1_n3593 ^ 1_n1455);
assign 1_n4881 = 1_n11235 & 1_n6113;
assign 1_n8154 = 1_n10158 | 1_n1583;
assign 1_n8509 = 1_n6119 & 1_n4432;
assign 1_n9932 = ~(1_n9407 ^ 1_n1933);
assign 1_n12806 = 1_n7532 | 1_n4724;
assign 1_n9853 = 1_n6215 | 1_n4453;
assign 1_n5150 = 1_n8030 | 1_n4640;
assign 1_n842 = 1_n1163 | 1_n3920;
assign 1_n2525 = ~(1_n8996 ^ 1_n6592);
assign 1_n8997 = 1_n10014 & 1_n8235;
assign 1_n8766 = 1_n12469 | 1_n8534;
assign 1_n8610 = 1_n3730 | 1_n12302;
assign 1_n11082 = ~(1_n10850 | 1_n1486);
assign 1_n3820 = 1_n3956 & 1_n13123;
assign 1_n1521 = ~1_n2690;
assign 1_n12232 = ~(1_n8074 ^ 1_n9615);
assign 1_n12909 = 1_n4771 & 1_n12332;
assign 1_n11026 = 1_n3719 & 1_n9958;
assign 1_n7534 = ~(1_n4842 ^ 1_n858);
assign 1_n2595 = 1_n2220 ^ 1_n2198;
assign 1_n11204 = 1_n4187 & 1_n10512;
assign 1_n289 = 1_n7927 & 1_n7456;
assign 1_n11176 = 1_n12227 & 1_n11286;
assign 1_n7518 = 1_n8583 | 1_n11524;
assign 1_n11924 = 1_n6112 | 1_n12623;
assign 1_n3137 = ~(1_n3283 ^ 1_n4281);
assign 1_n9132 = ~1_n7115;
assign 1_n8018 = ~(1_n8297 | 1_n13055);
assign 1_n5516 = 1_n1939 | 1_n8116;
assign 1_n1628 = 1_n7516 & 1_n1236;
assign 1_n615 = 1_n6875 | 1_n12847;
assign 1_n8388 = 1_n3344 | 1_n8609;
assign 1_n12865 = ~(1_n6424 ^ 1_n6884);
assign 1_n5135 = 1_n6175 | 1_n1192;
assign 1_n9857 = ~(1_n3255 ^ 1_n12672);
assign 1_n1959 = 1_n1215 | 1_n8511;
assign 1_n3243 = ~1_n11396;
assign 1_n11399 = 1_n3636 | 1_n10341;
assign 1_n11567 = 1_n12990 ^ 1_n1024;
assign 1_n3796 = ~(1_n4334 ^ 1_n12958);
assign 1_n521 = ~1_n11873;
assign 1_n963 = ~1_n6611;
assign 1_n3827 = 1_n12512 | 1_n10249;
assign 1_n10450 = ~(1_n2282 ^ 1_n5940);
assign 1_n1213 = 1_n12604 | 1_n2449;
assign 1_n8608 = ~(1_n7199 ^ 1_n10924);
assign 1_n6944 = ~1_n834;
assign 1_n5431 = ~(1_n9993 ^ 1_n6275);
assign 1_n413 = ~1_n3623;
assign 1_n6524 = ~1_n7417;
assign 1_n1339 = ~(1_n810 ^ 1_n8138);
assign 1_n61 = ~1_n11091;
assign 1_n1537 = ~(1_n12530 ^ 1_n797);
assign 1_n9990 = ~(1_n6614 ^ 1_n6996);
assign 1_n5200 = ~1_n12589;
assign 1_n3634 = ~1_n8860;
assign 1_n7200 = ~(1_n82 | 1_n2481);
assign 1_n12236 = 1_n7234 | 1_n206;
assign 1_n8426 = 1_n11729 | 1_n5797;
assign 1_n9532 = ~(1_n10704 ^ 1_n778);
assign 1_n11034 = ~(1_n9826 | 1_n8261);
assign 1_n9055 = ~1_n11089;
assign 1_n5648 = ~(1_n6534 | 1_n3474);
assign 1_n4193 = 1_n7322 & 1_n730;
assign 1_n2872 = ~1_n9531;
assign 1_n4198 = ~1_n3769;
assign 1_n3624 = ~(1_n8311 ^ 1_n6836);
assign 1_n4749 = 1_n8665 | 1_n12655;
assign 1_n12333 = 1_n11157 | 1_n8030;
assign 1_n2797 = ~(1_n973 ^ 1_n2281);
assign 1_n59 = 1_n3531 | 1_n4230;
assign 1_n9719 = ~(1_n8429 ^ 1_n11443);
assign 1_n11316 = 1_n10215 & 1_n5929;
assign 1_n2899 = ~1_n817;
assign 1_n5709 = ~1_n11974;
assign 1_n9567 = 1_n2129 | 1_n4373;
assign 1_n4371 = ~1_n7128;
assign 1_n3422 = 1_n1496 & 1_n5844;
assign 1_n10301 = 1_n12166 | 1_n1197;
assign 1_n11980 = 1_n10931 & 1_n1903;
assign 1_n3557 = 1_n8362 | 1_n6181;
assign 1_n2494 = ~(1_n8004 ^ 1_n2981);
assign 1_n4906 = 1_n3507 & 1_n5717;
assign 1_n53 = ~1_n761;
assign 1_n2299 = 1_n7129 | 1_n2617;
assign 1_n3303 = 1_n10770 & 1_n287;
assign 1_n10190 = 1_n333 | 1_n12967;
assign 1_n8529 = ~1_n5969;
assign 1_n4130 = ~(1_n5934 ^ 1_n12002);
assign 1_n11188 = 1_n10849 & 1_n7784;
assign 1_n9059 = 1_n5947 | 1_n12695;
assign 1_n1410 = 1_n10642 & 1_n7720;
assign 1_n8268 = 1_n765;
assign 1_n6354 = 1_n7608 | 1_n206;
assign 1_n2230 = ~(1_n12141 ^ 1_n12407);
assign 1_n6362 = 1_n4349 ^ 1_n2419;
assign 1_n3250 = ~(1_n1121 ^ 1_n12125);
assign 1_n1767 = ~1_n12950;
assign 1_n9235 = ~(1_n12237 | 1_n2512);
assign 1_n6264 = ~1_n2754;
assign 1_n4836 = 1_n7719 | 1_n275;
assign 1_n6325 = 1_n13201 & 1_n3085;
assign 1_n6842 = ~(1_n4684 | 1_n12927);
assign 1_n8653 = 1_n11103 | 1_n5388;
assign 1_n6207 = ~(1_n8773 | 1_n4345);
assign 1_n745 = 1_n5569 | 1_n7221;
assign 1_n6729 = 1_n3517 & 1_n3571;
assign 1_n7703 = 1_n12416 | 1_n9159;
assign 1_n13115 = 1_n11450 | 1_n4757;
assign 1_n5865 = ~1_n11835;
assign 1_n4951 = ~(1_n5793 ^ 1_n1990);
assign 1_n9772 = ~1_n1342;
assign 1_n2324 = 1_n10565 & 1_n5585;
assign 1_n810 = 1_n12671 | 1_n10430;
assign 1_n7488 = ~(1_n11883 | 1_n9598);
assign 1_n2056 = ~1_n5451;
assign 1_n11055 = 1_n379 | 1_n2816;
assign 1_n928 = 1_n4052 & 1_n109;
assign 1_n1563 = ~(1_n4509 ^ 1_n875);
assign 1_n7546 = 1_n6680 | 1_n2890;
assign 1_n1593 = 1_n8011 | 1_n2772;
assign 1_n7034 = ~(1_n94 ^ 1_n6935);
assign 1_n10518 = ~(1_n10671 ^ 1_n1317);
assign 1_n8866 = 1_n13013 | 1_n0;
assign 1_n7874 = 1_n3826 | 1_n10106;
assign 1_n1073 = ~1_n7749;
assign 1_n11219 = 1_n5113 & 1_n9133;
assign 1_n5757 = ~(1_n1077 ^ 1_n11598);
assign 1_n8979 = 1_n2484 | 1_n10552;
assign 1_n9053 = 1_n2391 | 1_n2531;
assign 1_n6971 = 1_n1107 & 1_n10571;
assign 1_n12539 = 1_n8153 & 1_n11275;
assign 1_n11668 = 1_n9280;
assign 1_n238 = 1_n1206 | 1_n11490;
assign 1_n1879 = 1_n8665 | 1_n1720;
assign 1_n6945 = 1_n3796 | 1_n12724;
assign 1_n2812 = 1_n9098 | 1_n6002;
assign 1_n7724 = ~(1_n1338 ^ 1_n4471);
assign 1_n173 = ~1_n10906;
assign 1_n10039 = ~1_n7144;
assign 1_n4078 = 1_n12348 & 1_n5065;
assign 1_n4533 = 1_n10078 & 1_n11040;
assign 1_n2350 = ~1_n10301;
assign 1_n4829 = 1_n12951 | 1_n7988;
assign 1_n4885 = 1_n9882 | 1_n11300;
assign 1_n12183 = ~1_n6242;
assign 1_n4354 = 1_n3982 & 1_n752;
assign 1_n7072 = ~1_n4399;
assign 1_n148 = ~(1_n10377 ^ 1_n3608);
assign 1_n10350 = 1_n5516 & 1_n6976;
assign 1_n5097 = ~1_n7605;
assign 1_n2827 = 1_n767 & 1_n3832;
assign 1_n1806 = ~(1_n10455 ^ 1_n1147);
assign 1_n5487 = ~(1_n4558 ^ 1_n1811);
assign 1_n5656 = 1_n5530 & 1_n1068;
assign 1_n10612 = ~(1_n5391 | 1_n9231);
assign 1_n1018 = ~1_n9313;
assign 1_n5003 = ~(1_n953 ^ 1_n8746);
assign 1_n12692 = ~(1_n3607 ^ 1_n2525);
assign 1_n1749 = 1_n6913 | 1_n9650;
assign 1_n208 = 1_n11980 | 1_n8375;
assign 1_n490 = ~1_n2869;
assign 1_n7106 = 1_n8766 | 1_n2647;
assign 1_n9105 = ~(1_n1141 ^ 1_n10521);
assign 1_n7515 = 1_n3613 ^ 1_n12527;
assign 1_n6112 = ~1_n8332;
assign 1_n873 = 1_n4173 & 1_n7275;
assign 1_n4817 = ~(1_n3502 | 1_n3857);
assign 1_n4467 = 1_n3208 | 1_n7221;
assign 1_n2126 = 1_n4659 & 1_n3151;
assign 1_n12792 = 1_n3818 | 1_n12040;
assign 1_n9611 = 1_n2008 & 1_n12318;
assign 1_n11284 = ~1_n11222;
assign 1_n3899 = ~(1_n4568 ^ 1_n2693);
assign 1_n2887 = 1_n1416 | 1_n4967;
assign 1_n7519 = 1_n4478 | 1_n1599;
assign 1_n2424 = 1_n6769 | 1_n7935;
assign 1_n3619 = ~1_n12661;
assign 1_n10277 = 1_n2424 | 1_n6729;
assign 1_n9558 = ~1_n12750;
assign 1_n9173 = ~(1_n9200 | 1_n5471);
assign 1_n6719 = 1_n12607 | 1_n8041;
assign 1_n11161 = ~(1_n7375 | 1_n10819);
assign 1_n9946 = ~(1_n1871 ^ 1_n10868);
assign 1_n2644 = 1_n6488 | 1_n6265;
assign 1_n1022 = 1_n10318 ^ 1_n11196;
assign 1_n1679 = 1_n10966 | 1_n9075;
assign 1_n9042 = 1_n9575 | 1_n1500;
assign 1_n657 = ~1_n2841;
assign 1_n1 = 1_n8430 & 1_n10255;
assign 1_n4177 = ~(1_n6292 ^ 1_n10418);
assign 1_n8635 = ~(1_n12815 ^ 1_n3799);
assign 1_n2375 = 1_n1759 & 1_n11382;
assign 1_n4798 = 1_n9239 & 1_n487;
assign 1_n11112 = ~(1_n2144 ^ 1_n11001);
assign 1_n12210 = 1_n6129 | 1_n11144;
assign 1_n7016 = 1_n3444 & 1_n7652;
assign 1_n3058 = ~1_n2482;
assign 1_n9662 = 1_n8992 | 1_n541;
assign 1_n6154 = ~(1_n1540 ^ 1_n6221);
assign 1_n5133 = 1_n5842 | 1_n6033;
assign 1_n3869 = 1_n12465 | 1_n13086;
assign 1_n11090 = ~(1_n12791 ^ 1_n6666);
assign 1_n3872 = ~(1_n570 | 1_n3366);
assign 1_n6950 = 1_n103 & 1_n854;
assign 1_n5186 = 1_n7622 & 1_n8815;
assign 1_n10674 = 1_n4844 | 1_n9075;
assign 1_n5136 = ~1_n7214;
assign 1_n12504 = 1_n6476 | 1_n8663;
assign 1_n11681 = 1_n9417 & 1_n256;
assign 1_n11036 = ~(1_n8109 ^ 1_n3515);
assign 1_n6261 = ~(1_n2203 ^ 1_n7623);
assign 1_n3306 = ~(1_n11775 ^ 1_n665);
assign 1_n10938 = 1_n227 | 1_n6635;
assign 1_n12824 = 1_n8175 & 1_n7616;
assign 1_n2829 = 1_n5786 ^ 1_n1687;
assign 1_n10778 = 1_n5217 & 1_n12011;
assign 1_n11790 = ~1_n12134;
assign 1_n5599 = ~(1_n889 | 1_n7897);
assign 1_n7230 = 1_n4890 | 1_n4936;
assign 1_n11825 = 1_n7210 | 1_n12499;
assign 1_n10825 = ~(1_n6650 ^ 1_n3390);
assign 1_n9814 = 1_n11187 | 1_n8517;
assign 1_n7550 = ~(1_n4260 ^ 1_n2093);
assign 1_n6881 = ~1_n12539;
assign 1_n607 = ~(1_n4708 ^ 1_n10644);
assign 1_n11443 = 1_n6267 & 1_n3400;
assign 1_n11119 = 1_n8105 | 1_n13204;
assign 1_n5763 = ~(1_n5015 ^ 1_n11380);
assign 1_n8719 = ~1_n3828;
assign 1_n2394 = ~1_n9536;
assign 1_n1777 = 1_n2622 | 1_n8268;
assign 1_n2452 = ~1_n3409;
assign 1_n11968 = 1_n4791 & 1_n11517;
assign 1_n11997 = ~(1_n13134 ^ 1_n3935);
assign 1_n10603 = 1_n3225 | 1_n2675;
assign 1_n3728 = 1_n11114 | 1_n11522;
assign 1_n9652 = ~(1_n2294 ^ 1_n13017);
assign 1_n12211 = ~1_n3756;
assign 1_n5463 = ~(1_n7192 ^ 1_n8389);
assign 1_n277 = ~(1_n10323 ^ 1_n1955);
assign 1_n7773 = 1_n10462 | 1_n4230;
assign 1_n3648 = 1_n12264 & 1_n12355;
assign 1_n8913 = ~1_n2354;
assign 1_n2490 = 1_n12266 & 1_n11625;
assign 1_n4027 = ~(1_n369 ^ 1_n5339);
assign 1_n4387 = 1_n12987 ^ 1_n3141;
assign 1_n7925 = ~1_n443;
assign 1_n7533 = ~1_n9062;
assign 1_n4624 = 1_n9132 & 1_n770;
assign 1_n95 = 1_n2416 | 1_n8534;
assign 1_n3626 = ~(1_n11098 ^ 1_n4280);
assign 1_n1112 = ~(1_n13211 ^ 1_n8725);
assign 1_n1117 = ~1_n2591;
assign 1_n8054 = ~(1_n5370 ^ 1_n5983);
assign 1_n11445 = ~(1_n8836 ^ 1_n6953);
assign 1_n2567 = ~(1_n9654 ^ 1_n2866);
assign 1_n7511 = ~(1_n3807 ^ 1_n5624);
assign 1_n6735 = 1_n6028 | 1_n7723;
assign 1_n1615 = ~(1_n2699 ^ 1_n8946);
assign 1_n5680 = ~(1_n4400 | 1_n12285);
assign 1_n11221 = ~(1_n2237 ^ 1_n9081);
assign 1_n8511 = ~1_n3845;
assign 1_n7336 = 1_n879 & 1_n12413;
assign 1_n9976 = 1_n6354 | 1_n8707;
assign 1_n3141 = 1_n8259 & 1_n12511;
assign 1_n12611 = ~(1_n400 ^ 1_n8596);
assign 1_n10216 = ~(1_n5133 ^ 1_n10020);
assign 1_n2416 = ~1_n9570;
assign 1_n5734 = ~(1_n20 | 1_n732);
assign 1_n3065 = ~(1_n10191 | 1_n9414);
assign 1_n12324 = ~1_n7720;
assign 1_n9543 = 1_n684 & 1_n8617;
assign 1_n8884 = 1_n2640 ^ 1_n9983;
assign 1_n8851 = ~(1_n10600 ^ 1_n3897);
assign 1_n1847 = ~1_n4874;
assign 1_n4150 = ~(1_n5140 ^ 1_n6791);
assign 1_n12744 = 1_n971 | 1_n3981;
assign 1_n12748 = ~1_n12651;
assign 1_n12188 = 1_n9257;
assign 1_n7739 = 1_n3127 | 1_n3949;
assign 1_n2633 = 1_n349 & 1_n11283;
assign 1_n6384 = ~(1_n10602 ^ 1_n2771);
assign 1_n11149 = 1_n3544 ^ 1_n10553;
assign 1_n3616 = ~1_n2341;
assign 1_n4043 = ~(1_n10592 ^ 1_n12502);
assign 1_n11962 = ~(1_n8883 ^ 1_n9479);
assign 1_n5274 = 1_n4305 & 1_n407;
assign 1_n4294 = ~1_n12990;
assign 1_n868 = ~1_n11663;
assign 1_n5456 = 1_n6048 | 1_n5919;
assign 1_n12316 = ~1_n10142;
assign 1_n10089 = ~(1_n12339 | 1_n8342);
assign 1_n12425 = ~1_n1700;
assign 1_n119 = ~1_n3815;
assign 1_n5121 = 1_n10908 & 1_n5065;
assign 1_n1269 = ~1_n2388;
assign 1_n7803 = ~(1_n7613 | 1_n12303);
assign 1_n7759 = ~(1_n4858 ^ 1_n6896);
assign 1_n10817 = ~(1_n6694 ^ 1_n11017);
assign 1_n4423 = ~(1_n5424 ^ 1_n3838);
assign 1_n7187 = 1_n7263 | 1_n12492;
assign 1_n7439 = ~(1_n1048 ^ 1_n378);
assign 1_n2330 = ~1_n8267;
assign 1_n1569 = 1_n13147 & 1_n2602;
assign 1_n11931 = ~(1_n3533 ^ 1_n4754);
assign 1_n8043 = ~(1_n11386 ^ 1_n1497);
assign 1_n12443 = 1_n2273 & 1_n1598;
assign 1_n8130 = ~(1_n1471 | 1_n13033);
assign 1_n6518 = 1_n5626 | 1_n12291;
assign 1_n3581 = 1_n9897 & 1_n897;
assign 1_n12208 = ~(1_n6521 ^ 1_n7565);
assign 1_n7134 = ~(1_n4689 | 1_n4705);
assign 1_n1820 = ~1_n8290;
assign 1_n11613 = 1_n1965 & 1_n11784;
assign 1_n10120 = ~1_n12477;
assign 1_n7607 = 1_n10761 | 1_n2675;
assign 1_n2848 = ~1_n11111;
assign 1_n12024 = ~(1_n8432 ^ 1_n8045);
assign 1_n1967 = ~1_n9481;
assign 1_n2027 = 1_n9868 | 1_n1043;
assign 1_n12139 = ~(1_n12011 ^ 1_n4897);
assign 1_n9794 = ~(1_n8387 ^ 1_n10333);
assign 1_n10508 = ~1_n7384;
assign 1_n7831 = 1_n6880 & 1_n5072;
assign 1_n11663 = 1_n12478 & 1_n13139;
assign 1_n8816 = 1_n36 | 1_n1703;
assign 1_n6248 = 1_n372 & 1_n12572;
assign 1_n7049 = ~1_n10606;
assign 1_n6923 = 1_n7787 | 1_n6878;
assign 1_n10269 = 1_n12380 & 1_n5082;
assign 1_n1751 = 1_n6735 | 1_n9791;
assign 1_n4383 = ~(1_n897 ^ 1_n4126);
assign 1_n3328 = 1_n10771 & 1_n1878;
assign 1_n5469 = ~1_n9847;
assign 1_n9436 = ~1_n11012;
assign 1_n4132 = ~1_n2339;
assign 1_n11938 = ~(1_n8996 | 1_n3607);
assign 1_n12224 = ~1_n7659;
assign 1_n12254 = ~1_n2339;
assign 1_n2956 = ~1_n1344;
assign 1_n3966 = 1_n1354 | 1_n7723;
assign 1_n7822 = ~(1_n13145 ^ 1_n319);
assign 1_n5631 = 1_n5236 & 1_n9954;
assign 1_n10742 = 1_n8598 | 1_n4640;
assign 1_n3992 = 1_n9113 | 1_n10179;
assign 1_n2959 = 1_n6241 & 1_n1846;
assign 1_n5368 = 1_n4379 & 1_n2897;
assign 1_n10127 = ~1_n10876;
assign 1_n8492 = ~1_n6209;
assign 1_n5560 = ~(1_n2766 ^ 1_n7566);
assign 1_n11886 = ~(1_n5161 ^ 1_n6116);
assign 1_n3162 = ~(1_n6780 | 1_n8855);
assign 1_n7544 = ~1_n11372;
assign 1_n11530 = 1_n4620 | 1_n2675;
assign 1_n10520 = 1_n11392 | 1_n9760;
assign 1_n12733 = ~(1_n8057 | 1_n4415);
assign 1_n8399 = 1_n8954 ^ 1_n11294;
assign 1_n9113 = ~1_n10874;
assign 1_n10100 = 1_n2563 & 1_n1509;
assign 1_n7508 = 1_n7438 | 1_n3732;
assign 1_n11288 = 1_n7191 | 1_n1144;
assign 1_n12727 = ~(1_n12333 | 1_n12640);
assign 1_n10462 = ~1_n1916;
assign 1_n1673 = 1_n8426 | 1_n11754;
assign 1_n7614 = ~1_n9052;
assign 1_n8007 = ~(1_n2804 ^ 1_n10678);
assign 1_n1143 = 1_n10425 & 1_n10380;
assign 1_n9943 = ~(1_n2618 ^ 1_n11179);
assign 1_n2695 = 1_n10493 & 1_n9927;
assign 1_n5980 = 1_n11864 | 1_n7961;
assign 1_n12000 = ~1_n9591;
assign 1_n9748 = 1_n2759 | 1_n3653;
assign 1_n12999 = 1_n5296 | 1_n2277;
assign 1_n7674 = 1_n6854 | 1_n8268;
assign 1_n11398 = ~1_n13212;
assign 1_n1838 = 1_n10784 | 1_n10576;
assign 1_n7853 = ~(1_n8682 ^ 1_n9351);
assign 1_n1721 = ~(1_n9579 ^ 1_n7024);
assign 1_n11829 = 1_n8091 | 1_n10932;
assign 1_n793 = ~(1_n6965 | 1_n1626);
assign 1_n4859 = 1_n1150 | 1_n6005;
assign 1_n11418 = ~1_n10416;
assign 1_n9753 = ~(1_n8981 ^ 1_n598);
assign 1_n4257 = ~1_n2012;
assign 1_n9689 = ~(1_n4233 | 1_n5229);
assign 1_n5844 = 1_n1335 | 1_n3890;
assign 1_n3436 = ~(1_n7321 ^ 1_n11993);
assign 1_n10214 = 1_n11074 & 1_n8753;
assign 1_n5413 = 1_n9403 & 1_n4578;
assign 1_n1881 = ~1_n3910;
assign 1_n8264 = 1_n1618 | 1_n12273;
assign 1_n8877 = ~1_n1291;
assign 1_n245 = 1_n761 & 1_n5548;
assign 1_n10899 = ~(1_n5952 | 1_n205);
assign 1_n9646 = 1_n10501 | 1_n4373;
assign 1_n517 = 1_n5384 & 1_n6118;
assign 1_n2990 = ~(1_n12928 | 1_n2247);
assign 1_n2013 = ~1_n5952;
assign 1_n10536 = 1_n10637 | 1_n9234;
assign 1_n6724 = ~1_n12408;
assign 1_n6202 = 1_n8904 | 1_n10029;
assign 1_n1817 = 1_n4038 | 1_n9984;
assign 1_n835 = ~(1_n344 ^ 1_n6639);
assign 1_n8933 = ~(1_n2910 | 1_n1430);
assign 1_n2839 = ~(1_n12020 ^ 1_n964);
assign 1_n7253 = 1_n2097 | 1_n2917;
assign 1_n7915 = ~(1_n8805 ^ 1_n11623);
assign 1_n12532 = 1_n6369 & 1_n13167;
assign 1_n764 = 1_n8228 & 1_n5920;
assign 1_n12950 = ~(1_n1125 ^ 1_n12488);
assign 1_n7730 = ~1_n5167;
assign 1_n3864 = ~(1_n5294 | 1_n8289);
assign 1_n4167 = 1_n9113 | 1_n177;
assign 1_n3398 = 1_n8877 & 1_n11133;
assign 1_n7268 = ~(1_n8923 ^ 1_n7479);
assign 1_n973 = 1_n13026 | 1_n177;
assign 1_n7464 = 1_n9303 & 1_n11029;
assign 1_n944 = 1_n9371 | 1_n12016;
assign 1_n6550 = 1_n1586 & 1_n2253;
assign 1_n10437 = ~1_n1302;
assign 1_n4485 = 1_n1529 | 1_n604;
assign 1_n5418 = ~(1_n9221 ^ 1_n12344);
assign 1_n11716 = ~(1_n6952 ^ 1_n8149);
assign 1_n12541 = ~(1_n7349 | 1_n12447);
assign 1_n6017 = ~(1_n12821 ^ 1_n9452);
assign 1_n12531 = ~(1_n10088 ^ 1_n12494);
assign 1_n1183 = 1_n6168 & 1_n12853;
assign 1_n9744 = 1_n13041 & 1_n3661;
assign 1_n7953 = 1_n1261 | 1_n177;
assign 1_n13142 = ~(1_n9588 ^ 1_n10708);
assign 1_n190 = 1_n9983 | 1_n8246;
assign 1_n1690 = ~(1_n11837 | 1_n913);
assign 1_n5112 = 1_n6100 & 1_n10389;
assign 1_n13036 = ~1_n9187;
assign 1_n4449 = ~(1_n3923 ^ 1_n261);
assign 1_n2082 = 1_n7990 & 1_n3609;
assign 1_n6696 = ~(1_n4988 ^ 1_n9686);
assign 1_n12198 = 1_n1947 | 1_n8018;
assign 1_n9342 = 1_n1334 | 1_n7926;
assign 1_n128 = ~1_n13011;
assign 1_n881 = ~1_n10951;
assign 1_n8401 = 1_n1727 | 1_n8083;
assign 1_n717 = ~(1_n475 ^ 1_n10012);
assign 1_n9324 = 1_n8948 & 1_n8786;
assign 1_n11234 = ~(1_n10186 | 1_n10206);
assign 1_n888 = 1_n8295 & 1_n6694;
assign 1_n1353 = ~1_n4748;
assign 1_n5901 = ~(1_n3973 ^ 1_n11389);
assign 1_n4570 = ~(1_n1426 ^ 1_n3751);
assign 1_n11352 = ~1_n7411;
assign 1_n12446 = 1_n1068 | 1_n5530;
assign 1_n9008 = ~1_n7164;
assign 1_n1835 = ~(1_n175 ^ 1_n9377);
assign 1_n5253 = ~(1_n625 | 1_n9390);
assign 1_n3461 = 1_n10676 & 1_n1091;
assign 1_n6704 = ~(1_n633 ^ 1_n1000);
assign 1_n5744 = 1_n9739 | 1_n10106;
assign 1_n7219 = 1_n11256 | 1_n9657;
assign 1_n12394 = 1_n1315 & 1_n10174;
assign 1_n5023 = ~(1_n3179 ^ 1_n11465);
assign 1_n2647 = ~(1_n8428 ^ 1_n11341);
assign 1_n6730 = ~(1_n6498 ^ 1_n4246);
assign 1_n1507 = 1_n734 | 1_n10956;
assign 1_n8731 = ~(1_n962 ^ 1_n11405);
assign 1_n9389 = 1_n11007 | 1_n2675;
assign 1_n11556 = ~(1_n9823 ^ 1_n2704);
assign 1_n5420 = ~1_n3181;
assign 1_n11338 = 1_n21 & 1_n2740;
assign 1_n7777 = 1_n2217 | 1_n10871;
assign 1_n9039 = 1_n6068 ^ 1_n5834;
assign 1_n10432 = 1_n3161 & 1_n3249;
assign 1_n7627 = ~(1_n9678 | 1_n5171);
assign 1_n10731 = 1_n992 | 1_n7239;
assign 1_n8012 = ~1_n3283;
assign 1_n3816 = ~1_n5062;
assign 1_n8481 = ~1_n3939;
assign 1_n5702 = ~(1_n7096 ^ 1_n7458);
assign 1_n2963 = 1_n9226 | 1_n9521;
assign 1_n7972 = 1_n10919 | 1_n4765;
assign 1_n1449 = ~(1_n12894 ^ 1_n6459);
assign 1_n10968 = ~(1_n11710 ^ 1_n11702);
assign 1_n8703 = 1_n7900 | 1_n10106;
assign 1_n2430 = ~1_n10458;
assign 1_n11056 = 1_n5400 & 1_n4047;
assign 1_n3959 = ~(1_n7542 ^ 1_n3710);
assign 1_n9205 = 1_n11965 | 1_n4844;
assign 1_n9619 = 1_n4382 & 1_n11109;
assign 1_n2106 = 1_n3327 | 1_n926;
assign 1_n7672 = ~1_n12579;
assign 1_n10985 = 1_n9135 & 1_n12548;
assign 1_n5770 = 1_n3311 & 1_n6085;
assign 1_n9524 = ~(1_n4851 | 1_n2998);
assign 1_n9153 = 1_n4213 | 1_n4255;
assign 1_n10119 = ~(1_n6268 ^ 1_n4358);
assign 1_n8400 = ~1_n11109;
assign 1_n8 = 1_n8645 | 1_n8563;
assign 1_n5378 = 1_n11430 & 1_n7519;
assign 1_n2364 = ~(1_n8638 ^ 1_n10679);
assign 1_n5978 = 1_n818 & 1_n6563;
assign 1_n10621 = ~(1_n12851 ^ 1_n13112);
assign 1_n2062 = 1_n4198 | 1_n4373;
assign 1_n8723 = ~1_n105;
assign 1_n6638 = ~1_n7374;
assign 1_n8433 = 1_n325 & 1_n3739;
assign 1_n2385 = ~1_n7802;
assign 1_n13231 = ~(1_n4785 ^ 1_n4120);
assign 1_n9318 = 1_n6841 | 1_n8129;
assign 1_n3372 = 1_n4485 & 1_n5936;
assign 1_n7604 = ~(1_n3032 ^ 1_n847);
assign 1_n11169 = 1_n9707 & 1_n8888;
assign 1_n8540 = ~1_n10787;
assign 1_n6148 = ~(1_n11742 ^ 1_n3098);
assign 1_n8833 = 1_n3724 | 1_n7959;
assign 1_n6526 = 1_n3395 ^ 1_n11402;
assign 1_n2944 = 1_n11592 & 1_n4491;
assign 1_n3694 = ~(1_n6176 ^ 1_n13062);
assign 1_n9617 = 1_n7069 | 1_n1694;
assign 1_n2897 = 1_n12758 | 1_n5797;
assign 1_n5842 = ~1_n951;
assign 1_n4545 = ~(1_n12897 | 1_n5133);
assign 1_n9388 = ~(1_n5323 | 1_n4094);
assign 1_n9124 = 1_n8082 | 1_n1026;
assign 1_n10556 = ~(1_n29 ^ 1_n7029);
assign 1_n7345 = ~(1_n10762 ^ 1_n363);
assign 1_n6462 = 1_n11702 & 1_n11710;
assign 1_n10744 = ~(1_n4232 ^ 1_n5137);
assign 1_n4983 = ~(1_n2951 | 1_n4369);
assign 1_n11785 = 1_n2465 & 1_n1868;
assign 1_n5875 = ~1_n5920;
assign 1_n5171 = 1_n10727 & 1_n1967;
assign 1_n2883 = 1_n2068 & 1_n12284;
assign 1_n8984 = 1_n11102 | 1_n2280;
assign 1_n1055 = ~1_n2791;
assign 1_n3238 = ~(1_n6892 | 1_n9952);
assign 1_n13219 = ~(1_n2370 ^ 1_n13161);
assign 1_n6832 = ~(1_n5627 ^ 1_n9009);
assign 1_n4398 = ~1_n7059;
assign 1_n4797 = ~(1_n6352 ^ 1_n9616);
assign 1_n9508 = ~(1_n12988 ^ 1_n2012);
assign 1_n4482 = 1_n3209 & 1_n8760;
assign 1_n1412 = ~(1_n3666 ^ 1_n10218);
assign 1_n11976 = ~(1_n12097 ^ 1_n1375);
assign 1_n7073 = ~1_n3199;
assign 1_n9467 = ~(1_n4602 ^ 1_n11487);
assign 1_n8119 = ~(1_n402 ^ 1_n12679);
assign 1_n813 = ~1_n9528;
assign 1_n8326 = 1_n7319 & 1_n12764;
assign 1_n5474 = 1_n5993 | 1_n1298;
assign 1_n6535 = ~(1_n2088 ^ 1_n11731);
assign 1_n6929 = 1_n7730 | 1_n3825;
assign 1_n8675 = 1_n6522 ^ 1_n11840;
assign 1_n4640 = 1_n12128;
assign 1_n9061 = 1_n525 & 1_n10753;
assign 1_n1092 = ~(1_n7363 ^ 1_n11216);
assign 1_n9326 = 1_n2046 | 1_n12637;
assign 1_n12784 = 1_n5823 & 1_n5381;
assign 1_n11666 = 1_n5522 & 1_n11056;
assign 1_n733 = ~(1_n8424 ^ 1_n2225);
assign 1_n2597 = ~(1_n12590 ^ 1_n4410);
assign 1_n6378 = 1_n4983 | 1_n553;
assign 1_n1821 = 1_n8950 | 1_n12695;
assign 1_n1366 = ~1_n10869;
assign 1_n7569 = 1_n6749 | 1_n7076;
assign 1_n5187 = 1_n12458 | 1_n4303;
assign 1_n9941 = ~(1_n10312 ^ 1_n4353);
assign 1_n1711 = 1_n1158 | 1_n1713;
assign 1_n5090 = 1_n9913 | 1_n11868;
assign 1_n12826 = ~(1_n7442 | 1_n12464);
assign 1_n12061 = ~(1_n7694 ^ 1_n9438);
assign 1_n4827 = 1_n2462 | 1_n10319;
assign 1_n5460 = ~1_n3769;
assign 1_n2607 = 1_n294 | 1_n11164;
assign 1_n11084 = 1_n3527;
assign 1_n1134 = ~1_n2619;
assign 1_n8878 = 1_n10332 | 1_n1344;
assign 1_n671 = 1_n3957 | 1_n11273;
assign 1_n3213 = 1_n9383 | 1_n3981;
assign 1_n13233 = ~(1_n11973 | 1_n12163);
assign 1_n3345 = 1_n2723 | 1_n4209;
assign 1_n7275 = 1_n10999 | 1_n10342;
assign 1_n9500 = ~(1_n4403 | 1_n1828);
assign 1_n8259 = ~1_n2966;
assign 1_n4565 = 1_n10920 & 1_n5497;
assign 1_n7172 = ~(1_n8606 ^ 1_n3342);
assign 1_n6795 = 1_n6136 & 1_n8022;
assign 1_n10829 = ~(1_n2995 ^ 1_n2840);
assign 1_n8800 = ~1_n5722;
assign 1_n3116 = ~1_n2647;
assign 1_n7532 = ~1_n497;
assign 1_n5849 = ~(1_n13070 | 1_n6840);
assign 1_n1997 = 1_n7770 | 1_n8066;
assign 1_n9020 = 1_n10149 | 1_n9413;
assign 1_n5242 = 1_n1750;
assign 1_n7468 = 1_n719 | 1_n290;
assign 1_n9773 = 1_n1912 & 1_n13060;
assign 1_n2704 = ~(1_n10766 ^ 1_n7287);
assign 1_n5364 = ~(1_n10390 ^ 1_n12034);
assign 1_n7784 = ~1_n13223;
assign 1_n6963 = ~(1_n5800 | 1_n1624);
assign 1_n3571 = 1_n9162 | 1_n12328;
assign 1_n5533 = ~1_n3043;
assign 1_n2135 = ~1_n1982;
assign 1_n2380 = 1_n5465 | 1_n6861;
assign 1_n7191 = ~1_n12651;
assign 1_n11626 = 1_n8584 & 1_n4814;
assign 1_n10769 = 1_n8731 ^ 1_n9437;
assign 1_n7107 = ~(1_n8457 ^ 1_n6903);
assign 1_n13085 = 1_n2789 | 1_n8029;
assign 1_n3615 = 1_n12933 & 1_n3526;
assign 1_n3118 = ~1_n12217;
assign 1_n10170 = 1_n12202 | 1_n2042;
assign 1_n6457 = 1_n6614 | 1_n6996;
assign 1_n2849 = ~1_n10395;
assign 1_n10721 = ~(1_n4266 ^ 1_n483);
assign 1_n7927 = 1_n11407 | 1_n4787;
assign 1_n5943 = 1_n121 | 1_n9118;
assign 1_n9371 = ~(1_n454 ^ 1_n1179);
assign 1_n12112 = 1_n63 | 1_n479;
assign 1_n4849 = ~(1_n1508 ^ 1_n4955);
assign 1_n4400 = 1_n12295 | 1_n10319;
assign 1_n7943 = ~(1_n9498 ^ 1_n6217);
assign 1_n4987 = 1_n8680 & 1_n222;
assign 1_n2822 = ~1_n11809;
assign 1_n12559 = ~(1_n8497 ^ 1_n10634);
assign 1_n5280 = 1_n4042 & 1_n1646;
assign 1_n2886 = 1_n10550 | 1_n6258;
assign 1_n12817 = 1_n9174 & 1_n9250;
assign 1_n10944 = ~1_n10850;
assign 1_n10530 = 1_n10357 | 1_n409;
assign 1_n11942 = ~1_n3014;
assign 1_n2579 = ~1_n12429;
assign 1_n3079 = 1_n8378 & 1_n12080;
assign 1_n7355 = 1_n1320 | 1_n9223;
assign 1_n4692 = 1_n4465 | 1_n8534;
assign 1_n5520 = ~1_n5758;
assign 1_n418 = ~1_n12622;
assign 1_n4845 = ~(1_n914 ^ 1_n6840);
assign 1_n5938 = 1_n1602 ^ 1_n1612;
assign 1_n10929 = ~1_n9846;
assign 1_n3893 = ~(1_n12199 ^ 1_n13004);
assign 1_n293 = 1_n2743 & 1_n1620;
assign 1_n5967 = 1_n3006 & 1_n5729;
assign 1_n8458 = ~1_n12614;
assign 1_n3261 = ~(1_n6016 ^ 1_n8782);
assign 1_n4391 = 1_n10877 | 1_n4936;
assign 1_n1893 = ~1_n2882;
assign 1_n2413 = 1_n4171 | 1_n10516;
assign 1_n12827 = ~(1_n2177 ^ 1_n7571);
assign 1_n12428 = 1_n5420 & 1_n10980;
assign 1_n11743 = 1_n2409 & 1_n12026;
assign 1_n3429 = ~1_n13188;
assign 1_n4924 = ~(1_n10745 | 1_n5457);
assign 1_n6222 = ~(1_n5016 ^ 1_n1238);
assign 1_n12852 = ~(1_n4978 ^ 1_n5236);
assign 1_n9707 = 1_n3311 & 1_n13058;
assign 1_n3621 = 1_n6629 | 1_n12188;
assign 1_n3150 = ~(1_n4934 ^ 1_n23);
assign 1_n3857 = ~(1_n1060 | 1_n5860);
assign 1_n4256 = ~1_n1836;
assign 1_n1850 = 1_n5009 & 1_n7632;
assign 1_n10696 = ~1_n411;
assign 1_n8311 = ~(1_n6744 ^ 1_n5263);
assign 1_n2045 = ~1_n10751;
assign 1_n3627 = 1_n11449 | 1_n12847;
assign 1_n7481 = ~1_n4708;
assign 1_n9474 = 1_n7068 | 1_n2544;
assign 1_n5083 = ~(1_n7418 ^ 1_n3015);
assign 1_n12603 = ~(1_n3695 ^ 1_n4774);
assign 1_n6805 = 1_n10045 | 1_n2675;
assign 1_n9378 = ~1_n12850;
assign 1_n3934 = ~(1_n7368 | 1_n11916);
assign 1_n6883 = ~1_n10606;
assign 1_n1191 = ~1_n1231;
assign 1_n5794 = ~(1_n12479 ^ 1_n2655);
assign 1_n7876 = 1_n9112 | 1_n2671;
assign 1_n5407 = 1_n4366 | 1_n2970;
assign 1_n11991 = ~(1_n5207 ^ 1_n1708);
assign 1_n5040 = ~1_n6826;
assign 1_n5521 = ~1_n11030;
assign 1_n1791 = 1_n2940 | 1_n11756;
assign 1_n4489 = 1_n10798 | 1_n6404;
assign 1_n7209 = ~(1_n8517 ^ 1_n6324);
assign 1_n6717 = 1_n10137 | 1_n8268;
assign 1_n1678 = 1_n4701 & 1_n10507;
assign 1_n7825 = ~1_n9093;
assign 1_n10660 = 1_n10266 | 1_n1695;
assign 1_n13205 = ~(1_n11716 ^ 1_n873);
assign 1_n9851 = ~(1_n6001 | 1_n10866);
assign 1_n3156 = 1_n5163 | 1_n3981;
assign 1_n7060 = 1_n8659 & 1_n2153;
assign 1_n11165 = ~1_n5311;
assign 1_n2107 = 1_n2296 | 1_n2387;
assign 1_n1780 = ~(1_n4417 ^ 1_n12156);
assign 1_n9347 = 1_n11509 & 1_n1254;
assign 1_n7653 = ~(1_n1169 ^ 1_n10401);
assign 1_n12161 = 1_n12109 | 1_n206;
assign 1_n7567 = ~1_n11416;
assign 1_n9759 = ~(1_n13104 | 1_n8566);
assign 1_n12546 = ~(1_n8914 ^ 1_n12231);
assign 1_n7245 = ~(1_n9347 | 1_n13030);
assign 1_n11715 = ~(1_n649 ^ 1_n5691);
assign 1_n11002 = ~1_n9401;
assign 1_n9257 = ~1_n7772;
assign 1_n9390 = 1_n11365 & 1_n6531;
assign 1_n1627 = 1_n4583 & 1_n2925;
assign 1_n225 = ~(1_n11026 | 1_n661);
assign 1_n13204 = 1_n2613 & 1_n12233;
assign 1_n5567 = ~(1_n5872 | 1_n1170);
assign 1_n12336 = 1_n9794 | 1_n9681;
assign 1_n8331 = 1_n8875 & 1_n8491;
assign 1_n12975 = 1_n5206 & 1_n9789;
assign 1_n6166 = ~1_n11030;
assign 1_n9236 = 1_n4278 ^ 1_n1879;
assign 1_n12415 = 1_n2479 & 1_n8292;
assign 1_n10429 = 1_n2487 | 1_n9075;
assign 1_n12270 = 1_n6220 | 1_n8225;
assign 1_n4841 = ~1_n9824;
assign 1_n8200 = 1_n6231 | 1_n5797;
assign 1_n3424 = 1_n109 | 1_n4052;
assign 1_n475 = 1_n1893 | 1_n206;
assign 1_n9670 = 1_n98 | 1_n10286;
assign 1_n9601 = ~1_n4423;
assign 1_n1800 = 1_n8837 | 1_n5100;
assign 1_n167 = 1_n9330 & 1_n11357;
assign 1_n720 = 1_n785 | 1_n4373;
assign 1_n3022 = 1_n10412 | 1_n5262;
assign 1_n6053 = ~(1_n13024 | 1_n6887);
assign 1_n7423 = ~(1_n10546 ^ 1_n2277);
assign 1_n9019 = ~1_n1916;
assign 1_n6172 = 1_n11781 | 1_n8505;
assign 1_n10792 = ~1_n6409;
assign 1_n2125 = ~(1_n819 | 1_n2324);
assign 1_n11212 = ~1_n7974;
assign 1_n12829 = 1_n10830 | 1_n7530;
assign 1_n82 = 1_n8645 | 1_n3981;
assign 1_n2611 = 1_n8576 & 1_n8825;
assign 1_n2444 = 1_n1571 | 1_n11668;
assign 1_n11558 = 1_n11400 | 1_n111;
assign 1_n7896 = ~(1_n6382 ^ 1_n5183);
assign 1_n1171 = 1_n11132 & 1_n1854;
assign 1_n6349 = 1_n7805 | 1_n11144;
assign 1_n12203 = ~1_n8468;
assign 1_n6277 = ~(1_n5563 ^ 1_n1118);
assign 1_n3091 = ~1_n2376;
assign 1_n925 = 1_n4846 & 1_n7678;
assign 1_n7449 = ~(1_n5091 ^ 1_n907);
assign 1_n8192 = ~(1_n4445 ^ 1_n6970);
assign 1_n8407 = ~(1_n8385 ^ 1_n3406);
assign 1_n7509 = ~(1_n13053 ^ 1_n1851);
assign 1_n2562 = 1_n7557 & 1_n3430;
assign 1_n6279 = 1_n13106 | 1_n6963;
assign 1_n4907 = 1_n2118 | 1_n4230;
assign 1_n11874 = 1_n1323 | 1_n13238;
assign 1_n2916 = 1_n3026 | 1_n13209;
assign 1_n2572 = ~1_n10744;
assign 1_n10830 = ~1_n8163;
assign 1_n12544 = ~1_n7428;
assign 1_n5968 = ~1_n11574;
assign 1_n7585 = 1_n10041 & 1_n11741;
assign 1_n1078 = 1_n821 | 1_n10904;
assign 1_n8926 = 1_n7930 | 1_n7935;
assign 1_n2979 = ~(1_n2091 ^ 1_n5580);
assign 1_n6834 = 1_n3313 & 1_n14;
assign 1_n8886 = ~(1_n5250 ^ 1_n11345);
assign 1_n11955 = ~(1_n9254 ^ 1_n5635);
assign 1_n12393 = 1_n8325 | 1_n12695;
assign 1_n12863 = 1_n9891 ^ 1_n4997;
assign 1_n13103 = 1_n1688 | 1_n10871;
assign 1_n3090 = ~(1_n3563 ^ 1_n12460);
assign 1_n2711 = ~1_n11109;
assign 1_n11933 = ~1_n2341;
assign 1_n3821 = 1_n319 & 1_n13145;
assign 1_n5590 = 1_n4132 | 1_n7723;
assign 1_n3759 = ~(1_n3042 | 1_n12403);
assign 1_n13189 = 1_n9724 & 1_n11956;
assign 1_n12620 = ~1_n11181;
assign 1_n4503 = 1_n12017 & 1_n2474;
assign 1_n1723 = ~(1_n6948 ^ 1_n4395);
assign 1_n2198 = 1_n3178 & 1_n834;
assign 1_n10942 = ~(1_n9624 ^ 1_n5710);
assign 1_n8384 = ~1_n4713;
assign 1_n3136 = 1_n9345 & 1_n4003;
assign 1_n2003 = 1_n5321 | 1_n1013;
assign 1_n11584 = ~(1_n59 ^ 1_n12209);
assign 1_n2563 = 1_n8143 | 1_n12328;
assign 1_n6580 = ~1_n6632;
assign 1_n11557 = 1_n11237 | 1_n8494;
assign 1_n4468 = 1_n713 | 1_n8319;
assign 1_n7274 = ~(1_n10653 ^ 1_n7397);
assign 1_n5525 = ~(1_n4896 | 1_n7910);
assign 1_n93 = ~1_n7161;
assign 1_n3668 = ~(1_n9960 | 1_n9393);
assign 1_n4153 = 1_n2148 | 1_n2133;
assign 1_n13091 = 1_n5122 & 1_n35;
assign 1_n3035 = 1_n5586 & 1_n2498;
assign 1_n9614 = 1_n7966 | 1_n177;
assign 1_n13243 = 1_n5347 | 1_n5373;
assign 1_n96 = ~1_n9039;
assign 1_n10876 = 1_n2691 & 1_n8363;
assign 1_n8266 = 1_n1783 | 1_n2757;
assign 1_n7207 = ~(1_n2987 | 1_n2822);
assign 1_n13010 = 1_n5704 | 1_n10194;
assign 1_n6374 = 1_n12212 | 1_n3379;
assign 1_n1617 = ~(1_n7064 ^ 1_n11317);
assign 1_n5776 = ~(1_n1722 ^ 1_n12103);
assign 1_n7139 = 1_n575 | 1_n12870;
assign 1_n8917 = 1_n5048 | 1_n8702;
assign 1_n3003 = 1_n11893 & 1_n11705;
assign 1_n5914 = 1_n7518 & 1_n7112;
assign 1_n2687 = 1_n12178 | 1_n7840;
assign 1_n6135 = 1_n2312 | 1_n7820;
assign 1_n8657 = 1_n5055 & 1_n5593;
assign 1_n4932 = ~(1_n6757 | 1_n11000);
assign 1_n10824 = 1_n3595 & 1_n9109;
assign 1_n634 = 1_n1237 & 1_n3216;
assign 1_n11996 = 1_n9527 | 1_n4469;
assign 1_n2137 = ~(1_n4831 ^ 1_n13034);
assign 1_n10325 = 1_n10989 & 1_n1226;
assign 1_n6676 = 1_n6347 | 1_n12377;
assign 1_n10828 = ~(1_n8584 ^ 1_n4119);
assign 1_n12238 = ~(1_n310 ^ 1_n6503);
assign 1_n1852 = ~(1_n9695 ^ 1_n8305);
assign 1_n7378 = 1_n4516 & 1_n5121;
assign 1_n11917 = 1_n12834 | 1_n7950;
assign 1_n2901 = 1_n4566 | 1_n8719;
assign 1_n6157 = 1_n7564 | 1_n11415;
assign 1_n5634 = ~1_n1084;
assign 1_n10867 = 1_n3239 & 1_n3037;
assign 1_n11146 = 1_n9969 & 1_n7732;
assign 1_n1604 = ~(1_n12076 ^ 1_n13162);
assign 1_n7466 = ~(1_n7250 | 1_n1822);
assign 1_n9787 = 1_n4619 & 1_n5288;
assign 1_n6020 = ~(1_n9094 ^ 1_n431);
assign 1_n8521 = 1_n3870 & 1_n5584;
assign 1_n3576 = 1_n7418 & 1_n11744;
assign 1_n3101 = 1_n1621 | 1_n8534;
assign 1_n7734 = 1_n4288 & 1_n10503;
assign 1_n6612 = 1_n1868 | 1_n2465;
assign 1_n3485 = 1_n940 & 1_n568;
assign 1_n1539 = 1_n5857 | 1_n6177;
assign 1_n1026 = 1_n8160;
assign 1_n13148 = ~1_n8183;
assign 1_n7697 = 1_n9639 & 1_n9168;
assign 1_n10333 = ~(1_n1163 ^ 1_n5022);
assign 1_n4215 = 1_n3940 | 1_n8038;
assign 1_n10934 = ~(1_n920 ^ 1_n11282);
assign 1_n2817 = ~(1_n2350 | 1_n1073);
assign 1_n6915 = ~(1_n1393 | 1_n7708);
assign 1_n6958 = 1_n11719 & 1_n8158;
assign 1_n6291 = 1_n12806 | 1_n2589;
assign 1_n6071 = ~(1_n2285 ^ 1_n5304);
assign 1_n13225 = 1_n5032 & 1_n6426;
assign 1_n1391 = ~(1_n387 ^ 1_n10887);
assign 1_n10221 = ~1_n6794;
assign 1_n12230 = 1_n12023 | 1_n3698;
assign 1_n8258 = ~(1_n7503 ^ 1_n3794);
assign 1_n10800 = 1_n937 & 1_n3769;
assign 1_n880 = 1_n7661 | 1_n11668;
assign 1_n7280 = ~(1_n10048 ^ 1_n12842);
assign 1_n12739 = ~(1_n6526 ^ 1_n8066);
assign 1_n5829 = 1_n7607 | 1_n3501;
assign 1_n12617 = ~1_n3832;
assign 1_n2173 = 1_n7167 | 1_n12657;
assign 1_n9556 = ~(1_n5335 ^ 1_n3453);
assign 1_n278 = ~1_n8714;
assign 1_n9445 = 1_n8243 | 1_n11267;
assign 1_n8649 = 1_n351 & 1_n9764;
assign 1_n3265 = 1_n9711 | 1_n1463;
assign 1_n12143 = 1_n6515 & 1_n2393;
assign 1_n12595 = ~1_n9666;
assign 1_n5307 = 1_n3995 & 1_n9899;
assign 1_n12896 = ~(1_n1617 | 1_n5596);
assign 1_n8557 = ~(1_n12883 ^ 1_n8441);
assign 1_n4505 = 1_n6492 & 1_n11464;
assign 1_n4668 = 1_n114 | 1_n121;
assign 1_n3262 = ~(1_n1361 ^ 1_n4849);
assign 1_n5716 = 1_n8926 & 1_n5736;
assign 1_n7190 = 1_n710 | 1_n11500;
assign 1_n580 = ~(1_n8112 ^ 1_n7940);
assign 1_n10121 = ~(1_n8127 ^ 1_n9298);
assign 1_n8173 = ~1_n12284;
assign 1_n1447 = ~1_n3076;
assign 1_n12028 = ~(1_n4389 ^ 1_n4746);
assign 1_n2973 = 1_n829 | 1_n5242;
assign 1_n9332 = 1_n3013 | 1_n2398;
assign 1_n13237 = ~(1_n7697 | 1_n11172);
assign 1_n884 = 1_n3096 | 1_n12383;
assign 1_n10093 = 1_n3584 | 1_n376;
assign 1_n12778 = ~1_n7882;
assign 1_n7898 = 1_n4653 & 1_n2514;
assign 1_n6713 = ~(1_n3385 ^ 1_n6485);
assign 1_n10345 = ~1_n1148;
assign 1_n11129 = ~(1_n2754 ^ 1_n11458);
assign 1_n11481 = 1_n740 | 1_n4847;
assign 1_n524 = 1_n5788 | 1_n12811;
assign 1_n11954 = 1_n445 | 1_n121;
assign 1_n584 = ~1_n2771;
assign 1_n6669 = 1_n1571 | 1_n13086;
assign 1_n2740 = 1_n3005 | 1_n13017;
assign 1_n6498 = ~(1_n8604 ^ 1_n11030);
assign 1_n4494 = 1_n6371 | 1_n10071;
assign 1_n6856 = 1_n12431 | 1_n8385;
assign 1_n3385 = 1_n1152 | 1_n9195;
assign 1_n5635 = ~(1_n2532 ^ 1_n8140);
assign 1_n12082 = ~1_n32;
assign 1_n11333 = ~1_n772;
assign 1_n6445 = ~(1_n8009 ^ 1_n6628);
assign 1_n6293 = ~1_n2771;
assign 1_n1064 = 1_n937 & 1_n8233;
assign 1_n5007 = 1_n10641 | 1_n6635;
assign 1_n11914 = ~1_n5012;
assign 1_n11701 = 1_n2546 | 1_n8076;
assign 1_n7930 = ~1_n3085;
assign 1_n4270 = ~(1_n12047 | 1_n5346);
assign 1_n1932 = 1_n11910 | 1_n4490;
assign 1_n9005 = ~1_n7087;
assign 1_n5261 = ~1_n12912;
assign 1_n8514 = ~1_n2071;
assign 1_n12952 = ~1_n10544;
assign 1_n3046 = 1_n2518 & 1_n5331;
assign 1_n6106 = ~(1_n11637 | 1_n2432);
assign 1_n12426 = 1_n11373 & 1_n8829;
assign 1_n9740 = 1_n10066 | 1_n6690;
assign 1_n10617 = ~(1_n1233 | 1_n13213);
assign 1_n1289 = ~1_n2656;
assign 1_n2925 = ~(1_n12167 ^ 1_n11586);
assign 1_n8072 = ~(1_n505 ^ 1_n3377);
assign 1_n5899 = ~1_n11561;
assign 1_n4260 = ~1_n6920;
assign 1_n12142 = ~(1_n8745 ^ 1_n919);
assign 1_n7154 = ~1_n3567;
assign 1_n10304 = 1_n2868 | 1_n10350;
assign 1_n2091 = 1_n542 | 1_n6404;
assign 1_n4337 = 1_n2122 & 1_n7388;
assign 1_n6424 = ~(1_n3775 ^ 1_n3756);
assign 1_n12533 = 1_n2449 | 1_n2675;
assign 1_n5251 = ~1_n3226;
assign 1_n4823 = 1_n12795 | 1_n4453;
assign 1_n6214 = 1_n2456 | 1_n13233;
assign 1_n1379 = 1_n10920 | 1_n5497;
assign 1_n6440 = ~(1_n4154 ^ 1_n898);
assign 1_n3514 = ~1_n1038;
assign 1_n234 = 1_n6299 & 1_n8064;
assign 1_n7615 = 1_n11080 & 1_n10155;
assign 1_n4945 = 1_n1873 | 1_n12074;
assign 1_n2857 = ~(1_n4436 ^ 1_n642);
assign 1_n1947 = ~(1_n10211 | 1_n3734);
assign 1_n6155 = ~(1_n4742 ^ 1_n11084);
assign 1_n8029 = ~1_n12520;
assign 1_n12740 = ~(1_n12720 ^ 1_n12175);
assign 1_n1206 = 1_n5595 | 1_n12388;
assign 1_n5965 = 1_n956 | 1_n12188;
assign 1_n11117 = ~(1_n1319 ^ 1_n957);
assign 1_n6684 = 1_n4364 & 1_n12165;
assign 1_n2657 = ~1_n5920;
assign 1_n6133 = ~1_n4335;
assign 1_n9967 = 1_n10929 | 1_n6635;
assign 1_n10881 = ~(1_n3753 ^ 1_n6819);
assign 1_n5942 = ~(1_n7984 ^ 1_n12261);
assign 1_n8821 = ~(1_n8474 ^ 1_n1827);
assign 1_n6517 = 1_n44 | 1_n4947;
assign 1_n9594 = ~(1_n6473 | 1_n10694);
assign 1_n9667 = ~(1_n7931 ^ 1_n915);
assign 1_n2381 = ~(1_n3631 ^ 1_n10841);
assign 1_n12356 = 1_n2605 & 1_n5245;
assign 1_n10992 = ~(1_n1658 ^ 1_n7233);
assign 1_n2311 = 1_n1740 & 1_n9881;
assign 1_n10017 = ~1_n5969;
assign 1_n10814 = ~1_n13060;
assign 1_n4605 = 1_n9625 | 1_n1767;
assign 1_n970 = 1_n11236 & 1_n6937;
assign 1_n12596 = ~1_n854;
assign 1_n7500 = ~(1_n9996 ^ 1_n1721);
assign 1_n454 = 1_n3972 | 1_n8534;
assign 1_n13170 = ~1_n3085;
assign 1_n7923 = 1_n4885 & 1_n585;
assign 1_n1217 = ~(1_n8771 ^ 1_n3842);
assign 1_n12241 = ~1_n6009;
assign 1_n8306 = ~1_n9906;
assign 1_n4777 = ~(1_n4449 ^ 1_n9077);
assign 1_n6911 = 1_n4387 | 1_n726;
assign 1_n9710 = ~1_n7208;
assign 1_n6296 = ~(1_n12386 ^ 1_n6261);
assign 1_n9348 = ~(1_n3684 ^ 1_n9189);
assign 1_n3171 = 1_n795 | 1_n12930;
assign 1_n5768 = 1_n10770 & 1_n6392;
assign 1_n8103 = ~(1_n4617 | 1_n5162);
assign 1_n11140 = 1_n1344 ^ 1_n3950;
assign 1_n6345 = 1_n5176 | 1_n3640;
assign 1_n6401 = 1_n5841 | 1_n542;
assign 1_n11930 = ~(1_n2555 ^ 1_n11479);
assign 1_n7235 = 1_n11723 | 1_n2893;
assign 1_n8794 = ~(1_n10472 ^ 1_n12148);
assign 1_n10474 = ~1_n11324;
assign 1_n3177 = 1_n13068 & 1_n7361;
assign 1_n4725 = 1_n10023 | 1_n11042;
assign 1_n9299 = 1_n1989 | 1_n7805;
assign 1_n4549 = ~(1_n3592 ^ 1_n11811);
assign 1_n9784 = ~1_n1364;
assign 1_n8923 = ~(1_n3441 ^ 1_n3277);
assign 1_n8372 = 1_n9421 | 1_n6732;
assign 1_n11866 = 1_n5801 & 1_n10408;
assign 1_n7350 = 1_n2733 | 1_n1272;
assign 1_n9909 = 1_n24 & 1_n1593;
assign 1_n13098 = 1_n3646 | 1_n6635;
assign 1_n10495 = 1_n8518 | 1_n11750;
assign 1_n4311 = ~(1_n729 ^ 1_n1071);
assign 1_n12227 = 1_n7363 | 1_n10;
assign 1_n5786 = 1_n10814 | 1_n2675;
assign 1_n9446 = ~(1_n6483 ^ 1_n8991);
assign 1_n8815 = 1_n8529 | 1_n8702;
assign 1_n8686 = ~(1_n2283 ^ 1_n3762);
assign 1_n6391 = 1_n8390 | 1_n2076;
assign 1_n6104 = ~(1_n9320 ^ 1_n10449);
assign 1_n7617 = ~(1_n67 ^ 1_n5587);
assign 1_n2317 = ~(1_n6468 ^ 1_n8599);
assign 1_n1874 = 1_n2279 | 1_n9126;
assign 1_n5558 = 1_n2346 | 1_n12695;
assign 1_n5992 = ~1_n10738;
assign 1_n11834 = ~(1_n1642 ^ 1_n12280);
assign 1_n9316 = 1_n2720 ^ 1_n12645;
assign 1_n9311 = ~1_n1405;
assign 1_n5000 = ~(1_n8710 ^ 1_n10933);
assign 1_n13024 = 1_n737 | 1_n8702;
assign 1_n8735 = ~(1_n5321 ^ 1_n6351);
assign 1_n6465 = 1_n3516 | 1_n3126;
assign 1_n4923 = 1_n10546 | 1_n4667;
assign 1_n11718 = 1_n3222 | 1_n4925;
assign 1_n786 = 1_n4758 & 1_n6420;
assign 1_n9453 = ~1_n12842;
assign 1_n11655 = 1_n12969 & 1_n12686;
assign 1_n2660 = ~1_n8867;
assign 1_n13168 = ~1_n4330;
assign 1_n270 = 1_n3241 & 1_n601;
assign 1_n4115 = ~(1_n1343 | 1_n11047);
assign 1_n2706 = ~(1_n3879 | 1_n4115);
assign 1_n13021 = ~1_n4074;
assign 1_n10838 = 1_n10762 & 1_n1675;
assign 1_n1853 = ~(1_n13162 | 1_n3883);
assign 1_n9154 = ~1_n8522;
assign 1_n738 = 1_n9029 & 1_n7679;
assign 1_n2588 = ~(1_n12161 ^ 1_n12455);
assign 1_n4396 = ~1_n4698;
assign 1_n10749 = 1_n12448 | 1_n7838;
assign 1_n4127 = ~(1_n5499 | 1_n5363);
assign 1_n8708 = 1_n6268 | 1_n4358;
assign 1_n186 = 1_n9792 & 1_n4995;
assign 1_n13053 = 1_n8508 & 1_n13235;
assign 1_n9680 = ~(1_n12928 ^ 1_n2247);
assign 1_n3111 = ~1_n2431;
assign 1_n8234 = ~1_n10763;
assign 1_n1097 = ~(1_n7716 ^ 1_n7103);
assign 1_n4092 = ~(1_n1968 ^ 1_n9572);
assign 1_n3331 = ~(1_n7286 | 1_n8798);
assign 1_n286 = 1_n3767 | 1_n11257;
assign 1_n11534 = ~(1_n5199 ^ 1_n2039);
assign 1_n10670 = 1_n6289 | 1_n1614;
assign 1_n611 = ~(1_n610 ^ 1_n1275);
assign 1_n7056 = 1_n3268 | 1_n6270;
assign 1_n8968 = ~(1_n120 | 1_n12028);
assign 1_n7573 = 1_n9627 | 1_n12195;
assign 1_n7356 = ~1_n9750;
assign 1_n11121 = ~1_n691;
assign 1_n8395 = ~(1_n1385 ^ 1_n10554);
assign 1_n11802 = ~(1_n13217 ^ 1_n6550);
assign 1_n8510 = ~1_n817;
assign 1_n446 = ~(1_n5075 ^ 1_n1430);
assign 1_n5518 = 1_n4473 | 1_n7935;
assign 1_n1914 = 1_n3273 | 1_n1780;
assign 1_n658 = ~(1_n2259 ^ 1_n949);
assign 1_n12302 = 1_n1933 & 1_n9407;
assign 1_n6205 = 1_n1783 | 1_n2958;
assign 1_n6183 = ~1_n4591;
assign 1_n512 = ~(1_n10645 | 1_n7583);
assign 1_n3285 = 1_n12598 & 1_n1003;
assign 1_n4515 = ~1_n9475;
assign 1_n11656 = ~(1_n1805 ^ 1_n8694);
assign 1_n10455 = 1_n3729 & 1_n11006;
assign 1_n7498 = 1_n596 | 1_n1825;
assign 1_n2984 = ~(1_n3009 ^ 1_n10488);
assign 1_n8412 = 1_n11858 | 1_n5873;
assign 1_n6334 = ~(1_n10335 ^ 1_n3966);
assign 1_n6548 = ~(1_n3188 ^ 1_n4002);
assign 1_n13207 = 1_n5360 | 1_n6601;
assign 1_n10903 = ~1_n4623;
assign 1_n7826 = ~(1_n5255 | 1_n10436);
assign 1_n9416 = 1_n9374 & 1_n3389;
assign 1_n12147 = ~(1_n1003 | 1_n12598);
assign 1_n11127 = 1_n4793 | 1_n10165;
assign 1_n4187 = ~1_n5827;
assign 1_n4592 = ~(1_n12532 ^ 1_n1330);
assign 1_n6513 = 1_n11975 & 1_n8408;
assign 1_n8356 = 1_n6689 | 1_n10049;
assign 1_n11661 = 1_n13 | 1_n2127;
assign 1_n8830 = ~(1_n329 ^ 1_n8479);
assign 1_n9663 = 1_n2791 ^ 1_n4138;
assign 1_n2097 = 1_n2205 & 1_n5095;
assign 1_n3358 = 1_n6808 & 1_n1289;
assign 1_n1268 = 1_n10768 & 1_n10154;
assign 1_n2154 = 1_n5872 & 1_n1170;
assign 1_n13215 = 1_n10895 | 1_n9014;
assign 1_n12077 = 1_n11060 & 1_n5633;
assign 1_n8596 = ~(1_n11903 ^ 1_n5765);
assign 1_n6798 = ~(1_n12805 ^ 1_n4);
assign 1_n3942 = ~(1_n3230 | 1_n10486);
assign 1_n6395 = ~(1_n277 ^ 1_n7050);
assign 1_n8316 = 1_n9668 | 1_n5242;
assign 1_n10797 = 1_n13011 ^ 1_n13219;
assign 1_n2099 = 1_n7037 & 1_n5337;
assign 1_n7348 = 1_n12109 | 1_n6732;
assign 1_n12374 = 1_n3243 | 1_n206;
assign 1_n9395 = 1_n8576 | 1_n8825;
assign 1_n10546 = ~(1_n3722 ^ 1_n3903);
assign 1_n7581 = ~(1_n13152 | 1_n5950);
assign 1_n7164 = 1_n12722 & 1_n2134;
assign 1_n1699 = 1_n11680 | 1_n2542;
assign 1_n3399 = 1_n8892 & 1_n4522;
assign 1_n2455 = ~1_n1774;
assign 1_n11289 = ~(1_n4853 ^ 1_n12337);
assign 1_n6877 = 1_n4584 | 1_n7723;
assign 1_n5632 = ~(1_n1865 ^ 1_n7922);
assign 1_n1340 = ~(1_n12855 ^ 1_n1670);
assign 1_n9863 = ~(1_n3471 | 1_n11287);
assign 1_n3397 = 1_n10830 | 1_n6265;
assign 1_n8105 = 1_n8759 | 1_n9075;
assign 1_n243 = 1_n9581 | 1_n8348;
assign 1_n3922 = 1_n1284 | 1_n10885;
assign 1_n9714 = 1_n9477 & 1_n12611;
assign 1_n6137 = 1_n7505 | 1_n8278;
assign 1_n2514 = 1_n4780 & 1_n10623;
assign 1_n8218 = 1_n2211 & 1_n7772;
assign 1_n12098 = 1_n7251 | 1_n9229;
assign 1_n1411 = ~(1_n11297 ^ 1_n4100);
assign 1_n11057 = ~(1_n2377 ^ 1_n2147);
assign 1_n4179 = ~1_n411;
assign 1_n3610 = ~(1_n11625 ^ 1_n12266);
assign 1_n8993 = 1_n12785 | 1_n12900;
assign 1_n3473 = 1_n6280 | 1_n742;
assign 1_n12290 = 1_n1113 | 1_n8030;
assign 1_n9387 = 1_n13181 | 1_n9444;
assign 1_n1472 = 1_n1035 | 1_n8702;
assign 1_n4848 = 1_n10223 | 1_n2082;
assign 1_n10403 = 1_n12105 & 1_n10129;
assign 1_n11853 = ~1_n11968;
assign 1_n12941 = 1_n11611 & 1_n3985;
assign 1_n5602 = 1_n5342 | 1_n2609;
assign 1_n8564 = ~(1_n390 ^ 1_n6328);
assign 1_n1653 = ~(1_n5757 ^ 1_n10119);
assign 1_n1715 = 1_n0 | 1_n8348;
assign 1_n4333 = ~1_n851;
assign 1_n10647 = ~(1_n2780 ^ 1_n7314);
assign 1_n9260 = ~(1_n5469 ^ 1_n8470);
assign 1_n3739 = 1_n8466 & 1_n5536;
assign 1_n2205 = ~(1_n10662 ^ 1_n8303);
assign 1_n1739 = 1_n12619 | 1_n5344;
assign 1_n6272 = ~(1_n6363 | 1_n6582);
assign 1_n10131 = ~1_n12845;
assign 1_n4584 = ~1_n11350;
assign 1_n7849 = ~(1_n11188 ^ 1_n7387);
assign 1_n6129 = ~1_n443;
assign 1_n2545 = ~1_n12267;
assign 1_n7051 = ~(1_n11275 ^ 1_n8459);
assign 1_n7687 = ~(1_n3327 ^ 1_n10729);
assign 1_n2729 = 1_n9842 & 1_n4275;
assign 1_n4331 = ~(1_n2721 ^ 1_n9343);
assign 1_n11187 = 1_n4166 | 1_n7530;
assign 1_n12889 = ~1_n11290;
assign 1_n10394 = ~(1_n3174 ^ 1_n10136);
assign 1_n10117 = ~1_n12005;
assign 1_n12330 = ~1_n11715;
assign 1_n11815 = ~1_n3378;
assign 1_n1089 = ~1_n3669;
assign 1_n3411 = 1_n6174 ^ 1_n4003;
assign 1_n7694 = 1_n6557 | 1_n13108;
assign 1_n7405 = ~(1_n11938 | 1_n6592);
assign 1_n6250 = ~1_n12651;
assign 1_n8858 = ~1_n5981;
assign 1_n2233 = ~(1_n5160 ^ 1_n6510);
assign 1_n583 = ~1_n962;
assign 1_n12201 = ~(1_n13138 ^ 1_n564);
assign 1_n5419 = ~(1_n12866 ^ 1_n9214);
assign 1_n7870 = ~(1_n5113 | 1_n9133);
assign 1_n12127 = ~(1_n3642 | 1_n11913);
assign 1_n8172 = ~(1_n8543 ^ 1_n582);
assign 1_n9608 = 1_n2786 & 1_n8972;
assign 1_n2654 = ~(1_n5095 ^ 1_n2917);
assign 1_n10933 = 1_n10301;
assign 1_n9073 = ~(1_n8507 ^ 1_n9852);
assign 1_n4617 = 1_n8006 | 1_n6178;
assign 1_n8152 = 1_n1200 & 1_n7645;
assign 1_n3276 = 1_n9451 & 1_n5366;
assign 1_n5120 = 1_n6755 | 1_n2556;
assign 1_n7381 = ~(1_n12147 | 1_n4733);
assign 1_n7555 = ~1_n3303;
assign 1_n9244 = 1_n12777 | 1_n1034;
assign 1_n8583 = ~(1_n11027 ^ 1_n11693);
assign 1_n5912 = ~(1_n739 ^ 1_n11488);
assign 1_n2408 = 1_n10208 & 1_n8683;
assign 1_n1167 = ~(1_n8512 ^ 1_n7658);
assign 1_n1937 = ~(1_n491 ^ 1_n9680);
assign 1_n6120 = ~1_n9893;
assign 1_n8791 = ~(1_n3785 ^ 1_n12185);
assign 1_n3185 = ~1_n11058;
assign 1_n6238 = ~1_n342;
assign 1_n12499 = ~(1_n10572 ^ 1_n2703);
assign 1_n12843 = 1_n1194 | 1_n206;
assign 1_n5601 = 1_n12102 | 1_n2197;
assign 1_n1894 = 1_n4811 & 1_n8787;
assign 1_n10028 = 1_n8355 & 1_n2663;
assign 1_n13033 = ~(1_n2644 | 1_n2803);
assign 1_n1585 = 1_n45 | 1_n9075;
assign 1_n268 = ~(1_n7564 ^ 1_n11415);
assign 1_n11836 = ~(1_n5293 ^ 1_n4409);
assign 1_n2504 = ~1_n12965;
assign 1_n7844 = 1_n11175 & 1_n6612;
assign 1_n9700 = 1_n8562 | 1_n1985;
assign 1_n7908 = ~1_n10538;
assign 1_n1180 = 1_n8391 & 1_n5762;
assign 1_n12855 = 1_n12483 | 1_n10573;
assign 1_n7323 = 1_n4293 ^ 1_n7877;
assign 1_n253 = 1_n9434 & 1_n3466;
assign 1_n11266 = 1_n3225 | 1_n4936;
assign 1_n9989 = 1_n7072 & 1_n12243;
assign 1_n3907 = 1_n8275 | 1_n11712;
assign 1_n2268 = 1_n2944 | 1_n7733;
assign 1_n5710 = 1_n5511 & 1_n7913;
assign 1_n5922 = 1_n6751 | 1_n5076;
assign 1_n4663 = 1_n6769 | 1_n2675;
assign 1_n10173 = 1_n9699 & 1_n1230;
assign 1_n11745 = ~1_n4086;
assign 1_n6086 = ~1_n9747;
assign 1_n3097 = 1_n5214 & 1_n9669;
assign 1_n12810 = ~(1_n568 ^ 1_n7246);
assign 1_n9485 = 1_n4750 | 1_n2460;
assign 1_n12169 = ~1_n1494;
assign 1_n2241 = ~(1_n5908 ^ 1_n11469);
assign 1_n7138 = ~(1_n3291 ^ 1_n9198);
assign 1_n10324 = 1_n11680 | 1_n11078;
assign 1_n7836 = 1_n2861 | 1_n1026;
assign 1_n12501 = 1_n9257;
assign 1_n9780 = 1_n6447 | 1_n5987;
assign 1_n12830 = 1_n8446 & 1_n6413;
assign 1_n12758 = ~1_n6023;
assign 1_n508 = 1_n4531 | 1_n12909;
assign 1_n4943 = 1_n10911 | 1_n2181;
assign 1_n9078 = 1_n1892 & 1_n1679;
assign 1_n5362 = ~(1_n1859 ^ 1_n7816);
assign 1_n8337 = 1_n9436 | 1_n3411;
assign 1_n13232 = ~(1_n1427 ^ 1_n5591);
assign 1_n12403 = ~1_n10207;
assign 1_n7080 = 1_n11015 & 1_n7955;
assign 1_n7745 = ~(1_n6170 ^ 1_n11181);
assign 1_n514 = ~(1_n1625 | 1_n1829);
assign 1_n2379 = 1_n4396 & 1_n6893;
assign 1_n8759 = ~1_n6826;
assign 1_n2249 = 1_n8685 & 1_n3780;
assign 1_n7250 = 1_n504 & 1_n7356;
assign 1_n2354 = 1_n11457 ^ 1_n5991;
assign 1_n2627 = 1_n4497 & 1_n8619;
assign 1_n3928 = ~1_n11734;
assign 1_n8640 = ~1_n7529;
assign 1_n13089 = 1_n10069 & 1_n5419;
assign 1_n3531 = ~1_n510;
assign 1_n8914 = 1_n8985 & 1_n6585;
assign 1_n11674 = 1_n10898 | 1_n12695;
assign 1_n9919 = ~1_n4335;
assign 1_n12115 = ~1_n10497;
assign 1_n4281 = ~(1_n4457 ^ 1_n4925);
assign 1_n7104 = 1_n1893 | 1_n1570;
assign 1_n3280 = 1_n7745 | 1_n418;
assign 1_n12106 = ~(1_n6812 ^ 1_n6548);
assign 1_n13026 = ~1_n12263;
assign 1_n1775 = 1_n8646 | 1_n6404;
assign 1_n3159 = 1_n121 | 1_n2890;
assign 1_n11849 = 1_n1835 | 1_n8509;
assign 1_n5760 = 1_n1700 | 1_n11045;
assign 1_n4754 = 1_n6743 | 1_n8702;
assign 1_n4809 = 1_n12039 & 1_n8245;
assign 1_n9156 = ~(1_n1760 ^ 1_n8451);
assign 1_n7299 = 1_n1601 | 1_n10508;
assign 1_n10295 = ~(1_n5846 ^ 1_n5597);
assign 1_n10420 = ~(1_n6342 | 1_n4093);
assign 1_n3700 = 1_n8428 | 1_n8530;
assign 1_n8765 = ~(1_n9845 ^ 1_n7800);
assign 1_n6167 = 1_n12629 | 1_n6732;
assign 1_n7536 = ~(1_n95 ^ 1_n4579);
assign 1_n9086 = 1_n11570 & 1_n4239;
assign 1_n10199 = 1_n4628 | 1_n12205;
assign 1_n12932 = 1_n9216 & 1_n10606;
assign 1_n6069 = ~(1_n9837 | 1_n7290);
assign 1_n2141 = ~1_n3631;
assign 1_n5990 = ~1_n8290;
assign 1_n372 = 1_n1281 | 1_n2672;
assign 1_n9565 = 1_n1857 & 1_n9096;
assign 1_n12914 = ~1_n4113;
assign 1_n1646 = 1_n2592 & 1_n497;
assign 1_n12728 = 1_n11920 | 1_n237;
assign 1_n8630 = ~1_n4325;
assign 1_n1958 = 1_n10894 & 1_n2503;
assign 1_n12869 = ~(1_n8157 | 1_n9086);
assign 1_n1188 = ~1_n11222;
assign 1_n7941 = ~(1_n7045 | 1_n4069);
assign 1_n8507 = ~(1_n7654 ^ 1_n8555);
assign 1_n5712 = 1_n390 & 1_n9439;
assign 1_n13234 = 1_n5013 | 1_n84;
assign 1_n2629 = ~(1_n3136 ^ 1_n587);
assign 1_n5340 = 1_n5528 & 1_n11377;
assign 1_n1950 = ~(1_n2603 ^ 1_n10224);
assign 1_n2953 = ~(1_n5192 ^ 1_n722);
assign 1_n4049 = ~(1_n7609 | 1_n11924);
assign 1_n10471 = ~1_n12965;
assign 1_n7416 = 1_n189 | 1_n5875;
assign 1_n8392 = ~1_n10594;
assign 1_n6545 = ~(1_n12880 | 1_n8478);
assign 1_n10815 = ~(1_n247 ^ 1_n7995);
assign 1_n8969 = 1_n4837 & 1_n6740;
assign 1_n4402 = 1_n11567 | 1_n7526;
assign 1_n10406 = ~(1_n335 ^ 1_n10349);
assign 1_n1424 = 1_n3965 | 1_n8941;
assign 1_n10839 = ~(1_n3579 ^ 1_n6998);
assign 1_n3008 = 1_n11236 & 1_n10408;
assign 1_n6307 = ~(1_n10415 ^ 1_n6415);
assign 1_n3437 = ~1_n10928;
assign 1_n12706 = ~(1_n7413 | 1_n8220);
assign 1_n13018 = ~(1_n5625 | 1_n9539);
assign 1_n3249 = ~(1_n12819 ^ 1_n7960);
assign 1_n11780 = 1_n2018 & 1_n411;
assign 1_n5148 = ~1_n10162;
assign 1_n9331 = 1_n2639 | 1_n2675;
assign 1_n6531 = ~(1_n6888 ^ 1_n4671);
assign 1_n2739 = ~(1_n6363 ^ 1_n2328);
assign 1_n5881 = 1_n4660 & 1_n6633;
assign 1_n1173 = 1_n12578 & 1_n7163;
assign 1_n964 = ~(1_n3939 ^ 1_n9006);
assign 1_n4984 = 1_n891 | 1_n1092;
assign 1_n12381 = ~(1_n10867 ^ 1_n10648);
assign 1_n2121 = ~(1_n8750 ^ 1_n12481);
assign 1_n2659 = ~(1_n12091 ^ 1_n9752);
assign 1_n6646 = ~(1_n5030 ^ 1_n11547);
assign 1_n5192 = ~(1_n4699 ^ 1_n13101);
assign 1_n3183 = 1_n6790 & 1_n10398;
assign 1_n2698 = 1_n7534 & 1_n7427;
assign 1_n9811 = ~(1_n4609 | 1_n2461);
assign 1_n1015 = 1_n1427 | 1_n5591;
assign 1_n1467 = 1_n2636 & 1_n7815;
assign 1_n8684 = 1_n3781 & 1_n9485;
assign 1_n7978 = ~(1_n3735 ^ 1_n8484);
assign 1_n10175 = 1_n9025 & 1_n11374;
assign 1_n5344 = 1_n252 & 1_n10429;
assign 1_n246 = ~(1_n4562 ^ 1_n1384);
assign 1_n2446 = ~1_n7012;
assign 1_n5624 = 1_n4657 | 1_n1605;
assign 1_n12025 = 1_n2228 | 1_n12604;
assign 1_n1599 = 1_n1438 | 1_n479;
assign 1_n1738 = 1_n10724 & 1_n9880;
assign 1_n572 = 1_n9723 | 1_n12501;
assign 1_n12384 = ~1_n5068;
assign 1_n4838 = ~(1_n4920 | 1_n6049);
assign 1_n5502 = ~1_n5477;
assign 1_n4160 = ~(1_n12276 | 1_n5244);
assign 1_n8869 = 1_n6977 & 1_n5007;
assign 1_n9755 = ~(1_n359 ^ 1_n7905);
assign 1_n3800 = ~1_n5570;
assign 1_n906 = ~1_n7569;
assign 1_n10059 = ~1_n3815;
assign 1_n4138 = ~(1_n7728 ^ 1_n12956);
assign 1_n32 = ~(1_n6212 ^ 1_n6406);
assign 1_n3537 = ~1_n1198;
assign 1_n2977 = 1_n5248 ^ 1_n1689;
assign 1_n10687 = ~(1_n6080 ^ 1_n3463);
assign 1_n3173 = ~1_n10482;
assign 1_n2051 = 1_n1029 & 1_n10252;
assign 1_n5163 = ~1_n1392;
assign 1_n1883 = ~1_n9915;
assign 1_n11514 = ~1_n4452;
assign 1_n6823 = 1_n10599 ^ 1_n5117;
assign 1_n11983 = 1_n11514 | 1_n7430;
assign 1_n10082 = ~(1_n47 ^ 1_n1728);
assign 1_n9418 = 1_n11020 & 1_n2727;
assign 1_n5546 = ~(1_n11719 ^ 1_n5629);
assign 1_n8081 = ~1_n4395;
assign 1_n1389 = ~1_n246;
assign 1_n785 = ~1_n12408;
assign 1_n6942 = ~1_n7285;
assign 1_n503 = 1_n3008 & 1_n9005;
assign 1_n9888 = ~1_n2062;
assign 1_n10132 = 1_n5588 | 1_n4640;
assign 1_n11282 = 1_n613 & 1_n4137;
assign 1_n11949 = ~(1_n1762 ^ 1_n11003);
assign 1_n8717 = 1_n4453 | 1_n3225;
assign 1_n724 = ~(1_n10873 ^ 1_n4512);
assign 1_n6520 = 1_n8020 | 1_n10179;
assign 1_n4779 = ~1_n9230;
assign 1_n4063 = ~1_n9732;
assign 1_n2618 = 1_n8033 & 1_n2949;
assign 1_n5620 = 1_n6524 & 1_n5380;
assign 1_n10344 = ~(1_n10064 ^ 1_n12549);
assign 1_n5785 = 1_n7683 & 1_n4592;
assign 1_n7386 = 1_n8966 | 1_n9689;
assign 1_n11389 = ~(1_n1278 ^ 1_n2031);
assign 1_n3718 = ~(1_n7794 ^ 1_n9114);
assign 1_n12444 = 1_n5146 | 1_n2958;
assign 1_n693 = 1_n5199 | 1_n2039;
assign 1_n8613 = ~1_n12936;
assign 1_n11092 = 1_n10439 | 1_n7530;
assign 1_n7492 = ~(1_n11776 ^ 1_n3290);
assign 1_n6720 = ~(1_n5907 | 1_n5785);
assign 1_n11710 = 1_n3616 | 1_n10179;
assign 1_n10182 = ~1_n1330;
assign 1_n5996 = 1_n8609 | 1_n9919;
assign 1_n10163 = 1_n11777 & 1_n10774;
assign 1_n4736 = 1_n371 | 1_n5186;
assign 1_n5282 = ~(1_n535 | 1_n8274);
assign 1_n12349 = 1_n12199 | 1_n9582;
assign 1_n8207 = 1_n1051 | 1_n5076;
assign 1_n1296 = ~1_n3815;
assign 1_n1926 = 1_n11212 | 1_n8702;
assign 1_n5445 = 1_n75 | 1_n4936;
assign 1_n10 = 1_n11768 & 1_n7836;
assign 1_n12441 = ~1_n1636;
assign 1_n12079 = ~(1_n11777 ^ 1_n12761);
assign 1_n2601 = 1_n2434 | 1_n2036;
assign 1_n9360 = ~(1_n4681 | 1_n1313);
assign 1_n11998 = 1_n6699 | 1_n6265;
assign 1_n6554 = ~(1_n2665 | 1_n4759);
assign 1_n5173 = 1_n6981 & 1_n1020;
assign 1_n3312 = 1_n673 & 1_n366;
assign 1_n170 = 1_n7350 & 1_n4180;
assign 1_n13055 = 1_n7213 & 1_n8961;
assign 1_n6096 = 1_n11557 & 1_n3375;
assign 1_n9288 = 1_n12122 | 1_n6091;
assign 1_n9837 = ~1_n336;
assign 1_n5748 = 1_n8778 | 1_n1999;
assign 1_n1935 = 1_n6219 & 1_n6734;
assign 1_n12911 = 1_n3225 | 1_n6404;
assign 1_n8676 = 1_n6810 | 1_n10871;
assign 1_n4594 = 1_n2018 & 1_n13058;
assign 1_n10331 = ~1_n13064;
assign 1_n8066 = 1_n12349 & 1_n8444;
assign 1_n11173 = 1_n1850 & 1_n8882;
assign 1_n1647 = 1_n4999 | 1_n5652;
assign 1_n1166 = ~(1_n6712 | 1_n6578);
assign 1_n1911 = ~(1_n11024 ^ 1_n3156);
assign 1_n5913 = ~(1_n5228 ^ 1_n3330);
assign 1_n10019 = 1_n1431 & 1_n10856;
assign 1_n11005 = 1_n11929 | 1_n9268;
assign 1_n10999 = 1_n6063 | 1_n1463;
assign 1_n7551 = 1_n1305 & 1_n747;
assign 1_n8726 = 1_n7134 | 1_n8247;
assign 1_n6647 = ~(1_n5584 ^ 1_n825);
assign 1_n11216 = ~(1_n7836 ^ 1_n11768);
assign 1_n9448 = 1_n909 & 1_n4805;
assign 1_n6619 = ~(1_n5702 ^ 1_n12201);
assign 1_n7802 = ~(1_n8549 ^ 1_n5804);
assign 1_n7779 = 1_n11559 ^ 1_n8542;
assign 1_n5225 = ~(1_n9037 | 1_n7599);
assign 1_n9286 = ~1_n7;
assign 1_n1919 = ~1_n8290;
assign 1_n2661 = 1_n7741 | 1_n9159;
assign 1_n11213 = 1_n718 | 1_n12862;
assign 1_n12168 = 1_n5565 | 1_n1144;
assign 1_n7359 = ~(1_n13031 ^ 1_n3073);
assign 1_n6747 = ~(1_n8 ^ 1_n4401);
assign 1_n9277 = 1_n1325 | 1_n3825;
assign 1_n5740 = ~1_n8139;
assign 1_n11571 = 1_n7819 | 1_n2449;
assign 1_n9560 = ~(1_n10431 ^ 1_n9299);
assign 1_n6761 = ~(1_n2518 | 1_n5331);
assign 1_n8544 = ~(1_n5185 ^ 1_n9650);
assign 1_n2957 = ~(1_n5072 ^ 1_n9289);
assign 1_n6446 = 1_n10411 | 1_n11239;
assign 1_n2074 = 1_n6447 & 1_n5987;
assign 1_n6988 = ~1_n10657;
assign 1_n11864 = ~1_n3832;
assign 1_n1187 = 1_n6180 & 1_n1862;
assign 1_n8217 = ~(1_n11464 ^ 1_n11651);
assign 1_n4034 = 1_n11094 | 1_n4936;
assign 1_n2929 = ~(1_n10630 ^ 1_n2690);
assign 1_n5153 = 1_n11648 | 1_n8805;
assign 1_n7517 = 1_n6749 | 1_n2943;
assign 1_n11736 = ~(1_n12312 ^ 1_n12239);
assign 1_n10722 = ~(1_n223 ^ 1_n1590);
assign 1_n7873 = 1_n8915 & 1_n12012;
assign 1_n4897 = ~(1_n9138 ^ 1_n11254);
assign 1_n8565 = 1_n12254 | 1_n4230;
assign 1_n9530 = ~(1_n13171 ^ 1_n7536);
assign 1_n1870 = ~(1_n2388 ^ 1_n4186);
assign 1_n4499 = ~1_n5603;
assign 1_n5728 = ~(1_n13196 ^ 1_n4727);
assign 1_n3506 = 1_n1328 & 1_n6741;
assign 1_n12354 = 1_n6173 | 1_n4116;
assign 1_n8650 = ~1_n7725;
assign 1_n3594 = ~(1_n5324 ^ 1_n3074);
assign 1_n12773 = 1_n9580 | 1_n486;
assign 1_n5995 = 1_n5449 & 1_n5855;
assign 1_n593 = 1_n10351 | 1_n8448;
assign 1_n8124 = ~(1_n9247 ^ 1_n2979);
assign 1_n11719 = ~(1_n6926 ^ 1_n746);
assign 1_n5964 = 1_n6901 | 1_n11670;
assign 1_n10252 = 1_n745 | 1_n982;
assign 1_n4843 = ~(1_n1932 ^ 1_n7850);
assign 1_n10827 = ~(1_n3708 ^ 1_n5496);
assign 1_n12986 = ~1_n8520;
assign 1_n7545 = 1_n6086 | 1_n5076;
assign 1_n7921 = 1_n7862 | 1_n9861;
assign 1_n11096 = 1_n2416 | 1_n8348;
assign 1_n12864 = ~(1_n9878 | 1_n3030);
assign 1_n5096 = 1_n10147 & 1_n2564;
assign 1_n7445 = ~(1_n5431 ^ 1_n4429);
assign 1_n1254 = 1_n8183 & 1_n854;
assign 1_n6901 = 1_n8953 & 1_n3880;
assign 1_n9384 = 1_n10509 | 1_n11928;
assign 1_n9600 = 1_n5233 | 1_n9579;
assign 1_n7726 = ~(1_n3161 ^ 1_n251);
assign 1_n8177 = 1_n6492 | 1_n11464;
assign 1_n3344 = ~1_n10162;
assign 1_n12670 = 1_n12615 & 1_n7667;
assign 1_n2119 = ~(1_n4187 ^ 1_n2216);
assign 1_n3152 = ~(1_n6607 ^ 1_n7116);
assign 1_n12087 = 1_n2194 & 1_n5109;
assign 1_n11548 = ~1_n9093;
assign 1_n6479 = 1_n10798 | 1_n10179;
assign 1_n4787 = 1_n8264 & 1_n10834;
assign 1_n8443 = 1_n12894 | 1_n2969;
assign 1_n3988 = ~(1_n12652 ^ 1_n10076);
assign 1_n6351 = ~(1_n615 ^ 1_n8386);
assign 1_n11228 = 1_n3928 | 1_n12501;
assign 1_n4882 = ~(1_n3886 ^ 1_n8899);
assign 1_n1630 = 1_n2823 | 1_n566;
assign 1_n8959 = 1_n11761 | 1_n6874;
assign 1_n12223 = ~(1_n5615 | 1_n805);
assign 1_n11134 = ~(1_n3006 ^ 1_n5568);
assign 1_n12468 = ~(1_n5616 ^ 1_n5332);
assign 1_n6059 = ~(1_n11203 ^ 1_n3926);
assign 1_n2265 = 1_n11084 | 1_n3479;
assign 1_n10489 = 1_n5923 | 1_n8188;
assign 1_n8082 = ~1_n2295;
assign 1_n8283 = ~(1_n2437 ^ 1_n691);
assign 1_n6553 = ~(1_n1450 ^ 1_n703);
assign 1_n8996 = 1_n3903 & 1_n3722;
assign 1_n2736 = ~(1_n2137 ^ 1_n342);
assign 1_n5738 = 1_n9019 | 1_n8348;
assign 1_n7854 = 1_n5671 & 1_n4335;
assign 1_n5333 = 1_n11745 & 1_n1920;
assign 1_n1133 = 1_n13127 & 1_n452;
assign 1_n11614 = ~1_n6857;
assign 1_n13159 = ~1_n6818;
assign 1_n10055 = ~(1_n9384 ^ 1_n2401);
assign 1_n7945 = ~1_n12391;
assign 1_n5771 = 1_n5544 | 1_n3372;
assign 1_n10150 = 1_n2062 ^ 1_n6394;
assign 1_n1400 = 1_n11928 | 1_n2958;
assign 1_n14 = 1_n6672 | 1_n1043;
assign 1_n8321 = 1_n1997 & 1_n4054;
assign 1_n11434 = 1_n11324 & 1_n12284;
assign 1_n5501 = ~(1_n2536 ^ 1_n982);
assign 1_n9675 = ~1_n353;
assign 1_n3286 = 1_n629 & 1_n5153;
assign 1_n901 = ~(1_n7545 ^ 1_n4276);
assign 1_n5549 = ~(1_n2569 ^ 1_n4590);
assign 1_n5137 = ~(1_n3974 ^ 1_n11906);
assign 1_n13032 = 1_n1009 & 1_n8296;
assign 1_n6478 = 1_n9032 & 1_n3235;
assign 1_n6624 = ~(1_n9190 ^ 1_n9503);
assign 1_n8185 = 1_n9776 | 1_n8587;
assign 1_n8238 = ~(1_n6513 | 1_n2475);
assign 1_n6771 = ~(1_n6310 ^ 1_n9950);
assign 1_n296 = ~(1_n12649 ^ 1_n11983);
assign 1_n7942 = ~1_n2043;
assign 1_n1124 = ~(1_n5649 | 1_n8695);
assign 1_n2655 = 1_n10168 & 1_n3832;
assign 1_n4286 = 1_n3413 & 1_n9708;
assign 1_n2833 = 1_n3062 | 1_n542;
assign 1_n4169 = 1_n4133 & 1_n11915;
assign 1_n5250 = 1_n2688 | 1_n6265;
assign 1_n5458 = ~(1_n3683 ^ 1_n9832);
assign 1_n5817 = 1_n12077 & 1_n5125;
assign 1_n12321 = 1_n9474 ^ 1_n11854;
assign 1_n8383 = ~1_n2771;
assign 1_n1345 = ~1_n2758;
assign 1_n4365 = 1_n304 | 1_n10079;
assign 1_n5044 = 1_n13075 & 1_n2390;
assign 1_n11696 = ~1_n12560;
assign 1_n5848 = 1_n6543 & 1_n13187;
assign 1_n12121 = ~(1_n8242 ^ 1_n10209);
assign 1_n991 = ~1_n12306;
assign 1_n9865 = ~(1_n8238 | 1_n725);
assign 1_n6273 = 1_n4888 & 1_n6579;
assign 1_n3221 = ~(1_n8989 | 1_n3);
assign 1_n6084 = 1_n4462 | 1_n8702;
assign 1_n3049 = ~1_n9732;
assign 1_n1559 = 1_n10481 | 1_n8563;
assign 1_n3799 = 1_n3795 & 1_n1736;
assign 1_n2448 = 1_n11105 & 1_n9355;
assign 1_n7791 = ~1_n3029;
assign 1_n9969 = 1_n4536 | 1_n10057;
assign 1_n2677 = 1_n7291 | 1_n5076;
assign 1_n6600 = ~(1_n11587 ^ 1_n2684);
assign 1_n10605 = 1_n12235 & 1_n12204;
assign 1_n11784 = ~1_n4703;
assign 1_n12935 = 1_n10950 | 1_n8268;
assign 1_n564 = 1_n3867 & 1_n442;
assign 1_n12420 = ~(1_n11501 | 1_n7630);
assign 1_n1011 = 1_n536 | 1_n6834;
assign 1_n8206 = ~1_n5962;
assign 1_n1137 = 1_n1428 & 1_n9191;
assign 1_n1736 = 1_n5447 | 1_n4861;
assign 1_n1036 = ~(1_n9958 ^ 1_n12461);
assign 1_n11951 = 1_n4716 | 1_n6055;
assign 1_n1131 = 1_n2449 | 1_n7935;
assign 1_n5006 = ~(1_n11774 | 1_n3828);
assign 1_n2166 = ~1_n4709;
assign 1_n10343 = 1_n7342;
assign 1_n7282 = ~(1_n434 ^ 1_n3787);
assign 1_n2131 = ~1_n8535;
assign 1_n12888 = 1_n3265 | 1_n2188;
assign 1_n2443 = ~1_n11553;
assign 1_n9304 = 1_n1484 | 1_n3432;
assign 1_n4077 = ~1_n3769;
assign 1_n12222 = 1_n3459 | 1_n3225;
assign 1_n4367 = ~(1_n12764 ^ 1_n7319);
assign 1_n853 = ~(1_n1523 | 1_n9002);
assign 1_n4364 = 1_n6803 | 1_n8763;
assign 1_n983 = 1_n1876 ^ 1_n9303;
assign 1_n683 = ~1_n7061;
assign 1_n1021 = 1_n8308 & 1_n3409;
assign 1_n5493 = ~(1_n11184 ^ 1_n8258);
assign 1_n12754 = 1_n6769 | 1_n1570;
assign 1_n4544 = 1_n13080 | 1_n4337;
assign 1_n12731 = ~(1_n9004 ^ 1_n11735);
assign 1_n6118 = ~(1_n970 ^ 1_n997);
assign 1_n12380 = ~1_n11814;
assign 1_n12955 = ~1_n103;
assign 1_n10635 = ~(1_n6929 ^ 1_n12664);
assign 1_n2776 = ~(1_n163 ^ 1_n3065);
assign 1_n4870 = 1_n5238 & 1_n5350;
assign 1_n4159 = 1_n10270 | 1_n9595;
assign 1_n10070 = ~(1_n3603 ^ 1_n1622);
assign 1_n2418 = ~(1_n9792 ^ 1_n11428);
assign 1_n7042 = 1_n5547 | 1_n3981;
assign 1_n7583 = 1_n1480 | 1_n905;
assign 1_n9065 = ~(1_n3477 ^ 1_n7861);
assign 1_n9550 = ~(1_n10834 ^ 1_n8264);
assign 1_n1308 = ~1_n13044;
assign 1_n9901 = ~(1_n4830 ^ 1_n10541);
assign 1_n715 = ~1_n11396;
assign 1_n10822 = 1_n3288 | 1_n5291;
assign 1_n962 = 1_n8840 & 1_n13157;
assign 1_n10299 = ~(1_n6574 | 1_n7614);
assign 1_n4088 = 1_n6960 | 1_n4723;
assign 1_n743 = ~(1_n11585 ^ 1_n12094);
assign 1_n8305 = 1_n9060 & 1_n8722;
assign 1_n10041 = ~1_n2535;
assign 1_n9000 = ~(1_n12411 ^ 1_n4745);
assign 1_n11179 = ~(1_n2896 ^ 1_n1061);
assign 1_n1234 = 1_n5973 | 1_n9075;
assign 1_n7955 = 1_n12481 | 1_n8750;
assign 1_n5054 = 1_n3296 | 1_n3114;
assign 1_n9562 = ~(1_n1827 | 1_n13059);
assign 1_n716 = 1_n9144 & 1_n6870;
assign 1_n1638 = ~1_n5729;
assign 1_n2463 = ~1_n12289;
assign 1_n10537 = 1_n2045 & 1_n1032;
assign 1_n9983 = ~(1_n4152 ^ 1_n2159);
assign 1_n10959 = 1_n511 | 1_n12162;
assign 1_n6613 = ~(1_n2495 | 1_n2026);
assign 1_n1526 = ~1_n2813;
assign 1_n12 = ~(1_n6593 ^ 1_n2511);
assign 1_n4719 = 1_n3040 ^ 1_n7761;
assign 1_n12276 = ~(1_n7898 ^ 1_n11285);
assign 1_n12174 = ~1_n6392;
assign 1_n1974 = ~(1_n12736 ^ 1_n1994);
assign 1_n9583 = ~(1_n1304 ^ 1_n4718);
assign 1_n1506 = 1_n12348 & 1_n469;
assign 1_n2484 = ~1_n10594;
assign 1_n5515 = 1_n5138 & 1_n8784;
assign 1_n3469 = 1_n8324 | 1_n8702;
assign 1_n10523 = ~(1_n9914 ^ 1_n697);
assign 1_n8148 = 1_n3070 | 1_n4930;
assign 1_n8943 = 1_n6156 | 1_n10207;
assign 1_n9699 = 1_n1011 & 1_n3350;
assign 1_n4675 = ~(1_n2010 | 1_n10661);
assign 1_n12452 = 1_n7608 | 1_n12388;
assign 1_n1017 = ~1_n5881;
assign 1_n7527 = ~(1_n3846 ^ 1_n6277);
assign 1_n10392 = 1_n6209 ^ 1_n11084;
assign 1_n5286 = ~1_n7573;
assign 1_n5 = ~1_n11511;
assign 1_n9335 = ~(1_n3988 | 1_n2445);
assign 1_n6615 = 1_n12390 & 1_n1075;
assign 1_n6502 = 1_n10150 | 1_n9512;
assign 1_n10167 = ~(1_n10746 ^ 1_n4712);
assign 1_n6634 = 1_n2230 | 1_n12120;
assign 1_n7574 = ~(1_n4391 ^ 1_n6102);
assign 1_n11351 = 1_n3420 & 1_n6123;
assign 1_n2495 = 1_n6755 | 1_n8374;
assign 1_n5621 = ~(1_n5391 ^ 1_n9231);
assign 1_n4819 = 1_n7947 & 1_n12601;
assign 1_n2862 = 1_n9484 | 1_n2842;
assign 1_n11598 = ~(1_n7227 ^ 1_n5231);
assign 1_n3201 = ~1_n7713;
assign 1_n3740 = ~(1_n11688 ^ 1_n5374);
assign 1_n2157 = ~1_n11692;
assign 1_n3855 = ~(1_n8331 | 1_n798);
assign 1_n1311 = 1_n2933 | 1_n13225;
assign 1_n3770 = 1_n2041 | 1_n1144;
assign 1_n1740 = 1_n787 | 1_n4947;
assign 1_n10705 = ~(1_n1321 | 1_n3144);
assign 1_n3383 = ~(1_n6107 | 1_n9988);
assign 1_n12008 = ~(1_n4754 | 1_n3533);
assign 1_n8743 = 1_n11291 | 1_n1026;
assign 1_n12365 = 1_n4227 | 1_n3418;
assign 1_n1790 = 1_n8469 ^ 1_n9473;
assign 1_n1274 = 1_n4308 | 1_n3820;
assign 1_n5904 = 1_n9659 | 1_n395;
assign 1_n702 = 1_n8234 & 1_n10820;
assign 1_n2743 = ~(1_n6153 ^ 1_n2392);
assign 1_n9830 = 1_n5079 | 1_n8030;
assign 1_n9149 = 1_n1158 & 1_n1713;
assign 1_n633 = ~1_n5309;
assign 1_n11022 = 1_n361 | 1_n3039;
assign 1_n265 = 1_n3847 & 1_n10065;
assign 1_n11048 = ~(1_n12458 ^ 1_n1151);
assign 1_n4771 = 1_n1919 | 1_n8348;
assign 1_n2843 = ~(1_n11720 ^ 1_n4045);
assign 1_n10565 = ~1_n8092;
assign 1_n7485 = ~1_n8518;
assign 1_n2757 = ~1_n9732;
assign 1_n4655 = ~1_n3188;
assign 1_n10485 = 1_n7040 ^ 1_n3763;
assign 1_n106 = ~(1_n9592 | 1_n2668);
assign 1_n3347 = ~(1_n9209 | 1_n6528);
assign 1_n6792 = ~(1_n3749 | 1_n46);
assign 1_n538 = 1_n1141 | 1_n8937;
assign 1_n773 = ~(1_n172 ^ 1_n4973);
assign 1_n5818 = 1_n4456 | 1_n5353;
assign 1_n8651 = ~(1_n3558 ^ 1_n11766);
assign 1_n12719 = ~(1_n9138 | 1_n11254);
assign 1_n3546 = ~(1_n8867 | 1_n9827);
assign 1_n520 = ~(1_n3236 ^ 1_n9197);
assign 1_n10935 = 1_n1102 & 1_n11908;
assign 1_n531 = ~(1_n12135 ^ 1_n6714);
assign 1_n2852 = ~(1_n11881 ^ 1_n6991);
assign 1_n5505 = 1_n146 & 1_n95;
assign 1_n1776 = ~(1_n12056 ^ 1_n446);
assign 1_n9735 = 1_n9152 & 1_n6457;
assign 1_n7160 = ~(1_n12949 ^ 1_n8818);
assign 1_n9561 = ~(1_n9220 | 1_n8333);
assign 1_n1149 = ~(1_n9496 ^ 1_n8034);
assign 1_n3580 = 1_n2838 & 1_n2388;
assign 1_n1482 = 1_n646 & 1_n47;
assign 1_n6965 = ~(1_n11279 ^ 1_n11454);
assign 1_n601 = ~(1_n8241 ^ 1_n7462);
assign 1_n5535 = 1_n3311 & 1_n10606;
assign 1_n10381 = ~1_n8284;
assign 1_n8248 = ~1_n9825;
assign 1_n4039 = ~(1_n5655 ^ 1_n2206);
assign 1_n10629 = ~(1_n4199 | 1_n6938);
assign 1_n12275 = ~(1_n2173 ^ 1_n3490);
assign 1_n5465 = 1_n5433 | 1_n4230;
assign 1_n10212 = 1_n12832 | 1_n1690;
assign 1_n9970 = 1_n9723 | 1_n10871;
assign 1_n3608 = ~(1_n4026 | 1_n1243);
assign 1_n1168 = ~1_n10162;
assign 1_n8144 = ~(1_n7578 ^ 1_n6775);
assign 1_n12845 = ~(1_n264 ^ 1_n6500);
assign 1_n10682 = 1_n856 | 1_n8602;
assign 1_n11487 = 1_n5226 | 1_n8024;
assign 1_n11077 = ~(1_n5073 ^ 1_n12962);
assign 1_n9098 = 1_n2932 & 1_n11182;
assign 1_n3708 = 1_n2346 | 1_n8348;
assign 1_n6490 = 1_n9066 | 1_n7681;
assign 1_n10566 = 1_n9444 | 1_n4373;
assign 1_n13047 = ~(1_n11338 ^ 1_n6609);
assign 1_n3650 = 1_n9864 & 1_n4224;
assign 1_n8702 = 1_n4013;
assign 1_n12291 = ~(1_n6583 ^ 1_n1142);
assign 1_n9855 = 1_n7673 & 1_n1223;
assign 1_n5335 = 1_n11404 | 1_n12273;
assign 1_n9325 = ~1_n8827;
assign 1_n6223 = ~1_n4006;
assign 1_n5750 = 1_n11969 & 1_n4560;
assign 1_n6076 = 1_n10220 | 1_n12215;
assign 1_n1004 = 1_n570 & 1_n3366;
assign 1_n8295 = ~1_n11017;
assign 1_n2005 = 1_n7828 & 1_n3888;
assign 1_n12067 = ~(1_n7734 ^ 1_n1374);
assign 1_n2040 = ~(1_n11722 ^ 1_n7502);
assign 1_n12615 = ~1_n12961;
assign 1_n487 = 1_n2590 & 1_n7720;
assign 1_n1120 = ~(1_n10160 ^ 1_n10625);
assign 1_n4734 = ~(1_n4094 ^ 1_n5323);
assign 1_n4869 = 1_n3095 | 1_n2983;
assign 1_n9653 = 1_n3480 | 1_n3119;
assign 1_n8023 = ~(1_n8801 ^ 1_n12509);
assign 1_n5110 = ~(1_n11456 ^ 1_n7589);
assign 1_n7070 = ~(1_n2065 ^ 1_n1565);
assign 1_n9458 = ~(1_n8547 ^ 1_n416);
assign 1_n10500 = 1_n5782 | 1_n10319;
assign 1_n3883 = 1_n12270 & 1_n12076;
assign 1_n1726 = ~(1_n6372 ^ 1_n10624);
assign 1_n806 = ~(1_n271 ^ 1_n12647);
assign 1_n1170 = 1_n5105 | 1_n8505;
assign 1_n1691 = 1_n385 | 1_n13056;
assign 1_n6964 = ~(1_n2564 ^ 1_n10147);
assign 1_n4393 = 1_n7748 | 1_n2133;
assign 1_n12589 = 1_n12705 & 1_n9051;
assign 1_n9825 = ~(1_n2677 ^ 1_n6708);
assign 1_n687 = ~(1_n2886 ^ 1_n8854);
assign 1_n3275 = 1_n9559 | 1_n4690;
assign 1_n9045 = ~(1_n5439 | 1_n10315);
assign 1_n6477 = ~(1_n1509 ^ 1_n2563);
assign 1_n1606 = 1_n10498 | 1_n10889;
assign 1_n5534 = ~(1_n8825 ^ 1_n8576);
assign 1_n5857 = ~(1_n9625 ^ 1_n12950);
assign 1_n602 = ~1_n2824;
assign 1_n2093 = ~(1_n6697 ^ 1_n1842);
assign 1_n5603 = 1_n8941 | 1_n5797;
assign 1_n13078 = 1_n840 & 1_n6667;
assign 1_n427 = 1_n3006 & 1_n4470;
assign 1_n12813 = ~1_n11897;
assign 1_n4789 = 1_n8940 & 1_n11222;
assign 1_n8028 = 1_n9761 | 1_n1570;
assign 1_n4305 = ~1_n10111;
assign 1_n8346 = 1_n9502 | 1_n2719;
assign 1_n3760 = 1_n10908 & 1_n10408;
assign 1_n11102 = ~(1_n6426 ^ 1_n5032);
assign 1_n6616 = ~(1_n109 ^ 1_n3287);
assign 1_n3232 = ~1_n62;
assign 1_n126 = 1_n2488 | 1_n793;
assign 1_n7227 = 1_n2825 | 1_n6404;
assign 1_n4068 = ~(1_n9630 | 1_n12359);
assign 1_n12253 = 1_n3333 | 1_n6715;
assign 1_n4102 = 1_n1978 ^ 1_n3168;
assign 1_n10977 = ~1_n2174;
assign 1_n11673 = 1_n11236 & 1_n854;
assign 1_n9923 = ~(1_n12389 | 1_n7539);
assign 1_n3930 = ~(1_n11913 ^ 1_n8409);
assign 1_n3896 = ~(1_n10969 ^ 1_n2843);
assign 1_n9628 = 1_n2625 | 1_n4386;
assign 1_n9754 = ~(1_n7833 | 1_n791);
assign 1_n2209 = 1_n12141 & 1_n10513;
assign 1_n3630 = ~1_n22;
assign 1_n3655 = ~1_n3123;
assign 1_n5705 = 1_n8817 | 1_n10106;
assign 1_n10391 = 1_n898 | 1_n4154;
assign 1_n4959 = 1_n2860 & 1_n10125;
assign 1_n1062 = 1_n6038 | 1_n1468;
assign 1_n1707 = ~(1_n9248 ^ 1_n6872);
assign 1_n1384 = ~(1_n7201 ^ 1_n11337);
assign 1_n2226 = ~1_n12605;
assign 1_n7283 = ~1_n1307;
assign 1_n8370 = 1_n2444 | 1_n11461;
assign 1_n2114 = 1_n11094 | 1_n7530;
assign 1_n6442 = 1_n1452 & 1_n5503;
assign 1_n13030 = ~(1_n4097 | 1_n12876);
assign 1_n12279 = ~(1_n6573 ^ 1_n9671);
assign 1_n9420 = 1_n3974 | 1_n9018;
assign 1_n5353 = 1_n8498 | 1_n4373;
assign 1_n8609 = ~1_n11061;
assign 1_n9737 = 1_n6024 & 1_n4915;
assign 1_n9340 = ~1_n13161;
assign 1_n8439 = ~(1_n11444 | 1_n12430);
assign 1_n5850 = 1_n9679 | 1_n9118;
assign 1_n5894 = ~(1_n11332 ^ 1_n4240);
assign 1_n11586 = ~(1_n10316 ^ 1_n12022);
assign 1_n12772 = ~1_n4293;
assign 1_n11126 = ~(1_n7796 ^ 1_n4829);
assign 1_n3391 = ~(1_n6778 ^ 1_n12110);
assign 1_n187 = ~(1_n11005 ^ 1_n1896);
assign 1_n8849 = ~1_n12482;
assign 1_n6969 = ~(1_n155 ^ 1_n9806);
assign 1_n9440 = ~(1_n8536 ^ 1_n3896);
assign 1_n9346 = 1_n3425 | 1_n1028;
assign 1_n11645 = 1_n2888 & 1_n3764;
assign 1_n10697 = 1_n5483 & 1_n6889;
assign 1_n1553 = 1_n583 | 1_n11405;
assign 1_n2927 = 1_n12022 & 1_n10316;
assign 1_n2594 = ~(1_n691 | 1_n1874);
assign 1_n8196 = 1_n1751 & 1_n9801;
assign 1_n1924 = ~(1_n10054 | 1_n10651);
assign 1_n1386 = ~(1_n9944 ^ 1_n1898);
assign 1_n8696 = 1_n8124 & 1_n4262;
assign 1_n10743 = ~(1_n6943 ^ 1_n7030);
assign 1_n9823 = ~(1_n12021 ^ 1_n11695);
assign 1_n4915 = 1_n7597 | 1_n6732;
assign 1_n596 = 1_n10286 | 1_n6944;
assign 1_n6305 = 1_n10898 | 1_n12847;
assign 1_n11095 = 1_n9400 | 1_n8030;
assign 1_n18 = ~1_n4357;
assign 1_n3566 = 1_n13096 & 1_n6146;
assign 1_n11566 = 1_n8431 | 1_n12666;
assign 1_n2116 = 1_n7891 & 1_n8048;
assign 1_n9574 = ~(1_n6513 ^ 1_n725);
assign 1_n9734 = ~(1_n3964 | 1_n6879);
assign 1_n3453 = 1_n0 | 1_n4230;
assign 1_n1430 = 1_n6444 & 1_n11489;
assign 1_n12178 = 1_n11171 | 1_n12847;
assign 1_n8280 = ~1_n4368;
assign 1_n10241 = 1_n12312 | 1_n12781;
assign 1_n3925 = ~(1_n4953 ^ 1_n8119);
assign 1_n556 = ~(1_n8313 ^ 1_n1715);
assign 1_n13051 = ~1_n9669;
assign 1_n10232 = 1_n7677 | 1_n12048;
assign 1_n1044 = 1_n11951 & 1_n11936;
assign 1_n2985 = 1_n4690 & 1_n9559;
assign 1_n7397 = ~(1_n11875 ^ 1_n11755);
assign 1_n6575 = ~1_n4695;
assign 1_n5371 = 1_n1183 & 1_n7747;
assign 1_n6134 = ~(1_n8867 ^ 1_n2382);
assign 1_n10813 = 1_n8208 & 1_n12375;
assign 1_n4548 = ~(1_n2208 ^ 1_n3402);
assign 1_n9512 = ~1_n2334;
assign 1_n3393 = 1_n4655 | 1_n6924;
assign 1_n8049 = ~(1_n10878 ^ 1_n8308);
assign 1_n361 = 1_n1510 & 1_n12816;
assign 1_n2008 = 1_n8090 | 1_n11282;
assign 1_n8225 = ~1_n5729;
assign 1_n8924 = 1_n4967 | 1_n3981;
assign 1_n3567 = 1_n1499 & 1_n1210;
assign 1_n11427 = ~1_n12937;
assign 1_n4348 = 1_n12003 & 1_n11109;
assign 1_n9201 = ~(1_n6131 ^ 1_n9757);
assign 1_n4684 = 1_n4977 & 1_n6864;
assign 1_n3644 = 1_n12920 & 1_n9727;
assign 1_n7695 = 1_n12477 | 1_n8231;
assign 1_n3586 = ~1_n3263;
assign 1_n9429 = ~1_n9528;
assign 1_n36 = 1_n3049 | 1_n5264;
assign 1_n473 = ~1_n4459;
assign 1_n7125 = 1_n11588 | 1_n8748;
assign 1_n12247 = ~(1_n7671 | 1_n8078);
assign 1_n430 = 1_n10138 | 1_n9386;
assign 1_n3289 = ~(1_n8944 ^ 1_n6567);
assign 1_n2803 = 1_n7650 & 1_n3657;
assign 1_n6329 = 1_n345 | 1_n1961;
assign 1_n1590 = ~(1_n10294 ^ 1_n13222);
assign 1_n4051 = ~(1_n10992 ^ 1_n8015);
assign 1_n7600 = 1_n3564 | 1_n10029;
assign 1_n8554 = ~(1_n3204 ^ 1_n4729);
assign 1_n4699 = ~(1_n7161 | 1_n8030);
assign 1_n11704 = 1_n2262 | 1_n4865;
assign 1_n290 = ~1_n5457;
assign 1_n6366 = ~1_n3625;
assign 1_n10699 = ~(1_n4086 ^ 1_n1920);
assign 1_n2026 = 1_n889 & 1_n7897;
assign 1_n1329 = ~1_n11429;
assign 1_n1451 = ~1_n9906;
assign 1_n3318 = ~1_n6604;
assign 1_n763 = ~(1_n1170 ^ 1_n5872);
assign 1_n2196 = ~(1_n5128 ^ 1_n6200);
assign 1_n2783 = 1_n987 | 1_n10319;
assign 1_n2039 = ~(1_n4467 ^ 1_n12142);
assign 1_n482 = ~1_n2777;
assign 1_n6865 = ~(1_n346 ^ 1_n5755);
assign 1_n2528 = 1_n3726 | 1_n2133;
assign 1_n3494 = ~(1_n8476 ^ 1_n10689);
assign 1_n788 = ~(1_n9892 ^ 1_n10526);
assign 1_n3756 = ~(1_n13 ^ 1_n11687);
assign 1_n4579 = 1_n5832 & 1_n3303;
assign 1_n12436 = ~(1_n4508 ^ 1_n11432);
assign 1_n11947 = 1_n4715 | 1_n6561;
assign 1_n11926 = ~1_n9127;
assign 1_n7033 = ~1_n9093;
assign 1_n6985 = ~(1_n11393 ^ 1_n2997);
assign 1_n1551 = ~(1_n12247 | 1_n10754);
assign 1_n12571 = ~(1_n4525 ^ 1_n7684);
assign 1_n979 = 1_n4931 & 1_n11084;
assign 1_n7846 = ~1_n2590;
assign 1_n3190 = ~(1_n8747 ^ 1_n10737);
assign 1_n11807 = ~1_n8359;
assign 1_n328 = ~(1_n6525 ^ 1_n8232);
assign 1_n12401 = 1_n6995 & 1_n8690;
assign 1_n2306 = ~1_n2979;
assign 1_n6062 = 1_n11263 & 1_n13081;
assign 1_n13192 = 1_n6830 & 1_n3786;
assign 1_n1297 = 1_n8197 & 1_n10245;
assign 1_n10413 = 1_n13146 | 1_n8564;
assign 1_n1811 = ~(1_n6700 ^ 1_n5277);
assign 1_n7162 = ~(1_n9553 ^ 1_n6059);
assign 1_n5679 = ~1_n6655;
assign 1_n11205 = ~(1_n3699 ^ 1_n4976);
assign 1_n4831 = 1_n8111 & 1_n2967;
assign 1_n370 = ~(1_n12453 ^ 1_n7766);
assign 1_n5228 = 1_n1737 | 1_n9638;
assign 1_n3155 = 1_n925 & 1_n8199;
assign 1_n3103 = ~1_n11332;
assign 1_n10681 = ~1_n3130;
assign 1_n12438 = ~1_n6251;
assign 1_n1766 = 1_n12568 | 1_n8534;
assign 1_n7811 = 1_n829 | 1_n9075;
assign 1_n4988 = 1_n6986 | 1_n10430;
assign 1_n123 = 1_n991 | 1_n12501;
assign 1_n4350 = 1_n9662 & 1_n10386;
assign 1_n4359 = 1_n1536 | 1_n2675;
assign 1_n5205 = 1_n2044 & 1_n12293;
assign 1_n12639 = ~(1_n3542 ^ 1_n5418);
assign 1_n9292 = 1_n7434 & 1_n8185;
assign 1_n7040 = 1_n2163 & 1_n2618;
assign 1_n9775 = ~(1_n5689 ^ 1_n2467);
assign 1_n12655 = ~1_n10408;
assign 1_n13174 = 1_n2698 | 1_n9203;
assign 1_n1621 = ~1_n10162;
assign 1_n11087 = ~1_n5470;
assign 1_n9790 = ~1_n9965;
assign 1_n2436 = 1_n2407 & 1_n2578;
assign 1_n8277 = 1_n1571 | 1_n7935;
assign 1_n3396 = 1_n10884 & 1_n5926;
assign 1_n9841 = ~(1_n12074 ^ 1_n11767);
assign 1_n7409 = 1_n11490 & 1_n1206;
assign 1_n6259 = 1_n13182 | 1_n1985;
assign 1_n2327 = 1_n794 | 1_n2980;
assign 1_n7182 = 1_n3336 & 1_n5685;
assign 1_n11177 = ~(1_n752 ^ 1_n3982);
assign 1_n13097 = ~1_n9049;
assign 1_n3887 = ~(1_n3836 ^ 1_n11892);
assign 1_n2676 = 1_n7722 & 1_n11485;
assign 1_n5843 = 1_n1987 | 1_n285;
assign 1_n13092 = ~(1_n6712 ^ 1_n12186);
assign 1_n10958 = 1_n7010 & 1_n2752;
assign 1_n8758 = ~(1_n9609 ^ 1_n3134);
assign 1_n2626 = ~(1_n12942 ^ 1_n717);
assign 1_n12182 = ~(1_n10109 ^ 1_n3232);
assign 1_n7231 = 1_n560 | 1_n8490;
assign 1_n3927 = 1_n7231 | 1_n6583;
assign 1_n1352 = ~(1_n12816 | 1_n1510);
assign 1_n9684 = 1_n3102 & 1_n10385;
assign 1_n2083 = ~1_n791;
assign 1_n1342 = 1_n6137 & 1_n6379;
assign 1_n1944 = ~(1_n3357 ^ 1_n3012);
assign 1_n9281 = ~1_n11508;
assign 1_n886 = ~(1_n8122 ^ 1_n8995);
assign 1_n7303 = 1_n5076 | 1_n10106;
assign 1_n5532 = ~(1_n1391 ^ 1_n3737);
assign 1_n11958 = 1_n12493 | 1_n177;
assign 1_n6644 = 1_n10761 | 1_n206;
assign 1_n6298 = ~(1_n7161 | 1_n5076);
assign 1_n3392 = 1_n9353 & 1_n10063;
assign 1_n1700 = ~(1_n9074 ^ 1_n4799);
assign 1_n414 = ~(1_n9939 ^ 1_n2356);
assign 1_n3366 = 1_n8174 | 1_n2958;
assign 1_n12732 = ~1_n12965;
assign 1_n9870 = ~(1_n6053 | 1_n3080);
assign 1_n4765 = ~(1_n6661 ^ 1_n6675);
assign 1_n4581 = ~(1_n14 ^ 1_n3313);
assign 1_n7284 = 1_n3505 | 1_n6689;
assign 1_n6180 = ~1_n1283;
assign 1_n2453 = ~1_n11890;
assign 1_n380 = ~(1_n8240 ^ 1_n5373);
assign 1_n6433 = 1_n1912 & 1_n2498;
assign 1_n11060 = 1_n12660 | 1_n4881;
assign 1_n11873 = 1_n5768 & 1_n10563;
assign 1_n5682 = ~(1_n8823 ^ 1_n4434);
assign 1_n2782 = 1_n1250 | 1_n3113;
assign 1_n7011 = 1_n12395 | 1_n4960;
assign 1_n6701 = ~(1_n8207 ^ 1_n1106);
assign 1_n8963 = 1_n8847 & 1_n3007;
assign 1_n5979 = ~(1_n12279 ^ 1_n9210);
assign 1_n10140 = 1_n848 & 1_n10620;
assign 1_n7379 = 1_n10196 & 1_n10104;
assign 1_n8700 = ~1_n4813;
assign 1_n9764 = 1_n5770 | 1_n4312;
assign 1_n11541 = ~(1_n4639 ^ 1_n1457);
assign 1_n4919 = 1_n7468 & 1_n8442;
assign 1_n12347 = ~(1_n7910 ^ 1_n11358);
assign 1_n7115 = ~(1_n5126 ^ 1_n1363);
assign 1_n5870 = 1_n4964 & 1_n510;
assign 1_n13088 = ~1_n6537;
assign 1_n4413 = 1_n5661 & 1_n7174;
assign 1_n6786 = 1_n5092 & 1_n12462;
assign 1_n7738 = 1_n2829 | 1_n228;
assign 1_n10627 = ~(1_n4661 ^ 1_n8713);
assign 1_n4874 = 1_n11288 ^ 1_n8408;
assign 1_n5084 = 1_n2643 & 1_n4629;
assign 1_n7455 = 1_n4828 ^ 1_n8197;
assign 1_n11683 = ~1_n6937;
assign 1_n6070 = 1_n10792 | 1_n542;
assign 1_n8530 = 1_n4863 & 1_n243;
assign 1_n667 = 1_n11239 | 1_n8030;
assign 1_n7003 = 1_n8240 | 1_n9123;
assign 1_n141 = ~(1_n7289 ^ 1_n5463);
assign 1_n10484 = ~(1_n1756 ^ 1_n6380);
assign 1_n8456 = ~(1_n9871 ^ 1_n9350);
assign 1_n2036 = ~(1_n5810 ^ 1_n10720);
assign 1_n9407 = 1_n2582 | 1_n6635;
assign 1_n4053 = 1_n4201 | 1_n11144;
assign 1_n5433 = ~1_n9887;
assign 1_n8129 = ~1_n5962;
assign 1_n11238 = 1_n1053 | 1_n9491;
assign 1_n11004 = ~(1_n9433 ^ 1_n5628);
assign 1_n7222 = 1_n6651 | 1_n2658;
assign 1_n9659 = 1_n8585 | 1_n4640;
assign 1_n4116 = ~1_n3130;
assign 1_n13096 = 1_n3069 | 1_n8365;
assign 1_n7909 = ~(1_n9602 ^ 1_n2870);
assign 1_n3723 = 1_n8900 & 1_n5284;
assign 1_n85 = ~(1_n8256 ^ 1_n5582);
assign 1_n6405 = ~1_n124;
assign 1_n9245 = ~1_n9214;
assign 1_n2515 = ~1_n8924;
assign 1_n10725 = 1_n12007 & 1_n2066;
assign 1_n677 = 1_n1558 | 1_n1692;
assign 1_n13028 = ~1_n9732;
assign 1_n12687 = ~(1_n4458 | 1_n9091);
assign 1_n4701 = 1_n2214 | 1_n10589;
assign 1_n395 = 1_n11466 | 1_n479;
assign 1_n5258 = ~(1_n6009 | 1_n11089);
assign 1_n5372 = ~1_n6998;
assign 1_n10430 = ~1_n3130;
assign 1_n3970 = ~1_n11306;
assign 1_n2994 = ~(1_n13144 ^ 1_n4911);
assign 1_n12619 = ~(1_n2767 ^ 1_n6617);
assign 1_n8135 = ~(1_n10623 ^ 1_n1902);
assign 1_n1547 = ~(1_n986 ^ 1_n9471);
assign 1_n1882 = ~(1_n8064 ^ 1_n3843);
assign 1_n1573 = ~(1_n7476 ^ 1_n11948);
assign 1_n13241 = 1_n11915 | 1_n4133;
assign 1_n7586 = ~1_n8398;
assign 1_n6011 = 1_n590 & 1_n11168;
assign 1_n6539 = ~(1_n7100 | 1_n9045);
assign 1_n6145 = ~(1_n10785 | 1_n429);
assign 1_n12361 = ~(1_n9901 ^ 1_n1350);
assign 1_n6107 = ~(1_n9344 ^ 1_n5735);
assign 1_n11006 = ~1_n1065;
assign 1_n10809 = 1_n864 & 1_n8458;
assign 1_n1350 = ~(1_n11801 ^ 1_n6216);
assign 1_n11680 = ~1_n11891;
assign 1_n2763 = 1_n1280 | 1_n12907;
assign 1_n8718 = 1_n1346 & 1_n5839;
assign 1_n13015 = ~(1_n1537 ^ 1_n5464);
assign 1_n8623 = ~(1_n2323 | 1_n183);
assign 1_n8046 = 1_n937 & 1_n287;
assign 1_n212 = 1_n5257 & 1_n8425;
assign 1_n11158 = ~(1_n11108 ^ 1_n887);
assign 1_n153 = ~1_n1721;
assign 1_n8022 = 1_n5231 | 1_n7227;
assign 1_n1445 = 1_n3780 | 1_n8685;
assign 1_n2186 = 1_n3639 & 1_n503;
assign 1_n9213 = ~(1_n10540 ^ 1_n8343);
assign 1_n3459 = ~1_n3669;
assign 1_n3906 = ~1_n11881;
assign 1_n6466 = 1_n7604 | 1_n4585;
assign 1_n6927 = ~(1_n659 ^ 1_n1591);
assign 1_n1802 = ~(1_n5465 ^ 1_n7760);
assign 1_n2755 = 1_n7986 | 1_n8540;
assign 1_n6859 = 1_n8776 | 1_n10761;
assign 1_n1979 = 1_n10221 | 1_n2977;
assign 1_n8158 = 1_n12953 ^ 1_n6140;
assign 1_n2462 = ~1_n13058;
assign 1_n7194 = 1_n6971 | 1_n3798;
assign 1_n11274 = ~(1_n3224 ^ 1_n340);
assign 1_n8606 = 1_n9353 & 1_n9915;
assign 1_n13146 = ~1_n3868;
assign 1_n5014 = ~(1_n9858 ^ 1_n618);
assign 1_n6295 = ~1_n2758;
assign 1_n5124 = ~(1_n10167 ^ 1_n4643);
assign 1_n5213 = ~(1_n11572 | 1_n1584);
assign 1_n10970 = ~(1_n7887 ^ 1_n626);
assign 1_n3964 = ~(1_n9938 ^ 1_n8184);
assign 1_n8577 = 1_n9797 & 1_n12584;
assign 1_n9527 = ~(1_n2541 | 1_n11280);
assign 1_n12417 = 1_n48 | 1_n11144;
assign 1_n4206 = 1_n3755 | 1_n2845;
assign 1_n7933 = 1_n13168 | 1_n1985;
assign 1_n2466 = 1_n2861 | 1_n12388;
assign 1_n4414 = 1_n12734 & 1_n2441;
assign 1_n10761 = 1_n6405;
assign 1_n6379 = 1_n5700 | 1_n9975;
assign 1_n3527 = 1_n12596 | 1_n5242;
assign 1_n7900 = ~1_n9747;
assign 1_n1778 = 1_n12745 & 1_n1968;
assign 1_n11511 = 1_n10343 | 1_n6983;
assign 1_n11676 = ~(1_n6296 ^ 1_n11073);
assign 1_n7089 = ~1_n6286;
assign 1_n8621 = ~1_n9415;
assign 1_n7123 = ~(1_n11004 ^ 1_n5994);
assign 1_n12423 = ~(1_n90 ^ 1_n6262);
assign 1_n8377 = ~(1_n5447 ^ 1_n2367);
assign 1_n7226 = 1_n6011 | 1_n13105;
assign 1_n5035 = ~1_n13040;
assign 1_n474 = ~(1_n11930 ^ 1_n9316);
assign 1_n12766 = 1_n595 | 1_n3221;
assign 1_n7660 = ~(1_n1490 ^ 1_n54);
assign 1_n1854 = 1_n3017 & 1_n6921;
assign 1_n12969 = ~1_n7229;
assign 1_n7731 = 1_n6638 | 1_n1043;
assign 1_n2156 = 1_n10000 | 1_n10534;
assign 1_n1505 = ~1_n7779;
assign 1_n7238 = 1_n4957 ^ 1_n8452;
assign 1_n10441 = ~(1_n17 | 1_n11460);
assign 1_n12486 = ~(1_n10502 ^ 1_n7617);
assign 1_n8140 = ~(1_n11765 ^ 1_n8851);
assign 1_n12959 = ~1_n10770;
assign 1_n249 = 1_n1680 | 1_n451;
assign 1_n1415 = ~(1_n3434 ^ 1_n5211);
assign 1_n4936 = 1_n2623;
assign 1_n10923 = 1_n1378 & 1_n9835;
assign 1_n7689 = 1_n12757 | 1_n225;
assign 1_n6557 = ~1_n8332;
assign 1_n4908 = 1_n6668 & 1_n10451;
assign 1_n12433 = 1_n7575 | 1_n6624;
assign 1_n796 = ~(1_n12506 ^ 1_n4631);
assign 1_n10821 = 1_n7857 & 1_n1396;
assign 1_n4763 = ~(1_n9555 | 1_n1830);
assign 1_n1224 = ~(1_n2166 | 1_n3862);
assign 1_n899 = ~1_n9187;
assign 1_n467 = ~1_n10572;
assign 1_n7269 = 1_n822 | 1_n11176;
assign 1_n1278 = 1_n5334 ^ 1_n9215;
assign 1_n4980 = ~1_n11634;
assign 1_n2615 = 1_n11051 & 1_n7953;
assign 1_n13132 = 1_n1682 & 1_n1306;
assign 1_n10360 = 1_n3302 & 1_n8133;
assign 1_n2920 = 1_n12814 | 1_n5740;
assign 1_n8930 = ~(1_n484 | 1_n7618);
assign 1_n9599 = ~(1_n9853 ^ 1_n12044);
assign 1_n2933 = ~(1_n3589 | 1_n7217);
assign 1_n4253 = ~1_n10770;
assign 1_n335 = ~(1_n688 | 1_n9816);
assign 1_n769 = ~(1_n10919 ^ 1_n4765);
assign 1_n9409 = 1_n5441 | 1_n4164;
assign 1_n11041 = 1_n7769 | 1_n7162;
assign 1_n4032 = ~(1_n6530 | 1_n4950);
assign 1_n12476 = ~(1_n10499 | 1_n12269);
assign 1_n1963 = ~1_n9204;
assign 1_n9334 = 1_n11381 | 1_n1848;
assign 1_n11081 = ~(1_n4800 | 1_n2089);
assign 1_n578 = ~1_n7959;
assign 1_n4111 = 1_n7772 & 1_n12853;
assign 1_n10249 = 1_n944 & 1_n1673;
assign 1_n3588 = ~1_n6831;
assign 1_n1272 = ~(1_n4325 ^ 1_n1743);
assign 1_n2754 = 1_n2411 & 1_n757;
assign 1_n10112 = ~1_n10594;
assign 1_n3104 = 1_n11108 & 1_n5731;
assign 1_n9227 = ~(1_n9166 | 1_n4284);
assign 1_n6143 = 1_n1609 ^ 1_n8544;
assign 1_n9009 = ~(1_n8215 | 1_n270);
assign 1_n9665 = ~(1_n7843 ^ 1_n5151);
assign 1_n12647 = 1_n12316 | 1_n11960;
assign 1_n7342 = ~1_n9249;
assign 1_n2104 = ~1_n1202;
assign 1_n10901 = ~(1_n6559 | 1_n8071);
assign 1_n8142 = ~1_n1731;
assign 1_n12564 = ~(1_n6338 ^ 1_n9644);
assign 1_n11141 = 1_n759 & 1_n12035;
assign 1_n1367 = ~1_n3558;
assign 1_n2100 = 1_n9931 | 1_n8348;
assign 1_n3672 = ~(1_n7769 ^ 1_n2959);
assign 1_n8938 = 1_n7201 | 1_n10725;
assign 1_n6323 = 1_n9378 | 1_n2632;
assign 1_n8427 = ~(1_n7514 ^ 1_n10305);
assign 1_n10317 = ~(1_n1148 ^ 1_n13003);
assign 1_n8227 = ~(1_n7973 ^ 1_n5014);
assign 1_n7862 = 1_n10256 | 1_n9159;
assign 1_n11123 = 1_n1869 | 1_n3981;
assign 1_n11950 = ~1_n13058;
assign 1_n12690 = ~(1_n12449 ^ 1_n7104);
assign 1_n11631 = ~(1_n3109 ^ 1_n5275);
assign 1_n6300 = 1_n2767 | 1_n10584;
assign 1_n2171 = ~(1_n8847 | 1_n3007);
assign 1_n6404 = 1_n5041;
assign 1_n9616 = ~(1_n1669 ^ 1_n4820);
assign 1_n8369 = ~(1_n12771 ^ 1_n5813);
assign 1_n4916 = 1_n12411 | 1_n4745;
assign 1_n8937 = ~(1_n4690 ^ 1_n11435);
assign 1_n13117 = ~1_n9531;
assign 1_n3994 = ~(1_n12285 ^ 1_n82);
assign 1_n8486 = ~1_n12987;
assign 1_n7340 = 1_n10929 | 1_n12273;
assign 1_n5453 = ~(1_n1245 ^ 1_n6386);
assign 1_n8485 = ~1_n4798;
assign 1_n91 = 1_n6796 & 1_n8984;
assign 1_n6210 = ~1_n13201;
assign 1_n12267 = 1_n5554 & 1_n11321;
assign 1_n10105 = ~1_n9125;
assign 1_n9062 = 1_n12626 & 1_n1562;
assign 1_n12212 = ~1_n3448;
assign 1_n6 = ~(1_n5791 | 1_n2517);
assign 1_n1341 = ~(1_n8654 ^ 1_n2457);
assign 1_n13072 = 1_n10977 | 1_n4230;
assign 1_n12608 = ~(1_n4649 | 1_n10866);
assign 1_n5345 = ~(1_n5206 | 1_n9789);
assign 1_n6872 = ~(1_n3828 ^ 1_n4566);
assign 1_n358 = ~(1_n530 ^ 1_n1022);
assign 1_n3279 = 1_n2474 | 1_n12017;
assign 1_n12762 = 1_n785 | 1_n8534;
assign 1_n8359 = 1_n6341 & 1_n9244;
assign 1_n4477 = ~(1_n9824 ^ 1_n13078);
assign 1_n11343 = 1_n11929 | 1_n2958;
assign 1_n1830 = 1_n6873 & 1_n7555;
assign 1_n6682 = ~(1_n3599 ^ 1_n773);
assign 1_n3508 = ~1_n7702;
assign 1_n5594 = ~(1_n7296 ^ 1_n12546);
assign 1_n958 = ~1_n13065;
assign 1_n698 = 1_n4114 & 1_n510;
assign 1_n7383 = 1_n1672 & 1_n6321;
assign 1_n6611 = 1_n12324 | 1_n4724;
assign 1_n2841 = 1_n11771 & 1_n128;
assign 1_n7246 = ~(1_n8055 ^ 1_n712);
assign 1_n5667 = ~1_n9906;
assign 1_n1623 = 1_n6228 & 1_n12774;
assign 1_n8170 = 1_n6630 | 1_n8005;
assign 1_n5612 = ~(1_n5140 | 1_n6791);
assign 1_n10447 = ~1_n4006;
assign 1_n5276 = ~(1_n11301 ^ 1_n5444);
assign 1_n4898 = 1_n12465 | 1_n644;
assign 1_n12562 = ~(1_n5052 ^ 1_n11325);
assign 1_n4156 = 1_n5044 ^ 1_n1444;
assign 1_n12409 = ~(1_n3905 ^ 1_n9111);
assign 1_n6274 = ~1_n10560;
assign 1_n11684 = 1_n9148 & 1_n282;
assign 1_n464 = ~1_n11448;
assign 1_n9645 = 1_n18 | 1_n6732;
assign 1_n12898 = ~(1_n5558 ^ 1_n9941);
assign 1_n3133 = 1_n6541 & 1_n9519;
assign 1_n6643 = 1_n153 & 1_n9996;
assign 1_n8590 = 1_n2057 & 1_n1198;
assign 1_n4259 = 1_n5559 & 1_n1526;
assign 1_n1305 = 1_n9318 | 1_n10532;
assign 1_n10671 = 1_n8925 & 1_n2930;
assign 1_n9104 = 1_n11170 | 1_n5575;
assign 1_n2080 = ~1_n7812;
assign 1_n3208 = ~1_n9846;
assign 1_n2780 = ~(1_n8338 | 1_n4200);
assign 1_n2441 = ~1_n3097;
assign 1_n9812 = 1_n13009 & 1_n7105;
assign 1_n6002 = ~(1_n10133 | 1_n8052);
assign 1_n639 = 1_n1050 & 1_n11728;
assign 1_n3560 = 1_n9868 | 1_n7846;
assign 1_n5647 = 1_n11807 & 1_n1366;
assign 1_n3938 = 1_n8720 | 1_n1554;
assign 1_n947 = ~1_n11324;
assign 1_n10563 = 1_n10770 & 1_n3769;
assign 1_n5639 = 1_n495 | 1_n6853;
assign 1_n2090 = 1_n947 | 1_n11950;
assign 1_n11622 = ~(1_n8994 ^ 1_n6847);
assign 1_n1694 = ~(1_n10167 | 1_n11158);
assign 1_n5855 = 1_n7852 | 1_n1449;
assign 1_n5238 = 1_n3032 | 1_n12244;
assign 1_n1550 = 1_n9867 | 1_n5076;
assign 1_n4476 = ~(1_n3358 ^ 1_n5927);
assign 1_n1429 = ~(1_n8180 | 1_n2667);
assign 1_n11658 = ~(1_n2248 ^ 1_n462);
assign 1_n619 = 1_n8919 | 1_n8549;
assign 1_n10258 = ~1_n9875;
assign 1_n9189 = ~(1_n10945 ^ 1_n3969);
assign 1_n3245 = 1_n4491 | 1_n11592;
assign 1_n8965 = 1_n2773 & 1_n6380;
assign 1_n9529 = 1_n11864 | 1_n8079;
assign 1_n12130 = 1_n6968 | 1_n10761;
assign 1_n12836 = ~(1_n13037 ^ 1_n12865);
assign 1_n6779 = ~(1_n1839 | 1_n7182);
assign 1_n8755 = ~1_n2393;
assign 1_n5956 = 1_n8249 | 1_n7723;
assign 1_n8430 = 1_n1082 | 1_n12258;
assign 1_n12580 = 1_n12837 | 1_n4230;
assign 1_n6731 = ~1_n10809;
assign 1_n457 = 1_n2941 | 1_n9822;
assign 1_n2138 = ~(1_n1068 ^ 1_n11538);
assign 1_n3548 = ~(1_n9775 ^ 1_n4282);
assign 1_n4250 = 1_n2284 & 1_n8770;
assign 1_n848 = ~1_n1569;
assign 1_n9726 = ~(1_n2359 ^ 1_n4871);
assign 1_n7319 = 1_n3805 | 1_n2675;
assign 1_n4109 = ~(1_n9838 | 1_n12943);
assign 1_n12591 = ~(1_n10310 ^ 1_n12414);
assign 1_n2733 = ~(1_n12272 | 1_n10455);
assign 1_n11280 = ~(1_n8285 ^ 1_n5481);
assign 1_n7096 = 1_n3572 | 1_n9080;
assign 1_n9955 = 1_n5306 | 1_n12544;
assign 1_n7631 = ~(1_n7648 | 1_n11208);
assign 1_n8941 = ~1_n4335;
assign 1_n11240 = 1_n9035 | 1_n3794;
assign 1_n1745 = 1_n3104 | 1_n11093;
assign 1_n8956 = 1_n8277 | 1_n2337;
assign 1_n9232 = 1_n2136 & 1_n13069;
assign 1_n1201 = ~(1_n2925 ^ 1_n4583);
assign 1_n2016 = ~(1_n10152 ^ 1_n8810);
assign 1_n7834 = 1_n4530 & 1_n7256;
assign 1_n957 = ~(1_n3984 ^ 1_n12964);
assign 1_n9367 = 1_n1064 & 1_n12952;
assign 1_n7897 = 1_n6271 | 1_n8754;
assign 1_n12488 = ~(1_n1535 ^ 1_n5775);
assign 1_n1747 = 1_n542 | 1_n1570;
assign 1_n8406 = 1_n2705 | 1_n5387;
assign 1_n13212 = 1_n7396 | 1_n7723;
assign 1_n1659 = ~1_n11327;
assign 1_n5747 = ~(1_n6537 ^ 1_n7670);
assign 1_n2536 = ~1_n6917;
assign 1_n10611 = 1_n10795 | 1_n5992;
assign 1_n2707 = 1_n3684 & 1_n11672;
assign 1_n7562 = 1_n5696 & 1_n538;
assign 1_n11425 = 1_n6512 & 1_n11189;
assign 1_n919 = 1_n11240 & 1_n2322;
assign 1_n6547 = 1_n7098 & 1_n9349;
assign 1_n9538 = ~1_n5995;
assign 1_n6439 = ~1_n8233;
assign 1_n10030 = 1_n12455 & 1_n12161;
assign 1_n10582 = 1_n5343 & 1_n2821;
assign 1_n1960 = ~(1_n7340 ^ 1_n9287);
assign 1_n3617 = 1_n3255 | 1_n6823;
assign 1_n9011 = 1_n368 & 1_n10839;
assign 1_n5504 = 1_n7772 & 1_n9093;
assign 1_n5231 = 1_n3225 | 1_n1570;
assign 1_n7152 = ~1_n3815;
assign 1_n2669 = ~1_n2174;
assign 1_n10688 = ~(1_n3191 ^ 1_n8588);
assign 1_n3343 = 1_n4961 | 1_n7292;
assign 1_n10253 = 1_n126 & 1_n5783;
assign 1_n6606 = ~1_n10785;
assign 1_n8457 = 1_n6846 | 1_n8534;
assign 1_n7108 = 1_n12711 | 1_n11259;
assign 1_n8452 = 1_n8228 & 1_n5962;
assign 1_n3647 = 1_n10761 | 1_n7935;
assign 1_n8754 = ~1_n2590;
assign 1_n606 = ~(1_n5441 ^ 1_n4164);
assign 1_n915 = ~(1_n1028 ^ 1_n3425);
assign 1_n12326 = 1_n12558 | 1_n11397;
assign 1_n2513 = 1_n12304 & 1_n12574;
assign 1_n4526 = ~(1_n10317 ^ 1_n3023);
assign 1_n3176 = 1_n2402 & 1_n12451;
assign 1_n11597 = 1_n1634 | 1_n12997;
assign 1_n1458 = 1_n5452 & 1_n12681;
assign 1_n2906 = ~(1_n13110 ^ 1_n5005);
assign 1_n6075 = ~(1_n11500 ^ 1_n4769);
assign 1_n7237 = ~(1_n3776 ^ 1_n1551);
assign 1_n146 = ~1_n4579;
assign 1_n8631 = ~1_n12091;
assign 1_n10491 = 1_n5839 | 1_n1346;
assign 1_n352 = 1_n7621 | 1_n2077;
assign 1_n11400 = ~1_n12260;
assign 1_n8774 = ~(1_n6436 ^ 1_n6735);
assign 1_n4947 = 1_n9709;
assign 1_n11770 = ~(1_n9621 | 1_n7888);
assign 1_n7300 = 1_n11210 | 1_n2116;
assign 1_n1426 = 1_n12371 & 1_n12297;
assign 1_n10084 = ~(1_n10358 ^ 1_n3574);
assign 1_n4481 = ~1_n3579;
assign 1_n3252 = ~(1_n8369 ^ 1_n3286);
assign 1_n9979 = ~(1_n6233 ^ 1_n5598);
assign 1_n1266 = ~(1_n1797 ^ 1_n4676);
assign 1_n627 = 1_n5134 & 1_n6311;
assign 1_n2245 = ~(1_n9763 | 1_n11812);
assign 1_n5615 = 1_n6639 & 1_n12031;
assign 1_n10601 = 1_n9484 & 1_n2842;
assign 1_n8241 = ~(1_n9597 ^ 1_n7531);
assign 1_n8881 = 1_n2095 | 1_n2599;
assign 1_n10368 = 1_n5395 | 1_n7915;
assign 1_n10779 = ~(1_n7378 ^ 1_n3202);
assign 1_n863 = 1_n7263 & 1_n12492;
assign 1_n10802 = ~(1_n13231 ^ 1_n7644);
assign 1_n6326 = 1_n1456 & 1_n11610;
assign 1_n11827 = 1_n12090 | 1_n2611;
assign 1_n10857 = 1_n6590 | 1_n10029;
assign 1_n768 = 1_n633 | 1_n1600;
assign 1_n8320 = ~(1_n7355 ^ 1_n9259);
assign 1_n1892 = 1_n8129 | 1_n10319;
assign 1_n4228 = ~(1_n4015 | 1_n7465);
assign 1_n12268 = ~(1_n2403 | 1_n11348);
assign 1_n1645 = 1_n6110 | 1_n5691;
assign 1_n7173 = ~(1_n6165 ^ 1_n2448);
assign 1_n5305 = 1_n863 | 1_n7559;
assign 1_n4815 = ~1_n6017;
assign 1_n2778 = 1_n2955 | 1_n8145;
assign 1_n674 = 1_n8325 | 1_n7221;
assign 1_n6063 = ~1_n6655;
assign 1_n1969 = ~(1_n10406 ^ 1_n11126);
assign 1_n13236 = ~(1_n88 ^ 1_n11411);
assign 1_n8602 = 1_n7917 & 1_n2049;
assign 1_n5302 = ~(1_n661 ^ 1_n1036);
assign 1_n13235 = ~1_n2948;
assign 1_n2775 = ~(1_n3977 ^ 1_n7175);
assign 1_n10974 = ~1_n1916;
assign 1_n7819 = ~1_n12352;
assign 1_n12508 = ~1_n9151;
assign 1_n7477 = ~(1_n7091 ^ 1_n10440);
assign 1_n9368 = ~(1_n10876 ^ 1_n6645);
assign 1_n7384 = ~(1_n4586 ^ 1_n1431);
assign 1_n4647 = ~(1_n9997 ^ 1_n9387);
assign 1_n8367 = ~(1_n3511 | 1_n11738);
assign 1_n10034 = 1_n10230 & 1_n8525;
assign 1_n5064 = ~(1_n930 ^ 1_n2055);
assign 1_n321 = ~1_n6826;
assign 1_n568 = 1_n6190 | 1_n1861;
assign 1_n7646 = ~(1_n7399 ^ 1_n11984);
assign 1_n6614 = 1_n4980 | 1_n10179;
assign 1_n11890 = 1_n7772 & 1_n4470;
assign 1_n13063 = ~1_n3499;
assign 1_n9749 = 1_n5752 & 1_n2177;
assign 1_n6170 = 1_n5697 & 1_n10636;
assign 1_n9129 = ~1_n817;
assign 1_n4037 = ~(1_n12889 ^ 1_n171);
assign 1_n9713 = ~(1_n5112 | 1_n1180);
assign 1_n3542 = ~(1_n8901 ^ 1_n11552);
assign 1_n4830 = ~1_n6920;
assign 1_n3259 = ~1_n5969;
assign 1_n7801 = 1_n10571 | 1_n1107;
assign 1_n12781 = 1_n511 & 1_n12162;
assign 1_n248 = 1_n8349 | 1_n12823;
assign 1_n11178 = 1_n2590 & 1_n6392;
assign 1_n8362 = ~(1_n495 ^ 1_n461);
assign 1_n8600 = 1_n8263 & 1_n2988;
assign 1_n9621 = 1_n12348 & 1_n854;
assign 1_n9882 = ~1_n5536;
assign 1_n12213 = 1_n766 | 1_n129;
assign 1_n4600 = 1_n787 | 1_n9223;
assign 1_n12802 = 1_n4832 & 1_n820;
assign 1_n11920 = ~1_n8506;
assign 1_n12698 = ~1_n2389;
assign 1_n3505 = ~1_n12965;
assign 1_n9016 = ~1_n8332;
assign 1_n8182 = 1_n2449 | 1_n6265;
assign 1_n4509 = 1_n5671 & 1_n510;
assign 1_n8223 = 1_n6245 | 1_n2449;
assign 1_n7236 = ~(1_n8418 ^ 1_n1260);
assign 1_n6620 = ~(1_n1752 ^ 1_n12367);
assign 1_n5778 = ~(1_n7725 ^ 1_n13023);
assign 1_n9876 = ~(1_n216 ^ 1_n3772);
assign 1_n2286 = ~(1_n1409 ^ 1_n5657);
assign 1_n338 = ~1_n12853;
assign 1_n4041 = 1_n8079 | 1_n542;
assign 1_n11828 = 1_n2478 & 1_n10715;
assign 1_n4306 = 1_n8254 | 1_n12789;
assign 1_n6499 = ~1_n7270;
assign 1_n5798 = ~(1_n3183 ^ 1_n11445);
assign 1_n12519 = 1_n12689 & 1_n4103;
assign 1_n12299 = ~(1_n11189 | 1_n6512);
assign 1_n2845 = ~(1_n1365 ^ 1_n11162);
assign 1_n4126 = ~(1_n10366 ^ 1_n12474);
assign 1_n3918 = 1_n8168 & 1_n12944;
assign 1_n3877 = ~(1_n8689 | 1_n8630);
assign 1_n8680 = 1_n6957 | 1_n9370;
assign 1_n1354 = ~1_n6023;
assign 1_n4939 = 1_n8796 | 1_n10214;
assign 1_n7335 = 1_n4108 & 1_n3554;
assign 1_n2506 = 1_n10908 & 1_n411;
assign 1_n9913 = ~1_n7812;
assign 1_n4035 = ~(1_n11812 ^ 1_n1066);
assign 1_n10599 = 1_n8463 | 1_n12655;
assign 1_n7995 = ~(1_n5622 | 1_n10531);
assign 1_n2347 = ~(1_n2653 | 1_n13111);
assign 1_n10559 = ~(1_n12993 ^ 1_n6589);
assign 1_n1909 = ~(1_n4245 ^ 1_n5866);
assign 1_n2258 = ~(1_n8953 ^ 1_n10930);
assign 1_n8598 = ~1_n499;
assign 1_n7367 = ~(1_n3612 ^ 1_n9312);
assign 1_n1397 = ~(1_n8349 ^ 1_n10121);
assign 1_n678 = ~(1_n5056 ^ 1_n2819);
assign 1_n8720 = ~1_n10162;
assign 1_n11667 = ~(1_n11826 ^ 1_n8353);
assign 1_n5410 = ~(1_n6108 | 1_n4091);
assign 1_n11486 = ~(1_n4049 | 1_n11161);
assign 1_n2836 = ~(1_n3660 ^ 1_n8958);
assign 1_n6130 = 1_n10143 | 1_n13238;
assign 1_n10730 = ~1_n9528;
assign 1_n7147 = 1_n6825 & 1_n6467;
assign 1_n9139 = ~(1_n5774 ^ 1_n2236);
assign 1_n11335 = ~(1_n11652 ^ 1_n1446);
assign 1_n2646 = ~(1_n3310 ^ 1_n4909);
assign 1_n6738 = 1_n202 | 1_n10106;
assign 1_n307 = 1_n5520 | 1_n542;
assign 1_n2328 = ~(1_n4679 ^ 1_n8085);
assign 1_n3788 = ~(1_n1475 ^ 1_n12489);
assign 1_n9322 = ~(1_n4810 ^ 1_n3936);
assign 1_n1687 = 1_n2057 & 1_n2295;
assign 1_n7151 = 1_n1136 | 1_n716;
assign 1_n10553 = ~(1_n12936 ^ 1_n7312);
assign 1_n3423 = 1_n119 | 1_n6404;
assign 1_n7866 = 1_n6764 & 1_n13138;
assign 1_n4420 = ~1_n10642;
assign 1_n10061 = ~(1_n11820 ^ 1_n9979);
assign 1_n751 = ~(1_n5868 ^ 1_n5805);
assign 1_n10909 = 1_n12775 & 1_n4359;
assign 1_n10580 = ~(1_n9856 | 1_n6101);
assign 1_n5181 = 1_n8858 & 1_n8194;
assign 1_n12250 = 1_n8557 & 1_n12756;
assign 1_n6458 = ~(1_n1087 ^ 1_n9546);
assign 1_n4263 = ~(1_n10853 ^ 1_n1311);
assign 1_n4791 = 1_n5028 | 1_n2735;
assign 1_n8153 = ~1_n8459;
assign 1_n12366 = ~(1_n9833 | 1_n5746);
assign 1_n9805 = 1_n10034 ^ 1_n2951;
assign 1_n11191 = 1_n11677 | 1_n2572;
assign 1_n4031 = ~(1_n12984 ^ 1_n9646);
assign 1_n10470 = ~1_n11885;
assign 1_n7277 = 1_n1331 | 1_n11107;
assign 1_n2464 = 1_n3854 | 1_n11668;
assign 1_n4511 = ~(1_n4552 ^ 1_n3324);
assign 1_n3968 = 1_n9940 & 1_n8397;
assign 1_n4028 = ~1_n7792;
assign 1_n9365 = 1_n13084 | 1_n479;
assign 1_n10700 = 1_n5794 | 1_n3512;
assign 1_n4161 = ~1_n287;
assign 1_n5669 = 1_n5168 | 1_n11107;
assign 1_n73 = 1_n3129 | 1_n3143;
assign 1_n5954 = ~1_n1978;
assign 1_n6221 = ~(1_n1745 ^ 1_n3349);
assign 1_n10709 = ~(1_n368 ^ 1_n5891);
assign 1_n506 = ~(1_n3314 ^ 1_n9583);
assign 1_n2142 = ~(1_n5621 ^ 1_n3043);
assign 1_n1907 = 1_n10835 | 1_n10843;
assign 1_n9359 = ~(1_n8627 ^ 1_n12694);
assign 1_n6597 = ~(1_n8573 ^ 1_n12096);
assign 1_n9076 = 1_n7506 & 1_n10543;
assign 1_n9049 = 1_n10626 & 1_n8271;
assign 1_n5688 = ~1_n4748;
assign 1_n12360 = 1_n11115 & 1_n2509;
assign 1_n11331 = ~1_n2751;
assign 1_n789 = ~1_n9216;
assign 1_n11277 = ~(1_n12577 | 1_n2055);
assign 1_n7805 = ~1_n13058;
assign 1_n12214 = ~(1_n12260 ^ 1_n3142);
assign 1_n1096 = 1_n9668 | 1_n10886;
assign 1_n1256 = 1_n1058 | 1_n3817;
assign 1_n13080 = ~1_n5556;
assign 1_n8151 = ~(1_n6964 ^ 1_n4539);
assign 1_n6685 = 1_n10263 | 1_n7221;
assign 1_n4347 = ~(1_n1306 ^ 1_n7753);
assign 1_n4376 = 1_n6040 | 1_n10179;
assign 1_n8805 = 1_n8410 ^ 1_n10800;
assign 1_n6758 = 1_n8308 & 1_n4330;
assign 1_n2670 = ~1_n10103;
assign 1_n6759 = ~(1_n2638 ^ 1_n415);
assign 1_n4096 = 1_n2527 | 1_n2030;
assign 1_n12473 = ~(1_n7299 ^ 1_n4082);
assign 1_n12682 = 1_n3225 | 1_n6041;
assign 1_n626 = 1_n2889 | 1_n121;
assign 1_n8240 = 1_n6419 | 1_n11107;
assign 1_n1639 = 1_n3982 | 1_n752;
assign 1_n7310 = 1_n9383 | 1_n2958;
assign 1_n7271 = 1_n10400 | 1_n8348;
assign 1_n13068 = 1_n1235 | 1_n8673;
assign 1_n11552 = 1_n12416 | 1_n10029;
assign 1_n9087 = ~(1_n2948 ^ 1_n8155);
assign 1_n12150 = 1_n3866 | 1_n2675;
assign 1_n10160 = 1_n6438 | 1_n7530;
assign 1_n7431 = ~(1_n4304 ^ 1_n11885);
assign 1_n11842 = ~1_n10615;
assign 1_n6027 = ~(1_n11896 ^ 1_n7120);
assign 1_n8216 = 1_n3302 | 1_n8133;
assign 1_n13181 = ~1_n937;
assign 1_n244 = ~(1_n13093 | 1_n4338);
assign 1_n349 = 1_n9919 | 1_n6635;
assign 1_n4523 = 1_n2520 & 1_n255;
assign 1_n934 = 1_n5914 | 1_n3356;
assign 1_n10208 = 1_n11628 | 1_n8563;
assign 1_n5316 = ~(1_n5943 ^ 1_n12929);
assign 1_n5019 = ~(1_n12422 | 1_n10198);
assign 1_n7390 = 1_n1214 | 1_n9418;
assign 1_n6968 = ~1_n3669;
assign 1_n5971 = ~1_n11766;
assign 1_n3282 = 1_n11319 | 1_n4067;
assign 1_n9195 = 1_n11418;
assign 1_n8131 = ~1_n2252;
assign 1_n84 = 1_n6503 & 1_n310;
assign 1_n136 = 1_n9339 | 1_n10029;
assign 1_n7261 = 1_n10136 | 1_n3174;
assign 1_n2267 = 1_n5835 | 1_n3488;
assign 1_n3903 = 1_n5586 & 1_n3832;
assign 1_n8371 = ~(1_n229 | 1_n651);
assign 1_n11975 = ~1_n11288;
assign 1_n5735 = ~(1_n6566 ^ 1_n6969);
assign 1_n6451 = 1_n13106 ^ 1_n7447;
assign 1_n9219 = ~(1_n3711 ^ 1_n8294);
assign 1_n11268 = ~(1_n10254 | 1_n4730);
assign 1_n1034 = ~(1_n1835 ^ 1_n11349);
assign 1_n10953 = ~(1_n12259 | 1_n3048);
assign 1_n10228 = 1_n122 | 1_n6062;
assign 1_n11893 = 1_n12614 ^ 1_n864;
assign 1_n3991 = ~(1_n404 ^ 1_n6759);
assign 1_n8418 = 1_n8790 & 1_n10312;
assign 1_n8235 = 1_n5954 & 1_n3168;
assign 1_n11375 = 1_n2677 & 1_n10912;
assign 1_n2878 = ~(1_n9387 | 1_n9997);
assign 1_n6721 = ~1_n11891;
assign 1_n6853 = 1_n1779 & 1_n10132;
assign 1_n1087 = 1_n7234 | 1_n8702;
assign 1_n530 = ~1_n4987;
assign 1_n12793 = 1_n6191 | 1_n1894;
assign 1_n8339 = ~1_n11559;
assign 1_n2864 = ~(1_n2100 ^ 1_n12220);
assign 1_n670 = 1_n1220 & 1_n3878;
assign 1_n12038 = ~(1_n664 ^ 1_n3968);
assign 1_n6955 = ~(1_n3265 ^ 1_n1433);
assign 1_n7818 = ~(1_n9065 ^ 1_n3332);
assign 1_n1239 = 1_n12281 & 1_n1698;
assign 1_n5959 = ~1_n7806;
assign 1_n10002 = 1_n9732 & 1_n854;
assign 1_n3732 = 1_n6414 & 1_n12770;
assign 1_n7946 = 1_n8327 | 1_n3374;
assign 1_n13023 = 1_n7022 & 1_n3656;
assign 1_n9746 = ~(1_n10395 ^ 1_n102);
assign 1_n8357 = ~(1_n10294 ^ 1_n8283);
assign 1_n10613 = ~(1_n10549 ^ 1_n3693);
assign 1_n10949 = 1_n406 | 1_n7998;
assign 1_n7281 = 1_n11218 | 1_n2059;
assign 1_n2697 = ~(1_n10475 ^ 1_n7021);
assign 1_n6340 = ~(1_n10718 ^ 1_n10124);
assign 1_n9223 = 1_n12954;
assign 1_n10723 = ~(1_n12152 | 1_n7735);
assign 1_n2224 = 1_n12754 | 1_n11714;
assign 1_n10849 = ~1_n12822;
assign 1_n10767 = ~(1_n9101 ^ 1_n2214);
assign 1_n125 = 1_n9039 | 1_n10466;
assign 1_n2465 = 1_n3361 ^ 1_n4908;
assign 1_n1146 = ~(1_n5727 ^ 1_n13175);
assign 1_n3983 = 1_n11352 | 1_n10029;
assign 1_n1466 = 1_n12613 & 1_n375;
assign 1_n13158 = ~(1_n12296 ^ 1_n10096);
assign 1_n4438 = 1_n12493 | 1_n11668;
assign 1_n10027 = ~(1_n6992 ^ 1_n10297);
assign 1_n7308 = ~(1_n9240 ^ 1_n10659);
assign 1_n3911 = ~1_n11180;
assign 1_n12913 = 1_n121 | 1_n4960;
assign 1_n8498 = ~1_n10162;
assign 1_n3244 = ~(1_n1524 ^ 1_n6873);
assign 1_n6509 = 1_n13168 | 1_n2544;
assign 1_n12981 = ~(1_n8085 | 1_n4679);
assign 1_n3028 = 1_n75 | 1_n8024;
assign 1_n11249 = 1_n7970 | 1_n3075;
assign 1_n4329 = ~(1_n8273 ^ 1_n4156);
assign 1_n11606 = 1_n9199 & 1_n11192;
assign 1_n12938 = 1_n3489 | 1_n3715;
assign 1_n10364 = 1_n9987 & 1_n7901;
assign 1_n10917 = ~(1_n6240 ^ 1_n7211);
assign 1_n11024 = 1_n11514 | 1_n8777;
assign 1_n984 = ~(1_n3123 ^ 1_n9212);
assign 1_n2182 = 1_n1515 | 1_n7004;
assign 1_n4233 = ~(1_n11133 ^ 1_n1291);
assign 1_n707 = ~(1_n2811 ^ 1_n11250);
assign 1_n13210 = 1_n11704 & 1_n2348;
assign 1_n7610 = 1_n3636 & 1_n10341;
assign 1_n8342 = ~(1_n2476 | 1_n2510);
assign 1_n6182 = ~1_n6937;
assign 1_n1450 = ~(1_n2616 | 1_n5285);
assign 1_n1058 = ~1_n510;
assign 1_n1030 = ~1_n4017;
assign 1_n9160 = ~1_n12892;
assign 1_n2460 = ~(1_n9099 ^ 1_n245);
assign 1_n11202 = 1_n11236 & 1_n411;
assign 1_n1936 = ~1_n3566;
assign 1_n7634 = 1_n5733 | 1_n10474;
assign 1_n2960 = 1_n7038 | 1_n1833;
assign 1_n13090 = 1_n10112 | 1_n5076;
assign 1_n8282 = ~(1_n11804 ^ 1_n4548);
assign 1_n6328 = ~(1_n2659 ^ 1_n2736);
assign 1_n11086 = 1_n1747 & 1_n11423;
assign 1_n12118 = ~(1_n7637 ^ 1_n5038);
assign 1_n11493 = 1_n10857 | 1_n8793;
assign 1_n9002 = ~(1_n10796 | 1_n12058);
assign 1_n5078 = ~(1_n8292 ^ 1_n13090);
assign 1_n9238 = ~1_n469;
assign 1_n2684 = ~(1_n12974 ^ 1_n10038);
assign 1_n3862 = 1_n5490 & 1_n10740;
assign 1_n5075 = ~(1_n9324 ^ 1_n4090);
assign 1_n1840 = ~(1_n12873 | 1_n8756);
assign 1_n6844 = 1_n1323 | 1_n12062;
assign 1_n258 = 1_n3019 & 1_n11987;
assign 1_n1990 = 1_n2899 | 1_n11910;
assign 1_n4631 = ~(1_n1276 ^ 1_n184);
assign 1_n507 = 1_n2243 & 1_n4311;
assign 1_n2546 = 1_n7056 & 1_n7432;
assign 1_n6688 = 1_n12032 | 1_n8490;
assign 1_n7223 = ~1_n3677;
assign 1_n8352 = 1_n2530 & 1_n12473;
assign 1_n6422 = 1_n6881 | 1_n10702;
assign 1_n9146 = 1_n13190 | 1_n206;
assign 1_n1875 = 1_n4135 ^ 1_n12612;
assign 1_n11330 = 1_n9698 | 1_n4023;
assign 1_n10989 = ~1_n12939;
assign 1_n10013 = 1_n9429 | 1_n4640;
assign 1_n1371 = 1_n6934 & 1_n3871;
assign 1_n2875 = ~1_n11537;
assign 1_n12525 = 1_n7566 | 1_n2766;
assign 1_n1885 = ~1_n3977;
assign 1_n11172 = ~1_n4102;
assign 1_n5970 = ~1_n5786;
assign 1_n10823 = 1_n3957 & 1_n11273;
assign 1_n11372 = 1_n2449 | 1_n8490;
assign 1_n7158 = ~1_n6085;
assign 1_n4508 = 1_n8974 & 1_n10726;
assign 1_n2981 = ~(1_n1373 ^ 1_n10721);
assign 1_n7153 = 1_n7073 & 1_n1477;
assign 1_n5132 = 1_n10527 | 1_n11107;
assign 1_n12624 = ~1_n10238;
assign 1_n2976 = ~(1_n9502 ^ 1_n2719);
assign 1_n8374 = ~1_n510;
assign 1_n5686 = ~(1_n4171 ^ 1_n5173);
assign 1_n7077 = ~(1_n8279 | 1_n802);
assign 1_n145 = 1_n12058 & 1_n10796;
assign 1_n9575 = 1_n11996 & 1_n12650;
assign 1_n7670 = ~(1_n2006 ^ 1_n6325);
assign 1_n10741 = 1_n12775 | 1_n4359;
assign 1_n12715 = ~(1_n10671 ^ 1_n1927);
assign 1_n12934 = 1_n1791 & 1_n1886;
assign 1_n9067 = 1_n11614 & 1_n3536;
assign 1_n7247 = ~1_n5470;
assign 1_n373 = 1_n10824 | 1_n9923;
assign 1_n7137 = 1_n4361 & 1_n4563;
assign 1_n11021 = 1_n3458 & 1_n4475;
assign 1_n8643 = ~(1_n8923 | 1_n7479);
assign 1_n9804 = ~1_n11567;
assign 1_n1438 = ~1_n10594;
assign 1_n2162 = 1_n1513 | 1_n2298;
assign 1_n5489 = ~1_n5590;
assign 1_n7886 = 1_n12353 | 1_n8316;
assign 1_n10370 = 1_n6231 | 1_n12273;
assign 1_n4120 = ~(1_n10155 ^ 1_n11080);
assign 1_n2459 = ~(1_n2854 ^ 1_n2853);
assign 1_n8541 = 1_n10897 | 1_n1856;
assign 1_n10502 = 1_n8664 & 1_n10161;
assign 1_n3474 = ~(1_n4538 | 1_n12450);
assign 1_n1145 = ~1_n4681;
assign 1_n10555 = 1_n2614 | 1_n5076;
assign 1_n4044 = 1_n6823 & 1_n3255;
assign 1_n5753 = 1_n11515 & 1_n1542;
assign 1_n3574 = ~(1_n3131 | 1_n7627);
assign 1_n1734 = ~(1_n4706 ^ 1_n7851);
assign 1_n10305 = ~1_n7778;
assign 1_n7037 = 1_n10608 | 1_n3618;
assign 1_n11935 = ~(1_n10282 | 1_n5859);
assign 1_n6160 = ~1_n3774;
assign 1_n11476 = 1_n8384 | 1_n10098;
assign 1_n11912 = ~(1_n10328 | 1_n10366);
assign 1_n5889 = 1_n5773 & 1_n12600;
assign 1_n5524 = 1_n8120 & 1_n9334;
assign 1_n12102 = 1_n3110 ^ 1_n7083;
assign 1_n6607 = 1_n6046 & 1_n2333;
assign 1_n4637 = ~(1_n6844 | 1_n11085);
assign 1_n7612 = 1_n845 | 1_n9075;
assign 1_n3699 = 1_n6506 | 1_n7865;
assign 1_n10463 = ~(1_n12850 ^ 1_n2632);
assign 1_n9179 = ~(1_n3387 | 1_n12115);
assign 1_n2501 = 1_n10997 & 1_n3996;
assign 1_n9982 = ~(1_n6075 ^ 1_n10821);
assign 1_n11379 = ~1_n8291;
assign 1_n10948 = ~1_n10172;
assign 1_n12660 = 1_n11982 | 1_n10764;
assign 1_n1753 = ~(1_n4489 ^ 1_n10968);
assign 1_n8932 = 1_n2757 | 1_n6001;
assign 1_n6254 = 1_n6769 | 1_n12388;
assign 1_n12713 = ~1_n10378;
assign 1_n9950 = ~(1_n5371 ^ 1_n2441);
assign 1_n5836 = ~(1_n7527 | 1_n8913);
assign 1_n11910 = ~1_n951;
assign 1_n6105 = ~(1_n544 ^ 1_n6025);
assign 1_n5975 = ~(1_n5497 ^ 1_n1387);
assign 1_n10404 = ~(1_n5998 | 1_n3173);
assign 1_n7656 = 1_n7415 & 1_n3436;
assign 1_n337 = 1_n3647 | 1_n5098;
assign 1_n8031 = ~(1_n2798 ^ 1_n4670);
assign 1_n1842 = 1_n4808 | 1_n8534;
assign 1_n2280 = 1_n10422 & 1_n12773;
assign 1_n12659 = 1_n10471 | 1_n5242;
assign 1_n3056 = 1_n3900 | 1_n5443;
assign 1_n4712 = ~(1_n7534 ^ 1_n7212);
assign 1_n7086 = ~1_n8824;
assign 1_n2891 = 1_n2471 & 1_n165;
assign 1_n11348 = ~(1_n2475 ^ 1_n9574);
assign 1_n5963 = 1_n1261 | 1_n7935;
assign 1_n1735 = 1_n6770 | 1_n10319;
assign 1_n5853 = ~1_n5140;
assign 1_n7948 = ~(1_n1368 ^ 1_n10042);
assign 1_n12588 = ~(1_n215 | 1_n10629);
assign 1_n2577 = ~(1_n11845 ^ 1_n7057);
assign 1_n7858 = ~(1_n3480 ^ 1_n2859);
assign 1_n1046 = 1_n3539 & 1_n12446;
assign 1_n2565 = ~(1_n3980 ^ 1_n3714);
assign 1_n297 = 1_n6517 | 1_n6493;
assign 1_n12720 = 1_n4166 | 1_n1570;
assign 1_n215 = ~(1_n2024 | 1_n6508);
assign 1_n10994 = 1_n1989 | 1_n6770;
assign 1_n1986 = 1_n10889 & 1_n10498;
assign 1_n4720 = 1_n9637 | 1_n5188;
assign 1_n12184 = 1_n7783 | 1_n6265;
assign 1_n7393 = ~(1_n4345 ^ 1_n12570);
assign 1_n11237 = ~1_n6701;
assign 1_n2287 = ~1_n8230;
assign 1_n5232 = ~(1_n7896 ^ 1_n851);
assign 1_n4498 = ~1_n5546;
assign 1_n9151 = 1_n4638 & 1_n7453;
assign 1_n1434 = ~1_n8332;
assign 1_n9704 = 1_n867 & 1_n9326;
assign 1_n1876 = 1_n11548 | 1_n1985;
assign 1_n3817 = ~1_n2590;
assign 1_n3455 = ~(1_n4600 ^ 1_n1723);
assign 1_n12631 = ~(1_n7439 | 1_n10963);
assign 1_n6819 = ~(1_n12845 ^ 1_n13087);
assign 1_n6880 = 1_n13039 | 1_n2133;
assign 1_n5976 = 1_n1875 | 1_n12366;
assign 1_n2403 = ~1_n13121;
assign 1_n12400 = ~(1_n1774 | 1_n8413);
assign 1_n13155 = ~(1_n10547 ^ 1_n7689);
assign 1_n9897 = ~1_n4126;
assign 1_n12832 = 1_n3662 & 1_n6664;
assign 1_n12427 = 1_n3091 | 1_n2083;
assign 1_n1579 = ~1_n10075;
assign 1_n12838 = ~1_n10582;
assign 1_n7377 = ~1_n5962;
assign 1_n3692 = 1_n13025 | 1_n2059;
assign 1_n10872 = ~1_n4906;
assign 1_n12179 = 1_n11779 | 1_n7254;
assign 1_n11306 = ~(1_n5357 ^ 1_n3887);
assign 1_n713 = ~1_n6647;
assign 1_n5577 = 1_n9564 | 1_n5029;
assign 1_n6007 = ~(1_n6388 ^ 1_n6243);
assign 1_n236 = ~(1_n1334 ^ 1_n11176);
assign 1_n1309 = ~(1_n9066 ^ 1_n7681);
assign 1_n9172 = ~1_n2073;
assign 1_n5072 = 1_n9069 | 1_n8268;
assign 1_n4349 = 1_n4376 ^ 1_n11813;
assign 1_n1844 = ~(1_n7754 ^ 1_n775);
assign 1_n12598 = ~(1_n9922 ^ 1_n6031);
assign 1_n12439 = ~(1_n9083 ^ 1_n4390);
assign 1_n5554 = ~1_n748;
assign 1_n5001 = ~1_n8559;
assign 1_n5693 = 1_n12573 | 1_n4640;
assign 1_n9579 = ~(1_n6079 ^ 1_n1293);
assign 1_n11353 = ~(1_n7067 ^ 1_n5979);
assign 1_n6976 = 1_n6657 | 1_n265;
assign 1_n8897 = ~(1_n5693 ^ 1_n667);
assign 1_n12535 = ~1_n4042;
assign 1_n384 = ~(1_n12933 ^ 1_n6158);
assign 1_n1452 = 1_n8610 & 1_n12521;
assign 1_n7004 = ~(1_n2251 | 1_n665);
assign 1_n932 = 1_n5655 | 1_n2206;
assign 1_n5666 = ~1_n6392;
assign 1_n1035 = ~1_n353;
assign 1_n1603 = 1_n3570 & 1_n7898;
assign 1_n10281 = ~1_n1650;
assign 1_n4535 = ~(1_n300 ^ 1_n10619);
assign 1_n6677 = 1_n6956 ^ 1_n2583;
assign 1_n451 = 1_n11779 | 1_n4640;
assign 1_n11031 = ~(1_n5421 ^ 1_n11806);
assign 1_n11405 = ~(1_n3747 ^ 1_n999);
assign 1_n8093 = 1_n3550 | 1_n5059;
assign 1_n13133 = ~1_n7465;
assign 1_n4353 = 1_n1867 & 1_n1448;
assign 1_n11459 = 1_n161 | 1_n12328;
assign 1_n557 = ~(1_n12448 ^ 1_n7838);
assign 1_n6652 = ~1_n4645;
assign 1_n3861 = ~1_n3913;
assign 1_n10551 = 1_n10094 & 1_n147;
assign 1_n5645 = ~1_n10805;
assign 1_n2087 = ~(1_n9797 | 1_n12584);
assign 1_n3296 = ~(1_n7891 ^ 1_n6693);
assign 1_n315 = 1_n12585 & 1_n6315;
assign 1_n6678 = ~(1_n12235 ^ 1_n1253);
assign 1_n9800 = ~(1_n5933 ^ 1_n6670);
assign 1_n12953 = 1_n1035 | 1_n6732;
assign 1_n4261 = 1_n4974 | 1_n5076;
assign 1_n1654 = 1_n3587 | 1_n4947;
assign 1_n7279 = 1_n8139 & 1_n10606;
assign 1_n8520 = 1_n3316 & 1_n5411;
assign 1_n11273 = 1_n2639 | 1_n8490;
assign 1_n5206 = 1_n9131 | 1_n10871;
assign 1_n8165 = 1_n2109 | 1_n488;
assign 1_n6716 = ~1_n68;
assign 1_n4180 = 1_n983 | 1_n9177;
assign 1_n7914 = ~1_n8818;
assign 1_n4930 = 1_n8335 | 1_n2675;
assign 1_n1282 = ~(1_n11556 ^ 1_n3745);
assign 1_n6664 = 1_n12241 | 1_n9055;
assign 1_n9136 = ~(1_n9565 ^ 1_n4597);
assign 1_n735 = ~1_n1528;
assign 1_n4314 = 1_n4610 | 1_n479;
assign 1_n12166 = ~1_n11324;
assign 1_n6443 = ~(1_n12167 | 1_n2927);
assign 1_n7290 = 1_n72 ^ 1_n9250;
assign 1_n3113 = 1_n7780 | 1_n1144;
assign 1_n8099 = ~(1_n5327 | 1_n4421);
assign 1_n11959 = 1_n1311 & 1_n10853;
assign 1_n67 = ~(1_n3899 ^ 1_n4195);
assign 1_n7935 = 1_n9558;
assign 1_n1373 = 1_n8727 | 1_n6824;
assign 1_n8829 = 1_n2236 | 1_n5774;
assign 1_n10577 = 1_n13028 | 1_n6173;
assign 1_n1695 = ~1_n7720;
assign 1_n10151 = ~(1_n13188 ^ 1_n1288);
assign 1_n2042 = ~(1_n2486 | 1_n979);
assign 1_n7480 = ~1_n11129;
assign 1_n10021 = ~1_n11891;
assign 1_n5564 = 1_n11099 | 1_n10689;
assign 1_n9152 = 1_n10688 | 1_n10759;
assign 1_n2890 = ~1_n13058;
assign 1_n11366 = 1_n6751 | 1_n1463;
assign 1_n6078 = ~(1_n8476 | 1_n10027);
assign 1_n3999 = ~1_n5962;
assign 1_n5690 = ~(1_n7457 | 1_n3117);
assign 1_n10586 = ~1_n11411;
assign 1_n11971 = ~(1_n11199 ^ 1_n4601);
assign 1_n7244 = 1_n5166 & 1_n10536;
assign 1_n1601 = 1_n5616 | 1_n4055;
assign 1_n3810 = ~(1_n5763 ^ 1_n459);
assign 1_n4670 = ~(1_n7265 ^ 1_n12100);
assign 1_n12054 = 1_n8715 ^ 1_n6921;
assign 1_n8873 = 1_n3802 | 1_n12189;
assign 1_n1493 = ~1_n2169;
assign 1_n5556 = 1_n9904 ^ 1_n12915;
assign 1_n8090 = 1_n9079 & 1_n920;
assign 1_n8537 = 1_n5090 & 1_n7638;
assign 1_n7744 = ~(1_n1262 ^ 1_n5235);
assign 1_n10941 = ~1_n8422;
assign 1_n12573 = ~1_n11891;
assign 1_n12377 = ~1_n8798;
assign 1_n10478 = ~(1_n5556 ^ 1_n6073);
assign 1_n272 = 1_n9399 | 1_n13031;
assign 1_n3060 = 1_n11790 | 1_n7574;
assign 1_n9681 = ~1_n12810;
assign 1_n1369 = ~(1_n2289 ^ 1_n4569);
assign 1_n10145 = 1_n8457 | 1_n9972;
assign 1_n9287 = 1_n6922 | 1_n6635;
assign 1_n8171 = 1_n10287 | 1_n12847;
assign 1_n12652 = 1_n1447 | 1_n6404;
assign 1_n4586 = ~(1_n1233 ^ 1_n10632);
assign 1_n1291 = ~(1_n941 ^ 1_n4071);
assign 1_n6302 = 1_n6383 | 1_n1570;
assign 1_n4203 = ~1_n9841;
assign 1_n1334 = ~(1_n6167 ^ 1_n5981);
assign 1_n11695 = ~(1_n1742 | 1_n8475);
assign 1_n11813 = 1_n8466 & 1_n8506;
assign 1_n13120 = ~(1_n7752 ^ 1_n9274);
assign 1_n4795 = 1_n5561 | 1_n2315;
assign 1_n3687 = 1_n3331 | 1_n952;
assign 1_n5266 = ~(1_n13040 ^ 1_n859);
assign 1_n12309 = 1_n10492 | 1_n6138;
assign 1_n8769 = 1_n9298 | 1_n8127;
assign 1_n4542 = 1_n10929 | 1_n7723;
assign 1_n8437 = 1_n204 & 1_n5572;
assign 1_n8752 = ~(1_n5546 ^ 1_n13044);
assign 1_n8780 = 1_n8329 | 1_n5797;
assign 1_n10315 = 1_n980 & 1_n11297;
assign 1_n2717 = ~1_n10541;
assign 1_n5387 = 1_n842 & 1_n4274;
assign 1_n3515 = 1_n946 | 1_n12501;
assign 1_n6282 = ~(1_n1206 ^ 1_n2714);
assign 1_n612 = ~(1_n2743 | 1_n1620);
assign 1_n7320 = 1_n8142 & 1_n4443;
assign 1_n12047 = 1_n8759 | 1_n13148;
assign 1_n4112 = 1_n6495 & 1_n12315;
assign 1_n6174 = ~(1_n12151 ^ 1_n12540);
assign 1_n9924 = 1_n5271 | 1_n6404;
assign 1_n3001 = 1_n10411 | 1_n4208;
assign 1_n1194 = ~1_n8163;
assign 1_n5464 = ~(1_n12638 ^ 1_n736);
assign 1_n7578 = ~(1_n8538 | 1_n12200);
assign 1_n7188 = ~1_n510;
assign 1_n11472 = ~(1_n5913 ^ 1_n10379);
assign 1_n13173 = 1_n761 & 1_n3085;
assign 1_n8693 = ~1_n5307;
assign 1_n5793 = 1_n5107 | 1_n119;
assign 1_n12756 = 1_n8123 & 1_n3373;
assign 1_n8945 = ~(1_n3578 ^ 1_n4766);
assign 1_n4633 = ~(1_n12127 | 1_n5196);
assign 1_n6732 = 1_n8160;
assign 1_n8483 = ~(1_n3397 ^ 1_n11459);
assign 1_n7361 = 1_n6205 | 1_n425;
assign 1_n891 = 1_n12629 | 1_n4936;
assign 1_n1306 = 1_n12576 & 1_n7817;
assign 1_n7084 = ~1_n817;
assign 1_n8573 = ~(1_n12485 ^ 1_n1309);
assign 1_n9690 = 1_n11499 | 1_n10909;
assign 1_n9584 = 1_n9499 | 1_n1381;
assign 1_n1437 = ~1_n11376;
assign 1_n2331 = 1_n5809 | 1_n9759;
assign 1_n7883 = ~1_n10620;
assign 1_n3256 = 1_n3295 | 1_n4751;
assign 1_n1463 = 1_n3058;
assign 1_n1403 = ~(1_n10324 ^ 1_n7202);
assign 1_n13050 = ~(1_n9863 ^ 1_n11128);
assign 1_n11628 = ~1_n5920;
assign 1_n134 = ~(1_n68 ^ 1_n6246);
assign 1_n669 = ~(1_n8972 ^ 1_n6125);
assign 1_n7698 = ~(1_n2340 ^ 1_n1386);
assign 1_n6496 = 1_n7629 & 1_n3197;
assign 1_n5361 = 1_n11705 | 1_n11893;
assign 1_n9994 = 1_n10714 | 1_n10319;
assign 1_n6427 = ~(1_n2372 ^ 1_n9785);
assign 1_n823 = ~(1_n12660 ^ 1_n6435);
assign 1_n8317 = ~1_n3379;
assign 1_n11992 = ~(1_n9037 ^ 1_n7599);
assign 1_n12998 = ~1_n10873;
assign 1_n757 = ~1_n4417;
assign 1_n10475 = ~(1_n11676 ^ 1_n2483);
assign 1_n11143 = ~1_n8564;
assign 1_n9140 = 1_n6384 | 1_n10417;
assign 1_n5452 = 1_n12786 | 1_n8268;
assign 1_n8387 = 1_n10590 & 1_n10483;
assign 1_n956 = ~1_n10451;
assign 1_n8762 = 1_n8728 & 1_n4518;
assign 1_n10630 = ~(1_n9466 ^ 1_n13120);
assign 1_n10728 = ~(1_n12356 ^ 1_n3734);
assign 1_n9986 = 1_n3172 & 1_n1773;
assign 1_n4135 = 1_n4465 | 1_n4373;
assign 1_n6119 = 1_n7215 & 1_n249;
assign 1_n2115 = 1_n692 & 1_n12676;
assign 1_n2129 = ~1_n8860;
assign 1_n11641 = 1_n7772 & 1_n9531;
assign 1_n11572 = ~(1_n8180 ^ 1_n4872);
assign 1_n9872 = ~(1_n259 ^ 1_n10227);
assign 1_n5736 = 1_n2581 | 1_n12328;
assign 1_n12448 = 1_n11757 | 1_n8490;
assign 1_n8585 = ~1_n2758;
assign 1_n3142 = ~(1_n1608 ^ 1_n12398);
assign 1_n331 = 1_n11054 | 1_n12188;
assign 1_n4326 = 1_n8599 & 1_n6468;
assign 1_n9559 = 1_n6112 | 1_n7935;
assign 1_n2502 = ~(1_n11022 ^ 1_n3343);
assign 1_n1473 = ~(1_n12390 ^ 1_n1300);
assign 1_n7676 = 1_n4991 & 1_n10066;
assign 1_n774 = ~(1_n10949 ^ 1_n7122);
assign 1_n3947 = ~(1_n9956 ^ 1_n10775);
assign 1_n5523 = 1_n4080 | 1_n11300;
assign 1_n11861 = ~(1_n4866 ^ 1_n908);
assign 1_n3268 = ~(1_n112 ^ 1_n10003);
assign 1_n6352 = 1_n12114 & 1_n2186;
assign 1_n7296 = ~(1_n12601 ^ 1_n9036);
assign 1_n766 = ~(1_n9992 | 1_n10630);
assign 1_n5714 = ~1_n7183;
assign 1_n4504 = ~(1_n8137 | 1_n4740);
assign 1_n11650 = 1_n10381 | 1_n7824;
assign 1_n730 = 1_n7272 | 1_n3918;
assign 1_n11555 = 1_n5953 & 1_n12712;
assign 1_n10840 = ~(1_n6797 | 1_n3294);
assign 1_n7501 = 1_n9304 & 1_n6475;
assign 1_n12176 = 1_n1440 & 1_n8741;
assign 1_n7863 = ~(1_n888 ^ 1_n2765);
assign 1_n10512 = ~1_n3412;
assign 1_n3447 = 1_n1520 & 1_n10145;
assign 1_n6052 = ~1_n8319;
assign 1_n8811 = 1_n10577 ^ 1_n3995;
assign 1_n10898 = ~1_n1307;
assign 1_n1798 = 1_n11030 & 1_n9531;
assign 1_n5585 = ~(1_n5234 ^ 1_n11201);
assign 1_n7842 = ~(1_n10973 ^ 1_n2761);
assign 1_n8310 = 1_n9626 | 1_n130;
assign 1_n13084 = ~1_n5884;
assign 1_n5273 = ~(1_n12442 ^ 1_n9839);
assign 1_n3662 = 1_n8102 | 1_n5258;
assign 1_n6670 = 1_n1138 & 1_n8125;
assign 1_n9102 = 1_n10545 | 1_n11639;
assign 1_n12074 = ~(1_n6823 ^ 1_n9857);
assign 1_n8999 = 1_n3758 | 1_n164;
assign 1_n1113 = ~1_n4006;
assign 1_n4554 = ~(1_n1877 | 1_n1429);
assign 1_n8975 = 1_n6305 | 1_n984;
assign 1_n5472 = 1_n9150 & 1_n8743;
assign 1_n7305 = 1_n7566 & 1_n2766;
assign 1_n630 = 1_n5307 & 1_n4036;
assign 1_n4618 = ~1_n10946;
assign 1_n8916 = ~(1_n9648 ^ 1_n955);
assign 1_n8853 = 1_n7523 | 1_n7975;
assign 1_n2651 = 1_n9605 & 1_n1054;
assign 1_n2377 = 1_n10260 & 1_n5916;
assign 1_n6714 = 1_n1257 & 1_n6845;
assign 1_n7969 = 1_n4875 | 1_n12328;
assign 1_n2874 = ~(1_n4578 ^ 1_n4150);
assign 1_n4708 = 1_n906 & 1_n2056;
assign 1_n4178 = 1_n12552 | 1_n10213;
assign 1_n5380 = ~(1_n10023 ^ 1_n11042);
assign 1_n1204 = ~(1_n5918 ^ 1_n811);
assign 1_n11700 = ~1_n7491;
assign 1_n7797 = 1_n11751 | 1_n617;
assign 1_n4247 = ~(1_n12321 ^ 1_n5781);
assign 1_n6659 = 1_n8009 | 1_n6628;
assign 1_n3528 = 1_n7049 | 1_n8563;
assign 1_n11945 = 1_n3307 | 1_n5566;
assign 1_n11064 = ~(1_n2451 ^ 1_n9034);
assign 1_n8118 = 1_n3822 & 1_n3339;
assign 1_n9819 = 1_n8817 | 1_n9159;
assign 1_n13082 = ~1_n2174;
assign 1_n1362 = ~(1_n4968 ^ 1_n756);
assign 1_n4475 = 1_n13183 | 1_n177;
assign 1_n3666 = ~(1_n9269 ^ 1_n515);
assign 1_n4887 = ~(1_n12606 | 1_n7020);
assign 1_n5508 = 1_n10452 | 1_n6243;
assign 1_n8491 = ~1_n10979;
assign 1_n2489 = ~(1_n3959 | 1_n4286);
assign 1_n9077 = ~(1_n6852 ^ 1_n6307);
assign 1_n11494 = 1_n9546 & 1_n1087;
assign 1_n3990 = ~(1_n3606 | 1_n7869);
assign 1_n6093 = 1_n10351 & 1_n8448;
assign 1_n803 = ~1_n11990;
assign 1_n9442 = 1_n4855 | 1_n10319;
assign 1_n3418 = ~1_n3319;
assign 1_n9847 = 1_n8139 & 1_n12965;
assign 1_n10584 = 1_n1741 | 1_n9537;
assign 1_n9668 = ~1_n6826;
assign 1_n9114 = 1_n7498 & 1_n4225;
assign 1_n6290 = ~1_n1421;
assign 1_n12808 = ~1_n6607;
assign 1_n927 = ~(1_n12784 ^ 1_n6620);
assign 1_n4158 = 1_n1663 | 1_n2415;
assign 1_n6153 = ~(1_n5274 ^ 1_n11296);
assign 1_n10798 = ~1_n2295;
assign 1_n8900 = ~1_n818;
assign 1_n11326 = ~(1_n11414 ^ 1_n12354);
assign 1_n7847 = ~1_n10575;
assign 1_n10587 = ~1_n5729;
assign 1_n9777 = ~(1_n9796 ^ 1_n2040);
assign 1_n1399 = ~(1_n11125 ^ 1_n10249);
assign 1_n3746 = ~(1_n5711 ^ 1_n6895);
assign 1_n12193 = ~(1_n1137 ^ 1_n6899);
assign 1_n3148 = ~(1_n2053 | 1_n7834);
assign 1_n10538 = ~(1_n5509 ^ 1_n12875);
assign 1_n12257 = 1_n8732 | 1_n3882;
assign 1_n11062 = ~(1_n10640 ^ 1_n3382);
assign 1_n12679 = 1_n1634 | 1_n9745;
assign 1_n4792 = ~1_n10451;
assign 1_n5764 = ~(1_n8008 ^ 1_n12113);
assign 1_n9215 = 1_n5031 & 1_n510;
assign 1_n1624 = ~1_n5796;
assign 1_n5055 = 1_n5568 & 1_n5729;
assign 1_n3117 = 1_n2582 | 1_n2816;
assign 1_n9411 = 1_n6416 | 1_n9075;
assign 1_n8739 = ~1_n4978;
assign 1_n9612 = 1_n7748 | 1_n4373;
assign 1_n11561 = ~(1_n5306 ^ 1_n7428);
assign 1_n9196 = ~(1_n4263 ^ 1_n11816);
assign 1_n7156 = 1_n8776 | 1_n6769;
assign 1_n2560 = ~(1_n2049 ^ 1_n7917);
assign 1_n4103 = 1_n12236 | 1_n4835;
assign 1_n4629 = 1_n6215 | 1_n10433;
assign 1_n4013 = ~1_n2057;
assign 1_n2255 = 1_n10248 & 1_n5369;
assign 1_n12725 = 1_n5826 & 1_n2831;
assign 1_n7719 = ~1_n7439;
assign 1_n5060 = ~(1_n9048 ^ 1_n6105);
assign 1_n3204 = 1_n3634 | 1_n1043;
assign 1_n12569 = 1_n11117 | 1_n8445;
assign 1_n3878 = 1_n3176 | 1_n10652;
assign 1_n3696 = ~1_n1432;
assign 1_n3937 = 1_n4475 | 1_n3458;
assign 1_n5252 = 1_n10153 | 1_n3650;
assign 1_n4711 = ~(1_n9955 ^ 1_n3562);
assign 1_n4303 = 1_n1719 ^ 1_n2423;
assign 1_n2006 = 1_n5671 & 1_n8506;
assign 1_n11995 = 1_n3922 & 1_n2428;
assign 1_n1086 = ~(1_n31 ^ 1_n8872);
assign 1_n12964 = 1_n11960 | 1_n9075;
assign 1_n2044 = ~(1_n5451 ^ 1_n7569);
assign 1_n9874 = ~(1_n6151 | 1_n5033);
assign 1_n6904 = ~(1_n11692 ^ 1_n7309);
assign 1_n7743 = 1_n1087 | 1_n9546;
assign 1_n1002 = 1_n1909 | 1_n3955;
assign 1_n7987 = 1_n4739 | 1_n4675;
assign 1_n3923 = ~(1_n7875 ^ 1_n4856);
assign 1_n9131 = ~1_n1302;
assign 1_n1865 = ~(1_n9423 | 1_n3206);
assign 1_n11786 = 1_n7062 | 1_n12273;
assign 1_n12977 = ~(1_n11168 ^ 1_n13105);
assign 1_n6414 = 1_n7042 | 1_n9078;
assign 1_n6525 = 1_n803 & 1_n8558;
assign 1_n3889 = ~(1_n5678 ^ 1_n8684);
assign 1_n7009 = ~1_n10457;
assign 1_n1697 = ~1_n1938;
assign 1_n8428 = ~1_n10398;
assign 1_n2574 = ~(1_n7529 | 1_n7715);
assign 1_n931 = 1_n4564 | 1_n3949;
assign 1_n10071 = ~(1_n9903 ^ 1_n3644);
assign 1_n7309 = 1_n542 | 1_n11668;
assign 1_n10995 = ~(1_n4057 ^ 1_n10994);
assign 1_n4450 = 1_n6029 & 1_n2179;
assign 1_n10465 = ~1_n7659;
assign 1_n11474 = ~(1_n7330 ^ 1_n11760);
assign 1_n5428 = 1_n7142 | 1_n6265;
assign 1_n7556 = 1_n812 & 1_n9717;
assign 1_n16 = ~1_n12348;
assign 1_n7540 = ~(1_n8827 ^ 1_n6378);
assign 1_n3123 = ~(1_n10828 ^ 1_n5651);
assign 1_n807 = ~(1_n3274 ^ 1_n49);
assign 1_n6515 = 1_n4908 & 1_n11545;
assign 1_n2544 = 1_n8640;
assign 1_n6034 = 1_n1453 & 1_n8216;
assign 1_n10218 = ~(1_n2054 ^ 1_n4575);
assign 1_n10038 = 1_n5893 & 1_n3124;
assign 1_n6407 = ~1_n834;
assign 1_n4048 = ~(1_n8483 ^ 1_n3881);
assign 1_n10482 = 1_n13071 & 1_n2419;
assign 1_n1864 = 1_n6967 | 1_n12328;
assign 1_n8008 = 1_n1511 | 1_n1026;
assign 1_n2146 = 1_n1544 & 1_n7611;
assign 1_n8450 = ~(1_n5568 | 1_n8308);
assign 1_n13067 = 1_n8020 | 1_n7530;
assign 1_n6891 = ~(1_n8141 ^ 1_n11510);
assign 1_n6695 = ~(1_n8559 ^ 1_n1623);
assign 1_n7618 = 1_n80 | 1_n1571;
assign 1_n9433 = ~(1_n8224 ^ 1_n7449);
assign 1_n2234 = 1_n2155 & 1_n6291;
assign 1_n6813 = 1_n6587 | 1_n2675;
assign 1_n994 = 1_n2188 & 1_n3265;
assign 1_n3434 = ~(1_n7038 ^ 1_n10621);
assign 1_n7398 = ~(1_n4210 ^ 1_n1473);
assign 1_n1497 = 1_n7146 | 1_n8030;
assign 1_n6475 = 1_n6244 | 1_n9043;
assign 1_n12747 = ~1_n11518;
assign 1_n12103 = ~(1_n4393 ^ 1_n4073);
assign 1_n3402 = ~(1_n2360 ^ 1_n9128);
assign 1_n8575 = ~(1_n5494 | 1_n9578);
assign 1_n11672 = 1_n3969 | 1_n10945;
assign 1_n2503 = 1_n6566 | 1_n155;
assign 1_n11961 = ~(1_n2887 ^ 1_n8244);
assign 1_n5359 = ~1_n5030;
assign 1_n11012 = ~(1_n3549 ^ 1_n11151);
assign 1_n9385 = ~(1_n3152 | 1_n4815);
assign 1_n397 = ~(1_n3401 ^ 1_n1555);
assign 1_n7415 = ~1_n1157;
assign 1_n9306 = ~(1_n5292 | 1_n8213);
assign 1_n9180 = 1_n6740 | 1_n4837;
assign 1_n5540 = ~1_n9777;
assign 1_n3242 = ~(1_n1277 ^ 1_n11627);
assign 1_n3032 = 1_n2449 | 1_n12388;
assign 1_n2511 = ~(1_n3223 ^ 1_n1518);
assign 1_n10109 = ~1_n13220;
assign 1_n4588 = 1_n5466 | 1_n11025;
assign 1_n5109 = 1_n6118 | 1_n5384;
assign 1_n9660 = 1_n13128 | 1_n10858;
assign 1_n11720 = ~(1_n3414 | 1_n5708);
assign 1_n9981 = 1_n6602 & 1_n9255;
assign 1_n6233 = ~(1_n4579 | 1_n4763);
assign 1_n12825 = 1_n5854 | 1_n13172;
assign 1_n11300 = ~1_n10770;
assign 1_n5473 = ~(1_n7289 | 1_n9285);
assign 1_n9987 = 1_n1208 | 1_n7264;
assign 1_n9717 = 1_n5341 & 1_n9108;
assign 1_n3706 = 1_n8696 | 1_n12351;
assign 1_n3401 = ~(1_n12090 ^ 1_n5534);
assign 1_n4435 = ~(1_n10469 ^ 1_n4404);
assign 1_n8870 = ~(1_n1753 ^ 1_n1915);
assign 1_n5480 = 1_n11582 ^ 1_n751;
assign 1_n3609 = 1_n10533 | 1_n12919;
assign 1_n10655 = 1_n2506 & 1_n5093;
assign 1_n740 = ~1_n3511;
assign 1_n11859 = 1_n3208 | 1_n8268;
assign 1_n1972 = 1_n7188 | 1_n5797;
assign 1_n4437 = ~(1_n1003 ^ 1_n4733);
assign 1_n2541 = ~1_n10343;
assign 1_n6540 = 1_n6733 | 1_n8702;
assign 1_n10012 = 1_n2168 & 1_n1445;
assign 1_n12051 = 1_n10604 | 1_n1516;
assign 1_n1209 = 1_n10670 & 1_n5172;
assign 1_n7118 = ~(1_n13136 ^ 1_n702);
assign 1_n7979 = 1_n8940 & 1_n8233;
assign 1_n10152 = 1_n1188 | 1_n8348;
assign 1_n7294 = ~(1_n4052 ^ 1_n6616);
assign 1_n3639 = ~1_n9820;
assign 1_n10727 = ~1_n10024;
assign 1_n1730 = ~(1_n12946 | 1_n2508);
assign 1_n3464 = 1_n2272 & 1_n4704;
assign 1_n2366 = ~(1_n6476 ^ 1_n555);
assign 1_n890 = 1_n3456 & 1_n5355;
assign 1_n6641 = ~(1_n7094 ^ 1_n1086);
assign 1_n4755 = 1_n9557 | 1_n2958;
assign 1_n10766 = ~(1_n948 ^ 1_n9211);
assign 1_n6683 = ~(1_n2697 ^ 1_n12160);
assign 1_n10631 = 1_n10001 | 1_n5209;
assign 1_n11076 = ~(1_n9193 ^ 1_n2797);
assign 1_n700 = ~(1_n13188 | 1_n1288);
assign 1_n2169 = 1_n11165 & 1_n3201;
assign 1_n3067 = 1_n13151 & 1_n2598;
assign 1_n11872 = 1_n80 | 1_n542;
assign 1_n7830 = 1_n10170 & 1_n12221;
assign 1_n366 = ~(1_n141 ^ 1_n607);
assign 1_n7753 = 1_n2702 & 1_n5057;
assign 1_n8057 = ~(1_n2774 | 1_n67);
assign 1_n629 = 1_n6126 | 1_n2627;
assign 1_n11011 = ~(1_n9664 | 1_n6047);
assign 1_n3803 = ~(1_n1048 | 1_n9106);
assign 1_n10750 = 1_n7510 & 1_n3812;
assign 1_n10983 = ~(1_n3267 ^ 1_n33);
assign 1_n1349 = ~1_n3682;
assign 1_n1984 = 1_n4385 | 1_n7930;
assign 1_n7570 = 1_n7355 | 1_n9259;
assign 1_n11401 = ~(1_n9829 ^ 1_n423);
assign 1_n7078 = 1_n973 | 1_n2281;
assign 1_n6436 = 1_n11122 | 1_n8268;
assign 1_n2696 = 1_n946 | 1_n479;
assign 1_n11414 = 1_n1422 | 1_n2059;
assign 1_n214 = ~(1_n32 | 1_n4020);
assign 1_n12574 = 1_n12211 & 1_n3775;
assign 1_n1957 = ~1_n744;
assign 1_n11907 = ~(1_n12650 ^ 1_n11996);
assign 1_n3910 = 1_n1638 | 1_n12188;
assign 1_n1495 = 1_n10057 | 1_n4947;
assign 1_n2892 = ~(1_n8310 ^ 1_n3081);
assign 1_n5300 = ~(1_n11597 ^ 1_n1483);
assign 1_n3346 = ~(1_n5590 ^ 1_n12935);
assign 1_n1275 = ~(1_n8144 ^ 1_n1666);
assign 1_n12167 = 1_n12203 | 1_n3949;
assign 1_n2995 = 1_n5177 & 1_n8098;
assign 1_n7903 = ~1_n9620;
assign 1_n8929 = ~(1_n4331 | 1_n1151);
assign 1_n5348 = ~1_n9241;
assign 1_n2172 = ~(1_n12233 ^ 1_n8105);
assign 1_n9953 = 1_n8580 & 1_n6242;
assign 1_n10835 = 1_n11446 | 1_n3949;
assign 1_n7579 = 1_n6728 & 1_n2027;
assign 1_n130 = 1_n7433 & 1_n9107;
assign 1_n4123 = ~(1_n3113 ^ 1_n1250);
assign 1_n3445 = ~1_n9362;
assign 1_n3680 = ~(1_n4388 ^ 1_n11246);
assign 1_n13079 = 1_n8517 & 1_n11187;
assign 1_n1518 = ~(1_n9524 ^ 1_n2947);
assign 1_n2520 = 1_n6865 | 1_n5792;
assign 1_n6591 = 1_n6686 | 1_n6786;
assign 1_n13114 = ~(1_n6679 ^ 1_n9573);
assign 1_n3763 = ~(1_n3016 ^ 1_n4501);
assign 1_n11517 = 1_n12916 | 1_n657;
assign 1_n3160 = 1_n11979 | 1_n9360;
assign 1_n4861 = ~(1_n7924 ^ 1_n7994);
assign 1_n5324 = 1_n958 & 1_n11681;
assign 1_n8036 = 1_n10903 & 1_n5215;
assign 1_n10273 = 1_n10276 & 1_n12183;
assign 1_n479 = 1_n917;
assign 1_n4536 = ~1_n8183;
assign 1_n8656 = ~(1_n12947 | 1_n9568);
assign 1_n1070 = ~1_n9297;
assign 1_n11144 = 1_n6274;
assign 1_n10418 = 1_n11308 & 1_n9321;
assign 1_n6124 = ~(1_n1892 ^ 1_n4297);
assign 1_n8603 = ~(1_n989 ^ 1_n11575);
assign 1_n9886 = ~(1_n11844 | 1_n9076);
assign 1_n12942 = ~(1_n6686 ^ 1_n2760);
assign 1_n7867 = 1_n8890 | 1_n5955;
assign 1_n10686 = 1_n10802 & 1_n2785;
assign 1_n6772 = 1_n11310 | 1_n6827;
assign 1_n3129 = 1_n5945 & 1_n2950;
assign 1_n3977 = 1_n7847 & 1_n5170;
assign 1_n2213 = ~1_n6532;
assign 1_n8742 = ~(1_n4563 ^ 1_n1228);
assign 1_n11349 = ~(1_n4432 ^ 1_n6119);
assign 1_n12962 = ~(1_n9095 ^ 1_n11103);
assign 1_n10118 = ~(1_n7633 ^ 1_n77);
assign 1_n1203 = ~(1_n2495 ^ 1_n9246);
assign 1_n7940 = 1_n6854 | 1_n8754;
assign 1_n152 = 1_n12882 | 1_n8268;
assign 1_n1899 = 1_n2912 & 1_n672;
assign 1_n5944 = 1_n8499 | 1_n1144;
assign 1_n5477 = ~(1_n6337 ^ 1_n10881);
assign 1_n11451 = 1_n10293 | 1_n2038;
assign 1_n2181 = 1_n3622 & 1_n7230;
assign 1_n3664 = 1_n2176 & 1_n881;
assign 1_n10186 = 1_n1437 & 1_n10200;
assign 1_n11133 = 1_n9145 & 1_n6036;
assign 1_n12891 = ~(1_n1227 | 1_n4024);
assign 1_n3403 = ~(1_n4821 ^ 1_n4268);
assign 1_n4237 = ~1_n11324;
assign 1_n6841 = ~1_n8139;
assign 1_n3495 = ~(1_n4735 ^ 1_n2972);
assign 1_n6285 = 1_n5803 & 1_n3193;
assign 1_n2058 = 1_n10117 & 1_n10005;
assign 1_n2043 = ~(1_n3135 ^ 1_n4989);
assign 1_n7991 = 1_n3727 | 1_n118;
assign 1_n8745 = ~(1_n5776 ^ 1_n9457);
assign 1_n3419 = ~1_n9134;
assign 1_n7018 = 1_n10977 | 1_n5797;
assign 1_n9960 = 1_n10861 & 1_n5071;
assign 1_n2818 = 1_n13082 | 1_n8534;
assign 1_n4566 = ~1_n11774;
assign 1_n5385 = 1_n9917 | 1_n2943;
assign 1_n2243 = 1_n436 | 1_n9453;
assign 1_n9671 = 1_n9335 | 1_n8524;
assign 1_n3912 = ~(1_n1411 | 1_n476);
assign 1_n2784 = ~(1_n954 | 1_n1996);
assign 1_n5906 = ~(1_n630 | 1_n12753);
assign 1_n2124 = 1_n7230 | 1_n3622;
assign 1_n8885 = 1_n4143 | 1_n9195;
assign 1_n9043 = ~1_n2820;
assign 1_n1783 = ~1_n12284;
assign 1_n7140 = ~(1_n2094 | 1_n738);
assign 1_n11325 = 1_n7315 & 1_n238;
assign 1_n4099 = 1_n3401 | 1_n9233;
assign 1_n2690 = ~(1_n2676 ^ 1_n6868);
assign 1_n3488 = 1_n8405 & 1_n936;
assign 1_n12453 = ~(1_n2365 ^ 1_n9007);
assign 1_n34 = 1_n7842 | 1_n176;
assign 1_n2988 = 1_n1327 | 1_n9375;
assign 1_n2880 = ~1_n2762;
assign 1_n5283 = ~(1_n3382 | 1_n10640);
assign 1_n9012 = 1_n5901 & 1_n12119;
assign 1_n8467 = 1_n9382 & 1_n10361;
assign 1_n4985 = 1_n5565 | 1_n9195;
assign 1_n10185 = ~(1_n13104 ^ 1_n8566);
assign 1_n9194 = ~(1_n2409 ^ 1_n6358);
assign 1_n5997 = 1_n2158 & 1_n11271;
assign 1_n9750 = 1_n7700 | 1_n1570;
assign 1_n12940 = ~1_n9981;
assign 1_n2333 = 1_n6942 & 1_n13240;
assign 1_n11432 = 1_n6501 & 1_n272;
assign 1_n6742 = 1_n7277 | 1_n5378;
assign 1_n5661 = 1_n12709 | 1_n431;
assign 1_n2989 = 1_n4652 & 1_n9700;
assign 1_n8709 = ~(1_n1230 ^ 1_n9699);
assign 1_n2140 = ~(1_n9585 | 1_n3766);
assign 1_n2247 = ~(1_n6850 ^ 1_n8553);
assign 1_n5866 = ~(1_n12591 ^ 1_n10047);
assign 1_n8588 = ~(1_n3423 ^ 1_n2357);
assign 1_n6642 = ~(1_n136 ^ 1_n9744);
assign 1_n339 = 1_n7699 & 1_n8703;
assign 1_n11787 = 1_n10077 | 1_n4994;
assign 1_n10928 = 1_n6575 | 1_n9504;
assign 1_n4899 = 1_n2091 & 1_n3597;
assign 1_n9261 = ~(1_n4752 ^ 1_n10561);
assign 1_n8904 = ~1_n12853;
assign 1_n6425 = 1_n5161 & 1_n9119;
assign 1_n13153 = ~(1_n11504 | 1_n10262);
assign 1_n640 = ~1_n405;
assign 1_n5229 = ~1_n4315;
assign 1_n6571 = 1_n11149 | 1_n8352;
assign 1_n6522 = 1_n10352 | 1_n11107;
assign 1_n2285 = 1_n1047 & 1_n963;
assign 1_n9738 = 1_n11829 & 1_n6940;
assign 1_n5434 = ~1_n7726;
assign 1_n3051 = 1_n45 | 1_n8563;
assign 1_n2958 = 1_n12954;
assign 1_n6722 = 1_n4564 | 1_n6370;
assign 1_n1160 = 1_n7044 & 1_n12368;
assign 1_n6983 = ~1_n9885;
assign 1_n10380 = ~1_n465;
assign 1_n11776 = ~(1_n9205 ^ 1_n5425);
assign 1_n12092 = ~1_n12715;
assign 1_n5440 = 1_n899 | 1_n11107;
assign 1_n665 = 1_n8252 & 1_n3120;
assign 1_n11691 = ~(1_n6927 ^ 1_n3107);
assign 1_n5689 = ~(1_n4912 ^ 1_n7773);
assign 1_n8538 = 1_n5961 & 1_n4244;
assign 1_n9795 = ~1_n12269;
assign 1_n8838 = 1_n8460 & 1_n2291;
assign 1_n10480 = 1_n5351 | 1_n12659;
assign 1_n9489 = ~1_n8468;
assign 1_n4418 = 1_n9450 | 1_n1570;
assign 1_n3412 = ~1_n11248;
assign 1_n11200 = 1_n695 & 1_n7483;
assign 1_n9898 = 1_n1246 & 1_n10597;
assign 1_n3501 = 1_n12795 | 1_n8702;
assign 1_n7992 = ~(1_n9207 ^ 1_n12207);
assign 1_n2277 = 1_n500 & 1_n13241;
assign 1_n6209 = 1_n1972 ^ 1_n10015;
assign 1_n1262 = ~(1_n4805 ^ 1_n909);
assign 1_n4487 = ~1_n9904;
assign 1_n12961 = ~(1_n10511 ^ 1_n706);
assign 1_n779 = ~(1_n8731 | 1_n3175);
assign 1_n7198 = ~(1_n6717 | 1_n9812);
assign 1_n10036 = 1_n489 & 1_n12206;
assign 1_n3440 = ~(1_n3309 | 1_n4513);
assign 1_n6996 = 1_n2292 & 1_n2362;
assign 1_n5085 = 1_n7774 | 1_n11355;
assign 1_n4495 = ~1_n6168;
assign 1_n5831 = ~(1_n4924 | 1_n4919);
assign 1_n7665 = 1_n3978 | 1_n8270;
assign 1_n5611 = ~1_n7659;
assign 1_n4518 = 1_n8228 & 1_n6085;
assign 1_n1065 = 1_n1152 | 1_n1463;
assign 1_n8814 = ~(1_n12608 ^ 1_n7310);
assign 1_n8986 = 1_n5159 & 1_n10496;
assign 1_n8549 = ~(1_n1107 ^ 1_n9541);
assign 1_n12044 = 1_n12741 | 1_n13086;
assign 1_n7701 = 1_n12754 & 1_n11714;
assign 1_n5652 = ~(1_n7728 | 1_n9804);
assign 1_n189 = ~1_n103;
assign 1_n3583 = 1_n1017 | 1_n8281;
assign 1_n543 = 1_n9348 & 1_n4271;
assign 1_n3894 = ~1_n7436;
assign 1_n2709 = ~(1_n6987 ^ 1_n6646);
assign 1_n7440 = 1_n2090 & 1_n3834;
assign 1_n7620 = ~1_n4748;
assign 1_n4569 = ~(1_n3417 ^ 1_n12432);
assign 1_n4264 = ~(1_n7023 ^ 1_n11497);
assign 1_n9147 = 1_n4358 & 1_n6268;
assign 1_n12633 = 1_n9385 | 1_n670;
assign 1_n6960 = ~1_n6535;
assign 1_n12132 = 1_n5666 | 1_n2133;
assign 1_n8982 = 1_n10208 | 1_n8683;
assign 1_n8296 = 1_n3111 | 1_n11169;
assign 1_n3851 = 1_n9411 | 1_n7440;
assign 1_n5592 = 1_n8028 | 1_n2746;
assign 1_n8133 = 1_n2183 | 1_n12695;
assign 1_n560 = ~1_n353;
assign 1_n1681 = 1_n136 | 1_n5816;
assign 1_n3305 = ~(1_n6203 ^ 1_n763);
assign 1_n11104 = 1_n4948 | 1_n11362;
assign 1_n5691 = ~(1_n1034 ^ 1_n12925);
assign 1_n12382 = 1_n2090 | 1_n3834;
assign 1_n12623 = ~1_n9620;
assign 1_n7453 = 1_n1508 | 1_n5454;
assign 1_n6111 = 1_n115 | 1_n479;
assign 1_n3787 = ~(1_n6213 ^ 1_n7144);
assign 1_n2066 = 1_n11519 | 1_n5242;
assign 1_n6947 = 1_n700 | 1_n6284;
assign 1_n5622 = ~(1_n3188 | 1_n4002);
assign 1_n11573 = ~(1_n9500 | 1_n1492);
assign 1_n4018 = ~(1_n11715 | 1_n5289);
assign 1_n1961 = 1_n5983 & 1_n5370;
assign 1_n6864 = 1_n4714 & 1_n3690;
assign 1_n5792 = ~(1_n8357 | 1_n8134);
assign 1_n10202 = 1_n7892 & 1_n11599;
assign 1_n5272 = ~(1_n6453 ^ 1_n11647);
assign 1_n7513 = ~(1_n3868 ^ 1_n8564);
assign 1_n4868 = ~(1_n11230 | 1_n799);
assign 1_n122 = 1_n5423 | 1_n8348;
assign 1_n2059 = 1_n11148;
assign 1_n5101 = ~(1_n547 ^ 1_n8676);
assign 1_n8167 = 1_n7299 | 1_n4082;
assign 1_n10407 = 1_n6374 & 1_n3933;
assign 1_n1992 = ~(1_n6014 ^ 1_n5754);
assign 1_n6889 = ~1_n828;
assign 1_n3106 = 1_n10113 & 1_n2252;
assign 1_n2705 = 1_n12215 & 1_n10220;
assign 1_n12035 = ~(1_n5027 ^ 1_n9446);
assign 1_n11327 = ~(1_n8550 ^ 1_n1114);
assign 1_n1013 = 1_n8386 & 1_n615;
assign 1_n7400 = 1_n1538 & 1_n641;
assign 1_n2518 = 1_n13117 | 1_n2387;
assign 1_n8278 = 1_n7461 & 1_n8148;
assign 1_n9596 = ~1_n13138;
assign 1_n13037 = 1_n13216 & 1_n6502;
assign 1_n7491 = 1_n9978 & 1_n4322;
assign 1_n10393 = ~(1_n3845 ^ 1_n1215);
assign 1_n10799 = ~(1_n549 ^ 1_n4441);
assign 1_n2798 = 1_n4744 & 1_n10244;
assign 1_n2304 = 1_n13047 & 1_n8394;
assign 1_n2679 = 1_n1319 & 1_n3984;
assign 1_n3642 = 1_n4440 & 1_n8846;
assign 1_n6590 = ~1_n4470;
assign 1_n1504 = 1_n871 | 1_n8514;
assign 1_n7066 = ~(1_n11725 ^ 1_n3052);
assign 1_n11915 = 1_n12617 | 1_n8702;
assign 1_n2965 = 1_n6918 & 1_n4061;
assign 1_n8002 = ~1_n2310;
assign 1_n3873 = ~(1_n9601 ^ 1_n8934);
assign 1_n7414 = 1_n10402 | 1_n3981;
assign 1_n8952 = 1_n4827 | 1_n2240;
assign 1_n5808 = 1_n11990 ^ 1_n8558;
assign 1_n9197 = ~(1_n9084 ^ 1_n12744);
assign 1_n10010 = ~1_n11266;
assign 1_n3771 = ~(1_n4867 ^ 1_n10995);
assign 1_n11730 = ~(1_n12022 | 1_n10316);
assign 1_n1976 = ~1_n1190;
assign 1_n3416 = 1_n618 & 1_n9858;
assign 1_n8946 = 1_n9696 | 1_n11011;
assign 1_n4657 = ~1_n8332;
assign 1_n8447 = 1_n13137 | 1_n5130;
assign 1_n11125 = 1_n11242 | 1_n5797;
assign 1_n4315 = 1_n6320 & 1_n127;
assign 1_n8488 = 1_n75 | 1_n7530;
assign 1_n10458 = 1_n12921 & 1_n9600;
assign 1_n9243 = ~(1_n7126 | 1_n2227);
assign 1_n2903 = ~(1_n8461 ^ 1_n6007);
assign 1_n2055 = ~1_n10463;
assign 1_n11612 = ~1_n817;
assign 1_n12472 = 1_n1194 | 1_n2675;
assign 1_n12258 = ~1_n295;
assign 1_n320 = ~1_n8432;
assign 1_n941 = ~(1_n2230 ^ 1_n11726);
assign 1_n4000 = ~(1_n8931 ^ 1_n10416);
assign 1_n10892 = ~1_n1313;
assign 1_n11232 = ~1_n10442;
assign 1_n12897 = 1_n12023 | 1_n2449;
assign 1_n12237 = 1_n7963 & 1_n3334;
assign 1_n13209 = 1_n8443 & 1_n132;
assign 1_n10209 = ~(1_n1491 ^ 1_n1109);
assign 1_n3593 = ~(1_n257 ^ 1_n4190);
assign 1_n4469 = 1_n910 & 1_n178;
assign 1_n3657 = 1_n11212 | 1_n206;
assign 1_n4642 = ~1_n11666;
assign 1_n251 = ~(1_n3249 ^ 1_n10403);
assign 1_n10257 = ~(1_n13018 | 1_n355);
assign 1_n4893 = 1_n11514 | 1_n11244;
assign 1_n12460 = ~(1_n2076 ^ 1_n8390);
assign 1_n1442 = 1_n6922 | 1_n4724;
assign 1_n6226 = 1_n12997 | 1_n5797;
assign 1_n13145 = 1_n9008 & 1_n3118;
assign 1_n4488 = ~1_n10821;
assign 1_n7839 = ~1_n4033;
assign 1_n4416 = ~(1_n8605 | 1_n112);
assign 1_n11722 = 1_n5806 | 1_n3981;
assign 1_n203 = 1_n6337 | 1_n10881;
assign 1_n2369 = ~(1_n11671 ^ 1_n9062);
assign 1_n1804 = ~(1_n1134 | 1_n3283);
assign 1_n7800 = ~(1_n11304 | 1_n4463);
assign 1_n4200 = ~(1_n9494 | 1_n2996);
assign 1_n1846 = 1_n3530 | 1_n5676;
assign 1_n755 = ~1_n8820;
assign 1_n2773 = ~1_n1756;
assign 1_n9056 = ~(1_n4641 | 1_n6817);
assign 1_n4986 = ~(1_n5504 ^ 1_n5732);
assign 1_n1192 = 1_n12027 & 1_n11502;
assign 1_n10287 = ~1_n4075;
assign 1_n12613 = 1_n1224 | 1_n7781;
assign 1_n5921 = ~1_n925;
assign 1_n7626 = ~(1_n7806 | 1_n11290);
assign 1_n10357 = ~(1_n9293 ^ 1_n6400);
assign 1_n13048 = ~(1_n12293 ^ 1_n2907);
assign 1_n9517 = 1_n12599 | 1_n941;
assign 1_n12566 = 1_n6073 & 1_n4544;
assign 1_n31 = ~(1_n1789 ^ 1_n2908);
assign 1_n8536 = ~(1_n8205 ^ 1_n11834);
assign 1_n10486 = ~(1_n4328 | 1_n12320);
assign 1_n1205 = ~(1_n7156 ^ 1_n4843);
assign 1_n4300 = 1_n3820 & 1_n4308;
assign 1_n7837 = ~1_n2771;
assign 1_n4750 = 1_n11612 | 1_n7935;
assign 1_n6827 = 1_n5301 & 1_n422;
assign 1_n11258 = 1_n11431 | 1_n4435;
assign 1_n2134 = 1_n383 | 1_n11899;
assign 1_n1075 = 1_n767 & 1_n2498;
assign 1_n3042 = ~(1_n1917 ^ 1_n9777);
assign 1_n12358 = 1_n2722 & 1_n2146;
assign 1_n1277 = ~(1_n8799 ^ 1_n1665);
assign 1_n13126 = 1_n11226 | 1_n4640;
assign 1_n11549 = 1_n11450 & 1_n4757;
assign 1_n7993 = ~(1_n7876 ^ 1_n3692);
assign 1_n12378 = ~1_n5161;
assign 1_n7312 = ~1_n12538;
assign 1_n4516 = 1_n10560 & 1_n1636;
assign 1_n9024 = ~(1_n6867 ^ 1_n2454);
assign 1_n2391 = 1_n8527 & 1_n2143;
assign 1_n3458 = ~(1_n11159 ^ 1_n3952);
assign 1_n11883 = ~(1_n11702 | 1_n11710);
assign 1_n9761 = ~1_n834;
assign 1_n12873 = 1_n10876 & 1_n3645;
assign 1_n495 = 1_n2701 | 1_n10029;
assign 1_n5275 = 1_n6723 & 1_n2327;
assign 1_n4981 = 1_n10047 & 1_n12591;
assign 1_n3168 = 1_n13201 & 1_n3815;
assign 1_n2854 = 1_n10814 | 1_n11668;
assign 1_n12277 = ~(1_n12765 ^ 1_n11346);
assign 1_n7373 = ~(1_n437 ^ 1_n10028);
assign 1_n952 = 1_n6676 & 1_n9869;
assign 1_n10693 = ~(1_n11798 | 1_n551);
assign 1_n11013 = ~(1_n1531 ^ 1_n2001);
assign 1_n1582 = 1_n9490 | 1_n9618;
assign 1_n10390 = 1_n12095 & 1_n6464;
assign 1_n10016 = ~1_n10642;
assign 1_n5683 = ~1_n6085;
assign 1_n1216 = ~1_n4957;
assign 1_n5034 = 1_n9762 & 1_n3038;
assign 1_n12590 = 1_n8414 | 1_n4124;
assign 1_n11854 = 1_n7715 & 1_n9669;
assign 1_n5382 = ~1_n7419;
assign 1_n4338 = ~(1_n12559 ^ 1_n6026);
assign 1_n8161 = ~1_n1356;
assign 1_n10784 = ~(1_n7025 | 1_n6994);
assign 1_n13012 = ~1_n5715;
assign 1_n4199 = 1_n715 | 1_n4936;
assign 1_n8442 = ~(1_n6754 ^ 1_n4009);
assign 1_n10789 = ~(1_n122 ^ 1_n10303);
assign 1_n4464 = ~1_n4330;
assign 1_n488 = ~1_n6085;
assign 1_n7054 = 1_n11600 & 1_n2610;
assign 1_n9902 = ~(1_n12541 ^ 1_n3680);
assign 1_n6032 = ~(1_n11139 ^ 1_n10393);
assign 1_n10452 = 1_n8461 & 1_n6388;
assign 1_n2847 = ~(1_n8567 ^ 1_n12176);
assign 1_n8911 = 1_n6967 | 1_n11871;
assign 1_n5467 = ~1_n3627;
assign 1_n12872 = ~(1_n2888 ^ 1_n11066);
assign 1_n11788 = ~(1_n10807 ^ 1_n12656);
assign 1_n11447 = ~(1_n6669 ^ 1_n11872);
assign 1_n9896 = ~(1_n11270 ^ 1_n6899);
assign 1_n72 = 1_n7949 & 1_n3215;
assign 1_n7526 = ~1_n7728;
assign 1_n4163 = ~(1_n9306 ^ 1_n6430);
assign 1_n12653 = ~(1_n6930 | 1_n377);
assign 1_n6342 = ~(1_n1753 | 1_n1915);
assign 1_n749 = 1_n8500 & 1_n3860;
assign 1_n9192 = 1_n7681 & 1_n9066;
assign 1_n9218 = ~(1_n1173 ^ 1_n8347);
assign 1_n10058 = ~(1_n4308 ^ 1_n3820);
assign 1_n3721 = 1_n2048 | 1_n121;
assign 1_n8067 = ~(1_n5096 ^ 1_n9536);
assign 1_n9938 = 1_n10730 | 1_n5076;
assign 1_n4241 = 1_n392 | 1_n6041;
assign 1_n9729 = 1_n8131 | 1_n4640;
assign 1_n975 = ~(1_n13069 ^ 1_n1130);
assign 1_n9498 = ~(1_n2102 | 1_n4838);
assign 1_n11052 = 1_n4588 & 1_n1914;
assign 1_n8035 = ~(1_n4316 ^ 1_n3573);
assign 1_n11182 = ~(1_n2949 ^ 1_n10789);
assign 1_n3811 = ~(1_n3664 | 1_n6408);
assign 1_n8887 = 1_n813 | 1_n10871;
assign 1_n10139 = ~(1_n8998 ^ 1_n4076);
assign 1_n10313 = 1_n10439 | 1_n1026;
assign 1_n2065 = ~(1_n11730 | 1_n6443);
assign 1_n5565 = ~1_n2252;
assign 1_n10268 = 1_n7529 & 1_n2252;
assign 1_n3543 = 1_n6630 | 1_n4230;
assign 1_n6885 = ~(1_n10925 | 1_n4256);
assign 1_n13213 = 1_n563 & 1_n9677;
assign 1_n1828 = 1_n9421 | 1_n8490;
assign 1_n7989 = ~(1_n2087 | 1_n10557);
assign 1_n4751 = 1_n5934 & 1_n4461;
assign 1_n1142 = ~(1_n7231 ^ 1_n12519);
assign 1_n3153 = ~(1_n5139 ^ 1_n5518);
assign 1_n5028 = ~(1_n8626 | 1_n2841);
assign 1_n2072 = 1_n912 ^ 1_n3831;
assign 1_n11724 = ~(1_n1172 ^ 1_n6681);
assign 1_n1077 = 1_n12069 | 1_n9761;
assign 1_n10925 = ~(1_n12539 ^ 1_n10702);
assign 1_n9711 = ~1_n9528;
assign 1_n5869 = 1_n3586 | 1_n1771;
assign 1_n11647 = 1_n1012 | 1_n956;
assign 1_n923 = ~(1_n2013 ^ 1_n205);
assign 1_n11903 = ~(1_n12134 ^ 1_n7574);
assign 1_n10991 = ~1_n772;
assign 1_n9921 = ~1_n7572;
assign 1_n7782 = ~(1_n11499 ^ 1_n6784);
assign 1_n2187 = ~(1_n8717 | 1_n3869);
assign 1_n6411 = ~(1_n7483 ^ 1_n4332);
assign 1_n3367 = 1_n2226 | 1_n9622;
assign 1_n2273 = 1_n3311 & 1_n411;
assign 1_n2130 = ~1_n12567;
assign 1_n1238 = ~1_n5768;
assign 1_n5049 = ~(1_n9842 ^ 1_n12803);
assign 1_n8527 = ~(1_n11015 ^ 1_n2121);
assign 1_n1698 = 1_n2482 & 1_n2758;
assign 1_n2671 = ~1_n3130;
assign 1_n7654 = ~(1_n901 ^ 1_n4775);
assign 1_n9481 = 1_n2777 & 1_n8860;
assign 1_n726 = 1_n12475 ^ 1_n5488;
assign 1_n6866 = 1_n10733 | 1_n10331;
assign 1_n7085 = 1_n11553 ^ 1_n11641;
assign 1_n1215 = ~1_n6445;
assign 1_n3837 = 1_n1579 & 1_n11307;
assign 1_n5851 = 1_n3784 | 1_n9075;
assign 1_n11045 = ~1_n600;
assign 1_n4953 = ~(1_n10660 ^ 1_n7351);
assign 1_n9094 = 1_n7620 | 1_n1985;
assign 1_n1968 = 1_n5733 | 1_n5242;
assign 1_n8589 = ~(1_n11541 ^ 1_n3742);
assign 1_n1114 = ~(1_n13119 ^ 1_n5499);
assign 1_n8548 = 1_n4610 | 1_n5169;
assign 1_n6361 = ~(1_n12857 ^ 1_n7804);
assign 1_n8335 = ~1_n5969;
assign 1_n6507 = 1_n490 & 1_n6389;
assign 1_n6382 = 1_n11284 | 1_n12273;
assign 1_n11510 = ~(1_n7359 ^ 1_n3199);
assign 1_n4800 = ~(1_n5120 ^ 1_n8821);
assign 1_n3790 = ~(1_n10897 ^ 1_n4996);
assign 1_n13125 = 1_n3284 & 1_n6813;
assign 1_n3021 = ~(1_n385 ^ 1_n3523);
assign 1_n10768 = 1_n4001 | 1_n12177;
assign 1_n9929 = 1_n4818 & 1_n1602;
assign 1_n12992 = 1_n10638 | 1_n8983;
assign 1_n10349 = ~(1_n10578 | 1_n5282);
assign 1_n2163 = ~1_n11179;
assign 1_n8179 = 1_n870 & 1_n11655;
assign 1_n3868 = ~(1_n7382 ^ 1_n10461);
assign 1_n359 = ~(1_n8967 ^ 1_n12163);
assign 1_n1259 = 1_n3090 | 1_n990;
assign 1_n2351 = 1_n1715 & 1_n8313;
assign 1_n6165 = ~(1_n4645 ^ 1_n2447);
assign 1_n5629 = ~(1_n8158 ^ 1_n12360);
assign 1_n869 = 1_n5902 | 1_n11606;
assign 1_n9592 = ~1_n7085;
assign 1_n9233 = 1_n10289 & 1_n4755;
assign 1_n8690 = ~(1_n13121 ^ 1_n11348);
assign 1_n987 = ~1_n12065;
assign 1_n11229 = 1_n11751 | 1_n1820;
assign 1_n1499 = 1_n10962 | 1_n10473;
assign 1_n513 = ~1_n229;
assign 1_n4727 = 1_n1101 | 1_n10871;
assign 1_n8612 = ~(1_n690 ^ 1_n6893);
assign 1_n4952 = ~(1_n5071 | 1_n10861);
assign 1_n2718 = ~1_n9620;
assign 1_n7971 = 1_n9515 | 1_n2569;
assign 1_n10654 = ~1_n3095;
assign 1_n3157 = ~1_n103;
assign 1_n5673 = ~1_n7153;
assign 1_n4824 = 1_n5965 ^ 1_n485;
assign 1_n570 = 1_n7925 | 1_n8563;
assign 1_n1395 = 1_n10479 & 1_n11434;
assign 1_n7815 = ~(1_n9989 ^ 1_n12692);
assign 1_n2450 = ~(1_n9235 | 1_n9506);
assign 1_n4713 = ~(1_n9150 ^ 1_n2397);
assign 1_n9482 = 1_n11845 | 1_n4658;
assign 1_n13193 = ~(1_n11361 ^ 1_n13016);
assign 1_n12765 = 1_n10085 | 1_n1570;
assign 1_n10595 = 1_n8717 & 1_n3869;
assign 1_n2893 = ~1_n8230;
assign 1_n6789 = 1_n6066 & 1_n3706;
assign 1_n1385 = ~(1_n10446 ^ 1_n10939);
assign 1_n3145 = 1_n7443 & 1_n12442;
assign 1_n9028 = ~(1_n10046 ^ 1_n5259);
assign 1_n2079 = 1_n7872 | 1_n8744;
assign 1_n4737 = 1_n3348 | 1_n11748;
assign 1_n1995 = ~(1_n2440 | 1_n13163);
assign 1_n3842 = 1_n3733 | 1_n11426;
assign 1_n8005 = ~1_n2590;
assign 1_n7166 = ~(1_n9861 ^ 1_n1207);
assign 1_n5846 = 1_n1168 | 1_n8348;
assign 1_n7276 = 1_n1757 & 1_n4330;
assign 1_n11211 = ~(1_n2261 ^ 1_n7061);
assign 1_n7901 = 1_n1633 | 1_n5524;
assign 1_n10911 = ~(1_n12754 ^ 1_n7451);
assign 1_n10454 = ~(1_n705 | 1_n9208);
assign 1_n11072 = ~(1_n2730 ^ 1_n11440);
assign 1_n12471 = ~1_n767;
assign 1_n9679 = ~1_n5320;
assign 1_n10411 = ~1_n1982;
assign 1_n6164 = ~1_n8917;
assign 1_n1346 = ~1_n6836;
assign 1_n2795 = 1_n6054 | 1_n5290;
assign 1_n12185 = 1_n8670 | 1_n2707;
assign 1_n388 = ~(1_n6195 ^ 1_n12886);
assign 1_n11270 = ~1_n691;
assign 1_n11569 = 1_n8642 & 1_n8488;
assign 1_n7664 = ~(1_n7671 ^ 1_n8078);
assign 1_n9916 = ~(1_n8718 | 1_n11531);
assign 1_n10846 = ~(1_n7593 ^ 1_n10701);
assign 1_n8543 = 1_n104 & 1_n6911;
assign 1_n11833 = ~(1_n7500 | 1_n3681);
assign 1_n9150 = 1_n4166 | 1_n6404;
assign 1_n9225 = 1_n12361 & 1_n10317;
assign 1_n2923 = ~(1_n12217 ^ 1_n7164);
assign 1_n6850 = 1_n4966 | 1_n9714;
assign 1_n10987 = ~(1_n4750 ^ 1_n11475);
assign 1_n9267 = ~(1_n3309 ^ 1_n11534);
assign 1_n4440 = 1_n11665 & 1_n8860;
assign 1_n4669 = 1_n8736 & 1_n7081;
assign 1_n8852 = ~1_n5214;
assign 1_n2293 = ~(1_n6722 ^ 1_n7416);
assign 1_n8909 = 1_n9634 | 1_n12029;
assign 1_n10816 = ~(1_n10331 ^ 1_n13226);
assign 1_n7068 = ~1_n9528;
assign 1_n2089 = 1_n5268 & 1_n7012;
assign 1_n9275 = ~(1_n7715 | 1_n2458);
assign 1_n1710 = 1_n5442 & 1_n181;
assign 1_n10785 = ~(1_n10804 ^ 1_n1573);
assign 1_n3288 = 1_n11320 | 1_n10871;
assign 1_n1920 = ~1_n6064;
assign 1_n2781 = 1_n12565 | 1_n5067;
assign 1_n13029 = ~(1_n6780 ^ 1_n2111);
assign 1_n11602 = ~(1_n2058 | 1_n6907);
assign 1_n4059 = ~(1_n2731 ^ 1_n5880);
assign 1_n3191 = 1_n2449 | 1_n1570;
assign 1_n4461 = 1_n4348 | 1_n7813;
assign 1_n8009 = 1_n3025 | 1_n4510;
assign 1_n4733 = 1_n5129 & 1_n9180;
assign 1_n9206 = ~(1_n7118 ^ 1_n12480);
assign 1_n6861 = 1_n10544 ^ 1_n1064;
assign 1_n12667 = ~1_n6950;
assign 1_n4832 = ~(1_n2821 ^ 1_n5343);
assign 1_n7980 = ~1_n6277;
assign 1_n1877 = ~(1_n4205 | 1_n1351);
assign 1_n6871 = 1_n12522 | 1_n5775;
assign 1_n3981 = 1_n789;
assign 1_n2824 = ~1_n5833;
assign 1_n9451 = 1_n2384 | 1_n3396;
assign 1_n11085 = 1_n7797 & 1_n5996;
assign 1_n3818 = 1_n6086 | 1_n12188;
assign 1_n800 = ~(1_n8587 ^ 1_n4707);
assign 1_n2768 = ~1_n4335;
assign 1_n4739 = 1_n5784 ^ 1_n7722;
assign 1_n8137 = ~(1_n2361 ^ 1_n11897);
assign 1_n4890 = ~1_n3832;
assign 1_n12949 = 1_n2583 & 1_n10673;
assign 1_n1762 = 1_n2472 & 1_n11593;
assign 1_n7960 = 1_n11665 & 1_n9570;
assign 1_n7932 = ~(1_n3739 ^ 1_n325);
assign 1_n8778 = ~1_n3988;
assign 1_n9736 = ~1_n11474;
assign 1_n10469 = 1_n4855 | 1_n2958;
assign 1_n11355 = ~(1_n52 ^ 1_n11923);
assign 1_n2014 = ~(1_n8411 ^ 1_n807);
assign 1_n6981 = 1_n7177 | 1_n10551;
assign 1_n4587 = 1_n6884 & 1_n6424;
assign 1_n6737 = ~(1_n10047 | 1_n12591);
assign 1_n4724 = 1_n3858;
assign 1_n2678 = ~1_n11734;
assign 1_n8239 = 1_n2576 | 1_n8262;
assign 1_n12833 = 1_n13190 | 1_n6265;
assign 1_n1480 = ~1_n11734;
assign 1_n10711 = ~1_n3715;
assign 1_n10771 = 1_n2896 | 1_n10311;
assign 1_n9361 = 1_n7878 | 1_n10552;
assign 1_n10650 = 1_n4649 | 1_n2059;
assign 1_n12716 = 1_n11965 | 1_n10764;
assign 1_n10624 = 1_n5645 | 1_n6732;
assign 1_n11867 = 1_n12648 | 1_n8561;
assign 1_n12231 = 1_n417 & 1_n7109;
assign 1_n13099 = 1_n881 | 1_n2176;
assign 1_n11083 = ~(1_n11572 ^ 1_n1584);
assign 1_n4322 = 1_n12020 | 1_n3210;
assign 1_n10658 = 1_n12010 & 1_n11451;
assign 1_n12315 = ~1_n2374;
assign 1_n12187 = ~(1_n3862 ^ 1_n571);
assign 1_n6434 = ~(1_n824 ^ 1_n1318);
assign 1_n13144 = ~(1_n5874 ^ 1_n10468);
assign 1_n4752 = ~(1_n3615 | 1_n5507);
assign 1_n4721 = ~(1_n9645 ^ 1_n10056);
assign 1_n4778 = ~1_n382;
assign 1_n7924 = ~(1_n4217 ^ 1_n3029);
assign 1_n10561 = 1_n1360 | 1_n9511;
assign 1_n11340 = ~1_n11199;
assign 1_n2396 = 1_n9593 | 1_n8806;
assign 1_n1554 = ~1_n937;
assign 1_n5222 = ~1_n299;
assign 1_n11105 = 1_n9341 | 1_n2594;
assign 1_n6572 = ~(1_n3802 ^ 1_n2459);
assign 1_n12431 = 1_n9339 | 1_n9159;
assign 1_n710 = ~(1_n4576 ^ 1_n9773);
assign 1_n8323 = ~(1_n8426 ^ 1_n11754);
assign 1_n8515 = ~(1_n9534 ^ 1_n3268);
assign 1_n10459 = ~1_n9901;
assign 1_n8107 = 1_n13205 | 1_n4310;
assign 1_n3967 = 1_n7470 & 1_n3020;
assign 1_n4290 = ~1_n9531;
assign 1_n2548 = ~(1_n6067 ^ 1_n1076);
assign 1_n8756 = ~(1_n3305 | 1_n5662);
assign 1_n845 = ~1_n7729;
assign 1_n723 = 1_n3429 | 1_n4030;
assign 1_n7785 = 1_n3936 & 1_n4810;
assign 1_n2382 = ~(1_n9535 ^ 1_n2852);
assign 1_n5796 = ~(1_n9107 ^ 1_n4520);
assign 1_n11408 = 1_n10593 | 1_n3063;
assign 1_n12561 = ~(1_n5309 | 1_n1000);
assign 1_n1228 = ~(1_n2128 ^ 1_n8403);
assign 1_n2832 = ~1_n12422;
assign 1_n6039 = 1_n9252 | 1_n3464;
assign 1_n8027 = ~(1_n10913 ^ 1_n3746);
assign 1_n1789 = ~1_n3253;
assign 1_n8314 = 1_n53 | 1_n6769;
assign 1_n2825 = ~1_n5189;
assign 1_n11919 = 1_n6043 | 1_n327;
assign 1_n9951 = ~(1_n10514 ^ 1_n7293);
assign 1_n11413 = ~(1_n1991 ^ 1_n8603);
assign 1_n7362 = ~1_n13128;
assign 1_n12543 = 1_n12992 & 1_n9409;
assign 1_n9539 = 1_n4665 | 1_n1985;
assign 1_n5695 = 1_n1511 | 1_n11668;
assign 1_n10879 = ~1_n5031;
assign 1_n10092 = 1_n7258 | 1_n12234;
assign 1_n5617 = ~(1_n9874 ^ 1_n6397);
assign 1_n5491 = 1_n10354 | 1_n12763;
assign 1_n8584 = ~(1_n487 ^ 1_n9239);
assign 1_n6218 = 1_n11318 | 1_n8880;
assign 1_n9752 = 1_n3583 & 1_n13010;
assign 1_n2348 = 1_n300 | 1_n10619;
assign 1_n4744 = ~1_n1595;
assign 1_n5036 = 1_n10346 & 1_n2534;
assign 1_n11362 = 1_n11415 & 1_n7564;
assign 1_n5966 = 1_n7984 | 1_n11470;
assign 1_n2067 = ~1_n7137;
assign 1_n4802 = ~(1_n11142 ^ 1_n11762);
assign 1_n7419 = 1_n10188 | 1_n4947;
assign 1_n7887 = 1_n5667 | 1_n11144;
assign 1_n5676 = 1_n3022 & 1_n12807;
assign 1_n12344 = 1_n12224 | 1_n4979;
assign 1_n12011 = ~(1_n12081 ^ 1_n9936);
assign 1_n11633 = 1_n1265 | 1_n2552;
assign 1_n2673 = ~1_n1552;
assign 1_n9877 = 1_n5079 | 1_n1144;
assign 1_n9661 = 1_n898 & 1_n4154;
assign 1_n11649 = ~(1_n244 | 1_n2436);
assign 1_n9313 = 1_n4796 | 1_n4947;
assign 1_n7751 = 1_n2118 | 1_n12273;
assign 1_n12735 = ~(1_n4508 | 1_n7686);
assign 1_n10339 = 1_n11339 & 1_n1080;
assign 1_n9198 = ~(1_n12061 ^ 1_n753);
assign 1_n12375 = 1_n8934 | 1_n4423;
assign 1_n1351 = 1_n3898 | 1_n9223;
assign 1_n10690 = ~(1_n3254 | 1_n3979);
assign 1_n1292 = 1_n581 & 1_n8957;
assign 1_n11742 = 1_n12242 | 1_n5087;
assign 1_n5285 = ~(1_n3138 | 1_n11316);
assign 1_n3643 = 1_n2451 & 1_n2799;
assign 1_n11771 = ~1_n13219;
assign 1_n12928 = ~(1_n10197 ^ 1_n10615);
assign 1_n9520 = 1_n278 | 1_n11968;
assign 1_n11987 = 1_n12748 | 1_n10871;
assign 1_n6287 = ~(1_n11229 ^ 1_n7758);
assign 1_n13221 = 1_n10761 | 1_n13242;
assign 1_n9269 = ~(1_n9683 | 1_n5849);
assign 1_n2034 = 1_n97 | 1_n4373;
assign 1_n12831 = ~(1_n11653 ^ 1_n13042);
assign 1_n5379 = 1_n12129 & 1_n10960;
assign 1_n6494 = ~(1_n3518 | 1_n1069);
assign 1_n3860 = 1_n11986 & 1_n10376;
assign 1_n4567 = ~(1_n4568 | 1_n3353);
assign 1_n4837 = ~(1_n6861 ^ 1_n1802);
assign 1_n6269 = 1_n2590 & 1_n8290;
assign 1_n9827 = ~1_n6317;
assign 1_n11898 = 1_n11994 & 1_n331;
assign 1_n1532 = ~(1_n12584 ^ 1_n3045);
assign 1_n4409 = ~(1_n7788 ^ 1_n8007);
assign 1_n6426 = 1_n11819 & 1_n8775;
assign 1_n6775 = 1_n6710 | 1_n5782;
assign 1_n11402 = 1_n5568 & 1_n4748;
assign 1_n10426 = 1_n4235 | 1_n3576;
assign 1_n5177 = ~1_n12557;
assign 1_n10891 = 1_n9011 | 1_n3559;
assign 1_n841 = ~(1_n12796 ^ 1_n8308);
assign 1_n8523 = 1_n3944 & 1_n3541;
assign 1_n10402 = ~1_n1636;
assign 1_n4772 = ~(1_n7849 ^ 1_n5543);
assign 1_n7558 = ~(1_n8830 ^ 1_n10181);
assign 1_n171 = ~(1_n7806 ^ 1_n11377);
assign 1_n9317 = ~(1_n5744 ^ 1_n7715);
assign 1_n12172 = 1_n13006 ^ 1_n10268;
assign 1_n6569 = ~(1_n250 | 1_n2492);
assign 1_n7233 = ~(1_n9543 | 1_n2489);
assign 1_n5544 = ~(1_n4559 ^ 1_n5675);
assign 1_n6817 = ~(1_n4573 | 1_n10838);
assign 1_n714 = 1_n8324 | 1_n2675;
assign 1_n4471 = 1_n2405 | 1_n8614;
assign 1_n4459 = ~(1_n5197 ^ 1_n6600);
assign 1_n5030 = ~(1_n8657 ^ 1_n9127);
assign 1_n10166 = ~(1_n7560 | 1_n6600);
assign 1_n6239 = 1_n1607 & 1_n9780;
assign 1_n12345 = ~(1_n4768 ^ 1_n3943);
assign 1_n11660 = 1_n6183 | 1_n3977;
assign 1_n8804 = ~(1_n3501 ^ 1_n7607);
assign 1_n9214 = ~(1_n536 ^ 1_n4581);
assign 1_n6438 = ~1_n1165;
assign 1_n5381 = 1_n6314 | 1_n2354;
assign 1_n1125 = 1_n10558 | 1_n4724;
assign 1_n9117 = 1_n4211 ^ 1_n10485;
assign 1_n5151 = 1_n1101 | 1_n2387;
assign 1_n11449 = ~1_n6392;
assign 1_n10652 = 1_n1460 & 1_n5506;
assign 1_n12328 = 1_n9280;
assign 1_n2368 = ~(1_n11035 ^ 1_n1439);
assign 1_n9920 = 1_n100 & 1_n9725;
assign 1_n3417 = 1_n10128 | 1_n11107;
assign 1_n11407 = 1_n935 | 1_n4230;
assign 1_n6314 = ~1_n7527;
assign 1_n8995 = ~1_n4788;
assign 1_n11707 = ~1_n2409;
assign 1_n9505 = ~(1_n12769 ^ 1_n2909);
assign 1_n8474 = 1_n8912 | 1_n2622;
assign 1_n10623 = 1_n12915 & 1_n4487;
assign 1_n4231 = 1_n1024 & 1_n4294;
assign 1_n6854 = ~1_n12482;
assign 1_n5787 = ~1_n7240;
assign 1_n12745 = ~(1_n6816 ^ 1_n7332);
assign 1_n10669 = ~(1_n8317 ^ 1_n12212);
assign 1_n10861 = ~(1_n6353 ^ 1_n7431);
assign 1_n4351 = ~(1_n2830 ^ 1_n10833);
assign 1_n10086 = ~(1_n7416 | 1_n6722);
assign 1_n2472 = ~1_n3390;
assign 1_n1098 = 1_n9489 | 1_n2059;
assign 1_n6725 = 1_n2662 | 1_n6863;
assign 1_n8582 = ~(1_n696 ^ 1_n9000);
assign 1_n9999 = ~(1_n10024 ^ 1_n1967);
assign 1_n6812 = ~(1_n7345 ^ 1_n8895);
assign 1_n3353 = 1_n9460 & 1_n12452;
assign 1_n1132 = 1_n715 | 1_n11668;
assign 1_n10286 = ~1_n9620;
assign 1_n3949 = 1_n6274;
assign 1_n11467 = ~(1_n9843 ^ 1_n6528);
assign 1_n7347 = ~(1_n6720 ^ 1_n2584);
assign 1_n4507 = ~(1_n4538 ^ 1_n8667);
assign 1_n11473 = 1_n8350 & 1_n6000;
assign 1_n660 = ~(1_n4630 | 1_n5312);
assign 1_n428 = ~1_n10599;
assign 1_n6169 = ~(1_n9926 ^ 1_n5175);
assign 1_n6949 = 1_n7476 & 1_n2301;
assign 1_n2811 = 1_n9478 | 1_n1144;
assign 1_n1714 = ~(1_n9975 ^ 1_n7482);
assign 1_n4693 = ~(1_n3885 | 1_n6499);
assign 1_n10468 = ~(1_n9122 ^ 1_n7674);
assign 1_n12416 = ~1_n2252;
assign 1_n4069 = ~(1_n12598 ^ 1_n4437);
assign 1_n11711 = ~(1_n4081 | 1_n9186);
assign 1_n5360 = ~1_n12381;
assign 1_n11579 = ~(1_n4065 ^ 1_n3226);
assign 1_n6587 = ~1_n10805;
assign 1_n5830 = 1_n13202 | 1_n7016;
assign 1_n11263 = 1_n6133 | 1_n4373;
assign 1_n10883 = ~1_n5920;
assign 1_n9191 = 1_n11121 | 1_n6899;
assign 1_n8771 = ~(1_n4992 | 1_n2399);
assign 1_n322 = 1_n2546 ^ 1_n7477;
assign 1_n13104 = ~(1_n2700 ^ 1_n3575);
assign 1_n7497 = 1_n6670 & 1_n7346;
assign 1_n2656 = ~(1_n1954 ^ 1_n1488);
assign 1_n9107 = 1_n5008 | 1_n4110;
assign 1_n4871 = 1_n9383 | 1_n5242;
assign 1_n4213 = 1_n6014 & 1_n6359;
assign 1_n5312 = ~1_n376;
assign 1_n3441 = 1_n9711 | 1_n8030;
assign 1_n2322 = 1_n7503 | 1_n11184;
assign 1_n11332 = ~(1_n8070 ^ 1_n8735);
assign 1_n9873 = 1_n248 & 1_n8769;
assign 1_n9962 = ~1_n5729;
assign 1_n1809 = 1_n12229 & 1_n4941;
assign 1_n10836 = ~(1_n8130 ^ 1_n3190);
assign 1_n330 = ~(1_n8866 | 1_n8620);
assign 1_n4676 = ~(1_n25 ^ 1_n5901);
assign 1_n6201 = ~(1_n4922 ^ 1_n365);
assign 1_n12903 = ~(1_n12558 ^ 1_n12426);
assign 1_n9940 = 1_n8104 | 1_n7528;
assign 1_n9320 = 1_n4519 | 1_n7080;
assign 1_n8340 = 1_n11504 & 1_n10262;
assign 1_n1703 = 1_n8594 & 1_n12804;
assign 1_n7770 = 1_n1951 & 1_n6526;
assign 1_n4691 = 1_n1630 & 1_n5807;
assign 1_n8324 = ~1_n9300;
assign 1_n12749 = ~(1_n12301 ^ 1_n2180);
assign 1_n10372 = ~(1_n7676 | 1_n1209);
assign 1_n7232 = 1_n175 | 1_n9369;
assign 1_n2315 = 1_n10712 & 1_n1864;
assign 1_n11832 = ~(1_n9855 | 1_n7063);
assign 1_n10382 = ~(1_n1841 ^ 1_n10938);
assign 1_n4595 = 1_n4967 | 1_n8563;
assign 1_n4366 = ~1_n8233;
assign 1_n2559 = 1_n7170 | 1_n2631;
assign 1_n8420 = 1_n10225 ^ 1_n10322;
assign 1_n4238 = 1_n7783 | 1_n12388;
assign 1_n9350 = ~1_n1826;
assign 1_n2480 = 1_n9275 | 1_n5744;
assign 1_n2581 = ~1_n10805;
assign 1_n3307 = 1_n4063 | 1_n1218;
assign 1_n10680 = 1_n1563 ^ 1_n2951;
assign 1_n8525 = 1_n423 | 1_n9179;
assign 1_n2691 = ~1_n10190;
assign 1_n6358 = ~1_n12026;
assign 1_n10400 = ~1_n9846;
assign 1_n3804 = ~1_n1992;
assign 1_n8761 = 1_n3726 | 1_n7723;
assign 1_n11253 = 1_n3911 | 1_n9075;
assign 1_n1785 = 1_n7658 | 1_n8512;
assign 1_n11430 = 1_n9648 | 1_n8677;
assign 1_n3414 = 1_n10258 & 1_n7823;
assign 1_n12782 = ~(1_n11773 | 1_n10116);
assign 1_n11257 = ~(1_n3954 ^ 1_n1792);
assign 1_n8431 = 1_n9554 & 1_n4252;
assign 1_n2952 = 1_n10624 | 1_n11708;
assign 1_n3192 = 1_n3877 | 1_n8874;
assign 1_n8740 = 1_n12316 | 1_n1422;
assign 1_n3534 = ~1_n1636;
assign 1_n347 = 1_n8681 | 1_n7723;
assign 1_n12002 = ~(1_n7813 ^ 1_n5742);
assign 1_n1555 = ~(1_n4755 ^ 1_n10289);
assign 1_n10831 = ~(1_n2512 ^ 1_n131);
assign 1_n8856 = 1_n11068 & 1_n9308;
assign 1_n3105 = ~(1_n8380 ^ 1_n7596);
assign 1_n8652 = ~(1_n11295 ^ 1_n1982);
assign 1_n11826 = ~(1_n10983 ^ 1_n12154);
assign 1_n11648 = 1_n5148 | 1_n4230;
assign 1_n9903 = ~(1_n10516 ^ 1_n5686);
assign 1_n8262 = 1_n9169 & 1_n1796;
assign 1_n8517 = ~(1_n5902 ^ 1_n6092);
assign 1_n3975 = 1_n10650 | 1_n921;
assign 1_n920 = 1_n12254 | 1_n1043;
assign 1_n12129 = 1_n6828 | 1_n11796;
assign 1_n12244 = 1_n12150 & 1_n4145;
assign 1_n1965 = ~1_n4557;
assign 1_n4346 = 1_n1073 & 1_n6983;
assign 1_n6560 = ~(1_n12470 | 1_n7656);
assign 1_n180 = ~(1_n5329 ^ 1_n5701);
assign 1_n12850 = 1_n3804 & 1_n12941;
assign 1_n11490 = 1_n1202 ^ 1_n10808;
assign 1_n2451 = ~(1_n4719 ^ 1_n11412);
assign 1_n7938 = 1_n10977 | 1_n8348;
assign 1_n5391 = ~(1_n11907 ^ 1_n12327);
assign 1_n11320 = ~1_n4330;
assign 1_n21 = 1_n2255 | 1_n9314;
assign 1_n7603 = ~(1_n8331 ^ 1_n1046);
assign 1_n1904 = 1_n755 | 1_n3598;
assign 1_n6900 = 1_n12630 | 1_n1240;
assign 1_n8906 = 1_n10423 | 1_n264;
assign 1_n10724 = 1_n10854 | 1_n837;
assign 1_n12632 = 1_n6633 ^ 1_n11607;
assign 1_n8361 = 1_n6630 | 1_n4373;
assign 1_n5043 = ~(1_n6212 | 1_n11219);
assign 1_n314 = ~(1_n12688 | 1_n4270);
assign 1_n2505 = ~(1_n12840 ^ 1_n4611);
assign 1_n7973 = 1_n305 | 1_n5724;
assign 1_n37 = 1_n7358 | 1_n1571;
assign 1_n3254 = ~(1_n2284 | 1_n8770);
assign 1_n805 = ~(1_n1716 | 1_n11438);
assign 1_n10231 = 1_n11910 | 1_n2449;
assign 1_n8868 = ~1_n13058;
assign 1_n66 = 1_n2595 ^ 1_n8760;
assign 1_n58 = ~(1_n8766 ^ 1_n6874);
assign 1_n11868 = ~1_n10451;
assign 1_n10133 = ~(1_n2932 | 1_n11182);
assign 1_n12996 = ~(1_n2417 ^ 1_n4319);
assign 1_n12108 = ~(1_n2522 | 1_n9998);
assign 1_n8954 = 1_n6099 | 1_n1043;
assign 1_n9355 = 1_n11121 | 1_n5802;
assign 1_n11731 = ~(1_n5851 ^ 1_n7413);
assign 1_n1154 = 1_n8307 & 1_n4940;
assign 1_n5510 = 1_n8447 & 1_n12292;
assign 1_n12790 = 1_n3676 | 1_n3640;
assign 1_n11773 = 1_n10266 | 1_n9745;
assign 1_n12537 = ~1_n4964;
assign 1_n3572 = ~1_n1982;
assign 1_n5499 = 1_n6486 | 1_n12501;
assign 1_n13002 = ~(1_n11190 ^ 1_n10740);
assign 1_n11863 = ~(1_n740 ^ 1_n11738);
assign 1_n2693 = ~(1_n12452 ^ 1_n9115);
assign 1_n7593 = ~(1_n9124 ^ 1_n7229);
assign 1_n10868 = ~(1_n2710 ^ 1_n541);
assign 1_n6875 = ~1_n9591;
assign 1_n8168 = 1_n8876 | 1_n12487;
assign 1_n8701 = ~(1_n2280 ^ 1_n2185);
assign 1_n4140 = ~(1_n7999 ^ 1_n8171);
assign 1_n690 = 1_n10611 & 1_n11307;
assign 1_n2312 = ~(1_n6172 ^ 1_n5756);
assign 1_n11259 = 1_n1062 & 1_n12310;
assign 1_n11639 = 1_n6329 & 1_n4883;
assign 1_n3844 = ~(1_n8235 ^ 1_n3100);
assign 1_n11160 = ~(1_n5123 ^ 1_n2029);
assign 1_n756 = ~(1_n4759 ^ 1_n5116);
assign 1_n5481 = ~(1_n2651 ^ 1_n10933);
assign 1_n312 = ~1_n12112;
assign 1_n12367 = 1_n8838 ^ 1_n3494;
assign 1_n13161 = ~(1_n7979 ^ 1_n3392);
assign 1_n2978 = 1_n2874 & 1_n12815;
assign 1_n3126 = ~1_n12965;
assign 1_n3014 = ~(1_n13014 ^ 1_n12751);
assign 1_n11203 = 1_n10143 | 1_n4373;
assign 1_n8432 = 1_n9171 | 1_n6257;
assign 1_n10574 = ~1_n394;
assign 1_n12376 = ~(1_n7485 | 1_n4889);
assign 1_n294 = 1_n5157 | 1_n12049;
assign 1_n5052 = ~(1_n6065 ^ 1_n1120);
assign 1_n7010 = 1_n9497 & 1_n6330;
assign 1_n6397 = ~(1_n12879 ^ 1_n2494);
assign 1_n8446 = 1_n2022 | 1_n1193;
assign 1_n8114 = ~(1_n10915 ^ 1_n10226);
assign 1_n9419 = ~(1_n3088 ^ 1_n7121);
assign 1_n8260 = 1_n12738 & 1_n3543;
assign 1_n10529 = 1_n7953 | 1_n11051;
assign 1_n9413 = 1_n3372 & 1_n5544;
assign 1_n1713 = 1_n12465 | 1_n11668;
assign 1_n6878 = ~1_n9293;
assign 1_n9607 = ~1_n5647;
assign 1_n76 = 1_n11104 & 1_n6157;
assign 1_n8614 = 1_n3326 & 1_n387;
assign 1_n2756 = ~(1_n9522 ^ 1_n10635);
assign 1_n8552 = 1_n9930 & 1_n3980;
assign 1_n11371 = ~(1_n686 ^ 1_n2885);
assign 1_n3599 = 1_n2067 | 1_n8096;
assign 1_n4558 = 1_n8977 | 1_n10179;
assign 1_n840 = 1_n1778 | 1_n9572;
assign 1_n4690 = ~(1_n12025 ^ 1_n8314);
assign 1_n5949 = ~1_n6392;
assign 1_n662 = 1_n11225 | 1_n2133;
assign 1_n6931 = ~(1_n3101 ^ 1_n2290);
assign 1_n12096 = ~(1_n6753 ^ 1_n4812);
assign 1_n6455 = 1_n1333 & 1_n8842;
assign 1_n5882 = ~(1_n7379 ^ 1_n9165);
assign 1_n11690 = 1_n5498 | 1_n8800;
assign 1_n12984 = 1_n11404 | 1_n5797;
assign 1_n2859 = ~(1_n10221 ^ 1_n5812);
assign 1_n6656 = ~(1_n9374 | 1_n3389);
assign 1_n6820 = ~(1_n1242 ^ 1_n12173);
assign 1_n9956 = ~(1_n4459 ^ 1_n1662);
assign 1_n6030 = ~(1_n8813 ^ 1_n2470);
assign 1_n10740 = 1_n3006 & 1_n10451;
assign 1_n10641 = ~1_n2737;
assign 1_n3570 = ~1_n11285;
assign 1_n9875 = ~(1_n11334 ^ 1_n9359);
assign 1_n5550 = ~1_n11665;
assign 1_n6067 = 1_n795 | 1_n10135;
assign 1_n2316 = ~(1_n10150 ^ 1_n12054);
assign 1_n6564 = ~(1_n9526 | 1_n10146);
assign 1_n7682 = 1_n11345 & 1_n5250;
assign 1_n3277 = ~(1_n7776 ^ 1_n518);
assign 1_n12878 = 1_n10991 | 1_n8268;
assign 1_n10220 = 1_n12295 | 1_n3981;
assign 1_n1665 = 1_n11370 | 1_n4724;
assign 1_n13177 = 1_n398 | 1_n10813;
assign 1_n3460 = ~1_n9570;
assign 1_n11497 = 1_n10137 | 1_n2133;
assign 1_n7332 = ~(1_n1419 ^ 1_n30);
assign 1_n391 = ~(1_n2072 | 1_n8481);
assign 1_n8044 = ~1_n1762;
assign 1_n858 = ~(1_n6975 ^ 1_n7871);
assign 1_n10159 = ~(1_n4033 ^ 1_n3552);
assign 1_n496 = 1_n9328 & 1_n5948;
assign 1_n9185 = ~(1_n10844 ^ 1_n5042);
assign 1_n2358 = 1_n12648 | 1_n9962;
assign 1_n3408 = 1_n3259 | 1_n6732;
assign 1_n1358 = ~1_n976;
assign 1_n6636 = 1_n10039 & 1_n11110;
assign 1_n11763 = ~(1_n1299 ^ 1_n5397);
assign 1_n7988 = 1_n4085 & 1_n10348;
assign 1_n11953 = ~(1_n6821 ^ 1_n1369);
assign 1_n5774 = 1_n69 | 1_n12273;
assign 1_n7462 = ~(1_n2466 ^ 1_n11068);
assign 1_n12570 = ~(1_n5419 ^ 1_n10069);
assign 1_n9088 = 1_n12630 & 1_n1240;
assign 1_n3600 = 1_n11818 & 1_n10022;
assign 1_n12207 = ~(1_n4284 ^ 1_n9166);
assign 1_n1061 = ~(1_n7193 ^ 1_n9933);
assign 1_n3776 = ~(1_n242 | 1_n6941);
assign 1_n11783 = ~1_n10025;
assign 1_n2357 = 1_n9129 | 1_n1026;
assign 1_n12567 = 1_n12370 & 1_n12824;
assign 1_n13163 = ~(1_n3907 ^ 1_n7513);
assign 1_n4534 = 1_n7114 & 1_n4192;
assign 1_n12146 = ~(1_n9049 ^ 1_n1577);
assign 1_n8208 = 1_n7997 | 1_n4959;
assign 1_n11803 = 1_n3836 | 1_n1103;
assign 1_n10328 = 1_n5372 & 1_n4481;
assign 1_n1848 = ~(1_n7952 | 1_n9571);
assign 1_n13206 = ~(1_n8389 | 1_n7192);
assign 1_n11692 = 1_n1571 | 1_n8490;
assign 1_n7435 = ~(1_n6148 ^ 1_n6458);
assign 1_n11642 = 1_n10499 | 1_n11843;
assign 1_n3368 = ~(1_n10477 ^ 1_n10484);
assign 1_n6396 = ~(1_n9928 ^ 1_n12314);
assign 1_n8094 = 1_n7765 & 1_n10906;
assign 1_n10242 = ~(1_n7156 | 1_n1932);
assign 1_n11281 = 1_n1489 & 1_n10806;
assign 1_n2334 = 1_n7544 & 1_n198;
assign 1_n7053 = ~(1_n3543 ^ 1_n9367);
assign 1_n11988 = 1_n9216 & 1_n9475;
assign 1_n4967 = ~1_n6085;
assign 1_n11956 = 1_n3249 | 1_n3161;
assign 1_n12017 = 1_n7475 & 1_n8982;
assign 1_n8788 = 1_n6367 | 1_n10319;
assign 1_n1108 = ~(1_n7885 | 1_n1187);
assign 1_n8947 = ~(1_n8567 | 1_n6718);
assign 1_n8691 = ~(1_n7136 ^ 1_n10698);
assign 1_n12947 = ~(1_n7375 ^ 1_n12618);
assign 1_n6743 = ~1_n22;
assign 1_n6990 = ~1_n5475;
assign 1_n13160 = ~(1_n5316 ^ 1_n8320);
assign 1_n10527 = ~1_n10122;
assign 1_n12153 = ~1_n11411;
assign 1_n10589 = 1_n7669 & 1_n9101;
assign 1_n1119 = ~(1_n8299 ^ 1_n11752);
assign 1_n1052 = ~1_n6826;
assign 1_n6504 = ~1_n498;
assign 1_n7418 = 1_n8615 | 1_n8268;
assign 1_n12151 = ~(1_n1977 ^ 1_n849);
assign 1_n9339 = ~1_n11891;
assign 1_n4860 = ~(1_n3148 ^ 1_n4902);
assign 1_n4722 = ~1_n3677;
assign 1_n2071 = 1_n5811 & 1_n8202;
assign 1_n913 = ~1_n6561;
assign 1_n6566 = 1_n11868 | 1_n5076;
assign 1_n7928 = ~(1_n4480 ^ 1_n10598);
assign 1_n3442 = 1_n567 | 1_n11833;
assign 1_n437 = ~(1_n720 ^ 1_n5600);
assign 1_n12217 = ~(1_n1456 ^ 1_n9333);
assign 1_n3214 = 1_n1367 | 1_n5971;
assign 1_n13039 = ~1_n3769;
assign 1_n8493 = 1_n8034 & 1_n9496;
assign 1_n2308 = 1_n2607 & 1_n6640;
assign 1_n8016 = 1_n9418 & 1_n1214;
assign 1_n4922 = ~(1_n3872 | 1_n9301);
assign 1_n12876 = 1_n4441 & 1_n2600;
assign 1_n4033 = 1_n8046 & 1_n1410;
assign 1_n12967 = ~1_n4470;
assign 1_n801 = ~(1_n10965 ^ 1_n2826);
assign 1_n5657 = ~(1_n6494 ^ 1_n4438);
assign 1_n5587 = ~(1_n2774 ^ 1_n4415);
assign 1_n5051 = ~(1_n11039 ^ 1_n11873);
assign 1_n1105 = ~1_n587;
assign 1_n792 = 1_n4138 & 1_n239;
assign 1_n3431 = ~(1_n6206 ^ 1_n2170);
assign 1_n11871 = ~1_n761;
assign 1_n8553 = ~(1_n4271 ^ 1_n9348);
assign 1_n12221 = ~1_n8156;
assign 1_n8042 = 1_n2296 | 1_n7254;
assign 1_n5209 = 1_n655 & 1_n2914;
assign 1_n8075 = ~(1_n4439 | 1_n2956);
assign 1_n12388 = 1_n7424;
assign 1_n1684 = 1_n5039 | 1_n7821;
assign 1_n12516 = 1_n1651 | 1_n6265;
assign 1_n9068 = ~1_n3709;
assign 1_n12498 = 1_n12013 & 1_n1632;
assign 1_n908 = 1_n10293 ^ 1_n5480;
assign 1_n10222 = ~(1_n12715 | 1_n11027);
assign 1_n3100 = ~(1_n12533 ^ 1_n3694);
assign 1_n4962 = 1_n2692 | 1_n3981;
assign 1_n4277 = 1_n734 | 1_n493;
assign 1_n7092 = ~(1_n1974 ^ 1_n1595);
assign 1_n12874 = 1_n5795 | 1_n5510;
assign 1_n2352 = ~1_n10657;
assign 1_n1196 = ~(1_n4651 ^ 1_n12118);
assign 1_n8710 = ~1_n10343;
assign 1_n8892 = ~1_n10479;
assign 1_n6753 = 1_n10018 | 1_n3981;
assign 1_n8120 = 1_n9350 | 1_n10627;
assign 1_n3957 = 1_n3225 | 1_n11668;
assign 1_n12301 = ~(1_n9516 ^ 1_n11789);
assign 1_n8746 = ~(1_n13205 ^ 1_n4310);
assign 1_n11313 = 1_n3696 | 1_n447;
assign 1_n9635 = ~1_n1603;
assign 1_n9276 = ~1_n9685;
assign 1_n7289 = 1_n1416 | 1_n10696;
assign 1_n8360 = ~1_n6826;
assign 1_n10379 = ~(1_n6412 ^ 1_n12763);
assign 1_n6671 = 1_n5749 | 1_n8534;
assign 1_n8574 = 1_n440 | 1_n5431;
assign 1_n12160 = ~(1_n7123 ^ 1_n1119);
assign 1_n11079 = 1_n5508 & 1_n861;
assign 1_n7804 = ~(1_n8276 ^ 1_n2905);
assign 1_n7489 = ~(1_n11873 | 1_n4529);
assign 1_n7947 = 1_n12713 | 1_n7082;
assign 1_n12305 = ~(1_n10077 ^ 1_n9229);
assign 1_n4583 = 1_n2353 & 1_n5542;
assign 1_n12101 = 1_n10575 ^ 1_n5170;
assign 1_n3462 = ~(1_n10152 | 1_n5368);
assign 1_n1612 = ~(1_n590 ^ 1_n12977);
assign 1_n6773 = ~(1_n7645 ^ 1_n1200);
assign 1_n11132 = ~1_n1273;
assign 1_n8212 = ~1_n7051;
assign 1_n11392 = 1_n5271 | 1_n8490;
assign 1_n9881 = 1_n5634 | 1_n5242;
assign 1_n10289 = 1_n1705 & 1_n2788;
assign 1_n9457 = ~(1_n924 ^ 1_n2938);
assign 1_n4796 = ~1_n13058;
assign 1_n12780 = 1_n5581 | 1_n5173;
assign 1_n6324 = ~(1_n11187 ^ 1_n6474);
assign 1_n10775 = ~(1_n6809 ^ 1_n11000);
assign 1_n8393 = 1_n4022 | 1_n177;
assign 1_n12703 = ~(1_n733 ^ 1_n2200);
assign 1_n3792 = 1_n10650 & 1_n921;
assign 1_n1535 = ~(1_n11472 ^ 1_n11949);
assign 1_n2918 = 1_n3318 & 1_n5714;
assign 1_n1564 = 1_n11411 & 1_n6168;
assign 1_n2109 = ~1_n10142;
assign 1_n7019 = 1_n1185 | 1_n1669;
assign 1_n11279 = 1_n12086 & 1_n11988;
assign 1_n11896 = ~(1_n1205 ^ 1_n12146);
assign 1_n4937 = 1_n9080 | 1_n9159;
assign 1_n827 = ~(1_n9726 ^ 1_n8962);
assign 1_n9927 = 1_n13051 | 1_n2544;
assign 1_n6973 = 1_n7386 & 1_n5745;
assign 1_n2278 = ~1_n8940;
assign 1_n5918 = ~(1_n11961 ^ 1_n12571);
assign 1_n13105 = 1_n2713 & 1_n7325;
assign 1_n2332 = ~1_n3076;
assign 1_n6994 = ~(1_n10306 ^ 1_n8678);
assign 1_n11168 = 1_n13082 | 1_n7221;
assign 1_n4834 = ~(1_n1410 ^ 1_n8046);
assign 1_n4627 = 1_n5329 | 1_n4503;
assign 1_n10260 = 1_n756 | 1_n5221;
assign 1_n11186 = ~(1_n6838 | 1_n12587);
assign 1_n11043 = ~(1_n1730 ^ 1_n7077);
assign 1_n11290 = 1_n10201 & 1_n7204;
assign 1_n2001 = ~(1_n4556 ^ 1_n135);
assign 1_n12322 = 1_n3630 | 1_n12328;
assign 1_n4608 = 1_n3986 | 1_n5716;
assign 1_n3489 = ~1_n10613;
assign 1_n8874 = 1_n6516 & 1_n9085;
assign 1_n5659 = 1_n10696 | 1_n9075;
assign 1_n142 = ~1_n2370;
assign 1_n5207 = ~(1_n7668 ^ 1_n12232);
assign 1_n8864 = ~1_n9270;
assign 1_n10147 = 1_n2057 & 1_n10063;
assign 1_n9728 = 1_n4080 | 1_n7723;
assign 1_n5352 = 1_n9309 | 1_n8005;
assign 1_n5113 = 1_n5694 | 1_n4947;
assign 1_n6437 = ~(1_n2358 | 1_n8462);
assign 1_n11482 = 1_n10928 ^ 1_n4155;
assign 1_n1895 = 1_n7301 & 1_n1274;
assign 1_n4807 = 1_n2800 & 1_n2466;
assign 1_n1032 = 1_n11815 & 1_n191;
assign 1_n8737 = ~(1_n9173 ^ 1_n13100);
assign 1_n8064 = 1_n6557 | 1_n1570;
assign 1_n10847 = ~(1_n11384 | 1_n11141);
assign 1_n2469 = 1_n8639 | 1_n10935;
assign 1_n3206 = 1_n13085 & 1_n12696;
assign 1_n9949 = 1_n5358 | 1_n5011;
assign 1_n10423 = ~(1_n8628 ^ 1_n1021);
assign 1_n11065 = 1_n5757 | 1_n9147;
assign 1_n4757 = 1_n3158 | 1_n4724;
assign 1_n9708 = 1_n9934 | 1_n12388;
assign 1_n5660 = 1_n338 | 1_n5076;
assign 1_n7530 = 1_n6210;
assign 1_n108 = ~(1_n3841 ^ 1_n1829);
assign 1_n8215 = ~(1_n4507 | 1_n1342);
assign 1_n12526 = 1_n8416 & 1_n12590;
assign 1_n650 = ~1_n8233;
assign 1_n6388 = 1_n7865 | 1_n3149;
assign 1_n6793 = 1_n1353 | 1_n9159;
assign 1_n1357 = ~1_n3543;
assign 1_n12068 = 1_n5676 & 1_n3530;
assign 1_n7922 = ~(1_n2621 | 1_n3220);
assign 1_n4996 = ~(1_n11799 ^ 1_n8669);
assign 1_n866 = 1_n1248 | 1_n10878;
assign 1_n5541 = ~(1_n966 | 1_n7336);
assign 1_n7257 = ~1_n5277;
assign 1_n11608 = ~(1_n12682 ^ 1_n9362);
assign 1_n5301 = 1_n11742 | 1_n13125;
assign 1_n12510 = 1_n5415 | 1_n167;
assign 1_n5168 = ~1_n11734;
assign 1_n6338 = 1_n4370 | 1_n8348;
assign 1_n1502 = ~(1_n4383 ^ 1_n3566);
assign 1_n11723 = ~1_n4330;
assign 1_n7531 = ~(1_n5224 ^ 1_n37);
assign 1_n9427 = ~(1_n9879 | 1_n12983);
assign 1_n10803 = ~(1_n5100 ^ 1_n10185);
assign 1_n7807 = 1_n8064 | 1_n6299;
assign 1_n11635 = ~1_n7161;
assign 1_n1376 = 1_n2301 | 1_n7476;
assign 1_n11841 = 1_n6139 & 1_n6490;
assign 1_n2553 = 1_n1067 | 1_n1195;
assign 1_n12528 = 1_n5265 | 1_n10871;
assign 1_n9613 = ~(1_n10219 ^ 1_n11411);
assign 1_n8738 = ~(1_n3357 | 1_n3012);
assign 1_n3377 = 1_n6726 | 1_n10179;
assign 1_n2180 = ~(1_n2395 ^ 1_n1615);
assign 1_n10032 = ~1_n11734;
assign 1_n1359 = 1_n318 | 1_n1985;
assign 1_n4004 = 1_n6572 & 1_n5888;
assign 1_n10717 = 1_n4000 | 1_n4223;
assign 1_n4098 = ~1_n11640;
assign 1_n13149 = 1_n4161 | 1_n2970;
assign 1_n11250 = 1_n4665 | 1_n10871;
assign 1_n4142 = ~(1_n1575 ^ 1_n8622);
assign 1_n3493 = ~1_n10860;
assign 1_n6025 = ~1_n322;
assign 1_n1320 = ~1_n11109;
assign 1_n231 = 1_n4969 | 1_n3276;
assign 1_n10180 = 1_n6518 | 1_n557;
assign 1_n7069 = 1_n654 & 1_n230;
assign 1_n2747 = ~1_n1397;
assign 1_n13122 = ~1_n4376;
assign 1_n10735 = ~(1_n2297 | 1_n3421);
assign 1_n2585 = ~(1_n3941 ^ 1_n12658);
assign 1_n13007 = 1_n12846 & 1_n12486;
assign 1_n10278 = 1_n11232 & 1_n7243;
assign 1_n6393 = 1_n4771 | 1_n12332;
assign 1_n2356 = 1_n12249 | 1_n8563;
assign 1_n5773 = 1_n11010 | 1_n9046;
assign 1_n1774 = 1_n11294 & 1_n10748;
assign 1_n1443 = ~(1_n4825 ^ 1_n7165);
assign 1_n2170 = ~(1_n12236 ^ 1_n4835);
assign 1_n882 = ~1_n6965;
assign 1_n10248 = 1_n8600 | 1_n1804;
assign 1_n10864 = ~(1_n5130 ^ 1_n10113);
assign 1_n9159 = 1_n2406;
assign 1_n3933 = 1_n4587 | 1_n9251;
assign 1_n13102 = 1_n9416 | 1_n7203;
assign 1_n5265 = ~1_n9669;
assign 1_n6242 = 1_n9934 | 1_n1570;
assign 1_n10358 = ~(1_n2878 | 1_n12891);
assign 1_n12556 = 1_n5404 | 1_n5721;
assign 1_n2726 = ~1_n9475;
assign 1_n11286 = 1_n7836 | 1_n11768;
assign 1_n12197 = ~(1_n314 ^ 1_n11253);
assign 1_n1461 = ~(1_n5567 | 1_n11563);
assign 1_n1609 = 1_n8449 & 1_n1533;
assign 1_n9071 = 1_n12843 | 1_n8988;
assign 1_n4066 = ~1_n7745;
assign 1_n175 = 1_n2041 | 1_n584;
assign 1_n3793 = ~(1_n10765 | 1_n852);
assign 1_n1898 = ~(1_n5861 | 1_n7548);
assign 1_n4934 = 1_n3364 | 1_n11007;
assign 1_n6402 = ~1_n11339;
assign 1_n1091 = 1_n4108 | 1_n3554;
assign 1_n3986 = 1_n10761 | 1_n6265;
assign 1_n2002 = 1_n5725 & 1_n4451;
assign 1_n2392 = 1_n10180 & 1_n10749;
assign 1_n2485 = ~1_n624;
assign 1_n3730 = 1_n8615 | 1_n4230;
assign 1_n10616 = ~1_n2513;
assign 1_n12064 = 1_n12342 & 1_n9977;
assign 1_n4007 = ~(1_n976 | 1_n260);
assign 1_n11457 = 1_n2570 & 1_n6923;
assign 1_n12314 = ~(1_n12809 ^ 1_n11267);
assign 1_n1509 = 1_n9016 | 1_n206;
assign 1_n11512 = 1_n12859 | 1_n10971;
assign 1_n4977 = ~(1_n1470 ^ 1_n10614);
assign 1_n4405 = 1_n10598 & 1_n4480;
assign 1_n12957 = ~1_n937;
assign 1_n1264 = 1_n11799 | 1_n3187;
assign 1_n6177 = ~(1_n6196 ^ 1_n12831);
assign 1_n8408 = 1_n10113 & 1_n7411;
assign 1_n4955 = ~1_n5454;
assign 1_n8889 = ~(1_n4692 ^ 1_n556);
assign 1_n11502 = 1_n544 | 1_n322;
assign 1_n7131 = 1_n3522 | 1_n8086;
assign 1_n3009 = 1_n2226 | 1_n9309;
assign 1_n10926 = 1_n6027 & 1_n6898;
assign 1_n625 = 1_n5638 & 1_n6888;
assign 1_n1214 = ~(1_n1297 ^ 1_n6984);
assign 1_n11944 = ~(1_n903 ^ 1_n12197);
assign 1_n8178 = ~(1_n2936 ^ 1_n9356);
assign 1_n6060 = 1_n1238 & 1_n3819;
assign 1_n2609 = 1_n5613 & 1_n12555;
assign 1_n967 = ~1_n5322;
assign 1_n12218 = ~(1_n2101 ^ 1_n4794);
assign 1_n11769 = ~(1_n11971 ^ 1_n12102);
assign 1_n3602 = 1_n8980 | 1_n7509;
assign 1_n8378 = 1_n8862 | 1_n12072;
assign 1_n11993 = ~(1_n10861 ^ 1_n6736);
assign 1_n4853 = 1_n1725 | 1_n12948;
assign 1_n2117 = 1_n3837 & 1_n6327;
assign 1_n406 = ~1_n10657;
assign 1_n12152 = ~(1_n7929 | 1_n12106);
assign 1_n11819 = ~(1_n783 ^ 1_n8893);
assign 1_n10776 = ~(1_n8135 ^ 1_n11536);
assign 1_n8645 = ~1_n11835;
assign 1_n9486 = 1_n7951 & 1_n7921;
assign 1_n5022 = ~(1_n7414 ^ 1_n8845);
assign 1_n237 = ~1_n10642;
assign 1_n2240 = 1_n10883 | 1_n9075;
assign 1_n9437 = 1_n10419 ^ 1_n2000;
assign 1_n1669 = ~(1_n9676 ^ 1_n11367);
assign 1_n6191 = 1_n202 | 1_n1985;
assign 1_n3690 = ~1_n880;
assign 1_n8880 = 1_n10591 | 1_n7723;
assign 1_n1658 = ~(1_n11496 | 1_n7893);
assign 1_n3866 = ~1_n3815;
assign 1_n11536 = ~(1_n12140 ^ 1_n3989);
assign 1_n434 = 1_n1651 | 1_n4936;
assign 1_n10101 = 1_n10392 ^ 1_n9655;
assign 1_n6961 = 1_n9154 | 1_n12501;
assign 1_n13022 = ~(1_n9637 ^ 1_n3649);
assign 1_n4074 = 1_n3335 & 1_n11178;
assign 1_n2432 = ~(1_n4521 ^ 1_n2497);
assign 1_n7553 = ~(1_n2841 ^ 1_n11528);
assign 1_n3181 = ~(1_n11592 ^ 1_n4656);
assign 1_n1462 = ~(1_n7552 | 1_n10793);
assign 1_n2088 = 1_n6375 | 1_n10319;
assign 1_n11484 = ~(1_n12581 ^ 1_n12905);
assign 1_n5037 = ~1_n4413;
assign 1_n17 = 1_n11683 | 1_n10319;
assign 1_n4888 = 1_n9353 & 1_n3085;
assign 1_n5219 = ~(1_n12804 ^ 1_n8594);
assign 1_n11151 = ~(1_n1758 ^ 1_n6034);
assign 1_n7967 = ~(1_n1810 ^ 1_n1755);
assign 1_n11664 = ~1_n5375;
assign 1_n9034 = ~(1_n2799 ^ 1_n6544);
assign 1_n2183 = ~1_n9591;
assign 1_n4164 = 1_n1906 & 1_n6095;
assign 1_n10683 = 1_n9917 | 1_n11446;
assign 1_n9835 = 1_n4370 | 1_n4724;
assign 1_n3039 = ~(1_n1352 | 1_n8037);
assign 1_n5782 = ~1_n411;
assign 1_n12357 = ~1_n4015;
assign 1_n250 = 1_n11356 | 1_n8702;
assign 1_n10897 = 1_n5456 & 1_n8833;
assign 1_n4695 = 1_n1889 & 1_n4320;
assign 1_n4607 = 1_n12911 | 1_n2792;
assign 1_n10511 = ~(1_n10217 ^ 1_n2837);
assign 1_n1824 = ~(1_n8067 | 1_n10817);
assign 1_n9954 = 1_n8739 | 1_n8036;
assign 1_n8201 = ~(1_n7230 ^ 1_n3622);
assign 1_n11374 = 1_n12758 | 1_n4724;
assign 1_n6765 = ~(1_n1601 ^ 1_n7384);
assign 1_n9161 = 1_n12768 | 1_n1570;
assign 1_n3266 = 1_n1772 | 1_n7701;
assign 1_n6702 = ~(1_n7852 ^ 1_n1770);
assign 1_n1546 = 1_n6381 | 1_n4947;
assign 1_n12609 = 1_n4891 & 1_n6360;
assign 1_n11183 = 1_n1638 | 1_n10029;
assign 1_n5095 = ~(1_n5121 ^ 1_n4516);
assign 1_n7354 = 1_n542 | 1_n6265;
assign 1_n7912 = ~(1_n11709 | 1_n3447);
assign 1_n6400 = ~(1_n5453 ^ 1_n12836);
assign 1_n3492 = 1_n5407 | 1_n3648;
assign 1_n8417 = ~(1_n6535 | 1_n4064);
assign 1_n9254 = ~(1_n12467 | 1_n9561);
assign 1_n5277 = 1_n6894 & 1_n6980;
assign 1_n4810 = 1_n5182 | 1_n11521;
assign 1_n4249 = 1_n5526 & 1_n1691;
assign 1_n12449 = 1_n12617 | 1_n9808;
assign 1_n10342 = ~(1_n7802 ^ 1_n5336);
assign 1_n2101 = ~(1_n267 ^ 1_n12762);
assign 1_n8727 = ~(1_n5251 | 1_n4065);
assign 1_n3606 = ~(1_n890 ^ 1_n7209);
assign 1_n968 = 1_n11113 | 1_n9223;
assign 1_n3784 = ~1_n12065;
assign 1_n176 = ~(1_n1349 | 1_n4259);
assign 1_n2206 = ~(1_n6371 ^ 1_n10071);
assign 1_n3530 = 1_n3460 | 1_n12695;
assign 1_n6047 = 1_n7554 & 1_n591;
assign 1_n719 = ~1_n10745;
assign 1_n10900 = ~1_n1364;
assign 1_n2102 = 1_n7514 & 1_n7778;
assign 1_n12467 = ~(1_n5005 | 1_n13110);
assign 1_n8348 = 1_n3671;
assign 1_n9310 = ~1_n5470;
assign 1_n6447 = ~(1_n7256 ^ 1_n832);
assign 1_n651 = ~1_n9027;
assign 1_n3633 = ~1_n6973;
assign 1_n3854 = ~1_n353;
assign 1_n5784 = 1_n3225 | 1_n8490;
assign 1_n8275 = ~(1_n9033 | 1_n5722);
assign 1_n5847 = ~1_n6820;
assign 1_n4756 = 1_n9248 | 1_n5006;
assign 1_n1613 = ~(1_n3339 ^ 1_n12878);
assign 1_n3336 = ~1_n6189;
assign 1_n4378 = 1_n5911 & 1_n3603;
assign 1_n9839 = ~(1_n2994 ^ 1_n8110);
assign 1_n5531 = 1_n10139 | 1_n8101;
assign 1_n4430 = ~1_n1225;
assign 1_n11913 = ~(1_n11936 ^ 1_n3252);
assign 1_n10706 = ~(1_n1640 | 1_n1704);
assign 1_n10075 = 1_n10738 & 1_n11673;
assign 1_n11416 = ~(1_n10385 ^ 1_n3863);
assign 1_n1258 = ~1_n6597;
assign 1_n2806 = 1_n872 | 1_n7252;
assign 1_n11943 = 1_n7546 | 1_n2490;
assign 1_n9166 = ~(1_n10325 ^ 1_n1929);
assign 1_n445 = ~1_n5065;
assign 1_n4716 = ~1_n8369;
assign 1_n6150 = 1_n11927 & 1_n1300;
assign 1_n3915 = 1_n11263 | 1_n13081;
assign 1_n6752 = ~(1_n3171 | 1_n5154);
assign 1_n5694 = ~1_n3677;
assign 1_n3143 = 1_n3359 & 1_n7570;
assign 1_n784 = 1_n930 | 1_n10463;
assign 1_n5255 = ~(1_n4304 | 1_n11885);
assign 1_n7155 = 1_n316 & 1_n4084;
assign 1_n12414 = ~(1_n11793 ^ 1_n11177);
assign 1_n1468 = ~(1_n11534 | 1_n3440);
assign 1_n1402 = ~1_n10606;
assign 1_n7736 = ~(1_n12013 ^ 1_n8222);
assign 1_n9807 = 1_n6672 | 1_n4420;
assign 1_n875 = 1_n13201 & 1_n834;
assign 1_n3225 = 1_n6193;
assign 1_n8950 = ~1_n11429;
assign 1_n3563 = 1_n13028 | 1_n8777;
assign 1_n3438 = ~(1_n11900 ^ 1_n10816);
assign 1_n3808 = ~(1_n2286 ^ 1_n647);
assign 1_n8068 = 1_n7637 | 1_n12171;
assign 1_n6082 = 1_n3800 & 1_n10269;
assign 1_n13176 = 1_n11408 & 1_n7911;
assign 1_n9293 = 1_n8865 | 1_n8819;
assign 1_n5719 = 1_n5932 | 1_n2633;
assign 1_n351 = 1_n4537 & 1_n5962;
assign 1_n4251 = 1_n48 | 1_n3981;
assign 1_n4689 = ~1_n3797;
assign 1_n12337 = 1_n332 | 1_n12733;
assign 1_n1560 = 1_n787 | 1_n2059;
assign 1_n3273 = 1_n987 | 1_n5242;
assign 1_n10054 = ~(1_n11070 | 1_n3503);
assign 1_n9858 = ~(1_n8616 ^ 1_n799);
assign 1_n4484 = ~1_n919;
assign 1_n11779 = ~1_n7659;
assign 1_n8473 = ~(1_n2347 ^ 1_n12346);
assign 1_n5184 = 1_n4356 & 1_n4010;
assign 1_n12069 = ~1_n11537;
assign 1_n2748 = ~(1_n6750 | 1_n7572);
assign 1_n6141 = 1_n11247 & 1_n2812;
assign 1_n1587 = ~1_n2498;
assign 1_n9497 = ~1_n1563;
assign 1_n12340 = 1_n3498 | 1_n10106;
assign 1_n9405 = ~(1_n11215 | 1_n2375);
assign 1_n10955 = ~(1_n7882 ^ 1_n1923);
assign 1_n3551 = 1_n6731 & 1_n11901;
assign 1_n6821 = 1_n11513 & 1_n312;
assign 1_n9487 = 1_n98 | 1_n8702;
assign 1_n1786 = 1_n1645 | 1_n6169;
assign 1_n6467 = 1_n3760 & 1_n5446;
assign 1_n4024 = 1_n9387 & 1_n9997;
assign 1_n8080 = ~(1_n12270 ^ 1_n1604);
assign 1_n7127 = ~1_n7452;
assign 1_n2022 = ~1_n5052;
assign 1_n5529 = 1_n7176 | 1_n8366;
assign 1_n12256 = 1_n8891 | 1_n3961;
assign 1_n4208 = ~1_n12289;
assign 1_n2159 = 1_n7272 ^ 1_n195;
assign 1_n1845 = ~(1_n6322 ^ 1_n10649);
assign 1_n3388 = ~(1_n10829 | 1_n6071);
assign 1_n4662 = 1_n11 & 1_n8956;
assign 1_n12905 = ~(1_n6314 ^ 1_n8913);
assign 1_n7696 = 1_n10212 & 1_n11947;
assign 1_n7710 = ~1_n7906;
assign 1_n4546 = 1_n2795 & 1_n11654;
assign 1_n2421 = 1_n4836 & 1_n12883;
assign 1_n3255 = 1_n3505 | 1_n9537;
assign 1_n500 = 1_n7782 | 1_n4169;
assign 1_n528 = 1_n8940 & 1_n8290;
assign 1_n605 = 1_n11914 & 1_n12760;
assign 1_n4121 = 1_n3006 & 1_n12853;
assign 1_n3605 = 1_n13154 | 1_n6635;
assign 1_n3679 = 1_n5478 | 1_n6293;
assign 1_n1439 = 1_n10974 | 1_n8534;
assign 1_n242 = ~(1_n7699 | 1_n8703);
assign 1_n8480 = 1_n12942 & 1_n475;
assign 1_n12286 = ~(1_n9642 ^ 1_n714);
assign 1_n2264 = ~1_n10606;
assign 1_n7754 = ~(1_n27 ^ 1_n11353);
assign 1_n1765 = 1_n4221 | 1_n3225;
assign 1_n4696 = ~1_n4114;
assign 1_n12524 = ~(1_n12829 ^ 1_n6461);
assign 1_n2910 = ~1_n5075;
assign 1_n10097 = 1_n12024 | 1_n8568;
assign 1_n3231 = 1_n6168 & 1_n4470;
assign 1_n10497 = 1_n11218 | 1_n2958;
assign 1_n5102 = ~(1_n8807 ^ 1_n12275);
assign 1_n1427 = 1_n5679 | 1_n11107;
assign 1_n2009 = ~(1_n2533 ^ 1_n8042);
assign 1_n1151 = ~1_n4303;
assign 1_n5218 = 1_n6926 & 1_n4418;
assign 1_n5872 = 1_n10893 | 1_n6364;
assign 1_n385 = 1_n12032 | 1_n12388;
assign 1_n12039 = ~(1_n6828 ^ 1_n4917);
assign 1_n12390 = 1_n7371 & 1_n8438;
assign 1_n6941 = ~(1_n4965 | 1_n339);
assign 1_n2850 = 1_n877 | 1_n11898;
assign 1_n7094 = ~(1_n707 ^ 1_n4307);
assign 1_n8848 = ~1_n6021;
assign 1_n11830 = ~(1_n11584 ^ 1_n9738);
assign 1_n11532 = ~(1_n7236 | 1_n2099);
assign 1_n960 = ~(1_n7618 ^ 1_n4617);
assign 1_n638 = 1_n1896 & 1_n11005;
assign 1_n3124 = 1_n924 | 1_n5776;
assign 1_n775 = ~(1_n11046 ^ 1_n6030);
assign 1_n8661 = ~1_n7161;
assign 1_n3847 = 1_n572 | 1_n11375;
assign 1_n6348 = 1_n12878 | 1_n8118;
assign 1_n5911 = 1_n12082 | 1_n4786;
assign 1_n6778 = 1_n8681 | 1_n5797;
assign 1_n13196 = 1_n11054 | 1_n1463;
assign 1_n12383 = ~1_n834;
assign 1_n10753 = 1_n9674 | 1_n1255;
assign 1_n4480 = 1_n2487 | 1_n5242;
assign 1_n3332 = ~(1_n3139 ^ 1_n9470);
assign 1_n9463 = ~(1_n5737 | 1_n7643);
assign 1_n9290 = 1_n9259 & 1_n7355;
assign 1_n10895 = 1_n12768 | 1_n6265;
assign 1_n3044 = ~1_n10102;
assign 1_n1795 = ~1_n7500;
assign 1_n256 = 1_n2394 & 1_n5096;
assign 1_n12440 = ~(1_n7403 ^ 1_n4034);
assign 1_n35 = 1_n3707 | 1_n5207;
assign 1_n9605 = 1_n549 | 1_n5;
assign 1_n1155 = ~1_n1910;
assign 1_n6368 = 1_n10828 & 1_n3346;
assign 1_n11875 = ~(1_n8302 ^ 1_n7366);
assign 1_n8502 = 1_n11493 & 1_n5529;
assign 1_n1090 = ~(1_n371 ^ 1_n439);
assign 1_n7671 = ~(1_n7699 ^ 1_n874);
assign 1_n11397 = 1_n11055 ^ 1_n139;
assign 1_n11870 = 1_n8390 & 1_n2076;
assign 1_n4181 = ~(1_n1166 | 1_n5525);
assign 1_n9625 = 1_n12808 | 1_n8857;
assign 1_n12674 = 1_n10217 | 1_n6442;
assign 1_n11851 = 1_n12084 & 1_n13054;
assign 1_n6353 = ~(1_n1716 ^ 1_n835);
assign 1_n13054 = ~(1_n12941 ^ 1_n1992);
assign 1_n1626 = 1_n10404 | 1_n3997;
assign 1_n6339 = ~(1_n3388 | 1_n12140);
assign 1_n9400 = ~1_n2252;
assign 1_n9396 = ~1_n4797;
assign 1_n9833 = 1_n2809 & 1_n9013;
assign 1_n2487 = ~1_n1724;
assign 1_n11260 = 1_n968 | 1_n2923;
assign 1_n3037 = 1_n9160 & 1_n2335;
assign 1_n9618 = ~1_n9952;
assign 1_n7450 = 1_n5313 | 1_n12973;
assign 1_n8905 = ~1_n3644;
assign 1_n6710 = ~1_n4452;
assign 1_n2132 = 1_n4600 | 1_n1723;
assign 1_n12918 = 1_n1425 | 1_n11689;
assign 1_n8347 = 1_n9003 & 1_n1606;
assign 1_n11966 = ~(1_n3427 | 1_n3949);
assign 1_n8935 = ~1_n12553;
assign 1_n12421 = 1_n3528 & 1_n10918;
assign 1_n9852 = ~(1_n11206 ^ 1_n1845);
assign 1_n11120 = 1_n2538 | 1_n2059;
assign 1_n11404 = ~1_n12482;
assign 1_n11015 = 1_n4228 | 1_n12684;
assign 1_n8224 = ~(1_n9860 ^ 1_n1761);
assign 1_n4195 = ~(1_n3061 ^ 1_n13192);
assign 1_n6031 = ~(1_n12603 ^ 1_n1910);
assign 1_n3719 = ~1_n12461;
assign 1_n10005 = ~1_n5319;
assign 1_n3452 = ~(1_n11964 | 1_n10766);
assign 1_n1285 = ~(1_n11736 ^ 1_n12015);
assign 1_n10421 = ~1_n9915;
assign 1_n6936 = 1_n3822 | 1_n3339;
assign 1_n369 = ~(1_n5514 ^ 1_n7916);
assign 1_n659 = ~(1_n12690 ^ 1_n7511);
assign 1_n4086 = 1_n93 & 1_n10113;
assign 1_n11581 = 1_n3016 & 1_n7018;
assign 1_n1989 = ~1_n9041;
assign 1_n7823 = 1_n10794 & 1_n10131;
assign 1_n4194 = ~1_n8230;
assign 1_n2834 = 1_n10731 | 1_n5485;
assign 1_n1253 = ~(1_n5475 ^ 1_n974);
assign 1_n5263 = ~(1_n347 ^ 1_n6797);
assign 1_n12435 = 1_n6970 | 1_n4445;
assign 1_n2437 = ~1_n1055;
assign 1_n6370 = ~1_n9732;
assign 1_n1530 = 1_n4380 & 1_n10093;
assign 1_n8639 = 1_n9190 & 1_n3532;
assign 1_n9398 = 1_n12580 | 1_n4834;
assign 1_n12020 = ~(1_n4084 ^ 1_n316);
assign 1_n12192 = 1_n3281 | 1_n4116;
assign 1_n1918 = 1_n8926 | 1_n5736;
assign 1_n5114 = 1_n4371 & 1_n4078;
assign 1_n924 = ~(1_n7706 ^ 1_n679);
assign 1_n6131 = 1_n5271 | 1_n1026;
assign 1_n11811 = 1_n10274 | 1_n11527;
assign 1_n3109 = 1_n7872 | 1_n8563;
assign 1_n3522 = 1_n5482 | 1_n1303;
assign 1_n7370 = 1_n6106 | 1_n5986;
assign 1_n11299 = ~(1_n11832 ^ 1_n4040);
assign 1_n2407 = 1_n10517 | 1_n11735;
assign 1_n10428 = 1_n10029 | 1_n8030;
assign 1_n8687 = 1_n1975 | 1_n6454;
assign 1_n6852 = ~(1_n2519 ^ 1_n8591);
assign 1_n10457 = 1_n2458 & 1_n12306;
assign 1_n9177 = ~1_n10455;
assign 1_n8973 = 1_n9635 | 1_n3455;
assign 1_n4107 = ~1_n5962;
assign 1_n9593 = ~(1_n11783 | 1_n12079);
assign 1_n4023 = 1_n4580 & 1_n12844;
assign 1_n7301 = 1_n9364 | 1_n4300;
assign 1_n7966 = ~1_n4357;
assign 1_n11376 = 1_n6769 | 1_n177;
assign 1_n8634 = 1_n5679 | 1_n8030;
assign 1_n787 = ~1_n6818;
assign 1_n12976 = ~(1_n3375 ^ 1_n480);
assign 1_n362 = ~(1_n6930 ^ 1_n9031);
assign 1_n6083 = ~(1_n13227 ^ 1_n2770);
assign 1_n7891 = 1_n2276 | 1_n5430;
assign 1_n12767 = 1_n8593 & 1_n565;
assign 1_n4005 = 1_n6438 | 1_n11668;
assign 1_n11339 = 1_n1963 & 1_n1008;
assign 1_n2805 = ~(1_n6831 ^ 1_n5967);
assign 1_n2410 = ~(1_n3705 | 1_n13177);
assign 1_n2793 = ~1_n102;
assign 1_n9914 = 1_n7647 | 1_n10387;
assign 1_n12513 = ~(1_n9807 ^ 1_n12790);
assign 1_n2343 = ~(1_n2146 ^ 1_n9163);
assign 1_n1871 = 1_n7792 ^ 1_n6851;
assign 1_n11619 = ~(1_n1169 | 1_n5620);
assign 1_n2658 = ~(1_n3696 ^ 1_n4885);
assign 1_n782 = 1_n4480 | 1_n10598;
assign 1_n2086 = 1_n4772 | 1_n12495;
assign 1_n10618 = 1_n7313 | 1_n2931;
assign 1_n8156 = ~(1_n577 ^ 1_n780);
assign 1_n2914 = 1_n11729 | 1_n7723;
assign 1_n9074 = 1_n5671 & 1_n5536;
assign 1_n143 = ~(1_n562 ^ 1_n6398);
assign 1_n10493 = 1_n5103 & 1_n3768;
assign 1_n9961 = ~(1_n12989 ^ 1_n7143);
assign 1_n410 = 1_n7205 | 1_n9985;
assign 1_n12515 = ~(1_n8647 ^ 1_n4168);
assign 1_n1625 = ~1_n3841;
assign 1_n8313 = 1_n9931 | 1_n4373;
assign 1_n1759 = 1_n5679 | 1_n10871;
assign 1_n4312 = 1_n8139 & 1_n9906;
assign 1_n7293 = 1_n5261 | 1_n9223;
assign 1_n832 = 1_n6659 & 1_n9071;
assign 1_n1541 = ~(1_n2182 ^ 1_n5278);
assign 1_n235 = ~1_n8742;
assign 1_n5091 = 1_n13026 | 1_n7961;
assign 1_n5156 = ~(1_n2598 ^ 1_n10985);
assign 1_n10346 = 1_n9843 | 1_n11394;
assign 1_n41 = ~(1_n12771 | 1_n5538);
assign 1_n9036 = ~(1_n10378 ^ 1_n4249);
assign 1_n3024 = 1_n11328 | 1_n3763;
assign 1_n4856 = ~(1_n10639 ^ 1_n2921);
assign 1_n3027 = ~(1_n12222 | 1_n4336);
assign 1_n7263 = ~(1_n9294 ^ 1_n212);
assign 1_n10193 = ~(1_n4978 | 1_n9821);
assign 1_n1484 = 1_n10060 & 1_n6866;
assign 1_n10978 = ~1_n9609;
assign 1_n2049 = 1_n5148 | 1_n4724;
assign 1_n6997 = ~(1_n3934 ^ 1_n2414);
assign 1_n527 = 1_n6245 | 1_n6769;
assign 1_n13239 = ~1_n6487;
assign 1_n12292 = 1_n1144 | 1_n10871;
assign 1_n6126 = 1_n8805 & 1_n11648;
assign 1_n4243 = ~1_n2258;
assign 1_n9459 = ~(1_n870 ^ 1_n11604);
assign 1_n12797 = ~(1_n8546 ^ 1_n1585);
assign 1_n955 = ~(1_n1599 ^ 1_n4478);
assign 1_n6371 = 1_n8757 | 1_n8490;
assign 1_n10282 = ~(1_n518 | 1_n7776);
assign 1_n139 = 1_n937 & 1_n8506;
assign 1_n11824 = 1_n4065 & 1_n5251;
assign 1_n5010 = 1_n12475 | 1_n3759;
assign 1_n831 = ~(1_n3953 ^ 1_n796);
assign 1_n262 = ~(1_n6993 | 1_n3506);
assign 1_n3108 = ~(1_n1067 ^ 1_n12303);
assign 1_n7044 = 1_n11061 & 1_n8506;
assign 1_n6232 = ~1_n12255;
assign 1_n9217 = 1_n10705 | 1_n2561;
assign 1_n11283 = 1_n97 | 1_n1043;
assign 1_n12043 = ~1_n10091;
assign 1_n12729 = ~(1_n5158 ^ 1_n3861);
assign 1_n11226 = ~1_n5884;
assign 1_n6905 = 1_n8196 & 1_n11269;
assign 1_n1577 = ~1_n2827;
assign 1_n9370 = ~(1_n5062 | 1_n7262);
assign 1_n11939 = ~(1_n1653 ^ 1_n10307);
assign 1_n109 = 1_n2464 ^ 1_n8123;
assign 1_n10533 = 1_n2689 | 1_n10179;
assign 1_n3858 = ~1_n5671;
assign 1_n5675 = ~(1_n336 ^ 1_n7290);
assign 1_n12085 = ~(1_n5738 ^ 1_n7365);
assign 1_n8281 = ~(1_n5704 ^ 1_n10194);
assign 1_n591 = ~1_n140;
assign 1_n4559 = 1_n4155 & 1_n3437;
assign 1_n12714 = ~(1_n10873 | 1_n8419);
assign 1_n1110 = ~(1_n5452 ^ 1_n12307);
assign 1_n12657 = ~1_n1364;
assign 1_n7295 = 1_n3194 | 1_n4680;
assign 1_n1983 = ~(1_n7772 ^ 1_n7529);
assign 1_n5321 = 1_n4454 | 1_n8268;
assign 1_n12297 = ~1_n11589;
assign 1_n654 = 1_n1719 | 1_n2686;
assign 1_n691 = 1_n11966;
assign 1_n819 = 1_n10203 & 1_n5234;
assign 1_n10240 = ~1_n5548;
assign 1_n1147 = ~(1_n983 ^ 1_n1272);
assign 1_n3073 = ~(1_n9399 ^ 1_n11841);
assign 1_n10645 = ~(1_n6168 | 1_n11411);
assign 1_n2175 = ~1_n40;
assign 1_n12847 = 1_n11940;
assign 1_n341 = 1_n52 & 1_n144;
assign 1_n10708 = 1_n866 & 1_n10428;
assign 1_n2804 = ~(1_n11659 | 1_n12945);
assign 1_n6163 = ~(1_n38 | 1_n7923);
assign 1_n2876 = ~(1_n2991 ^ 1_n9440);
assign 1_n791 = ~(1_n9684 ^ 1_n12691);
assign 1_n3578 = ~(1_n5789 ^ 1_n5437);
assign 1_n11506 = ~(1_n2982 ^ 1_n11764);
assign 1_n12816 = 1_n9773 & 1_n4576;
assign 1_n6115 = ~(1_n10429 ^ 1_n252);
assign 1_n5561 = 1_n542 | 1_n7935;
assign 1_n12884 = 1_n12897 & 1_n5133;
assign 1_n9638 = ~1_n10642;
assign 1_n11792 = ~(1_n4188 ^ 1_n427);
assign 1_n5357 = 1_n11202 & 1_n1117;
assign 1_n9495 = ~(1_n5018 ^ 1_n4477);
assign 1_n10608 = 1_n10978 | 1_n11008;
assign 1_n154 = ~1_n8820;
assign 1_n3134 = ~(1_n11303 ^ 1_n8572);
assign 1_n2846 = ~(1_n5440 ^ 1_n2244);
assign 1_n8931 = ~(1_n2298 ^ 1_n1757);
assign 1_n3427 = ~1_n854;
assign 1_n7755 = ~(1_n9769 ^ 1_n11388);
assign 1_n3102 = ~1_n3863;
assign 1_n7828 = 1_n7825 | 1_n1144;
assign 1_n11019 = ~(1_n7759 ^ 1_n3200);
assign 1_n11304 = ~(1_n10395 | 1_n102);
assign 1_n1860 = ~(1_n3144 ^ 1_n9090);
assign 1_n6803 = 1_n8315 | 1_n12847;
assign 1_n5304 = ~(1_n4317 ^ 1_n5405);
assign 1_n3638 = 1_n5191 | 1_n4070;
assign 1_n10852 = 1_n10625 & 1_n10160;
assign 1_n10745 = ~(1_n11215 ^ 1_n8214);
assign 1_n6365 = ~(1_n6954 ^ 1_n1556);
assign 1_n5462 = ~1_n873;
assign 1_n8122 = ~1_n7863;
assign 1_n6887 = 1_n2329 | 1_n177;
assign 1_n10675 = ~(1_n6123 ^ 1_n3420);
assign 1_n11247 = 1_n2832 | 1_n9943;
assign 1_n3082 = ~1_n1466;
assign 1_n3762 = ~(1_n9841 ^ 1_n12219);
assign 1_n3224 = ~(1_n11178 ^ 1_n3335);
assign 1_n6674 = 1_n5158 | 1_n3913;
assign 1_n11687 = ~(1_n11877 ^ 1_n10566);
assign 1_n5977 = 1_n8909 & 1_n3004;
assign 1_n8109 = 1_n2080 | 1_n13117;
assign 1_n3745 = ~(1_n3611 ^ 1_n13155);
assign 1_n8817 = ~1_n7113;
assign 1_n731 = ~(1_n1424 ^ 1_n1693);
assign 1_n13027 = 1_n6416 | 1_n121;
assign 1_n12419 = ~(1_n11397 ^ 1_n12903);
assign 1_n2767 = 1_n4536 | 1_n7430;
assign 1_n5220 = 1_n8188 | 1_n2738;
assign 1_n10223 = 1_n1092 & 1_n891;
assign 1_n2753 = ~(1_n11608 ^ 1_n4894);
assign 1_n8475 = ~(1_n9211 | 1_n8767);
assign 1_n4671 = ~(1_n12730 ^ 1_n328);
assign 1_n7580 = 1_n11723 | 1_n2222;
assign 1_n12702 = 1_n12765 | 1_n11447;
assign 1_n6757 = ~1_n6809;
assign 1_n675 = ~(1_n8779 ^ 1_n5828);
assign 1_n3670 = ~(1_n6229 ^ 1_n6263);
assign 1_n10932 = 1_n10938 & 1_n1841;
assign 1_n3226 = ~(1_n11129 ^ 1_n11052);
assign 1_n7026 = 1_n6202 | 1_n721;
assign 1_n10375 = 1_n5016 | 1_n4172;
assign 1_n12862 = ~(1_n8036 ^ 1_n12852);
assign 1_n4774 = 1_n602 ^ 1_n10654;
assign 1_n8074 = 1_n12732 | 1_n121;
assign 1_n12359 = 1_n12780 & 1_n2413;
assign 1_n3449 = ~(1_n12078 ^ 1_n4798);
assign 1_n10509 = ~1_n10142;
assign 1_n494 = 1_n7819 | 1_n12383;
assign 1_n7317 = 1_n10195 | 1_n12691;
assign 1_n6044 = ~(1_n6811 | 1_n11364);
assign 1_n2602 = 1_n8230 & 1_n12289;
assign 1_n4828 = 1_n10068 | 1_n12173;
assign 1_n11625 = 1_n6986 | 1_n2059;
assign 1_n9866 = ~(1_n12341 ^ 1_n8027);
assign 1_n12506 = ~(1_n2865 ^ 1_n3548);
assign 1_n8155 = 1_n7541 ^ 1_n1953;
assign 1_n2856 = 1_n4890 | 1_n6265;
assign 1_n10760 = 1_n4412 | 1_n8679;
assign 1_n10880 = 1_n8802 | 1_n6235;
assign 1_n5437 = 1_n9501 | 1_n1044;
assign 1_n11812 = ~(1_n3317 ^ 1_n7812);
assign 1_n7401 = 1_n4107 | 1_n11144;
assign 1_n8519 = ~(1_n1610 | 1_n10605);
assign 1_n7407 = ~1_n12746;
assign 1_n7606 = 1_n10941 | 1_n12746;
assign 1_n11110 = ~1_n6213;
assign 1_n12890 = ~(1_n12019 ^ 1_n620);
assign 1_n4895 = ~(1_n10815 ^ 1_n8791);
assign 1_n11755 = ~(1_n6785 ^ 1_n8691);
assign 1_n11852 = ~(1_n7711 ^ 1_n9756);
assign 1_n7329 = 1_n5328 | 1_n1463;
assign 1_n8276 = ~(1_n3405 | 1_n6752);
assign 1_n8143 = ~1_n9915;
assign 1_n6265 = 1_n138;
assign 1_n9504 = ~(1_n2974 ^ 1_n788);
assign 1_n13200 = 1_n6189 & 1_n9092;
assign 1_n12429 = ~(1_n5384 ^ 1_n4296);
assign 1_n1260 = ~(1_n8203 ^ 1_n315);
assign 1_n7504 = 1_n1250 & 1_n3113;
assign 1_n10334 = ~1_n8163;
assign 1_n11685 = 1_n8533 & 1_n2515;
assign 1_n3216 = 1_n11091 | 1_n12665;
assign 1_n4466 = 1_n5808 | 1_n3135;
assign 1_n3463 = ~(1_n9856 ^ 1_n313);
assign 1_n5436 = 1_n1747 | 1_n11423;
assign 1_n11345 = 1_n2738 | 1_n7935;
assign 1_n6584 = 1_n4937 | 1_n978;
assign 1_n1081 = ~(1_n8647 | 1_n3702);
assign 1_n11215 = 1_n813 | 1_n1144;
assign 1_n7343 = ~(1_n8043 ^ 1_n814);
assign 1_n5833 = 1_n3509 | 1_n6635;
assign 1_n5471 = ~(1_n7751 | 1_n7093);
assign 1_n5512 = 1_n12135 | 1_n6714;
assign 1_n2300 = ~(1_n6747 ^ 1_n6553);
assign 1_n198 = ~1_n1667;
assign 1_n6456 = 1_n6428 & 1_n839;
assign 1_n305 = 1_n3594 & 1_n4632;
assign 1_n7395 = ~1_n10567;
assign 1_n10921 = ~(1_n5982 ^ 1_n10827);
assign 1_n11689 = 1_n7640 & 1_n12697;
assign 1_n9072 = 1_n5892 | 1_n5942;
assign 1_n2760 = ~(1_n12462 ^ 1_n5092);
assign 1_n5883 = 1_n2734 | 1_n9921;
assign 1_n11322 = 1_n6837 | 1_n11166;
assign 1_n6916 = 1_n13227 | 1_n11028;
assign 1_n13190 = ~1_n4357;
assign 1_n10326 = ~(1_n3725 ^ 1_n263);
assign 1_n8050 = ~1_n10782;
assign 1_n4621 = ~1_n5920;
assign 1_n4374 = ~(1_n8433 ^ 1_n441);
assign 1_n28 = ~(1_n6624 ^ 1_n4993);
assign 1_n10444 = 1_n5100 & 1_n8837;
assign 1_n11749 = 1_n8053 | 1_n7935;
assign 1_n420 = 1_n11488 & 1_n12853;
assign 1_n11705 = 1_n8529 | 1_n7935;
assign 1_n11623 = ~(1_n11648 ^ 1_n2627);
assign 1_n656 = ~1_n3713;
assign 1_n3554 = 1_n12573 | 1_n1463;
assign 1_n7685 = ~(1_n5404 ^ 1_n4739);
assign 1_n8497 = ~(1_n2358 ^ 1_n2009);
assign 1_n6018 = 1_n3158 | 1_n12957;
assign 1_n11957 = 1_n640 | 1_n1808;
assign 1_n12331 = ~(1_n13208 ^ 1_n7070);
assign 1_n1063 = ~(1_n9271 ^ 1_n3925);
assign 1_n7404 = 1_n1290 | 1_n9151;
assign 1_n2769 = 1_n10825 | 1_n6869;
assign 1_n9111 = ~(1_n9488 ^ 1_n2114);
assign 1_n8925 = ~1_n209;
assign 1_n8251 = ~1_n9452;
assign 1_n11218 = ~1_n854;
assign 1_n5955 = ~(1_n12429 ^ 1_n5815);
assign 1_n2318 = 1_n4191 | 1_n5074;
assign 1_n7471 = ~1_n6644;
assign 1_n1938 = 1_n5562 | 1_n9075;
assign 1_n1038 = 1_n3164 & 1_n8928;
assign 1_n4568 = ~(1_n4710 ^ 1_n2313);
assign 1_n3195 = ~1_n4304;
assign 1_n9280 = ~1_n6333;
assign 1_n3675 = ~(1_n11082 | 1_n627);
assign 1_n10791 = ~(1_n451 ^ 1_n1680);
assign 1_n8806 = ~(1_n8650 | 1_n13023);
assign 1_n4323 = ~(1_n5203 | 1_n309);
assign 1_n4217 = 1_n6225 | 1_n12717;
assign 1_n2635 = ~(1_n11363 | 1_n10539);
assign 1_n371 = 1_n542 | 1_n12388;
assign 1_n10178 = ~1_n11169;
assign 1_n7087 = 1_n2264 | 1_n5242;
assign 1_n12088 = ~1_n13069;
assign 1_n5325 = ~(1_n2971 ^ 1_n6684);
assign 1_n8405 = 1_n2968 | 1_n4018;
assign 1_n3919 = 1_n3002 & 1_n11223;
assign 1_n13049 = 1_n4317 | 1_n11549;
assign 1_n4408 = ~(1_n7364 | 1_n219);
assign 1_n3487 = ~(1_n4994 ^ 1_n12305);
assign 1_n6689 = ~1_n3130;
assign 1_n1900 = 1_n1484 ^ 1_n9771;
assign 1_n6493 = 1_n12597 & 1_n9834;
assign 1_n13057 = ~(1_n11709 ^ 1_n3447);
assign 1_n5457 = 1_n7194 & 1_n7801;
assign 1_n8692 = ~(1_n11577 | 1_n9408);
assign 1_n9640 = ~(1_n9467 ^ 1_n13158);
assign 1_n4356 = 1_n10075 | 1_n7737;
assign 1_n7679 = 1_n7593 | 1_n2753;
assign 1_n7954 = 1_n10336 & 1_n6771;
assign 1_n11417 = ~(1_n7066 ^ 1_n9156);
assign 1_n9926 = 1_n9478 | 1_n479;
assign 1_n7718 = ~1_n9475;
assign 1_n1221 = ~(1_n6864 ^ 1_n7562);
assign 1_n13076 = 1_n12098 & 1_n11787;
assign 1_n9246 = ~(1_n7897 ^ 1_n889);
assign 1_n4265 = 1_n3178 & 1_n1007;
assign 1_n7641 = 1_n1649 & 1_n4263;
assign 1_n2622 = ~1_n5536;
assign 1_n42 = ~1_n3527;
assign 1_n8797 = ~(1_n8908 | 1_n8376);
assign 1_n7443 = ~1_n9839;
assign 1_n7766 = ~(1_n7380 ^ 1_n10156);
assign 1_n5862 = 1_n1888 | 1_n3224;
assign 1_n8243 = ~1_n12809;
assign 1_n1314 = 1_n11651 | 1_n4505;
assign 1_n9922 = ~(1_n3659 ^ 1_n7053);
assign 1_n6423 = 1_n12496 | 1_n6093;
assign 1_n2305 = 1_n12266 | 1_n11625;
assign 1_n151 = 1_n9193 | 1_n12287;
assign 1_n2447 = 1_n9358 ^ 1_n3720;
assign 1_n5421 = ~(1_n992 ^ 1_n12319);
assign 1_n10539 = 1_n12652 & 1_n12699;
assign 1_n10787 = ~(1_n1326 ^ 1_n11406);
assign 1_n11000 = 1_n4784 & 1_n4493;
assign 1_n5288 = ~(1_n5403 ^ 1_n9800);
assign 1_n9889 = ~1_n13078;
assign 1_n465 = ~(1_n2903 ^ 1_n10922);
assign 1_n254 = 1_n9926 | 1_n5175;
assign 1_n8422 = ~(1_n12117 ^ 1_n12594);
assign 1_n5892 = 1_n7661 | 1_n4936;
assign 1_n8464 = 1_n6223 | 1_n10871;
assign 1_n13179 = ~(1_n5881 ^ 1_n8281);
assign 1_n483 = ~(1_n12826 ^ 1_n5761);
assign 1_n3351 = ~(1_n1592 ^ 1_n3850);
assign 1_n6930 = ~(1_n8230 ^ 1_n6668);
assign 1_n1631 = 1_n5541 | 1_n6234;
assign 1_n1686 = 1_n7871 & 1_n6975;
assign 1_n5025 = 1_n3564 | 1_n11107;
assign 1_n4009 = ~(1_n10906 ^ 1_n9905);
assign 1_n8307 = 1_n13144 | 1_n6905;
assign 1_n3375 = ~(1_n10765 ^ 1_n6662);
assign 1_n10501 = ~1_n7720;
assign 1_n344 = 1_n2877 | 1_n12388;
assign 1_n4030 = ~1_n1288;
assign 1_n5638 = ~1_n4671;
assign 1_n261 = ~(1_n9222 ^ 1_n1348);
assign 1_n9015 = 1_n1262 | 1_n2986;
assign 1_n7376 = ~(1_n6611 ^ 1_n3605);
assign 1_n2838 = ~1_n4186;
assign 1_n3164 = 1_n1872 | 1_n11995;
assign 1_n4216 = 1_n1480 | 1_n902;
assign 1_n13017 = ~1_n12228;
assign 1_n13136 = ~(1_n2749 | 1_n10515);
assign 1_n11378 = 1_n1930 | 1_n8268;
assign 1_n13188 = ~(1_n5428 ^ 1_n9774);
assign 1_n33 = ~(1_n6395 ^ 1_n7148);
assign 1_n6330 = ~1_n11544;
assign 1_n1080 = ~1_n9918;
assign 1_n12063 = 1_n137 | 1_n4636;
assign 1_n3711 = ~(1_n503 ^ 1_n9820);
assign 1_n2623 = ~1_n3178;
assign 1_n7796 = ~(1_n1033 | 1_n4127);
assign 1_n7136 = ~(1_n3993 | 1_n2007);
assign 1_n5164 = 1_n2657 | 1_n3949;
assign 1_n5197 = 1_n4484 & 1_n11540;
assign 1_n211 = 1_n10680 ^ 1_n4121;
assign 1_n1135 = ~1_n9041;
assign 1_n2217 = ~1_n1231;
assign 1_n11456 = ~(1_n4954 | 1_n8162);
assign 1_n3170 = ~(1_n10855 ^ 1_n3547);
assign 1_n10568 = ~(1_n668 ^ 1_n2543);
assign 1_n518 = 1_n3908 | 1_n4640;
assign 1_n7062 = ~1_n7374;
assign 1_n8764 = 1_n5660 | 1_n2319;
assign 1_n5279 = ~1_n7514;
assign 1_n9127 = ~(1_n8060 ^ 1_n10169);
assign 1_n11386 = 1_n8729 | 1_n4640;
assign 1_n2823 = 1_n11941 | 1_n2133;
assign 1_n3360 = 1_n10383 | 1_n4724;
assign 1_n291 = ~(1_n7105 ^ 1_n13009);
assign 1_n12353 = 1_n7718 | 1_n4947;
assign 1_n9449 = ~(1_n11289 ^ 1_n13114);
assign 1_n12288 = 1_n9496 | 1_n8034;
assign 1_n11694 = ~(1_n6965 ^ 1_n2488);
assign 1_n9774 = ~(1_n1828 ^ 1_n4403);
assign 1_n10115 = ~(1_n2643 | 1_n4629);
assign 1_n6902 = 1_n3035 & 1_n8590;
assign 1_n10490 = 1_n9131 | 1_n1144;
assign 1_n4188 = 1_n9849 ^ 1_n11866;
assign 1_n9844 = ~(1_n7594 ^ 1_n7512);
assign 1_n6245 = ~1_n4419;
assign 1_n3838 = ~(1_n4291 ^ 1_n2256);
assign 1_n333 = ~1_n11488;
assign 1_n6862 = ~(1_n12051 ^ 1_n7663);
assign 1_n11463 = 1_n12293 | 1_n2044;
assign 1_n13140 = 1_n4339 | 1_n170;
assign 1_n4273 = ~(1_n3535 ^ 1_n393);
assign 1_n11905 = 1_n8385 & 1_n12431;
assign 1_n184 = ~(1_n13197 ^ 1_n8945);
assign 1_n7288 = ~(1_n3933 ^ 1_n10669);
assign 1_n8048 = 1_n2657 | 1_n3149;
assign 1_n6041 = ~1_n11537;
assign 1_n7675 = ~1_n7411;
assign 1_n12717 = ~1_n2590;
assign 1_n3015 = ~(1_n11744 ^ 1_n4235);
assign 1_n4822 = 1_n8113 | 1_n7032;
assign 1_n12392 = 1_n12441 | 1_n6814;
assign 1_n8741 = 1_n8420 | 1_n1866;
assign 1_n12084 = ~(1_n11508 ^ 1_n6623);
assign 1_n12091 = ~(1_n7829 ^ 1_n5532);
assign 1_n3735 = ~(1_n781 ^ 1_n4582);
assign 1_n8569 = ~1_n1757;
assign 1_n6208 = ~(1_n9243 | 1_n2245);
assign 1_n3754 = ~(1_n12484 ^ 1_n1957);
assign 1_n4867 = ~(1_n5539 ^ 1_n12444);
assign 1_n3072 = ~(1_n3389 ^ 1_n9374);
assign 1_n11097 = 1_n4835 & 1_n12236;
assign 1_n12269 = ~(1_n4396 ^ 1_n8612);
assign 1_n1949 = 1_n4754 & 1_n3533;
assign 1_n7566 = 1_n8561 | 1_n10871;
assign 1_n8899 = 1_n13130 | 1_n8828;
assign 1_n3120 = 1_n8158 | 1_n11719;
assign 1_n4517 = ~1_n10113;
assign 1_n10702 = ~(1_n968 ^ 1_n2923);
assign 1_n3900 = 1_n2892 & 1_n108;
assign 1_n8985 = ~1_n160;
assign 1_n10890 = ~1_n9324;
assign 1_n10873 = 1_n13122 & 1_n11813;
assign 1_n6501 = 1_n7327 | 1_n11841;
assign 1_n8669 = ~1_n3187;
assign 1_n8257 = 1_n10313 | 1_n1782;
assign 1_n5591 = ~(1_n2750 ^ 1_n8824);
assign 1_n5576 = ~(1_n2238 ^ 1_n12248);
assign 1_n3712 = ~1_n3973;
assign 1_n10483 = 1_n5527 & 1_n3831;
assign 1_n8102 = 1_n10668 & 1_n5141;
assign 1_n1596 = 1_n7427 | 1_n7534;
assign 1_n11925 = 1_n7159 & 1_n4928;
assign 1_n8744 = ~1_n8139;
assign 1_n8966 = ~(1_n2534 ^ 1_n11467);
assign 1_n9715 = 1_n10891 & 1_n5653;
assign 1_n10967 = 1_n7960 & 1_n12819;
assign 1_n3920 = 1_n8845 & 1_n7414;
assign 1_n9200 = ~(1_n9967 | 1_n1442);
assign 1_n10226 = ~(1_n7937 | 1_n7721);
assign 1_n5527 = ~1_n912;
assign 1_n8175 = ~1_n6083;
assign 1_n5323 = 1_n5713 | 1_n10029;
assign 1_n5310 = ~1_n13047;
assign 1_n7178 = ~(1_n9701 ^ 1_n7009);
assign 1_n12868 = 1_n5044 | 1_n12860;
assign 1_n2510 = 1_n3493 & 1_n1085;
assign 1_n2294 = ~1_n3005;
assign 1_n12858 = ~1_n4350;
endmodule
