.INIT_D0({INIT[15*4+0], INIT[14*4+0], INIT[13*4+0], INIT[12*4+0],
	  INIT[11*4+0], INIT[10*4+0], INIT[9*4+0], INIT[8*4+0],
	  INIT[7*4+0], INIT[6*4+0], INIT[5*4+0], INIT[4*4+0],
	  INIT[3*4+0], INIT[2*4+0], INIT[1*4+0], INIT[0*4+0]}),
.INIT_D1({INIT[15*4+1], INIT[14*4+1], INIT[13*4+1], INIT[12*4+1],
	  INIT[11*4+1], INIT[10*4+1], INIT[9*4+1], INIT[8*4+1],
	  INIT[7*4+1], INIT[6*4+1], INIT[5*4+1], INIT[4*4+1],
	  INIT[3*4+1], INIT[2*4+1], INIT[1*4+1], INIT[0*4+1]}),
.INIT_D2({INIT[15*4+2], INIT[14*4+2], INIT[13*4+2], INIT[12*4+2],
	  INIT[11*4+2], INIT[10*4+2], INIT[9*4+2], INIT[8*4+2],
	  INIT[7*4+2], INIT[6*4+2], INIT[5*4+2], INIT[4*4+2],
	  INIT[3*4+2], INIT[2*4+2], INIT[1*4+2], INIT[0*4+2]}),
.INIT_D3({INIT[15*4+3], INIT[14*4+3], INIT[13*4+3], INIT[12*4+3],
	  INIT[11*4+3], INIT[10*4+3], INIT[9*4+3], INIT[8*4+3],
	  INIT[7*4+3], INIT[6*4+3], INIT[5*4+3], INIT[4*4+3],
	  INIT[3*4+3], INIT[2*4+3], INIT[1*4+3], INIT[0*4+3]})
