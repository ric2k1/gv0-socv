module top( 1_n2 , 1_n11 , 1_n13 , 1_n16 , 1_n21 , 1_n44 , 1_n45 , 1_n46 , 1_n55 , 1_n74 , 1_n75 , 1_n81 , 1_n84 , 1_n85 , 1_n87 , 1_n93 , 1_n96 , 1_n98 , 1_n101 , 1_n105 , 1_n111 , 1_n123 , 1_n128 , 1_n131 , 1_n134 , 1_n139 , 1_n148 , 1_n153 , 1_n159 , 1_n163 , 1_n177 , 1_n191 , 1_n196 , 1_n199 , 1_n206 , 1_n211 , 1_n216 , 1_n223 , 1_n226 , 1_n240 , 1_n243 , 1_n254 , 1_n260 , 1_n264 , 1_n266 , 1_n280 , 1_n282 , 1_n283 , 1_n287 , 1_n290 , 1_n291 , 1_n299 , 1_n309 , 1_n336 , 1_n346 , 1_n349 , 1_n360 , 1_n368 , 1_n369 , 1_n377 , 1_n388 , 1_n394 , 1_n409 , 1_n428 , 1_n435 , 1_n442 , 1_n447 , 1_n449 , 1_n454 , 1_n457 , 1_n468 , 1_n471 , 1_n481 , 1_n484 , 1_n494 , 1_n500 , 1_n507 , 1_n511 , 1_n518 , 1_n519 , 1_n525 , 1_n534 , 1_n542 , 1_n547 , 1_n557 , 1_n561 , 1_n568 , 1_n569 , 1_n571 , 1_n575 , 1_n581 , 1_n582 , 1_n583 , 1_n587 , 1_n600 , 1_n603 , 1_n609 , 1_n613 , 1_n614 , 1_n616 , 1_n627 , 1_n635 , 1_n646 , 1_n659 , 1_n661 , 1_n664 , 1_n672 , 1_n673 );
    input 1_n2 , 1_n11 , 1_n13 , 1_n16 , 1_n21 , 1_n45 , 1_n46 , 1_n55 , 1_n74 , 1_n75 , 1_n81 , 1_n84 , 1_n85 , 1_n93 , 1_n96 , 1_n98 , 1_n101 , 1_n111 , 1_n128 , 1_n131 , 1_n134 , 1_n139 , 1_n153 , 1_n159 , 1_n177 , 1_n199 , 1_n206 , 1_n211 , 1_n216 , 1_n223 , 1_n243 , 1_n264 , 1_n266 , 1_n280 , 1_n282 , 1_n287 , 1_n290 , 1_n309 , 1_n336 , 1_n346 , 1_n349 , 1_n360 , 1_n368 , 1_n369 , 1_n377 , 1_n388 , 1_n394 , 1_n409 , 1_n428 , 1_n435 , 1_n447 , 1_n454 , 1_n457 , 1_n468 , 1_n471 , 1_n481 , 1_n494 , 1_n500 , 1_n507 , 1_n511 , 1_n519 , 1_n525 , 1_n557 , 1_n561 , 1_n569 , 1_n571 , 1_n575 , 1_n581 , 1_n582 , 1_n583 , 1_n587 , 1_n600 , 1_n603 , 1_n609 , 1_n613 , 1_n614 , 1_n616 , 1_n646 , 1_n659 , 1_n661 , 1_n664 , 1_n673 ;
    output 1_n44 , 1_n87 , 1_n105 , 1_n123 , 1_n148 , 1_n163 , 1_n191 , 1_n196 , 1_n226 , 1_n240 , 1_n254 , 1_n260 , 1_n283 , 1_n291 , 1_n299 , 1_n442 , 1_n449 , 1_n484 , 1_n518 , 1_n534 , 1_n542 , 1_n547 , 1_n568 , 1_n627 , 1_n635 , 1_n672 ;
    wire 1_n0 , 1_n1 , 1_n3 , 1_n4 , 1_n5 , 1_n6 , 1_n7 , 1_n8 , 1_n9 , 1_n10 , 1_n12 , 1_n14 , 1_n15 , 1_n17 , 1_n18 , 1_n19 , 1_n20 , 1_n22 , 1_n23 , 1_n24 , 1_n25 , 1_n26 , 1_n27 , 1_n28 , 1_n29 , 1_n30 , 1_n31 , 1_n32 , 1_n33 , 1_n34 , 1_n35 , 1_n36 , 1_n37 , 1_n38 , 1_n39 , 1_n40 , 1_n41 , 1_n42 , 1_n43 , 1_n47 , 1_n48 , 1_n49 , 1_n50 , 1_n51 , 1_n52 , 1_n53 , 1_n54 , 1_n56 , 1_n57 , 1_n58 , 1_n59 , 1_n60 , 1_n61 , 1_n62 , 1_n63 , 1_n64 , 1_n65 , 1_n66 , 1_n67 , 1_n68 , 1_n69 , 1_n70 , 1_n71 , 1_n72 , 1_n73 , 1_n76 , 1_n77 , 1_n78 , 1_n79 , 1_n80 , 1_n82 , 1_n83 , 1_n86 , 1_n88 , 1_n89 , 1_n90 , 1_n91 , 1_n92 , 1_n94 , 1_n95 , 1_n97 , 1_n99 , 1_n100 , 1_n102 , 1_n103 , 1_n104 , 1_n106 , 1_n107 , 1_n108 , 1_n109 , 1_n110 , 1_n112 , 1_n113 , 1_n114 , 1_n115 , 1_n116 , 1_n117 , 1_n118 , 1_n119 , 1_n120 , 1_n121 , 1_n122 , 1_n124 , 1_n125 , 1_n126 , 1_n127 , 1_n129 , 1_n130 , 1_n132 , 1_n133 , 1_n135 , 1_n136 , 1_n137 , 1_n138 , 1_n140 , 1_n141 , 1_n142 , 1_n143 , 1_n144 , 1_n145 , 1_n146 , 1_n147 , 1_n149 , 1_n150 , 1_n151 , 1_n152 , 1_n154 , 1_n155 , 1_n156 , 1_n157 , 1_n158 , 1_n160 , 1_n161 , 1_n162 , 1_n164 , 1_n165 , 1_n166 , 1_n167 , 1_n168 , 1_n169 , 1_n170 , 1_n171 , 1_n172 , 1_n173 , 1_n174 , 1_n175 , 1_n176 , 1_n178 , 1_n179 , 1_n180 , 1_n181 , 1_n182 , 1_n183 , 1_n184 , 1_n185 , 1_n186 , 1_n187 , 1_n188 , 1_n189 , 1_n190 , 1_n192 , 1_n193 , 1_n194 , 1_n195 , 1_n197 , 1_n198 , 1_n200 , 1_n201 , 1_n202 , 1_n203 , 1_n204 , 1_n205 , 1_n207 , 1_n208 , 1_n209 , 1_n210 , 1_n212 , 1_n213 , 1_n214 , 1_n215 , 1_n217 , 1_n218 , 1_n219 , 1_n220 , 1_n221 , 1_n222 , 1_n224 , 1_n225 , 1_n227 , 1_n228 , 1_n229 , 1_n230 , 1_n231 , 1_n232 , 1_n233 , 1_n234 , 1_n235 , 1_n236 , 1_n237 , 1_n238 , 1_n239 , 1_n241 , 1_n242 , 1_n244 , 1_n245 , 1_n246 , 1_n247 , 1_n248 , 1_n249 , 1_n250 , 1_n251 , 1_n252 , 1_n253 , 1_n255 , 1_n256 , 1_n257 , 1_n258 , 1_n259 , 1_n261 , 1_n262 , 1_n263 , 1_n265 , 1_n267 , 1_n268 , 1_n269 , 1_n270 , 1_n271 , 1_n272 , 1_n273 , 1_n274 , 1_n275 , 1_n276 , 1_n277 , 1_n278 , 1_n279 , 1_n281 , 1_n284 , 1_n285 , 1_n286 , 1_n288 , 1_n289 , 1_n292 , 1_n293 , 1_n294 , 1_n295 , 1_n296 , 1_n297 , 1_n298 , 1_n300 , 1_n301 , 1_n302 , 1_n303 , 1_n304 , 1_n305 , 1_n306 , 1_n307 , 1_n308 , 1_n310 , 1_n311 , 1_n312 , 1_n313 , 1_n314 , 1_n315 , 1_n316 , 1_n317 , 1_n318 , 1_n319 , 1_n320 , 1_n321 , 1_n322 , 1_n323 , 1_n324 , 1_n325 , 1_n326 , 1_n327 , 1_n328 , 1_n329 , 1_n330 , 1_n331 , 1_n332 , 1_n333 , 1_n334 , 1_n335 , 1_n337 , 1_n338 , 1_n339 , 1_n340 , 1_n341 , 1_n342 , 1_n343 , 1_n344 , 1_n345 , 1_n347 , 1_n348 , 1_n350 , 1_n351 , 1_n352 , 1_n353 , 1_n354 , 1_n355 , 1_n356 , 1_n357 , 1_n358 , 1_n359 , 1_n361 , 1_n362 , 1_n363 , 1_n364 , 1_n365 , 1_n366 , 1_n367 , 1_n370 , 1_n371 , 1_n372 , 1_n373 , 1_n374 , 1_n375 , 1_n376 , 1_n378 , 1_n379 , 1_n380 , 1_n381 , 1_n382 , 1_n383 , 1_n384 , 1_n385 , 1_n386 , 1_n387 , 1_n389 , 1_n390 , 1_n391 , 1_n392 , 1_n393 , 1_n395 , 1_n396 , 1_n397 , 1_n398 , 1_n399 , 1_n400 , 1_n401 , 1_n402 , 1_n403 , 1_n404 , 1_n405 , 1_n406 , 1_n407 , 1_n408 , 1_n410 , 1_n411 , 1_n412 , 1_n413 , 1_n414 , 1_n415 , 1_n416 , 1_n417 , 1_n418 , 1_n419 , 1_n420 , 1_n421 , 1_n422 , 1_n423 , 1_n424 , 1_n425 , 1_n426 , 1_n427 , 1_n429 , 1_n430 , 1_n431 , 1_n432 , 1_n433 , 1_n434 , 1_n436 , 1_n437 , 1_n438 , 1_n439 , 1_n440 , 1_n441 , 1_n443 , 1_n444 , 1_n445 , 1_n446 , 1_n448 , 1_n450 , 1_n451 , 1_n452 , 1_n453 , 1_n455 , 1_n456 , 1_n458 , 1_n459 , 1_n460 , 1_n461 , 1_n462 , 1_n463 , 1_n464 , 1_n465 , 1_n466 , 1_n467 , 1_n469 , 1_n470 , 1_n472 , 1_n473 , 1_n474 , 1_n475 , 1_n476 , 1_n477 , 1_n478 , 1_n479 , 1_n480 , 1_n482 , 1_n483 , 1_n485 , 1_n486 , 1_n487 , 1_n488 , 1_n489 , 1_n490 , 1_n491 , 1_n492 , 1_n493 , 1_n495 , 1_n496 , 1_n497 , 1_n498 , 1_n499 , 1_n501 , 1_n502 , 1_n503 , 1_n504 , 1_n505 , 1_n506 , 1_n508 , 1_n509 , 1_n510 , 1_n512 , 1_n513 , 1_n514 , 1_n515 , 1_n516 , 1_n517 , 1_n520 , 1_n521 , 1_n522 , 1_n523 , 1_n524 , 1_n526 , 1_n527 , 1_n528 , 1_n529 , 1_n530 , 1_n531 , 1_n532 , 1_n533 , 1_n535 , 1_n536 , 1_n537 , 1_n538 , 1_n539 , 1_n540 , 1_n541 , 1_n543 , 1_n544 , 1_n545 , 1_n546 , 1_n548 , 1_n549 , 1_n550 , 1_n551 , 1_n552 , 1_n553 , 1_n554 , 1_n555 , 1_n556 , 1_n558 , 1_n559 , 1_n560 , 1_n562 , 1_n563 , 1_n564 , 1_n565 , 1_n566 , 1_n567 , 1_n570 , 1_n572 , 1_n573 , 1_n574 , 1_n576 , 1_n577 , 1_n578 , 1_n579 , 1_n580 , 1_n584 , 1_n585 , 1_n586 , 1_n588 , 1_n589 , 1_n590 , 1_n591 , 1_n592 , 1_n593 , 1_n594 , 1_n595 , 1_n596 , 1_n597 , 1_n598 , 1_n599 , 1_n601 , 1_n602 , 1_n604 , 1_n605 , 1_n606 , 1_n607 , 1_n608 , 1_n610 , 1_n611 , 1_n612 , 1_n615 , 1_n617 , 1_n618 , 1_n619 , 1_n620 , 1_n621 , 1_n622 , 1_n623 , 1_n624 , 1_n625 , 1_n626 , 1_n628 , 1_n629 , 1_n630 , 1_n631 , 1_n632 , 1_n633 , 1_n634 , 1_n636 , 1_n637 , 1_n638 , 1_n639 , 1_n640 , 1_n641 , 1_n642 , 1_n643 , 1_n644 , 1_n645 , 1_n647 , 1_n648 , 1_n649 , 1_n650 , 1_n651 , 1_n652 , 1_n653 , 1_n654 , 1_n655 , 1_n656 , 1_n657 , 1_n658 , 1_n660 , 1_n662 , 1_n663 , 1_n665 , 1_n666 , 1_n667 , 1_n668 , 1_n669 , 1_n670 , 1_n671 ;
assign 1_n657 = 1_n356 & 1_n451;
assign 1_n203 = 1_n224 & 1_n349;
assign 1_n660 = 1_n340 & 1_n25;
assign 1_n347 = ~(1_n468 | 1_n417);
assign 1_n253 = ~1_n54;
assign 1_n6 = 1_n48 | 1_n383;
assign 1_n291 = ~(1_n339 ^ 1_n668);
assign 1_n308 = 1_n515 & 1_n168;
assign 1_n629 = 1_n253 | 1_n652;
assign 1_n187 = ~(1_n2 | 1_n159);
assign 1_n585 = ~1_n434;
assign 1_n570 = 1_n389;
assign 1_n47 = ~(1_n414 | 1_n467);
assign 1_n393 = ~(1_n444 ^ 1_n216);
assign 1_n391 = ~1_n531;
assign 1_n443 = ~1_n176;
assign 1_n76 = ~(1_n556 ^ 1_n16);
assign 1_n390 = ~(1_n598 ^ 1_n290);
assign 1_n38 = ~1_n499;
assign 1_n426 = 1_n524 | 1_n62;
assign 1_n117 = ~(1_n93 | 1_n396);
assign 1_n89 = 1_n9 & 1_n72;
assign 1_n628 = ~(1_n107 ^ 1_n531);
assign 1_n550 = ~1_n159;
assign 1_n365 = 1_n321 & 1_n253;
assign 1_n163 = ~(1_n0 ^ 1_n479);
assign 1_n61 = ~(1_n7 ^ 1_n613);
assign 1_n648 = 1_n127 & 1_n125;
assign 1_n283 = ~(1_n31 ^ 1_n648);
assign 1_n608 = ~1_n31;
assign 1_n327 = 1_n638 & 1_n367;
assign 1_n444 = 1_n285 | 1_n412;
assign 1_n373 = ~1_n639;
assign 1_n602 = 1_n570 & 1_n101;
assign 1_n251 = ~1_n75;
assign 1_n107 = ~1_n520;
assign 1_n427 = 1_n608 | 1_n125;
assign 1_n480 = ~(1_n349 | 1_n322);
assign 1_n359 = 1_n137 & 1_n604;
assign 1_n95 = ~(1_n13 | 1_n2);
assign 1_n118 = ~(1_n623 | 1_n540);
assign 1_n474 = ~1_n613;
assign 1_n115 = ~(1_n93 | 1_n37);
assign 1_n398 = ~1_n0;
assign 1_n289 = ~(1_n280 ^ 1_n287);
assign 1_n543 = 1_n390 & 1_n266;
assign 1_n60 = ~(1_n624 ^ 1_n464);
assign 1_n141 = 1_n538 | 1_n452;
assign 1_n572 = ~1_n466;
assign 1_n339 = 1_n5 | 1_n492;
assign 1_n31 = 1_n559 | 1_n424;
assign 1_n514 = ~1_n206;
assign 1_n234 = 1_n198 & 1_n326;
assign 1_n258 = 1_n19 & 1_n266;
assign 1_n300 = ~1_n428;
assign 1_n651 = 1_n526 & 1_n570;
assign 1_n197 = ~1_n138;
assign 1_n351 = ~1_n508;
assign 1_n649 = ~1_n225;
assign 1_n100 = 1_n413 | 1_n179;
assign 1_n670 = ~(1_n203 | 1_n611);
assign 1_n30 = 1_n318 | 1_n342;
assign 1_n144 = 1_n385 | 1_n445;
assign 1_n453 = 1_n539 | 1_n344;
assign 1_n78 = ~1_n365;
assign 1_n496 = 1_n233 & 1_n93;
assign 1_n179 = ~(1_n570 | 1_n330);
assign 1_n39 = ~(1_n490 | 1_n480);
assign 1_n149 = ~1_n144;
assign 1_n182 = ~(1_n183 | 1_n370);
assign 1_n9 = 1_n513 & 1_n551;
assign 1_n152 = ~(1_n356 ^ 1_n616);
assign 1_n576 = ~1_n100;
assign 1_n662 = 1_n580 & 1_n264;
assign 1_n123 = ~(1_n182 ^ 1_n463);
assign 1_n65 = 1_n201 | 1_n439;
assign 1_n259 = 1_n58 | 1_n1;
assign 1_n591 = ~(1_n590 | 1_n275);
assign 1_n200 = 1_n136 & 1_n266;
assign 1_n399 = ~1_n573;
assign 1_n558 = 1_n64 | 1_n453;
assign 1_n434 = 1_n450 | 1_n86;
assign 1_n618 = 1_n537 | 1_n18;
assign 1_n140 = 1_n333 & 1_n654;
assign 1_n553 = ~(1_n6 ^ 1_n432);
assign 1_n34 = 1_n375 | 1_n116;
assign 1_n5 = 1_n570 & 1_n500;
assign 1_n530 = ~(1_n472 | 1_n327);
assign 1_n626 = 1_n384 | 1_n642;
assign 1_n401 = ~(1_n582 ^ 1_n2);
assign 1_n450 = 1_n190 | 1_n307;
assign 1_n106 = 1_n465 & 1_n608;
assign 1_n40 = 1_n421 & 1_n93;
assign 1_n520 = ~1_n248;
assign 1_n299 = ~(1_n395 ^ 1_n175);
assign 1_n501 = ~1_n171;
assign 1_n420 = ~1_n45;
assign 1_n169 = 1_n319 | 1_n629;
assign 1_n637 = 1_n124 & 1_n335;
assign 1_n621 = ~1_n380;
assign 1_n267 = ~(1_n570 | 1_n140);
assign 1_n105 = ~(1_n54 ^ 1_n615);
assign 1_n533 = 1_n331 | 1_n52;
assign 1_n355 = 1_n71 | 1_n591;
assign 1_n260 = ~(1_n508 ^ 1_n669);
assign 1_n594 = 1_n514 | 1_n516;
assign 1_n395 = ~(1_n431 | 1_n663);
assign 1_n302 = ~(1_n453 ^ 1_n336);
assign 1_n363 = 1_n526 | 1_n239;
assign 1_n238 = 1_n42 & 1_n93;
assign 1_n424 = 1_n61 & 1_n266;
assign 1_n567 = 1_n77 & 1_n569;
assign 1_n79 = 1_n29 & 1_n266;
assign 1_n598 = 1_n298 | 1_n460;
assign 1_n620 = ~(1_n632 ^ 1_n392);
assign 1_n479 = ~(1_n185 | 1_n425);
assign 1_n143 = ~1_n339;
assign 1_n77 = 1_n389;
assign 1_n624 = 1_n285 | 1_n305;
assign 1_n218 = 1_n249 & 1_n266;
assign 1_n3 = 1_n147 & 1_n266;
assign 1_n88 = ~(1_n199 | 1_n85);
assign 1_n249 = ~(1_n426 ^ 1_n282);
assign 1_n380 = 1_n358 | 1_n597;
assign 1_n654 = 1_n58 | 1_n562;
assign 1_n165 = 1_n201 | 1_n660;
assign 1_n212 = ~(1_n75 | 1_n131);
assign 1_n623 = ~1_n577;
assign 1_n7 = 1_n636 | 1_n477;
assign 1_n340 = ~(1_n170 | 1_n418);
assign 1_n114 = 1_n482 | 1_n444;
assign 1_n560 = ~1_n209;
assign 1_n580 = 1_n666 & 1_n43;
assign 1_n274 = 1_n570 & 1_n603;
assign 1_n1 = ~1_n381;
assign 1_n484 = ~(1_n180 ^ 1_n584);
assign 1_n592 = 1_n606 | 1_n503;
assign 1_n222 = 1_n26 & 1_n436;
assign 1_n335 = 1_n397 | 1_n517;
assign 1_n461 = ~1_n13;
assign 1_n650 = ~(1_n665 | 1_n15);
assign 1_n552 = 1_n220 | 1_n461;
assign 1_n475 = 1_n227 | 1_n637;
assign 1_n386 = 1_n231 | 1_n323;
assign 1_n130 = 1_n440 | 1_n548;
assign 1_n312 = ~(1_n77 | 1_n637);
assign 1_n463 = 1_n566 | 1_n543;
assign 1_n497 = 1_n538 | 1_n278;
assign 1_n655 = 1_n470 | 1_n324;
assign 1_n257 = 1_n387 | 1_n200;
assign 1_n110 = 1_n65 & 1_n601;
assign 1_n478 = 1_n570 & 1_n153;
assign 1_n90 = 1_n653 | 1_n459;
assign 1_n658 = 1_n302 & 1_n266;
assign 1_n262 = ~(1_n177 ^ 1_n75);
assign 1_n155 = ~1_n521;
assign 1_n383 = ~1_n468;
assign 1_n167 = 1_n359 | 1_n219;
assign 1_n15 = ~1_n373;
assign 1_n247 = 1_n662 | 1_n404;
assign 1_n640 = 1_n284 & 1_n552;
assign 1_n201 = ~1_n352;
assign 1_n415 = ~(1_n194 | 1_n133);
assign 1_n367 = 1_n625 | 1_n209;
assign 1_n635 = ~(1_n12 ^ 1_n4);
assign 1_n207 = ~1_n641;
assign 1_n344 = 1_n429 | 1_n353;
assign 1_n192 = ~(1_n34 | 1_n517);
assign 1_n189 = 1_n235 & 1_n487;
assign 1_n261 = 1_n428 | 1_n48;
assign 1_n389 = ~1_n266;
assign 1_n148 = ~(1_n36 ^ 1_n17);
assign 1_n372 = 1_n57 & 1_n266;
assign 1_n579 = 1_n586 | 1_n78;
assign 1_n374 = 1_n393 & 1_n206;
assign 1_n124 = 1_n334 | 1_n140;
assign 1_n174 = ~1_n51;
assign 1_n4 = 1_n434 & 1_n52;
assign 1_n588 = ~1_n388;
assign 1_n269 = 1_n564 & 1_n126;
assign 1_n156 = 1_n63 | 1_n495;
assign 1_n286 = 1_n455 & 1_n482;
assign 1_n161 = ~(1_n657 | 1_n438);
assign 1_n483 = ~1_n6;
assign 1_n509 = ~1_n368;
assign 1_n541 = ~(1_n472 | 1_n39);
assign 1_n43 = ~1_n93;
assign 1_n64 = ~1_n336;
assign 1_n284 = 1_n95 | 1_n294;
assign 1_n328 = ~1_n631;
assign 1_n464 = ~(1_n511 ^ 1_n454);
assign 1_n433 = 1_n158 & 1_n441;
assign 1_n563 = ~1_n511;
assign 1_n71 = 1_n2 & 1_n582;
assign 1_n67 = 1_n94 & 1_n35;
assign 1_n456 = 1_n251 | 1_n8;
assign 1_n217 = ~(1_n135 | 1_n419);
assign 1_n448 = ~1_n595;
assign 1_n310 = ~1_n533;
assign 1_n265 = ~(1_n289 | 1_n316);
assign 1_n151 = 1_n286 | 1_n408;
assign 1_n281 = 1_n221 | 1_n593;
assign 1_n568 = ~(1_n217 ^ 1_n406);
assign 1_n644 = 1_n570 & 1_n614;
assign 1_n73 = ~1_n450;
assign 1_n154 = ~(1_n459 ^ 1_n583);
assign 1_n532 = 1_n475 & 1_n167;
assign 1_n607 = ~(1_n355 ^ 1_n97);
assign 1_n256 = 1_n553 & 1_n93;
assign 1_n150 = 1_n570 & 1_n519;
assign 1_n304 = ~(1_n107 | 1_n219);
assign 1_n80 = ~1_n352;
assign 1_n667 = 1_n639 & 1_n174;
assign 1_n248 = ~1_n359;
assign 1_n87 = ~(1_n156 ^ 1_n49);
assign 1_n168 = 1_n359 | 1_n271;
assign 1_n403 = 1_n451 | 1_n295;
assign 1_n324 = ~1_n560;
assign 1_n593 = 1_n546 & 1_n527;
assign 1_n215 = ~1_n235;
assign 1_n32 = 1_n659 & 1_n93;
assign 1_n458 = ~(1_n294 ^ 1_n112);
assign 1_n513 = 1_n187 | 1_n632;
assign 1_n467 = 1_n206 | 1_n509;
assign 1_n385 = 1_n237 | 1_n129;
assign 1_n72 = 1_n251 | 1_n121;
assign 1_n517 = ~1_n197;
assign 1_n8 = ~1_n177;
assign 1_n482 = ~1_n216;
assign 1_n337 = ~(1_n443 | 1_n269);
assign 1_n476 = 1_n650 | 1_n50;
assign 1_n638 = ~(1_n229 | 1_n265);
assign 1_n319 = ~1_n586;
assign 1_n157 = 1_n212 | 1_n89;
assign 1_n240 = ~(1_n341 ^ 1_n402);
assign 1_n24 = ~1_n491;
assign 1_n295 = 1_n493 | 1_n114;
assign 1_n627 = ~(1_n130 ^ 1_n366);
assign 1_n625 = ~1_n664;
assign 1_n178 = 1_n616 | 1_n66;
assign 1_n642 = 1_n505 | 1_n90;
assign 1_n311 = 1_n228 | 1_n363;
assign 1_n33 = ~(1_n620 | 1_n623);
assign 1_n18 = ~(1_n77 | 1_n60);
assign 1_n171 = 1_n351 | 1_n169;
assign 1_n341 = 1_n343 | 1_n345;
assign 1_n68 = 1_n570 & 1_n581;
assign 1_n556 = 1_n102 | 1_n329;
assign 1_n437 = ~(1_n119 | 1_n293);
assign 1_n606 = ~1_n646;
assign 1_n565 = ~1_n624;
assign 1_n412 = ~1_n454;
assign 1_n473 = ~1_n432;
assign 1_n462 = ~1_n381;
assign 1_n503 = 1_n315 | 1_n426;
assign 1_n48 = ~1_n409;
assign 1_n285 = ~1_n659;
assign 1_n27 = ~(1_n119 | 1_n356);
assign 1_n263 = ~(1_n626 ^ 1_n388);
assign 1_n430 = ~1_n579;
assign 1_n112 = ~(1_n13 ^ 1_n2);
assign 1_n536 = ~1_n561;
assign 1_n527 = 1_n478 | 1_n574;
assign 1_n358 = ~(1_n20 | 1_n43);
assign 1_n632 = 1_n276 | 1_n120;
assign 1_n505 = ~1_n55;
assign 1_n313 = 1_n386 & 1_n259;
assign 1_n104 = 1_n511 | 1_n659;
assign 1_n296 = ~(1_n435 | 1_n75);
assign 1_n146 = 1_n454 & 1_n511;
assign 1_n307 = 1_n272 & 1_n266;
assign 1_n321 = ~1_n656;
assign 1_n554 = ~1_n555;
assign 1_n276 = ~1_n287;
assign 1_n442 = ~(1_n172 ^ 1_n382);
assign 1_n619 = ~(1_n6 | 1_n473);
assign 1_n396 = 1_n165 & 1_n522;
assign 1_n566 = 1_n77 & 1_n74;
assign 1_n22 = ~1_n425;
assign 1_n120 = ~1_n96;
assign 1_n323 = ~(1_n306 | 1_n562);
assign 1_n224 = 1_n275 ^ 1_n401;
assign 1_n315 = ~1_n282;
assign 1_n23 = 1_n596 & 1_n155;
assign 1_n172 = 1_n274 | 1_n325;
assign 1_n306 = ~1_n576;
assign 1_n241 = 1_n506 | 1_n592;
assign 1_n528 = 1_n405 | 1_n427;
assign 1_n63 = 1_n570 & 1_n139;
assign 1_n183 = 1_n242 & 1_n555;
assign 1_n378 = ~(1_n292 | 1_n193);
assign 1_n20 = ~(1_n428 ^ 1_n454);
assign 1_n666 = ~(1_n80 | 1_n209);
assign 1_n669 = 1_n579 & 1_n169;
assign 1_n353 = 1_n634 | 1_n612;
assign 1_n126 = ~1_n350;
assign 1_n548 = 1_n622 & 1_n266;
assign 1_n42 = ~(1_n10 ^ 1_n202);
assign 1_n508 = 1_n166 | 1_n258;
assign 1_n488 = 1_n279 & 1_n77;
assign 1_n498 = ~(1_n423 ^ 1_n45);
assign 1_n116 = ~(1_n77 | 1_n76);
assign 1_n489 = 1_n437 | 1_n10;
assign 1_n37 = 1_n273 & 1_n594;
assign 1_n510 = ~1_n211;
assign 1_n278 = ~1_n38;
assign 1_n460 = 1_n230 | 1_n558;
assign 1_n226 = ~(1_n213 ^ 1_n245);
assign 1_n397 = ~1_n448;
assign 1_n559 = 1_n77 & 1_n609;
assign 1_n371 = 1_n77 & 1_n11;
assign 1_n405 = ~1_n172;
assign 1_n555 = 1_n486 | 1_n647;
assign 1_n268 = ~1_n629;
assign 1_n589 = 1_n106 & 1_n405;
assign 1_n205 = 1_n422 | 1_n241;
assign 1_n665 = ~1_n51;
assign 1_n421 = ~(1_n455 ^ 1_n103);
assign 1_n186 = 1_n580 & 1_n21;
assign 1_n417 = 1_n409 & 1_n428;
assign 1_n209 = 1_n85 | 1_n349;
assign 1_n293 = ~(1_n261 ^ 1_n468);
assign 1_n516 = ~(1_n214 ^ 1_n114);
assign 1_n135 = 1_n231 & 1_n77;
assign 1_n518 = ~(1_n555 ^ 1_n195);
assign 1_n633 = 1_n624 & 1_n104;
assign 1_n438 = 1_n489 & 1_n178;
assign 1_n663 = ~(1_n570 | 1_n532);
assign 1_n12 = 1_n602 | 1_n3;
assign 1_n82 = ~(1_n160 | 1_n312);
assign 1_n504 = ~(1_n296 | 1_n91);
assign 1_n250 = ~(1_n177 | 1_n75);
assign 1_n384 = ~1_n128;
assign 1_n142 = 1_n236 & 1_n497;
assign 1_n599 = ~1_n216;
assign 1_n645 = 1_n59 | 1_n228;
assign 1_n436 = 1_n485 | 1_n23;
assign 1_n564 = ~1_n132;
assign 1_n162 = ~(1_n514 | 1_n643);
assign 1_n108 = 1_n210 & 1_n85;
assign 1_n173 = 1_n317 & 1_n266;
assign 1_n596 = 1_n32 | 1_n332;
assign 1_n50 = ~(1_n667 | 1_n532);
assign 1_n230 = ~1_n494;
assign 1_n305 = ~1_n511;
assign 1_n298 = ~1_n223;
assign 1_n350 = 1_n68 | 1_n529;
assign 1_n160 = 1_n67 & 1_n77;
assign 1_n326 = 1_n599 | 1_n305;
assign 1_n366 = 1_n144 & 1_n184;
assign 1_n485 = ~1_n618;
assign 1_n577 = ~1_n467;
assign 1_n109 = ~1_n527;
assign 1_n522 = ~(1_n374 | 1_n118);
assign 1_n615 = 1_n656 & 1_n652;
assign 1_n537 = 1_n77 & 1_n46;
assign 1_n431 = 1_n308 & 1_n570;
assign 1_n254 = 1_n411 | 1_n281;
assign 1_n597 = ~(1_n93 | 1_n110);
assign 1_n147 = ~(1_n344 ^ 1_n369);
assign 1_n499 = 1_n40 | 1_n117;
assign 1_n121 = ~1_n131;
assign 1_n601 = ~(1_n33 | 1_n162);
assign 1_n127 = ~1_n465;
assign 1_n26 = 1_n380 | 1_n354;
assign 1_n17 = ~(1_n448 ^ 1_n138);
assign 1_n231 = 1_n181 & 1_n141;
assign 1_n198 = ~1_n288;
assign 1_n387 = 1_n570 & 1_n457;
assign 1_n653 = ~1_n583;
assign 1_n590 = ~(1_n582 | 1_n2);
assign 1_n361 = 1_n28 & 1_n53;
assign 1_n136 = ~(1_n288 ^ 1_n113);
assign 1_n652 = 1_n266 | 1_n415;
assign 1_n531 = 1_n186 | 1_n256;
assign 1_n166 = 1_n570 & 1_n571;
assign 1_n610 = ~1_n138;
assign 1_n297 = 1_n498 & 1_n266;
assign 1_n94 = 1_n192 | 1_n313;
assign 1_n145 = ~1_n130;
assign 1_n193 = 1_n47 | 1_n530;
assign 1_n232 = ~1_n377;
assign 1_n342 = 1_n145 | 1_n184;
assign 1_n138 = 1_n247 | 1_n496;
assign 1_n470 = ~1_n525;
assign 1_n213 = ~(1_n488 | 1_n362);
assign 1_n325 = 1_n154 & 1_n266;
assign 1_n382 = 1_n446 & 1_n427;
assign 1_n429 = ~1_n575;
assign 1_n538 = ~1_n207;
assign 1_n449 = ~(1_n155 ^ 1_n596);
assign 1_n418 = 1_n607 & 1_n349;
assign 1_n176 = 1_n126 | 1_n30;
assign 1_n605 = 1_n570 & 1_n84;
assign 1_n70 = 1_n143 | 1_n171;
assign 1_n370 = 1_n411 & 1_n554;
assign 1_n86 = ~1_n269;
assign 1_n119 = ~1_n616;
assign 1_n273 = ~(1_n502 | 1_n541);
assign 1_n441 = ~1_n239;
assign 1_n316 = 1_n349 | 1_n92;
assign 1_n630 = 1_n149 & 1_n145;
assign 1_n294 = 1_n276 | 1_n545;
assign 1_n318 = ~1_n341;
assign 1_n219 = ~1_n391;
assign 1_n604 = 1_n266 | 1_n232;
assign 1_n402 = ~(1_n416 | 1_n630);
assign 1_n672 = ~(1_n385 ^ 1_n400);
assign 1_n208 = ~1_n528;
assign 1_n272 = ~(1_n353 ^ 1_n575);
assign 1_n320 = ~1_n600;
assign 1_n376 = ~(1_n511 ^ 1_n616);
assign 1_n52 = 1_n73 | 1_n176;
assign 1_n314 = ~1_n109;
assign 1_n92 = ~1_n85;
assign 1_n611 = ~(1_n458 | 1_n316);
assign 1_n181 = 1_n122 | 1_n279;
assign 1_n53 = ~1_n180;
assign 1_n338 = 1_n75 & 1_n435;
assign 1_n245 = ~(1_n207 ^ 1_n499);
assign 1_n244 = ~(1_n558 ^ 1_n494);
assign 1_n521 = ~1_n526;
assign 1_n14 = ~1_n23;
assign 1_n540 = ~(1_n9 ^ 1_n164);
assign 1_n574 = 1_n244 & 1_n266;
assign 1_n303 = 1_n77 & 1_n346;
assign 1_n132 = 1_n341 | 1_n56;
assign 1_n422 = ~1_n557;
assign 1_n529 = 1_n469 & 1_n266;
assign 1_n671 = 1_n313 & 1_n77;
assign 1_n419 = ~(1_n77 | 1_n142);
assign 1_n354 = ~(1_n618 | 1_n14);
assign 1_n255 = 1_n563 | 1_n348;
assign 1_n221 = ~(1_n527 | 1_n225);
assign 1_n54 = 1_n605 | 1_n79;
assign 1_n102 = ~(1_n563 | 1_n214);
assign 1_n25 = 1_n510 | 1_n324;
assign 1_n204 = ~(1_n257 | 1_n452);
assign 1_n362 = ~(1_n570 | 1_n222);
assign 1_n636 = ~1_n471;
assign 1_n252 = 1_n599 | 1_n455;
assign 1_n356 = 1_n483 | 1_n347;
assign 1_n524 = ~1_n111;
assign 1_n413 = 1_n77 & 1_n507;
assign 1_n292 = ~(1_n659 | 1_n493);
assign 1_n357 = ~(1_n241 ^ 1_n557);
assign 1_n133 = ~(1_n99 | 1_n308);
assign 1_n647 = 1_n410 & 1_n266;
assign 1_n639 = 1_n277 | 1_n549;
assign 1_n495 = 1_n357 & 1_n266;
assign 1_n36 = ~(1_n671 | 1_n267);
assign 1_n329 = ~1_n234;
assign 1_n35 = 1_n397 | 1_n610;
assign 1_n526 = 1_n24 & 1_n270;
assign 1_n0 = 1_n303 | 1_n173;
assign 1_n379 = ~1_n156;
assign 1_n586 = 1_n371 | 1_n218;
assign 1_n28 = 1_n585 & 1_n331;
assign 1_n57 = ~(1_n477 ^ 1_n471);
assign 1_n472 = 1_n368 | 1_n206;
assign 1_n180 = 1_n567 | 1_n658;
assign 1_n535 = ~(1_n90 ^ 1_n55);
assign 1_n656 = 1_n77 | 1_n476;
assign 1_n91 = ~(1_n338 | 1_n355);
assign 1_n44 = ~(1_n466 ^ 1_n189);
assign 1_n41 = ~1_n16;
assign 1_n381 = 1_n238 | 1_n115;
assign 1_n56 = ~1_n630;
assign 1_n451 = ~1_n616;
assign 1_n99 = 1_n373 & 1_n174;
assign 1_n348 = ~1_n423;
assign 1_n322 = 1_n88 | 1_n108;
assign 1_n233 = ~(1_n438 ^ 1_n152);
assign 1_n220 = ~1_n2;
assign 1_n506 = ~1_n243;
assign 1_n235 = 1_n0 | 1_n22;
assign 1_n184 = 1_n69 | 1_n528;
assign 1_n539 = ~1_n369;
assign 1_n270 = 1_n266 | 1_n83;
assign 1_n551 = 1_n220 | 1_n550;
assign 1_n188 = ~(1_n268 | 1_n365);
assign 1_n465 = 1_n215 & 1_n572;
assign 1_n410 = ~(1_n460 ^ 1_n223);
assign 1_n195 = ~(1_n242 | 1_n411);
assign 1_n122 = ~(1_n257 | 1_n278);
assign 1_n288 = 1_n146 | 1_n565;
assign 1_n408 = ~(1_n428 ^ 1_n409);
assign 1_n49 = 1_n573 & 1_n70;
assign 1_n578 = 1_n640 & 1_n456;
assign 1_n547 = ~(1_n82 ^ 1_n628);
assign 1_n493 = ~1_n206;
assign 1_n331 = ~1_n12;
assign 1_n400 = ~(1_n208 | 1_n589);
assign 1_n66 = ~1_n293;
assign 1_n51 = 1_n150 | 1_n297;
assign 1_n631 = 1_n430 & 1_n351;
assign 1_n214 = ~1_n616;
assign 1_n236 = 1_n204 | 1_n222;
assign 1_n343 = 1_n77 & 1_n360;
assign 1_n668 = ~(1_n501 | 1_n631);
assign 1_n137 = 1_n77 | 1_n255;
assign 1_n406 = ~(1_n306 ^ 1_n381);
assign 1_n185 = ~1_n544;
assign 1_n641 = ~1_n257;
assign 1_n62 = 1_n420 | 1_n423;
assign 1_n246 = ~(1_n640 ^ 1_n262);
assign 1_n229 = 1_n364 & 1_n349;
assign 1_n59 = 1_n491 | 1_n651;
assign 1_n271 = ~1_n531;
assign 1_n227 = ~(1_n248 | 1_n271);
assign 1_n158 = 1_n407 | 1_n621;
assign 1_n242 = 1_n649 & 1_n314;
assign 1_n277 = 1_n580 & 1_n98;
assign 1_n29 = ~(1_n62 ^ 1_n111);
assign 1_n190 = 1_n570 & 1_n134;
assign 1_n491 = 1_n633 & 1_n266;
assign 1_n549 = 1_n619 & 1_n93;
assign 1_n634 = ~1_n661;
assign 1_n333 = 1_n617 | 1_n142;
assign 1_n202 = ~(1_n293 ^ 1_n616);
assign 1_n196 = ~(1_n645 ^ 1_n433);
assign 1_n58 = ~1_n100;
assign 1_n459 = 1_n474 | 1_n7;
assign 1_n364 = 1_n600 ^ 1_n287;
assign 1_n622 = ~(1_n642 ^ 1_n128);
assign 1_n643 = ~(1_n659 ^ 1_n454);
assign 1_n486 = 1_n77 & 1_n309;
assign 1_n515 = 1_n304 | 1_n67;
assign 1_n414 = ~(1_n287 ^ 1_n96);
assign 1_n194 = 1_n15 & 1_n51;
assign 1_n490 = 1_n504 & 1_n349;
assign 1_n584 = ~(1_n310 | 1_n28);
assign 1_n446 = ~1_n106;
assign 1_n191 = ~(1_n350 ^ 1_n523);
assign 1_n125 = 1_n572 | 1_n487;
assign 1_n103 = ~(1_n408 ^ 1_n216);
assign 1_n469 = ~(1_n612 ^ 1_n661);
assign 1_n228 = ~1_n596;
assign 1_n332 = ~(1_n93 | 1_n378);
assign 1_n502 = ~(1_n467 | 1_n157);
assign 1_n10 = 1_n151 & 1_n252;
assign 1_n512 = ~1_n556;
assign 1_n237 = 1_n570 & 1_n447;
assign 1_n573 = 1_n339 | 1_n328;
assign 1_n164 = ~(1_n75 ^ 1_n131);
assign 1_n69 = ~1_n385;
assign 1_n225 = 1_n53 | 1_n533;
assign 1_n239 = 1_n621 & 1_n407;
assign 1_n466 = 1_n644 | 1_n372;
assign 1_n407 = ~1_n618;
assign 1_n523 = 1_n132 & 1_n30;
assign 1_n175 = 1_n99 | 1_n194;
assign 1_n440 = 1_n570 & 1_n394;
assign 1_n544 = 1_n379 | 1_n70;
assign 1_n487 = 1_n398 | 1_n544;
assign 1_n545 = ~1_n280;
assign 1_n534 = ~(1_n586 ^ 1_n188);
assign 1_n210 = 1_n250 | 1_n578;
assign 1_n542 = ~(1_n450 ^ 1_n337);
assign 1_n279 = 1_n311 & 1_n158;
assign 1_n275 = 1_n276 | 1_n320;
assign 1_n330 = ~(1_n234 ^ 1_n376);
assign 1_n416 = ~1_n342;
assign 1_n546 = ~(1_n649 | 1_n361);
assign 1_n477 = 1_n536 | 1_n205;
assign 1_n411 = 1_n361 & 1_n109;
assign 1_n352 = ~1_n472;
assign 1_n612 = 1_n588 | 1_n626;
assign 1_n452 = ~1_n499;
assign 1_n423 = 1_n41 | 1_n512;
assign 1_n375 = 1_n77 & 1_n81;
assign 1_n492 = 1_n301 & 1_n266;
assign 1_n392 = ~(1_n2 ^ 1_n159);
assign 1_n129 = 1_n535 & 1_n266;
assign 1_n562 = ~1_n462;
assign 1_n334 = ~(1_n34 | 1_n610);
assign 1_n113 = ~(1_n511 ^ 1_n216);
assign 1_n439 = 1_n670 & 1_n655;
assign 1_n455 = 1_n300 | 1_n412;
assign 1_n345 = 1_n263 & 1_n266;
assign 1_n617 = ~(1_n100 | 1_n1);
assign 1_n97 = ~(1_n435 ^ 1_n75);
assign 1_n425 = 1_n399 & 1_n379;
assign 1_n432 = 1_n27 | 1_n161;
assign 1_n301 = ~(1_n592 ^ 1_n243);
assign 1_n445 = ~1_n589;
assign 1_n317 = ~(1_n205 ^ 1_n561);
assign 1_n19 = ~(1_n503 ^ 1_n646);
assign 1_n595 = ~1_n34;
assign 1_n404 = ~(1_n93 | 1_n403);
assign 1_n170 = ~(1_n316 | 1_n246);
assign 1_n83 = ~1_n673;
endmodule
