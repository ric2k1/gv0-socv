module a;
parameter integer real x=0;
endmodule
