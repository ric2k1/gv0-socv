module top( n0 , n3 , n4 , n10 , n11 , n15 , n21 , n33 , n35 , n36 , n37 , n39 , n41 , n61 , n66 , n70 , n71 , n73 , n79 , n80 );
    input n0 , n3 , n11 , n15 , n21 , n35 , n36 , n37 , n41 , n61 , n73 , n80 ;
    output n4 , n10 , n33 , n39 , n66 , n70 , n71 , n79 ;
    wire n1 , n2 , n5 , n6 , n7 , n8 , n9 , n12 , n13 , n14 , n16 , n17 , n18 , n19 , n20 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n34 , n38 , n40 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n62 , n63 , n64 , n65 , n67 , n68 , n69 , n72 , n74 , n75 , n76 , n77 , n78 , n81 , n82 , n83 ;
assign n72 = ~n74;
assign n76 = ~(n3 | n21);
assign n53 = ~(n73 | n34);
assign n58 = n31 & n19;
assign n19 = ~n36;
assign n67 = n18 & n43;
assign n59 = n69 | n50;
assign n66 = ~(n77 ^ n20);
assign n32 = n13 | n28;
assign n60 = n66 & n70;
assign n10 = ~(n33 & n71);
assign n47 = ~n15;
assign n29 = n65 | n24;
assign n48 = ~n80;
assign n16 = n46 | n42;
assign n44 = n72 | n55;
assign n22 = n68 | n53;
assign n64 = ~(n0 | n21);
assign n43 = n78 | n48;
assign n9 = n39 & n60;
assign n79 = n4 & n9;
assign n17 = n59 & n58;
assign n81 = n64 | n63;
assign n52 = ~(n44 | n5);
assign n40 = ~(n72 | n58);
assign n83 = ~n11;
assign n46 = n67 & n47;
assign n6 = ~n3;
assign n69 = ~n37;
assign n8 = ~n41;
assign n68 = ~(n61 | n21);
assign n55 = ~n59;
assign n74 = n19 | n22;
assign n39 = ~(n16 ^ n40);
assign n49 = n59 & n75;
assign n25 = ~(n17 | n52);
assign n56 = n58 | n51;
assign n26 = n34 | n48;
assign n13 = ~n77;
assign n57 = ~n41;
assign n77 = n83 | n29;
assign n34 = ~n61;
assign n5 = ~(n46 | n82);
assign n65 = ~(n35 | n21);
assign n24 = ~(n73 | n45);
assign n20 = ~(n28 | n46);
assign n31 = n7 & n26;
assign n70 = n77 & n12;
assign n1 = n14 & n27;
assign n38 = n62 | n54;
assign n75 = n37 | n38;
assign n82 = n23 & n2;
assign n63 = ~(n73 | n78);
assign n54 = ~(n3 | n57);
assign n78 = ~n0;
assign n7 = n61 | n57;
assign n30 = ~(n73 | n6);
assign n4 = ~(n49 ^ n56);
assign n27 = n45 | n48;
assign n28 = ~n23;
assign n23 = n47 | n81;
assign n50 = n76 | n30;
assign n14 = n35 | n8;
assign n51 = n16 & n74;
assign n2 = n1 & n83;
assign n45 = ~n35;
assign n33 = n25 & n75;
assign n42 = ~n32;
assign n12 = ~n2;
assign n71 = n32 | n44;
assign n62 = n80 & n3;
assign n18 = n0 | n8;
endmodule
